

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6508, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934;

  CLKBUF_X1 U7256 ( .A(n11242), .Z(n15648) );
  NAND2_X1 U7257 ( .A1(n10176), .A2(n10175), .ZN(n14329) );
  CLKBUF_X2 U7258 ( .A(n9834), .Z(n12571) );
  AND2_X1 U7259 ( .A1(n8464), .A2(n8463), .ZN(n11601) );
  INV_X2 U7260 ( .A(n9953), .ZN(n6513) );
  CLKBUF_X2 U7261 ( .A(n9101), .Z(n9356) );
  NAND2_X1 U7262 ( .A1(n11137), .A2(n9620), .ZN(n9621) );
  AND2_X2 U7263 ( .A1(n14075), .A2(n14176), .ZN(n11791) );
  INV_X2 U7264 ( .A(n9953), .ZN(n10108) );
  INV_X1 U7266 ( .A(n10185), .ZN(n10275) );
  INV_X2 U7267 ( .A(n10643), .ZN(n13968) );
  AND2_X2 U7268 ( .A1(n11209), .A2(n14075), .ZN(n11714) );
  INV_X1 U7269 ( .A(n8763), .ZN(n8750) );
  INV_X1 U7270 ( .A(n15648), .ZN(n6508) );
  INV_X1 U7271 ( .A(n6508), .ZN(P2_U3088) );
  INV_X1 U7272 ( .A(n6508), .ZN(n6510) );
  INV_X1 U7273 ( .A(n13006), .ZN(n13011) );
  INV_X2 U7275 ( .A(n6560), .ZN(n13991) );
  NAND3_X1 U7276 ( .A1(n10189), .A2(n7695), .A3(n7694), .ZN(n10165) );
  AND2_X1 U7277 ( .A1(n11633), .A2(n9085), .ZN(n11537) );
  AND2_X1 U7278 ( .A1(n9778), .A2(n13028), .ZN(n13006) );
  INV_X1 U7279 ( .A(n10091), .ZN(n9996) );
  AND2_X1 U7280 ( .A1(n15427), .A2(n8111), .ZN(n8765) );
  NAND2_X1 U7282 ( .A1(n8186), .A2(SI_22_), .ZN(n8189) );
  AND2_X2 U7283 ( .A1(n8216), .A2(n6594), .ZN(n7475) );
  NAND2_X1 U7285 ( .A1(n11936), .A2(n7911), .ZN(n12054) );
  INV_X2 U7286 ( .A(n15767), .ZN(n14481) );
  INV_X1 U7287 ( .A(n13843), .ZN(n15806) );
  INV_X1 U7288 ( .A(n10111), .ZN(n10123) );
  NAND2_X1 U7289 ( .A1(n12904), .A2(n12910), .ZN(n12879) );
  NAND2_X1 U7290 ( .A1(n7403), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9027) );
  NAND2_X2 U7291 ( .A1(n10235), .A2(n10234), .ZN(n14605) );
  NAND2_X1 U7292 ( .A1(n10799), .A2(n11398), .ZN(n11271) );
  NAND2_X1 U7293 ( .A1(n13706), .A2(n12634), .ZN(n13776) );
  AND2_X1 U7294 ( .A1(n11791), .A2(n14066), .ZN(n15780) );
  INV_X1 U7295 ( .A(n11905), .ZN(n7648) );
  INV_X2 U7296 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n10189) );
  NAND2_X1 U7297 ( .A1(n8333), .A2(n8332), .ZN(n11700) );
  INV_X2 U7298 ( .A(n8088), .ZN(n8768) );
  XNOR2_X1 U7299 ( .A(n10073), .B(n14839), .ZN(n15064) );
  OR2_X1 U7300 ( .A1(n10139), .A2(n8971), .ZN(n15571) );
  NAND3_X1 U7302 ( .A1(n8290), .A2(n8292), .A3(n8041), .ZN(n14855) );
  INV_X2 U7303 ( .A(n15232), .ZN(n15262) );
  INV_X1 U7304 ( .A(n8111), .ZN(n15431) );
  INV_X1 U7305 ( .A(n11839), .ZN(n6959) );
  NAND2_X2 U7306 ( .A1(n8890), .A2(n8889), .ZN(n12000) );
  XNOR2_X1 U7307 ( .A(n10189), .B(n10183), .ZN(n15609) );
  BUF_X2 U7309 ( .A(n9547), .Z(n9548) );
  AOI21_X2 U7310 ( .B1(n9729), .B2(n10922), .A(n9702), .ZN(n9735) );
  INV_X1 U7311 ( .A(n11677), .ZN(n14849) );
  INV_X2 U7312 ( .A(n14104), .ZN(n13816) );
  INV_X1 U7313 ( .A(n8764), .ZN(n8623) );
  NAND2_X2 U7314 ( .A1(n11712), .A2(n7679), .ZN(n11758) );
  NAND2_X1 U7315 ( .A1(n11421), .A2(n11427), .ZN(n11712) );
  NAND3_X2 U7317 ( .A1(n7751), .A2(n8979), .A3(n10868), .ZN(n10724) );
  AOI21_X2 U7318 ( .B1(n13081), .B2(n9629), .A(n9628), .ZN(n9630) );
  INV_X2 U7319 ( .A(n6560), .ZN(n6511) );
  NAND2_X2 U7321 ( .A1(n7039), .A2(n7521), .ZN(n9622) );
  NAND2_X4 U7322 ( .A1(n6981), .A2(n6980), .ZN(n8125) );
  NAND4_X2 U7323 ( .A1(n6983), .A2(n6982), .A3(P2_ADDR_REG_19__SCAN_IN), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n6980) );
  NAND4_X2 U7324 ( .A1(n8117), .A2(n7204), .A3(P3_ADDR_REG_19__SCAN_IN), .A4(
        n6957), .ZN(n6981) );
  NAND2_X2 U7325 ( .A1(n10813), .A2(n10812), .ZN(n11457) );
  OR2_X2 U7326 ( .A1(n9055), .A2(n15852), .ZN(n12903) );
  NAND2_X2 U7327 ( .A1(n8445), .A2(n8444), .ZN(n8965) );
  XNOR2_X2 U7328 ( .A(n14605), .B(n14095), .ZN(n14047) );
  NAND2_X4 U7329 ( .A1(n8010), .A2(n10229), .ZN(n13870) );
  NAND2_X2 U7330 ( .A1(n7130), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9046) );
  NAND2_X2 U7331 ( .A1(n8641), .A2(n8640), .ZN(n10073) );
  OR2_X2 U7332 ( .A1(n12656), .A2(n8075), .ZN(n6575) );
  AOI211_X1 U7333 ( .C1(n10816), .C2(n10815), .A(n13796), .B(n10814), .ZN(
        n10829) );
  BUF_X4 U7334 ( .A(n8765), .Z(n6514) );
  AOI211_X1 U7335 ( .C1(n14505), .C2(n14187), .A(n14481), .B(n14186), .ZN(
        n14504) );
  NAND2_X1 U7336 ( .A1(n14308), .A2(n6612), .ZN(n14301) );
  NAND2_X1 U7337 ( .A1(n10294), .A2(n10293), .ZN(n14217) );
  NAND2_X1 U7338 ( .A1(n7672), .A2(n7671), .ZN(n13707) );
  NAND2_X1 U7339 ( .A1(n12608), .A2(n12607), .ZN(n13634) );
  NAND2_X1 U7340 ( .A1(n8934), .A2(n8939), .ZN(n15210) );
  NAND2_X1 U7341 ( .A1(n8614), .A2(n8613), .ZN(n15319) );
  NAND2_X1 U7342 ( .A1(n10258), .A2(n10257), .ZN(n14580) );
  XNOR2_X1 U7343 ( .A(n8566), .B(n8565), .ZN(n11779) );
  AND3_X1 U7344 ( .A1(n11571), .A2(n7855), .A3(n7853), .ZN(n11920) );
  NAND2_X1 U7345 ( .A1(n11368), .A2(n11370), .ZN(n11369) );
  XNOR2_X1 U7346 ( .A(n8347), .B(n8346), .ZN(n10911) );
  NAND2_X2 U7347 ( .A1(n7156), .A2(n12900), .ZN(n11660) );
  INV_X1 U7348 ( .A(n13039), .ZN(n11772) );
  INV_X1 U7349 ( .A(n13041), .ZN(n7251) );
  INV_X2 U7350 ( .A(n13813), .ZN(n15800) );
  BUF_X2 U7351 ( .A(n11714), .Z(n15767) );
  INV_X4 U7352 ( .A(n8261), .ZN(n8779) );
  NAND4_X1 U7353 ( .A1(n8270), .A2(n8269), .A3(n8268), .A4(n8267), .ZN(n14854)
         );
  BUF_X1 U7354 ( .A(n7880), .Z(n6522) );
  CLKBUF_X2 U7355 ( .A(n9041), .Z(n9346) );
  NOR2_X1 U7356 ( .A1(n9058), .A2(n11777), .ZN(n9112) );
  INV_X4 U7357 ( .A(n12858), .ZN(n9466) );
  NOR2_X1 U7358 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n7327) );
  NAND2_X1 U7359 ( .A1(n7287), .A2(n14027), .ZN(n14079) );
  OAI21_X1 U7360 ( .B1(n6763), .B2(n6762), .A(n7698), .ZN(n7227) );
  AOI21_X1 U7361 ( .B1(n14213), .B2(n15770), .A(n14212), .ZN(n7308) );
  NAND2_X1 U7362 ( .A1(n7219), .A2(n7220), .ZN(n13783) );
  AND2_X1 U7363 ( .A1(n12564), .A2(n14490), .ZN(n10360) );
  AND2_X1 U7364 ( .A1(n8038), .A2(n8037), .ZN(n15287) );
  NOR2_X1 U7365 ( .A1(n14504), .A2(n7261), .ZN(n14506) );
  OAI21_X1 U7366 ( .B1(n14763), .B2(n7004), .A(n7739), .ZN(n14811) );
  OR3_X1 U7367 ( .A1(n15305), .A2(n15304), .A3(n15303), .ZN(n15406) );
  OAI21_X1 U7368 ( .B1(n14224), .B2(n6524), .A(n14058), .ZN(n7341) );
  AND2_X1 U7369 ( .A1(n14223), .A2(n14222), .ZN(n14224) );
  NOR2_X1 U7370 ( .A1(n13747), .A2(n12657), .ZN(n7266) );
  OAI21_X1 U7371 ( .B1(n14301), .B2(n14032), .A(n14031), .ZN(n14281) );
  XNOR2_X1 U7372 ( .A(n12653), .B(n12652), .ZN(n13747) );
  NAND2_X1 U7373 ( .A1(n7687), .A2(n12639), .ZN(n13725) );
  NAND2_X1 U7374 ( .A1(n13231), .A2(n8073), .ZN(n13216) );
  OR2_X1 U7375 ( .A1(n13776), .A2(n13775), .ZN(n7687) );
  NAND2_X1 U7376 ( .A1(n7760), .A2(n7759), .ZN(n14772) );
  NAND2_X1 U7377 ( .A1(n6916), .A2(n6915), .ZN(n14243) );
  AND2_X1 U7378 ( .A1(n10675), .A2(n13193), .ZN(n12867) );
  AND2_X1 U7379 ( .A1(n14283), .A2(n6564), .ZN(n14231) );
  XNOR2_X1 U7380 ( .A(n14217), .B(n14088), .ZN(n14222) );
  NAND2_X1 U7381 ( .A1(n12854), .A2(n12853), .ZN(n13183) );
  XNOR2_X1 U7382 ( .A(n8739), .B(n8738), .ZN(n12558) );
  CLKBUF_X1 U7383 ( .A(n9632), .Z(n9633) );
  NAND2_X1 U7384 ( .A1(n8681), .A2(n8680), .ZN(n15289) );
  NAND2_X1 U7385 ( .A1(n10299), .A2(n10298), .ZN(n14184) );
  OR2_X1 U7386 ( .A1(n10623), .A2(n14244), .ZN(n10628) );
  NAND2_X1 U7387 ( .A1(n6963), .A2(n6961), .ZN(n15149) );
  AOI22_X1 U7388 ( .A1(n12844), .A2(n7262), .B1(SI_30_), .B2(n12863), .ZN(
        n13507) );
  NAND2_X1 U7389 ( .A1(n8678), .A2(n8677), .ZN(n15437) );
  NAND2_X1 U7390 ( .A1(n8671), .A2(n8670), .ZN(n15030) );
  AND2_X1 U7391 ( .A1(n10506), .A2(n14051), .ZN(n7313) );
  XNOR2_X1 U7392 ( .A(n8639), .B(n8638), .ZN(n12036) );
  NAND2_X1 U7393 ( .A1(n6765), .A2(n6609), .ZN(n14390) );
  OAI21_X1 U7394 ( .B1(n12552), .B2(n12551), .A(n12550), .ZN(n12706) );
  NAND2_X1 U7395 ( .A1(n7151), .A2(n9289), .ZN(n13357) );
  NAND2_X1 U7396 ( .A1(n8649), .A2(n8648), .ZN(n12162) );
  NAND2_X1 U7397 ( .A1(n8248), .A2(n15441), .ZN(n15090) );
  NAND2_X1 U7398 ( .A1(n7843), .A2(n7847), .ZN(n15235) );
  NAND2_X1 U7399 ( .A1(n8933), .A2(n8484), .ZN(n8897) );
  AND2_X1 U7400 ( .A1(n8967), .A2(n7844), .ZN(n7843) );
  AOI21_X1 U7401 ( .B1(n9526), .B2(n12989), .A(n7872), .ZN(n7871) );
  OR2_X1 U7402 ( .A1(n8647), .A2(n8646), .ZN(n8648) );
  NAND2_X1 U7403 ( .A1(n8647), .A2(n8646), .ZN(n8649) );
  XNOR2_X1 U7404 ( .A(n8627), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15441) );
  NAND2_X1 U7405 ( .A1(n7514), .A2(n7513), .ZN(n13075) );
  NAND2_X1 U7406 ( .A1(n10262), .A2(n10261), .ZN(n14393) );
  NAND2_X2 U7407 ( .A1(n8511), .A2(n8510), .ZN(n15339) );
  NAND2_X1 U7408 ( .A1(n10277), .A2(n10276), .ZN(n14351) );
  NAND2_X1 U7409 ( .A1(n10279), .A2(n10278), .ZN(n14544) );
  OR2_X1 U7410 ( .A1(n8965), .A2(n15213), .ZN(n8933) );
  NAND2_X1 U7411 ( .A1(n8187), .A2(n8189), .ZN(n10283) );
  OAI22_X1 U7412 ( .A1(n6605), .A2(n6785), .B1(n13872), .B2(n13871), .ZN(
        n13875) );
  NAND2_X1 U7413 ( .A1(n6845), .A2(n8563), .ZN(n8566) );
  NAND2_X1 U7414 ( .A1(n7226), .A2(n10265), .ZN(n14568) );
  NAND2_X1 U7415 ( .A1(n12108), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n12107) );
  NAND2_X1 U7416 ( .A1(n9425), .A2(n9413), .ZN(n9426) );
  XNOR2_X1 U7417 ( .A(n8469), .B(n8468), .ZN(n11319) );
  AND2_X1 U7418 ( .A1(n7678), .A2(n12585), .ZN(n7677) );
  AND2_X1 U7419 ( .A1(n10445), .A2(n12069), .ZN(n12026) );
  AND2_X1 U7420 ( .A1(n6769), .A2(n6768), .ZN(n13862) );
  NAND2_X1 U7421 ( .A1(n7821), .A2(n7819), .ZN(n8591) );
  NAND2_X1 U7422 ( .A1(n8401), .A2(n8400), .ZN(n15391) );
  AOI21_X1 U7423 ( .B1(n9375), .B2(n6697), .A(n7805), .ZN(n9411) );
  OAI21_X1 U7424 ( .B1(n8519), .B2(n8518), .A(n8517), .ZN(n8521) );
  NAND2_X1 U7425 ( .A1(n9322), .A2(n9321), .ZN(n13538) );
  NOR2_X1 U7426 ( .A1(n9594), .A2(n9662), .ZN(n9595) );
  NAND2_X1 U7427 ( .A1(n12017), .A2(n14038), .ZN(n12016) );
  NAND2_X1 U7428 ( .A1(n11457), .A2(n7309), .ZN(n11456) );
  NOR2_X1 U7429 ( .A1(n11549), .A2(n7354), .ZN(n9594) );
  XNOR2_X1 U7430 ( .A(n8395), .B(n8394), .ZN(n10949) );
  OAI22_X1 U7431 ( .A1(n13851), .A2(n6767), .B1(n13852), .B2(n6766), .ZN(n6772) );
  NAND2_X1 U7432 ( .A1(n8393), .A2(n8392), .ZN(n8395) );
  NAND2_X1 U7433 ( .A1(n8461), .A2(n8085), .ZN(n7818) );
  NAND2_X1 U7434 ( .A1(n7510), .A2(n7509), .ZN(n7032) );
  XNOR2_X1 U7435 ( .A(n8391), .B(n8389), .ZN(n10222) );
  XNOR2_X1 U7436 ( .A(n9370), .B(n12359), .ZN(n9369) );
  NAND2_X1 U7437 ( .A1(n8158), .A2(n8157), .ZN(n8461) );
  OAI21_X1 U7438 ( .B1(n13846), .B2(n7697), .A(n7696), .ZN(n13851) );
  NAND2_X1 U7439 ( .A1(n11295), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n11547) );
  XNOR2_X1 U7440 ( .A(n15764), .B(n13855), .ZN(n15765) );
  NAND2_X1 U7441 ( .A1(n8375), .A2(n8374), .ZN(n8391) );
  NOR2_X1 U7442 ( .A1(n9593), .A2(n6736), .ZN(n11295) );
  OAI21_X1 U7443 ( .B1(n9302), .B2(n7791), .A(n7788), .ZN(n9332) );
  NAND2_X1 U7444 ( .A1(n6979), .A2(n8220), .ZN(n11500) );
  XNOR2_X1 U7445 ( .A(n12924), .B(n9834), .ZN(n11955) );
  INV_X1 U7446 ( .A(n8881), .ZN(n6515) );
  CLKBUF_X1 U7448 ( .A(n9886), .Z(n10098) );
  CLKBUF_X1 U7449 ( .A(n10798), .Z(n14479) );
  NAND4_X1 U7450 ( .A1(n10395), .A2(n10394), .A3(n10393), .A4(n10392), .ZN(
        n14101) );
  OAI211_X1 U7451 ( .C1(n7381), .C2(SI_4_), .A(n7095), .B(n7094), .ZN(n15885)
         );
  INV_X8 U7452 ( .A(n6520), .ZN(n14022) );
  AND3_X1 U7453 ( .A1(n9126), .A2(n9125), .A3(n9124), .ZN(n15896) );
  INV_X2 U7454 ( .A(n7381), .ZN(n12863) );
  NAND2_X1 U7455 ( .A1(n11151), .A2(n11152), .ZN(n7120) );
  NAND2_X2 U7456 ( .A1(n6632), .A2(n9045), .ZN(n9055) );
  INV_X1 U7457 ( .A(n8299), .ZN(n6516) );
  INV_X2 U7458 ( .A(n9064), .ZN(n7262) );
  AND4_X2 U7459 ( .A1(n8233), .A2(n8232), .A3(n8231), .A4(n8230), .ZN(n11489)
         );
  NAND4_X1 U7460 ( .A1(n9034), .A2(n9033), .A3(n9032), .A4(n9031), .ZN(n13042)
         );
  NAND2_X1 U7461 ( .A1(n8960), .A2(n8959), .ZN(n15545) );
  NAND2_X1 U7462 ( .A1(n13812), .A2(n11791), .ZN(n13811) );
  OR2_X1 U7463 ( .A1(n15571), .A2(n15199), .ZN(n15138) );
  NAND4_X1 U7464 ( .A1(n8245), .A2(n8244), .A3(n8243), .A4(n8242), .ZN(n14856)
         );
  CLKBUF_X3 U7465 ( .A(n9089), .Z(n12847) );
  INV_X1 U7466 ( .A(n10643), .ZN(n6521) );
  XNOR2_X1 U7467 ( .A(n9338), .B(n9486), .ZN(n13170) );
  INV_X1 U7468 ( .A(n10315), .ZN(n13812) );
  AOI21_X1 U7469 ( .B1(n7730), .B2(n9727), .A(n9699), .ZN(n9701) );
  CLKBUF_X1 U7470 ( .A(n10350), .Z(n14076) );
  INV_X1 U7471 ( .A(n8970), .ZN(n8958) );
  NAND2_X1 U7472 ( .A1(n9019), .A2(n9021), .ZN(n12858) );
  NAND2_X4 U7473 ( .A1(n14669), .A2(n10314), .ZN(n10184) );
  XNOR2_X1 U7474 ( .A(n8213), .B(n8212), .ZN(n8969) );
  CLKBUF_X1 U7475 ( .A(n8821), .Z(n14874) );
  NAND2_X1 U7476 ( .A1(n11138), .A2(n11139), .ZN(n11137) );
  AND2_X2 U7477 ( .A1(n8110), .A2(n15431), .ZN(n8764) );
  XNOR2_X1 U7478 ( .A(n7166), .B(P3_IR_REG_30__SCAN_IN), .ZN(n9021) );
  XNOR2_X1 U7479 ( .A(n8208), .B(P1_IR_REG_20__SCAN_IN), .ZN(n8971) );
  AND2_X1 U7480 ( .A1(n7398), .A2(n7396), .ZN(n7395) );
  XNOR2_X1 U7481 ( .A(n10319), .B(n14657), .ZN(n12560) );
  OR2_X1 U7482 ( .A1(n9016), .A2(n9015), .ZN(n9018) );
  NAND2_X1 U7483 ( .A1(n10344), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6758) );
  NAND2_X1 U7484 ( .A1(n14660), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10319) );
  NAND2_X1 U7485 ( .A1(n10310), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10312) );
  OAI21_X1 U7486 ( .B1(n8816), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8207) );
  AND2_X1 U7487 ( .A1(n9258), .A2(n12489), .ZN(n9260) );
  XNOR2_X1 U7488 ( .A(n7446), .B(n8209), .ZN(n15163) );
  AND2_X1 U7489 ( .A1(n10173), .A2(n7726), .ZN(n10305) );
  NAND2_X1 U7490 ( .A1(n7117), .A2(n7116), .ZN(n14660) );
  XNOR2_X1 U7491 ( .A(n7659), .B(P1_IR_REG_29__SCAN_IN), .ZN(n8111) );
  NAND2_X2 U7492 ( .A1(n10879), .A2(n6510), .ZN(n14671) );
  AND2_X1 U7493 ( .A1(n6680), .A2(n7118), .ZN(n7117) );
  NAND2_X2 U7494 ( .A1(n10879), .A2(P1_U3086), .ZN(n15438) );
  INV_X1 U7495 ( .A(n10833), .ZN(n11124) );
  XNOR2_X1 U7496 ( .A(n8126), .B(SI_2_), .ZN(n8280) );
  NAND2_X1 U7497 ( .A1(n7393), .A2(n6734), .ZN(n9102) );
  INV_X1 U7498 ( .A(n8474), .ZN(n6517) );
  AND2_X1 U7499 ( .A1(n7119), .A2(n10166), .ZN(n7115) );
  NOR2_X1 U7500 ( .A1(n9014), .A2(n7921), .ZN(n7918) );
  NOR2_X1 U7501 ( .A1(n10163), .A2(n10333), .ZN(n10167) );
  NAND4_X1 U7502 ( .A1(n7475), .A2(n6581), .A3(n8103), .A4(n7474), .ZN(n8109)
         );
  NAND2_X1 U7503 ( .A1(n10171), .A2(n10159), .ZN(n10163) );
  CLKBUF_X1 U7504 ( .A(n10171), .Z(n10172) );
  NAND2_X1 U7505 ( .A1(n9218), .A2(n9013), .ZN(n9014) );
  AND2_X1 U7506 ( .A1(n7150), .A2(n7149), .ZN(n8080) );
  NAND2_X1 U7507 ( .A1(n7129), .A2(n7128), .ZN(n7130) );
  AND3_X1 U7508 ( .A1(n7670), .A2(n7669), .A3(n7668), .ZN(n10224) );
  AND2_X1 U7509 ( .A1(n7320), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n9721) );
  NAND4_X1 U7510 ( .A1(n10162), .A2(n10161), .A3(n7327), .A4(n10160), .ZN(
        n10333) );
  AND3_X1 U7511 ( .A1(n6903), .A2(n6902), .A3(n6901), .ZN(n10171) );
  NOR2_X1 U7512 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n9012) );
  NOR2_X1 U7513 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n9011) );
  NOR2_X1 U7514 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n6901) );
  INV_X1 U7515 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n10160) );
  NOR2_X1 U7516 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n9010) );
  NOR2_X1 U7517 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n6902) );
  INV_X1 U7518 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n6983) );
  NOR2_X1 U7519 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6903) );
  NOR3_X1 U7520 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), .A3(
        P3_IR_REG_5__SCAN_IN), .ZN(n9013) );
  INV_X1 U7521 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n9335) );
  INV_X1 U7522 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n10177) );
  NOR2_X1 U7523 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n10161) );
  NOR2_X1 U7524 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n10162) );
  INV_X1 U7525 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n10318) );
  INV_X1 U7526 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7129) );
  INV_X1 U7527 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7128) );
  INV_X1 U7528 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8440) );
  INV_X1 U7529 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7652) );
  INV_X4 U7530 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U7531 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n7670) );
  NOR2_X1 U7532 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n7669) );
  NOR2_X1 U7533 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n7668) );
  INV_X1 U7534 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n12301) );
  INV_X1 U7535 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8210) );
  INV_X1 U7536 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9541) );
  INV_X1 U7537 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9544) );
  NOR2_X1 U7538 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n7150) );
  INV_X1 U7539 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7204) );
  INV_X1 U7540 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8117) );
  INV_X4 U7541 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7542 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8329) );
  NOR2_X1 U7543 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), .ZN(
        n9006) );
  NOR2_X1 U7544 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), .ZN(
        n9007) );
  INV_X1 U7545 ( .A(n8125), .ZN(n8132) );
  OR2_X2 U7546 ( .A1(n9634), .A2(n13101), .ZN(n6623) );
  INV_X1 U7547 ( .A(n12858), .ZN(n6518) );
  OAI21_X1 U7548 ( .B1(n13075), .B2(n13480), .A(n7511), .ZN(n13081) );
  INV_X1 U7549 ( .A(n11714), .ZN(n14311) );
  XNOR2_X2 U7550 ( .A(n9625), .B(n10903), .ZN(n12108) );
  OAI21_X2 U7551 ( .B1(n13390), .B2(n9288), .A(n9287), .ZN(n7151) );
  XNOR2_X2 U7552 ( .A(n9764), .B(P3_ADDR_REG_17__SCAN_IN), .ZN(n15468) );
  XNOR2_X2 U7553 ( .A(n9763), .B(P1_ADDR_REG_17__SCAN_IN), .ZN(n9764) );
  AOI21_X2 U7554 ( .B1(n11885), .B2(n11886), .A(n7508), .ZN(n9625) );
  AOI22_X2 U7555 ( .A1(n11196), .A2(P3_REG1_REG_5__SCAN_IN), .B1(n11202), .B2(
        n9623), .ZN(n11176) );
  NAND2_X1 U7556 ( .A1(n10184), .A2(n10879), .ZN(n6519) );
  OAI211_X1 U7557 ( .C1(n11145), .C2(n9605), .A(n9054), .B(n9053), .ZN(n15852)
         );
  BUF_X4 U7558 ( .A(n6561), .Z(n6520) );
  NAND2_X1 U7559 ( .A1(n15780), .A2(n13812), .ZN(n6561) );
  NOR2_X4 U7560 ( .A1(n10651), .A2(n13992), .ZN(n10722) );
  XNOR2_X2 U7561 ( .A(n6756), .B(n10318), .ZN(n10314) );
  NAND2_X1 U7562 ( .A1(n10572), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n10639) );
  INV_X1 U7563 ( .A(n10573), .ZN(n10572) );
  AND2_X1 U7564 ( .A1(n10647), .A2(n10646), .ZN(n14196) );
  NAND2_X1 U7565 ( .A1(n13894), .A2(n7724), .ZN(n7723) );
  AND2_X1 U7566 ( .A1(n13926), .A2(n7704), .ZN(n7703) );
  OR2_X1 U7567 ( .A1(n13928), .A2(n13927), .ZN(n7704) );
  NOR2_X1 U7568 ( .A1(n13929), .A2(n7239), .ZN(n13926) );
  AND2_X1 U7569 ( .A1(n13930), .A2(n13931), .ZN(n7239) );
  NOR2_X2 U7570 ( .A1(n13811), .A2(n14077), .ZN(n6560) );
  OR2_X1 U7571 ( .A1(n9806), .A2(n7963), .ZN(n7962) );
  INV_X1 U7572 ( .A(n7946), .ZN(n7939) );
  INV_X1 U7573 ( .A(n9019), .ZN(n9020) );
  NAND2_X1 U7574 ( .A1(n7120), .A2(n6604), .ZN(n7625) );
  OR2_X1 U7575 ( .A1(n13438), .A2(n12756), .ZN(n13012) );
  OR2_X1 U7576 ( .A1(n13037), .A2(n6956), .ZN(n12928) );
  CLKBUF_X1 U7577 ( .A(n9775), .Z(n11101) );
  OR2_X1 U7578 ( .A1(n13526), .A2(n12745), .ZN(n12992) );
  OR2_X1 U7579 ( .A1(n9557), .A2(n9569), .ZN(n10684) );
  AND2_X1 U7580 ( .A1(n7777), .A2(n9201), .ZN(n7776) );
  NAND2_X1 U7581 ( .A1(n7778), .A2(n9189), .ZN(n7777) );
  INV_X1 U7582 ( .A(n9187), .ZN(n7778) );
  NAND2_X1 U7583 ( .A1(n7472), .A2(n6600), .ZN(n8202) );
  AND2_X1 U7584 ( .A1(n8103), .A2(n8205), .ZN(n7472) );
  AND2_X1 U7585 ( .A1(n8106), .A2(n7279), .ZN(n7473) );
  OR2_X1 U7586 ( .A1(n8591), .A2(n11698), .ZN(n8607) );
  INV_X1 U7587 ( .A(n9058), .ZN(n9497) );
  NAND2_X1 U7588 ( .A1(n12557), .A2(n9019), .ZN(n9089) );
  OR2_X1 U7589 ( .A1(n13240), .A2(n13249), .ZN(n8073) );
  OR2_X1 U7591 ( .A1(n9778), .A2(n13028), .ZN(n15901) );
  NAND2_X1 U7592 ( .A1(n13603), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7166) );
  OR2_X1 U7593 ( .A1(n14219), .A2(n7879), .ZN(n10579) );
  NAND2_X1 U7594 ( .A1(n14191), .A2(n10710), .ZN(n14496) );
  NAND2_X1 U7595 ( .A1(n6918), .A2(n6917), .ZN(n10714) );
  AND2_X1 U7596 ( .A1(n6674), .A2(n10634), .ZN(n6917) );
  AOI21_X1 U7597 ( .B1(n7984), .B2(n7982), .A(n14244), .ZN(n7980) );
  NAND2_X1 U7598 ( .A1(n14032), .A2(n14031), .ZN(n7105) );
  AOI21_X1 U7599 ( .B1(n6528), .B2(n10619), .A(n6640), .ZN(n7914) );
  NAND2_X1 U7600 ( .A1(n10454), .A2(n12025), .ZN(n8008) );
  NAND2_X1 U7601 ( .A1(n11238), .A2(n10648), .ZN(n14472) );
  NAND2_X1 U7602 ( .A1(n10296), .A2(n10295), .ZN(n13992) );
  INV_X1 U7603 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7695) );
  INV_X1 U7604 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n7694) );
  AND4_X1 U7605 ( .A1(n7203), .A2(n7202), .A3(n7201), .A4(n7200), .ZN(n8103)
         );
  NOR2_X1 U7606 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n7203) );
  NOR2_X1 U7607 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n7202) );
  NOR2_X1 U7608 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n7200) );
  NAND2_X1 U7609 ( .A1(n7199), .A2(n6593), .ZN(n7388) );
  NOR2_X1 U7610 ( .A1(n7198), .A2(n6590), .ZN(n7197) );
  OAI22_X1 U7611 ( .A1(n9757), .A2(n9756), .B1(P1_ADDR_REG_15__SCAN_IN), .B2(
        n13104), .ZN(n9762) );
  NAND2_X1 U7612 ( .A1(n13818), .A2(n13817), .ZN(n13824) );
  OR2_X1 U7613 ( .A1(n13816), .A2(n6520), .ZN(n13818) );
  MUX2_X1 U7614 ( .A(n9892), .B(n14709), .S(n8261), .Z(n8264) );
  INV_X1 U7615 ( .A(n7633), .ZN(n8250) );
  OR2_X1 U7616 ( .A1(n8309), .A2(n11500), .ZN(n7171) );
  OAI21_X1 U7617 ( .B1(n8780), .B2(n14852), .A(n11500), .ZN(n7170) );
  NAND2_X1 U7618 ( .A1(n7587), .A2(n6569), .ZN(n7585) );
  NAND2_X1 U7619 ( .A1(n8402), .A2(n7459), .ZN(n7458) );
  NAND2_X1 U7620 ( .A1(n8383), .A2(n7173), .ZN(n8404) );
  OAI21_X1 U7621 ( .B1(n8382), .B2(n8381), .A(n8380), .ZN(n7173) );
  AND2_X1 U7622 ( .A1(n12955), .A2(n7078), .ZN(n7077) );
  NAND2_X1 U7623 ( .A1(n7079), .A2(n7081), .ZN(n7078) );
  INV_X1 U7624 ( .A(n7084), .ZN(n7081) );
  AND2_X1 U7625 ( .A1(n8545), .A2(n8068), .ZN(n8546) );
  NAND2_X1 U7626 ( .A1(n13307), .A2(n12982), .ZN(n7091) );
  NOR2_X1 U7627 ( .A1(n12990), .A2(n13273), .ZN(n7092) );
  MUX2_X1 U7628 ( .A(n15098), .B(n15127), .S(n8261), .Z(n8596) );
  NAND2_X1 U7629 ( .A1(n13948), .A2(n13918), .ZN(n13951) );
  AND2_X1 U7630 ( .A1(n7723), .A2(n13889), .ZN(n7722) );
  OR4_X1 U7631 ( .A1(n11673), .A2(n11581), .A3(n8831), .A4(n11568), .ZN(n8832)
         );
  NAND2_X1 U7632 ( .A1(n6969), .A2(n6968), .ZN(n10629) );
  NAND2_X1 U7633 ( .A1(n10649), .A2(n14217), .ZN(n6968) );
  INV_X1 U7634 ( .A(n10625), .ZN(n6969) );
  NAND3_X1 U7635 ( .A1(n7180), .A2(n6654), .A3(n7177), .ZN(n7464) );
  AOI21_X1 U7636 ( .B1(n7961), .B2(n7963), .A(n9813), .ZN(n7960) );
  NAND2_X1 U7637 ( .A1(n11124), .A2(n15910), .ZN(n7526) );
  OR2_X1 U7638 ( .A1(n10833), .A2(n11124), .ZN(n7529) );
  AND2_X1 U7639 ( .A1(n10872), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7508) );
  NAND2_X1 U7640 ( .A1(n7629), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7138) );
  AND2_X1 U7641 ( .A1(n6699), .A2(n9281), .ZN(n7041) );
  INV_X1 U7642 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n9281) );
  AND2_X1 U7643 ( .A1(n6677), .A2(n7161), .ZN(n7160) );
  NAND2_X1 U7644 ( .A1(n7162), .A2(n9184), .ZN(n7161) );
  INV_X1 U7645 ( .A(n7164), .ZN(n7162) );
  INV_X1 U7646 ( .A(n9511), .ZN(n7894) );
  NAND2_X1 U7647 ( .A1(n15896), .A2(n13038), .ZN(n12923) );
  AND2_X1 U7648 ( .A1(n13511), .A2(n12868), .ZN(n12873) );
  NOR2_X1 U7649 ( .A1(n9368), .A2(n13307), .ZN(n13281) );
  AND2_X1 U7650 ( .A1(n12843), .A2(n13382), .ZN(n12961) );
  OR2_X1 U7651 ( .A1(n12148), .A2(n11950), .ZN(n9184) );
  AND2_X1 U7652 ( .A1(n9605), .A2(n9609), .ZN(n9505) );
  NAND2_X1 U7653 ( .A1(n8080), .A2(n7922), .ZN(n7921) );
  INV_X1 U7654 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7922) );
  INV_X1 U7655 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9575) );
  AND2_X1 U7656 ( .A1(n7972), .A2(n7971), .ZN(n7970) );
  NAND2_X1 U7657 ( .A1(n9334), .A2(n9320), .ZN(n9370) );
  INV_X1 U7658 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n12489) );
  NOR2_X1 U7659 ( .A1(n9137), .A2(n7786), .ZN(n7785) );
  INV_X1 U7660 ( .A(n9119), .ZN(n7786) );
  NAND2_X1 U7661 ( .A1(n10883), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n9136) );
  INV_X1 U7662 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9098) );
  XNOR2_X1 U7663 ( .A(n14580), .B(n11713), .ZN(n12613) );
  AND2_X1 U7664 ( .A1(n13928), .A2(n13927), .ZN(n7705) );
  INV_X1 U7665 ( .A(n12560), .ZN(n6907) );
  NAND2_X1 U7666 ( .A1(n6779), .A2(n6778), .ZN(n10651) );
  AND2_X1 U7667 ( .A1(n6780), .A2(n14626), .ZN(n6779) );
  INV_X1 U7668 ( .A(n14294), .ZN(n6778) );
  AND2_X1 U7669 ( .A1(n6564), .A2(n14619), .ZN(n6780) );
  XNOR2_X1 U7670 ( .A(n13870), .B(n8009), .ZN(n10597) );
  NOR2_X1 U7671 ( .A1(n7205), .A2(n13870), .ZN(n7656) );
  INV_X1 U7672 ( .A(n7905), .ZN(n7904) );
  OAI21_X1 U7673 ( .B1(n7908), .B2(n6562), .A(n7910), .ZN(n7905) );
  NAND2_X1 U7674 ( .A1(n7911), .A2(n14097), .ZN(n7910) );
  INV_X1 U7675 ( .A(n10810), .ZN(n11238) );
  NAND2_X1 U7676 ( .A1(n14656), .A2(n10301), .ZN(n10302) );
  AND2_X1 U7677 ( .A1(n7727), .A2(n10311), .ZN(n7726) );
  NAND2_X1 U7678 ( .A1(n7025), .A2(n6701), .ZN(n7026) );
  NAND2_X1 U7679 ( .A1(n7764), .A2(n11865), .ZN(n7017) );
  NAND2_X1 U7680 ( .A1(n7300), .A2(n7299), .ZN(n7139) );
  NAND2_X1 U7681 ( .A1(n10006), .A2(n14682), .ZN(n7299) );
  NAND2_X1 U7682 ( .A1(n10008), .A2(n10007), .ZN(n7300) );
  NAND2_X1 U7683 ( .A1(n7667), .A2(n8659), .ZN(n7666) );
  AND2_X1 U7684 ( .A1(n8057), .A2(n10653), .ZN(n8051) );
  NAND2_X1 U7685 ( .A1(n15289), .A2(n8956), .ZN(n8060) );
  NAND2_X1 U7686 ( .A1(n6651), .A2(n8943), .ZN(n6850) );
  NOR2_X1 U7687 ( .A1(n15108), .A2(n7544), .ZN(n7543) );
  INV_X1 U7688 ( .A(n8907), .ZN(n7544) );
  AOI22_X1 U7689 ( .A1(n15210), .A2(n8899), .B1(n15228), .B2(n15218), .ZN(
        n8900) );
  INV_X1 U7690 ( .A(n8888), .ZN(n8026) );
  NOR2_X1 U7691 ( .A1(n11839), .A2(n7487), .ZN(n7486) );
  OR2_X1 U7692 ( .A1(n15581), .A2(n11832), .ZN(n8926) );
  AOI21_X1 U7693 ( .B1(n8034), .B2(n8905), .A(n6652), .ZN(n8033) );
  AND2_X1 U7694 ( .A1(n8827), .A2(n8924), .ZN(n8061) );
  INV_X1 U7695 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8211) );
  OAI21_X1 U7696 ( .B1(n8649), .B2(n7830), .A(n7827), .ZN(n8702) );
  INV_X1 U7697 ( .A(n7833), .ZN(n7830) );
  AOI21_X1 U7698 ( .B1(n7829), .B2(n7833), .A(n7828), .ZN(n7827) );
  INV_X1 U7699 ( .A(n8197), .ZN(n7828) );
  NAND2_X1 U7700 ( .A1(n7818), .A2(n8162), .ZN(n8519) );
  AOI21_X1 U7701 ( .B1(n7013), .B2(n6855), .A(n6854), .ZN(n6856) );
  INV_X1 U7702 ( .A(n8153), .ZN(n6854) );
  INV_X1 U7703 ( .A(n6574), .ZN(n6855) );
  XNOR2_X1 U7704 ( .A(n9701), .B(P3_ADDR_REG_5__SCAN_IN), .ZN(n9729) );
  AOI21_X1 U7705 ( .B1(n7562), .B2(n7561), .A(n9710), .ZN(n9748) );
  INV_X1 U7706 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n7561) );
  INV_X1 U7707 ( .A(n9745), .ZN(n7562) );
  CLKBUF_X1 U7708 ( .A(n9047), .Z(n9605) );
  INV_X1 U7709 ( .A(n13358), .ZN(n12810) );
  NOR2_X1 U7710 ( .A1(n7059), .A2(n13273), .ZN(n12887) );
  NAND2_X1 U7711 ( .A1(n7067), .A2(n7060), .ZN(n7059) );
  NAND2_X1 U7712 ( .A1(n11115), .A2(n9589), .ZN(n11151) );
  INV_X1 U7713 ( .A(n7615), .ZN(n9589) );
  AND2_X1 U7714 ( .A1(n9592), .A2(n9591), .ZN(n11152) );
  NAND2_X1 U7715 ( .A1(n7029), .A2(n7028), .ZN(n11150) );
  NAND2_X1 U7716 ( .A1(n11158), .A2(n9073), .ZN(n7028) );
  OR2_X1 U7717 ( .A1(n11158), .A2(n9073), .ZN(n7029) );
  INV_X1 U7718 ( .A(n11180), .ZN(n7355) );
  OAI21_X1 U7719 ( .B1(n7125), .B2(n7124), .A(n7123), .ZN(n9597) );
  INV_X1 U7720 ( .A(n13045), .ZN(n7124) );
  AOI21_X1 U7721 ( .B1(n13047), .B2(n13045), .A(n6708), .ZN(n7123) );
  NAND2_X1 U7722 ( .A1(n7135), .A2(n13111), .ZN(n7134) );
  XNOR2_X1 U7723 ( .A(n9632), .B(n11066), .ZN(n13153) );
  OAI21_X1 U7724 ( .B1(n13223), .B2(n9530), .A(n13005), .ZN(n10675) );
  OR2_X1 U7725 ( .A1(n9447), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9464) );
  NAND2_X1 U7726 ( .A1(n13244), .A2(n9424), .ZN(n13233) );
  NAND2_X1 U7727 ( .A1(n9341), .A2(n12303), .ZN(n9343) );
  NOR2_X1 U7728 ( .A1(n9323), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9359) );
  NAND2_X1 U7729 ( .A1(n7864), .A2(n7863), .ZN(n12147) );
  AOI21_X1 U7730 ( .B1(n7866), .B2(n7868), .A(n12939), .ZN(n7863) );
  INV_X1 U7731 ( .A(n7867), .ZN(n7866) );
  NAND2_X1 U7732 ( .A1(n11847), .A2(n7606), .ZN(n12090) );
  NOR2_X1 U7733 ( .A1(n12930), .A2(n7607), .ZN(n7606) );
  INV_X1 U7734 ( .A(n9146), .ZN(n7607) );
  NAND2_X1 U7735 ( .A1(n11631), .A2(n12881), .ZN(n6822) );
  AOI21_X1 U7736 ( .B1(n12700), .B2(n9497), .A(n9484), .ZN(n13201) );
  NAND2_X1 U7737 ( .A1(n12866), .A2(n13013), .ZN(n13194) );
  INV_X1 U7738 ( .A(n13422), .ZN(n15861) );
  OR2_X1 U7739 ( .A1(n13568), .A2(n13382), .ZN(n9289) );
  AND2_X1 U7740 ( .A1(n13006), .A2(n9505), .ZN(n13422) );
  INV_X1 U7741 ( .A(n9047), .ZN(n9101) );
  INV_X1 U7742 ( .A(n15859), .ZN(n13420) );
  OR2_X1 U7743 ( .A1(n10686), .A2(n9570), .ZN(n9860) );
  OR2_X1 U7744 ( .A1(n9375), .A2(n9374), .ZN(n9386) );
  OAI21_X1 U7745 ( .B1(n9489), .B2(P3_IR_REG_20__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9488) );
  OAI21_X1 U7746 ( .B1(n9238), .B2(n7813), .A(n7811), .ZN(n9300) );
  INV_X1 U7747 ( .A(n7812), .ZN(n7811) );
  OAI21_X1 U7748 ( .B1(n7814), .B2(n7813), .A(n9292), .ZN(n7812) );
  AND2_X1 U7749 ( .A1(n7773), .A2(n6694), .ZN(n6807) );
  NAND2_X1 U7750 ( .A1(n6800), .A2(n9162), .ZN(n9186) );
  AND2_X1 U7751 ( .A1(n6804), .A2(n6803), .ZN(n6801) );
  OAI21_X1 U7752 ( .B1(n11271), .B2(n13762), .A(n10800), .ZN(n10801) );
  OR2_X1 U7753 ( .A1(n10563), .A2(n10562), .ZN(n10573) );
  INV_X1 U7754 ( .A(n14090), .ZN(n13717) );
  AND2_X1 U7755 ( .A1(n14075), .A2(n14076), .ZN(n14070) );
  NAND2_X1 U7756 ( .A1(n12698), .A2(n6907), .ZN(n7880) );
  INV_X1 U7757 ( .A(n7880), .ZN(n13969) );
  OAI22_X1 U7758 ( .A1(n7879), .A2(n7878), .B1(n11218), .B2(n7880), .ZN(n6906)
         );
  OAI21_X1 U7759 ( .B1(n15614), .B2(n6876), .A(n6874), .ZN(n15626) );
  INV_X1 U7760 ( .A(n6875), .ZN(n6874) );
  INV_X1 U7761 ( .A(n11254), .ZN(n6876) );
  AOI21_X1 U7762 ( .B1(n15653), .B2(n7496), .A(n6583), .ZN(n7495) );
  INV_X1 U7763 ( .A(n11260), .ZN(n7496) );
  OR2_X1 U7764 ( .A1(n7497), .A2(n14131), .ZN(n7494) );
  INV_X1 U7765 ( .A(n15653), .ZN(n7497) );
  NOR2_X1 U7766 ( .A1(n14060), .A2(n7646), .ZN(n7645) );
  INV_X1 U7767 ( .A(n7647), .ZN(n7646) );
  NAND2_X1 U7768 ( .A1(n7275), .A2(n10300), .ZN(n14505) );
  NAND2_X1 U7769 ( .A1(n7325), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n10563) );
  INV_X1 U7770 ( .A(n10620), .ZN(n7915) );
  AND2_X1 U7771 ( .A1(n6912), .A2(n10615), .ZN(n6911) );
  OR2_X1 U7772 ( .A1(n14432), .A2(n14448), .ZN(n7979) );
  NAND2_X1 U7773 ( .A1(n8008), .A2(n6626), .ZN(n14468) );
  NAND2_X1 U7774 ( .A1(n12016), .A2(n6904), .ZN(n10592) );
  NOR2_X1 U7775 ( .A1(n11786), .A2(n6905), .ZN(n6904) );
  INV_X1 U7776 ( .A(n10591), .ZN(n6905) );
  INV_X1 U7777 ( .A(n14472), .ZN(n14451) );
  AND2_X1 U7778 ( .A1(n13812), .A2(n14077), .ZN(n11209) );
  NOR2_X1 U7779 ( .A1(n7999), .A2(n6627), .ZN(n7996) );
  XNOR2_X1 U7780 ( .A(n14505), .B(n14059), .ZN(n14494) );
  BUF_X1 U7781 ( .A(n10188), .Z(n10251) );
  INV_X1 U7782 ( .A(n10184), .ZN(n10274) );
  INV_X1 U7783 ( .A(n10292), .ZN(n10188) );
  AND2_X1 U7784 ( .A1(n10347), .A2(n10346), .ZN(n15784) );
  INV_X1 U7785 ( .A(n10333), .ZN(n7119) );
  INV_X1 U7786 ( .A(n10163), .ZN(n7118) );
  NAND2_X1 U7787 ( .A1(n6757), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6756) );
  XNOR2_X1 U7788 ( .A(n10351), .B(n12438), .ZN(n12037) );
  OR2_X1 U7789 ( .A1(n10227), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n10230) );
  NAND2_X1 U7790 ( .A1(n10164), .A2(n10177), .ZN(n10182) );
  NAND2_X1 U7791 ( .A1(n8132), .A2(n8119), .ZN(n10180) );
  NAND2_X1 U7792 ( .A1(n8098), .A2(n6558), .ZN(n8682) );
  NAND2_X1 U7793 ( .A1(n10017), .A2(n10016), .ZN(n7328) );
  NOR2_X1 U7794 ( .A1(n8084), .A2(n10000), .ZN(n10009) );
  NAND2_X1 U7795 ( .A1(n8093), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8367) );
  INV_X1 U7796 ( .A(n8354), .ZN(n8093) );
  OR2_X1 U7797 ( .A1(n10132), .A2(n10865), .ZN(n10138) );
  OR2_X1 U7798 ( .A1(n8808), .A2(n8788), .ZN(n8801) );
  INV_X1 U7799 ( .A(n6514), .ZN(n8688) );
  AND4_X1 U7800 ( .A1(n8433), .A2(n8432), .A3(n8431), .A4(n8430), .ZN(n14785)
         );
  AND4_X1 U7801 ( .A1(n8388), .A2(n8387), .A3(n8386), .A4(n8385), .ZN(n12169)
         );
  NAND2_X1 U7802 ( .A1(n14835), .A2(n15256), .ZN(n8962) );
  INV_X1 U7803 ( .A(n8912), .ZN(n8957) );
  AND2_X1 U7804 ( .A1(n14989), .A2(n14995), .ZN(n8912) );
  INV_X1 U7805 ( .A(n7555), .ZN(n7554) );
  OAI21_X1 U7806 ( .B1(n15021), .B2(n6559), .A(n8040), .ZN(n7555) );
  NAND2_X1 U7807 ( .A1(n15289), .A2(n15032), .ZN(n8040) );
  OR2_X1 U7808 ( .A1(n15319), .A2(n15117), .ZN(n7545) );
  OR2_X1 U7809 ( .A1(n15571), .A2(n15163), .ZN(n10140) );
  NOR2_X1 U7810 ( .A1(n15339), .A2(n15140), .ZN(n8905) );
  NAND2_X1 U7811 ( .A1(n11992), .A2(n8930), .ZN(n12192) );
  AND2_X1 U7812 ( .A1(n10758), .A2(n10888), .ZN(n15257) );
  NAND2_X1 U7813 ( .A1(n10724), .A2(n10876), .ZN(n10865) );
  NOR2_X1 U7814 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n8105) );
  NOR2_X1 U7815 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n8104) );
  NAND2_X1 U7816 ( .A1(n8013), .A2(n8012), .ZN(n8110) );
  NAND2_X1 U7817 ( .A1(n8109), .A2(n8018), .ZN(n8012) );
  OAI21_X1 U7818 ( .B1(n8109), .B2(n8019), .A(n8014), .ZN(n8011) );
  NAND2_X1 U7819 ( .A1(n8109), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7659) );
  NAND2_X1 U7820 ( .A1(n8607), .A2(n8592), .ZN(n8610) );
  NAND2_X1 U7821 ( .A1(n8502), .A2(n8501), .ZN(n6845) );
  CLKBUF_X1 U7822 ( .A(n8125), .Z(n10879) );
  NAND2_X1 U7823 ( .A1(n10180), .A2(n8247), .ZN(n7816) );
  XNOR2_X1 U7824 ( .A(n6746), .B(n9721), .ZN(n9724) );
  NAND2_X1 U7825 ( .A1(n7335), .A2(n6747), .ZN(n6746) );
  NAND2_X1 U7826 ( .A1(n12249), .A2(P1_ADDR_REG_1__SCAN_IN), .ZN(n6747) );
  NAND2_X1 U7827 ( .A1(n6742), .A2(n6741), .ZN(n9731) );
  NAND2_X1 U7828 ( .A1(n15919), .A2(n6585), .ZN(n6742) );
  OAI21_X1 U7829 ( .B1(n7181), .B2(n6578), .A(n6752), .ZN(n15444) );
  INV_X1 U7830 ( .A(n6753), .ZN(n6752) );
  OAI21_X1 U7831 ( .B1(n6578), .B2(n7183), .A(n7563), .ZN(n6753) );
  NAND2_X1 U7832 ( .A1(n15468), .A2(n7564), .ZN(n7563) );
  NOR2_X1 U7833 ( .A1(n9766), .A2(n9765), .ZN(n9770) );
  OR2_X1 U7834 ( .A1(n6950), .A2(n6584), .ZN(n6946) );
  INV_X1 U7835 ( .A(n6949), .ZN(n6948) );
  NAND2_X1 U7836 ( .A1(n9478), .A2(n9477), .ZN(n13196) );
  AND4_X1 U7837 ( .A1(n9153), .A2(n9152), .A3(n9151), .A4(n9150), .ZN(n11944)
         );
  INV_X1 U7838 ( .A(n13336), .ZN(n12792) );
  INV_X1 U7839 ( .A(n13808), .ZN(n13733) );
  OR2_X1 U7840 ( .A1(n10721), .A2(n12673), .ZN(n6976) );
  AOI211_X1 U7841 ( .C1(n14496), .C2(n10715), .A(n14425), .B(n14192), .ZN(
        n10721) );
  AOI21_X1 U7842 ( .B1(n10650), .B2(n15759), .A(n13631), .ZN(n14211) );
  AND2_X1 U7843 ( .A1(n15500), .A2(n15256), .ZN(n14773) );
  NOR2_X1 U7844 ( .A1(n8810), .A2(n8762), .ZN(n8790) );
  OAI21_X1 U7845 ( .B1(n10668), .B2(n8750), .A(n8116), .ZN(n14837) );
  NAND2_X1 U7846 ( .A1(n15451), .A2(n15452), .ZN(n15448) );
  NAND2_X1 U7847 ( .A1(n6738), .A2(n7296), .ZN(n15450) );
  INV_X1 U7848 ( .A(n9725), .ZN(n7296) );
  INV_X1 U7849 ( .A(n6739), .ZN(n6738) );
  NAND2_X1 U7850 ( .A1(n6755), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n9746) );
  NAND2_X1 U7851 ( .A1(n7388), .A2(n7387), .ZN(n9747) );
  INV_X1 U7852 ( .A(n15464), .ZN(n7387) );
  NAND2_X1 U7853 ( .A1(n15483), .A2(n6751), .ZN(n15489) );
  NAND2_X1 U7854 ( .A1(n7167), .A2(n9755), .ZN(n6751) );
  OR2_X1 U7855 ( .A1(n15489), .A2(n15488), .ZN(n7729) );
  INV_X1 U7856 ( .A(n7290), .ZN(n7289) );
  OAI21_X1 U7857 ( .B1(n8311), .B2(n8883), .A(n8310), .ZN(n7290) );
  NAND2_X1 U7858 ( .A1(n7171), .A2(n7170), .ZN(n8310) );
  INV_X1 U7859 ( .A(n13854), .ZN(n6766) );
  NOR2_X1 U7860 ( .A1(n13853), .A2(n13854), .ZN(n6767) );
  INV_X1 U7861 ( .A(n13857), .ZN(n6771) );
  OAI21_X1 U7862 ( .B1(n12923), .B2(n13011), .A(n12924), .ZN(n7100) );
  NAND2_X1 U7863 ( .A1(n6786), .A2(n7718), .ZN(n6785) );
  NAND2_X1 U7864 ( .A1(n13872), .A2(n13871), .ZN(n6786) );
  AOI21_X1 U7865 ( .B1(n7460), .B2(n7458), .A(n7457), .ZN(n7456) );
  NOR2_X1 U7866 ( .A1(n7459), .A2(n8402), .ZN(n7460) );
  AND2_X1 U7867 ( .A1(n7458), .A2(n7457), .ZN(n7172) );
  AOI21_X1 U7868 ( .B1(n7580), .B2(n7581), .A(n7579), .ZN(n7578) );
  NAND2_X1 U7869 ( .A1(n7101), .A2(n7097), .ZN(n12931) );
  NAND2_X1 U7870 ( .A1(n7077), .A2(n7075), .ZN(n7074) );
  INV_X1 U7871 ( .A(n7079), .ZN(n7075) );
  INV_X1 U7872 ( .A(n13370), .ZN(n7082) );
  NAND2_X1 U7873 ( .A1(n7092), .A2(n7090), .ZN(n7087) );
  AOI21_X1 U7874 ( .B1(n7092), .B2(n6616), .A(n13263), .ZN(n7086) );
  NAND2_X1 U7875 ( .A1(n7090), .A2(n7089), .ZN(n7088) );
  NAND2_X1 U7876 ( .A1(n13884), .A2(n13886), .ZN(n7720) );
  NOR2_X1 U7877 ( .A1(n8596), .A2(n8595), .ZN(n7452) );
  NOR2_X1 U7878 ( .A1(n7453), .A2(n7454), .ZN(n7449) );
  AND2_X1 U7879 ( .A1(n8596), .A2(n8595), .ZN(n7454) );
  NAND2_X1 U7880 ( .A1(n7265), .A2(n6625), .ZN(n13955) );
  NAND2_X1 U7881 ( .A1(n6546), .A2(n7723), .ZN(n6783) );
  INV_X1 U7882 ( .A(n13894), .ZN(n7725) );
  INV_X1 U7883 ( .A(n9808), .ZN(n7963) );
  NAND2_X1 U7884 ( .A1(n13369), .A2(n7064), .ZN(n7063) );
  NOR2_X1 U7885 ( .A1(n13391), .A2(n7065), .ZN(n7064) );
  NOR3_X1 U7886 ( .A1(n12880), .A2(n12878), .A3(n7068), .ZN(n12882) );
  NAND2_X1 U7887 ( .A1(n9508), .A2(n7069), .ZN(n7068) );
  AND2_X1 U7888 ( .A1(n13001), .A2(n13002), .ZN(n7772) );
  INV_X1 U7889 ( .A(n9409), .ZN(n7806) );
  NOR2_X1 U7890 ( .A1(n10456), .A2(n10446), .ZN(n6967) );
  INV_X1 U7891 ( .A(n10447), .ZN(n10362) );
  INV_X1 U7892 ( .A(n8952), .ZN(n6847) );
  NOR2_X1 U7893 ( .A1(n15134), .A2(n8035), .ZN(n8034) );
  INV_X1 U7894 ( .A(n8181), .ZN(n6990) );
  NAND2_X1 U7895 ( .A1(n8182), .A2(SI_21_), .ZN(n8185) );
  NAND2_X1 U7896 ( .A1(n8150), .A2(n10901), .ZN(n8153) );
  NAND2_X1 U7897 ( .A1(n7384), .A2(n6873), .ZN(n8137) );
  NAND2_X1 U7898 ( .A1(n10878), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7384) );
  OR2_X1 U7899 ( .A1(n10878), .A2(n9118), .ZN(n6873) );
  OAI21_X1 U7900 ( .B1(n9719), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6649), .ZN(
        n7569) );
  INV_X1 U7901 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n9697) );
  NOR2_X1 U7902 ( .A1(n7967), .A2(n7966), .ZN(n7965) );
  INV_X1 U7903 ( .A(n12749), .ZN(n7966) );
  OAI21_X1 U7904 ( .B1(n7612), .B2(n7611), .A(n10833), .ZN(n7613) );
  NAND2_X1 U7905 ( .A1(n7525), .A2(n7533), .ZN(n7039) );
  INV_X1 U7906 ( .A(n11174), .ZN(n7435) );
  NAND2_X1 U7907 ( .A1(n11893), .A2(n6706), .ZN(n7383) );
  NAND2_X1 U7908 ( .A1(n7243), .A2(n6737), .ZN(n7125) );
  AND2_X1 U7909 ( .A1(n7620), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n6737) );
  INV_X1 U7910 ( .A(n9681), .ZN(n7418) );
  INV_X1 U7911 ( .A(n6720), .ZN(n7412) );
  OR2_X1 U7912 ( .A1(n13443), .A2(n13249), .ZN(n13004) );
  AND2_X1 U7913 ( .A1(n13004), .A2(n13008), .ZN(n13002) );
  INV_X1 U7914 ( .A(n9397), .ZN(n7153) );
  NOR2_X1 U7915 ( .A1(n13245), .A2(n7925), .ZN(n7924) );
  NOR2_X1 U7916 ( .A1(n12988), .A2(n12986), .ZN(n7869) );
  INV_X1 U7917 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n12303) );
  INV_X1 U7918 ( .A(n9362), .ZN(n9341) );
  INV_X1 U7919 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n9250) );
  AND2_X1 U7920 ( .A1(n7046), .A2(n9177), .ZN(n7045) );
  INV_X1 U7921 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n7046) );
  INV_X1 U7922 ( .A(n9128), .ZN(n7052) );
  AND2_X1 U7923 ( .A1(n12878), .A2(n9108), .ZN(n7608) );
  NAND2_X1 U7924 ( .A1(n12919), .A2(n12923), .ZN(n12878) );
  INV_X1 U7925 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n9074) );
  OAI21_X1 U7926 ( .B1(n11660), .B2(n12897), .A(n7156), .ZN(n15851) );
  NAND2_X1 U7927 ( .A1(n13042), .A2(n11661), .ZN(n12900) );
  AOI21_X1 U7928 ( .B1(n7899), .B2(n7897), .A(n12963), .ZN(n7896) );
  INV_X1 U7929 ( .A(n7899), .ZN(n7898) );
  INV_X1 U7930 ( .A(n9517), .ZN(n7897) );
  AND2_X1 U7931 ( .A1(n7876), .A2(n13405), .ZN(n7875) );
  NAND2_X1 U7932 ( .A1(n13416), .A2(n9512), .ZN(n7876) );
  NOR2_X1 U7933 ( .A1(n6831), .A2(n12945), .ZN(n6828) );
  INV_X1 U7934 ( .A(n7875), .ZN(n6831) );
  AOI21_X1 U7935 ( .B1(n7875), .B2(n12948), .A(n12949), .ZN(n7873) );
  NAND2_X1 U7936 ( .A1(n11634), .A2(n12905), .ZN(n11633) );
  NAND2_X1 U7937 ( .A1(n9411), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9425) );
  INV_X1 U7938 ( .A(n7797), .ZN(n7790) );
  AND2_X1 U7939 ( .A1(n6599), .A2(n8079), .ZN(n7588) );
  INV_X1 U7940 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n9336) );
  NOR2_X1 U7941 ( .A1(n9315), .A2(n7798), .ZN(n7797) );
  AND2_X1 U7942 ( .A1(n12251), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n9315) );
  INV_X1 U7943 ( .A(n9301), .ZN(n7798) );
  NOR2_X1 U7944 ( .A1(n10910), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n7780) );
  AND2_X1 U7945 ( .A1(n13637), .A2(n13633), .ZN(n12618) );
  INV_X1 U7946 ( .A(n12649), .ZN(n7682) );
  AOI22_X1 U7947 ( .A1(n6570), .A2(n7711), .B1(n7708), .B2(n7709), .ZN(n7706)
         );
  NOR2_X1 U7948 ( .A1(n6570), .A2(n7708), .ZN(n7707) );
  INV_X1 U7949 ( .A(n13904), .ZN(n6764) );
  INV_X1 U7950 ( .A(n7703), .ZN(n7700) );
  AND2_X1 U7951 ( .A1(n14017), .A2(n13990), .ZN(n14004) );
  NOR2_X1 U7952 ( .A1(n14505), .A2(n14184), .ZN(n7647) );
  OR2_X1 U7953 ( .A1(n10639), .A2(n10638), .ZN(n10716) );
  INV_X1 U7954 ( .A(n14030), .ZN(n7990) );
  AND2_X1 U7955 ( .A1(n7326), .A2(n6977), .ZN(n7325) );
  AND2_X1 U7956 ( .A1(n6978), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6977) );
  NAND2_X1 U7957 ( .A1(n7108), .A2(n10528), .ZN(n7107) );
  INV_X1 U7958 ( .A(n10519), .ZN(n7108) );
  INV_X1 U7959 ( .A(n14335), .ZN(n7109) );
  NOR2_X1 U7960 ( .A1(n10495), .A2(n6971), .ZN(n6970) );
  INV_X1 U7961 ( .A(n10491), .ZN(n10363) );
  INV_X1 U7962 ( .A(n14390), .ZN(n7664) );
  INV_X1 U7963 ( .A(n10593), .ZN(n7906) );
  NOR2_X1 U7964 ( .A1(n8004), .A2(n8000), .ZN(n7999) );
  OR2_X1 U7965 ( .A1(n10223), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n10199) );
  INV_X1 U7966 ( .A(n8228), .ZN(n6927) );
  INV_X1 U7967 ( .A(n8630), .ZN(n8098) );
  NOR2_X1 U7968 ( .A1(n8582), .A2(n8569), .ZN(n6933) );
  INV_X1 U7969 ( .A(n8570), .ZN(n8097) );
  NAND2_X1 U7970 ( .A1(n10724), .A2(n9877), .ZN(n10059) );
  NAND2_X1 U7971 ( .A1(n8743), .A2(n11828), .ZN(n7195) );
  OR2_X1 U7972 ( .A1(n8970), .A2(n8743), .ZN(n7196) );
  AND2_X1 U7973 ( .A1(n7376), .A2(n15134), .ZN(n7375) );
  NOR2_X1 U7974 ( .A1(n10659), .A2(n8055), .ZN(n8054) );
  INV_X1 U7975 ( .A(n8058), .ZN(n8055) );
  OR2_X1 U7976 ( .A1(n14984), .A2(n14982), .ZN(n14989) );
  OR2_X1 U7977 ( .A1(n8682), .A2(n14817), .ZN(n8684) );
  AND2_X1 U7978 ( .A1(n15045), .A2(n15044), .ZN(n15046) );
  NOR2_X1 U7979 ( .A1(n8063), .A2(n15076), .ZN(n6849) );
  NAND2_X1 U7980 ( .A1(n15224), .A2(n6628), .ZN(n8943) );
  AND2_X1 U7981 ( .A1(n15153), .A2(n8941), .ZN(n8942) );
  AND2_X1 U7982 ( .A1(n15134), .A2(n8944), .ZN(n8064) );
  NAND2_X1 U7983 ( .A1(n8096), .A2(n6929), .ZN(n8570) );
  AND2_X1 U7984 ( .A1(n6930), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6929) );
  INV_X1 U7985 ( .A(n7548), .ZN(n7547) );
  OAI21_X1 U7986 ( .B1(n6572), .B2(n7549), .A(n8903), .ZN(n7548) );
  NAND2_X1 U7987 ( .A1(n8901), .A2(n8902), .ZN(n7549) );
  NOR2_X1 U7988 ( .A1(n15350), .A2(n15342), .ZN(n7850) );
  NAND2_X1 U7989 ( .A1(n6871), .A2(n6870), .ZN(n8940) );
  AND2_X1 U7990 ( .A1(n15173), .A2(n15174), .ZN(n6870) );
  NAND2_X1 U7991 ( .A1(n8938), .A2(n6872), .ZN(n6871) );
  INV_X1 U7992 ( .A(n8939), .ZN(n6872) );
  NAND2_X1 U7993 ( .A1(n8898), .A2(n15228), .ZN(n8939) );
  NOR2_X1 U7994 ( .A1(n11996), .A2(n7845), .ZN(n7844) );
  NAND2_X1 U7995 ( .A1(n15372), .A2(n7846), .ZN(n7845) );
  INV_X1 U7996 ( .A(n15581), .ZN(n7855) );
  NOR2_X1 U7997 ( .A1(n11576), .A2(n11700), .ZN(n7856) );
  NAND2_X1 U7998 ( .A1(n11828), .A2(n8958), .ZN(n9877) );
  NAND2_X1 U7999 ( .A1(n8918), .A2(n8829), .ZN(n8917) );
  NOR2_X1 U8000 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n7201) );
  NAND2_X1 U8001 ( .A1(n8758), .A2(n8757), .ZN(n8735) );
  OAI21_X1 U8002 ( .B1(n8774), .B2(n8773), .A(n8708), .ZN(n8758) );
  NOR2_X1 U8003 ( .A1(n8668), .A2(n7832), .ZN(n7831) );
  INV_X1 U8004 ( .A(n8194), .ZN(n7832) );
  NAND2_X1 U8005 ( .A1(n7247), .A2(n7246), .ZN(n8187) );
  INV_X1 U8006 ( .A(n8186), .ZN(n7247) );
  NAND2_X1 U8007 ( .A1(n7822), .A2(n7826), .ZN(n8562) );
  NAND2_X1 U8008 ( .A1(n8165), .A2(n11014), .ZN(n8520) );
  NAND2_X1 U8009 ( .A1(n8519), .A2(n11044), .ZN(n6869) );
  NAND2_X1 U8010 ( .A1(n6866), .A2(SI_14_), .ZN(n6868) );
  INV_X1 U8011 ( .A(n8394), .ZN(n7014) );
  AND2_X1 U8012 ( .A1(n7009), .A2(n8147), .ZN(n7008) );
  NAND2_X1 U8013 ( .A1(n8145), .A2(n6676), .ZN(n7009) );
  NAND2_X1 U8014 ( .A1(n8136), .A2(n8135), .ZN(n8214) );
  XNOR2_X1 U8015 ( .A(n8137), .B(SI_5_), .ZN(n8215) );
  NAND2_X1 U8016 ( .A1(n9721), .A2(n9695), .ZN(n7336) );
  XNOR2_X1 U8017 ( .A(n14877), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n9720) );
  NAND2_X1 U8018 ( .A1(n6748), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7335) );
  XNOR2_X1 U8019 ( .A(n7569), .B(n9697), .ZN(n7730) );
  OAI22_X1 U8020 ( .A1(n9735), .A2(n9704), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n9703), .ZN(n9705) );
  INV_X1 U8021 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n9703) );
  OAI21_X1 U8022 ( .B1(n7930), .B2(n6950), .A(n12806), .ZN(n6949) );
  NAND2_X1 U8023 ( .A1(n12742), .A2(n7952), .ZN(n7948) );
  NAND2_X1 U8024 ( .A1(n12789), .A2(n12788), .ZN(n7950) );
  NAND2_X1 U8025 ( .A1(n9224), .A2(n9223), .ZN(n12954) );
  NAND2_X1 U8026 ( .A1(n7933), .A2(n7936), .ZN(n7932) );
  AND2_X1 U8027 ( .A1(n9791), .A2(n9787), .ZN(n7968) );
  NOR2_X1 U8028 ( .A1(n9825), .A2(n12792), .ZN(n7942) );
  INV_X1 U8029 ( .A(n13421), .ZN(n12531) );
  NAND2_X1 U8030 ( .A1(n6944), .A2(n6943), .ZN(n6942) );
  INV_X1 U8031 ( .A(n9832), .ZN(n6943) );
  AOI21_X1 U8032 ( .B1(n7930), .B2(n12761), .A(n6641), .ZN(n7929) );
  NAND2_X1 U8033 ( .A1(n12752), .A2(n9846), .ZN(n12818) );
  OAI21_X1 U8034 ( .B1(n13191), .B2(n7238), .A(n7294), .ZN(n7293) );
  NOR2_X1 U8035 ( .A1(n12870), .A2(n7295), .ZN(n7294) );
  NOR2_X1 U8036 ( .A1(n13032), .A2(n13507), .ZN(n7295) );
  NAND2_X1 U8037 ( .A1(n13018), .A2(n13019), .ZN(n7575) );
  INV_X1 U8038 ( .A(n9346), .ZN(n12855) );
  NOR2_X1 U8039 ( .A1(n9112), .A2(n6614), .ZN(n7071) );
  NAND2_X1 U8040 ( .A1(n9466), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9024) );
  NAND2_X1 U8041 ( .A1(n11132), .A2(n11133), .ZN(n11131) );
  INV_X1 U8042 ( .A(n7613), .ZN(n7617) );
  NOR2_X1 U8043 ( .A1(n9641), .A2(n9640), .ZN(n7441) );
  INV_X1 U8044 ( .A(n11148), .ZN(n7443) );
  NAND3_X1 U8045 ( .A1(n7625), .A2(n7622), .A3(n6733), .ZN(n11197) );
  INV_X1 U8046 ( .A(n7623), .ZN(n7622) );
  OAI21_X1 U8047 ( .B1(n7624), .B2(n9592), .A(P3_REG2_REG_5__SCAN_IN), .ZN(
        n7623) );
  NAND2_X1 U8048 ( .A1(n11185), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7619) );
  AND2_X1 U8049 ( .A1(n7618), .A2(n11297), .ZN(n9593) );
  NOR2_X1 U8050 ( .A1(n11175), .A2(n7271), .ZN(n9624) );
  NOR2_X1 U8051 ( .A1(n9644), .A2(n15915), .ZN(n7271) );
  AOI21_X1 U8052 ( .B1(n11547), .B2(n11545), .A(n11546), .ZN(n11549) );
  NAND2_X1 U8053 ( .A1(n7127), .A2(n7126), .ZN(n11893) );
  INV_X1 U8054 ( .A(n11890), .ZN(n7126) );
  NAND2_X1 U8055 ( .A1(n11891), .A2(n11889), .ZN(n7127) );
  NAND2_X1 U8056 ( .A1(n7420), .A2(n7419), .ZN(n13059) );
  NAND2_X1 U8057 ( .A1(n7422), .A2(n7429), .ZN(n7419) );
  INV_X1 U8058 ( .A(n13055), .ZN(n7036) );
  OR2_X1 U8059 ( .A1(n13054), .A2(n6553), .ZN(n7513) );
  AND2_X1 U8060 ( .A1(n13055), .A2(n10998), .ZN(n7515) );
  NAND2_X1 U8061 ( .A1(n13083), .A2(n13066), .ZN(n6731) );
  OR2_X1 U8062 ( .A1(n9599), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n6730) );
  XNOR2_X1 U8063 ( .A(n9630), .B(n7404), .ZN(n13113) );
  XNOR2_X1 U8064 ( .A(n9677), .B(n7404), .ZN(n13107) );
  AND2_X1 U8065 ( .A1(n13124), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7133) );
  NAND2_X1 U8066 ( .A1(n13125), .A2(n13124), .ZN(n7132) );
  NAND2_X1 U8067 ( .A1(n13113), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n13112) );
  INV_X1 U8068 ( .A(n13148), .ZN(n7413) );
  AOI21_X1 U8069 ( .B1(n6529), .B2(n6720), .A(n7416), .ZN(n7415) );
  INV_X1 U8070 ( .A(n13118), .ZN(n7416) );
  NAND2_X1 U8071 ( .A1(n7137), .A2(n9602), .ZN(n7628) );
  INV_X1 U8072 ( .A(n7138), .ZN(n7137) );
  NAND2_X1 U8073 ( .A1(n7136), .A2(n9604), .ZN(n13159) );
  OAI21_X1 U8074 ( .B1(n13153), .B2(n13468), .A(n7536), .ZN(n13177) );
  NAND2_X1 U8075 ( .A1(n9633), .A2(n11066), .ZN(n7536) );
  OR2_X1 U8076 ( .A1(n9479), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n13186) );
  NAND2_X1 U8077 ( .A1(n9463), .A2(n9867), .ZN(n9479) );
  INV_X1 U8078 ( .A(n9464), .ZN(n9463) );
  NAND2_X1 U8079 ( .A1(n9473), .A2(n13010), .ZN(n12890) );
  NAND2_X1 U8080 ( .A1(n6826), .A2(n13004), .ZN(n13223) );
  OAI21_X1 U8081 ( .B1(n13262), .B2(n6825), .A(n6824), .ZN(n6826) );
  AOI21_X1 U8082 ( .B1(n7924), .B2(n13263), .A(n6659), .ZN(n6824) );
  INV_X1 U8083 ( .A(n7924), .ZN(n6825) );
  INV_X1 U8084 ( .A(n13215), .ZN(n13224) );
  NAND2_X1 U8085 ( .A1(n9431), .A2(n9430), .ZN(n9447) );
  INV_X1 U8086 ( .A(n9432), .ZN(n9431) );
  INV_X1 U8087 ( .A(n13002), .ZN(n13232) );
  NAND2_X1 U8088 ( .A1(n13262), .A2(n12888), .ZN(n9528) );
  NAND2_X1 U8089 ( .A1(n9528), .A2(n7924), .ZN(n13250) );
  NAND2_X1 U8090 ( .A1(n13272), .A2(n9397), .ZN(n7155) );
  AND2_X1 U8091 ( .A1(n7155), .A2(n6598), .ZN(n13258) );
  NAND2_X1 U8092 ( .A1(n9251), .A2(n6705), .ZN(n9323) );
  INV_X1 U8093 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n7040) );
  NAND2_X1 U8094 ( .A1(n9251), .A2(n7041), .ZN(n9294) );
  AOI21_X1 U8095 ( .B1(n7160), .B2(n7163), .A(n6657), .ZN(n7158) );
  INV_X1 U8096 ( .A(n9184), .ZN(n7163) );
  CLKBUF_X1 U8097 ( .A(n11847), .Z(n7324) );
  INV_X1 U8098 ( .A(n12913), .ZN(n6821) );
  AOI21_X1 U8099 ( .B1(n7893), .B2(n7892), .A(n7891), .ZN(n7890) );
  INV_X1 U8100 ( .A(n12923), .ZN(n7891) );
  INV_X1 U8101 ( .A(n9510), .ZN(n7892) );
  NOR2_X1 U8102 ( .A1(n7894), .A2(n12922), .ZN(n7893) );
  CLKBUF_X1 U8103 ( .A(n11688), .Z(n11689) );
  INV_X1 U8104 ( .A(n12878), .ZN(n12918) );
  NAND2_X1 U8105 ( .A1(n6822), .A2(n12913), .ZN(n11535) );
  CLKBUF_X1 U8106 ( .A(n11536), .Z(n7321) );
  NAND2_X1 U8107 ( .A1(n9075), .A2(n9074), .ZN(n9087) );
  XNOR2_X1 U8108 ( .A(n13040), .B(n15885), .ZN(n12905) );
  INV_X1 U8109 ( .A(n13170), .ZN(n12895) );
  INV_X1 U8110 ( .A(n11092), .ZN(n11661) );
  OR2_X1 U8111 ( .A1(n11327), .A2(n13044), .ZN(n12897) );
  NAND2_X1 U8112 ( .A1(n9446), .A2(n9445), .ZN(n13438) );
  NAND2_X1 U8113 ( .A1(n9415), .A2(n9414), .ZN(n9835) );
  NAND2_X1 U8114 ( .A1(n6796), .A2(n6795), .ZN(n13272) );
  NAND2_X1 U8115 ( .A1(n13346), .A2(n13345), .ZN(n9314) );
  AOI21_X1 U8116 ( .B1(n13281), .B2(n7604), .A(n7603), .ZN(n7602) );
  INV_X1 U8117 ( .A(n8078), .ZN(n7604) );
  NAND2_X1 U8118 ( .A1(n13281), .A2(n13282), .ZN(n9383) );
  INV_X1 U8119 ( .A(n13281), .ZN(n7605) );
  NAND2_X1 U8120 ( .A1(n13302), .A2(n12983), .ZN(n13280) );
  NAND2_X1 U8121 ( .A1(n9526), .A2(n9525), .ZN(n13286) );
  NAND2_X1 U8122 ( .A1(n6840), .A2(n9524), .ZN(n13302) );
  NAND2_X1 U8123 ( .A1(n13295), .A2(n9519), .ZN(n6840) );
  NAND2_X1 U8124 ( .A1(n13006), .A2(n9504), .ZN(n15859) );
  NAND2_X1 U8125 ( .A1(n9314), .A2(n8078), .ZN(n13331) );
  NAND2_X1 U8126 ( .A1(n7159), .A2(n9184), .ZN(n12146) );
  NAND2_X1 U8127 ( .A1(n12090), .A2(n7164), .ZN(n7159) );
  NAND2_X1 U8128 ( .A1(n12147), .A2(n12942), .ZN(n6832) );
  INV_X1 U8129 ( .A(n15901), .ZN(n13499) );
  OR2_X1 U8130 ( .A1(n13023), .A2(n13028), .ZN(n15886) );
  NOR2_X1 U8131 ( .A1(n10878), .A2(n10837), .ZN(n6842) );
  OAI21_X1 U8132 ( .B1(n9557), .B2(P3_D_REG_0__SCAN_IN), .A(n9559), .ZN(n9775)
         );
  NAND2_X1 U8133 ( .A1(n7800), .A2(n7799), .ZN(n12552) );
  AOI21_X1 U8134 ( .B1(n7801), .B2(n9457), .A(n6719), .ZN(n7799) );
  NOR2_X1 U8135 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), .ZN(
        n7401) );
  NOR2_X1 U8136 ( .A1(n7921), .A2(n9102), .ZN(n7402) );
  NOR2_X1 U8137 ( .A1(n9102), .A2(n7919), .ZN(n7292) );
  INV_X1 U8138 ( .A(n8080), .ZN(n7919) );
  AND2_X1 U8139 ( .A1(n7970), .A2(n9575), .ZN(n7969) );
  AOI21_X1 U8140 ( .B1(n7808), .B2(n9374), .A(n6713), .ZN(n7807) );
  NOR2_X1 U8141 ( .A1(n9398), .A2(n7809), .ZN(n7808) );
  INV_X1 U8142 ( .A(n9385), .ZN(n7809) );
  NOR2_X1 U8143 ( .A1(n9492), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n7972) );
  NAND2_X1 U8144 ( .A1(n9372), .A2(n9371), .ZN(n9375) );
  NAND2_X1 U8145 ( .A1(n9332), .A2(n9331), .ZN(n9334) );
  NOR2_X1 U8146 ( .A1(n9354), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n9487) );
  INV_X1 U8147 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9486) );
  AND2_X1 U8148 ( .A1(n7793), .A2(n7795), .ZN(n7792) );
  INV_X1 U8149 ( .A(n9350), .ZN(n7793) );
  NAND2_X1 U8150 ( .A1(n9302), .A2(n7797), .ZN(n7794) );
  NAND2_X1 U8151 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n7796), .ZN(n7795) );
  AND2_X1 U8152 ( .A1(n9274), .A2(n9273), .ZN(n9275) );
  NAND2_X1 U8153 ( .A1(n6806), .A2(n6621), .ZN(n9238) );
  INV_X1 U8154 ( .A(n9234), .ZN(n7334) );
  NOR2_X1 U8155 ( .A1(n9276), .A2(n7815), .ZN(n7814) );
  INV_X1 U8156 ( .A(n9237), .ZN(n7815) );
  NAND2_X1 U8157 ( .A1(n9258), .A2(n6577), .ZN(n9493) );
  AOI21_X1 U8158 ( .B1(n7776), .B2(n7779), .A(n6650), .ZN(n7773) );
  INV_X1 U8159 ( .A(n9189), .ZN(n7779) );
  XNOR2_X1 U8160 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n9201) );
  NAND2_X1 U8161 ( .A1(n6661), .A2(n7782), .ZN(n6804) );
  INV_X1 U8162 ( .A(n7780), .ZN(n6802) );
  XNOR2_X1 U8163 ( .A(n9139), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n9154) );
  INV_X1 U8164 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9139) );
  INV_X1 U8165 ( .A(n7785), .ZN(n7784) );
  AOI21_X1 U8166 ( .B1(n7785), .B2(n9115), .A(n7783), .ZN(n7782) );
  INV_X1 U8167 ( .A(n9136), .ZN(n7783) );
  AND2_X1 U8168 ( .A1(n9136), .A2(n9120), .ZN(n9135) );
  INV_X1 U8169 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n9121) );
  OAI211_X1 U8170 ( .C1(n6793), .C2(n6790), .A(n6788), .B(n9096), .ZN(n9100)
         );
  INV_X1 U8171 ( .A(n9082), .ZN(n6790) );
  NOR2_X1 U8172 ( .A1(n9083), .A2(n6792), .ZN(n6791) );
  AND2_X1 U8173 ( .A1(n10839), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9083) );
  INV_X1 U8174 ( .A(n9067), .ZN(n6792) );
  XNOR2_X1 U8175 ( .A(n9098), .B(P1_DATAO_REG_4__SCAN_IN), .ZN(n9095) );
  INV_X1 U8176 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7282) );
  XNOR2_X1 U8177 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .ZN(n9049) );
  NAND2_X1 U8178 ( .A1(n10178), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9048) );
  NOR3_X1 U8179 ( .A1(n14674), .A2(n12548), .A3(n12160), .ZN(n10725) );
  OR2_X1 U8180 ( .A1(n10381), .A2(n15804), .ZN(n10382) );
  OR2_X1 U8181 ( .A1(n7879), .A2(n7274), .ZN(n10384) );
  OR2_X1 U8182 ( .A1(n10509), .A2(n10508), .ZN(n10521) );
  NAND2_X1 U8183 ( .A1(n7217), .A2(n7215), .ZN(n13625) );
  AOI21_X1 U8184 ( .B1(n7364), .B2(n7218), .A(n6545), .ZN(n7217) );
  NAND2_X1 U8185 ( .A1(n7208), .A2(n12634), .ZN(n7207) );
  INV_X1 U8186 ( .A(n13708), .ZN(n7208) );
  NAND2_X1 U8187 ( .A1(n12644), .A2(n13669), .ZN(n7689) );
  AOI21_X1 U8188 ( .B1(n7673), .B2(n7674), .A(n6580), .ZN(n7671) );
  AND2_X1 U8189 ( .A1(n12716), .A2(n12118), .ZN(n12119) );
  AND2_X1 U8190 ( .A1(n13686), .A2(n7221), .ZN(n7220) );
  NAND2_X1 U8191 ( .A1(n12659), .A2(n13714), .ZN(n7221) );
  AND2_X1 U8192 ( .A1(n10570), .A2(n10569), .ZN(n13718) );
  AND4_X1 U8193 ( .A1(n10419), .A2(n10418), .A3(n10417), .A4(n10416), .ZN(
        n13855) );
  NAND2_X1 U8194 ( .A1(n7494), .A2(n6601), .ZN(n15667) );
  INV_X1 U8195 ( .A(n15664), .ZN(n7493) );
  OR2_X1 U8196 ( .A1(n14140), .A2(n7498), .ZN(n6897) );
  NOR2_X1 U8197 ( .A1(n15732), .A2(n7502), .ZN(n14144) );
  AND2_X1 U8198 ( .A1(n15738), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7502) );
  OR2_X1 U8199 ( .A1(n14144), .A2(n14143), .ZN(n7501) );
  NAND2_X1 U8200 ( .A1(n10639), .A2(n10574), .ZN(n14219) );
  INV_X1 U8201 ( .A(n10628), .ZN(n10624) );
  INV_X1 U8202 ( .A(n14282), .ZN(n7988) );
  NOR2_X1 U8203 ( .A1(n14626), .A2(n13671), .ZN(n7986) );
  AND2_X1 U8204 ( .A1(n10558), .A2(n10557), .ZN(n14262) );
  OR2_X1 U8205 ( .A1(n14033), .A2(n14032), .ZN(n14300) );
  NAND2_X1 U8206 ( .A1(n10518), .A2(n10517), .ZN(n10519) );
  NAND2_X1 U8207 ( .A1(n6914), .A2(n10613), .ZN(n14337) );
  NAND2_X1 U8208 ( .A1(n14358), .A2(n14359), .ZN(n6914) );
  INV_X1 U8209 ( .A(n10609), .ZN(n7888) );
  NAND2_X1 U8210 ( .A1(n14573), .A2(n14093), .ZN(n7889) );
  OR2_X1 U8211 ( .A1(n14034), .A2(n6547), .ZN(n14409) );
  INV_X1 U8212 ( .A(n14428), .ZN(n7978) );
  NAND2_X1 U8213 ( .A1(n7655), .A2(n7656), .ZN(n6759) );
  INV_X1 U8214 ( .A(n10428), .ZN(n7111) );
  NOR2_X1 U8215 ( .A1(n7909), .A2(n15765), .ZN(n7908) );
  XNOR2_X1 U8216 ( .A(n13858), .B(n13859), .ZN(n11934) );
  NOR2_X1 U8217 ( .A1(n12013), .A2(n15813), .ZN(n11797) );
  OAI21_X1 U8218 ( .B1(n10185), .B2(n7693), .A(n7692), .ZN(n7691) );
  NAND2_X1 U8219 ( .A1(n11977), .A2(n11905), .ZN(n12012) );
  INV_X1 U8220 ( .A(n14474), .ZN(n14449) );
  NAND2_X1 U8221 ( .A1(n10314), .A2(n11238), .ZN(n14474) );
  AND2_X1 U8222 ( .A1(n10636), .A2(n10635), .ZN(n14425) );
  NAND2_X1 U8223 ( .A1(n7273), .A2(n14191), .ZN(n14193) );
  AND2_X1 U8224 ( .A1(n14505), .A2(n15812), .ZN(n7261) );
  AND2_X1 U8225 ( .A1(n14494), .A2(n14496), .ZN(n14495) );
  AND2_X1 U8226 ( .A1(n14501), .A2(n14500), .ZN(n14502) );
  NAND2_X1 U8227 ( .A1(n14494), .A2(n14499), .ZN(n14500) );
  NAND2_X1 U8228 ( .A1(n7305), .A2(n10301), .ZN(n10281) );
  NAND2_X1 U8229 ( .A1(n11319), .A2(n10251), .ZN(n10258) );
  AND2_X1 U8230 ( .A1(n11209), .A2(n13966), .ZN(n15812) );
  OAI21_X1 U8231 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(n6923), .A(n10320), .ZN(
        n6922) );
  NAND2_X1 U8232 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n6923), .ZN(n10320) );
  NAND2_X1 U8233 ( .A1(n10338), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10351) );
  INV_X1 U8234 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n12438) );
  AND2_X2 U8235 ( .A1(n7366), .A2(n10232), .ZN(n10173) );
  AND2_X1 U8236 ( .A1(n10172), .A2(n10267), .ZN(n7366) );
  AND2_X1 U8237 ( .A1(n10228), .A2(n10230), .ZN(n11263) );
  AND2_X1 U8238 ( .A1(n10204), .A2(n10208), .ZN(n11255) );
  INV_X1 U8239 ( .A(n8083), .ZN(n7747) );
  NAND2_X1 U8240 ( .A1(n6926), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8455) );
  INV_X1 U8241 ( .A(n8453), .ZN(n6926) );
  AND2_X1 U8242 ( .A1(n9964), .A2(n9963), .ZN(n12175) );
  NAND2_X1 U8243 ( .A1(n8092), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8354) );
  INV_X1 U8244 ( .A(n8335), .ZN(n8092) );
  AND2_X1 U8245 ( .A1(n7747), .A2(n11702), .ZN(n7746) );
  AOI21_X1 U8246 ( .B1(n14772), .B2(n14771), .A(n7350), .ZN(n14718) );
  AND2_X1 U8247 ( .A1(n10050), .A2(n10049), .ZN(n7350) );
  AND2_X1 U8248 ( .A1(n7005), .A2(n10097), .ZN(n14735) );
  INV_X1 U8249 ( .A(n14762), .ZN(n7003) );
  NOR2_X1 U8250 ( .A1(n9926), .A2(n11346), .ZN(n7000) );
  NAND2_X1 U8251 ( .A1(n9926), .A2(n11346), .ZN(n6999) );
  NAND2_X1 U8252 ( .A1(n8098), .A2(n6928), .ZN(n8660) );
  NAND2_X1 U8253 ( .A1(n6865), .A2(n14691), .ZN(n14763) );
  NAND2_X1 U8254 ( .A1(n6860), .A2(n6859), .ZN(n6865) );
  AND2_X1 U8255 ( .A1(n6861), .A2(n10068), .ZN(n6859) );
  INV_X1 U8256 ( .A(n9877), .ZN(n7750) );
  INV_X1 U8257 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8366) );
  AND2_X1 U8258 ( .A1(n14700), .A2(n6582), .ZN(n6853) );
  NAND2_X1 U8259 ( .A1(n14718), .A2(n6863), .ZN(n6860) );
  NOR2_X1 U8260 ( .A1(n14792), .A2(n6864), .ZN(n6863) );
  INV_X1 U8261 ( .A(n14717), .ZN(n6864) );
  OR2_X1 U8262 ( .A1(n8367), .A2(n8366), .ZN(n8407) );
  NAND2_X1 U8263 ( .A1(n7018), .A2(n9955), .ZN(n11862) );
  AND2_X1 U8264 ( .A1(n7762), .A2(n7017), .ZN(n7016) );
  AND2_X1 U8265 ( .A1(n9982), .A2(n9971), .ZN(n7762) );
  NAND2_X1 U8266 ( .A1(n6924), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8512) );
  INV_X1 U8267 ( .A(n8479), .ZN(n6924) );
  NOR2_X1 U8268 ( .A1(n8695), .A2(n8692), .ZN(n7194) );
  AND2_X1 U8269 ( .A1(n7468), .A2(n8673), .ZN(n7467) );
  OR2_X1 U8270 ( .A1(n8673), .A2(n7468), .ZN(n7288) );
  NAND2_X1 U8271 ( .A1(n8692), .A2(n8695), .ZN(n7193) );
  INV_X1 U8272 ( .A(n8980), .ZN(n7751) );
  AND4_X1 U8273 ( .A1(n8360), .A2(n8359), .A3(n8358), .A4(n8357), .ZN(n11832)
         );
  OR2_X1 U8274 ( .A1(n8750), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8269) );
  OR2_X1 U8275 ( .A1(n10954), .A2(n10955), .ZN(n10952) );
  OR2_X1 U8276 ( .A1(n11595), .A2(n11596), .ZN(n11593) );
  NAND2_X1 U8277 ( .A1(n8741), .A2(n8740), .ZN(n14977) );
  NAND2_X1 U8278 ( .A1(n8099), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n15005) );
  INV_X1 U8279 ( .A(n8684), .ZN(n8099) );
  OR2_X1 U8280 ( .A1(n7841), .A2(n14984), .ZN(n15002) );
  AND2_X1 U8281 ( .A1(n7554), .A2(n10659), .ZN(n7552) );
  NAND2_X1 U8282 ( .A1(n8955), .A2(n8060), .ZN(n8058) );
  NAND2_X1 U8283 ( .A1(n7301), .A2(n8060), .ZN(n8057) );
  NAND2_X1 U8284 ( .A1(n8059), .A2(n15021), .ZN(n7301) );
  AND2_X1 U8285 ( .A1(n8667), .A2(n8666), .ZN(n14815) );
  OR2_X1 U8286 ( .A1(n15033), .A2(n8750), .ZN(n8667) );
  NOR2_X2 U8287 ( .A1(n15046), .A2(n8954), .ZN(n15040) );
  AND2_X1 U8288 ( .A1(n7858), .A2(n15031), .ZN(n8954) );
  XNOR2_X1 U8289 ( .A(n15053), .B(n15031), .ZN(n15044) );
  NAND2_X1 U8290 ( .A1(n6850), .A2(n6849), .ZN(n15082) );
  NAND2_X1 U8291 ( .A1(n15123), .A2(n7543), .ZN(n7539) );
  INV_X1 U8292 ( .A(n7541), .ZN(n7540) );
  INV_X1 U8293 ( .A(n7545), .ZN(n7542) );
  NAND2_X1 U8294 ( .A1(n8943), .A2(n8942), .ZN(n15155) );
  NAND2_X1 U8295 ( .A1(n15206), .A2(n8895), .ZN(n6966) );
  AOI21_X1 U8296 ( .B1(n8044), .B2(n8046), .A(n6639), .ZN(n8042) );
  NOR2_X1 U8297 ( .A1(n8932), .A2(n8045), .ZN(n8044) );
  NOR2_X1 U8298 ( .A1(n12191), .A2(n8046), .ZN(n8045) );
  INV_X1 U8299 ( .A(n8931), .ZN(n8046) );
  NAND2_X1 U8300 ( .A1(n7559), .A2(n7558), .ZN(n15246) );
  AOI21_X1 U8301 ( .B1(n12189), .B2(n8030), .A(n6638), .ZN(n7558) );
  NAND2_X1 U8302 ( .A1(n12192), .A2(n12191), .ZN(n12190) );
  OAI21_X1 U8303 ( .B1(n11676), .B2(n7484), .A(n7480), .ZN(n11992) );
  NAND2_X1 U8304 ( .A1(n7486), .A2(n8929), .ZN(n7484) );
  NOR2_X1 U8305 ( .A1(n8047), .A2(n7481), .ZN(n7480) );
  NAND2_X1 U8306 ( .A1(n11830), .A2(n6571), .ZN(n11918) );
  INV_X1 U8307 ( .A(n8024), .ZN(n6960) );
  NAND2_X1 U8308 ( .A1(n11674), .A2(n7486), .ZN(n11830) );
  INV_X1 U8309 ( .A(n8926), .ZN(n7487) );
  NAND2_X1 U8310 ( .A1(n11676), .A2(n11675), .ZN(n11674) );
  AND4_X1 U8311 ( .A1(n8318), .A2(n8317), .A3(n8316), .A4(n8315), .ZN(n11703)
         );
  INV_X1 U8312 ( .A(n15257), .ZN(n15225) );
  INV_X1 U8313 ( .A(n15256), .ZN(n15227) );
  AND2_X1 U8314 ( .A1(n10758), .A2(n14874), .ZN(n15256) );
  INV_X1 U8315 ( .A(n14856), .ZN(n7631) );
  NAND2_X1 U8316 ( .A1(n8725), .A2(n8724), .ZN(n15269) );
  OR2_X1 U8317 ( .A1(n15437), .A2(n8679), .ZN(n8681) );
  OR2_X1 U8318 ( .A1(n11913), .A2(n8679), .ZN(n8614) );
  NAND2_X1 U8319 ( .A1(n11779), .A2(n8775), .ZN(n8568) );
  INV_X1 U8320 ( .A(n10907), .ZN(n8253) );
  NAND2_X1 U8321 ( .A1(n8995), .A2(n10875), .ZN(n10654) );
  OR2_X1 U8322 ( .A1(n10867), .A2(P1_D_REG_0__SCAN_IN), .ZN(n8995) );
  AND3_X1 U8323 ( .A1(n10118), .A2(n10140), .A3(n10655), .ZN(n9002) );
  NOR2_X1 U8324 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n8107) );
  INV_X1 U8325 ( .A(n8815), .ZN(n7474) );
  INV_X1 U8326 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8199) );
  INV_X1 U8327 ( .A(n8202), .ZN(n7278) );
  AND2_X1 U8328 ( .A1(n7834), .A2(n6698), .ZN(n7833) );
  NAND2_X1 U8329 ( .A1(n8649), .A2(n7831), .ZN(n7835) );
  INV_X1 U8330 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U8331 ( .A1(n7231), .A2(n7230), .ZN(n10285) );
  INV_X1 U8332 ( .A(n10282), .ZN(n7230) );
  INV_X1 U8333 ( .A(n10283), .ZN(n7231) );
  AOI21_X1 U8334 ( .B1(n7823), .B2(n7825), .A(n7820), .ZN(n7819) );
  INV_X1 U8335 ( .A(n8180), .ZN(n7820) );
  AND2_X1 U8336 ( .A1(n8607), .A2(n8606), .ZN(n8608) );
  NAND2_X1 U8337 ( .A1(n6517), .A2(n7757), .ZN(n8816) );
  AND2_X1 U8338 ( .A1(n7758), .A2(n8209), .ZN(n7757) );
  XNOR2_X1 U8339 ( .A(n8562), .B(SI_18_), .ZN(n8502) );
  OR2_X1 U8340 ( .A1(n8419), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8435) );
  OR2_X1 U8341 ( .A1(n8321), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n8328) );
  XNOR2_X1 U8342 ( .A(n8214), .B(n8215), .ZN(n10863) );
  INV_X1 U8343 ( .A(n8274), .ZN(n8276) );
  CLKBUF_X1 U8344 ( .A(n8273), .Z(n8274) );
  NOR2_X2 U8345 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n8283) );
  INV_X1 U8346 ( .A(P1_RD_REG_SCAN_IN), .ZN(n6957) );
  NAND2_X1 U8347 ( .A1(n7386), .A2(n6603), .ZN(n6739) );
  XNOR2_X1 U8348 ( .A(n7730), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n9728) );
  NOR2_X1 U8349 ( .A1(n15453), .A2(n9737), .ZN(n9739) );
  XNOR2_X1 U8350 ( .A(n9705), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n9718) );
  AOI21_X1 U8351 ( .B1(n9740), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n9707), .ZN(
        n9716) );
  XNOR2_X1 U8352 ( .A(n9709), .B(n14932), .ZN(n9745) );
  NAND2_X1 U8353 ( .A1(n9711), .A2(n7567), .ZN(n9751) );
  NAND2_X1 U8354 ( .A1(P3_ADDR_REG_12__SCAN_IN), .A2(n7568), .ZN(n7567) );
  INV_X1 U8355 ( .A(n7565), .ZN(n9757) );
  OAI21_X1 U8356 ( .B1(n9754), .B2(n9753), .A(n7566), .ZN(n7565) );
  NAND2_X1 U8357 ( .A1(n11623), .A2(P3_ADDR_REG_14__SCAN_IN), .ZN(n7566) );
  AND4_X1 U8358 ( .A1(n9270), .A2(n9269), .A3(n9268), .A4(n9267), .ZN(n13403)
         );
  NAND2_X1 U8359 ( .A1(n9401), .A2(n9400), .ZN(n12728) );
  AND2_X1 U8360 ( .A1(n9358), .A2(n9357), .ZN(n12811) );
  AND2_X1 U8361 ( .A1(n9280), .A2(n9279), .ZN(n12843) );
  OR2_X1 U8362 ( .A1(n9870), .A2(n13027), .ZN(n12836) );
  AND2_X1 U8363 ( .A1(n9851), .A2(n10683), .ZN(n12832) );
  INV_X1 U8364 ( .A(n13323), .ZN(n13288) );
  NAND2_X1 U8365 ( .A1(n9349), .A2(n9348), .ZN(n13336) );
  NAND4_X1 U8366 ( .A1(n9215), .A2(n9214), .A3(n9213), .A4(n9212), .ZN(n13034)
         );
  AND2_X1 U8367 ( .A1(n9132), .A2(n9134), .ZN(n6955) );
  AND2_X1 U8368 ( .A1(n7531), .A2(n6726), .ZN(n11149) );
  NOR2_X1 U8369 ( .A1(n13102), .A2(n13374), .ZN(n13126) );
  NAND2_X1 U8370 ( .A1(n7134), .A2(n9601), .ZN(n13102) );
  XNOR2_X1 U8371 ( .A(n6729), .B(n13165), .ZN(n6728) );
  NAND2_X1 U8372 ( .A1(n13159), .A2(n13158), .ZN(n6729) );
  AOI21_X1 U8373 ( .B1(n13177), .B2(n13176), .A(n7534), .ZN(n13179) );
  NOR2_X1 U8374 ( .A1(n13160), .A2(n7535), .ZN(n7534) );
  NOR2_X1 U8375 ( .A1(n13043), .A2(n9686), .ZN(n13173) );
  OR2_X1 U8376 ( .A1(n13513), .A2(n13431), .ZN(n7252) );
  NAND2_X1 U8377 ( .A1(n13220), .A2(n13219), .ZN(n13221) );
  NAND2_X1 U8378 ( .A1(n12089), .A2(n12930), .ZN(n7865) );
  INV_X1 U8379 ( .A(n11327), .ZN(n11662) );
  AND3_X1 U8380 ( .A1(n11110), .A2(n11109), .A3(n11108), .ZN(n13428) );
  AND2_X1 U8381 ( .A1(n7597), .A2(n7601), .ZN(n7596) );
  NAND2_X1 U8382 ( .A1(n10706), .A2(n13435), .ZN(n7601) );
  OR2_X1 U8383 ( .A1(n13204), .A2(n7598), .ZN(n7597) );
  XNOR2_X1 U8384 ( .A(n7054), .B(n13200), .ZN(n7600) );
  OAI211_X1 U8385 ( .C1(n13199), .C2(n13198), .A(n13197), .B(n6653), .ZN(n7054) );
  NAND2_X1 U8386 ( .A1(n12865), .A2(n12864), .ZN(n13511) );
  OR2_X1 U8387 ( .A1(n13513), .A2(n13593), .ZN(n7253) );
  AOI21_X1 U8388 ( .B1(n7600), .B2(n15864), .A(n13204), .ZN(n13509) );
  NAND2_X1 U8389 ( .A1(n12699), .A2(n9540), .ZN(n10707) );
  NOR2_X1 U8390 ( .A1(n12702), .A2(n13599), .ZN(n9581) );
  NAND2_X1 U8391 ( .A1(n9388), .A2(n9387), .ZN(n13526) );
  NAND2_X1 U8392 ( .A1(n6799), .A2(n9377), .ZN(n13532) );
  NAND2_X1 U8393 ( .A1(n7263), .A2(n7262), .ZN(n6799) );
  INV_X1 U8394 ( .A(n11751), .ZN(n7263) );
  NAND2_X1 U8395 ( .A1(n9308), .A2(n9307), .ZN(n13556) );
  NAND2_X1 U8396 ( .A1(n9249), .A2(n9248), .ZN(n13574) );
  AND2_X1 U8397 ( .A1(n11271), .A2(n13762), .ZN(n7310) );
  NOR2_X1 U8398 ( .A1(n13625), .A2(n13624), .ZN(n13623) );
  NAND2_X1 U8399 ( .A1(n11213), .A2(n10301), .ZN(n7226) );
  INV_X1 U8400 ( .A(n14092), .ZN(n10517) );
  NAND2_X1 U8401 ( .A1(n10250), .A2(n10249), .ZN(n14432) );
  NAND2_X1 U8402 ( .A1(n10238), .A2(n10237), .ZN(n14483) );
  OAI211_X2 U8403 ( .C1(n10292), .C2(n10881), .A(n10187), .B(n10186), .ZN(
        n13813) );
  AND3_X1 U8404 ( .A1(n10504), .A2(n10503), .A3(n10502), .ZN(n14376) );
  INV_X1 U8405 ( .A(n13750), .ZN(n13804) );
  AND2_X1 U8406 ( .A1(n13784), .A2(n12665), .ZN(n7364) );
  NAND2_X1 U8407 ( .A1(n10825), .A2(n15776), .ZN(n13808) );
  INV_X1 U8408 ( .A(n14082), .ZN(n7315) );
  INV_X1 U8409 ( .A(n7317), .ZN(n7316) );
  OAI21_X1 U8410 ( .B1(n14081), .B2(n14080), .A(n14078), .ZN(n7317) );
  NOR3_X1 U8411 ( .A1(n14063), .A2(n14066), .A3(n14073), .ZN(n14064) );
  INV_X1 U8412 ( .A(n14196), .ZN(n14183) );
  NAND2_X1 U8413 ( .A1(n10552), .A2(n10551), .ZN(n14090) );
  OR2_X1 U8414 ( .A1(n14261), .A2(n7879), .ZN(n10552) );
  NAND2_X1 U8415 ( .A1(n10545), .A2(n10544), .ZN(n14263) );
  AND2_X1 U8416 ( .A1(n10372), .A2(n10371), .ZN(n13909) );
  INV_X1 U8417 ( .A(n6906), .ZN(n7877) );
  NAND2_X1 U8418 ( .A1(n14122), .A2(n11252), .ZN(n15614) );
  NAND2_X1 U8419 ( .A1(n15614), .A2(n15615), .ZN(n15613) );
  INV_X1 U8420 ( .A(n6883), .ZN(n6881) );
  NAND2_X1 U8421 ( .A1(n15752), .A2(n14076), .ZN(n6882) );
  NOR2_X1 U8422 ( .A1(n15733), .A2(n14076), .ZN(n6886) );
  AOI21_X1 U8423 ( .B1(n15745), .B2(n14166), .A(P2_REG1_REG_19__SCAN_IN), .ZN(
        n6889) );
  NOR2_X1 U8424 ( .A1(n15733), .A2(n14176), .ZN(n6883) );
  AOI21_X1 U8425 ( .B1(n6885), .B2(n14176), .A(n7503), .ZN(n6884) );
  INV_X1 U8426 ( .A(n7504), .ZN(n6885) );
  AOI21_X1 U8427 ( .B1(n14175), .B2(n15752), .A(n15739), .ZN(n7504) );
  OR2_X1 U8428 ( .A1(n10722), .A2(n14025), .ZN(n7644) );
  NAND2_X1 U8429 ( .A1(n7998), .A2(n8004), .ZN(n10709) );
  XNOR2_X1 U8430 ( .A(n7359), .B(n7358), .ZN(n14514) );
  INV_X1 U8431 ( .A(n14222), .ZN(n7358) );
  AOI21_X1 U8432 ( .B1(n14230), .B2(n10571), .A(n8072), .ZN(n7359) );
  OR2_X1 U8433 ( .A1(n11658), .A2(n10292), .ZN(n10277) );
  AND2_X1 U8434 ( .A1(n15781), .A2(n14076), .ZN(n15770) );
  NAND2_X1 U8435 ( .A1(n10824), .A2(n15796), .ZN(n15776) );
  INV_X1 U8436 ( .A(n10823), .ZN(n10824) );
  NAND2_X1 U8437 ( .A1(n7285), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n7379) );
  NAND2_X1 U8438 ( .A1(n7635), .A2(n11249), .ZN(n7634) );
  INV_X1 U8439 ( .A(n6976), .ZN(n14206) );
  NAND2_X1 U8440 ( .A1(n7330), .A2(n10301), .ZN(n10294) );
  INV_X1 U8441 ( .A(n15437), .ZN(n7330) );
  NAND2_X1 U8442 ( .A1(n10357), .A2(n10356), .ZN(n15792) );
  AND3_X1 U8443 ( .A1(n7119), .A2(n10166), .A3(n6689), .ZN(n7116) );
  INV_X1 U8444 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11873) );
  INV_X1 U8445 ( .A(n10150), .ZN(n7352) );
  AND2_X1 U8446 ( .A1(n7339), .A2(n7340), .ZN(n14757) );
  AOI21_X1 U8447 ( .B1(n10019), .B2(n7329), .A(n14754), .ZN(n7340) );
  NAND2_X1 U8448 ( .A1(n8594), .A2(n8593), .ZN(n15324) );
  NOR2_X1 U8449 ( .A1(n10138), .A2(n10136), .ZN(n15500) );
  NOR2_X2 U8450 ( .A1(n10138), .A2(n10120), .ZN(n14813) );
  INV_X1 U8451 ( .A(n15503), .ZN(n14830) );
  NAND2_X1 U8452 ( .A1(n8801), .A2(n8802), .ZN(n8803) );
  NAND2_X1 U8453 ( .A1(n7371), .A2(n7370), .ZN(n7369) );
  INV_X1 U8454 ( .A(n8869), .ZN(n7370) );
  NAND2_X1 U8455 ( .A1(n8870), .A2(n12005), .ZN(n7371) );
  NAND2_X1 U8456 ( .A1(n8637), .A2(n8636), .ZN(n14839) );
  OR2_X1 U8457 ( .A1(n15068), .A2(n8750), .ZN(n8637) );
  NAND2_X1 U8458 ( .A1(n8604), .A2(n8603), .ZN(n15117) );
  INV_X1 U8459 ( .A(n14785), .ZN(n15258) );
  NAND2_X1 U8460 ( .A1(n8764), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8258) );
  NAND2_X1 U8461 ( .A1(n6514), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8259) );
  AOI21_X1 U8462 ( .B1(n8964), .B2(n15545), .A(n8963), .ZN(n12692) );
  NAND2_X1 U8463 ( .A1(n8962), .A2(n8961), .ZN(n8963) );
  NAND2_X1 U8464 ( .A1(n14837), .A2(n15257), .ZN(n8961) );
  NOR2_X2 U8465 ( .A1(n10865), .A2(n10140), .ZN(n15513) );
  OR2_X1 U8466 ( .A1(n11658), .A2(n8679), .ZN(n8511) );
  OR2_X1 U8467 ( .A1(n15262), .A2(n11384), .ZN(n15267) );
  INV_X1 U8468 ( .A(n15513), .ZN(n15259) );
  OAI21_X1 U8469 ( .B1(n8474), .B2(n8206), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n7446) );
  XNOR2_X1 U8470 ( .A(n9724), .B(n9723), .ZN(n15933) );
  OR2_X1 U8471 ( .A1(n15933), .A2(n15934), .ZN(n7386) );
  NAND2_X1 U8472 ( .A1(n6739), .A2(n9725), .ZN(n15451) );
  XNOR2_X1 U8473 ( .A(n9728), .B(n15625), .ZN(n15919) );
  NAND2_X1 U8474 ( .A1(n9726), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n6744) );
  INV_X1 U8475 ( .A(n15919), .ZN(n6740) );
  OR2_X1 U8476 ( .A1(n15926), .A2(n15927), .ZN(n6749) );
  XNOR2_X1 U8477 ( .A(n6750), .B(n9741), .ZN(n15457) );
  NAND2_X1 U8478 ( .A1(n15457), .A2(n15663), .ZN(n15456) );
  INV_X1 U8479 ( .A(n7388), .ZN(n15463) );
  INV_X1 U8480 ( .A(n9750), .ZN(n7342) );
  NAND2_X1 U8481 ( .A1(n9746), .A2(n9747), .ZN(n7175) );
  NAND2_X1 U8482 ( .A1(n15485), .A2(n15484), .ZN(n15483) );
  OR2_X1 U8483 ( .A1(n15493), .A2(n15742), .ZN(n7182) );
  NAND2_X1 U8484 ( .A1(n15493), .A2(n15742), .ZN(n7183) );
  XNOR2_X1 U8485 ( .A(n9767), .B(n9770), .ZN(n15445) );
  NAND2_X1 U8486 ( .A1(n7447), .A2(n8266), .ZN(n8297) );
  INV_X1 U8487 ( .A(n7156), .ZN(n12902) );
  OR2_X1 U8488 ( .A1(n13844), .A2(n13847), .ZN(n7696) );
  NAND2_X1 U8489 ( .A1(n13006), .A2(n12902), .ZN(n7591) );
  NAND2_X1 U8490 ( .A1(n12899), .A2(n12900), .ZN(n7593) );
  AND2_X1 U8491 ( .A1(n7291), .A2(n7189), .ZN(n7188) );
  AOI21_X1 U8492 ( .B1(n12906), .B2(n13006), .A(n12905), .ZN(n12912) );
  INV_X1 U8493 ( .A(n12904), .ZN(n12906) );
  AOI21_X1 U8494 ( .B1(n7594), .B2(n7592), .A(n7590), .ZN(n12908) );
  NAND2_X1 U8495 ( .A1(n13006), .A2(n7593), .ZN(n7592) );
  NAND2_X1 U8496 ( .A1(n12876), .A2(n7591), .ZN(n7590) );
  NAND2_X1 U8497 ( .A1(n12900), .A2(n12901), .ZN(n7594) );
  NAND2_X1 U8498 ( .A1(n12929), .A2(n12930), .ZN(n7587) );
  OR2_X1 U8499 ( .A1(n6772), .A2(n6771), .ZN(n6768) );
  NAND2_X1 U8500 ( .A1(n6770), .A2(n13856), .ZN(n6769) );
  AOI21_X1 U8501 ( .B1(n7583), .B2(n7586), .A(n12946), .ZN(n7582) );
  INV_X1 U8502 ( .A(n6569), .ZN(n7586) );
  NAND2_X1 U8503 ( .A1(n13867), .A2(n13866), .ZN(n7717) );
  OR2_X1 U8504 ( .A1(n13866), .A2(n13867), .ZN(n7718) );
  NAND2_X1 U8505 ( .A1(n7102), .A2(n6596), .ZN(n7101) );
  OAI21_X1 U8506 ( .B1(n12926), .B2(n13039), .A(n12919), .ZN(n7102) );
  INV_X1 U8507 ( .A(n7098), .ZN(n7097) );
  OAI21_X1 U8508 ( .B1(n12926), .B2(n12925), .A(n7099), .ZN(n7098) );
  INV_X1 U8509 ( .A(n7100), .ZN(n7099) );
  INV_X1 U8510 ( .A(n7582), .ZN(n7581) );
  INV_X1 U8511 ( .A(n12950), .ZN(n7579) );
  AOI21_X1 U8512 ( .B1(n7582), .B2(n7584), .A(n13416), .ZN(n7580) );
  AOI21_X1 U8513 ( .B1(n7084), .B2(n7080), .A(n6634), .ZN(n7079) );
  INV_X1 U8514 ( .A(n12952), .ZN(n7080) );
  INV_X1 U8515 ( .A(n12981), .ZN(n12974) );
  AOI21_X1 U8516 ( .B1(n13875), .B2(n13874), .A(n13873), .ZN(n13877) );
  OAI21_X1 U8517 ( .B1(n8404), .B2(n7460), .A(n7172), .ZN(n8426) );
  AND2_X1 U8518 ( .A1(n15241), .A2(n7651), .ZN(n7650) );
  AOI21_X1 U8519 ( .B1(n8437), .B2(n8439), .A(n6644), .ZN(n7651) );
  MUX2_X1 U8520 ( .A(n15140), .B(n15339), .S(n8779), .Z(n8547) );
  AOI21_X1 U8521 ( .B1(n6533), .B2(n7076), .A(n6660), .ZN(n7073) );
  INV_X1 U8522 ( .A(n7077), .ZN(n7076) );
  INV_X1 U8523 ( .A(n7093), .ZN(n7089) );
  INV_X1 U8524 ( .A(n8491), .ZN(n7639) );
  NAND2_X1 U8525 ( .A1(n8546), .A2(n7637), .ZN(n7636) );
  NOR2_X1 U8526 ( .A1(n8939), .A2(n8779), .ZN(n7637) );
  INV_X1 U8527 ( .A(n8581), .ZN(n7453) );
  NAND2_X1 U8528 ( .A1(n7085), .A2(n6592), .ZN(n7235) );
  OAI21_X1 U8529 ( .B1(n12980), .B2(n7087), .A(n7086), .ZN(n7085) );
  NOR2_X1 U8530 ( .A1(n7716), .A2(n13900), .ZN(n7714) );
  NAND2_X1 U8531 ( .A1(n13900), .A2(n7716), .ZN(n7713) );
  INV_X1 U8532 ( .A(n7452), .ZN(n7450) );
  AOI21_X1 U8533 ( .B1(n12742), .B2(n7947), .A(n9830), .ZN(n7946) );
  NOR2_X1 U8534 ( .A1(n12788), .A2(n7951), .ZN(n7947) );
  NOR2_X1 U8535 ( .A1(n7948), .A2(n7942), .ZN(n7941) );
  INV_X1 U8536 ( .A(n7533), .ZN(n7523) );
  NAND2_X1 U8537 ( .A1(n9640), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7533) );
  AND2_X1 U8538 ( .A1(n7066), .A2(n7900), .ZN(n7899) );
  NAND2_X1 U8539 ( .A1(n6535), .A2(n9517), .ZN(n7900) );
  INV_X1 U8540 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9236) );
  AOI22_X1 U8541 ( .A1(n13948), .A2(n13947), .B1(n13946), .B2(n13945), .ZN(
        n13953) );
  AND2_X1 U8542 ( .A1(n13964), .A2(n13998), .ZN(n7228) );
  INV_X1 U8543 ( .A(n13896), .ZN(n6782) );
  AOI21_X1 U8544 ( .B1(n7713), .B2(n7714), .A(n7712), .ZN(n7708) );
  NAND2_X1 U8545 ( .A1(n7713), .A2(n7712), .ZN(n7711) );
  INV_X1 U8546 ( .A(n7713), .ZN(n7709) );
  INV_X1 U8547 ( .A(n10302), .ZN(n13983) );
  INV_X1 U8548 ( .A(n14012), .ZN(n7346) );
  INV_X1 U8549 ( .A(n7979), .ZN(n7975) );
  INV_X1 U8550 ( .A(n14044), .ZN(n7902) );
  NAND2_X1 U8551 ( .A1(n8650), .A2(n8679), .ZN(n7024) );
  NAND2_X1 U8552 ( .A1(n7140), .A2(n10001), .ZN(n10005) );
  AND2_X1 U8553 ( .A1(n15122), .A2(n15153), .ZN(n7376) );
  OR4_X1 U8554 ( .A1(n15210), .A2(n8835), .A3(n8897), .A4(n15172), .ZN(n8836)
         );
  NOR2_X1 U8555 ( .A1(n6932), .A2(n6931), .ZN(n6930) );
  INV_X1 U8556 ( .A(n8512), .ZN(n8096) );
  INV_X1 U8557 ( .A(n8902), .ZN(n7551) );
  INV_X1 U8558 ( .A(n7831), .ZN(n7829) );
  NAND2_X1 U8559 ( .A1(n8530), .A2(n11067), .ZN(n7826) );
  AOI21_X1 U8560 ( .B1(n8174), .B2(n6630), .A(n7022), .ZN(n7021) );
  INV_X1 U8561 ( .A(n8175), .ZN(n7022) );
  NOR2_X1 U8562 ( .A1(n8518), .A2(n8163), .ZN(n8164) );
  INV_X1 U8563 ( .A(n8174), .ZN(n7023) );
  INV_X1 U8564 ( .A(n8149), .ZN(n6857) );
  AND2_X1 U8565 ( .A1(n8392), .A2(n8374), .ZN(n8147) );
  AND2_X1 U8566 ( .A1(n8138), .A2(n8135), .ZN(n7141) );
  OAI21_X1 U8567 ( .B1(n10878), .B2(n10886), .A(n7145), .ZN(n8140) );
  NAND2_X1 U8568 ( .A1(n10878), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7145) );
  NOR2_X1 U8569 ( .A1(n13300), .A2(n7061), .ZN(n7060) );
  NOR2_X1 U8570 ( .A1(n7063), .A2(n13334), .ZN(n7062) );
  INV_X1 U8571 ( .A(n13286), .ZN(n7067) );
  AND2_X1 U8572 ( .A1(n13013), .A2(n7770), .ZN(n7769) );
  NOR2_X1 U8573 ( .A1(n7771), .A2(n13006), .ZN(n7770) );
  NOR2_X1 U8574 ( .A1(n7767), .A2(n7238), .ZN(n7237) );
  NAND2_X1 U8575 ( .A1(n12866), .A2(n7768), .ZN(n7767) );
  NAND2_X1 U8576 ( .A1(n13013), .A2(n13014), .ZN(n7768) );
  OR2_X1 U8577 ( .A1(n9621), .A2(n11124), .ZN(n7530) );
  NOR2_X1 U8578 ( .A1(n9657), .A2(n12095), .ZN(n7354) );
  INV_X1 U8579 ( .A(n11897), .ZN(n7430) );
  INV_X1 U8580 ( .A(n12102), .ZN(n7429) );
  AND2_X1 U8581 ( .A1(n7430), .A2(n11743), .ZN(n7424) );
  NAND2_X1 U8582 ( .A1(n13090), .A2(n9676), .ZN(n9677) );
  NAND2_X1 U8583 ( .A1(n13132), .A2(n9631), .ZN(n9632) );
  INV_X1 U8584 ( .A(n12999), .ZN(n7923) );
  NOR2_X1 U8585 ( .A1(n9402), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7053) );
  INV_X1 U8586 ( .A(n12995), .ZN(n7872) );
  AND2_X1 U8587 ( .A1(n7869), .A2(n6836), .ZN(n6835) );
  NAND2_X1 U8588 ( .A1(n9524), .A2(n6841), .ZN(n6836) );
  INV_X1 U8589 ( .A(n9519), .ZN(n6841) );
  AND2_X1 U8590 ( .A1(n12303), .A2(n7050), .ZN(n7049) );
  INV_X1 U8591 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n7050) );
  INV_X1 U8592 ( .A(n9264), .ZN(n9251) );
  INV_X1 U8593 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n7042) );
  AND2_X1 U8594 ( .A1(n7045), .A2(n7044), .ZN(n7043) );
  INV_X1 U8595 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n7044) );
  INV_X1 U8596 ( .A(n12932), .ZN(n7868) );
  OAI21_X1 U8597 ( .B1(n12930), .B2(n7868), .A(n12937), .ZN(n7867) );
  INV_X1 U8598 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n9177) );
  INV_X1 U8599 ( .A(n9178), .ZN(n7389) );
  INV_X1 U8600 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n9127) );
  NAND2_X1 U8601 ( .A1(n13196), .A2(n13201), .ZN(n13013) );
  NAND2_X1 U8602 ( .A1(n12792), .A2(n13544), .ZN(n12981) );
  NAND2_X1 U8603 ( .A1(n7392), .A2(n7391), .ZN(n13305) );
  INV_X1 U8604 ( .A(n13319), .ZN(n7391) );
  NAND2_X1 U8605 ( .A1(n12981), .A2(n13299), .ZN(n7392) );
  NAND2_X1 U8606 ( .A1(n13379), .A2(n13367), .ZN(n9288) );
  OR2_X1 U8607 ( .A1(n13574), .A2(n12837), .ZN(n12959) );
  AND2_X1 U8608 ( .A1(n13568), .A2(n12765), .ZN(n12966) );
  NOR2_X1 U8609 ( .A1(n7165), .A2(n9185), .ZN(n7164) );
  INV_X1 U8610 ( .A(n9161), .ZN(n7165) );
  NOR2_X1 U8611 ( .A1(n9474), .A2(n7802), .ZN(n7801) );
  INV_X1 U8612 ( .A(n9459), .ZN(n7802) );
  INV_X1 U8613 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7149) );
  OAI21_X1 U8614 ( .B1(n7807), .B2(n7806), .A(n6718), .ZN(n7805) );
  INV_X1 U8615 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n7589) );
  NAND2_X1 U8616 ( .A1(n9275), .A2(n9290), .ZN(n7813) );
  NOR2_X1 U8617 ( .A1(n7780), .A2(n9163), .ZN(n6803) );
  AND2_X1 U8618 ( .A1(n8144), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9163) );
  OR2_X1 U8619 ( .A1(n9157), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n9166) );
  INV_X1 U8620 ( .A(n9154), .ZN(n7781) );
  NAND2_X1 U8621 ( .A1(n6789), .A2(n9082), .ZN(n6788) );
  INV_X1 U8622 ( .A(n6791), .ZN(n6789) );
  NOR2_X1 U8623 ( .A1(n10389), .A2(n11714), .ZN(n10800) );
  INV_X1 U8624 ( .A(n12666), .ZN(n7348) );
  INV_X1 U8625 ( .A(n7220), .ZN(n7218) );
  NOR2_X1 U8626 ( .A1(n10521), .A2(n10520), .ZN(n7326) );
  NOR2_X1 U8627 ( .A1(n13672), .A2(n10364), .ZN(n6978) );
  AOI21_X1 U8628 ( .B1(n7234), .B2(n12619), .A(n7233), .ZN(n7673) );
  INV_X1 U8629 ( .A(n12620), .ZN(n7233) );
  AOI21_X1 U8630 ( .B1(n12623), .B2(n12621), .A(n12622), .ZN(n12620) );
  OR3_X1 U8631 ( .A1(n12621), .A2(n12622), .A3(n12623), .ZN(n12628) );
  NAND2_X1 U8632 ( .A1(n7501), .A2(n7500), .ZN(n6899) );
  NAND2_X1 U8633 ( .A1(n14167), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7500) );
  AND2_X1 U8634 ( .A1(n6899), .A2(n14170), .ZN(n14165) );
  AND2_X1 U8635 ( .A1(n10627), .A2(n10626), .ZN(n10630) );
  NOR2_X1 U8636 ( .A1(n14522), .A2(n14528), .ZN(n7653) );
  NOR2_X1 U8637 ( .A1(n6909), .A2(n14051), .ZN(n6908) );
  NAND2_X1 U8638 ( .A1(n10614), .A2(n6913), .ZN(n6912) );
  INV_X1 U8639 ( .A(n10613), .ZN(n6913) );
  OR2_X1 U8640 ( .A1(n14404), .A2(n14405), .ZN(n8074) );
  INV_X1 U8641 ( .A(n14394), .ZN(n7280) );
  NAND2_X1 U8642 ( .A1(n10362), .A2(n6554), .ZN(n10475) );
  NAND2_X1 U8643 ( .A1(n10362), .A2(n6967), .ZN(n10466) );
  NAND2_X1 U8644 ( .A1(n10362), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n10457) );
  INV_X1 U8645 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10437) );
  OR2_X1 U8646 ( .A1(n10438), .A2(n10437), .ZN(n10447) );
  INV_X1 U8647 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10430) );
  OR2_X1 U8648 ( .A1(n10431), .A2(n10430), .ZN(n10438) );
  NAND2_X1 U8649 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n10404) );
  NAND2_X1 U8650 ( .A1(n7635), .A2(n11253), .ZN(n7692) );
  AND2_X1 U8651 ( .A1(n14058), .A2(n8002), .ZN(n8001) );
  NAND2_X1 U8652 ( .A1(n14283), .A2(n14273), .ZN(n14251) );
  NAND2_X1 U8653 ( .A1(n7664), .A2(n7660), .ZN(n14362) );
  NOR2_X1 U8654 ( .A1(n14413), .A2(n14580), .ZN(n14414) );
  NOR2_X1 U8655 ( .A1(n14767), .A2(n14695), .ZN(n6928) );
  NOR2_X1 U8656 ( .A1(n7463), .A2(n8642), .ZN(n7461) );
  INV_X1 U8657 ( .A(n8672), .ZN(n7468) );
  AND2_X1 U8658 ( .A1(n15269), .A2(n8779), .ZN(n8856) );
  AND2_X1 U8659 ( .A1(n6565), .A2(n8855), .ZN(n8850) );
  NAND2_X1 U8660 ( .A1(n8096), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8538) );
  AND2_X1 U8661 ( .A1(n6848), .A2(n6846), .ZN(n15045) );
  NOR2_X1 U8662 ( .A1(n6588), .A2(n8953), .ZN(n6846) );
  NOR2_X1 U8663 ( .A1(n10073), .A2(n7861), .ZN(n7859) );
  OAI21_X1 U8664 ( .B1(n8064), .B2(n8946), .A(n6646), .ZN(n8063) );
  NAND2_X1 U8665 ( .A1(n8097), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8583) );
  NAND2_X1 U8666 ( .A1(n8096), .A2(n6930), .ZN(n8540) );
  INV_X1 U8667 ( .A(n8892), .ZN(n8030) );
  NOR2_X1 U8668 ( .A1(n7483), .A2(n7482), .ZN(n7481) );
  NAND2_X1 U8669 ( .A1(n8929), .A2(n11673), .ZN(n7482) );
  INV_X1 U8670 ( .A(n7486), .ZN(n7483) );
  NAND2_X1 U8671 ( .A1(n6927), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n8312) );
  NAND2_X1 U8672 ( .A1(n11348), .A2(n11472), .ZN(n8919) );
  NAND2_X1 U8673 ( .A1(n15535), .A2(n8262), .ZN(n8875) );
  AND2_X1 U8674 ( .A1(n15094), .A2(n15095), .ZN(n15115) );
  NAND2_X1 U8675 ( .A1(n15180), .A2(n15159), .ZN(n15161) );
  AND2_X1 U8676 ( .A1(n11828), .A2(n15163), .ZN(n8974) );
  NAND2_X1 U8677 ( .A1(n8016), .A2(n8015), .ZN(n8014) );
  NAND2_X1 U8678 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n8017), .ZN(n8016) );
  NAND2_X1 U8679 ( .A1(n15422), .A2(n8020), .ZN(n8015) );
  NAND2_X1 U8680 ( .A1(n8020), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n8017) );
  NAND2_X1 U8681 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(n7658), .ZN(n8019) );
  NOR2_X1 U8682 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(n15422), .ZN(n8018) );
  AOI21_X1 U8683 ( .B1(n8184), .B2(n6990), .A(n6989), .ZN(n6988) );
  INV_X1 U8684 ( .A(n8184), .ZN(n6991) );
  INV_X1 U8685 ( .A(n8185), .ZN(n6989) );
  NAND2_X1 U8686 ( .A1(n6517), .A2(n6523), .ZN(n8792) );
  AOI21_X1 U8687 ( .B1(n7021), .B2(n7023), .A(n7824), .ZN(n7020) );
  INV_X1 U8688 ( .A(n7826), .ZN(n7825) );
  NOR2_X1 U8689 ( .A1(n8470), .A2(n8169), .ZN(n8517) );
  NOR2_X1 U8690 ( .A1(n8168), .A2(n11044), .ZN(n8169) );
  NOR2_X1 U8691 ( .A1(n8468), .A2(SI_14_), .ZN(n8518) );
  OR2_X1 U8692 ( .A1(n8377), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n8415) );
  XNOR2_X1 U8693 ( .A(n8140), .B(n10857), .ZN(n8139) );
  INV_X1 U8694 ( .A(n8215), .ZN(n7146) );
  INV_X1 U8695 ( .A(P2_RD_REG_SCAN_IN), .ZN(n6982) );
  NAND2_X1 U8696 ( .A1(n6810), .A2(n6809), .ZN(n9696) );
  NAND2_X1 U8697 ( .A1(n6573), .A2(n9720), .ZN(n6809) );
  NAND3_X1 U8698 ( .A1(n7336), .A2(n7335), .A3(n6573), .ZN(n6810) );
  INV_X1 U8699 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n12335) );
  INV_X1 U8700 ( .A(n7569), .ZN(n9698) );
  AND2_X1 U8701 ( .A1(n6811), .A2(n6668), .ZN(n9706) );
  OR2_X1 U8702 ( .A1(n9718), .A2(n14916), .ZN(n6811) );
  XNOR2_X1 U8703 ( .A(n9706), .B(n7570), .ZN(n9740) );
  INV_X1 U8704 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n7570) );
  NAND2_X1 U8705 ( .A1(n6814), .A2(n6812), .ZN(n9709) );
  NAND2_X1 U8706 ( .A1(P3_ADDR_REG_9__SCAN_IN), .A2(n6813), .ZN(n6812) );
  NAND2_X1 U8707 ( .A1(n9716), .A2(n9717), .ZN(n6814) );
  OAI22_X1 U8708 ( .A1(n9762), .A2(n9713), .B1(P3_ADDR_REG_16__SCAN_IN), .B2(
        n9760), .ZN(n9763) );
  NAND2_X1 U8709 ( .A1(n12750), .A2(n9840), .ZN(n6936) );
  INV_X1 U8710 ( .A(n7929), .ZN(n6950) );
  AND2_X1 U8711 ( .A1(n12751), .A2(n9843), .ZN(n9844) );
  INV_X1 U8712 ( .A(n7053), .ZN(n9416) );
  NOR2_X1 U8713 ( .A1(n9795), .A2(n11958), .ZN(n9796) );
  NAND2_X1 U8714 ( .A1(n6953), .A2(n6952), .ZN(n6951) );
  INV_X1 U8715 ( .A(n11767), .ZN(n6953) );
  NAND2_X1 U8716 ( .A1(n6941), .A2(n9803), .ZN(n11854) );
  INV_X1 U8717 ( .A(n11819), .ZN(n6941) );
  NAND2_X1 U8718 ( .A1(n6939), .A2(n6610), .ZN(n12241) );
  NAND2_X1 U8719 ( .A1(n7961), .A2(n11820), .ZN(n6940) );
  NAND2_X1 U8720 ( .A1(n11855), .A2(n9808), .ZN(n12527) );
  INV_X1 U8721 ( .A(n12771), .ZN(n7931) );
  OR2_X1 U8722 ( .A1(n13024), .A2(n9573), .ZN(n9854) );
  AOI21_X1 U8723 ( .B1(n10848), .B2(n9615), .A(n9616), .ZN(n11033) );
  AOI21_X1 U8724 ( .B1(n10848), .B2(n9585), .A(n9586), .ZN(n7121) );
  NAND2_X1 U8725 ( .A1(n7121), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n11032) );
  NAND2_X1 U8726 ( .A1(n7394), .A2(n7399), .ZN(n9635) );
  NAND2_X1 U8727 ( .A1(n7403), .A2(n6615), .ZN(n7399) );
  NAND2_X1 U8728 ( .A1(n13612), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7394) );
  XNOR2_X1 U8729 ( .A(n11145), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n11133) );
  XNOR2_X1 U8730 ( .A(n9621), .B(n11124), .ZN(n11118) );
  INV_X1 U8731 ( .A(n7525), .ZN(n7520) );
  NAND2_X1 U8732 ( .A1(n11118), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7531) );
  AND2_X1 U8733 ( .A1(n11179), .A2(n7625), .ZN(n11198) );
  NAND2_X1 U8734 ( .A1(n7445), .A2(n9654), .ZN(n11555) );
  AOI21_X1 U8735 ( .B1(n7433), .B2(n7439), .A(n9655), .ZN(n7431) );
  NAND2_X1 U8736 ( .A1(n11552), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7509) );
  OAI21_X1 U8737 ( .B1(n11745), .B2(n11744), .A(n11743), .ZN(n11899) );
  NAND2_X1 U8738 ( .A1(n7426), .A2(n7430), .ZN(n7425) );
  INV_X1 U8739 ( .A(n7427), .ZN(n7426) );
  AOI21_X1 U8740 ( .B1(n11743), .B2(n11744), .A(n7428), .ZN(n7427) );
  INV_X1 U8741 ( .A(n11898), .ZN(n7428) );
  NAND2_X1 U8742 ( .A1(n7244), .A2(n12106), .ZN(n7243) );
  INV_X1 U8743 ( .A(n7383), .ZN(n7244) );
  NAND2_X1 U8744 ( .A1(n11745), .A2(n7424), .ZN(n7423) );
  NAND2_X1 U8745 ( .A1(n12107), .A2(n9626), .ZN(n13054) );
  NAND2_X1 U8746 ( .A1(n7409), .A2(n7408), .ZN(n7407) );
  INV_X1 U8747 ( .A(n13070), .ZN(n7408) );
  INV_X1 U8748 ( .A(n13069), .ZN(n7409) );
  NAND2_X1 U8749 ( .A1(n7406), .A2(n7405), .ZN(n13090) );
  NOR2_X1 U8750 ( .A1(n13087), .A2(n13088), .ZN(n7405) );
  AND2_X1 U8751 ( .A1(n13151), .A2(n6716), .ZN(n7626) );
  OAI21_X1 U8752 ( .B1(n6586), .B2(n7417), .A(n7410), .ZN(n13161) );
  NOR2_X1 U8753 ( .A1(n7412), .A2(n7417), .ZN(n7411) );
  NOR2_X1 U8754 ( .A1(n7418), .A2(n13151), .ZN(n7417) );
  AND2_X1 U8755 ( .A1(n9472), .A2(n9471), .ZN(n12823) );
  INV_X1 U8756 ( .A(n12890), .ZN(n13193) );
  AND2_X1 U8757 ( .A1(n13012), .A2(n13005), .ZN(n13215) );
  NAND2_X1 U8758 ( .A1(n13217), .A2(n13420), .ZN(n13220) );
  NAND2_X1 U8759 ( .A1(n7053), .A2(n12783), .ZN(n9432) );
  INV_X1 U8760 ( .A(n13251), .ZN(n13245) );
  NAND2_X1 U8761 ( .A1(n6794), .A2(n7152), .ZN(n13246) );
  AOI21_X1 U8762 ( .B1(n7154), .B2(n7153), .A(n6647), .ZN(n7152) );
  NAND2_X1 U8763 ( .A1(n13246), .A2(n13245), .ZN(n13244) );
  OR2_X1 U8764 ( .A1(n9389), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9402) );
  NAND2_X1 U8765 ( .A1(n9341), .A2(n7047), .ZN(n9389) );
  AND2_X1 U8766 ( .A1(n7049), .A2(n7048), .ZN(n7047) );
  INV_X1 U8767 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n7048) );
  NAND2_X1 U8768 ( .A1(n9341), .A2(n7049), .ZN(n9378) );
  NAND2_X1 U8769 ( .A1(n9251), .A2(n9250), .ZN(n9266) );
  NAND2_X1 U8770 ( .A1(n6591), .A2(n9225), .ZN(n9264) );
  INV_X1 U8771 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n9225) );
  NAND2_X1 U8772 ( .A1(n7389), .A2(n7045), .ZN(n9210) );
  NAND2_X1 U8773 ( .A1(n7389), .A2(n9177), .ZN(n9194) );
  NAND2_X1 U8774 ( .A1(n7052), .A2(n7051), .ZN(n9178) );
  AND2_X1 U8775 ( .A1(n9127), .A2(n7390), .ZN(n7051) );
  NOR2_X1 U8776 ( .A1(n12884), .A2(n6820), .ZN(n6816) );
  NAND2_X1 U8777 ( .A1(n7052), .A2(n9127), .ZN(n9147) );
  NAND2_X1 U8778 ( .A1(n7249), .A2(n7248), .ZN(n9128) );
  INV_X1 U8779 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n7248) );
  NAND3_X1 U8780 ( .A1(n9075), .A2(n9074), .A3(n9086), .ZN(n9109) );
  INV_X1 U8781 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9086) );
  NOR2_X1 U8782 ( .A1(n15901), .A2(n9852), .ZN(n11106) );
  NAND2_X1 U8783 ( .A1(n15851), .A2(n12876), .ZN(n6823) );
  INV_X1 U8784 ( .A(n9055), .ZN(n11668) );
  NAND2_X1 U8785 ( .A1(n15918), .A2(n13401), .ZN(n7598) );
  NAND2_X1 U8786 ( .A1(n10700), .A2(n12823), .ZN(n13192) );
  NAND2_X1 U8787 ( .A1(n9429), .A2(n9428), .ZN(n13443) );
  AND2_X1 U8788 ( .A1(n12983), .A2(n12984), .ZN(n13307) );
  INV_X1 U8789 ( .A(n7392), .ZN(n13318) );
  AND2_X1 U8790 ( .A1(n12959), .A2(n12958), .ZN(n13369) );
  NAND2_X1 U8791 ( .A1(n9263), .A2(n9262), .ZN(n12896) );
  INV_X1 U8792 ( .A(n12955), .ZN(n13391) );
  AND2_X1 U8793 ( .A1(n7873), .A2(n6830), .ZN(n6829) );
  NAND2_X1 U8794 ( .A1(n7875), .A2(n12944), .ZN(n6830) );
  NAND2_X1 U8795 ( .A1(n7324), .A2(n9146), .ZN(n12092) );
  INV_X1 U8796 ( .A(n9852), .ZN(n10683) );
  OAI22_X1 U8797 ( .A1(n12706), .A2(n12553), .B1(P2_DATAO_REG_29__SCAN_IN), 
        .B2(n12697), .ZN(n12850) );
  NAND2_X1 U8798 ( .A1(n9443), .A2(n9442), .ZN(n9458) );
  OAI21_X1 U8799 ( .B1(n9426), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n9425), .ZN(
        n9441) );
  XNOR2_X1 U8800 ( .A(n9576), .B(n9575), .ZN(n9855) );
  INV_X1 U8801 ( .A(n7792), .ZN(n7791) );
  AOI21_X1 U8802 ( .B1(n7790), .B2(n7792), .A(n7789), .ZN(n7788) );
  INV_X1 U8803 ( .A(n9318), .ZN(n7789) );
  AND2_X1 U8804 ( .A1(n9320), .A2(n9319), .ZN(n9331) );
  NAND2_X1 U8805 ( .A1(n9238), .A2(n9237), .ZN(n9277) );
  OR2_X1 U8806 ( .A1(n9220), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n9157) );
  AND2_X1 U8807 ( .A1(n12617), .A2(n12619), .ZN(n13637) );
  NAND2_X1 U8808 ( .A1(n13634), .A2(n12618), .ZN(n13635) );
  OR2_X1 U8809 ( .A1(n7683), .A2(n7682), .ZN(n7267) );
  NOR2_X1 U8810 ( .A1(n7686), .A2(n7682), .ZN(n7681) );
  INV_X1 U8811 ( .A(n7326), .ZN(n10523) );
  NAND2_X1 U8812 ( .A1(n7326), .A2(n6978), .ZN(n10538) );
  XNOR2_X1 U8813 ( .A(n14539), .B(n12669), .ZN(n12648) );
  AOI21_X1 U8814 ( .B1(n7224), .B2(n12235), .A(n7223), .ZN(n7222) );
  INV_X1 U8815 ( .A(n12600), .ZN(n7223) );
  NAND2_X1 U8816 ( .A1(n10363), .A2(n6555), .ZN(n10509) );
  NOR2_X1 U8817 ( .A1(n13715), .A2(n13714), .ZN(n13713) );
  XNOR2_X1 U8818 ( .A(n7205), .B(n12669), .ZN(n12586) );
  XNOR2_X1 U8819 ( .A(n14329), .B(n11713), .ZN(n13726) );
  NAND2_X1 U8820 ( .A1(n12126), .A2(n12125), .ZN(n12232) );
  NAND2_X1 U8821 ( .A1(n13707), .A2(n13708), .ZN(n13706) );
  NAND2_X1 U8822 ( .A1(n13635), .A2(n12619), .ZN(n13698) );
  AND3_X1 U8823 ( .A1(n7699), .A2(n14003), .A3(n14004), .ZN(n7698) );
  AOI21_X1 U8824 ( .B1(n13905), .B2(n13906), .A(n6764), .ZN(n6763) );
  OAI21_X1 U8825 ( .B1(n13905), .B2(n13906), .A(n7701), .ZN(n6762) );
  XNOR2_X1 U8826 ( .A(n14025), .B(n14085), .ZN(n14028) );
  NOR2_X1 U8827 ( .A1(n14496), .A2(n7837), .ZN(n7836) );
  NAND2_X1 U8828 ( .A1(n6534), .A2(n8000), .ZN(n7837) );
  AOI21_X1 U8829 ( .B1(n14209), .B2(n10720), .A(n10583), .ZN(n13993) );
  INV_X1 U8830 ( .A(n10389), .ZN(n11275) );
  NAND4_X1 U8831 ( .A1(n10378), .A2(n10377), .A3(n10375), .A4(n10376), .ZN(
        n10586) );
  OR2_X1 U8832 ( .A1(n7879), .A2(n7270), .ZN(n10378) );
  NAND2_X1 U8833 ( .A1(n13969), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10375) );
  OR2_X1 U8834 ( .A1(n15670), .A2(n15669), .ZN(n15672) );
  NAND2_X1 U8835 ( .A1(n15667), .A2(n6890), .ZN(n6891) );
  NOR2_X1 U8836 ( .A1(n15687), .A2(n6893), .ZN(n6890) );
  OR2_X1 U8837 ( .A1(n15683), .A2(n15684), .ZN(n15680) );
  AND2_X1 U8838 ( .A1(n11241), .A2(n11240), .ZN(n11244) );
  OR2_X1 U8839 ( .A1(n11235), .A2(n11236), .ZN(n11646) );
  NOR2_X1 U8840 ( .A1(n6527), .A2(n11265), .ZN(n11641) );
  AND2_X1 U8841 ( .A1(n15694), .A2(n11647), .ZN(n11650) );
  NAND2_X1 U8842 ( .A1(n6552), .A2(n7499), .ZN(n6895) );
  NAND2_X1 U8843 ( .A1(n15709), .A2(n6552), .ZN(n6894) );
  AND2_X1 U8844 ( .A1(n15718), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n15716) );
  NOR2_X1 U8845 ( .A1(n14165), .A2(n6898), .ZN(n15746) );
  NOR2_X1 U8846 ( .A1(n6899), .A2(n14170), .ZN(n6898) );
  NOR2_X1 U8847 ( .A1(n7645), .A2(n14025), .ZN(n7642) );
  AND2_X1 U8848 ( .A1(n7645), .A2(n14025), .ZN(n7643) );
  AND2_X1 U8849 ( .A1(n10640), .A2(n10716), .ZN(n14203) );
  INV_X1 U8850 ( .A(n8005), .ZN(n8004) );
  OAI21_X1 U8851 ( .B1(n14222), .B2(n8007), .A(n8006), .ZN(n8005) );
  NAND2_X1 U8852 ( .A1(n14217), .A2(n14088), .ZN(n8006) );
  NOR2_X1 U8853 ( .A1(n14222), .A2(n8003), .ZN(n8002) );
  INV_X1 U8854 ( .A(n10571), .ZN(n8003) );
  NAND2_X1 U8855 ( .A1(n14283), .A2(n7653), .ZN(n14252) );
  NOR2_X1 U8856 ( .A1(n7913), .A2(n6542), .ZN(n6915) );
  INV_X1 U8857 ( .A(n7325), .ZN(n10546) );
  AOI21_X1 U8858 ( .B1(n7109), .B2(n6608), .A(n7106), .ZN(n14310) );
  NAND2_X1 U8859 ( .A1(n7107), .A2(n6642), .ZN(n7106) );
  NAND2_X1 U8860 ( .A1(n14310), .A2(n14309), .ZN(n14308) );
  NOR2_X1 U8861 ( .A1(n14390), .A2(n6525), .ZN(n14348) );
  NAND2_X1 U8862 ( .A1(n14348), .A2(n14632), .ZN(n14325) );
  XNOR2_X1 U8863 ( .A(n14351), .B(n14092), .ZN(n14338) );
  INV_X1 U8864 ( .A(n7884), .ZN(n7883) );
  OAI21_X1 U8865 ( .B1(n7889), .B2(n7885), .A(n10612), .ZN(n7884) );
  NAND2_X1 U8866 ( .A1(n10363), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n10496) );
  NAND2_X1 U8867 ( .A1(n10363), .A2(n6970), .ZN(n10500) );
  NAND2_X1 U8868 ( .A1(n7664), .A2(n7663), .ZN(n14377) );
  NAND2_X1 U8869 ( .A1(n7114), .A2(n7280), .ZN(n14385) );
  INV_X1 U8870 ( .A(n14387), .ZN(n7114) );
  OR2_X1 U8871 ( .A1(n10475), .A2(n13741), .ZN(n10483) );
  INV_X1 U8872 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10482) );
  OR2_X1 U8873 ( .A1(n10483), .A2(n10482), .ZN(n10491) );
  OR2_X1 U8874 ( .A1(n14443), .A2(n14442), .ZN(n14445) );
  INV_X1 U8875 ( .A(n10597), .ZN(n14046) );
  OR2_X1 U8876 ( .A1(n12054), .A2(n7654), .ZN(n12083) );
  INV_X1 U8877 ( .A(n7656), .ZN(n7654) );
  NAND2_X1 U8878 ( .A1(n10429), .A2(n10428), .ZN(n12049) );
  NAND2_X1 U8879 ( .A1(n7657), .A2(n10221), .ZN(n12081) );
  INV_X1 U8880 ( .A(n12054), .ZN(n7657) );
  OAI21_X1 U8881 ( .B1(n10592), .B2(n6562), .A(n7904), .ZN(n12048) );
  NAND2_X1 U8882 ( .A1(n10216), .A2(n10215), .ZN(n13858) );
  NAND2_X1 U8883 ( .A1(n10361), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10414) );
  NAND2_X1 U8884 ( .A1(n10361), .A2(n6532), .ZN(n10422) );
  NAND2_X1 U8885 ( .A1(n11966), .A2(n11965), .ZN(n10588) );
  INV_X1 U8886 ( .A(n10184), .ZN(n7635) );
  CLKBUF_X1 U8887 ( .A(n10188), .Z(n10301) );
  AND2_X1 U8888 ( .A1(n6916), .A2(n6919), .ZN(n14266) );
  NAND2_X1 U8889 ( .A1(n7117), .A2(n7115), .ZN(n10344) );
  NAND2_X1 U8890 ( .A1(n10337), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10303) );
  NAND2_X1 U8891 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n10306), .ZN(n10307) );
  NOR2_X1 U8892 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n7727) );
  NAND2_X1 U8893 ( .A1(n6761), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6760) );
  NAND2_X1 U8894 ( .A1(n10173), .A2(n10160), .ZN(n6761) );
  OR2_X1 U8895 ( .A1(n10203), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n10208) );
  INV_X1 U8896 ( .A(n10182), .ZN(n10190) );
  INV_X1 U8897 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n10178) );
  NAND2_X1 U8898 ( .A1(n6927), .A2(n6637), .ZN(n8335) );
  NAND2_X1 U8899 ( .A1(n7749), .A2(n9942), .ZN(n7748) );
  AND2_X1 U8900 ( .A1(n10115), .A2(n10114), .ZN(n10130) );
  NAND2_X1 U8901 ( .A1(n9889), .A2(n10123), .ZN(n9890) );
  NAND2_X1 U8902 ( .A1(n8097), .A2(n6933), .ZN(n8598) );
  NOR2_X1 U8903 ( .A1(n7139), .A2(n7755), .ZN(n7754) );
  NOR2_X1 U8904 ( .A1(n10010), .A2(n14824), .ZN(n7755) );
  OAI21_X1 U8905 ( .B1(n14744), .B2(n10018), .A(n6587), .ZN(n10019) );
  NAND2_X1 U8906 ( .A1(n7752), .A2(n10020), .ZN(n14755) );
  INV_X1 U8907 ( .A(n10019), .ZN(n10020) );
  NAND2_X1 U8908 ( .A1(n7756), .A2(n7754), .ZN(n7752) );
  NAND2_X1 U8909 ( .A1(n8098), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U8910 ( .A1(n10086), .A2(n10087), .ZN(n7743) );
  NAND2_X1 U8911 ( .A1(n11862), .A2(n9958), .ZN(n12174) );
  XNOR2_X1 U8912 ( .A(n9995), .B(n10123), .ZN(n14677) );
  NAND2_X1 U8913 ( .A1(n7147), .A2(n9994), .ZN(n9995) );
  NAND2_X1 U8914 ( .A1(n14724), .A2(n9886), .ZN(n7147) );
  NAND2_X1 U8915 ( .A1(n6862), .A2(n10058), .ZN(n6861) );
  INV_X1 U8916 ( .A(n14792), .ZN(n6862) );
  NAND2_X1 U8917 ( .A1(n14718), .A2(n14717), .ZN(n14794) );
  NAND2_X1 U8918 ( .A1(n8097), .A2(n6557), .ZN(n8618) );
  OR2_X1 U8919 ( .A1(n8618), .A2(n14798), .ZN(n8630) );
  INV_X1 U8920 ( .A(n9958), .ZN(n7765) );
  OAI22_X1 U8921 ( .A1(n15535), .A2(n10059), .B1(n9953), .B2(n8262), .ZN(n7001) );
  OR2_X1 U8922 ( .A1(n14804), .A2(n14803), .ZN(n7761) );
  INV_X1 U8923 ( .A(n6999), .ZN(n6996) );
  OAI21_X1 U8924 ( .B1(n9932), .B2(n6998), .A(n6997), .ZN(n6993) );
  OR2_X1 U8925 ( .A1(n11354), .A2(n11353), .ZN(n6997) );
  INV_X1 U8926 ( .A(n10097), .ZN(n7740) );
  INV_X1 U8927 ( .A(n8820), .ZN(n10758) );
  INV_X1 U8928 ( .A(n7756), .ZN(n7753) );
  NAND2_X1 U8929 ( .A1(n6925), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8479) );
  INV_X1 U8930 ( .A(n8455), .ZN(n6925) );
  INV_X1 U8931 ( .A(n15255), .ZN(n15213) );
  AND2_X1 U8932 ( .A1(n7191), .A2(n7258), .ZN(n7190) );
  NAND2_X1 U8933 ( .A1(n7194), .A2(n7193), .ZN(n7191) );
  NOR2_X1 U8934 ( .A1(n7374), .A2(n8841), .ZN(n7373) );
  AND3_X1 U8935 ( .A1(n8728), .A2(n8727), .A3(n8726), .ZN(n14973) );
  AND4_X1 U8936 ( .A1(n8460), .A2(n8459), .A3(n8458), .A4(n8457), .ZN(n15226)
         );
  AND2_X1 U8937 ( .A1(n8289), .A2(n8291), .ZN(n8041) );
  NAND2_X1 U8938 ( .A1(n6514), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8292) );
  OR2_X1 U8939 ( .A1(n10920), .A2(n10921), .ZN(n10918) );
  OR2_X1 U8940 ( .A1(n10935), .A2(n10936), .ZN(n10933) );
  INV_X1 U8941 ( .A(n11164), .ZN(n7337) );
  INV_X1 U8942 ( .A(n11163), .ZN(n7338) );
  OR2_X1 U8943 ( .A1(n11311), .A2(n11310), .ZN(n11313) );
  OR2_X1 U8944 ( .A1(n11599), .A2(n11600), .ZN(n11597) );
  AND2_X1 U8945 ( .A1(n11593), .A2(n10743), .ZN(n11619) );
  OR2_X1 U8946 ( .A1(n12216), .A2(n12217), .ZN(n12213) );
  OR2_X1 U8947 ( .A1(n12221), .A2(n12222), .ZN(n12218) );
  NAND2_X1 U8948 ( .A1(n8760), .A2(n8759), .ZN(n15003) );
  INV_X1 U8949 ( .A(n14996), .ZN(n14993) );
  AOI21_X1 U8950 ( .B1(n8057), .B2(n8054), .A(n8053), .ZN(n8052) );
  NOR2_X1 U8951 ( .A1(n7840), .A2(n14837), .ZN(n8053) );
  NAND2_X1 U8952 ( .A1(n15005), .A2(n8100), .ZN(n10668) );
  NAND2_X1 U8953 ( .A1(n15029), .A2(n15020), .ZN(n15015) );
  AND2_X1 U8954 ( .A1(n8684), .A2(n8683), .ZN(n15018) );
  AND2_X1 U8955 ( .A1(n15113), .A2(n7860), .ZN(n15079) );
  NAND2_X1 U8956 ( .A1(n7859), .A2(n15113), .ZN(n15066) );
  NAND2_X1 U8957 ( .A1(n7540), .A2(n7542), .ZN(n7537) );
  AND2_X1 U8958 ( .A1(n6851), .A2(n6850), .ZN(n15081) );
  INV_X1 U8959 ( .A(n8063), .ZN(n6851) );
  AND2_X1 U8960 ( .A1(n15113), .A2(n15107), .ZN(n15102) );
  INV_X1 U8961 ( .A(n14840), .ZN(n15099) );
  NAND2_X1 U8962 ( .A1(n7848), .A2(n7849), .ZN(n15137) );
  NOR2_X1 U8963 ( .A1(n15339), .A2(n15330), .ZN(n7848) );
  INV_X1 U8964 ( .A(n7852), .ZN(n7849) );
  NAND2_X1 U8965 ( .A1(n15193), .A2(n8968), .ZN(n15194) );
  INV_X1 U8966 ( .A(n8940), .ZN(n15150) );
  NOR2_X1 U8967 ( .A1(n7477), .A2(n7476), .ZN(n8937) );
  INV_X1 U8968 ( .A(n8933), .ZN(n7476) );
  INV_X1 U8969 ( .A(n15224), .ZN(n7477) );
  INV_X1 U8970 ( .A(n8897), .ZN(n15241) );
  NAND2_X1 U8971 ( .A1(n15222), .A2(n15241), .ZN(n15224) );
  NOR2_X1 U8972 ( .A1(n14724), .A2(n7842), .ZN(n15252) );
  NOR2_X1 U8973 ( .A1(n14724), .A2(n6702), .ZN(n15251) );
  NAND2_X1 U8974 ( .A1(n8095), .A2(n8094), .ZN(n8428) );
  INV_X1 U8975 ( .A(n8407), .ZN(n8095) );
  OR2_X1 U8976 ( .A1(n8428), .A2(n12346), .ZN(n8453) );
  NAND2_X1 U8977 ( .A1(n8031), .A2(n8892), .ZN(n12188) );
  NAND2_X1 U8978 ( .A1(n12000), .A2(n8891), .ZN(n8031) );
  AND4_X1 U8979 ( .A1(n8412), .A2(n8411), .A3(n8410), .A4(n8409), .ZN(n14729)
         );
  AND4_X1 U8980 ( .A1(n8373), .A2(n8372), .A3(n8371), .A4(n8370), .ZN(n12183)
         );
  INV_X1 U8981 ( .A(n8022), .ZN(n8021) );
  OAI21_X1 U8982 ( .B1(n8026), .B2(n11581), .A(n11673), .ZN(n8022) );
  NOR2_X1 U8983 ( .A1(n15396), .A2(n7854), .ZN(n7853) );
  INV_X1 U8984 ( .A(n7856), .ZN(n7854) );
  NAND2_X1 U8985 ( .A1(n11571), .A2(n15570), .ZN(n11587) );
  AND4_X1 U8986 ( .A1(n8341), .A2(n8340), .A3(n8339), .A4(n8338), .ZN(n11677)
         );
  NAND2_X1 U8987 ( .A1(n11386), .A2(n8920), .ZN(n11488) );
  NAND2_X1 U8988 ( .A1(n7839), .A2(n15502), .ZN(n11391) );
  INV_X1 U8989 ( .A(n11504), .ZN(n7839) );
  NAND2_X1 U8990 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n8228) );
  NAND2_X1 U8991 ( .A1(n7470), .A2(n8918), .ZN(n11073) );
  NAND2_X1 U8992 ( .A1(n11505), .A2(n8299), .ZN(n11504) );
  AND2_X1 U8993 ( .A1(n15535), .A2(n9892), .ZN(n7632) );
  CLKBUF_X1 U8994 ( .A(n8874), .Z(n11439) );
  XNOR2_X1 U8995 ( .A(n15536), .B(n9892), .ZN(n11440) );
  AND2_X1 U8996 ( .A1(n8032), .A2(n8033), .ZN(n15124) );
  NAND2_X1 U8997 ( .A1(n8537), .A2(n8536), .ZN(n15342) );
  NAND2_X1 U8998 ( .A1(n8062), .A2(n8924), .ZN(n11582) );
  INV_X1 U8999 ( .A(n15580), .ZN(n15569) );
  AOI21_X1 U9000 ( .B1(n8721), .B2(n8091), .A(n8720), .ZN(n8722) );
  NAND2_X1 U9001 ( .A1(n8735), .A2(n8734), .ZN(n8739) );
  XNOR2_X1 U9002 ( .A(n8200), .B(n8199), .ZN(n8821) );
  NAND2_X1 U9003 ( .A1(n7259), .A2(n8704), .ZN(n8774) );
  XNOR2_X1 U9004 ( .A(n8702), .B(n8198), .ZN(n14668) );
  XNOR2_X1 U9005 ( .A(n8669), .B(n8668), .ZN(n12547) );
  NAND2_X1 U9006 ( .A1(n8816), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8208) );
  XNOR2_X1 U9007 ( .A(n8610), .B(n8605), .ZN(n11827) );
  NAND2_X1 U9008 ( .A1(n6867), .A2(n6869), .ZN(n8472) );
  NAND2_X1 U9009 ( .A1(n6868), .A2(n8168), .ZN(n6867) );
  NAND2_X1 U9010 ( .A1(n6858), .A2(n8149), .ZN(n8413) );
  OR2_X1 U9011 ( .A1(n8348), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n8377) );
  INV_X1 U9012 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8217) );
  OR2_X1 U9013 ( .A1(n8271), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n8236) );
  INV_X1 U9014 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n11405) );
  XNOR2_X1 U9015 ( .A(n9696), .B(n12335), .ZN(n9719) );
  NAND2_X1 U9016 ( .A1(n15921), .A2(n9733), .ZN(n9736) );
  NAND2_X1 U9017 ( .A1(n6749), .A2(n6622), .ZN(n6750) );
  INV_X1 U9018 ( .A(n7560), .ZN(n9714) );
  OAI21_X1 U9019 ( .B1(n9748), .B2(n9749), .A(n6717), .ZN(n7560) );
  AOI21_X1 U9020 ( .B1(n9751), .B2(n9712), .A(n6725), .ZN(n9754) );
  INV_X1 U9021 ( .A(n7732), .ZN(n7731) );
  NAND2_X1 U9022 ( .A1(n15481), .A2(n7733), .ZN(n7169) );
  OR2_X1 U9023 ( .A1(n15480), .A2(n7734), .ZN(n7733) );
  NOR2_X1 U9024 ( .A1(n6539), .A2(n7955), .ZN(n7954) );
  NAND2_X1 U9025 ( .A1(n7958), .A2(n7959), .ZN(n7956) );
  AND3_X1 U9026 ( .A1(n6936), .A2(n12801), .A3(n12780), .ZN(n12781) );
  INV_X1 U9027 ( .A(n13035), .ZN(n12148) );
  NAND2_X1 U9028 ( .A1(n11854), .A2(n9806), .ZN(n11855) );
  NAND2_X1 U9029 ( .A1(n9340), .A2(n9339), .ZN(n12735) );
  NAND2_X1 U9030 ( .A1(n7957), .A2(n9850), .ZN(n12583) );
  XNOR2_X1 U9031 ( .A(n9798), .B(n13036), .ZN(n11958) );
  XNOR2_X1 U9032 ( .A(n7069), .B(n9834), .ZN(n11095) );
  NAND2_X1 U9033 ( .A1(n9036), .A2(n7610), .ZN(n11092) );
  NAND2_X1 U9034 ( .A1(n9047), .A2(n7609), .ZN(n7610) );
  OAI22_X1 U9035 ( .A1(n10878), .A2(n10849), .B1(n10850), .B2(n8125), .ZN(
        n7609) );
  NAND2_X1 U9036 ( .A1(n7950), .A2(n7949), .ZN(n12740) );
  AND2_X1 U9037 ( .A1(n7950), .A2(n7952), .ZN(n12741) );
  INV_X1 U9038 ( .A(n7948), .ZN(n7949) );
  AND2_X1 U9039 ( .A1(n9454), .A2(n9453), .ZN(n12756) );
  AOI21_X1 U9040 ( .B1(n11052), .B2(n7262), .A(n9293), .ZN(n12769) );
  AOI21_X1 U9041 ( .B1(n12829), .B2(n12760), .A(n12761), .ZN(n12763) );
  AND2_X1 U9042 ( .A1(n7932), .A2(n7934), .ZN(n12772) );
  NAND2_X1 U9043 ( .A1(n7932), .A2(n7930), .ZN(n12770) );
  NAND2_X1 U9044 ( .A1(n12781), .A2(n6937), .ZN(n6934) );
  NAND2_X1 U9045 ( .A1(n6938), .A2(n6937), .ZN(n6935) );
  NAND2_X1 U9046 ( .A1(n7943), .A2(n7940), .ZN(n12789) );
  INV_X1 U9047 ( .A(n7942), .ZN(n7940) );
  NAND2_X1 U9048 ( .A1(n7945), .A2(n7944), .ZN(n7943) );
  OR3_X1 U9049 ( .A1(n9870), .A2(n9869), .A3(n15859), .ZN(n12822) );
  NAND2_X1 U9050 ( .A1(n6942), .A2(n9833), .ZN(n12797) );
  NAND2_X1 U9051 ( .A1(n6947), .A2(n7929), .ZN(n12807) );
  NAND2_X1 U9052 ( .A1(n12829), .A2(n7930), .ZN(n6947) );
  AND2_X1 U9053 ( .A1(n9439), .A2(n9438), .ZN(n13249) );
  INV_X1 U9054 ( .A(n13392), .ZN(n12837) );
  NAND2_X1 U9055 ( .A1(n9866), .A2(n9865), .ZN(n12839) );
  NAND2_X1 U9056 ( .A1(n13026), .A2(n13025), .ZN(n7058) );
  NAND2_X1 U9057 ( .A1(n7293), .A2(n6633), .ZN(n12871) );
  AOI21_X1 U9058 ( .B1(n7057), .B2(n9776), .A(n7056), .ZN(n7055) );
  XNOR2_X1 U9059 ( .A(n12894), .B(n12895), .ZN(n7057) );
  OAI21_X1 U9060 ( .B1(n7574), .B2(n13022), .A(n7573), .ZN(n7056) );
  AND2_X1 U9061 ( .A1(n12861), .A2(n9502), .ZN(n12868) );
  INV_X1 U9062 ( .A(n12823), .ZN(n13217) );
  INV_X1 U9063 ( .A(n13249), .ZN(n13218) );
  NAND2_X1 U9064 ( .A1(n9367), .A2(n9366), .ZN(n13349) );
  NAND2_X1 U9065 ( .A1(n9313), .A2(n9312), .ZN(n13358) );
  OAI211_X1 U9066 ( .C1(n12847), .C2(n13561), .A(n9297), .B(n9296), .ZN(n13373) );
  OAI211_X1 U9067 ( .C1(n12847), .C2(n13567), .A(n9284), .B(n9283), .ZN(n13382) );
  INV_X1 U9068 ( .A(n13403), .ZN(n13381) );
  INV_X1 U9069 ( .A(n11944), .ZN(n13036) );
  AND2_X1 U9070 ( .A1(n9113), .A2(n7071), .ZN(n7070) );
  NAND4_X1 U9071 ( .A1(n9081), .A2(n9080), .A3(n9079), .A4(n9078), .ZN(n13040)
         );
  OR2_X1 U9072 ( .A1(n9041), .A2(n15907), .ZN(n9033) );
  NAND4_X1 U9073 ( .A1(n9025), .A2(n9024), .A3(n9023), .A4(n9022), .ZN(n13044)
         );
  OR2_X2 U9074 ( .A1(n9856), .A2(n10972), .ZN(n13043) );
  NOR2_X1 U9075 ( .A1(n7617), .A2(n7614), .ZN(n11116) );
  INV_X1 U9076 ( .A(n7616), .ZN(n7614) );
  NAND2_X1 U9077 ( .A1(n7442), .A2(n7440), .ZN(n11195) );
  INV_X1 U9078 ( .A(n7441), .ZN(n7440) );
  NAND2_X1 U9079 ( .A1(n7444), .A2(n7443), .ZN(n7442) );
  INV_X1 U9080 ( .A(n7438), .ZN(n7437) );
  OAI21_X1 U9081 ( .B1(n7443), .B2(n7439), .A(n11192), .ZN(n7438) );
  NAND2_X1 U9082 ( .A1(n11147), .A2(n6526), .ZN(n7436) );
  NOR2_X1 U9083 ( .A1(n7618), .A2(n11297), .ZN(n6736) );
  NAND2_X1 U9084 ( .A1(n7423), .A2(n7425), .ZN(n11901) );
  NAND2_X1 U9085 ( .A1(n7243), .A2(n7620), .ZN(n12100) );
  NAND2_X1 U9086 ( .A1(n7125), .A2(n7620), .ZN(n7122) );
  NAND2_X1 U9087 ( .A1(n6732), .A2(n13083), .ZN(n13066) );
  AOI21_X1 U9088 ( .B1(n13053), .B2(n9627), .A(n7518), .ZN(n7512) );
  NAND2_X1 U9089 ( .A1(n7033), .A2(n13133), .ZN(n13132) );
  NAND2_X1 U9090 ( .A1(n7034), .A2(n13112), .ZN(n7033) );
  INV_X1 U9091 ( .A(n13135), .ZN(n7034) );
  AND2_X1 U9092 ( .A1(n7132), .A2(n7131), .ZN(n13128) );
  NOR2_X1 U9093 ( .A1(n13105), .A2(n6529), .ZN(n13120) );
  INV_X1 U9094 ( .A(n13112), .ZN(n13134) );
  NAND2_X1 U9095 ( .A1(n7629), .A2(n9602), .ZN(n13141) );
  NAND2_X1 U9096 ( .A1(n7414), .A2(n7415), .ZN(n13147) );
  AND2_X1 U9097 ( .A1(n6586), .A2(n7414), .ZN(n13145) );
  NAND2_X1 U9098 ( .A1(n13105), .A2(n6720), .ZN(n7414) );
  INV_X1 U9099 ( .A(n9604), .ZN(n7627) );
  XNOR2_X1 U9100 ( .A(n13177), .B(n7272), .ZN(n9634) );
  INV_X1 U9101 ( .A(n13176), .ZN(n7272) );
  NAND2_X1 U9102 ( .A1(n13186), .A2(n9480), .ZN(n12700) );
  NAND2_X1 U9103 ( .A1(n13250), .A2(n12999), .ZN(n13230) );
  NAND2_X1 U9104 ( .A1(n7155), .A2(n7154), .ZN(n13257) );
  NAND2_X1 U9105 ( .A1(n9343), .A2(n9342), .ZN(n13327) );
  CLKBUF_X1 U9106 ( .A(n13398), .Z(n13399) );
  NAND2_X1 U9107 ( .A1(n12090), .A2(n9161), .ZN(n11942) );
  NAND2_X1 U9108 ( .A1(n6819), .A2(n7890), .ZN(n11843) );
  NAND2_X1 U9109 ( .A1(n7321), .A2(n9108), .ZN(n11687) );
  NAND2_X1 U9110 ( .A1(n11535), .A2(n9510), .ZN(n7895) );
  AND3_X1 U9111 ( .A1(n9106), .A2(n9105), .A3(n9104), .ZN(n11614) );
  INV_X1 U9112 ( .A(n13428), .ZN(n13266) );
  INV_X1 U9113 ( .A(n13431), .ZN(n13411) );
  INV_X1 U9114 ( .A(n15855), .ZN(n13427) );
  INV_X1 U9115 ( .A(n13183), .ZN(n13504) );
  NAND2_X1 U9116 ( .A1(n13441), .A2(n13440), .ZN(n13514) );
  INV_X1 U9117 ( .A(n7870), .ZN(n13271) );
  AOI21_X1 U9118 ( .B1(n13280), .B2(n9525), .A(n12988), .ZN(n7870) );
  OAI21_X1 U9119 ( .B1(n9314), .B2(n7605), .A(n7602), .ZN(n13285) );
  INV_X1 U9120 ( .A(n12735), .ZN(n13544) );
  INV_X1 U9121 ( .A(n12811), .ZN(n13550) );
  INV_X1 U9122 ( .A(n12769), .ZN(n13562) );
  INV_X1 U9123 ( .A(n12843), .ZN(n13568) );
  NAND2_X1 U9124 ( .A1(n13415), .A2(n13418), .ZN(n7874) );
  NAND2_X1 U9125 ( .A1(n12146), .A2(n12941), .ZN(n7595) );
  OAI21_X1 U9126 ( .B1(n6842), .B2(n6843), .A(n9047), .ZN(n6844) );
  NOR2_X1 U9127 ( .A1(n8125), .A2(n10836), .ZN(n6843) );
  INV_X1 U9128 ( .A(n13601), .ZN(n10972) );
  AND2_X1 U9129 ( .A1(n9855), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13601) );
  XNOR2_X1 U9130 ( .A(n12552), .B(n9476), .ZN(n12568) );
  INV_X1 U9131 ( .A(n7401), .ZN(n7396) );
  XNOR2_X1 U9132 ( .A(n9545), .B(n9544), .ZN(n13620) );
  OAI21_X1 U9133 ( .B1(n9543), .B2(P3_IR_REG_24__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9545) );
  NAND2_X1 U9134 ( .A1(n9543), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9542) );
  NAND2_X1 U9135 ( .A1(n7804), .A2(n7807), .ZN(n9410) );
  NAND2_X1 U9136 ( .A1(n9375), .A2(n7808), .ZN(n7804) );
  NAND2_X1 U9137 ( .A1(n9386), .A2(n9385), .ZN(n9399) );
  AND2_X1 U9138 ( .A1(n9496), .A2(n6566), .ZN(n13028) );
  NAND2_X1 U9139 ( .A1(n9260), .A2(n7972), .ZN(n9495) );
  NAND2_X1 U9140 ( .A1(n9386), .A2(n9376), .ZN(n11751) );
  XNOR2_X1 U9141 ( .A(n9491), .B(n9490), .ZN(n11699) );
  NAND2_X1 U9142 ( .A1(n7794), .A2(n7792), .ZN(n9353) );
  NAND2_X1 U9143 ( .A1(n7794), .A2(n7795), .ZN(n9351) );
  NAND2_X1 U9144 ( .A1(n9302), .A2(n9301), .ZN(n9316) );
  INV_X1 U9145 ( .A(SI_16_), .ZN(n11053) );
  INV_X1 U9146 ( .A(SI_15_), .ZN(n11014) );
  NAND2_X1 U9147 ( .A1(n7810), .A2(n9275), .ZN(n9291) );
  NAND2_X1 U9148 ( .A1(n9238), .A2(n7814), .ZN(n7810) );
  OR2_X1 U9149 ( .A1(n9246), .A2(n9245), .ZN(n13095) );
  INV_X1 U9150 ( .A(SI_13_), .ZN(n10999) );
  NAND2_X1 U9151 ( .A1(n6806), .A2(n9216), .ZN(n9235) );
  INV_X1 U9152 ( .A(SI_11_), .ZN(n10901) );
  NAND2_X1 U9153 ( .A1(n7774), .A2(n7773), .ZN(n9217) );
  XNOR2_X1 U9154 ( .A(n9191), .B(n9190), .ZN(n10872) );
  NAND2_X1 U9155 ( .A1(n7775), .A2(n9189), .ZN(n9202) );
  NAND2_X1 U9156 ( .A1(n9188), .A2(n9187), .ZN(n7775) );
  NAND2_X1 U9157 ( .A1(n6805), .A2(n6629), .ZN(n9164) );
  OAI21_X1 U9158 ( .B1(n9117), .B2(n7784), .A(n7782), .ZN(n9155) );
  NAND2_X1 U9159 ( .A1(n7787), .A2(n9119), .ZN(n9138) );
  NAND2_X1 U9160 ( .A1(n9117), .A2(n9116), .ZN(n7787) );
  NAND2_X1 U9161 ( .A1(n6787), .A2(n9082), .ZN(n9097) );
  NAND2_X1 U9162 ( .A1(n6793), .A2(n6791), .ZN(n6787) );
  NAND2_X1 U9163 ( .A1(n9102), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7030) );
  NAND2_X1 U9164 ( .A1(n9063), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6735) );
  NAND2_X1 U9165 ( .A1(n6793), .A2(n9067), .ZN(n9084) );
  INV_X1 U9166 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n12295) );
  NAND2_X1 U9167 ( .A1(n12119), .A2(n12712), .ZN(n12721) );
  NAND2_X1 U9168 ( .A1(n11713), .A2(n13820), .ZN(n10799) );
  INV_X1 U9169 ( .A(n12634), .ZN(n7209) );
  AND2_X1 U9170 ( .A1(n12639), .A2(n7207), .ZN(n7206) );
  AND2_X1 U9171 ( .A1(n10564), .A2(n10573), .ZN(n14232) );
  AND2_X1 U9172 ( .A1(n10819), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13750) );
  XNOR2_X1 U9173 ( .A(n11417), .B(n11418), .ZN(n11459) );
  OR2_X1 U9174 ( .A1(n12119), .A2(n6531), .ZN(n7678) );
  INV_X1 U9175 ( .A(n14094), .ZN(n14475) );
  AND2_X1 U9176 ( .A1(n12232), .A2(n12131), .ZN(n12599) );
  NOR2_X1 U9177 ( .A1(n13789), .A2(n14474), .ZN(n13769) );
  NOR2_X1 U9178 ( .A1(n13789), .A2(n14472), .ZN(n13770) );
  INV_X1 U9179 ( .A(n13796), .ZN(n13798) );
  INV_X1 U9180 ( .A(n13770), .ZN(n13805) );
  NAND2_X1 U9181 ( .A1(n11712), .A2(n11711), .ZN(n11760) );
  CLKBUF_X1 U9182 ( .A(n11275), .Z(n14102) );
  INV_X2 U9183 ( .A(P2_U3947), .ZN(n14103) );
  NAND2_X1 U9184 ( .A1(n15613), .A2(n11254), .ZN(n15627) );
  NAND2_X1 U9185 ( .A1(n14131), .A2(n11260), .ZN(n15652) );
  NAND2_X1 U9186 ( .A1(n15652), .A2(n15653), .ZN(n15651) );
  NAND2_X1 U9187 ( .A1(n7494), .A2(n7495), .ZN(n15665) );
  NAND2_X1 U9188 ( .A1(n15667), .A2(n6892), .ZN(n15686) );
  NOR2_X1 U9189 ( .A1(n11641), .A2(n7505), .ZN(n15698) );
  AND2_X1 U9190 ( .A1(n11644), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7505) );
  NAND2_X1 U9191 ( .A1(n15698), .A2(n15699), .ZN(n15697) );
  INV_X1 U9192 ( .A(n15709), .ZN(n6896) );
  INV_X1 U9193 ( .A(n6897), .ZN(n15710) );
  INV_X1 U9194 ( .A(n7501), .ZN(n14164) );
  NAND2_X1 U9195 ( .A1(n10722), .A2(n7645), .ZN(n14178) );
  AOI21_X1 U9196 ( .B1(n6777), .B2(n15781), .A(n14199), .ZN(n6776) );
  INV_X1 U9197 ( .A(n14507), .ZN(n6777) );
  NAND2_X1 U9198 ( .A1(n7981), .A2(n7982), .ZN(n14250) );
  NAND2_X1 U9199 ( .A1(n7989), .A2(n7983), .ZN(n7981) );
  NAND2_X1 U9200 ( .A1(n7987), .A2(n7985), .ZN(n14271) );
  INV_X1 U9201 ( .A(n7986), .ZN(n7985) );
  NAND2_X1 U9202 ( .A1(n7988), .A2(n7989), .ZN(n7987) );
  NAND2_X1 U9203 ( .A1(n7912), .A2(n7914), .ZN(n14278) );
  NAND2_X1 U9204 ( .A1(n14305), .A2(n6528), .ZN(n7912) );
  NAND2_X1 U9205 ( .A1(n7916), .A2(n10620), .ZN(n14291) );
  OR2_X1 U9206 ( .A1(n14305), .A2(n10619), .ZN(n7916) );
  NAND2_X1 U9207 ( .A1(n14334), .A2(n10519), .ZN(n14324) );
  NAND2_X1 U9208 ( .A1(n10610), .A2(n7887), .ZN(n7886) );
  NAND2_X1 U9209 ( .A1(n10610), .A2(n10609), .ZN(n14395) );
  NAND2_X1 U9210 ( .A1(n7976), .A2(n7979), .ZN(n14402) );
  NAND2_X1 U9211 ( .A1(n7978), .A2(n7977), .ZN(n7976) );
  NAND2_X1 U9212 ( .A1(n10242), .A2(n10241), .ZN(n14588) );
  NAND2_X1 U9213 ( .A1(n8008), .A2(n10455), .ZN(n14466) );
  NAND2_X1 U9214 ( .A1(n7907), .A2(n10593), .ZN(n11931) );
  NAND2_X1 U9215 ( .A1(n10592), .A2(n7908), .ZN(n7907) );
  NAND2_X1 U9216 ( .A1(n10592), .A2(n11785), .ZN(n15757) );
  INV_X1 U9217 ( .A(n14436), .ZN(n15763) );
  INV_X1 U9218 ( .A(n12012), .ZN(n10198) );
  NOR3_X1 U9219 ( .A1(n14182), .A2(n14494), .A3(n14499), .ZN(n14509) );
  INV_X1 U9220 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n7993) );
  INV_X1 U9221 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n7362) );
  INV_X1 U9222 ( .A(n14432), .ZN(n14645) );
  INV_X1 U9223 ( .A(n14483), .ZN(n14653) );
  NAND2_X1 U9224 ( .A1(n10222), .A2(n10251), .ZN(n8010) );
  NAND2_X1 U9225 ( .A1(n10838), .A2(n10188), .ZN(n10195) );
  INV_X1 U9226 ( .A(n15789), .ZN(n15790) );
  AND2_X1 U9227 ( .A1(n12037), .A2(n10809), .ZN(n15796) );
  AND2_X1 U9228 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10808), .ZN(n10809) );
  INV_X1 U9229 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n14657) );
  NAND2_X1 U9230 ( .A1(n6920), .A2(n6921), .ZN(n10321) );
  INV_X1 U9231 ( .A(n6922), .ZN(n6921) );
  INV_X1 U9232 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n10340) );
  NAND2_X1 U9233 ( .A1(n10339), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10341) );
  NAND2_X1 U9234 ( .A1(n10351), .A2(n12438), .ZN(n10339) );
  NAND2_X1 U9235 ( .A1(n10285), .A2(n10284), .ZN(n11872) );
  INV_X1 U9236 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n12359) );
  NAND2_X1 U9237 ( .A1(n10232), .A2(n10172), .ZN(n10266) );
  INV_X1 U9238 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11217) );
  INV_X1 U9239 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n12274) );
  INV_X1 U9240 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11323) );
  INV_X1 U9241 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n11051) );
  AND2_X1 U9242 ( .A1(n10248), .A2(n10253), .ZN(n14149) );
  INV_X1 U9243 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10967) );
  INV_X1 U9244 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10945) );
  INV_X1 U9245 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10910) );
  INV_X1 U9246 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10883) );
  INV_X1 U9247 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10839) );
  NAND2_X1 U9248 ( .A1(n10182), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10183) );
  NAND2_X1 U9249 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n6900) );
  INV_X1 U9250 ( .A(P2_STATE_REG_SCAN_IN), .ZN(n11242) );
  NAND2_X1 U9251 ( .A1(n7748), .A2(n7746), .ZN(n11701) );
  AND2_X1 U9252 ( .A1(n9919), .A2(n9908), .ZN(n7737) );
  INV_X1 U9253 ( .A(n15497), .ZN(n9919) );
  AND2_X1 U9254 ( .A1(n7761), .A2(n6582), .ZN(n14701) );
  AND2_X1 U9255 ( .A1(n10131), .A2(n14813), .ZN(n7344) );
  AOI21_X1 U9256 ( .B1(n7746), .B2(n11513), .A(n6540), .ZN(n7744) );
  INV_X1 U9257 ( .A(n7746), .ZN(n7745) );
  NAND2_X1 U9258 ( .A1(n14763), .A2(n7742), .ZN(n7738) );
  AND3_X1 U9259 ( .A1(n8483), .A2(n8482), .A3(n8481), .ZN(n15228) );
  INV_X1 U9260 ( .A(n14773), .ZN(n14826) );
  AOI21_X1 U9261 ( .B1(n14763), .B2(n14762), .A(n7743), .ZN(n14765) );
  NAND2_X1 U9262 ( .A1(n9924), .A2(n9925), .ZN(n11345) );
  AND2_X1 U9263 ( .A1(n6852), .A2(n6691), .ZN(n7759) );
  OR2_X1 U9264 ( .A1(n14677), .A2(n10002), .ZN(n14782) );
  NAND2_X1 U9265 ( .A1(n8466), .A2(n8465), .ZN(n14788) );
  NAND2_X1 U9266 ( .A1(n6860), .A2(n6861), .ZN(n14796) );
  NAND2_X1 U9267 ( .A1(n7763), .A2(n9971), .ZN(n12165) );
  NAND2_X1 U9268 ( .A1(n11862), .A2(n7764), .ZN(n7763) );
  NAND2_X1 U9269 ( .A1(n8756), .A2(n8755), .ZN(n14835) );
  OR3_X1 U9270 ( .A1(n15005), .A2(n8750), .A3(n15004), .ZN(n8756) );
  NAND2_X1 U9271 ( .A1(n8772), .A2(n8771), .ZN(n14982) );
  INV_X1 U9272 ( .A(n14815), .ZN(n14838) );
  NAND2_X1 U9273 ( .A1(n8657), .A2(n8656), .ZN(n15031) );
  OR2_X1 U9274 ( .A1(n15056), .A2(n8750), .ZN(n8657) );
  NAND2_X1 U9275 ( .A1(n6514), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8245) );
  NAND2_X1 U9276 ( .A1(n10952), .A2(n10734), .ZN(n11003) );
  OR2_X1 U9277 ( .A1(n10751), .A2(n14961), .ZN(n10752) );
  INV_X1 U9278 ( .A(n12215), .ZN(n14954) );
  INV_X1 U9279 ( .A(n15269), .ZN(n14974) );
  INV_X1 U9280 ( .A(n14977), .ZN(n15274) );
  NAND2_X1 U9281 ( .A1(n7553), .A2(n7554), .ZN(n8039) );
  AOI21_X1 U9282 ( .B1(n10662), .B2(n15545), .A(n10661), .ZN(n15286) );
  NAND2_X1 U9283 ( .A1(n15082), .A2(n8952), .ZN(n15065) );
  OAI21_X1 U9284 ( .B1(n15123), .B2(n7542), .A(n7540), .ZN(n15075) );
  NAND2_X1 U9285 ( .A1(n7539), .A2(n7545), .ZN(n15077) );
  NAND2_X1 U9286 ( .A1(n15123), .A2(n8907), .ZN(n15109) );
  INV_X1 U9287 ( .A(n15319), .ZN(n15107) );
  AND2_X1 U9288 ( .A1(n15155), .A2(n8944), .ZN(n15135) );
  NAND2_X1 U9289 ( .A1(n8036), .A2(n8904), .ZN(n15133) );
  OR2_X1 U9290 ( .A1(n15149), .A2(n8905), .ZN(n8036) );
  NAND2_X1 U9291 ( .A1(n7546), .A2(n8902), .ZN(n15185) );
  OR2_X1 U9292 ( .A1(n15189), .A2(n8901), .ZN(n7546) );
  OAI21_X1 U9293 ( .B1(n12192), .B2(n8046), .A(n8044), .ZN(n15247) );
  NAND2_X1 U9294 ( .A1(n12190), .A2(n8931), .ZN(n15249) );
  NAND2_X1 U9295 ( .A1(n11918), .A2(n8929), .ZN(n11993) );
  NOR2_X1 U9296 ( .A1(n7485), .A2(n7487), .ZN(n11831) );
  INV_X1 U9297 ( .A(n11674), .ZN(n7485) );
  NAND2_X1 U9298 ( .A1(n11580), .A2(n11581), .ZN(n8025) );
  NAND2_X1 U9299 ( .A1(n10863), .A2(n8775), .ZN(n6979) );
  NAND2_X1 U9300 ( .A1(n9892), .A2(n15257), .ZN(n11028) );
  NAND2_X1 U9301 ( .A1(n9892), .A2(n15256), .ZN(n11450) );
  INV_X1 U9302 ( .A(n15267), .ZN(n15242) );
  AND2_X1 U9303 ( .A1(n12692), .A2(n8976), .ZN(n8977) );
  NOR2_X1 U9304 ( .A1(n8090), .A2(n8089), .ZN(n8976) );
  AOI21_X1 U9305 ( .B1(n7491), .B2(n15545), .A(n15023), .ZN(n15291) );
  AND2_X2 U9306 ( .A1(n9002), .A2(n9001), .ZN(n15588) );
  OAI21_X1 U9307 ( .B1(n8812), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8811) );
  NAND2_X1 U9308 ( .A1(n10867), .A2(n10866), .ZN(n15531) );
  AND2_X1 U9309 ( .A1(n7279), .A2(n8199), .ZN(n7471) );
  XNOR2_X1 U9310 ( .A(n8774), .B(n8773), .ZN(n10297) );
  NOR2_X1 U9311 ( .A1(n7278), .A2(n7277), .ZN(n7276) );
  NOR2_X1 U9312 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n7277) );
  NAND2_X1 U9313 ( .A1(n7835), .A2(n7833), .ZN(n8677) );
  INV_X1 U9314 ( .A(n8969), .ZN(n15440) );
  NAND2_X1 U9315 ( .A1(n6987), .A2(n8184), .ZN(n8611) );
  NAND2_X1 U9316 ( .A1(n8591), .A2(n8181), .ZN(n6987) );
  INV_X1 U9317 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11780) );
  INV_X1 U9318 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11657) );
  OR2_X1 U9319 ( .A1(n8502), .A2(n8501), .ZN(n8504) );
  INV_X1 U9320 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11214) );
  INV_X1 U9321 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n11320) );
  XNOR2_X1 U9322 ( .A(n8443), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11621) );
  INV_X1 U9323 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n11047) );
  INV_X1 U9324 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n12309) );
  AND2_X1 U9325 ( .A1(n8420), .A2(n8435), .ZN(n11166) );
  INV_X1 U9326 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n12483) );
  INV_X1 U9327 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n12296) );
  XNOR2_X1 U9328 ( .A(n8285), .B(P1_IR_REG_2__SCAN_IN), .ZN(n14879) );
  MUX2_X1 U9329 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n8125), .Z(n7838) );
  XNOR2_X1 U9330 ( .A(n8254), .B(P1_IR_REG_1__SCAN_IN), .ZN(n14859) );
  NAND2_X1 U9331 ( .A1(n15448), .A2(n15450), .ZN(n15929) );
  XNOR2_X1 U9332 ( .A(n9731), .B(n9732), .ZN(n15923) );
  NAND2_X1 U9333 ( .A1(n15923), .A2(n15922), .ZN(n15921) );
  XNOR2_X1 U9334 ( .A(n9736), .B(n7735), .ZN(n15455) );
  NOR2_X1 U9335 ( .A1(n15455), .A2(n15454), .ZN(n15453) );
  NAND2_X1 U9336 ( .A1(n6754), .A2(n7174), .ZN(n15477) );
  NAND2_X1 U9337 ( .A1(n7382), .A2(n15475), .ZN(n15481) );
  OAI21_X1 U9338 ( .B1(n15477), .B2(n15476), .A(n15705), .ZN(n7382) );
  NAND2_X1 U9339 ( .A1(n7169), .A2(n7732), .ZN(n15485) );
  OAI21_X1 U9340 ( .B1(n15444), .B2(n15445), .A(n15756), .ZN(n7256) );
  NAND2_X1 U9341 ( .A1(n11330), .A2(n9787), .ZN(n11526) );
  XNOR2_X1 U9342 ( .A(n13179), .B(n13178), .ZN(n7038) );
  NAND2_X1 U9343 ( .A1(n6728), .A2(n13097), .ZN(n6727) );
  OAI211_X1 U9344 ( .C1(n13509), .C2(n15873), .A(n6635), .B(n6808), .ZN(
        P3_U3204) );
  NAND2_X1 U9345 ( .A1(n15873), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n6808) );
  OAI21_X1 U9346 ( .B1(n7600), .B2(n7599), .A(n7596), .ZN(n13437) );
  OR2_X1 U9347 ( .A1(n13204), .A2(n10706), .ZN(n7599) );
  NAND2_X1 U9348 ( .A1(n13207), .A2(n13488), .ZN(n10695) );
  OAI211_X1 U9349 ( .C1(n13509), .C2(n15906), .A(n6544), .B(n6695), .ZN(
        P3_U3456) );
  NOR2_X1 U9350 ( .A1(n9581), .A2(n9582), .ZN(n9583) );
  AND2_X1 U9351 ( .A1(n13632), .A2(n6714), .ZN(n7322) );
  NAND2_X1 U9352 ( .A1(n13783), .A2(n7364), .ZN(n13795) );
  OAI21_X1 U9353 ( .B1(n14079), .B2(n14065), .A(n14064), .ZN(n14084) );
  AOI21_X1 U9354 ( .B1(n14079), .B2(n7316), .A(n7315), .ZN(n7314) );
  NAND2_X1 U9355 ( .A1(n6889), .A2(n6883), .ZN(n6877) );
  INV_X1 U9356 ( .A(n6880), .ZN(n6879) );
  NAND2_X1 U9357 ( .A1(n6774), .A2(n6773), .ZN(P2_U3236) );
  NAND2_X1 U9358 ( .A1(n14504), .A2(n15770), .ZN(n6773) );
  INV_X1 U9359 ( .A(n6775), .ZN(n6774) );
  OAI21_X1 U9360 ( .B1(n14200), .B2(n14421), .A(n6776), .ZN(n6775) );
  NAND2_X1 U9361 ( .A1(n6976), .A2(n15781), .ZN(n6975) );
  AOI21_X1 U9362 ( .B1(n7995), .B2(n15770), .A(n14207), .ZN(n6974) );
  NAND2_X1 U9363 ( .A1(n6597), .A2(n7306), .ZN(P2_U3238) );
  INV_X1 U9364 ( .A(n7307), .ZN(n7306) );
  OAI21_X1 U9365 ( .B1(n14214), .B2(n14421), .A(n7308), .ZN(n7307) );
  NAND2_X1 U9366 ( .A1(n7285), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7284) );
  NOR2_X1 U9367 ( .A1(n6707), .A2(n6541), .ZN(n7385) );
  INV_X1 U9368 ( .A(n7378), .ZN(n7377) );
  OAI21_X1 U9369 ( .B1(n14511), .B2(n14602), .A(n7379), .ZN(n7378) );
  AOI21_X1 U9370 ( .B1(n14217), .B2(n12142), .A(n7319), .ZN(n7318) );
  NOR2_X1 U9371 ( .A1(n15848), .A2(n14515), .ZN(n7319) );
  NAND2_X1 U9372 ( .A1(n7304), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7286) );
  NOR2_X1 U9373 ( .A1(n6607), .A2(n7992), .ZN(n7991) );
  NAND2_X1 U9374 ( .A1(n10723), .A2(n15838), .ZN(n7994) );
  NOR2_X1 U9375 ( .A1(n15838), .A2(n7993), .ZN(n7992) );
  NAND2_X1 U9376 ( .A1(n7363), .A2(n7360), .ZN(P2_U3494) );
  NOR2_X1 U9377 ( .A1(n6700), .A2(n7361), .ZN(n7360) );
  NAND2_X1 U9378 ( .A1(n14510), .A2(n15838), .ZN(n7363) );
  NOR2_X1 U9379 ( .A1(n15838), .A2(n7362), .ZN(n7361) );
  OAI21_X1 U9380 ( .B1(n14618), .B2(n7304), .A(n7302), .ZN(P2_U3493) );
  AND2_X1 U9381 ( .A1(n7367), .A2(n7303), .ZN(n7302) );
  NAND2_X1 U9382 ( .A1(n7304), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n7303) );
  NAND2_X1 U9383 ( .A1(n14217), .A2(n7368), .ZN(n7367) );
  OAI21_X1 U9384 ( .B1(n7840), .B2(n15503), .A(n10155), .ZN(n10156) );
  AOI22_X1 U9385 ( .A1(n14830), .A2(n11055), .B1(n14773), .B2(n9892), .ZN(
        n11059) );
  AOI21_X1 U9386 ( .B1(n7372), .B2(n12005), .A(n7369), .ZN(n8871) );
  NAND2_X1 U9387 ( .A1(n7479), .A2(n7478), .ZN(P1_U3561) );
  NAND2_X1 U9388 ( .A1(P1_U4016), .A2(n9892), .ZN(n7478) );
  OR2_X1 U9389 ( .A1(P1_U4016), .A2(n10847), .ZN(n7479) );
  NOR2_X1 U9390 ( .A1(n10797), .A2(n14704), .ZN(n7241) );
  NAND2_X1 U9391 ( .A1(n10793), .A2(n15199), .ZN(n7242) );
  NAND2_X1 U9392 ( .A1(n10792), .A2(n15163), .ZN(n7240) );
  NAND2_X1 U9393 ( .A1(n7492), .A2(n7489), .ZN(n7488) );
  NAND2_X1 U9394 ( .A1(n15023), .A2(n15232), .ZN(n7489) );
  INV_X1 U9395 ( .A(n7386), .ZN(n15932) );
  INV_X1 U9396 ( .A(n15450), .ZN(n15449) );
  INV_X1 U9397 ( .A(n6745), .ZN(n15920) );
  NAND2_X1 U9398 ( .A1(n6743), .A2(n6744), .ZN(n6745) );
  INV_X1 U9399 ( .A(n6749), .ZN(n15925) );
  NAND2_X1 U9400 ( .A1(n15460), .A2(n15459), .ZN(n15458) );
  NAND2_X1 U9401 ( .A1(n15456), .A2(n9743), .ZN(n15460) );
  INV_X1 U9402 ( .A(n9747), .ZN(n15462) );
  INV_X1 U9403 ( .A(n15472), .ZN(n15471) );
  INV_X1 U9404 ( .A(n7729), .ZN(n15487) );
  AND2_X1 U9405 ( .A1(n7728), .A2(n7729), .ZN(n15492) );
  NOR2_X1 U9406 ( .A1(n15467), .A2(n15468), .ZN(n15466) );
  INV_X1 U9407 ( .A(n15445), .ZN(n7332) );
  INV_X1 U9408 ( .A(n15881), .ZN(n7250) );
  AND4_X1 U9409 ( .A1(n8205), .A2(n8211), .A3(n8210), .A4(n8209), .ZN(n6523)
         );
  AND2_X1 U9410 ( .A1(n14619), .A2(n14088), .ZN(n6524) );
  NAND2_X1 U9412 ( .A1(n10281), .A2(n10280), .ZN(n14539) );
  INV_X1 U9413 ( .A(n14522), .ZN(n14257) );
  OAI21_X1 U9414 ( .B1(n12162), .B2(n8679), .A(n8650), .ZN(n15053) );
  OR2_X1 U9415 ( .A1(n14351), .A2(n7661), .ZN(n6525) );
  NOR2_X1 U9416 ( .A1(n7441), .A2(n11191), .ZN(n6526) );
  AND2_X1 U9417 ( .A1(n6891), .A2(n6711), .ZN(n6527) );
  NOR2_X1 U9418 ( .A1(n10621), .A2(n7915), .ZN(n6528) );
  XNOR2_X1 U9419 ( .A(n6735), .B(n6734), .ZN(n10833) );
  NAND2_X1 U9420 ( .A1(n15155), .A2(n8064), .ZN(n15094) );
  AND2_X1 U9421 ( .A1(n9678), .A2(n13111), .ZN(n6529) );
  OR2_X1 U9422 ( .A1(n12779), .A2(n9841), .ZN(n6530) );
  INV_X1 U9423 ( .A(n8929), .ZN(n8048) );
  XNOR2_X1 U9424 ( .A(n15289), .B(n15032), .ZN(n15021) );
  INV_X1 U9425 ( .A(n15021), .ZN(n7556) );
  AND2_X1 U9426 ( .A1(n6945), .A2(n9833), .ZN(n12750) );
  AND2_X1 U9427 ( .A1(n12121), .A2(n12120), .ZN(n6531) );
  INV_X1 U9428 ( .A(n8928), .ZN(n8049) );
  AND2_X1 U9429 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n6532) );
  AND2_X1 U9430 ( .A1(n6655), .A2(n7074), .ZN(n6533) );
  AND3_X1 U9431 ( .A1(n14222), .A2(n14057), .A3(n14235), .ZN(n6534) );
  OR2_X1 U9432 ( .A1(n9515), .A2(n12961), .ZN(n6535) );
  AND3_X1 U9433 ( .A1(n13370), .A2(n13418), .A3(n13405), .ZN(n6536) );
  INV_X1 U9434 ( .A(n13858), .ZN(n7911) );
  OR2_X1 U9435 ( .A1(n9892), .A2(n15535), .ZN(n6537) );
  OAI21_X1 U9436 ( .B1(n12761), .B2(n12760), .A(n6656), .ZN(n7935) );
  AND2_X1 U9437 ( .A1(n7973), .A2(n7113), .ZN(n6538) );
  NOR2_X1 U9438 ( .A1(n9850), .A2(n9848), .ZN(n6539) );
  AND2_X1 U9439 ( .A1(n9949), .A2(n9948), .ZN(n6540) );
  INV_X1 U9440 ( .A(n10073), .ZN(n15309) );
  INV_X1 U9441 ( .A(n14568), .ZN(n7663) );
  NOR2_X1 U9442 ( .A1(n14205), .A2(n14602), .ZN(n6541) );
  NOR2_X1 U9443 ( .A1(n14528), .A2(n13717), .ZN(n6542) );
  NAND2_X1 U9444 ( .A1(n9251), .A2(n6699), .ZN(n6543) );
  INV_X1 U9445 ( .A(n13532), .ZN(n6798) );
  INV_X1 U9446 ( .A(n7463), .ZN(n7462) );
  NOR2_X1 U9447 ( .A1(n8628), .A2(n8629), .ZN(n7463) );
  AND2_X1 U9448 ( .A1(n7253), .A2(n13512), .ZN(n6544) );
  INV_X1 U9449 ( .A(n8206), .ZN(n7758) );
  AND2_X1 U9450 ( .A1(n7348), .A2(n12664), .ZN(n6545) );
  INV_X1 U9451 ( .A(n15289), .ZN(n15020) );
  AND2_X1 U9452 ( .A1(n13893), .A2(n7725), .ZN(n6546) );
  NAND2_X1 U9453 ( .A1(n6798), .A2(n6797), .ZN(n9526) );
  INV_X1 U9454 ( .A(n9526), .ZN(n12988) );
  AND2_X1 U9455 ( .A1(n14580), .A2(n14397), .ZN(n6547) );
  AND2_X1 U9456 ( .A1(n14166), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6548) );
  OR2_X1 U9457 ( .A1(n7342), .A2(n15474), .ZN(n6549) );
  AND2_X1 U9458 ( .A1(n10168), .A2(n10318), .ZN(n6550) );
  NAND2_X1 U9459 ( .A1(n9200), .A2(n6673), .ZN(n6551) );
  INV_X2 U9460 ( .A(n15873), .ZN(n15870) );
  AND2_X2 U9461 ( .A1(n11107), .A2(n15855), .ZN(n15873) );
  NAND2_X1 U9462 ( .A1(n15713), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6552) );
  INV_X1 U9463 ( .A(n9842), .ZN(n7967) );
  OR2_X1 U9464 ( .A1(n10998), .A2(n7517), .ZN(n6553) );
  AND2_X1 U9465 ( .A1(n6967), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6554) );
  AND2_X1 U9466 ( .A1(n6970), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6555) );
  AND2_X1 U9467 ( .A1(n10579), .A2(n10578), .ZN(n10649) );
  INV_X1 U9468 ( .A(n10649), .ZN(n14088) );
  NAND2_X1 U9469 ( .A1(n11571), .A2(n7856), .ZN(n7857) );
  OR2_X1 U9470 ( .A1(n9924), .A2(n9925), .ZN(n6556) );
  INV_X1 U9471 ( .A(n13111), .ZN(n7404) );
  AND2_X1 U9472 ( .A1(n6933), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6557) );
  AND2_X1 U9473 ( .A1(n6928), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6558) );
  INV_X1 U9474 ( .A(n15053), .ZN(n7858) );
  INV_X1 U9475 ( .A(n6956), .ZN(n11815) );
  NAND2_X1 U9476 ( .A1(n9144), .A2(n6631), .ZN(n6956) );
  NAND2_X1 U9477 ( .A1(n9037), .A2(n11092), .ZN(n7156) );
  INV_X2 U9478 ( .A(n10316), .ZN(n14066) );
  NAND2_X1 U9479 ( .A1(n15030), .A2(n14838), .ZN(n6559) );
  OR2_X1 U9480 ( .A1(n10017), .A2(n10016), .ZN(n7329) );
  INV_X2 U9481 ( .A(n7879), .ZN(n10720) );
  NAND2_X1 U9482 ( .A1(n9066), .A2(n9065), .ZN(n6793) );
  INV_X1 U9483 ( .A(n15535), .ZN(n14709) );
  XNOR2_X1 U9484 ( .A(n9103), .B(n9121), .ZN(n11202) );
  OR2_X1 U9485 ( .A1(n10594), .A2(n7906), .ZN(n6562) );
  OR2_X1 U9486 ( .A1(n14325), .A2(n14544), .ZN(n6563) );
  XNOR2_X1 U9487 ( .A(n9488), .B(P3_IR_REG_21__SCAN_IN), .ZN(n9778) );
  INV_X1 U9488 ( .A(n13037), .ZN(n6954) );
  AND2_X1 U9489 ( .A1(n7653), .A2(n14234), .ZN(n6564) );
  AND2_X1 U9490 ( .A1(n9030), .A2(n6844), .ZN(n11327) );
  XOR2_X1 U9491 ( .A(n15269), .B(n14973), .Z(n6565) );
  NAND2_X1 U9492 ( .A1(n9260), .A2(n7970), .ZN(n6566) );
  INV_X1 U9493 ( .A(n14025), .ZN(n12561) );
  NAND2_X1 U9494 ( .A1(n10302), .A2(n13981), .ZN(n14025) );
  OR2_X1 U9495 ( .A1(n7753), .A2(n7139), .ZN(n6567) );
  XNOR2_X1 U9496 ( .A(n13194), .B(n9531), .ZN(n6568) );
  NAND3_X1 U9497 ( .A1(n7877), .A2(n6579), .A3(n10374), .ZN(n14104) );
  AND2_X1 U9498 ( .A1(n12934), .A2(n12935), .ZN(n6569) );
  INV_X1 U9499 ( .A(n12761), .ZN(n7936) );
  AND2_X1 U9500 ( .A1(n14184), .A2(n14183), .ZN(n14499) );
  AND2_X1 U9501 ( .A1(n7710), .A2(n7715), .ZN(n6570) );
  NOR2_X1 U9502 ( .A1(n7935), .A2(n7931), .ZN(n7930) );
  AND2_X1 U9503 ( .A1(n8049), .A2(n8927), .ZN(n6571) );
  AND2_X1 U9504 ( .A1(n15342), .A2(n14841), .ZN(n6572) );
  NAND2_X1 U9505 ( .A1(n14877), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n6573) );
  OR2_X1 U9506 ( .A1(n8414), .A2(n6857), .ZN(n6574) );
  NAND2_X1 U9507 ( .A1(n9300), .A2(n9299), .ZN(n9302) );
  NAND2_X1 U9508 ( .A1(n12205), .A2(n13402), .ZN(n6576) );
  AND2_X1 U9509 ( .A1(n9244), .A2(n12489), .ZN(n6577) );
  INV_X1 U9510 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n8020) );
  NOR2_X1 U9511 ( .A1(n15468), .A2(n7564), .ZN(n6578) );
  XNOR2_X1 U9512 ( .A(n10177), .B(n6900), .ZN(n14105) );
  INV_X1 U9513 ( .A(n11297), .ZN(n9650) );
  OAI21_X1 U9514 ( .B1(n7007), .B2(n7006), .A(n14735), .ZN(n7004) );
  OR2_X1 U9515 ( .A1(n10381), .A2(n7881), .ZN(n6579) );
  NAND2_X1 U9516 ( .A1(n12628), .A2(n13696), .ZN(n6580) );
  INV_X1 U9517 ( .A(n14060), .ZN(n14616) );
  NAND2_X1 U9518 ( .A1(n10170), .A2(n10169), .ZN(n14060) );
  AND4_X1 U9519 ( .A1(n10427), .A2(n10426), .A3(n10425), .A4(n10424), .ZN(
        n13859) );
  NAND2_X1 U9520 ( .A1(n9597), .A2(n10998), .ZN(n13083) );
  XNOR2_X1 U9521 ( .A(n8207), .B(n8210), .ZN(n8970) );
  INV_X1 U9522 ( .A(n14528), .ZN(n14273) );
  NAND2_X1 U9523 ( .A1(n10288), .A2(n10287), .ZN(n14528) );
  XNOR2_X1 U9524 ( .A(n6956), .B(n6954), .ZN(n12924) );
  AND3_X1 U9525 ( .A1(n8205), .A2(n7471), .A3(n8106), .ZN(n6581) );
  NAND2_X1 U9526 ( .A1(n10038), .A2(n10037), .ZN(n6582) );
  INV_X1 U9527 ( .A(n9834), .ZN(n9781) );
  INV_X1 U9528 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9244) );
  AND2_X1 U9529 ( .A1(n11262), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6583) );
  INV_X1 U9530 ( .A(n7952), .ZN(n7951) );
  NAND2_X1 U9531 ( .A1(n9828), .A2(n13288), .ZN(n7952) );
  AND2_X1 U9532 ( .A1(n9824), .A2(n13349), .ZN(n6584) );
  OR2_X1 U9533 ( .A1(n9728), .A2(n15625), .ZN(n6585) );
  NAND2_X1 U9534 ( .A1(n6966), .A2(n8900), .ZN(n15189) );
  AND2_X1 U9535 ( .A1(n7415), .A2(n7413), .ZN(n6586) );
  NAND2_X1 U9536 ( .A1(n7595), .A2(n9200), .ZN(n13417) );
  NAND2_X1 U9537 ( .A1(n7886), .A2(n7889), .ZN(n14373) );
  AND2_X1 U9538 ( .A1(n7329), .A2(n7328), .ZN(n6587) );
  AND2_X1 U9539 ( .A1(n15064), .A2(n6847), .ZN(n6588) );
  OR2_X1 U9540 ( .A1(n8530), .A2(n11067), .ZN(n6589) );
  AND2_X1 U9541 ( .A1(n15459), .A2(n9744), .ZN(n6590) );
  INV_X1 U9542 ( .A(n8904), .ZN(n8035) );
  AND2_X1 U9543 ( .A1(n7389), .A2(n7043), .ZN(n6591) );
  OAI21_X2 U9544 ( .B1(n11872), .B2(n10292), .A(n10286), .ZN(n14284) );
  AND2_X1 U9545 ( .A1(n13532), .A2(n9384), .ZN(n12989) );
  INV_X1 U9546 ( .A(n11785), .ZN(n7909) );
  OR2_X1 U9547 ( .A1(n12994), .A2(n13011), .ZN(n6592) );
  OR2_X1 U9548 ( .A1(n15459), .A2(n9744), .ZN(n6593) );
  NOR2_X1 U9549 ( .A1(n13038), .A2(n15896), .ZN(n12922) );
  INV_X1 U9550 ( .A(n14202), .ZN(n7995) );
  AND4_X1 U9551 ( .A1(n10443), .A2(n10442), .A3(n10441), .A4(n10440), .ZN(
        n13868) );
  INV_X1 U9552 ( .A(n13868), .ZN(n8009) );
  AND4_X1 U9553 ( .A1(n12301), .A2(n8329), .A3(n8440), .A4(n8102), .ZN(n6594)
         );
  INV_X1 U9554 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n9017) );
  AND2_X1 U9555 ( .A1(n14282), .A2(n6528), .ZN(n6595) );
  XNOR2_X1 U9556 ( .A(n9542), .B(n9541), .ZN(n9558) );
  INV_X1 U9557 ( .A(n8403), .ZN(n7459) );
  AND2_X1 U9558 ( .A1(n12923), .A2(n13011), .ZN(n6596) );
  INV_X1 U9559 ( .A(n14605), .ZN(n7655) );
  INV_X1 U9560 ( .A(n8697), .ZN(n7258) );
  OR2_X1 U9561 ( .A1(n14211), .A2(n15783), .ZN(n6597) );
  INV_X1 U9562 ( .A(n11055), .ZN(n8966) );
  NAND2_X1 U9563 ( .A1(n9396), .A2(n12745), .ZN(n6598) );
  AND2_X1 U9564 ( .A1(n6577), .A2(n7589), .ZN(n6599) );
  INV_X1 U9565 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7279) );
  NAND2_X1 U9566 ( .A1(n12560), .A2(n10366), .ZN(n10643) );
  AND3_X1 U9567 ( .A1(n7475), .A2(n7473), .A3(n7474), .ZN(n6600) );
  INV_X1 U9568 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n12249) );
  NAND2_X1 U9569 ( .A1(n13207), .A2(n12823), .ZN(n13010) );
  INV_X1 U9570 ( .A(n13010), .ZN(n7771) );
  AND2_X1 U9571 ( .A1(n8278), .A2(n8277), .ZN(n15502) );
  AND2_X1 U9572 ( .A1(n7495), .A2(n7493), .ZN(n6601) );
  INV_X1 U9573 ( .A(n12619), .ZN(n7674) );
  OR2_X1 U9574 ( .A1(n14225), .A2(n14425), .ZN(n6602) );
  OR2_X1 U9575 ( .A1(n9724), .A2(n9723), .ZN(n6603) );
  NAND2_X1 U9576 ( .A1(n7109), .A2(n10516), .ZN(n14334) );
  AND2_X1 U9577 ( .A1(n9592), .A2(n7624), .ZN(n6604) );
  AND3_X1 U9578 ( .A1(n13864), .A2(n13863), .A3(n7717), .ZN(n6605) );
  AND2_X1 U9579 ( .A1(n7058), .A2(n7055), .ZN(n6606) );
  NOR2_X1 U9580 ( .A1(n14205), .A2(n14652), .ZN(n6607) );
  AND2_X1 U9581 ( .A1(n10516), .A2(n10528), .ZN(n6608) );
  INV_X1 U9582 ( .A(n11202), .ZN(n7624) );
  INV_X1 U9583 ( .A(n14984), .ZN(n14983) );
  NAND2_X1 U9584 ( .A1(n8778), .A2(n8777), .ZN(n14984) );
  AND4_X1 U9585 ( .A1(n8227), .A2(n8226), .A3(n8225), .A4(n8224), .ZN(n11564)
         );
  INV_X1 U9586 ( .A(n11564), .ZN(n14852) );
  AND2_X1 U9587 ( .A1(n14573), .A2(n14418), .ZN(n6609) );
  AND2_X1 U9588 ( .A1(n7960), .A2(n6940), .ZN(n6610) );
  OR2_X1 U9589 ( .A1(n14284), .A2(n13671), .ZN(n6611) );
  OR2_X1 U9590 ( .A1(n14316), .A2(n13909), .ZN(n6612) );
  AOI21_X1 U9591 ( .B1(n7093), .B2(n13334), .A(n7091), .ZN(n7090) );
  AND2_X1 U9592 ( .A1(n8255), .A2(n8256), .ZN(n6613) );
  NOR2_X1 U9593 ( .A1(n9089), .A2(n9111), .ZN(n6614) );
  AND2_X1 U9594 ( .A1(n7398), .A2(n7397), .ZN(n6615) );
  OR2_X1 U9595 ( .A1(n13511), .A2(n12868), .ZN(n13015) );
  INV_X1 U9596 ( .A(n13015), .ZN(n7238) );
  OR2_X1 U9597 ( .A1(n12728), .A2(n12801), .ZN(n12998) );
  INV_X1 U9598 ( .A(n12998), .ZN(n7925) );
  NAND2_X1 U9599 ( .A1(n12991), .A2(n7088), .ZN(n6616) );
  AND2_X1 U9600 ( .A1(n13899), .A2(n13898), .ZN(n6617) );
  NAND2_X1 U9601 ( .A1(n7723), .A2(n13891), .ZN(n6618) );
  AND2_X1 U9602 ( .A1(n7738), .A2(n7741), .ZN(n6619) );
  AND2_X1 U9603 ( .A1(n9528), .A2(n12998), .ZN(n6620) );
  AND2_X1 U9604 ( .A1(n7334), .A2(n9216), .ZN(n6621) );
  INV_X1 U9605 ( .A(n7584), .ZN(n7583) );
  NAND2_X1 U9606 ( .A1(n12947), .A2(n7585), .ZN(n7584) );
  OR2_X1 U9607 ( .A1(n9739), .A2(n9738), .ZN(n6622) );
  OR2_X1 U9608 ( .A1(n8376), .A2(SI_9_), .ZN(n6624) );
  INV_X1 U9609 ( .A(n6526), .ZN(n7439) );
  NAND2_X1 U9610 ( .A1(n13950), .A2(n13949), .ZN(n6625) );
  AND2_X1 U9611 ( .A1(n10463), .A2(n10455), .ZN(n6626) );
  NOR2_X1 U9612 ( .A1(n14511), .A2(n13993), .ZN(n6627) );
  INV_X1 U9613 ( .A(n8050), .ZN(n15039) );
  NAND2_X1 U9614 ( .A1(n8825), .A2(n8955), .ZN(n8050) );
  AND2_X1 U9615 ( .A1(n8936), .A2(n8933), .ZN(n6628) );
  INV_X1 U9616 ( .A(n7913), .ZN(n6919) );
  OAI21_X1 U9617 ( .B1(n7988), .B2(n7914), .A(n6611), .ZN(n7913) );
  AND2_X1 U9618 ( .A1(n6804), .A2(n6802), .ZN(n6629) );
  NAND2_X1 U9619 ( .A1(n8164), .A2(n8162), .ZN(n6630) );
  AND2_X1 U9620 ( .A1(n9143), .A2(n9142), .ZN(n6631) );
  AND3_X1 U9621 ( .A1(n9044), .A2(n9043), .A3(n9042), .ZN(n6632) );
  INV_X1 U9622 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n6734) );
  INV_X1 U9623 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7658) );
  OAI21_X1 U9624 ( .B1(n6571), .B2(n8048), .A(n12001), .ZN(n8047) );
  AND4_X1 U9625 ( .A1(n10385), .A2(n10384), .A3(n10383), .A4(n10382), .ZN(
        n10389) );
  NAND2_X1 U9626 ( .A1(n14660), .A2(n10321), .ZN(n12698) );
  INV_X1 U9627 ( .A(n12698), .ZN(n10366) );
  OR2_X1 U9628 ( .A1(n12893), .A2(n13504), .ZN(n6633) );
  NOR3_X1 U9629 ( .A1(n12954), .A2(n13011), .A3(n13421), .ZN(n6634) );
  AND2_X1 U9630 ( .A1(n7252), .A2(n13206), .ZN(n6635) );
  NAND2_X1 U9631 ( .A1(n8204), .A2(n8203), .ZN(n15284) );
  INV_X1 U9632 ( .A(n15284), .ZN(n7840) );
  OR2_X1 U9633 ( .A1(n12956), .A2(n12957), .ZN(n6636) );
  AND2_X1 U9634 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_REG3_REG_6__SCAN_IN), 
        .ZN(n6637) );
  NOR2_X1 U9635 ( .A1(n14724), .A2(n15258), .ZN(n6638) );
  NOR2_X1 U9636 ( .A1(n14788), .A2(n15226), .ZN(n6639) );
  NOR2_X1 U9637 ( .A1(n14539), .A2(n13729), .ZN(n6640) );
  NOR2_X1 U9638 ( .A1(n9823), .A2(n12810), .ZN(n6641) );
  OR2_X1 U9639 ( .A1(n14329), .A2(n14340), .ZN(n6642) );
  XOR2_X1 U9640 ( .A(n9774), .B(n9773), .Z(n6643) );
  OR2_X1 U9641 ( .A1(n14184), .A2(n14196), .ZN(n14191) );
  INV_X1 U9642 ( .A(n8628), .ZN(n7466) );
  AND2_X1 U9643 ( .A1(n8486), .A2(n8485), .ZN(n6644) );
  XNOR2_X1 U9644 ( .A(n8146), .B(SI_8_), .ZN(n8346) );
  AND2_X1 U9645 ( .A1(n7464), .A2(n7461), .ZN(n6645) );
  NAND2_X1 U9646 ( .A1(n10711), .A2(n10584), .ZN(n14058) );
  INV_X1 U9647 ( .A(n14058), .ZN(n8000) );
  AOI21_X1 U9648 ( .B1(n7703), .B2(n7705), .A(n7702), .ZN(n7701) );
  INV_X1 U9649 ( .A(n13356), .ZN(n7066) );
  AND2_X1 U9650 ( .A1(n8950), .A2(n8949), .ZN(n6646) );
  NOR2_X1 U9651 ( .A1(n13523), .A2(n12801), .ZN(n6647) );
  NAND2_X1 U9652 ( .A1(n9258), .A2(n6599), .ZN(n6648) );
  INV_X1 U9653 ( .A(n7661), .ZN(n7660) );
  NAND2_X1 U9654 ( .A1(n7663), .A2(n7662), .ZN(n7661) );
  INV_X1 U9655 ( .A(n7861), .ZN(n7860) );
  NAND2_X1 U9656 ( .A1(n15107), .A2(n15090), .ZN(n7861) );
  INV_X1 U9657 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10886) );
  OR2_X1 U9658 ( .A1(n9696), .A2(n12335), .ZN(n6649) );
  INV_X1 U9659 ( .A(n7824), .ZN(n7823) );
  OAI21_X1 U9660 ( .B1(n6589), .B2(n7825), .A(n8176), .ZN(n7824) );
  AND2_X1 U9661 ( .A1(n9203), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n6650) );
  AND2_X1 U9662 ( .A1(n8951), .A2(n8942), .ZN(n6651) );
  INV_X1 U9663 ( .A(n7225), .ZN(n7224) );
  NAND2_X1 U9664 ( .A1(n12131), .A2(n12598), .ZN(n7225) );
  NOR2_X1 U9665 ( .A1(n15330), .A2(n15116), .ZN(n6652) );
  NAND2_X1 U9666 ( .A1(n13196), .A2(n13195), .ZN(n6653) );
  OR2_X1 U9667 ( .A1(n7465), .A2(n7466), .ZN(n6654) );
  AND2_X1 U9668 ( .A1(n13369), .A2(n6636), .ZN(n6655) );
  NAND2_X1 U9669 ( .A1(n9822), .A2(n12774), .ZN(n6656) );
  INV_X1 U9670 ( .A(n7984), .ZN(n7983) );
  NAND2_X1 U9671 ( .A1(n7988), .A2(n7990), .ZN(n7984) );
  INV_X1 U9672 ( .A(n8072), .ZN(n8007) );
  AND2_X1 U9673 ( .A1(n6551), .A2(n6576), .ZN(n6657) );
  INV_X1 U9674 ( .A(n7013), .ZN(n7011) );
  NAND2_X1 U9675 ( .A1(n7014), .A2(n6624), .ZN(n7013) );
  NAND2_X1 U9676 ( .A1(n10197), .A2(n7690), .ZN(n13843) );
  AND2_X1 U9677 ( .A1(n7887), .A2(n14374), .ZN(n6658) );
  OR2_X1 U9678 ( .A1(n9529), .A2(n7923), .ZN(n6659) );
  OR2_X1 U9679 ( .A1(n7083), .A2(n7082), .ZN(n6660) );
  AND2_X1 U9680 ( .A1(n8105), .A2(n8104), .ZN(n8205) );
  AND2_X1 U9681 ( .A1(n7784), .A2(n7781), .ZN(n6661) );
  OR2_X1 U9682 ( .A1(n13201), .A2(n13196), .ZN(n12866) );
  INV_X1 U9683 ( .A(n8891), .ZN(n12001) );
  AND2_X1 U9684 ( .A1(n6798), .A2(n9384), .ZN(n6662) );
  INV_X1 U9685 ( .A(n7422), .ZN(n7421) );
  NAND2_X1 U9686 ( .A1(n7425), .A2(n9669), .ZN(n7422) );
  INV_X1 U9687 ( .A(n8827), .ZN(n11581) );
  OR2_X1 U9688 ( .A1(n14029), .A2(n7986), .ZN(n6663) );
  INV_X1 U9689 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n15422) );
  INV_X1 U9690 ( .A(n11660), .ZN(n7069) );
  INV_X1 U9691 ( .A(n8425), .ZN(n7457) );
  INV_X1 U9692 ( .A(n8617), .ZN(n7178) );
  INV_X1 U9693 ( .A(n8342), .ZN(n7189) );
  NOR2_X1 U9694 ( .A1(n15581), .A2(n14848), .ZN(n6664) );
  INV_X1 U9695 ( .A(n13893), .ZN(n7724) );
  OR2_X1 U9696 ( .A1(n13884), .A2(n13886), .ZN(n6665) );
  AND3_X1 U9697 ( .A1(n7474), .A2(n8205), .A3(n8106), .ZN(n6666) );
  OR2_X1 U9698 ( .A1(n13538), .A2(n13323), .ZN(n12983) );
  OR2_X1 U9699 ( .A1(n13598), .A2(n13423), .ZN(n12943) );
  AND2_X1 U9700 ( .A1(n12124), .A2(n12123), .ZN(n6667) );
  OR2_X1 U9701 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n9705), .ZN(n6668) );
  AND2_X1 U9702 ( .A1(n7782), .A2(n7781), .ZN(n6669) );
  AND2_X1 U9703 ( .A1(n7336), .A2(n7335), .ZN(n6670) );
  AND2_X1 U9704 ( .A1(n7557), .A2(n6559), .ZN(n6671) );
  AND2_X1 U9705 ( .A1(n12672), .A2(n13798), .ZN(n6672) );
  NAND2_X1 U9706 ( .A1(n10291), .A2(n10290), .ZN(n14517) );
  INV_X1 U9707 ( .A(n14517), .ZN(n14234) );
  OR2_X1 U9708 ( .A1(n12205), .A2(n13402), .ZN(n6673) );
  INV_X1 U9709 ( .A(n10653), .ZN(n10659) );
  XNOR2_X1 U9710 ( .A(n14837), .B(n15284), .ZN(n10653) );
  OR2_X1 U9711 ( .A1(n10628), .A2(n10629), .ZN(n6674) );
  NOR3_X1 U9712 ( .A1(n8912), .A2(n7556), .A3(n8840), .ZN(n6675) );
  AND2_X1 U9713 ( .A1(n8143), .A2(SI_7_), .ZN(n6676) );
  AND2_X1 U9714 ( .A1(n6576), .A2(n12941), .ZN(n6677) );
  NOR2_X1 U9715 ( .A1(n15396), .A2(n14847), .ZN(n6678) );
  NOR2_X1 U9716 ( .A1(n9972), .A2(n7765), .ZN(n7764) );
  AND2_X1 U9717 ( .A1(n12932), .A2(n12933), .ZN(n12930) );
  NOR2_X1 U9718 ( .A1(n7452), .A2(n7178), .ZN(n6679) );
  AND2_X1 U9719 ( .A1(n10224), .A2(n7652), .ZN(n6680) );
  AND2_X1 U9720 ( .A1(n6887), .A2(n6886), .ZN(n6681) );
  AND2_X1 U9721 ( .A1(n13215), .A2(n13008), .ZN(n6682) );
  AND2_X1 U9722 ( .A1(n14011), .A2(n7345), .ZN(n6683) );
  INV_X1 U9723 ( .A(n7550), .ZN(n6965) );
  NOR2_X1 U9724 ( .A1(n6572), .A2(n7551), .ZN(n7550) );
  NAND2_X1 U9725 ( .A1(n10087), .A2(n7002), .ZN(n7007) );
  AND2_X1 U9726 ( .A1(n7429), .A2(n7424), .ZN(n6684) );
  AND2_X1 U9727 ( .A1(n7840), .A2(n15020), .ZN(n6685) );
  AND2_X1 U9728 ( .A1(n8069), .A2(n7286), .ZN(n6686) );
  AND2_X1 U9729 ( .A1(n8070), .A2(n7284), .ZN(n6687) );
  OR2_X1 U9730 ( .A1(n8437), .A2(n8439), .ZN(n6688) );
  AND2_X1 U9731 ( .A1(n6550), .A2(n6923), .ZN(n6689) );
  INV_X1 U9732 ( .A(n10481), .ZN(n7977) );
  NAND2_X1 U9733 ( .A1(n6663), .A2(n7990), .ZN(n7982) );
  AND2_X1 U9734 ( .A1(n7556), .A2(n8050), .ZN(n6690) );
  AND2_X1 U9735 ( .A1(n13263), .A2(n6598), .ZN(n7154) );
  INV_X1 U9736 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n10267) );
  INV_X1 U9737 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n10311) );
  OR2_X1 U9738 ( .A1(n10045), .A2(n10044), .ZN(n6691) );
  AND2_X1 U9739 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), .ZN(
        n6692) );
  AND2_X1 U9740 ( .A1(n9810), .A2(n7962), .ZN(n7961) );
  INV_X1 U9741 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9118) );
  INV_X1 U9742 ( .A(n7434), .ZN(n7433) );
  NAND2_X1 U9743 ( .A1(n7437), .A2(n7435), .ZN(n7434) );
  INV_X1 U9744 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n10306) );
  INV_X1 U9745 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n12308) );
  INV_X1 U9746 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n8144) );
  INV_X1 U9747 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n9026) );
  INV_X1 U9748 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6923) );
  INV_X1 U9749 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n10168) );
  INV_X1 U9750 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7971) );
  INV_X1 U9751 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10912) );
  NAND2_X1 U9752 ( .A1(n7631), .A2(n11055), .ZN(n7633) );
  INV_X1 U9753 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10840) );
  OR2_X1 U9754 ( .A1(n10674), .A2(n10673), .ZN(P1_U3266) );
  INV_X1 U9755 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n12482) );
  AND2_X2 U9756 ( .A1(n10359), .A2(n15792), .ZN(n15838) );
  INV_X1 U9757 ( .A(n15838), .ZN(n7304) );
  INV_X1 U9758 ( .A(n9384), .ZN(n6797) );
  NOR2_X1 U9759 ( .A1(n15262), .A2(n15360), .ZN(n7490) );
  INV_X1 U9760 ( .A(n15848), .ZN(n7285) );
  NAND2_X1 U9761 ( .A1(n6832), .A2(n12943), .ZN(n13415) );
  INV_X1 U9762 ( .A(n10173), .ZN(n10269) );
  NAND2_X1 U9763 ( .A1(n9554), .A2(n9553), .ZN(n9557) );
  NAND2_X1 U9764 ( .A1(n9462), .A2(n9461), .ZN(n13207) );
  NAND2_X1 U9765 ( .A1(n7148), .A2(n8436), .ZN(n14724) );
  INV_X1 U9766 ( .A(n14652), .ZN(n7368) );
  XNOR2_X1 U9767 ( .A(n8811), .B(P1_IR_REG_25__SCAN_IN), .ZN(n8979) );
  INV_X1 U9768 ( .A(n8971), .ZN(n11828) );
  AND2_X1 U9769 ( .A1(n14480), .A2(n14653), .ZN(n14457) );
  AND2_X1 U9770 ( .A1(n11797), .A2(n15824), .ZN(n11936) );
  NAND2_X1 U9771 ( .A1(n10167), .A2(n10232), .ZN(n10335) );
  INV_X2 U9772 ( .A(n15781), .ZN(n15783) );
  INV_X1 U9773 ( .A(n13902), .ZN(n7712) );
  INV_X1 U9774 ( .A(n15330), .ZN(n7851) );
  INV_X1 U9775 ( .A(n7620), .ZN(n13047) );
  NAND2_X1 U9776 ( .A1(n7383), .A2(n10903), .ZN(n7620) );
  OAI211_X1 U9777 ( .C1(n6817), .C2(n6822), .A(n12928), .B(n6815), .ZN(n12089)
         );
  NAND2_X1 U9778 ( .A1(n10429), .A2(n7110), .ZN(n12025) );
  INV_X1 U9779 ( .A(n9775), .ZN(n9777) );
  INV_X1 U9780 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7796) );
  INV_X1 U9781 ( .A(n15733), .ZN(n15744) );
  NAND2_X1 U9782 ( .A1(n6827), .A2(n6829), .ZN(n13388) );
  NAND2_X1 U9783 ( .A1(n7865), .A2(n12932), .ZN(n11943) );
  NAND2_X1 U9784 ( .A1(n7895), .A2(n9511), .ZN(n11692) );
  NAND2_X1 U9785 ( .A1(n7874), .A2(n9512), .ZN(n13404) );
  AND2_X1 U9786 ( .A1(n9216), .A2(n9204), .ZN(n6694) );
  OR2_X1 U9787 ( .A1(n15905), .A2(n13510), .ZN(n6695) );
  NAND2_X1 U9788 ( .A1(n12016), .A2(n10591), .ZN(n11794) );
  NAND2_X1 U9789 ( .A1(n8025), .A2(n8888), .ZN(n11672) );
  NAND2_X1 U9790 ( .A1(n8023), .A2(n8024), .ZN(n11838) );
  NOR2_X1 U9791 ( .A1(n13071), .A2(n7407), .ZN(n13089) );
  INV_X1 U9792 ( .A(n13089), .ZN(n7406) );
  NAND2_X2 U9793 ( .A1(n11390), .A2(n15259), .ZN(n15232) );
  INV_X1 U9794 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n9700) );
  INV_X1 U9795 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n12476) );
  AND2_X1 U9796 ( .A1(n7122), .A2(n13045), .ZN(n6696) );
  NOR2_X1 U9797 ( .A1(n13066), .A2(n13394), .ZN(n13086) );
  AND3_X1 U9798 ( .A1(n9012), .A2(n9011), .A3(n9010), .ZN(n9218) );
  AND2_X1 U9799 ( .A1(n7808), .A2(n9409), .ZN(n6697) );
  OR2_X1 U9800 ( .A1(n8195), .A2(SI_25_), .ZN(n6698) );
  AND2_X1 U9801 ( .A1(n9250), .A2(n7042), .ZN(n6699) );
  INV_X1 U9802 ( .A(n14356), .ZN(n7113) );
  NAND2_X1 U9803 ( .A1(n8691), .A2(n8690), .ZN(n15032) );
  NAND2_X1 U9804 ( .A1(n9423), .A2(n9422), .ZN(n13259) );
  AND2_X1 U9805 ( .A1(n13992), .A2(n7368), .ZN(n6700) );
  AND2_X1 U9806 ( .A1(n10098), .A2(n7024), .ZN(n6701) );
  OR2_X1 U9807 ( .A1(n11996), .A2(n15384), .ZN(n6702) );
  INV_X1 U9808 ( .A(n14724), .ZN(n7847) );
  AND2_X1 U9809 ( .A1(n7423), .A2(n7421), .ZN(n6703) );
  AND2_X1 U9810 ( .A1(n6897), .A2(n6896), .ZN(n6704) );
  INV_X1 U9811 ( .A(n6893), .ZN(n6892) );
  AND2_X1 U9812 ( .A1(n7041), .A2(n7040), .ZN(n6705) );
  NAND2_X1 U9813 ( .A1(n10872), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6706) );
  AND2_X1 U9814 ( .A1(n7285), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6707) );
  NOR2_X1 U9815 ( .A1(n13052), .A2(n9596), .ZN(n6708) );
  AND2_X1 U9816 ( .A1(n11830), .A2(n8927), .ZN(n6709) );
  INV_X1 U9817 ( .A(n7499), .ZN(n7498) );
  NAND2_X1 U9818 ( .A1(n14149), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7499) );
  INV_X1 U9819 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8446) );
  OR2_X1 U9820 ( .A1(n9627), .A2(n7518), .ZN(n6710) );
  INV_X1 U9821 ( .A(SI_14_), .ZN(n11044) );
  OR2_X1 U9822 ( .A1(n11232), .A2(n7506), .ZN(n6711) );
  NAND2_X1 U9823 ( .A1(n13562), .A2(n13373), .ZN(n6712) );
  AND2_X1 U9824 ( .A1(n11873), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6713) );
  INV_X1 U9825 ( .A(n14217), .ZN(n14619) );
  INV_X1 U9826 ( .A(n12963), .ZN(n12968) );
  AND2_X1 U9827 ( .A1(n13562), .A2(n12774), .ZN(n12963) );
  INV_X1 U9828 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n12251) );
  OR2_X1 U9829 ( .A1(n14511), .A2(n13733), .ZN(n6714) );
  INV_X1 U9830 ( .A(n9826), .ZN(n7944) );
  INV_X1 U9831 ( .A(n12745), .ZN(n13289) );
  AND2_X1 U9832 ( .A1(n9395), .A2(n9394), .ZN(n12745) );
  AND2_X1 U9833 ( .A1(n7748), .A2(n7747), .ZN(n6715) );
  OAI21_X1 U9834 ( .B1(n13055), .B2(n6553), .A(n6710), .ZN(n7516) );
  INV_X1 U9835 ( .A(n7935), .ZN(n7934) );
  INV_X1 U9836 ( .A(n9892), .ZN(n8262) );
  INV_X1 U9837 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6971) );
  NAND2_X1 U9838 ( .A1(n10272), .A2(n10271), .ZN(n14364) );
  INV_X1 U9839 ( .A(n14364), .ZN(n7662) );
  NAND4_X1 U9840 ( .A1(n9062), .A2(n9061), .A3(n9060), .A4(n9059), .ZN(n13041)
         );
  INV_X1 U9841 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7735) );
  NAND2_X1 U9842 ( .A1(n8422), .A2(n8421), .ZN(n15384) );
  INV_X1 U9843 ( .A(n15384), .ZN(n7846) );
  NAND2_X2 U9844 ( .A1(n10184), .A2(n10878), .ZN(n10292) );
  NAND2_X1 U9845 ( .A1(n9114), .A2(n7070), .ZN(n13038) );
  INV_X1 U9846 ( .A(n13038), .ZN(n6952) );
  NAND2_X1 U9847 ( .A1(n7621), .A2(n11202), .ZN(n11179) );
  NAND2_X1 U9848 ( .A1(n7736), .A2(n9908), .ZN(n15495) );
  OR2_X1 U9849 ( .A1(n9680), .A2(n13360), .ZN(n6716) );
  NAND2_X1 U9850 ( .A1(n11699), .A2(n12895), .ZN(n13023) );
  INV_X1 U9851 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6931) );
  INV_X1 U9852 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6972) );
  OR2_X1 U9853 ( .A1(P3_ADDR_REG_11__SCAN_IN), .A2(n12257), .ZN(n6717) );
  NAND2_X1 U9854 ( .A1(n12039), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6718) );
  NAND2_X1 U9855 ( .A1(n7436), .A2(n7433), .ZN(n7432) );
  AND2_X1 U9856 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n7803), .ZN(n6719) );
  INV_X1 U9857 ( .A(n12801), .ZN(n13274) );
  AND2_X1 U9858 ( .A1(n14479), .A2(n13811), .ZN(n15817) );
  INV_X1 U9859 ( .A(n15545), .ZN(n15360) );
  INV_X1 U9860 ( .A(n15163), .ZN(n15199) );
  INV_X1 U9861 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7506) );
  OR2_X1 U9862 ( .A1(n9680), .A2(n9679), .ZN(n6720) );
  INV_X1 U9863 ( .A(n10350), .ZN(n14176) );
  OR2_X1 U9864 ( .A1(n8109), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n6721) );
  NAND2_X1 U9865 ( .A1(n11753), .A2(n9571), .ZN(n13024) );
  AND2_X1 U9866 ( .A1(n14078), .A2(n14069), .ZN(n6722) );
  AND2_X1 U9867 ( .A1(n7520), .A2(n7519), .ZN(n6723) );
  AND2_X1 U9868 ( .A1(n6740), .A2(n6745), .ZN(n6724) );
  AND2_X1 U9869 ( .A1(n11603), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n6725) );
  NAND2_X1 U9870 ( .A1(n9621), .A2(n10833), .ZN(n6726) );
  INV_X1 U9871 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n9075) );
  INV_X1 U9872 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7274) );
  INV_X1 U9873 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n7390) );
  INV_X1 U9874 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7881) );
  INV_X1 U9875 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7878) );
  INV_X1 U9876 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6748) );
  INV_X1 U9877 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7270) );
  INV_X1 U9878 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7693) );
  INV_X1 U9879 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7803) );
  INV_X1 U9880 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7320) );
  INV_X1 U9881 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6813) );
  INV_X1 U9882 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7568) );
  INV_X1 U9883 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n7535) );
  INV_X1 U9884 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10847) );
  NAND2_X1 U9885 ( .A1(n8043), .A2(n8042), .ZN(n15222) );
  NAND2_X1 U9886 ( .A1(n11562), .A2(n11563), .ZN(n8062) );
  OAI21_X2 U9887 ( .B1(n8201), .B2(n7279), .A(n7276), .ZN(n15433) );
  OAI211_X1 U9888 ( .C1(n7038), .C2(n13101), .A(n13181), .B(n6727), .ZN(
        P3_U3201) );
  NAND3_X1 U9889 ( .A1(n6731), .A2(n9598), .A3(n6730), .ZN(n13084) );
  NAND2_X1 U9890 ( .A1(n7357), .A2(n7518), .ZN(n6732) );
  NAND3_X1 U9891 ( .A1(n11151), .A2(n11152), .A3(n11202), .ZN(n6733) );
  NAND2_X1 U9892 ( .A1(n11179), .A2(n11197), .ZN(n7356) );
  NAND3_X1 U9893 ( .A1(n7134), .A2(n7133), .A3(n9601), .ZN(n7131) );
  NAND3_X1 U9894 ( .A1(n7132), .A2(n7626), .A3(n7131), .ZN(n7629) );
  NAND3_X1 U9895 ( .A1(n6743), .A2(n6585), .A3(n6744), .ZN(n6741) );
  INV_X1 U9896 ( .A(n15928), .ZN(n6743) );
  INV_X1 U9897 ( .A(n6750), .ZN(n9742) );
  XNOR2_X1 U9898 ( .A(n9739), .B(n9738), .ZN(n15926) );
  NAND2_X1 U9899 ( .A1(n7181), .A2(n7183), .ZN(n15467) );
  INV_X1 U9900 ( .A(n15444), .ZN(n7333) );
  NAND3_X1 U9901 ( .A1(n9746), .A2(n6549), .A3(n9747), .ZN(n6754) );
  NAND2_X1 U9902 ( .A1(n15463), .A2(n15464), .ZN(n6755) );
  NAND4_X1 U9903 ( .A1(n10232), .A2(n10167), .A3(n10168), .A4(n7652), .ZN(
        n6757) );
  XNOR2_X2 U9904 ( .A(n6758), .B(n10168), .ZN(n14669) );
  NOR2_X2 U9905 ( .A1(n12054), .A2(n6759), .ZN(n14480) );
  XNOR2_X1 U9906 ( .A(n6760), .B(n10174), .ZN(n10350) );
  INV_X1 U9907 ( .A(n14413), .ZN(n6765) );
  NAND2_X1 U9908 ( .A1(n6772), .A2(n6771), .ZN(n6770) );
  NOR2_X2 U9909 ( .A1(n14294), .A2(n14284), .ZN(n14283) );
  NAND2_X1 U9910 ( .A1(n6781), .A2(n13895), .ZN(n13899) );
  NAND4_X1 U9911 ( .A1(n7721), .A2(n6782), .A3(n6783), .A4(n6784), .ZN(n6781)
         );
  OR2_X1 U9912 ( .A1(n13888), .A2(n6618), .ZN(n6784) );
  NAND3_X1 U9913 ( .A1(n7721), .A2(n6784), .A3(n6783), .ZN(n13897) );
  NAND3_X1 U9914 ( .A1(n11905), .A2(n15806), .A3(n11977), .ZN(n12013) );
  NOR2_X2 U9915 ( .A1(n11976), .A2(n13813), .ZN(n11977) );
  NAND2_X1 U9916 ( .A1(n11364), .A2(n13820), .ZN(n11976) );
  NAND3_X1 U9917 ( .A1(n6796), .A2(n6795), .A3(n7154), .ZN(n6794) );
  NAND2_X1 U9918 ( .A1(n9314), .A2(n7602), .ZN(n6795) );
  AOI21_X1 U9919 ( .B1(n7602), .B2(n7605), .A(n6662), .ZN(n6796) );
  NAND2_X1 U9920 ( .A1(n6669), .A2(n9117), .ZN(n6805) );
  INV_X1 U9921 ( .A(n9186), .ZN(n9188) );
  NAND2_X1 U9922 ( .A1(n6801), .A2(n6805), .ZN(n6800) );
  NAND2_X1 U9923 ( .A1(n7774), .A2(n6807), .ZN(n6806) );
  NAND2_X1 U9924 ( .A1(n6822), .A2(n6820), .ZN(n6819) );
  NAND2_X1 U9925 ( .A1(n7890), .A2(n6816), .ZN(n6815) );
  NAND2_X1 U9926 ( .A1(n7890), .A2(n12924), .ZN(n6817) );
  NOR2_X1 U9927 ( .A1(n7894), .A2(n6818), .ZN(n6820) );
  OR2_X1 U9928 ( .A1(n12922), .A2(n6821), .ZN(n6818) );
  INV_X1 U9929 ( .A(n12876), .ZN(n15857) );
  NAND2_X1 U9930 ( .A1(n6823), .A2(n12903), .ZN(n11476) );
  AND2_X2 U9931 ( .A1(n12903), .A2(n12909), .ZN(n12876) );
  NAND2_X1 U9932 ( .A1(n12147), .A2(n6828), .ZN(n6827) );
  AOI21_X2 U9933 ( .B1(n10678), .B2(n15864), .A(n6833), .ZN(n13214) );
  NAND2_X1 U9934 ( .A1(n6834), .A2(n10681), .ZN(n6833) );
  NAND2_X1 U9935 ( .A1(n10679), .A2(n12150), .ZN(n6834) );
  NAND2_X1 U9936 ( .A1(n10676), .A2(n7245), .ZN(n10679) );
  NAND2_X1 U9937 ( .A1(n13295), .A2(n6835), .ZN(n6839) );
  NAND3_X1 U9938 ( .A1(n6839), .A2(n7871), .A3(n6837), .ZN(n9527) );
  NAND2_X1 U9939 ( .A1(n7869), .A2(n6838), .ZN(n6837) );
  INV_X1 U9940 ( .A(n9524), .ZN(n6838) );
  NAND2_X2 U9941 ( .A1(n9503), .A2(n13612), .ZN(n9047) );
  NAND2_X2 U9942 ( .A1(n9047), .A2(n10879), .ZN(n9064) );
  NAND2_X1 U9943 ( .A1(n9047), .A2(n10878), .ZN(n9069) );
  NAND2_X1 U9944 ( .A1(n8504), .A2(n6845), .ZN(n11658) );
  NAND3_X1 U9945 ( .A1(n6850), .A2(n6849), .A3(n15064), .ZN(n6848) );
  NAND3_X1 U9946 ( .A1(n14700), .A2(n6582), .A3(n14803), .ZN(n6852) );
  NAND2_X1 U9947 ( .A1(n14804), .A2(n6853), .ZN(n7760) );
  NAND2_X1 U9948 ( .A1(n7761), .A2(n6853), .ZN(n14699) );
  NAND2_X1 U9949 ( .A1(n7012), .A2(n7011), .ZN(n6858) );
  OAI21_X2 U9950 ( .B1(n7012), .B2(n6574), .A(n6856), .ZN(n8434) );
  NAND2_X1 U9951 ( .A1(n8434), .A2(n8086), .ZN(n8158) );
  MUX2_X1 U9952 ( .A(n10840), .B(n12482), .S(n8125), .Z(n8126) );
  NAND2_X1 U9953 ( .A1(n6868), .A2(n6869), .ZN(n8469) );
  INV_X1 U9954 ( .A(n8519), .ZN(n6866) );
  OAI21_X1 U9955 ( .B1(n15615), .B2(n6876), .A(n15628), .ZN(n6875) );
  NAND4_X1 U9956 ( .A1(n6884), .A2(n6879), .A3(n6878), .A4(n6877), .ZN(
        P2_U3233) );
  NAND2_X1 U9957 ( .A1(n6888), .A2(n6681), .ZN(n6878) );
  OAI22_X1 U9958 ( .A1(n14175), .A2(n6882), .B1(n6887), .B2(n6881), .ZN(n6880)
         );
  NAND2_X1 U9959 ( .A1(n15745), .A2(n6548), .ZN(n6887) );
  INV_X1 U9960 ( .A(n6889), .ZN(n6888) );
  INV_X1 U9961 ( .A(n6891), .ZN(n15685) );
  NOR2_X1 U9962 ( .A1(n11263), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6893) );
  OAI21_X1 U9963 ( .B1(n14140), .B2(n6895), .A(n6894), .ZN(n14141) );
  XNOR2_X1 U9964 ( .A(n14141), .B(n14155), .ZN(n15718) );
  NAND2_X1 U9965 ( .A1(n10592), .A2(n7904), .ZN(n7903) );
  NAND2_X2 U9966 ( .A1(n10366), .A2(n6907), .ZN(n7879) );
  NAND2_X1 U9967 ( .A1(n14358), .A2(n6908), .ZN(n6910) );
  INV_X1 U9968 ( .A(n10614), .ZN(n6909) );
  NAND2_X1 U9969 ( .A1(n6910), .A2(n6911), .ZN(n14320) );
  NAND2_X1 U9970 ( .A1(n11339), .A2(n14035), .ZN(n11966) );
  XNOR2_X1 U9971 ( .A(n13816), .B(n11364), .ZN(n14035) );
  NAND2_X1 U9972 ( .A1(n14305), .A2(n6595), .ZN(n6916) );
  NAND2_X1 U9973 ( .A1(n14243), .A2(n10630), .ZN(n6918) );
  NAND4_X1 U9974 ( .A1(n7117), .A2(n7115), .A3(n6550), .A4(
        P2_IR_REG_29__SCAN_IN), .ZN(n6920) );
  INV_X1 U9975 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6932) );
  NAND3_X1 U9976 ( .A1(n6935), .A2(n12832), .A3(n6934), .ZN(n12787) );
  NAND2_X1 U9977 ( .A1(n12780), .A2(n12779), .ZN(n6938) );
  NAND2_X1 U9978 ( .A1(n6936), .A2(n12780), .ZN(n12724) );
  INV_X1 U9979 ( .A(n12782), .ZN(n6937) );
  NAND2_X1 U9980 ( .A1(n7961), .A2(n11819), .ZN(n6939) );
  NAND2_X1 U9981 ( .A1(n9831), .A2(n9832), .ZN(n9833) );
  INV_X1 U9982 ( .A(n6945), .ZN(n12796) );
  NAND3_X1 U9983 ( .A1(n6942), .A2(n12745), .A3(n9833), .ZN(n6945) );
  INV_X1 U9984 ( .A(n9831), .ZN(n6944) );
  NAND2_X1 U9985 ( .A1(n12733), .A2(n7941), .ZN(n7937) );
  OAI22_X2 U9986 ( .A1(n12829), .A2(n6946), .B1(n6584), .B2(n6948), .ZN(n12733) );
  NAND3_X1 U9987 ( .A1(n11765), .A2(n11955), .A3(n6951), .ZN(n9795) );
  NAND3_X1 U9988 ( .A1(n9131), .A2(n6955), .A3(n9133), .ZN(n13037) );
  OAI21_X2 U9989 ( .B1(n8023), .B2(n6959), .A(n6958), .ZN(n11917) );
  AOI21_X1 U9990 ( .B1(n6960), .B2(n11839), .A(n6678), .ZN(n6958) );
  NAND2_X1 U9991 ( .A1(n11917), .A2(n8928), .ZN(n8890) );
  INV_X1 U9992 ( .A(n6962), .ZN(n6961) );
  OAI21_X1 U9993 ( .B1(n8900), .B2(n6965), .A(n7547), .ZN(n6962) );
  NAND2_X1 U9994 ( .A1(n15206), .A2(n6964), .ZN(n6963) );
  AND2_X1 U9995 ( .A1(n8895), .A2(n7550), .ZN(n6964) );
  NAND3_X1 U9996 ( .A1(n6975), .A2(n6974), .A3(n6973), .ZN(P2_U3237) );
  OR2_X1 U9997 ( .A1(n14201), .A2(n14421), .ZN(n6973) );
  NAND2_X1 U9998 ( .A1(n7326), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n10529) );
  NAND3_X1 U9999 ( .A1(n10361), .A2(n6532), .A3(P2_REG3_REG_7__SCAN_IN), .ZN(
        n10431) );
  NAND3_X1 U10000 ( .A1(n6986), .A2(n8191), .A3(n6984), .ZN(n8647) );
  NAND2_X1 U10001 ( .A1(n7817), .A2(n6985), .ZN(n6984) );
  INV_X1 U10002 ( .A(n8189), .ZN(n6985) );
  NAND2_X1 U10003 ( .A1(n8187), .A2(n7817), .ZN(n6986) );
  OAI21_X2 U10004 ( .B1(n8591), .B2(n6991), .A(n6988), .ZN(n8186) );
  NAND2_X1 U10005 ( .A1(n9924), .A2(n6995), .ZN(n6994) );
  NAND2_X1 U10006 ( .A1(n6994), .A2(n6992), .ZN(n11515) );
  INV_X1 U10007 ( .A(n6993), .ZN(n6992) );
  OAI21_X1 U10008 ( .B1(n9924), .B2(n7000), .A(n6999), .ZN(n11356) );
  NOR2_X1 U10009 ( .A1(n9932), .A2(n6996), .ZN(n6995) );
  NAND2_X1 U10010 ( .A1(n7000), .A2(n6999), .ZN(n6998) );
  XNOR2_X1 U10011 ( .A(n7001), .B(n10111), .ZN(n9898) );
  AND2_X2 U10012 ( .A1(n6613), .A2(n8257), .ZN(n15535) );
  NAND2_X1 U10013 ( .A1(n10093), .A2(n10094), .ZN(n10097) );
  NAND3_X1 U10014 ( .A1(n10086), .A2(n10087), .A3(n7003), .ZN(n7002) );
  INV_X1 U10015 ( .A(n7007), .ZN(n7742) );
  INV_X1 U10016 ( .A(n7004), .ZN(n7741) );
  NAND2_X1 U10017 ( .A1(n10096), .A2(n10095), .ZN(n7005) );
  INV_X1 U10018 ( .A(n7743), .ZN(n7006) );
  NAND3_X1 U10019 ( .A1(n8326), .A2(n8145), .A3(n8142), .ZN(n7010) );
  NAND2_X1 U10020 ( .A1(n7214), .A2(n8141), .ZN(n8326) );
  NAND2_X1 U10021 ( .A1(n7010), .A2(n7008), .ZN(n7012) );
  INV_X1 U10022 ( .A(n11864), .ZN(n7018) );
  NAND2_X1 U10023 ( .A1(n7016), .A2(n7015), .ZN(n12163) );
  NAND2_X1 U10024 ( .A1(n11864), .A2(n7764), .ZN(n7015) );
  NAND2_X1 U10025 ( .A1(n7818), .A2(n7021), .ZN(n7019) );
  OAI21_X1 U10026 ( .B1(n7818), .B2(n7023), .A(n7021), .ZN(n8529) );
  NAND2_X1 U10027 ( .A1(n7019), .A2(n7020), .ZN(n7821) );
  NAND2_X1 U10028 ( .A1(n12162), .A2(n8650), .ZN(n7025) );
  NAND2_X1 U10029 ( .A1(n7026), .A2(n10079), .ZN(n10080) );
  INV_X4 U10030 ( .A(n8125), .ZN(n10878) );
  OAI21_X1 U10031 ( .B1(n8125), .B2(n10912), .A(n7027), .ZN(n8146) );
  NAND2_X1 U10032 ( .A1(n8125), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n7027) );
  XNOR2_X2 U10033 ( .A(n7030), .B(P3_IR_REG_4__SCAN_IN), .ZN(n11158) );
  OAI22_X2 U10034 ( .A1(n11736), .A2(n12462), .B1(n9662), .B2(n7031), .ZN(
        n11885) );
  INV_X1 U10035 ( .A(n7032), .ZN(n7031) );
  XNOR2_X2 U10036 ( .A(n7032), .B(n11740), .ZN(n11736) );
  OAI21_X1 U10037 ( .B1(n12108), .B2(n7037), .A(n7035), .ZN(n13053) );
  AOI21_X1 U10038 ( .B1(n9626), .B2(n13487), .A(n7036), .ZN(n7035) );
  INV_X1 U10039 ( .A(n9626), .ZN(n7037) );
  NAND3_X1 U10040 ( .A1(n7532), .A2(n7527), .A3(n7526), .ZN(n7525) );
  INV_X1 U10041 ( .A(n9109), .ZN(n7249) );
  NAND3_X1 U10042 ( .A1(n12886), .A2(n13318), .A3(n7062), .ZN(n7061) );
  NAND3_X1 U10043 ( .A1(n7066), .A2(n13348), .A3(n6536), .ZN(n7065) );
  XNOR2_X2 U10044 ( .A(n9018), .B(n9017), .ZN(n9019) );
  NAND2_X1 U10045 ( .A1(n7072), .A2(n7073), .ZN(n12965) );
  NAND2_X1 U10046 ( .A1(n12953), .A2(n6533), .ZN(n7072) );
  INV_X1 U10047 ( .A(n12960), .ZN(n7083) );
  NAND2_X1 U10048 ( .A1(n12951), .A2(n13006), .ZN(n7084) );
  OR2_X1 U10049 ( .A1(n12979), .A2(n12978), .ZN(n7093) );
  NAND2_X1 U10050 ( .A1(n9356), .A2(n9640), .ZN(n7094) );
  NAND2_X1 U10051 ( .A1(n7262), .A2(n7096), .ZN(n7095) );
  INV_X1 U10052 ( .A(n10830), .ZN(n7096) );
  NAND3_X1 U10053 ( .A1(n7103), .A2(n7105), .A3(n7982), .ZN(n7104) );
  NAND2_X1 U10054 ( .A1(n14301), .A2(n14031), .ZN(n7103) );
  NAND2_X1 U10055 ( .A1(n7104), .A2(n7980), .ZN(n14248) );
  NAND2_X2 U10056 ( .A1(n14248), .A2(n10560), .ZN(n14230) );
  NOR2_X1 U10057 ( .A1(n10444), .A2(n7111), .ZN(n7110) );
  NAND2_X1 U10058 ( .A1(n7311), .A2(n7973), .ZN(n14387) );
  NAND2_X1 U10059 ( .A1(n7313), .A2(n7112), .ZN(n7312) );
  NAND3_X1 U10060 ( .A1(n7280), .A2(n7311), .A3(n6538), .ZN(n7112) );
  AND2_X2 U10061 ( .A1(n10166), .A2(n10224), .ZN(n10232) );
  NAND2_X1 U10062 ( .A1(n7120), .A2(n9592), .ZN(n7621) );
  OAI21_X1 U10063 ( .B1(n11151), .B2(n11152), .A(n7120), .ZN(n11153) );
  OAI21_X1 U10064 ( .B1(n7121), .B2(P3_REG2_REG_1__SCAN_IN), .A(n11032), .ZN(
        n11035) );
  INV_X1 U10065 ( .A(n7125), .ZN(n13046) );
  INV_X1 U10066 ( .A(n7130), .ZN(n9614) );
  INV_X1 U10067 ( .A(n9600), .ZN(n7135) );
  NAND3_X1 U10068 ( .A1(n7132), .A2(n6716), .A3(n7131), .ZN(n7630) );
  NAND2_X1 U10069 ( .A1(n9602), .A2(n7138), .ZN(n7136) );
  INV_X1 U10070 ( .A(n7628), .ZN(n13140) );
  NAND2_X1 U10071 ( .A1(n14782), .A2(n14678), .ZN(n7140) );
  NAND3_X1 U10072 ( .A1(n10005), .A2(n10003), .A3(n10004), .ZN(n10007) );
  NAND2_X1 U10073 ( .A1(n8215), .A2(n8138), .ZN(n7142) );
  NAND2_X1 U10074 ( .A1(n8136), .A2(n7141), .ZN(n7143) );
  NAND3_X1 U10075 ( .A1(n7143), .A2(n8139), .A3(n7142), .ZN(n7214) );
  NAND2_X1 U10076 ( .A1(n7144), .A2(n8138), .ZN(n8319) );
  NAND2_X1 U10077 ( .A1(n8214), .A2(n7146), .ZN(n7144) );
  INV_X1 U10078 ( .A(n8139), .ZN(n8320) );
  NAND2_X1 U10079 ( .A1(n11001), .A2(n8775), .ZN(n7148) );
  NAND2_X1 U10080 ( .A1(n11537), .A2(n9107), .ZN(n11536) );
  NAND2_X1 U10081 ( .A1(n11477), .A2(n9072), .ZN(n11634) );
  OAI21_X2 U10082 ( .B1(n13357), .B2(n8077), .A(n6712), .ZN(n13346) );
  NAND2_X1 U10083 ( .A1(n12090), .A2(n7160), .ZN(n7157) );
  NAND2_X1 U10084 ( .A1(n7157), .A2(n7158), .ZN(n13398) );
  AND3_X1 U10085 ( .A1(n7917), .A2(n7918), .A3(n9547), .ZN(n9016) );
  NAND4_X1 U10086 ( .A1(n7917), .A2(n7918), .A3(n9547), .A4(n9017), .ZN(n13603) );
  NAND2_X1 U10087 ( .A1(n7168), .A2(n7169), .ZN(n7167) );
  NOR2_X1 U10088 ( .A1(n15484), .A2(n7731), .ZN(n7168) );
  NAND3_X1 U10089 ( .A1(n9746), .A2(n7342), .A3(n9747), .ZN(n15472) );
  OR2_X1 U10090 ( .A1(n9750), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7174) );
  NAND2_X1 U10091 ( .A1(n15473), .A2(n15474), .ZN(n15470) );
  NAND2_X1 U10092 ( .A1(n7175), .A2(n9750), .ZN(n15473) );
  NAND2_X1 U10093 ( .A1(n7176), .A2(n8642), .ZN(n8644) );
  NAND2_X1 U10094 ( .A1(n7464), .A2(n7462), .ZN(n7176) );
  NAND2_X1 U10095 ( .A1(n7179), .A2(n7178), .ZN(n7177) );
  NAND2_X1 U10096 ( .A1(n7451), .A2(n7450), .ZN(n7179) );
  NAND2_X1 U10097 ( .A1(n8616), .A2(n8615), .ZN(n7180) );
  NAND3_X1 U10098 ( .A1(n7728), .A2(n7182), .A3(n7729), .ZN(n7181) );
  NAND3_X1 U10099 ( .A1(n7728), .A2(n15493), .A3(n7729), .ZN(n15491) );
  NAND3_X1 U10100 ( .A1(n8325), .A2(n7291), .A3(n7289), .ZN(n7186) );
  NAND2_X1 U10101 ( .A1(n7184), .A2(n8345), .ZN(n8362) );
  NAND4_X1 U10102 ( .A1(n7186), .A2(n7187), .A3(n7185), .A4(n8827), .ZN(n7184)
         );
  NAND2_X1 U10103 ( .A1(n7188), .A2(n7289), .ZN(n7185) );
  NAND2_X1 U10104 ( .A1(n8325), .A2(n7189), .ZN(n7187) );
  OAI21_X1 U10105 ( .B1(n8693), .B2(n7194), .A(n7193), .ZN(n8699) );
  NAND2_X1 U10106 ( .A1(n7192), .A2(n7190), .ZN(n7257) );
  NAND2_X1 U10107 ( .A1(n8693), .A2(n7193), .ZN(n7192) );
  NAND2_X2 U10108 ( .A1(n7196), .A2(n7195), .ZN(n8261) );
  XNOR2_X1 U10109 ( .A(n15163), .B(n8969), .ZN(n8743) );
  INV_X1 U10110 ( .A(n9743), .ZN(n7198) );
  NAND2_X1 U10111 ( .A1(n15456), .A2(n7197), .ZN(n7199) );
  NAND2_X2 U10112 ( .A1(n7475), .A2(n8103), .ZN(n8474) );
  AND2_X2 U10113 ( .A1(n8283), .A2(n8101), .ZN(n8216) );
  OAI21_X1 U10114 ( .B1(n15755), .B2(n7204), .A(n14177), .ZN(n7503) );
  INV_X1 U10115 ( .A(n7205), .ZN(n10221) );
  XNOR2_X1 U10116 ( .A(n7205), .B(n14096), .ZN(n14044) );
  NAND2_X2 U10117 ( .A1(n10220), .A2(n10219), .ZN(n7205) );
  NAND2_X1 U10118 ( .A1(n7689), .A2(n12639), .ZN(n7686) );
  OAI211_X1 U10119 ( .C1(n13707), .C2(n7209), .A(n7689), .B(n7206), .ZN(n7685)
         );
  NAND2_X2 U10120 ( .A1(n7211), .A2(n7210), .ZN(n8347) );
  AOI21_X1 U10121 ( .B1(n8142), .B2(n7213), .A(n6676), .ZN(n7210) );
  NAND2_X1 U10122 ( .A1(n8319), .A2(n7212), .ZN(n7211) );
  AND2_X1 U10123 ( .A1(n8142), .A2(n8139), .ZN(n7212) );
  INV_X1 U10124 ( .A(n8141), .ZN(n7213) );
  NAND2_X1 U10125 ( .A1(n7216), .A2(n7364), .ZN(n7215) );
  INV_X1 U10126 ( .A(n7219), .ZN(n7216) );
  NAND2_X1 U10127 ( .A1(n13715), .A2(n12659), .ZN(n7219) );
  OAI21_X2 U10128 ( .B1(n12126), .B2(n7225), .A(n7222), .ZN(n13677) );
  NAND2_X1 U10129 ( .A1(n8868), .A2(n8867), .ZN(n7372) );
  NAND2_X1 U10130 ( .A1(n8842), .A2(n6565), .ZN(n7374) );
  NAND2_X1 U10131 ( .A1(n6675), .A2(n7373), .ZN(n8843) );
  NAND2_X1 U10132 ( .A1(n7227), .A2(n7268), .ZN(n7287) );
  NAND3_X1 U10133 ( .A1(n13965), .A2(n7229), .A3(n7228), .ZN(n7702) );
  NAND3_X1 U10134 ( .A1(n13934), .A2(n13932), .A3(n13933), .ZN(n7229) );
  INV_X1 U10135 ( .A(n13951), .ZN(n7265) );
  NAND2_X1 U10136 ( .A1(n10285), .A2(n8189), .ZN(n8639) );
  NAND2_X1 U10137 ( .A1(n9784), .A2(n11329), .ZN(n11330) );
  NAND2_X1 U10138 ( .A1(n11607), .A2(n11608), .ZN(n11766) );
  NAND2_X1 U10139 ( .A1(n12723), .A2(n12722), .ZN(n12780) );
  OAI21_X1 U10140 ( .B1(n13403), .B2(n9816), .A(n9815), .ZN(n12541) );
  NAND2_X1 U10141 ( .A1(n7232), .A2(n11093), .ZN(n11279) );
  NAND2_X1 U10142 ( .A1(n9783), .A2(n15860), .ZN(n7232) );
  NAND2_X1 U10143 ( .A1(n7937), .A2(n7938), .ZN(n9831) );
  NAND2_X2 U10144 ( .A1(n12830), .A2(n12831), .ZN(n12829) );
  AOI21_X1 U10145 ( .B1(n15858), .B2(n15857), .A(n9056), .ZN(n11478) );
  AOI21_X1 U10146 ( .B1(n13398), .B2(n9233), .A(n9232), .ZN(n13390) );
  INV_X1 U10147 ( .A(n12618), .ZN(n7234) );
  NAND2_X1 U10148 ( .A1(n9145), .A2(n12884), .ZN(n11847) );
  NAND2_X1 U10149 ( .A1(n9039), .A2(n9038), .ZN(n15858) );
  OAI211_X1 U10150 ( .C1(n7365), .C2(n7310), .A(n10802), .B(n10803), .ZN(
        n10816) );
  NAND3_X1 U10151 ( .A1(n7235), .A2(n12997), .A3(n13251), .ZN(n13003) );
  NAND2_X1 U10152 ( .A1(n7574), .A2(n15853), .ZN(n7573) );
  OAI211_X1 U10153 ( .C1(n13016), .C2(n13017), .A(n7237), .B(n7236), .ZN(
        n13021) );
  NAND2_X1 U10154 ( .A1(n7571), .A2(n7769), .ZN(n7236) );
  AOI21_X2 U10155 ( .B1(n13216), .B2(n9456), .A(n9455), .ZN(n13199) );
  NAND2_X1 U10156 ( .A1(n7256), .A2(n15443), .ZN(n7254) );
  NAND2_X1 U10157 ( .A1(n15444), .A2(n15445), .ZN(n15443) );
  NAND2_X1 U10158 ( .A1(n14503), .A2(n14502), .ZN(n14508) );
  NAND2_X1 U10159 ( .A1(n12163), .A2(n9983), .ZN(n14725) );
  INV_X1 U10160 ( .A(n11150), .ZN(n7532) );
  OAI21_X2 U10161 ( .B1(n12162), .B2(n10292), .A(n10289), .ZN(n14522) );
  AOI21_X1 U10162 ( .B1(n7741), .B2(n7007), .A(n7740), .ZN(n7739) );
  NAND3_X2 U10163 ( .A1(n7538), .A2(n7537), .A3(n8908), .ZN(n15063) );
  NAND2_X1 U10164 ( .A1(n7338), .A2(n7337), .ZN(n11161) );
  NAND2_X1 U10165 ( .A1(n7553), .A2(n7552), .ZN(n8038) );
  NAND3_X1 U10166 ( .A1(n7242), .A2(n7241), .A3(n7240), .ZN(P1_U3262) );
  NAND2_X1 U10167 ( .A1(n7588), .A2(n9258), .ZN(n9354) );
  NAND3_X1 U10168 ( .A1(n7129), .A2(n7128), .A3(n7282), .ZN(n9063) );
  AOI22_X2 U10169 ( .A1(n12541), .A2(n12540), .B1(n9818), .B2(n13392), .ZN(
        n12830) );
  NAND2_X1 U10170 ( .A1(n11456), .A2(n11419), .ZN(n11421) );
  NAND2_X2 U10171 ( .A1(n11727), .A2(n11726), .ZN(n12712) );
  NAND3_X1 U10172 ( .A1(n11131), .A2(n11124), .A3(n9588), .ZN(n7616) );
  NAND2_X1 U10173 ( .A1(n10713), .A2(n10714), .ZN(n7273) );
  INV_X1 U10174 ( .A(n7273), .ZN(n14192) );
  OR2_X1 U10175 ( .A1(n10675), .A2(n13193), .ZN(n7245) );
  OAI21_X2 U10176 ( .B1(n13364), .B2(n7898), .A(n7896), .ZN(n13295) );
  OAI21_X1 U10177 ( .B1(n13756), .B2(n13757), .A(n13761), .ZN(n7365) );
  NAND2_X1 U10178 ( .A1(n11935), .A2(n11934), .ZN(n10429) );
  INV_X1 U10179 ( .A(n12234), .ZN(n12126) );
  NAND2_X1 U10180 ( .A1(n7676), .A2(n7675), .ZN(n12234) );
  NOR2_X1 U10181 ( .A1(n13816), .A2(n11714), .ZN(n13762) );
  NAND2_X1 U10182 ( .A1(n8702), .A2(n8701), .ZN(n7259) );
  INV_X1 U10183 ( .A(SI_22_), .ZN(n7246) );
  NAND2_X1 U10184 ( .A1(n9359), .A2(n9324), .ZN(n9362) );
  NAND2_X1 U10185 ( .A1(n7251), .A2(n7250), .ZN(n12904) );
  NAND3_X2 U10186 ( .A1(n7402), .A2(n7920), .A3(n9548), .ZN(n7403) );
  INV_X1 U10187 ( .A(n10816), .ZN(n10813) );
  XNOR2_X1 U10188 ( .A(n11364), .B(n11420), .ZN(n13761) );
  NAND2_X1 U10189 ( .A1(n13668), .A2(n12649), .ZN(n12653) );
  XNOR2_X1 U10190 ( .A(n7254), .B(n6643), .ZN(SUB_1596_U4) );
  NOR2_X2 U10191 ( .A1(n14757), .A2(n10031), .ZN(n14804) );
  NAND2_X1 U10192 ( .A1(n7255), .A2(n12643), .ZN(n12644) );
  NAND3_X1 U10193 ( .A1(n13665), .A2(n13666), .A3(n13655), .ZN(n7255) );
  NAND2_X1 U10194 ( .A1(n11024), .A2(n11025), .ZN(n7736) );
  NAND2_X1 U10195 ( .A1(n14712), .A2(n14711), .ZN(n14710) );
  NAND2_X1 U10196 ( .A1(n7331), .A2(n15443), .ZN(n7260) );
  OAI21_X1 U10197 ( .B1(n8872), .B2(n8873), .A(n8871), .ZN(P1_U3242) );
  NAND2_X1 U10198 ( .A1(n7257), .A2(n8696), .ZN(n8698) );
  OAI21_X1 U10199 ( .B1(n8674), .B2(n7467), .A(n7288), .ZN(n8693) );
  NAND2_X1 U10200 ( .A1(n7333), .A2(n7332), .ZN(n7331) );
  XNOR2_X1 U10201 ( .A(n7260), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  INV_X1 U10202 ( .A(n8946), .ZN(n8951) );
  OAI21_X1 U10203 ( .B1(n15040), .B2(n8058), .A(n8057), .ZN(n10660) );
  AND2_X2 U10204 ( .A1(n10722), .A2(n7647), .ZN(n14186) );
  NAND2_X1 U10205 ( .A1(n11536), .A2(n7608), .ZN(n11688) );
  NAND2_X1 U10206 ( .A1(n11478), .A2(n12879), .ZN(n11477) );
  NOR2_X1 U10207 ( .A1(n9102), .A2(P3_IR_REG_28__SCAN_IN), .ZN(n7917) );
  NAND2_X2 U10208 ( .A1(n9021), .A2(n9020), .ZN(n9058) );
  NAND2_X1 U10209 ( .A1(n9051), .A2(n9050), .ZN(n9066) );
  NAND2_X1 U10210 ( .A1(n9100), .A2(n9099), .ZN(n9117) );
  NAND2_X1 U10211 ( .A1(n9369), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9372) );
  NAND2_X1 U10212 ( .A1(n7264), .A2(n13986), .ZN(n14017) );
  OAI22_X1 U10213 ( .A1(n14014), .A2(n14015), .B1(n14009), .B2(n14010), .ZN(
        n7264) );
  NAND2_X1 U10214 ( .A1(n14811), .A2(n14812), .ZN(n14810) );
  NOR2_X2 U10215 ( .A1(n7266), .A2(n6575), .ZN(n13715) );
  OAI21_X1 U10216 ( .B1(n8610), .B2(n8609), .A(n8608), .ZN(n8612) );
  INV_X1 U10217 ( .A(n11913), .ZN(n7305) );
  NAND2_X1 U10218 ( .A1(n12645), .A2(n7688), .ZN(n7684) );
  NAND3_X1 U10219 ( .A1(n7680), .A2(n12652), .A3(n7267), .ZN(n13645) );
  AOI21_X1 U10220 ( .B1(n12654), .B2(n13649), .A(n13645), .ZN(n12656) );
  NAND2_X1 U10221 ( .A1(n10585), .A2(n14076), .ZN(n10798) );
  INV_X1 U10222 ( .A(n14021), .ZN(n7268) );
  NAND2_X1 U10223 ( .A1(n12558), .A2(n10251), .ZN(n10170) );
  NAND2_X1 U10224 ( .A1(n7269), .A2(n6722), .ZN(n14083) );
  INV_X1 U10225 ( .A(n14079), .ZN(n7269) );
  NAND2_X1 U10226 ( .A1(n14468), .A2(n10464), .ZN(n14440) );
  NAND2_X1 U10227 ( .A1(n10412), .A2(n10411), .ZN(n15766) );
  NOR2_X2 U10228 ( .A1(n11176), .A2(n11177), .ZN(n11175) );
  NAND2_X1 U10229 ( .A1(n7530), .A2(n7522), .ZN(n7521) );
  NAND2_X1 U10230 ( .A1(n11544), .A2(n11543), .ZN(n7510) );
  NAND2_X1 U10231 ( .A1(n15477), .A2(n15476), .ZN(n15475) );
  AND2_X2 U10232 ( .A1(n9877), .A2(n8914), .ZN(n10111) );
  XNOR2_X1 U10233 ( .A(n7838), .B(n8252), .ZN(n10907) );
  NAND2_X1 U10234 ( .A1(n14810), .A2(n10107), .ZN(n10149) );
  NAND2_X1 U10235 ( .A1(n11973), .A2(n10390), .ZN(n11368) );
  NAND3_X1 U10236 ( .A1(n10587), .A2(n10388), .A3(n10387), .ZN(n11973) );
  NAND2_X1 U10237 ( .A1(n12696), .A2(n10301), .ZN(n7275) );
  NAND2_X1 U10238 ( .A1(n6517), .A2(n6666), .ZN(n8818) );
  NAND2_X1 U10239 ( .A1(n14725), .A2(n10009), .ZN(n7756) );
  AOI21_X1 U10240 ( .B1(n7974), .B2(n10481), .A(n6547), .ZN(n7973) );
  NAND2_X1 U10241 ( .A1(n14182), .A2(n14495), .ZN(n14503) );
  NAND2_X1 U10242 ( .A1(n10386), .A2(n10589), .ZN(n10587) );
  NAND2_X1 U10243 ( .A1(n7685), .A2(n7683), .ZN(n13668) );
  NAND2_X1 U10244 ( .A1(n13676), .A2(n12606), .ZN(n13740) );
  NAND2_X1 U10245 ( .A1(n13021), .A2(n13020), .ZN(n7576) );
  NAND2_X1 U10246 ( .A1(n7576), .A2(n7575), .ZN(n7574) );
  XNOR2_X1 U10247 ( .A(n11420), .B(n13843), .ZN(n11417) );
  INV_X1 U10248 ( .A(n7691), .ZN(n7690) );
  NAND2_X1 U10249 ( .A1(n13677), .A2(n13678), .ZN(n13676) );
  INV_X4 U10250 ( .A(n11420), .ZN(n11713) );
  OR2_X1 U10251 ( .A1(n11460), .A2(n10804), .ZN(n10805) );
  NAND2_X2 U10252 ( .A1(n10798), .A2(n14068), .ZN(n11420) );
  NAND3_X1 U10253 ( .A1(n13756), .A2(n11270), .A3(n7283), .ZN(n10802) );
  INV_X1 U10254 ( .A(n11271), .ZN(n7283) );
  OAI21_X1 U10255 ( .B1(n10360), .B2(n7285), .A(n6687), .ZN(P2_U3530) );
  OAI21_X1 U10256 ( .B1(n10360), .B2(n7304), .A(n6686), .ZN(P2_U3498) );
  NAND3_X1 U10257 ( .A1(n8308), .A2(n6515), .A3(n11487), .ZN(n7291) );
  NAND2_X1 U10258 ( .A1(n7448), .A2(n8263), .ZN(n7447) );
  NAND3_X1 U10259 ( .A1(n7920), .A2(n9547), .A3(n7292), .ZN(n9551) );
  NAND2_X1 U10260 ( .A1(n10618), .A2(n10617), .ZN(n14305) );
  OAI211_X2 U10261 ( .C1(n10907), .C2(n10292), .A(n7634), .B(n7297), .ZN(
        n10379) );
  OR2_X1 U10262 ( .A1(n6519), .A2(n10847), .ZN(n7297) );
  NAND2_X4 U10263 ( .A1(n8568), .A2(n8567), .ZN(n15330) );
  NAND2_X1 U10264 ( .A1(n7298), .A2(n14813), .ZN(n10158) );
  NAND2_X1 U10265 ( .A1(n7351), .A2(n10148), .ZN(n7298) );
  NAND2_X1 U10266 ( .A1(n8056), .A2(n8052), .ZN(n14986) );
  OAI211_X1 U10267 ( .C1(n15280), .C2(n15360), .A(n15282), .B(n15279), .ZN(
        n15402) );
  NAND3_X1 U10268 ( .A1(n7756), .A2(n7754), .A3(n7329), .ZN(n7339) );
  OAI21_X1 U10269 ( .B1(n6602), .B2(n14224), .A(n14226), .ZN(n14512) );
  AOI21_X1 U10270 ( .B1(n14243), .B2(n10627), .A(n10624), .ZN(n14236) );
  AOI211_X1 U10271 ( .C1(n14514), .C2(n15835), .A(n14513), .B(n14512), .ZN(
        n14618) );
  NAND2_X1 U10272 ( .A1(n7997), .A2(n7996), .ZN(n14182) );
  NAND2_X1 U10273 ( .A1(n7312), .A2(n10507), .ZN(n14335) );
  INV_X1 U10274 ( .A(n9588), .ZN(n7611) );
  NAND2_X1 U10275 ( .A1(n7903), .A2(n7901), .ZN(n10596) );
  NAND2_X1 U10276 ( .A1(n7862), .A2(n10600), .ZN(n14403) );
  NAND2_X1 U10277 ( .A1(n10599), .A2(n10598), .ZN(n12028) );
  NAND2_X1 U10278 ( .A1(n10714), .A2(n7341), .ZN(n10650) );
  AND2_X1 U10279 ( .A1(n11459), .A2(n11416), .ZN(n7309) );
  INV_X1 U10280 ( .A(n10800), .ZN(n13756) );
  NAND2_X1 U10281 ( .A1(n13775), .A2(n12639), .ZN(n7688) );
  NAND2_X1 U10282 ( .A1(n7684), .A2(n7689), .ZN(n7683) );
  NAND2_X1 U10283 ( .A1(n13623), .A2(n6672), .ZN(n12681) );
  NAND2_X1 U10284 ( .A1(n12560), .A2(n12698), .ZN(n10381) );
  NAND2_X1 U10285 ( .A1(n14428), .A2(n7974), .ZN(n7311) );
  NAND3_X1 U10286 ( .A1(n14083), .A2(n14084), .A3(n7314), .ZN(P2_U3328) );
  AOI21_X1 U10287 ( .B1(n14236), .B2(n14235), .A(n10625), .ZN(n14223) );
  NOR2_X2 U10288 ( .A1(n10182), .A2(n10165), .ZN(n10166) );
  OAI21_X1 U10289 ( .B1(n14618), .B2(n7285), .A(n7318), .ZN(P2_U3525) );
  NAND2_X1 U10290 ( .A1(n7737), .A2(n7736), .ZN(n15505) );
  INV_X1 U10291 ( .A(n11515), .ZN(n7749) );
  NAND2_X1 U10292 ( .A1(n7323), .A2(n7322), .ZN(P2_U3186) );
  NAND2_X1 U10293 ( .A1(n13627), .A2(n13626), .ZN(n7323) );
  AOI21_X2 U10294 ( .B1(n15063), .B2(n8910), .A(n8909), .ZN(n15043) );
  OAI22_X2 U10295 ( .A1(n15043), .A2(n15044), .B1(n15053), .B2(n15031), .ZN(
        n15027) );
  NAND2_X1 U10296 ( .A1(n7349), .A2(n6690), .ZN(n7553) );
  INV_X1 U10297 ( .A(n8038), .ZN(n15000) );
  XNOR2_X2 U10298 ( .A(n15330), .B(n15116), .ZN(n15134) );
  NAND3_X2 U10299 ( .A1(n8032), .A2(n8906), .A3(n8033), .ZN(n15123) );
  NOR2_X1 U10300 ( .A1(n15929), .A2(n15930), .ZN(n15928) );
  AOI21_X1 U10301 ( .B1(n7677), .B2(n6531), .A(n6667), .ZN(n7675) );
  NOR2_X1 U10302 ( .A1(n14034), .A2(n7975), .ZN(n7974) );
  NAND2_X1 U10303 ( .A1(n8347), .A2(n8145), .ZN(n8375) );
  NAND2_X1 U10304 ( .A1(n10723), .A2(n15848), .ZN(n7926) );
  NAND2_X1 U10305 ( .A1(n7835), .A2(n6698), .ZN(n8676) );
  NOR2_X1 U10306 ( .A1(n7928), .A2(n7995), .ZN(n7927) );
  NAND2_X1 U10307 ( .A1(n8645), .A2(n7666), .ZN(n7665) );
  OAI21_X1 U10308 ( .B1(n7258), .B2(n8699), .A(n8698), .ZN(n8789) );
  OAI211_X1 U10309 ( .C1(n8492), .C2(n7638), .A(n7636), .B(n8579), .ZN(n7640)
         );
  NAND2_X1 U10310 ( .A1(n7640), .A2(n7449), .ZN(n7451) );
  XNOR2_X1 U10311 ( .A(n9729), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n9730) );
  NAND2_X1 U10312 ( .A1(n7994), .A2(n7991), .ZN(P2_U3495) );
  NAND2_X1 U10313 ( .A1(n9188), .A2(n7776), .ZN(n7774) );
  NAND2_X1 U10314 ( .A1(n7926), .A2(n7385), .ZN(P2_U3527) );
  AND2_X1 U10315 ( .A1(n10606), .A2(n8074), .ZN(n10607) );
  NAND2_X1 U10316 ( .A1(n10147), .A2(n7343), .ZN(P1_U3220) );
  NAND2_X1 U10317 ( .A1(n10127), .A2(n7344), .ZN(n7343) );
  NAND2_X1 U10318 ( .A1(n14028), .A2(n6683), .ZN(n14016) );
  NAND2_X1 U10319 ( .A1(n7347), .A2(n7346), .ZN(n7345) );
  INV_X1 U10320 ( .A(n14013), .ZN(n7347) );
  NAND2_X1 U10321 ( .A1(n8723), .A2(n8722), .ZN(n14656) );
  INV_X1 U10322 ( .A(n15027), .ZN(n7349) );
  OAI21_X1 U10323 ( .B1(n7543), .B2(n7542), .A(n15076), .ZN(n7541) );
  INV_X1 U10324 ( .A(n14374), .ZN(n7885) );
  NAND2_X1 U10325 ( .A1(n7353), .A2(n7352), .ZN(n7351) );
  INV_X1 U10326 ( .A(n10149), .ZN(n7353) );
  OR2_X1 U10327 ( .A1(n13955), .A2(n13925), .ZN(n13929) );
  NAND2_X1 U10328 ( .A1(n7701), .A2(n7700), .ZN(n7699) );
  NAND2_X1 U10329 ( .A1(n7356), .A2(n7355), .ZN(n11182) );
  INV_X1 U10330 ( .A(n9597), .ZN(n7357) );
  NAND2_X1 U10331 ( .A1(n7630), .A2(n11066), .ZN(n9602) );
  NAND3_X1 U10332 ( .A1(n8837), .A2(n15108), .A3(n7375), .ZN(n8838) );
  AND2_X1 U10333 ( .A1(n11717), .A2(n11711), .ZN(n7679) );
  NAND2_X1 U10334 ( .A1(n7882), .A2(n7883), .ZN(n14358) );
  NAND2_X1 U10335 ( .A1(n7380), .A2(n7377), .ZN(P2_U3526) );
  NAND2_X1 U10336 ( .A1(n14510), .A2(n15848), .ZN(n7380) );
  NOR2_X1 U10337 ( .A1(n10611), .A2(n7888), .ZN(n7887) );
  NAND2_X1 U10338 ( .A1(n11665), .A2(n11660), .ZN(n9039) );
  NAND2_X1 U10339 ( .A1(n11662), .A2(n13044), .ZN(n11665) );
  NAND2_X1 U10340 ( .A1(n11737), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n11891) );
  NAND2_X1 U10341 ( .A1(n11182), .A2(n7619), .ZN(n7618) );
  NAND2_X1 U10342 ( .A1(n8131), .A2(n8130), .ZN(n8234) );
  NAND2_X1 U10343 ( .A1(n8124), .A2(n8123), .ZN(n8279) );
  NAND2_X1 U10344 ( .A1(n14206), .A2(n7927), .ZN(n10723) );
  NOR2_X1 U10345 ( .A1(n14201), .A2(n15817), .ZN(n7928) );
  NAND3_X1 U10346 ( .A1(n9383), .A2(n13286), .A3(n13283), .ZN(n7603) );
  NAND2_X1 U10347 ( .A1(n9035), .A2(P3_IR_REG_1__SCAN_IN), .ZN(n7507) );
  NAND2_X1 U10348 ( .A1(n9759), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n7728) );
  INV_X1 U10349 ( .A(n9063), .ZN(n7393) );
  NAND2_X4 U10350 ( .A1(n7395), .A2(n7403), .ZN(n13612) );
  NOR2_X1 U10351 ( .A1(n7401), .A2(n7400), .ZN(n7397) );
  NAND2_X1 U10352 ( .A1(n9551), .A2(n6692), .ZN(n7398) );
  INV_X1 U10353 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n7400) );
  NAND2_X1 U10354 ( .A1(n13105), .A2(n7411), .ZN(n7410) );
  NAND2_X1 U10355 ( .A1(n11745), .A2(n6684), .ZN(n7420) );
  OAI21_X1 U10356 ( .B1(n11147), .B2(n7434), .A(n7431), .ZN(n7445) );
  INV_X1 U10357 ( .A(n11147), .ZN(n7444) );
  NAND2_X1 U10358 ( .A1(n7436), .A2(n7437), .ZN(n11173) );
  INV_X1 U10359 ( .A(n7432), .ZN(n11298) );
  MUX2_X1 U10360 ( .A(n8250), .B(n8251), .S(n8261), .Z(n7448) );
  NAND2_X1 U10361 ( .A1(n7451), .A2(n6679), .ZN(n8616) );
  NAND2_X1 U10362 ( .A1(n8404), .A2(n7458), .ZN(n7455) );
  NAND2_X1 U10363 ( .A1(n7455), .A2(n7456), .ZN(n8424) );
  INV_X1 U10364 ( .A(n8629), .ZN(n7465) );
  NAND2_X1 U10365 ( .A1(n7470), .A2(n7469), .ZN(n15546) );
  OR2_X1 U10366 ( .A1(n11510), .A2(n11509), .ZN(n7469) );
  NAND2_X1 U10367 ( .A1(n11510), .A2(n11509), .ZN(n7470) );
  INV_X1 U10368 ( .A(n8937), .ZN(n15170) );
  AND2_X1 U10369 ( .A1(n8763), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n8071) );
  AND2_X2 U10370 ( .A1(n8111), .A2(n8110), .ZN(n8763) );
  XNOR2_X1 U10371 ( .A(n15022), .B(n15021), .ZN(n7491) );
  AOI21_X1 U10372 ( .B1(n7491), .B2(n7490), .A(n7488), .ZN(n15025) );
  AOI21_X1 U10373 ( .B1(n15288), .B2(n15254), .A(n15024), .ZN(n7492) );
  OAI21_X2 U10374 ( .B1(n9046), .B2(P3_IR_REG_1__SCAN_IN), .A(n7507), .ZN(
        n10848) );
  INV_X1 U10375 ( .A(n7512), .ZN(n7511) );
  AOI21_X1 U10376 ( .B1(n13054), .B2(n7515), .A(n7516), .ZN(n7514) );
  INV_X1 U10377 ( .A(n9627), .ZN(n7517) );
  INV_X1 U10378 ( .A(n10998), .ZN(n7518) );
  NAND2_X1 U10379 ( .A1(n7530), .A2(n7528), .ZN(n7519) );
  NOR2_X1 U10380 ( .A1(n7524), .A2(n7523), .ZN(n7522) );
  INV_X1 U10381 ( .A(n7528), .ZN(n7524) );
  OR2_X2 U10382 ( .A1(n9621), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7527) );
  NAND2_X1 U10383 ( .A1(n9621), .A2(n7529), .ZN(n7528) );
  NAND2_X1 U10384 ( .A1(n15123), .A2(n7540), .ZN(n7538) );
  OR2_X1 U10385 ( .A1(n15027), .A2(n15039), .ZN(n7557) );
  INV_X1 U10386 ( .A(n7557), .ZN(n15026) );
  NAND3_X1 U10387 ( .A1(n12000), .A2(n12189), .A3(n8891), .ZN(n7559) );
  INV_X1 U10388 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7564) );
  NAND2_X1 U10389 ( .A1(n7572), .A2(n13012), .ZN(n7571) );
  NAND2_X1 U10390 ( .A1(n13009), .A2(n6682), .ZN(n7572) );
  NAND2_X1 U10391 ( .A1(n13003), .A2(n7772), .ZN(n13009) );
  NAND2_X1 U10392 ( .A1(n7577), .A2(n7578), .ZN(n12953) );
  NAND2_X1 U10393 ( .A1(n12931), .A2(n7580), .ZN(n7577) );
  INV_X1 U10394 ( .A(n11131), .ZN(n7612) );
  NAND3_X1 U10395 ( .A1(n7613), .A2(P3_REG2_REG_3__SCAN_IN), .A3(n7616), .ZN(
        n11115) );
  AOI21_X1 U10396 ( .B1(n11131), .B2(n9588), .A(n11124), .ZN(n7615) );
  NAND3_X1 U10397 ( .A1(n9602), .A2(n7628), .A3(n7627), .ZN(n9612) );
  XNOR2_X2 U10398 ( .A(n9046), .B(P3_IR_REG_2__SCAN_IN), .ZN(n11145) );
  NAND2_X1 U10399 ( .A1(n7633), .A2(n9877), .ZN(n8249) );
  NAND2_X1 U10400 ( .A1(n7633), .A2(n8828), .ZN(n11453) );
  AOI21_X1 U10401 ( .B1(n6537), .B2(n7633), .A(n7632), .ZN(n11510) );
  INV_X2 U10402 ( .A(n10379), .ZN(n11364) );
  NAND2_X1 U10403 ( .A1(n8546), .A2(n7639), .ZN(n7638) );
  NAND2_X1 U10404 ( .A1(n7644), .A2(n7641), .ZN(n10313) );
  AOI21_X1 U10405 ( .B1(n10722), .B2(n7643), .A(n7642), .ZN(n7641) );
  NAND2_X1 U10406 ( .A1(n10722), .A2(n14205), .ZN(n14187) );
  NAND3_X1 U10407 ( .A1(n8427), .A2(n6688), .A3(n8426), .ZN(n7649) );
  NAND2_X1 U10408 ( .A1(n7649), .A2(n7650), .ZN(n8490) );
  OAI22_X1 U10409 ( .A1(n7665), .A2(n6645), .B1(n8659), .B2(n7667), .ZN(n8674)
         );
  INV_X1 U10410 ( .A(n8658), .ZN(n7667) );
  NAND2_X1 U10411 ( .A1(n13634), .A2(n7673), .ZN(n7672) );
  NAND2_X1 U10412 ( .A1(n12712), .A2(n7677), .ZN(n7676) );
  OAI21_X1 U10413 ( .B1(n12712), .B2(n6531), .A(n7677), .ZN(n12597) );
  NAND2_X1 U10414 ( .A1(n11758), .A2(n11725), .ZN(n11727) );
  NAND2_X1 U10415 ( .A1(n13776), .A2(n7681), .ZN(n7680) );
  NOR2_X1 U10416 ( .A1(n13845), .A2(n13848), .ZN(n7697) );
  OAI21_X1 U10417 ( .B1(n6617), .B2(n7707), .A(n7706), .ZN(n13905) );
  NAND3_X1 U10418 ( .A1(n7713), .A2(n7714), .A3(n7712), .ZN(n7710) );
  INV_X1 U10419 ( .A(n13903), .ZN(n7715) );
  INV_X1 U10420 ( .A(n13901), .ZN(n7716) );
  NAND2_X1 U10421 ( .A1(n7719), .A2(n7720), .ZN(n13888) );
  NAND3_X1 U10422 ( .A1(n13883), .A2(n6665), .A3(n13882), .ZN(n7719) );
  NAND2_X1 U10423 ( .A1(n13890), .A2(n7722), .ZN(n7721) );
  NAND2_X1 U10424 ( .A1(n10173), .A2(n7727), .ZN(n10310) );
  NOR2_X1 U10425 ( .A1(n15481), .A2(n15480), .ZN(n15479) );
  NAND2_X1 U10426 ( .A1(n15480), .A2(n7734), .ZN(n7732) );
  INV_X1 U10427 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7734) );
  NAND2_X2 U10428 ( .A1(n10184), .A2(n10879), .ZN(n10185) );
  OAI21_X1 U10429 ( .B1(n7749), .B2(n7745), .A(n7744), .ZN(n11864) );
  INV_X1 U10430 ( .A(n7761), .ZN(n14802) );
  INV_X1 U10431 ( .A(n9048), .ZN(n7766) );
  NAND2_X1 U10432 ( .A1(n7766), .A2(n9049), .ZN(n9051) );
  NAND2_X1 U10433 ( .A1(n9458), .A2(n7801), .ZN(n7800) );
  OAI21_X1 U10434 ( .B1(n9458), .B2(n9457), .A(n9459), .ZN(n9475) );
  NAND2_X1 U10435 ( .A1(n8121), .A2(n7816), .ZN(n8124) );
  XNOR2_X1 U10436 ( .A(n7816), .B(n10850), .ZN(n8252) );
  AOI21_X2 U10437 ( .B1(n8189), .B2(n10282), .A(n8638), .ZN(n7817) );
  NAND2_X1 U10438 ( .A1(n8529), .A2(n6589), .ZN(n7822) );
  NAND2_X1 U10439 ( .A1(n8649), .A2(n8194), .ZN(n8669) );
  INV_X1 U10440 ( .A(n8675), .ZN(n7834) );
  NAND4_X1 U10441 ( .A1(n14498), .A2(n14061), .A3(n7836), .A4(n14028), .ZN(
        n14062) );
  NOR2_X2 U10442 ( .A1(n11391), .A2(n15554), .ZN(n11497) );
  AND2_X1 U10443 ( .A1(n8966), .A2(n15535), .ZN(n11505) );
  NAND2_X1 U10444 ( .A1(n15029), .A2(n6685), .ZN(n7841) );
  INV_X1 U10445 ( .A(n7841), .ZN(n10665) );
  NOR2_X4 U10446 ( .A1(n15002), .A2(n15003), .ZN(n15001) );
  INV_X1 U10447 ( .A(n7844), .ZN(n7842) );
  NAND2_X1 U10448 ( .A1(n15193), .A2(n7850), .ZN(n7852) );
  INV_X1 U10449 ( .A(n7852), .ZN(n15180) );
  NAND3_X1 U10450 ( .A1(n7855), .A2(n11571), .A3(n7856), .ZN(n11834) );
  INV_X1 U10451 ( .A(n7857), .ZN(n11586) );
  NAND3_X1 U10452 ( .A1(n7859), .A2(n7858), .A3(n15113), .ZN(n15055) );
  NAND2_X1 U10453 ( .A1(n14403), .A2(n10604), .ZN(n10608) );
  NAND2_X1 U10454 ( .A1(n12028), .A2(n14047), .ZN(n7862) );
  NAND2_X1 U10455 ( .A1(n12089), .A2(n7866), .ZN(n7864) );
  NAND2_X1 U10456 ( .A1(n10610), .A2(n6658), .ZN(n7882) );
  OAI21_X1 U10457 ( .B1(n13364), .B2(n6535), .A(n9517), .ZN(n13355) );
  AOI21_X1 U10458 ( .B1(n7904), .B2(n6562), .A(n7902), .ZN(n7901) );
  INV_X1 U10459 ( .A(n9014), .ZN(n7920) );
  NOR2_X2 U10460 ( .A1(n9014), .A2(n9102), .ZN(n9258) );
  INV_X1 U10461 ( .A(n12829), .ZN(n7933) );
  INV_X1 U10462 ( .A(n12733), .ZN(n7945) );
  AOI21_X1 U10463 ( .B1(n7941), .B2(n9826), .A(n7939), .ZN(n7938) );
  OAI211_X1 U10464 ( .C1(n12817), .C2(n7956), .A(n12832), .B(n7953), .ZN(n9876) );
  NAND2_X1 U10465 ( .A1(n12817), .A2(n7954), .ZN(n7953) );
  INV_X1 U10466 ( .A(n7958), .ZN(n7955) );
  NAND2_X1 U10467 ( .A1(n12817), .A2(n9849), .ZN(n7957) );
  NAND2_X1 U10468 ( .A1(n9850), .A2(n9848), .ZN(n7958) );
  INV_X1 U10469 ( .A(n9850), .ZN(n7959) );
  OAI21_X1 U10470 ( .B1(n12796), .B2(n7964), .A(n9844), .ZN(n12752) );
  NAND2_X1 U10471 ( .A1(n9833), .A2(n7965), .ZN(n7964) );
  NAND2_X1 U10472 ( .A1(n11330), .A2(n7968), .ZN(n11523) );
  NAND2_X1 U10473 ( .A1(n7969), .A2(n9260), .ZN(n9543) );
  INV_X1 U10474 ( .A(n14281), .ZN(n7989) );
  NAND2_X1 U10475 ( .A1(n14230), .A2(n8001), .ZN(n7997) );
  NAND2_X1 U10476 ( .A1(n14230), .A2(n8002), .ZN(n7998) );
  INV_X1 U10477 ( .A(n8011), .ZN(n8013) );
  NAND2_X1 U10478 ( .A1(n11580), .A2(n8021), .ZN(n8023) );
  AOI21_X1 U10479 ( .B1(n8026), .B2(n11673), .A(n6664), .ZN(n8024) );
  NAND2_X1 U10480 ( .A1(n8880), .A2(n8879), .ZN(n11385) );
  NAND3_X1 U10481 ( .A1(n8028), .A2(n8883), .A3(n8027), .ZN(n8885) );
  NAND2_X1 U10482 ( .A1(n8882), .A2(n6515), .ZN(n8027) );
  NAND3_X1 U10483 ( .A1(n8880), .A2(n8882), .A3(n8879), .ZN(n8028) );
  NAND2_X1 U10484 ( .A1(n8029), .A2(n8882), .ZN(n11486) );
  NAND2_X1 U10485 ( .A1(n11385), .A2(n8881), .ZN(n8029) );
  NAND2_X1 U10486 ( .A1(n15149), .A2(n8034), .ZN(n8032) );
  NAND2_X1 U10487 ( .A1(n9893), .A2(n9892), .ZN(n9895) );
  NAND2_X1 U10488 ( .A1(n8039), .A2(n10653), .ZN(n8037) );
  NAND4_X1 U10489 ( .A1(n6516), .A2(n8290), .A3(n8292), .A4(n8041), .ZN(n8918)
         );
  NAND2_X1 U10490 ( .A1(n14855), .A2(n8299), .ZN(n8829) );
  NAND2_X1 U10491 ( .A1(n10108), .A2(n14855), .ZN(n9901) );
  NAND2_X1 U10492 ( .A1(n12192), .A2(n8044), .ZN(n8043) );
  NAND2_X1 U10493 ( .A1(n8050), .A2(n8955), .ZN(n8059) );
  NAND2_X1 U10494 ( .A1(n15040), .A2(n15039), .ZN(n15038) );
  NAND2_X1 U10495 ( .A1(n15040), .A2(n8051), .ZN(n8056) );
  NAND2_X1 U10496 ( .A1(n15038), .A2(n8955), .ZN(n15022) );
  NAND2_X1 U10497 ( .A1(n8062), .A2(n8061), .ZN(n11584) );
  OR2_X1 U10498 ( .A1(n14996), .A2(n10659), .ZN(n8841) );
  NAND2_X1 U10499 ( .A1(n8845), .A2(n8844), .ZN(n8868) );
  NOR2_X1 U10500 ( .A1(n8866), .A2(n8865), .ZN(n8867) );
  NAND2_X1 U10501 ( .A1(n8297), .A2(n8296), .ZN(n8306) );
  NAND2_X1 U10502 ( .A1(n8297), .A2(n8066), .ZN(n8307) );
  OR2_X1 U10503 ( .A1(n14403), .A2(n10463), .ZN(n14469) );
  NAND2_X1 U10504 ( .A1(n8806), .A2(n8805), .ZN(n8872) );
  OAI21_X1 U10505 ( .B1(n10707), .B2(n10706), .A(n10705), .ZN(n10708) );
  NAND2_X1 U10506 ( .A1(n10707), .A2(n15905), .ZN(n9584) );
  OAI21_X1 U10507 ( .B1(n12850), .B2(n12849), .A(n12848), .ZN(n12852) );
  INV_X1 U10508 ( .A(n13196), .ZN(n12702) );
  AOI21_X1 U10509 ( .B1(n14188), .B2(n10720), .A(n10719), .ZN(n14059) );
  XNOR2_X1 U10510 ( .A(n8758), .B(n8757), .ZN(n12696) );
  NAND2_X1 U10511 ( .A1(n10309), .A2(n10337), .ZN(n10316) );
  NAND2_X1 U10512 ( .A1(n10305), .A2(n10306), .ZN(n10337) );
  INV_X1 U10513 ( .A(n9730), .ZN(n9732) );
  CLKBUF_X1 U10514 ( .A(n14413), .Z(n14430) );
  INV_X1 U10515 ( .A(n14393), .ZN(n14573) );
  NAND2_X1 U10516 ( .A1(n9441), .A2(n9440), .ZN(n9443) );
  NAND2_X1 U10517 ( .A1(n15852), .A2(n9055), .ZN(n12909) );
  INV_X1 U10518 ( .A(n8735), .ZN(n8721) );
  OR2_X1 U10519 ( .A1(n10597), .A2(n12070), .ZN(n12069) );
  INV_X1 U10520 ( .A(n14184), .ZN(n14205) );
  OAI21_X1 U10521 ( .B1(n14020), .B2(n14019), .A(n14018), .ZN(n14021) );
  NAND2_X1 U10522 ( .A1(n8978), .A2(n8977), .ZN(n9003) );
  XNOR2_X1 U10523 ( .A(n8128), .B(SI_3_), .ZN(n8275) );
  OR2_X1 U10524 ( .A1(n8125), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8122) );
  AOI21_X1 U10525 ( .B1(P1_REG0_REG_1__SCAN_IN), .B2(n8088), .A(n8071), .ZN(
        n8260) );
  INV_X1 U10526 ( .A(n8917), .ZN(n11509) );
  INV_X1 U10527 ( .A(n8110), .ZN(n15427) );
  AND2_X1 U10528 ( .A1(n8303), .A2(n11070), .ZN(n8065) );
  NAND2_X1 U10529 ( .A1(n8295), .A2(n8294), .ZN(n8066) );
  NAND2_X1 U10530 ( .A1(n15342), .A2(n15196), .ZN(n8067) );
  AND2_X1 U10531 ( .A1(n8544), .A2(n15173), .ZN(n8068) );
  INV_X1 U10532 ( .A(n13207), .ZN(n10700) );
  INV_X1 U10533 ( .A(n13992), .ZN(n14511) );
  NAND2_X2 U10534 ( .A1(n11790), .A2(n15776), .ZN(n15781) );
  OR2_X1 U10535 ( .A1(n12561), .A2(n14652), .ZN(n8069) );
  OR2_X1 U10536 ( .A1(n12561), .A2(n14602), .ZN(n8070) );
  INV_X1 U10537 ( .A(n15122), .ZN(n8906) );
  INV_X1 U10538 ( .A(n14470), .ZN(n10463) );
  AND2_X1 U10539 ( .A1(n14517), .A2(n14089), .ZN(n8072) );
  AND2_X1 U10540 ( .A1(n13646), .A2(n12655), .ZN(n8075) );
  OR2_X1 U10541 ( .A1(n8126), .A2(n10854), .ZN(n8076) );
  AND2_X1 U10542 ( .A1(n12769), .A2(n12774), .ZN(n8077) );
  OR2_X1 U10543 ( .A1(n12778), .A2(n12810), .ZN(n8078) );
  AND2_X1 U10544 ( .A1(n9336), .A2(n9335), .ZN(n8079) );
  AND3_X1 U10545 ( .A1(n10129), .A2(n10128), .A3(n14813), .ZN(n8081) );
  OR2_X1 U10546 ( .A1(n12702), .A2(n13496), .ZN(n8082) );
  AND2_X1 U10547 ( .A1(n9941), .A2(n9940), .ZN(n8083) );
  AND2_X1 U10548 ( .A1(n14683), .A2(n10003), .ZN(n8084) );
  INV_X1 U10549 ( .A(n14262), .ZN(n10559) );
  AND2_X1 U10550 ( .A1(n8162), .A2(n8161), .ZN(n8085) );
  INV_X1 U10551 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9738) );
  INV_X1 U10552 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9727) );
  OR2_X1 U10553 ( .A1(n10724), .A2(n10869), .ZN(n14836) );
  AND2_X1 U10554 ( .A1(n8157), .A2(n8156), .ZN(n8086) );
  AND2_X1 U10555 ( .A1(n10438), .A2(n10432), .ZN(n8087) );
  INV_X1 U10556 ( .A(n15350), .ZN(n8968) );
  INV_X1 U10557 ( .A(n9089), .ZN(n9176) );
  AND2_X2 U10558 ( .A1(n15427), .A2(n15431), .ZN(n8088) );
  AND2_X1 U10559 ( .A1(n14984), .A2(n15580), .ZN(n8089) );
  AND2_X1 U10560 ( .A1(n15002), .A2(n8973), .ZN(n8090) );
  INV_X1 U10561 ( .A(n9835), .ZN(n13519) );
  AND2_X1 U10562 ( .A1(n8715), .A2(n8737), .ZN(n8091) );
  AND2_X1 U10563 ( .A1(n15866), .A2(n15886), .ZN(n13508) );
  NAND2_X1 U10564 ( .A1(n15918), .A2(n13499), .ZN(n13496) );
  AND2_X2 U10565 ( .A1(n11110), .A2(n10691), .ZN(n15918) );
  INV_X1 U10566 ( .A(n15918), .ZN(n10706) );
  INV_X1 U10567 ( .A(n14351), .ZN(n10518) );
  OR2_X1 U10568 ( .A1(n15906), .A2(n15901), .ZN(n13599) );
  INV_X1 U10569 ( .A(n13599), .ZN(n10701) );
  AND2_X1 U10570 ( .A1(n9580), .A2(n9579), .ZN(n15906) );
  INV_X1 U10571 ( .A(n14494), .ZN(n14498) );
  INV_X1 U10572 ( .A(n12916), .ZN(n9107) );
  INV_X1 U10573 ( .A(n13844), .ZN(n13845) );
  NOR2_X1 U10574 ( .A1(n8304), .A2(n8065), .ZN(n8305) );
  AND2_X1 U10575 ( .A1(n8578), .A2(n15134), .ZN(n8579) );
  NOR2_X1 U10576 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n8106) );
  INV_X1 U10577 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n8102) );
  OAI21_X1 U10578 ( .B1(n12526), .B2(n13034), .A(n12529), .ZN(n9809) );
  NAND2_X1 U10579 ( .A1(n14681), .A2(n9999), .ZN(n10000) );
  NAND2_X1 U10580 ( .A1(n8940), .A2(n8555), .ZN(n8941) );
  INV_X1 U10581 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8101) );
  NAND2_X1 U10582 ( .A1(n6530), .A2(n9842), .ZN(n9843) );
  OAI21_X1 U10583 ( .B1(n9812), .B2(n12530), .A(n9811), .ZN(n9813) );
  INV_X1 U10584 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10456) );
  INV_X1 U10585 ( .A(n14338), .ZN(n10516) );
  NAND2_X1 U10586 ( .A1(n10608), .A2(n10607), .ZN(n10610) );
  NAND2_X1 U10587 ( .A1(n14104), .A2(n10379), .ZN(n10387) );
  AND2_X1 U10588 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n8094) );
  INV_X1 U10589 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n12346) );
  NAND2_X1 U10590 ( .A1(n8170), .A2(n11053), .ZN(n8175) );
  OR2_X1 U10591 ( .A1(n12239), .A2(n13381), .ZN(n9814) );
  INV_X1 U10592 ( .A(n11525), .ZN(n9791) );
  NAND2_X1 U10593 ( .A1(n13199), .A2(n12890), .ZN(n10677) );
  OR2_X1 U10594 ( .A1(n10687), .A2(n13006), .ZN(n11104) );
  INV_X1 U10595 ( .A(n13346), .ZN(n13347) );
  INV_X1 U10596 ( .A(n13416), .ZN(n13418) );
  OR2_X1 U10597 ( .A1(n9370), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9371) );
  INV_X1 U10598 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9203) );
  INV_X1 U10599 ( .A(n11761), .ZN(n11717) );
  INV_X1 U10600 ( .A(n10815), .ZN(n10812) );
  INV_X1 U10601 ( .A(n12235), .ZN(n12125) );
  NAND2_X1 U10602 ( .A1(n13816), .A2(n11364), .ZN(n11972) );
  OR2_X1 U10603 ( .A1(n10817), .A2(n11242), .ZN(n11273) );
  OR2_X1 U10604 ( .A1(n10337), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n10338) );
  XNOR2_X1 U10605 ( .A(n9902), .B(n10111), .ZN(n9907) );
  INV_X1 U10606 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8478) );
  INV_X1 U10607 ( .A(n8775), .ZN(n8679) );
  NAND2_X1 U10608 ( .A1(n11319), .A2(n8775), .ZN(n8445) );
  AOI211_X1 U10609 ( .C1(n15278), .C2(n15555), .A(n15277), .B(n15276), .ZN(
        n15279) );
  INV_X1 U10610 ( .A(n15193), .ZN(n15211) );
  NOR2_X1 U10611 ( .A1(n8719), .A2(n8718), .ZN(n8720) );
  INV_X1 U10612 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n9744) );
  INV_X1 U10613 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n9755) );
  INV_X1 U10614 ( .A(n13349), .ZN(n13322) );
  NAND2_X1 U10615 ( .A1(n9856), .A2(n13601), .ZN(n9852) );
  AND2_X1 U10616 ( .A1(n9408), .A2(n9407), .ZN(n12801) );
  INV_X1 U10617 ( .A(n11740), .ZN(n9662) );
  INV_X1 U10618 ( .A(n15849), .ZN(n13144) );
  INV_X1 U10619 ( .A(n13612), .ZN(n13164) );
  INV_X1 U10620 ( .A(n13259), .ZN(n13237) );
  INV_X1 U10621 ( .A(n13034), .ZN(n13402) );
  INV_X1 U10622 ( .A(n12924), .ZN(n12884) );
  INV_X1 U10623 ( .A(n13023), .ZN(n15853) );
  OR2_X1 U10624 ( .A1(n11105), .A2(n11101), .ZN(n10686) );
  AND2_X1 U10625 ( .A1(n13307), .A2(n9523), .ZN(n9524) );
  INV_X1 U10626 ( .A(n15864), .ZN(n13401) );
  AND2_X1 U10627 ( .A1(n9539), .A2(n9538), .ZN(n15866) );
  INV_X1 U10628 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n13741) );
  OR2_X1 U10629 ( .A1(n10822), .A2(n10820), .ZN(n13789) );
  NAND2_X1 U10630 ( .A1(n11246), .A2(n11245), .ZN(n15749) );
  NAND2_X1 U10631 ( .A1(n15781), .A2(n11800), .ZN(n14436) );
  OAI21_X1 U10632 ( .B1(n10349), .B2(n10348), .A(n15784), .ZN(n10806) );
  NAND2_X1 U10633 ( .A1(n10308), .A2(n10307), .ZN(n10309) );
  OR2_X1 U10634 ( .A1(n10247), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n10253) );
  NAND2_X1 U10635 ( .A1(n9891), .A2(n9890), .ZN(n14711) );
  XNOR2_X1 U10636 ( .A(n9898), .B(n9896), .ZN(n14712) );
  XNOR2_X1 U10637 ( .A(n9892), .B(n15535), .ZN(n8874) );
  AND2_X1 U10638 ( .A1(n11019), .A2(n8975), .ZN(n15580) );
  OR2_X1 U10639 ( .A1(n11384), .A2(n15199), .ZN(n11493) );
  OR2_X1 U10640 ( .A1(n10867), .A2(n8994), .ZN(n10655) );
  INV_X1 U10641 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10932) );
  INV_X1 U10642 ( .A(n12822), .ZN(n12834) );
  INV_X1 U10643 ( .A(n12842), .ZN(n12803) );
  AND2_X1 U10644 ( .A1(n12861), .A2(n12860), .ZN(n13185) );
  AND2_X1 U10645 ( .A1(n9330), .A2(n9329), .ZN(n13323) );
  OR3_X1 U10646 ( .A1(n13620), .A2(n9558), .A3(n13616), .ZN(n9856) );
  OR2_X1 U10647 ( .A1(n9689), .A2(n9608), .ZN(n9687) );
  INV_X1 U10648 ( .A(n13182), .ZN(n13097) );
  INV_X1 U10649 ( .A(n13171), .ZN(n13152) );
  NAND2_X1 U10650 ( .A1(n11106), .A2(n15853), .ZN(n15855) );
  INV_X1 U10651 ( .A(n13496), .ZN(n13488) );
  AND2_X1 U10652 ( .A1(n10686), .A2(n10685), .ZN(n11110) );
  AND2_X1 U10653 ( .A1(n13015), .A2(n12874), .ZN(n13200) );
  INV_X1 U10654 ( .A(n13369), .ZN(n13379) );
  INV_X1 U10655 ( .A(n13508), .ZN(n15899) );
  NOR2_X1 U10656 ( .A1(n10973), .A2(n10972), .ZN(n10975) );
  INV_X1 U10657 ( .A(n13789), .ZN(n13730) );
  OR2_X1 U10658 ( .A1(n15792), .A2(n11787), .ZN(n10822) );
  INV_X1 U10659 ( .A(n11232), .ZN(n15690) );
  INV_X1 U10660 ( .A(n14152), .ZN(n15713) );
  AND2_X1 U10661 ( .A1(n11264), .A2(n14071), .ZN(n15752) );
  INV_X1 U10662 ( .A(n15776), .ZN(n15762) );
  INV_X1 U10663 ( .A(n14425), .ZN(n15759) );
  INV_X1 U10664 ( .A(n14421), .ZN(n15771) );
  AND2_X1 U10665 ( .A1(n14491), .A2(n14490), .ZN(n14613) );
  INV_X1 U10666 ( .A(n15817), .ZN(n15835) );
  AND2_X1 U10667 ( .A1(n10806), .A2(n10355), .ZN(n10359) );
  INV_X1 U10668 ( .A(n10232), .ZN(n10239) );
  AND2_X1 U10669 ( .A1(n8804), .A2(n8803), .ZN(n8805) );
  INV_X1 U10670 ( .A(n12220), .ZN(n14965) );
  INV_X1 U10671 ( .A(n12225), .ZN(n14962) );
  INV_X1 U10672 ( .A(n15571), .ZN(n15555) );
  OAI21_X1 U10673 ( .B1(n15286), .B2(n15262), .A(n10672), .ZN(n10673) );
  INV_X1 U10674 ( .A(n15172), .ZN(n15191) );
  INV_X1 U10675 ( .A(n15517), .ZN(n15239) );
  INV_X1 U10676 ( .A(n15578), .ZN(n15560) );
  INV_X1 U10677 ( .A(n11493), .ZN(n15552) );
  AND2_X1 U10678 ( .A1(n10654), .A2(n10656), .ZN(n9001) );
  NAND2_X1 U10679 ( .A1(n8982), .A2(n10868), .ZN(n10867) );
  AND2_X1 U10680 ( .A1(n8819), .A2(n8818), .ZN(n10868) );
  INV_X1 U10681 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8209) );
  INV_X1 U10682 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9723) );
  AND2_X1 U10683 ( .A1(n9689), .A2(n9688), .ZN(n15849) );
  INV_X1 U10684 ( .A(n12832), .ZN(n12815) );
  NAND2_X1 U10685 ( .A1(n9853), .A2(n11106), .ZN(n12842) );
  INV_X1 U10686 ( .A(n12756), .ZN(n13234) );
  INV_X1 U10687 ( .A(n13173), .ZN(n13146) );
  INV_X1 U10688 ( .A(n13180), .ZN(n13101) );
  NAND2_X1 U10689 ( .A1(n9611), .A2(n9610), .ZN(n13182) );
  AOI21_X1 U10690 ( .B1(n13222), .B2(n15864), .A(n13221), .ZN(n13440) );
  NAND2_X1 U10691 ( .A1(n15870), .A2(n11534), .ZN(n13431) );
  NAND2_X1 U10692 ( .A1(n15899), .A2(n15918), .ZN(n13491) );
  NAND2_X1 U10693 ( .A1(n13207), .A2(n10701), .ZN(n10702) );
  OR2_X1 U10694 ( .A1(n15906), .A2(n13508), .ZN(n13593) );
  NAND2_X1 U10695 ( .A1(n9193), .A2(n9192), .ZN(n13598) );
  INV_X2 U10696 ( .A(n15906), .ZN(n15905) );
  NAND2_X1 U10697 ( .A1(n9556), .A2(n9555), .ZN(n11105) );
  INV_X1 U10698 ( .A(SI_17_), .ZN(n11067) );
  INV_X1 U10699 ( .A(SI_12_), .ZN(n10915) );
  INV_X1 U10700 ( .A(n11928), .ZN(n13622) );
  INV_X1 U10701 ( .A(n14588), .ZN(n14458) );
  INV_X1 U10702 ( .A(n13769), .ZN(n13803) );
  INV_X1 U10703 ( .A(n13718), .ZN(n14089) );
  INV_X1 U10704 ( .A(n14376), .ZN(n14339) );
  INV_X1 U10705 ( .A(n15600), .ZN(n15755) );
  INV_X1 U10706 ( .A(n15770), .ZN(n14461) );
  INV_X1 U10707 ( .A(n12056), .ZN(n14489) );
  NAND2_X1 U10708 ( .A1(n15781), .A2(n11793), .ZN(n14421) );
  NAND2_X1 U10709 ( .A1(n15848), .A2(n15812), .ZN(n14602) );
  AND2_X2 U10710 ( .A1(n10359), .A2(n10358), .ZN(n15848) );
  INV_X1 U10711 ( .A(n14329), .ZN(n14632) );
  NAND2_X1 U10712 ( .A1(n15838), .A2(n15812), .ZN(n14652) );
  NOR2_X1 U10713 ( .A1(n15793), .A2(n15784), .ZN(n15789) );
  INV_X1 U10714 ( .A(n15796), .ZN(n15793) );
  XNOR2_X1 U10715 ( .A(n10341), .B(n10340), .ZN(n12160) );
  INV_X1 U10716 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n11023) );
  INV_X1 U10717 ( .A(n10156), .ZN(n10157) );
  NAND2_X1 U10718 ( .A1(n11029), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15508) );
  INV_X1 U10719 ( .A(n14813), .ZN(n15496) );
  OR2_X1 U10720 ( .A1(n10887), .A2(n14971), .ZN(n12215) );
  AND2_X1 U10721 ( .A1(n11995), .A2(n11994), .ZN(n15387) );
  OR2_X1 U10722 ( .A1(n15599), .A2(n8997), .ZN(n8998) );
  AND2_X2 U10723 ( .A1(n9002), .A2(n8996), .ZN(n15599) );
  INV_X1 U10724 ( .A(n15599), .ZN(n15597) );
  OR2_X1 U10725 ( .A1(n15383), .A2(n15382), .ZN(n15418) );
  INV_X1 U10726 ( .A(n15588), .ZN(n15587) );
  AND2_X1 U10727 ( .A1(n10757), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10876) );
  INV_X1 U10728 ( .A(n8979), .ZN(n12565) );
  INV_X1 U10729 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11377) );
  INV_X1 U10730 ( .A(n13043), .ZN(P3_U3897) );
  NAND2_X1 U10731 ( .A1(n9584), .A2(n9583), .ZN(P3_U3455) );
  AND2_X1 U10732 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11237), .ZN(P2_U3947) );
  INV_X1 U10733 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8493) );
  INV_X1 U10734 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8582) );
  INV_X1 U10735 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14798) );
  INV_X1 U10736 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14738) );
  INV_X1 U10737 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14817) );
  INV_X1 U10738 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n10153) );
  NAND2_X1 U10739 ( .A1(n8684), .A2(n10153), .ZN(n8100) );
  NOR2_X1 U10740 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n8108) );
  NAND4_X1 U10741 ( .A1(n8108), .A2(n8107), .A3(n8210), .A4(n8211), .ZN(n8815)
         );
  INV_X1 U10742 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n8114) );
  NAND2_X1 U10743 ( .A1(n8764), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8113) );
  NAND2_X1 U10744 ( .A1(n6514), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8112) );
  OAI211_X1 U10745 ( .C1(n8114), .C2(n8768), .A(n8113), .B(n8112), .ZN(n8115)
         );
  INV_X1 U10746 ( .A(n8115), .ZN(n8116) );
  INV_X1 U10747 ( .A(n14837), .ZN(n14816) );
  AND2_X1 U10748 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8118) );
  NAND2_X1 U10749 ( .A1(n8125), .A2(n8118), .ZN(n8247) );
  AND2_X1 U10750 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8119) );
  INV_X1 U10751 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10906) );
  NAND2_X1 U10752 ( .A1(n8132), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8120) );
  INV_X1 U10753 ( .A(SI_1_), .ZN(n10850) );
  OAI211_X1 U10754 ( .C1(n8132), .C2(n10906), .A(n8120), .B(n10850), .ZN(n8121) );
  OAI211_X1 U10755 ( .C1(P2_DATAO_REG_1__SCAN_IN), .C2(n8132), .A(n8122), .B(
        SI_1_), .ZN(n8123) );
  NAND2_X1 U10756 ( .A1(n8279), .A2(n8280), .ZN(n8127) );
  INV_X1 U10757 ( .A(SI_2_), .ZN(n10854) );
  NAND2_X1 U10758 ( .A1(n8127), .A2(n8076), .ZN(n8273) );
  MUX2_X1 U10759 ( .A(n12296), .B(n10839), .S(n8132), .Z(n8128) );
  NAND2_X1 U10760 ( .A1(n8273), .A2(n8275), .ZN(n8131) );
  INV_X1 U10761 ( .A(n8128), .ZN(n8129) );
  NAND2_X1 U10762 ( .A1(n8129), .A2(SI_3_), .ZN(n8130) );
  MUX2_X1 U10763 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n8132), .Z(n8134) );
  XNOR2_X1 U10764 ( .A(n8134), .B(SI_4_), .ZN(n8235) );
  INV_X1 U10765 ( .A(n8235), .ZN(n8133) );
  NAND2_X1 U10766 ( .A1(n8234), .A2(n8133), .ZN(n8136) );
  NAND2_X1 U10767 ( .A1(n8134), .A2(SI_4_), .ZN(n8135) );
  NAND2_X1 U10768 ( .A1(n8137), .A2(SI_5_), .ZN(n8138) );
  NAND2_X1 U10769 ( .A1(n8140), .A2(SI_6_), .ZN(n8141) );
  MUX2_X1 U10770 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n10878), .Z(n8143) );
  XNOR2_X1 U10771 ( .A(n8143), .B(SI_7_), .ZN(n8327) );
  INV_X1 U10772 ( .A(n8327), .ZN(n8142) );
  INV_X1 U10773 ( .A(n8346), .ZN(n8145) );
  MUX2_X1 U10774 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10878), .Z(n8376) );
  NAND2_X1 U10775 ( .A1(n8376), .A2(SI_9_), .ZN(n8392) );
  NAND2_X1 U10776 ( .A1(n8146), .A2(SI_8_), .ZN(n8374) );
  MUX2_X1 U10777 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10878), .Z(n8148) );
  XNOR2_X1 U10778 ( .A(n8148), .B(SI_10_), .ZN(n8394) );
  NAND2_X1 U10779 ( .A1(n8148), .A2(SI_10_), .ZN(n8149) );
  MUX2_X1 U10780 ( .A(n12309), .B(n10967), .S(n10878), .Z(n8150) );
  INV_X1 U10781 ( .A(n8150), .ZN(n8151) );
  NAND2_X1 U10782 ( .A1(n8151), .A2(SI_11_), .ZN(n8152) );
  NAND2_X1 U10783 ( .A1(n8153), .A2(n8152), .ZN(n8414) );
  MUX2_X1 U10784 ( .A(n9236), .B(n11023), .S(n10878), .Z(n8154) );
  NAND2_X1 U10785 ( .A1(n8154), .A2(n10915), .ZN(n8157) );
  INV_X1 U10786 ( .A(n8154), .ZN(n8155) );
  NAND2_X1 U10787 ( .A1(n8155), .A2(SI_12_), .ZN(n8156) );
  MUX2_X1 U10788 ( .A(n11047), .B(n11051), .S(n10878), .Z(n8159) );
  NAND2_X1 U10789 ( .A1(n8159), .A2(n10999), .ZN(n8162) );
  INV_X1 U10790 ( .A(n8159), .ZN(n8160) );
  NAND2_X1 U10791 ( .A1(n8160), .A2(SI_13_), .ZN(n8161) );
  MUX2_X1 U10792 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n10878), .Z(n8468) );
  MUX2_X1 U10793 ( .A(n11377), .B(n12274), .S(n10878), .Z(n8165) );
  INV_X1 U10794 ( .A(n8520), .ZN(n8163) );
  INV_X1 U10795 ( .A(n8165), .ZN(n8166) );
  NAND2_X1 U10796 ( .A1(n8166), .A2(SI_15_), .ZN(n8167) );
  NAND2_X1 U10797 ( .A1(n8520), .A2(n8167), .ZN(n8470) );
  INV_X1 U10798 ( .A(n8468), .ZN(n8168) );
  INV_X1 U10799 ( .A(n8517), .ZN(n8173) );
  MUX2_X1 U10800 ( .A(n11214), .B(n11217), .S(n10878), .Z(n8170) );
  INV_X1 U10801 ( .A(n8170), .ZN(n8171) );
  NAND2_X1 U10802 ( .A1(n8171), .A2(SI_16_), .ZN(n8172) );
  NAND2_X1 U10803 ( .A1(n8175), .A2(n8172), .ZN(n8522) );
  AOI21_X1 U10804 ( .B1(n8173), .B2(n8520), .A(n8522), .ZN(n8174) );
  MUX2_X1 U10805 ( .A(n12251), .B(n7796), .S(n10878), .Z(n8530) );
  MUX2_X1 U10806 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n10878), .Z(n8501) );
  MUX2_X1 U10807 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10878), .Z(n8564) );
  AOI22_X1 U10808 ( .A1(n8501), .A2(SI_18_), .B1(n8564), .B2(SI_19_), .ZN(
        n8176) );
  OAI21_X1 U10809 ( .B1(n8501), .B2(SI_18_), .A(SI_19_), .ZN(n8179) );
  INV_X1 U10810 ( .A(n8564), .ZN(n8178) );
  NOR2_X1 U10811 ( .A1(SI_18_), .A2(SI_19_), .ZN(n8177) );
  INV_X1 U10812 ( .A(n8501), .ZN(n8503) );
  AOI22_X1 U10813 ( .A1(n8179), .A2(n8178), .B1(n8177), .B2(n8503), .ZN(n8180)
         );
  MUX2_X1 U10814 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n10878), .Z(n8605) );
  NAND2_X1 U10815 ( .A1(n8605), .A2(SI_20_), .ZN(n8181) );
  MUX2_X1 U10816 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n10878), .Z(n8182) );
  OAI21_X1 U10817 ( .B1(n8182), .B2(SI_21_), .A(n8185), .ZN(n8606) );
  NOR2_X1 U10818 ( .A1(n8605), .A2(SI_20_), .ZN(n8183) );
  NOR2_X1 U10819 ( .A1(n8606), .A2(n8183), .ZN(n8184) );
  INV_X1 U10820 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8188) );
  MUX2_X1 U10821 ( .A(n8188), .B(n11873), .S(n10878), .Z(n10282) );
  MUX2_X1 U10822 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10878), .Z(n8190) );
  NAND2_X1 U10823 ( .A1(n8190), .A2(SI_23_), .ZN(n8191) );
  OAI21_X1 U10824 ( .B1(SI_23_), .B2(n8190), .A(n8191), .ZN(n8638) );
  MUX2_X1 U10825 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n10878), .Z(n8192) );
  NAND2_X1 U10826 ( .A1(n8192), .A2(SI_24_), .ZN(n8194) );
  OAI21_X1 U10827 ( .B1(n8192), .B2(SI_24_), .A(n8194), .ZN(n8193) );
  INV_X1 U10828 ( .A(n8193), .ZN(n8646) );
  MUX2_X1 U10829 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n10878), .Z(n8195) );
  XNOR2_X1 U10830 ( .A(n8195), .B(SI_25_), .ZN(n8668) );
  MUX2_X1 U10831 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n10878), .Z(n8196) );
  NAND2_X1 U10832 ( .A1(n8196), .A2(SI_26_), .ZN(n8197) );
  OAI21_X1 U10833 ( .B1(n8196), .B2(SI_26_), .A(n8197), .ZN(n8675) );
  MUX2_X1 U10834 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n10878), .Z(n8703) );
  XNOR2_X1 U10835 ( .A(n8703), .B(SI_27_), .ZN(n8198) );
  NAND2_X1 U10836 ( .A1(n8202), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8200) );
  NAND2_X1 U10837 ( .A1(n8818), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8201) );
  NAND2_X2 U10838 ( .A1(n8821), .A2(n15433), .ZN(n8248) );
  AND2_X4 U10839 ( .A1(n8248), .A2(n10879), .ZN(n8775) );
  NAND2_X1 U10840 ( .A1(n14668), .A2(n8775), .ZN(n8204) );
  AND2_X2 U10841 ( .A1(n8248), .A2(n10878), .ZN(n8282) );
  NAND2_X1 U10842 ( .A1(n8776), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8203) );
  INV_X1 U10843 ( .A(n8205), .ZN(n8206) );
  NAND2_X1 U10844 ( .A1(n8792), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8213) );
  INV_X1 U10845 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8212) );
  MUX2_X1 U10846 ( .A(n14816), .B(n7840), .S(n8779), .Z(n8697) );
  INV_X4 U10847 ( .A(n8248), .ZN(n10756) );
  INV_X1 U10848 ( .A(n8216), .ZN(n8271) );
  INV_X1 U10849 ( .A(n8236), .ZN(n8218) );
  NAND2_X1 U10850 ( .A1(n8218), .A2(n8217), .ZN(n8321) );
  NAND2_X1 U10851 ( .A1(n8321), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8219) );
  XNOR2_X1 U10852 ( .A(n8219), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10924) );
  AOI22_X1 U10853 ( .A1(n8282), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n10756), 
        .B2(n10924), .ZN(n8220) );
  NAND2_X1 U10854 ( .A1(n8088), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8227) );
  INV_X1 U10855 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n8221) );
  OR2_X1 U10856 ( .A1(n8688), .A2(n8221), .ZN(n8226) );
  INV_X1 U10857 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8222) );
  NAND2_X1 U10858 ( .A1(n8228), .A2(n8222), .ZN(n8223) );
  NAND2_X1 U10859 ( .A1(n8312), .A2(n8223), .ZN(n11494) );
  OR2_X1 U10860 ( .A1(n8750), .A2(n11494), .ZN(n8225) );
  INV_X1 U10861 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n11495) );
  OR2_X1 U10862 ( .A1(n8623), .A2(n11495), .ZN(n8224) );
  XNOR2_X1 U10863 ( .A(n11500), .B(n11564), .ZN(n8883) );
  NAND2_X1 U10864 ( .A1(n6514), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8233) );
  OAI21_X1 U10865 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(P1_REG3_REG_4__SCAN_IN), 
        .A(n8228), .ZN(n11392) );
  OR2_X1 U10866 ( .A1(n8750), .A2(n11392), .ZN(n8232) );
  INV_X1 U10867 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n8229) );
  OR2_X1 U10868 ( .A1(n8768), .A2(n8229), .ZN(n8231) );
  INV_X1 U10869 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11389) );
  OR2_X1 U10870 ( .A1(n8623), .A2(n11389), .ZN(n8230) );
  INV_X1 U10871 ( .A(n11489), .ZN(n14853) );
  XNOR2_X1 U10872 ( .A(n8234), .B(n8235), .ZN(n10859) );
  NAND2_X1 U10873 ( .A1(n10859), .A2(n8775), .ZN(n8239) );
  NAND2_X1 U10874 ( .A1(n8236), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8237) );
  XNOR2_X1 U10875 ( .A(n8237), .B(P1_IR_REG_4__SCAN_IN), .ZN(n14904) );
  AOI22_X1 U10876 ( .A1(n8282), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n10756), 
        .B2(n14904), .ZN(n8238) );
  NAND2_X1 U10877 ( .A1(n8239), .A2(n8238), .ZN(n15554) );
  INV_X1 U10878 ( .A(n15554), .ZN(n11393) );
  NAND3_X1 U10879 ( .A1(n14853), .A2(n11393), .A3(n8780), .ZN(n8241) );
  NAND3_X1 U10880 ( .A1(n11489), .A2(n8779), .A3(n15554), .ZN(n8240) );
  AND2_X1 U10881 ( .A1(n8241), .A2(n8240), .ZN(n8311) );
  NAND2_X1 U10882 ( .A1(n8763), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n8244) );
  NAND2_X1 U10883 ( .A1(n8088), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8243) );
  NAND2_X1 U10884 ( .A1(n8764), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8242) );
  INV_X1 U10885 ( .A(SI_0_), .ZN(n10836) );
  INV_X1 U10886 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9028) );
  OAI21_X1 U10887 ( .B1(n10878), .B2(n10836), .A(n9028), .ZN(n8246) );
  AND2_X1 U10888 ( .A1(n8247), .A2(n8246), .ZN(n15442) );
  MUX2_X1 U10889 ( .A(P1_IR_REG_0__SCAN_IN), .B(n15442), .S(n8248), .Z(n11055)
         );
  NAND2_X1 U10890 ( .A1(n14856), .A2(n8966), .ZN(n8828) );
  NAND2_X1 U10891 ( .A1(n8249), .A2(n8828), .ZN(n8251) );
  NAND2_X1 U10892 ( .A1(n8775), .A2(n8253), .ZN(n8257) );
  NAND2_X1 U10893 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8254) );
  NAND2_X1 U10894 ( .A1(n10756), .A2(n14859), .ZN(n8256) );
  NAND2_X1 U10895 ( .A1(n8282), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8255) );
  NAND3_X2 U10896 ( .A1(n8260), .A2(n8259), .A3(n8258), .ZN(n9892) );
  OAI21_X1 U10897 ( .B1(n15535), .B2(n8262), .A(n8264), .ZN(n8263) );
  INV_X1 U10898 ( .A(n8264), .ZN(n8265) );
  NAND2_X1 U10899 ( .A1(n8265), .A2(n8875), .ZN(n8266) );
  NAND2_X1 U10900 ( .A1(n6514), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8270) );
  NAND2_X1 U10901 ( .A1(n8088), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8268) );
  NAND2_X1 U10902 ( .A1(n8764), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8267) );
  INV_X1 U10903 ( .A(n14854), .ZN(n11348) );
  NAND2_X1 U10904 ( .A1(n8271), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8272) );
  XNOR2_X1 U10905 ( .A(n8272), .B(P1_IR_REG_3__SCAN_IN), .ZN(n14892) );
  AOI22_X1 U10906 ( .A1(n8282), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n10756), 
        .B2(n14892), .ZN(n8278) );
  XNOR2_X1 U10907 ( .A(n8275), .B(n8276), .ZN(n10838) );
  NAND2_X1 U10908 ( .A1(n10838), .A2(n8775), .ZN(n8277) );
  INV_X1 U10909 ( .A(n15502), .ZN(n11472) );
  XNOR2_X1 U10910 ( .A(n8279), .B(n8280), .ZN(n10881) );
  INV_X1 U10911 ( .A(n10881), .ZN(n8281) );
  NAND2_X1 U10912 ( .A1(n8775), .A2(n8281), .ZN(n8288) );
  NAND2_X1 U10913 ( .A1(n8282), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8287) );
  INV_X1 U10914 ( .A(n8283), .ZN(n8284) );
  NAND2_X1 U10915 ( .A1(n8284), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8285) );
  NAND2_X1 U10916 ( .A1(n10756), .A2(n14879), .ZN(n8286) );
  AND3_X2 U10917 ( .A1(n8288), .A2(n8287), .A3(n8286), .ZN(n8299) );
  NAND3_X1 U10918 ( .A1(n8919), .A2(n8299), .A3(n8780), .ZN(n8295) );
  NAND2_X1 U10919 ( .A1(n14854), .A2(n15502), .ZN(n8298) );
  NAND2_X1 U10920 ( .A1(n8763), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n8291) );
  NAND2_X1 U10921 ( .A1(n8088), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8290) );
  NAND2_X1 U10922 ( .A1(n8764), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n8289) );
  INV_X1 U10923 ( .A(n14855), .ZN(n8293) );
  NAND3_X1 U10924 ( .A1(n8298), .A2(n8293), .A3(n8779), .ZN(n8294) );
  AND4_X1 U10925 ( .A1(n8919), .A2(n8298), .A3(n14855), .A4(n6516), .ZN(n8296)
         );
  NAND2_X1 U10926 ( .A1(n8298), .A2(n8779), .ZN(n8301) );
  NAND4_X1 U10927 ( .A1(n8919), .A2(n8299), .A3(n8780), .A4(n14855), .ZN(n8300) );
  OAI21_X1 U10928 ( .B1(n8301), .B2(n8918), .A(n8300), .ZN(n8304) );
  NAND2_X1 U10929 ( .A1(n8919), .A2(n8780), .ZN(n8302) );
  NAND2_X1 U10930 ( .A1(n8302), .A2(n8301), .ZN(n8303) );
  XNOR2_X1 U10931 ( .A(n14854), .B(n15502), .ZN(n11070) );
  NAND3_X1 U10932 ( .A1(n8307), .A2(n8306), .A3(n8305), .ZN(n8308) );
  INV_X1 U10933 ( .A(n8883), .ZN(n11487) );
  XNOR2_X1 U10934 ( .A(n11489), .B(n15554), .ZN(n8881) );
  NOR2_X1 U10935 ( .A1(n11564), .A2(n8779), .ZN(n8309) );
  NAND2_X1 U10936 ( .A1(n6514), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8318) );
  INV_X1 U10937 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11574) );
  OR2_X1 U10938 ( .A1(n8623), .A2(n11574), .ZN(n8317) );
  INV_X1 U10939 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n11516) );
  NAND2_X1 U10940 ( .A1(n8312), .A2(n11516), .ZN(n8313) );
  NAND2_X1 U10941 ( .A1(n8335), .A2(n8313), .ZN(n11573) );
  OR2_X1 U10942 ( .A1(n8750), .A2(n11573), .ZN(n8316) );
  INV_X1 U10943 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n8314) );
  OR2_X1 U10944 ( .A1(n8768), .A2(n8314), .ZN(n8315) );
  INV_X1 U10945 ( .A(n11703), .ZN(n14851) );
  XNOR2_X1 U10946 ( .A(n8319), .B(n8320), .ZN(n10882) );
  NAND2_X1 U10947 ( .A1(n10882), .A2(n8775), .ZN(n8324) );
  NAND2_X1 U10948 ( .A1(n8328), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8322) );
  XNOR2_X1 U10949 ( .A(n8322), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10939) );
  AOI22_X1 U10950 ( .A1(n8282), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n10756), 
        .B2(n10939), .ZN(n8323) );
  NAND2_X1 U10951 ( .A1(n8324), .A2(n8323), .ZN(n11576) );
  MUX2_X1 U10952 ( .A(n14851), .B(n11576), .S(n8779), .Z(n8342) );
  MUX2_X1 U10953 ( .A(n14851), .B(n11576), .S(n8261), .Z(n8325) );
  XNOR2_X1 U10954 ( .A(n8326), .B(n8327), .ZN(n10904) );
  NAND2_X1 U10955 ( .A1(n10904), .A2(n8775), .ZN(n8333) );
  INV_X1 U10956 ( .A(n8328), .ZN(n8330) );
  NAND2_X1 U10957 ( .A1(n8330), .A2(n8329), .ZN(n8348) );
  NAND2_X1 U10958 ( .A1(n8348), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8331) );
  XNOR2_X1 U10959 ( .A(n8331), .B(P1_IR_REG_7__SCAN_IN), .ZN(n14918) );
  AOI22_X1 U10960 ( .A1(n8282), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n10756), 
        .B2(n14918), .ZN(n8332) );
  NAND2_X1 U10961 ( .A1(n6514), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8341) );
  INV_X1 U10962 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n8334) );
  OR2_X1 U10963 ( .A1(n8623), .A2(n8334), .ZN(n8340) );
  INV_X1 U10964 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n12302) );
  NAND2_X1 U10965 ( .A1(n8335), .A2(n12302), .ZN(n8336) );
  NAND2_X1 U10966 ( .A1(n8354), .A2(n8336), .ZN(n15512) );
  OR2_X1 U10967 ( .A1(n8750), .A2(n15512), .ZN(n8339) );
  INV_X1 U10968 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n8337) );
  OR2_X1 U10969 ( .A1(n8768), .A2(n8337), .ZN(n8338) );
  XNOR2_X1 U10970 ( .A(n11700), .B(n14849), .ZN(n8827) );
  NOR2_X1 U10971 ( .A1(n11677), .A2(n8779), .ZN(n8344) );
  OAI21_X1 U10972 ( .B1(n14849), .B2(n8261), .A(n11700), .ZN(n8343) );
  OAI21_X1 U10973 ( .B1(n8344), .B2(n11700), .A(n8343), .ZN(n8345) );
  NAND2_X1 U10974 ( .A1(n10911), .A2(n8775), .ZN(n8351) );
  NAND2_X1 U10975 ( .A1(n8377), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8349) );
  XNOR2_X1 U10976 ( .A(n8349), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U10977 ( .A1(n8282), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n10959), 
        .B2(n10756), .ZN(n8350) );
  NAND2_X2 U10978 ( .A1(n8351), .A2(n8350), .ZN(n15581) );
  NAND2_X1 U10979 ( .A1(n8764), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8360) );
  INV_X1 U10980 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n8352) );
  OR2_X1 U10981 ( .A1(n8688), .A2(n8352), .ZN(n8359) );
  INV_X1 U10982 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8353) );
  NAND2_X1 U10983 ( .A1(n8354), .A2(n8353), .ZN(n8355) );
  NAND2_X1 U10984 ( .A1(n8367), .A2(n8355), .ZN(n11868) );
  OR2_X1 U10985 ( .A1(n8750), .A2(n11868), .ZN(n8358) );
  INV_X1 U10986 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n8356) );
  OR2_X1 U10987 ( .A1(n8768), .A2(n8356), .ZN(n8357) );
  NAND2_X1 U10988 ( .A1(n15581), .A2(n11832), .ZN(n8826) );
  MUX2_X1 U10989 ( .A(n8826), .B(n8926), .S(n8779), .Z(n8361) );
  NAND2_X1 U10990 ( .A1(n8362), .A2(n8361), .ZN(n8365) );
  INV_X1 U10991 ( .A(n11832), .ZN(n14848) );
  MUX2_X1 U10992 ( .A(n14848), .B(n15581), .S(n8261), .Z(n8363) );
  OR2_X1 U10993 ( .A1(n6664), .A2(n8363), .ZN(n8364) );
  NAND2_X1 U10994 ( .A1(n8365), .A2(n8364), .ZN(n8382) );
  NAND2_X1 U10995 ( .A1(n8764), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n8373) );
  INV_X1 U10996 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10735) );
  OR2_X1 U10997 ( .A1(n8688), .A2(n10735), .ZN(n8372) );
  NAND2_X1 U10998 ( .A1(n8367), .A2(n8366), .ZN(n8368) );
  NAND2_X1 U10999 ( .A1(n8407), .A2(n8368), .ZN(n12065) );
  OR2_X1 U11000 ( .A1(n8750), .A2(n12065), .ZN(n8371) );
  INV_X1 U11001 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n8369) );
  OR2_X1 U11002 ( .A1(n8768), .A2(n8369), .ZN(n8370) );
  XNOR2_X1 U11003 ( .A(n8376), .B(SI_9_), .ZN(n8389) );
  NAND2_X1 U11004 ( .A1(n10222), .A2(n8775), .ZN(n8379) );
  NAND2_X1 U11005 ( .A1(n8415), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8397) );
  XNOR2_X1 U11006 ( .A(n8397), .B(P1_IR_REG_9__SCAN_IN), .ZN(n11006) );
  AOI22_X1 U11007 ( .A1(n11006), .A2(n10756), .B1(n8776), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n8378) );
  NAND2_X2 U11008 ( .A1(n8379), .A2(n8378), .ZN(n15396) );
  INV_X1 U11009 ( .A(n15396), .ZN(n11837) );
  MUX2_X1 U11010 ( .A(n12183), .B(n11837), .S(n8261), .Z(n8381) );
  INV_X1 U11011 ( .A(n12183), .ZN(n14847) );
  MUX2_X1 U11012 ( .A(n14847), .B(n15396), .S(n8779), .Z(n8380) );
  NAND2_X1 U11013 ( .A1(n8382), .A2(n8381), .ZN(n8383) );
  NAND2_X1 U11014 ( .A1(n6514), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8388) );
  INV_X1 U11015 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n8384) );
  OR2_X1 U11016 ( .A1(n8768), .A2(n8384), .ZN(n8387) );
  INV_X1 U11017 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8406) );
  XNOR2_X1 U11018 ( .A(n8407), .B(n8406), .ZN(n12182) );
  OR2_X1 U11019 ( .A1(n8750), .A2(n12182), .ZN(n8386) );
  INV_X1 U11020 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11923) );
  OR2_X1 U11021 ( .A1(n8623), .A2(n11923), .ZN(n8385) );
  INV_X1 U11022 ( .A(n12169), .ZN(n14846) );
  INV_X1 U11023 ( .A(n8389), .ZN(n8390) );
  NAND2_X1 U11024 ( .A1(n8391), .A2(n8390), .ZN(n8393) );
  NAND2_X1 U11025 ( .A1(n10949), .A2(n8775), .ZN(n8401) );
  INV_X1 U11026 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8396) );
  NAND2_X1 U11027 ( .A1(n8397), .A2(n8396), .ZN(n8398) );
  NAND2_X1 U11028 ( .A1(n8398), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8399) );
  XNOR2_X1 U11029 ( .A(n8399), .B(P1_IR_REG_10__SCAN_IN), .ZN(n14934) );
  AOI22_X1 U11030 ( .A1(n14934), .A2(n10756), .B1(n8776), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n8400) );
  MUX2_X1 U11031 ( .A(n14846), .B(n15391), .S(n8779), .Z(n8403) );
  MUX2_X1 U11032 ( .A(n14846), .B(n15391), .S(n8261), .Z(n8402) );
  NAND2_X1 U11033 ( .A1(n8088), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8412) );
  INV_X1 U11034 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n12415) );
  OR2_X1 U11035 ( .A1(n8688), .A2(n12415), .ZN(n8411) );
  INV_X1 U11036 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8405) );
  OAI21_X1 U11037 ( .B1(n8407), .B2(n8406), .A(n8405), .ZN(n8408) );
  NAND2_X1 U11038 ( .A1(n8428), .A2(n8408), .ZN(n12168) );
  OR2_X1 U11039 ( .A1(n8750), .A2(n12168), .ZN(n8410) );
  INV_X1 U11040 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10771) );
  OR2_X1 U11041 ( .A1(n8623), .A2(n10771), .ZN(n8409) );
  INV_X1 U11042 ( .A(n14729), .ZN(n14845) );
  XNOR2_X1 U11043 ( .A(n8413), .B(n8414), .ZN(n10966) );
  NAND2_X1 U11044 ( .A1(n10966), .A2(n8775), .ZN(n8422) );
  INV_X1 U11045 ( .A(n8415), .ZN(n8417) );
  NOR2_X1 U11046 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n8416) );
  NAND2_X1 U11047 ( .A1(n8417), .A2(n8416), .ZN(n8419) );
  NAND2_X1 U11048 ( .A1(n8419), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8418) );
  MUX2_X1 U11049 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8418), .S(
        P1_IR_REG_11__SCAN_IN), .Z(n8420) );
  AOI22_X1 U11050 ( .A1(n11166), .A2(n10756), .B1(n8776), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n8421) );
  MUX2_X1 U11051 ( .A(n14845), .B(n15384), .S(n8780), .Z(n8425) );
  MUX2_X1 U11052 ( .A(n14845), .B(n15384), .S(n8779), .Z(n8423) );
  NAND2_X1 U11053 ( .A1(n8424), .A2(n8423), .ZN(n8427) );
  NAND2_X1 U11054 ( .A1(n6514), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8433) );
  INV_X1 U11055 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n12198) );
  OR2_X1 U11056 ( .A1(n8623), .A2(n12198), .ZN(n8432) );
  NAND2_X1 U11057 ( .A1(n8428), .A2(n12346), .ZN(n8429) );
  NAND2_X1 U11058 ( .A1(n8453), .A2(n8429), .ZN(n14728) );
  OR2_X1 U11059 ( .A1(n8750), .A2(n14728), .ZN(n8431) );
  INV_X1 U11060 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n12454) );
  OR2_X1 U11061 ( .A1(n8768), .A2(n12454), .ZN(n8430) );
  XNOR2_X1 U11062 ( .A(n8434), .B(n8086), .ZN(n11001) );
  NAND2_X1 U11063 ( .A1(n8435), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8441) );
  XNOR2_X1 U11064 ( .A(n8441), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11316) );
  AOI22_X1 U11065 ( .A1(n11316), .A2(n10756), .B1(n8776), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n8436) );
  MUX2_X1 U11066 ( .A(n15258), .B(n14724), .S(n8779), .Z(n8438) );
  MUX2_X1 U11067 ( .A(n15258), .B(n14724), .S(n8780), .Z(n8437) );
  INV_X1 U11068 ( .A(n8438), .ZN(n8439) );
  NAND2_X1 U11069 ( .A1(n8441), .A2(n8440), .ZN(n8442) );
  NAND2_X1 U11070 ( .A1(n8442), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8462) );
  INV_X1 U11071 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n12256) );
  NAND2_X1 U11072 ( .A1(n8462), .A2(n12256), .ZN(n8464) );
  NAND2_X1 U11073 ( .A1(n8464), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8443) );
  AOI22_X1 U11074 ( .A1(n11621), .A2(n10756), .B1(n8776), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8444) );
  NAND2_X1 U11075 ( .A1(n8455), .A2(n8446), .ZN(n8447) );
  NAND2_X1 U11076 ( .A1(n8479), .A2(n8447), .ZN(n15229) );
  OR2_X1 U11077 ( .A1(n15229), .A2(n8750), .ZN(n8451) );
  INV_X1 U11078 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n12280) );
  OR2_X1 U11079 ( .A1(n8768), .A2(n12280), .ZN(n8450) );
  NAND2_X1 U11080 ( .A1(n8764), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8449) );
  NAND2_X1 U11081 ( .A1(n6514), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8448) );
  NAND4_X1 U11082 ( .A1(n8451), .A2(n8450), .A3(n8449), .A4(n8448), .ZN(n15255) );
  NAND2_X1 U11083 ( .A1(n8965), .A2(n15213), .ZN(n8484) );
  NAND2_X1 U11084 ( .A1(n6514), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8460) );
  INV_X1 U11085 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n12441) );
  OR2_X1 U11086 ( .A1(n8623), .A2(n12441), .ZN(n8459) );
  INV_X1 U11087 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8452) );
  NAND2_X1 U11088 ( .A1(n8453), .A2(n8452), .ZN(n8454) );
  NAND2_X1 U11089 ( .A1(n8455), .A2(n8454), .ZN(n15260) );
  OR2_X1 U11090 ( .A1(n8750), .A2(n15260), .ZN(n8458) );
  INV_X1 U11091 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n8456) );
  OR2_X1 U11092 ( .A1(n8768), .A2(n8456), .ZN(n8457) );
  INV_X1 U11093 ( .A(n15226), .ZN(n14844) );
  XNOR2_X1 U11094 ( .A(n8461), .B(n8085), .ZN(n11046) );
  NAND2_X1 U11095 ( .A1(n11046), .A2(n8775), .ZN(n8466) );
  OR2_X1 U11096 ( .A1(n8462), .A2(n12256), .ZN(n8463) );
  AOI22_X1 U11097 ( .A1(n11601), .A2(n10756), .B1(n8776), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n8465) );
  MUX2_X1 U11098 ( .A(n14844), .B(n14788), .S(n8780), .Z(n8486) );
  NOR2_X1 U11099 ( .A1(n15226), .A2(n8779), .ZN(n8467) );
  AOI21_X1 U11100 ( .B1(n14788), .B2(n8779), .A(n8467), .ZN(n8485) );
  INV_X1 U11101 ( .A(n8470), .ZN(n8471) );
  XNOR2_X1 U11102 ( .A(n8472), .B(n8471), .ZN(n10259) );
  NAND2_X1 U11103 ( .A1(n10259), .A2(n8775), .ZN(n8477) );
  NAND2_X1 U11104 ( .A1(n8474), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8473) );
  MUX2_X1 U11105 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8473), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n8475) );
  OR2_X1 U11106 ( .A1(n8474), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n8525) );
  AND2_X1 U11107 ( .A1(n8475), .A2(n8525), .ZN(n11881) );
  AOI22_X1 U11108 ( .A1(n8282), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n10756), 
        .B2(n11881), .ZN(n8476) );
  NAND2_X2 U11109 ( .A1(n8477), .A2(n8476), .ZN(n8898) );
  NAND2_X1 U11110 ( .A1(n8479), .A2(n8478), .ZN(n8480) );
  AND2_X1 U11111 ( .A1(n8512), .A2(n8480), .ZN(n15215) );
  NAND2_X1 U11112 ( .A1(n15215), .A2(n8763), .ZN(n8483) );
  AOI22_X1 U11113 ( .A1(n8088), .A2(P1_REG0_REG_15__SCAN_IN), .B1(n6514), .B2(
        P1_REG1_REG_15__SCAN_IN), .ZN(n8482) );
  NAND2_X1 U11114 ( .A1(n8764), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n8481) );
  NAND2_X1 U11115 ( .A1(n8939), .A2(n8484), .ZN(n8488) );
  NOR2_X1 U11116 ( .A1(n8486), .A2(n8485), .ZN(n8487) );
  AOI22_X1 U11117 ( .A1(n8779), .A2(n8488), .B1(n15241), .B2(n8487), .ZN(n8489) );
  OR2_X2 U11118 ( .A1(n8898), .A2(n15228), .ZN(n8934) );
  INV_X1 U11119 ( .A(n8934), .ZN(n15171) );
  AOI21_X1 U11120 ( .B1(n8490), .B2(n8489), .A(n15171), .ZN(n8492) );
  AOI21_X1 U11121 ( .B1(n8934), .B2(n8933), .A(n8779), .ZN(n8491) );
  NAND2_X1 U11122 ( .A1(n8540), .A2(n8493), .ZN(n8494) );
  AND2_X1 U11123 ( .A1(n8570), .A2(n8494), .ZN(n15162) );
  NAND2_X1 U11124 ( .A1(n15162), .A2(n8763), .ZN(n8500) );
  INV_X1 U11125 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n8497) );
  NAND2_X1 U11126 ( .A1(n8764), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8496) );
  NAND2_X1 U11127 ( .A1(n6514), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8495) );
  OAI211_X1 U11128 ( .C1(n8497), .C2(n8768), .A(n8496), .B(n8495), .ZN(n8498)
         );
  INV_X1 U11129 ( .A(n8498), .ZN(n8499) );
  NAND2_X1 U11130 ( .A1(n8500), .A2(n8499), .ZN(n15140) );
  INV_X1 U11131 ( .A(n8525), .ZN(n8506) );
  INV_X1 U11132 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8505) );
  NAND2_X1 U11133 ( .A1(n8506), .A2(n8505), .ZN(n8532) );
  INV_X1 U11134 ( .A(n8532), .ZN(n8508) );
  INV_X1 U11135 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8507) );
  NAND2_X1 U11136 ( .A1(n8508), .A2(n8507), .ZN(n8534) );
  NAND2_X1 U11137 ( .A1(n8534), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8509) );
  XNOR2_X1 U11138 ( .A(n8509), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14961) );
  AOI22_X1 U11139 ( .A1(n8282), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n10756), 
        .B2(n14961), .ZN(n8510) );
  NAND2_X1 U11140 ( .A1(n15339), .A2(n15140), .ZN(n8904) );
  NAND2_X1 U11141 ( .A1(n8547), .A2(n8904), .ZN(n8545) );
  INV_X1 U11142 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n8516) );
  NAND2_X1 U11143 ( .A1(n8512), .A2(n6931), .ZN(n8513) );
  NAND2_X1 U11144 ( .A1(n8538), .A2(n8513), .ZN(n14749) );
  OR2_X1 U11145 ( .A1(n14749), .A2(n8750), .ZN(n8515) );
  AOI22_X1 U11146 ( .A1(n8764), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n6514), .B2(
        P1_REG1_REG_16__SCAN_IN), .ZN(n8514) );
  OAI211_X1 U11147 ( .C1(n8768), .C2(n8516), .A(n8515), .B(n8514), .ZN(n14842)
         );
  NAND2_X1 U11148 ( .A1(n8521), .A2(n8520), .ZN(n8524) );
  INV_X1 U11149 ( .A(n8522), .ZN(n8523) );
  XNOR2_X2 U11150 ( .A(n8524), .B(n8523), .ZN(n11213) );
  NAND2_X1 U11151 ( .A1(n11213), .A2(n8775), .ZN(n8528) );
  NAND2_X1 U11152 ( .A1(n8525), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8526) );
  XNOR2_X1 U11153 ( .A(n8526), .B(P1_IR_REG_16__SCAN_IN), .ZN(n11212) );
  AOI22_X1 U11154 ( .A1(n8776), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n10756), 
        .B2(n11212), .ZN(n8527) );
  NAND2_X2 U11155 ( .A1(n8528), .A2(n8527), .ZN(n15350) );
  MUX2_X1 U11156 ( .A(n14842), .B(n15350), .S(n8261), .Z(n8552) );
  NOR2_X1 U11157 ( .A1(n14842), .A2(n8779), .ZN(n8551) );
  NOR2_X1 U11158 ( .A1(n15350), .A2(n8261), .ZN(n8548) );
  OR3_X1 U11159 ( .A1(n8552), .A2(n8551), .A3(n8548), .ZN(n8544) );
  XNOR2_X1 U11160 ( .A(n8530), .B(SI_17_), .ZN(n8531) );
  XNOR2_X1 U11161 ( .A(n8529), .B(n8531), .ZN(n11446) );
  NAND2_X1 U11162 ( .A1(n11446), .A2(n8775), .ZN(n8537) );
  NAND2_X1 U11163 ( .A1(n8532), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8533) );
  MUX2_X1 U11164 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8533), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n8535) );
  NAND2_X1 U11165 ( .A1(n8535), .A2(n8534), .ZN(n11448) );
  INV_X1 U11166 ( .A(n11448), .ZN(n14947) );
  AOI22_X1 U11167 ( .A1(n8282), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n10756), 
        .B2(n14947), .ZN(n8536) );
  INV_X1 U11168 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n8543) );
  NAND2_X1 U11169 ( .A1(n8538), .A2(n6932), .ZN(n8539) );
  NAND2_X1 U11170 ( .A1(n8540), .A2(n8539), .ZN(n14758) );
  OR2_X1 U11171 ( .A1(n14758), .A2(n8750), .ZN(n8542) );
  AOI22_X1 U11172 ( .A1(n8764), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n6514), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n8541) );
  OAI211_X1 U11173 ( .C1(n8768), .C2(n8543), .A(n8542), .B(n8541), .ZN(n14841)
         );
  XNOR2_X1 U11174 ( .A(n15342), .B(n14841), .ZN(n15173) );
  INV_X1 U11175 ( .A(n8547), .ZN(n8561) );
  INV_X1 U11176 ( .A(n15342), .ZN(n15183) );
  AND2_X1 U11177 ( .A1(n15183), .A2(n14841), .ZN(n15154) );
  NAND2_X1 U11178 ( .A1(n15154), .A2(n8779), .ZN(n8550) );
  INV_X1 U11179 ( .A(n14841), .ZN(n15196) );
  NAND3_X1 U11180 ( .A1(n8552), .A2(n8548), .A3(n8067), .ZN(n8549) );
  AND2_X1 U11181 ( .A1(n8550), .A2(n8549), .ZN(n8557) );
  NAND2_X1 U11182 ( .A1(n8552), .A2(n8551), .ZN(n8554) );
  OR2_X1 U11183 ( .A1(n8067), .A2(n8779), .ZN(n8553) );
  NAND2_X1 U11184 ( .A1(n8554), .A2(n8553), .ZN(n8556) );
  INV_X1 U11185 ( .A(n15154), .ZN(n8555) );
  NAND2_X1 U11186 ( .A1(n8556), .A2(n8555), .ZN(n8558) );
  NAND3_X1 U11187 ( .A1(n8905), .A2(n8557), .A3(n8558), .ZN(n8560) );
  NAND2_X1 U11188 ( .A1(n8558), .A2(n8557), .ZN(n8559) );
  AOI22_X1 U11189 ( .A1(n8561), .A2(n8560), .B1(n8035), .B2(n8559), .ZN(n8578)
         );
  INV_X1 U11190 ( .A(SI_18_), .ZN(n11127) );
  OR2_X1 U11191 ( .A1(n8562), .A2(n11127), .ZN(n8563) );
  XNOR2_X1 U11192 ( .A(n8564), .B(SI_19_), .ZN(n8565) );
  AOI22_X1 U11193 ( .A1(n8282), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10756), 
        .B2(n15199), .ZN(n8567) );
  INV_X1 U11194 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U11195 ( .A1(n8570), .A2(n8569), .ZN(n8571) );
  NAND2_X1 U11196 ( .A1(n8583), .A2(n8571), .ZN(n14702) );
  OR2_X1 U11197 ( .A1(n14702), .A2(n8750), .ZN(n8577) );
  INV_X1 U11198 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n8574) );
  NAND2_X1 U11199 ( .A1(n8088), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U11200 ( .A1(n6514), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n8572) );
  OAI211_X1 U11201 ( .C1(n8623), .C2(n8574), .A(n8573), .B(n8572), .ZN(n8575)
         );
  INV_X1 U11202 ( .A(n8575), .ZN(n8576) );
  NAND2_X1 U11203 ( .A1(n8577), .A2(n8576), .ZN(n15116) );
  INV_X1 U11204 ( .A(n15116), .ZN(n14776) );
  OR2_X1 U11205 ( .A1(n15330), .A2(n14776), .ZN(n8580) );
  NAND2_X1 U11206 ( .A1(n15330), .A2(n14776), .ZN(n15095) );
  MUX2_X1 U11207 ( .A(n8580), .B(n15095), .S(n8779), .Z(n8581) );
  NAND2_X1 U11208 ( .A1(n8583), .A2(n8582), .ZN(n8584) );
  AND2_X1 U11209 ( .A1(n8598), .A2(n8584), .ZN(n15125) );
  NAND2_X1 U11210 ( .A1(n15125), .A2(n8763), .ZN(n8590) );
  INV_X1 U11211 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n8587) );
  NAND2_X1 U11212 ( .A1(n6514), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n8586) );
  NAND2_X1 U11213 ( .A1(n8764), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8585) );
  OAI211_X1 U11214 ( .C1(n8768), .C2(n8587), .A(n8586), .B(n8585), .ZN(n8588)
         );
  INV_X1 U11215 ( .A(n8588), .ZN(n8589) );
  NAND2_X1 U11216 ( .A1(n8590), .A2(n8589), .ZN(n15139) );
  INV_X1 U11217 ( .A(n15139), .ZN(n15098) );
  INV_X1 U11218 ( .A(SI_20_), .ZN(n11698) );
  NAND2_X1 U11219 ( .A1(n8591), .A2(n11698), .ZN(n8592) );
  NAND2_X1 U11220 ( .A1(n11827), .A2(n8775), .ZN(n8594) );
  NAND2_X1 U11221 ( .A1(n8776), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8593) );
  INV_X1 U11222 ( .A(n15324), .ZN(n15127) );
  MUX2_X1 U11223 ( .A(n15139), .B(n15324), .S(n8779), .Z(n8595) );
  INV_X1 U11224 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U11225 ( .A1(n8598), .A2(n8597), .ZN(n8599) );
  NAND2_X1 U11226 ( .A1(n8618), .A2(n8599), .ZN(n15104) );
  OR2_X1 U11227 ( .A1(n15104), .A2(n8750), .ZN(n8604) );
  INV_X1 U11228 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n12358) );
  NAND2_X1 U11229 ( .A1(n8764), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8601) );
  NAND2_X1 U11230 ( .A1(n8088), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8600) );
  OAI211_X1 U11231 ( .C1(n8688), .C2(n12358), .A(n8601), .B(n8600), .ZN(n8602)
         );
  INV_X1 U11232 ( .A(n8602), .ZN(n8603) );
  INV_X1 U11233 ( .A(n8605), .ZN(n8609) );
  NAND2_X1 U11234 ( .A1(n8612), .A2(n8611), .ZN(n11913) );
  NAND2_X1 U11235 ( .A1(n8776), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8613) );
  MUX2_X1 U11236 ( .A(n15117), .B(n15319), .S(n8779), .Z(n8617) );
  MUX2_X1 U11237 ( .A(n15117), .B(n15319), .S(n8261), .Z(n8615) );
  NAND2_X1 U11238 ( .A1(n8618), .A2(n14798), .ZN(n8619) );
  AND2_X1 U11239 ( .A1(n8630), .A2(n8619), .ZN(n15088) );
  NAND2_X1 U11240 ( .A1(n15088), .A2(n8763), .ZN(n8626) );
  INV_X1 U11241 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n8622) );
  NAND2_X1 U11242 ( .A1(n8088), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8621) );
  NAND2_X1 U11243 ( .A1(n6514), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8620) );
  OAI211_X1 U11244 ( .C1(n8623), .C2(n8622), .A(n8621), .B(n8620), .ZN(n8624)
         );
  INV_X1 U11245 ( .A(n8624), .ZN(n8625) );
  NAND2_X1 U11246 ( .A1(n8626), .A2(n8625), .ZN(n14840) );
  OR2_X1 U11247 ( .A1(n10283), .A2(n10878), .ZN(n8627) );
  INV_X1 U11248 ( .A(n15090), .ZN(n15314) );
  MUX2_X1 U11249 ( .A(n14840), .B(n15314), .S(n8780), .Z(n8629) );
  MUX2_X1 U11250 ( .A(n15099), .B(n15090), .S(n8779), .Z(n8628) );
  INV_X1 U11251 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14695) );
  NAND2_X1 U11252 ( .A1(n8630), .A2(n14695), .ZN(n8631) );
  NAND2_X1 U11253 ( .A1(n8651), .A2(n8631), .ZN(n15068) );
  INV_X1 U11254 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n8634) );
  NAND2_X1 U11255 ( .A1(n6514), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8633) );
  NAND2_X1 U11256 ( .A1(n8764), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8632) );
  OAI211_X1 U11257 ( .C1(n8768), .C2(n8634), .A(n8633), .B(n8632), .ZN(n8635)
         );
  INV_X1 U11258 ( .A(n8635), .ZN(n8636) );
  NAND2_X1 U11259 ( .A1(n12036), .A2(n8775), .ZN(n8641) );
  NAND2_X1 U11260 ( .A1(n8776), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8640) );
  MUX2_X1 U11261 ( .A(n14839), .B(n10073), .S(n8779), .Z(n8642) );
  MUX2_X1 U11262 ( .A(n14839), .B(n10073), .S(n8780), .Z(n8643) );
  NAND2_X1 U11263 ( .A1(n8644), .A2(n8643), .ZN(n8645) );
  NAND2_X1 U11264 ( .A1(n8776), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8650) );
  INV_X1 U11265 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14767) );
  NAND2_X1 U11266 ( .A1(n8651), .A2(n14767), .ZN(n8652) );
  NAND2_X1 U11267 ( .A1(n8660), .A2(n8652), .ZN(n15056) );
  INV_X1 U11268 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n12468) );
  NAND2_X1 U11269 ( .A1(n8764), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8654) );
  NAND2_X1 U11270 ( .A1(n8088), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8653) );
  OAI211_X1 U11271 ( .C1(n8688), .C2(n12468), .A(n8654), .B(n8653), .ZN(n8655)
         );
  INV_X1 U11272 ( .A(n8655), .ZN(n8656) );
  MUX2_X1 U11273 ( .A(n15053), .B(n15031), .S(n8779), .Z(n8659) );
  MUX2_X1 U11274 ( .A(n15031), .B(n15053), .S(n8779), .Z(n8658) );
  NAND2_X1 U11275 ( .A1(n8660), .A2(n14738), .ZN(n8661) );
  NAND2_X1 U11276 ( .A1(n8682), .A2(n8661), .ZN(n15033) );
  INV_X1 U11277 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n8664) );
  NAND2_X1 U11278 ( .A1(n8764), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8663) );
  NAND2_X1 U11279 ( .A1(n6514), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8662) );
  OAI211_X1 U11280 ( .C1(n8664), .C2(n8768), .A(n8663), .B(n8662), .ZN(n8665)
         );
  INV_X1 U11281 ( .A(n8665), .ZN(n8666) );
  NAND2_X1 U11282 ( .A1(n12547), .A2(n8775), .ZN(n8671) );
  NAND2_X1 U11283 ( .A1(n8776), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8670) );
  MUX2_X1 U11284 ( .A(n14838), .B(n15030), .S(n8779), .Z(n8673) );
  MUX2_X1 U11285 ( .A(n14838), .B(n15030), .S(n8261), .Z(n8672) );
  NAND2_X1 U11286 ( .A1(n8676), .A2(n8675), .ZN(n8678) );
  NAND2_X1 U11287 ( .A1(n8776), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8680) );
  NAND2_X1 U11288 ( .A1(n8682), .A2(n14817), .ZN(n8683) );
  NAND2_X1 U11289 ( .A1(n15018), .A2(n8763), .ZN(n8691) );
  INV_X1 U11290 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8687) );
  NAND2_X1 U11291 ( .A1(n8764), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8686) );
  NAND2_X1 U11292 ( .A1(n8088), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8685) );
  OAI211_X1 U11293 ( .C1(n8688), .C2(n8687), .A(n8686), .B(n8685), .ZN(n8689)
         );
  INV_X1 U11294 ( .A(n8689), .ZN(n8690) );
  MUX2_X1 U11295 ( .A(n15289), .B(n15032), .S(n8779), .Z(n8694) );
  MUX2_X1 U11296 ( .A(n15032), .B(n15289), .S(n8779), .Z(n8692) );
  INV_X1 U11297 ( .A(n8694), .ZN(n8695) );
  MUX2_X1 U11298 ( .A(n14837), .B(n15284), .S(n8780), .Z(n8696) );
  INV_X1 U11299 ( .A(n8703), .ZN(n8700) );
  INV_X1 U11300 ( .A(SI_27_), .ZN(n13609) );
  NAND2_X1 U11301 ( .A1(n8700), .A2(n13609), .ZN(n8701) );
  NAND2_X1 U11302 ( .A1(n8703), .A2(SI_27_), .ZN(n8704) );
  INV_X1 U11303 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12684) );
  INV_X1 U11304 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14667) );
  MUX2_X1 U11305 ( .A(n12684), .B(n14667), .S(n10878), .Z(n8705) );
  INV_X1 U11306 ( .A(SI_28_), .ZN(n12570) );
  NAND2_X1 U11307 ( .A1(n8705), .A2(n12570), .ZN(n8708) );
  INV_X1 U11308 ( .A(n8705), .ZN(n8706) );
  NAND2_X1 U11309 ( .A1(n8706), .A2(SI_28_), .ZN(n8707) );
  NAND2_X1 U11310 ( .A1(n8708), .A2(n8707), .ZN(n8773) );
  INV_X1 U11311 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15432) );
  INV_X1 U11312 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n12697) );
  MUX2_X1 U11313 ( .A(n15432), .B(n12697), .S(n10878), .Z(n8710) );
  XNOR2_X1 U11314 ( .A(n8710), .B(SI_29_), .ZN(n8757) );
  MUX2_X1 U11315 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n10878), .Z(n8714) );
  INV_X1 U11316 ( .A(n8714), .ZN(n8709) );
  INV_X1 U11317 ( .A(SI_30_), .ZN(n12555) );
  NAND2_X1 U11318 ( .A1(n8709), .A2(n12555), .ZN(n8736) );
  INV_X1 U11319 ( .A(SI_29_), .ZN(n12708) );
  NAND2_X1 U11320 ( .A1(n8710), .A2(n12708), .ZN(n8734) );
  NAND2_X1 U11321 ( .A1(n8736), .A2(n8734), .ZN(n8716) );
  MUX2_X1 U11322 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10878), .Z(n8712) );
  INV_X1 U11323 ( .A(SI_31_), .ZN(n8711) );
  XNOR2_X1 U11324 ( .A(n8712), .B(n8711), .ZN(n8715) );
  NOR2_X1 U11325 ( .A1(n8716), .A2(n8715), .ZN(n8713) );
  NAND2_X1 U11326 ( .A1(n8735), .A2(n8713), .ZN(n8723) );
  NAND2_X1 U11327 ( .A1(n8714), .A2(SI_30_), .ZN(n8737) );
  INV_X1 U11328 ( .A(n8715), .ZN(n8717) );
  NOR2_X1 U11329 ( .A1(n8716), .A2(n8717), .ZN(n8719) );
  XNOR2_X1 U11330 ( .A(n8717), .B(n8737), .ZN(n8718) );
  NAND2_X1 U11331 ( .A1(n14656), .A2(n8775), .ZN(n8725) );
  NAND2_X1 U11332 ( .A1(n8776), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8724) );
  NAND2_X1 U11333 ( .A1(n14974), .A2(n8261), .ZN(n8852) );
  NAND2_X1 U11334 ( .A1(n6514), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8728) );
  NAND2_X1 U11335 ( .A1(n8764), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8727) );
  NAND2_X1 U11336 ( .A1(n8088), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8726) );
  OR2_X1 U11337 ( .A1(n9877), .A2(n15163), .ZN(n10658) );
  NAND2_X1 U11338 ( .A1(n8958), .A2(n15440), .ZN(n8820) );
  OAI21_X1 U11339 ( .B1(n8971), .B2(n15440), .A(n8820), .ZN(n8729) );
  NAND2_X1 U11340 ( .A1(n10658), .A2(n8729), .ZN(n8851) );
  NAND2_X1 U11341 ( .A1(n8970), .A2(n8971), .ZN(n8853) );
  AND2_X1 U11342 ( .A1(n8851), .A2(n8853), .ZN(n8857) );
  NAND2_X1 U11343 ( .A1(n8856), .A2(n14973), .ZN(n8730) );
  OAI211_X1 U11344 ( .C1(n8852), .C2(n14973), .A(n8857), .B(n8730), .ZN(n8863)
         );
  INV_X1 U11345 ( .A(n8863), .ZN(n8749) );
  NAND2_X1 U11346 ( .A1(n6514), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8733) );
  NAND2_X1 U11347 ( .A1(n8764), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8732) );
  NAND2_X1 U11348 ( .A1(n8088), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8731) );
  AND3_X1 U11349 ( .A1(n8733), .A2(n8732), .A3(n8731), .ZN(n15008) );
  AOI21_X1 U11350 ( .B1(n14973), .B2(n8971), .A(n15008), .ZN(n8742) );
  AND2_X1 U11351 ( .A1(n8737), .A2(n8736), .ZN(n8738) );
  NAND2_X1 U11352 ( .A1(n12558), .A2(n8775), .ZN(n8741) );
  NAND2_X1 U11353 ( .A1(n8776), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8740) );
  MUX2_X1 U11354 ( .A(n8742), .B(n14977), .S(n8779), .Z(n8846) );
  INV_X1 U11355 ( .A(n14973), .ZN(n14834) );
  NAND2_X1 U11356 ( .A1(n14834), .A2(n8779), .ZN(n8746) );
  INV_X1 U11357 ( .A(n8743), .ZN(n8744) );
  NAND2_X1 U11358 ( .A1(n8744), .A2(n8970), .ZN(n8745) );
  AOI21_X1 U11359 ( .B1(n8746), .B2(n8745), .A(n15008), .ZN(n8747) );
  AOI21_X1 U11360 ( .B1(n14977), .B2(n8261), .A(n8747), .ZN(n8847) );
  OR2_X1 U11361 ( .A1(n8846), .A2(n8847), .ZN(n8748) );
  NAND2_X1 U11362 ( .A1(n8749), .A2(n8748), .ZN(n8810) );
  INV_X1 U11363 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n15004) );
  INV_X1 U11364 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8753) );
  NAND2_X1 U11365 ( .A1(n8764), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8752) );
  NAND2_X1 U11366 ( .A1(n6514), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8751) );
  OAI211_X1 U11367 ( .C1(n8753), .C2(n8768), .A(n8752), .B(n8751), .ZN(n8754)
         );
  INV_X1 U11368 ( .A(n8754), .ZN(n8755) );
  NAND2_X1 U11369 ( .A1(n12696), .A2(n8775), .ZN(n8760) );
  NAND2_X1 U11370 ( .A1(n8776), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8759) );
  MUX2_X1 U11371 ( .A(n14835), .B(n15003), .S(n8779), .Z(n8786) );
  INV_X1 U11372 ( .A(n8786), .ZN(n8761) );
  MUX2_X1 U11373 ( .A(n14835), .B(n15003), .S(n8261), .Z(n8785) );
  NAND2_X1 U11374 ( .A1(n8761), .A2(n8785), .ZN(n8807) );
  INV_X1 U11375 ( .A(n8807), .ZN(n8762) );
  XNOR2_X1 U11376 ( .A(n15005), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n12685) );
  NAND2_X1 U11377 ( .A1(n12685), .A2(n8763), .ZN(n8772) );
  INV_X1 U11378 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n8769) );
  NAND2_X1 U11379 ( .A1(n8764), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8767) );
  NAND2_X1 U11380 ( .A1(n6514), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8766) );
  OAI211_X1 U11381 ( .C1(n8769), .C2(n8768), .A(n8767), .B(n8766), .ZN(n8770)
         );
  INV_X1 U11382 ( .A(n8770), .ZN(n8771) );
  INV_X1 U11383 ( .A(n14982), .ZN(n15009) );
  NAND2_X1 U11384 ( .A1(n10297), .A2(n8775), .ZN(n8778) );
  NAND2_X1 U11385 ( .A1(n8776), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8777) );
  MUX2_X1 U11386 ( .A(n15009), .B(n14983), .S(n8779), .Z(n8782) );
  MUX2_X1 U11387 ( .A(n14982), .B(n14984), .S(n8780), .Z(n8781) );
  AND2_X1 U11388 ( .A1(n8782), .A2(n8781), .ZN(n8802) );
  NOR3_X1 U11389 ( .A1(n8789), .A2(n8790), .A3(n8802), .ZN(n8873) );
  INV_X1 U11390 ( .A(n8781), .ZN(n8784) );
  INV_X1 U11391 ( .A(n8782), .ZN(n8783) );
  NAND2_X1 U11392 ( .A1(n8784), .A2(n8783), .ZN(n8791) );
  NAND2_X1 U11393 ( .A1(n8846), .A2(n8847), .ZN(n8864) );
  INV_X1 U11394 ( .A(n8851), .ZN(n8855) );
  NAND2_X1 U11395 ( .A1(n8864), .A2(n8850), .ZN(n8808) );
  INV_X1 U11396 ( .A(n8785), .ZN(n8787) );
  NAND2_X1 U11397 ( .A1(n8787), .A2(n8786), .ZN(n8809) );
  INV_X1 U11398 ( .A(n8809), .ZN(n8788) );
  NAND3_X1 U11399 ( .A1(n8789), .A2(n8791), .A3(n8801), .ZN(n8806) );
  INV_X1 U11400 ( .A(n8790), .ZN(n8800) );
  INV_X1 U11401 ( .A(n8791), .ZN(n8799) );
  NOR2_X2 U11402 ( .A1(n8792), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n8796) );
  INV_X1 U11403 ( .A(n8796), .ZN(n8793) );
  NAND2_X1 U11404 ( .A1(n8793), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8794) );
  MUX2_X1 U11405 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8794), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n8797) );
  NAND2_X1 U11406 ( .A1(n8796), .A2(n8795), .ZN(n8812) );
  NAND2_X1 U11407 ( .A1(n8797), .A2(n8812), .ZN(n10757) );
  INV_X1 U11408 ( .A(n10757), .ZN(n8798) );
  NAND2_X1 U11409 ( .A1(n8798), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10755) );
  AOI21_X1 U11410 ( .B1(n8800), .B2(n8799), .A(n10755), .ZN(n8804) );
  INV_X1 U11411 ( .A(n10755), .ZN(n12005) );
  OAI22_X1 U11412 ( .A1(n8810), .A2(n8809), .B1(n8808), .B2(n8807), .ZN(n8870)
         );
  INV_X1 U11413 ( .A(P1_B_REG_SCAN_IN), .ZN(n8823) );
  NAND2_X1 U11414 ( .A1(n8812), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8814) );
  INV_X1 U11415 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8813) );
  XNOR2_X1 U11416 ( .A(n8814), .B(n8813), .ZN(n8980) );
  OAI21_X1 U11417 ( .B1(n8816), .B2(n8815), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8817) );
  MUX2_X1 U11418 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8817), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n8819) );
  OR2_X1 U11419 ( .A1(n8820), .A2(n8974), .ZN(n10135) );
  AND3_X1 U11420 ( .A1(n10724), .A2(n10757), .A3(n10135), .ZN(n10133) );
  NAND2_X1 U11421 ( .A1(n10133), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9000) );
  INV_X1 U11422 ( .A(n14874), .ZN(n10888) );
  NOR3_X1 U11423 ( .A1(n9000), .A2(n15433), .A3(n15225), .ZN(n8822) );
  AOI211_X1 U11424 ( .C1(n12005), .C2(n8969), .A(n8823), .B(n8822), .ZN(n8869)
         );
  XOR2_X1 U11425 ( .A(n15008), .B(n14977), .Z(n8842) );
  INV_X1 U11426 ( .A(n14835), .ZN(n8824) );
  XNOR2_X1 U11427 ( .A(n15003), .B(n8824), .ZN(n14996) );
  NAND2_X1 U11428 ( .A1(n14984), .A2(n14982), .ZN(n14995) );
  NAND2_X1 U11429 ( .A1(n15030), .A2(n14815), .ZN(n8955) );
  OR2_X1 U11430 ( .A1(n15030), .A2(n14815), .ZN(n8825) );
  XNOR2_X1 U11431 ( .A(n15090), .B(n14840), .ZN(n15076) );
  XNOR2_X1 U11432 ( .A(n15319), .B(n15117), .ZN(n15108) );
  XNOR2_X1 U11433 ( .A(n15339), .B(n15140), .ZN(n15153) );
  XNOR2_X1 U11434 ( .A(n14788), .B(n15226), .ZN(n8932) );
  XNOR2_X1 U11435 ( .A(n14724), .B(n14785), .ZN(n12189) );
  XNOR2_X1 U11436 ( .A(n15384), .B(n14729), .ZN(n8891) );
  XNOR2_X1 U11437 ( .A(n15391), .B(n12169), .ZN(n8928) );
  XNOR2_X1 U11438 ( .A(n15396), .B(n12183), .ZN(n11839) );
  NAND2_X1 U11439 ( .A1(n8926), .A2(n8826), .ZN(n11673) );
  NOR3_X1 U11440 ( .A1(n11439), .A2(n11453), .A3(n8917), .ZN(n8830) );
  INV_X1 U11441 ( .A(n11070), .ZN(n11072) );
  NAND4_X1 U11442 ( .A1(n11487), .A2(n8830), .A3(n6515), .A4(n11072), .ZN(
        n8831) );
  XNOR2_X1 U11443 ( .A(n11576), .B(n11703), .ZN(n11568) );
  NOR2_X1 U11444 ( .A1(n11839), .A2(n8832), .ZN(n8833) );
  NAND3_X1 U11445 ( .A1(n12001), .A2(n8049), .A3(n8833), .ZN(n8834) );
  OR3_X1 U11446 ( .A1(n8932), .A2(n12189), .A3(n8834), .ZN(n8835) );
  INV_X1 U11447 ( .A(n14842), .ZN(n15214) );
  XNOR2_X1 U11448 ( .A(n15350), .B(n15214), .ZN(n15172) );
  INV_X1 U11449 ( .A(n15173), .ZN(n15184) );
  NOR2_X1 U11450 ( .A1(n8836), .A2(n15184), .ZN(n8837) );
  XNOR2_X1 U11451 ( .A(n15324), .B(n15139), .ZN(n15122) );
  NOR2_X1 U11452 ( .A1(n15076), .A2(n8838), .ZN(n8839) );
  NAND4_X1 U11453 ( .A1(n15039), .A2(n8839), .A3(n15044), .A4(n15064), .ZN(
        n8840) );
  XNOR2_X1 U11454 ( .A(n8843), .B(n15199), .ZN(n8845) );
  INV_X1 U11455 ( .A(n8853), .ZN(n8844) );
  INV_X1 U11456 ( .A(n8846), .ZN(n8849) );
  INV_X1 U11457 ( .A(n8847), .ZN(n8848) );
  NAND3_X1 U11458 ( .A1(n8850), .A2(n8849), .A3(n8848), .ZN(n8862) );
  XNOR2_X1 U11459 ( .A(n8852), .B(n8851), .ZN(n8854) );
  NAND4_X1 U11460 ( .A1(n8854), .A2(n14974), .A3(n14834), .A4(n8853), .ZN(
        n8861) );
  NAND3_X1 U11461 ( .A1(n8856), .A2(n14973), .A3(n8855), .ZN(n8860) );
  INV_X1 U11462 ( .A(n8856), .ZN(n8858) );
  NAND4_X1 U11463 ( .A1(n8858), .A2(n14973), .A3(n8857), .A4(n15269), .ZN(
        n8859) );
  NAND4_X1 U11464 ( .A1(n8862), .A2(n8861), .A3(n8860), .A4(n8859), .ZN(n8866)
         );
  NOR2_X1 U11465 ( .A1(n8864), .A2(n8863), .ZN(n8865) );
  NAND2_X1 U11466 ( .A1(n14856), .A2(n11055), .ZN(n11434) );
  NAND2_X1 U11467 ( .A1(n8874), .A2(n11434), .ZN(n8876) );
  NAND2_X1 U11468 ( .A1(n8876), .A2(n8875), .ZN(n11503) );
  NAND2_X1 U11469 ( .A1(n11503), .A2(n8917), .ZN(n8878) );
  OR2_X1 U11470 ( .A1(n14855), .A2(n6516), .ZN(n8877) );
  NAND2_X1 U11471 ( .A1(n8878), .A2(n8877), .ZN(n11069) );
  NAND2_X1 U11472 ( .A1(n11069), .A2(n11070), .ZN(n8880) );
  NAND2_X1 U11473 ( .A1(n11348), .A2(n15502), .ZN(n8879) );
  NAND2_X1 U11474 ( .A1(n11393), .A2(n11489), .ZN(n8882) );
  OR2_X1 U11475 ( .A1(n11500), .A2(n14852), .ZN(n8884) );
  NAND2_X1 U11476 ( .A1(n8885), .A2(n8884), .ZN(n11567) );
  NAND2_X1 U11477 ( .A1(n11567), .A2(n11568), .ZN(n8887) );
  OR2_X1 U11478 ( .A1(n11576), .A2(n14851), .ZN(n8886) );
  NAND2_X1 U11479 ( .A1(n8887), .A2(n8886), .ZN(n11580) );
  OR2_X1 U11480 ( .A1(n11700), .A2(n14849), .ZN(n8888) );
  OR2_X1 U11481 ( .A1(n15391), .A2(n14846), .ZN(n8889) );
  OR2_X1 U11482 ( .A1(n15384), .A2(n14845), .ZN(n8892) );
  NAND2_X1 U11483 ( .A1(n15246), .A2(n8932), .ZN(n8894) );
  OR2_X1 U11484 ( .A1(n14788), .A2(n14844), .ZN(n8893) );
  NAND2_X1 U11485 ( .A1(n8894), .A2(n8893), .ZN(n15206) );
  NAND2_X1 U11486 ( .A1(n8965), .A2(n15255), .ZN(n8896) );
  AND2_X1 U11487 ( .A1(n15210), .A2(n8896), .ZN(n8895) );
  INV_X1 U11488 ( .A(n8896), .ZN(n15207) );
  NOR2_X1 U11489 ( .A1(n8897), .A2(n15207), .ZN(n8899) );
  INV_X1 U11490 ( .A(n8898), .ZN(n15218) );
  NOR2_X1 U11491 ( .A1(n15350), .A2(n14842), .ZN(n8901) );
  NAND2_X1 U11492 ( .A1(n15350), .A2(n14842), .ZN(n8902) );
  OR2_X1 U11493 ( .A1(n15342), .A2(n14841), .ZN(n8903) );
  NAND2_X1 U11494 ( .A1(n15324), .A2(n15139), .ZN(n8907) );
  NAND2_X1 U11495 ( .A1(n15090), .A2(n15099), .ZN(n8908) );
  NAND2_X1 U11496 ( .A1(n10073), .A2(n14839), .ZN(n8910) );
  NOR2_X1 U11497 ( .A1(n10073), .A2(n14839), .ZN(n8909) );
  INV_X1 U11498 ( .A(n15032), .ZN(n8956) );
  NOR2_X1 U11499 ( .A1(n15284), .A2(n14837), .ZN(n14988) );
  NOR2_X1 U11500 ( .A1(n15000), .A2(n14988), .ZN(n8911) );
  NAND2_X1 U11501 ( .A1(n8911), .A2(n8912), .ZN(n12689) );
  INV_X1 U11502 ( .A(n8911), .ZN(n8913) );
  NAND2_X1 U11503 ( .A1(n8913), .A2(n8957), .ZN(n12688) );
  NAND2_X1 U11504 ( .A1(n15440), .A2(n15163), .ZN(n8914) );
  OR2_X1 U11505 ( .A1(n9877), .A2(n8969), .ZN(n8915) );
  NAND2_X1 U11506 ( .A1(n10123), .A2(n8915), .ZN(n11384) );
  AND2_X1 U11507 ( .A1(n15199), .A2(n8969), .ZN(n8916) );
  NAND2_X1 U11508 ( .A1(n11828), .A2(n8916), .ZN(n15548) );
  NAND2_X1 U11509 ( .A1(n11493), .A2(n15548), .ZN(n15578) );
  NAND3_X1 U11510 ( .A1(n12689), .A2(n12688), .A3(n15578), .ZN(n8978) );
  NAND2_X1 U11511 ( .A1(n11073), .A2(n11072), .ZN(n11071) );
  NAND2_X1 U11512 ( .A1(n11071), .A2(n8919), .ZN(n11387) );
  NAND2_X1 U11513 ( .A1(n11387), .A2(n6515), .ZN(n11386) );
  NAND2_X1 U11514 ( .A1(n11489), .A2(n15554), .ZN(n8920) );
  OR2_X1 U11515 ( .A1(n11500), .A2(n11564), .ZN(n8921) );
  NAND2_X1 U11516 ( .A1(n11488), .A2(n8921), .ZN(n8923) );
  NAND2_X1 U11517 ( .A1(n11500), .A2(n11564), .ZN(n8922) );
  NAND2_X1 U11518 ( .A1(n8923), .A2(n8922), .ZN(n11562) );
  INV_X1 U11519 ( .A(n11568), .ZN(n11563) );
  NAND2_X1 U11520 ( .A1(n11576), .A2(n11703), .ZN(n8924) );
  OR2_X1 U11521 ( .A1(n11700), .A2(n11677), .ZN(n8925) );
  NAND2_X1 U11522 ( .A1(n11584), .A2(n8925), .ZN(n11676) );
  INV_X1 U11523 ( .A(n11673), .ZN(n11675) );
  NAND2_X1 U11524 ( .A1(n15396), .A2(n12183), .ZN(n8927) );
  OR2_X1 U11525 ( .A1(n15391), .A2(n12169), .ZN(n8929) );
  OR2_X1 U11526 ( .A1(n15384), .A2(n14729), .ZN(n8930) );
  INV_X1 U11527 ( .A(n12189), .ZN(n12191) );
  OR2_X1 U11528 ( .A1(n14724), .A2(n14785), .ZN(n8931) );
  INV_X1 U11529 ( .A(n8932), .ZN(n15248) );
  OR2_X1 U11530 ( .A1(n15350), .A2(n15214), .ZN(n8938) );
  NAND2_X1 U11531 ( .A1(n8934), .A2(n8938), .ZN(n15151) );
  INV_X1 U11532 ( .A(n15151), .ZN(n8935) );
  AND2_X1 U11533 ( .A1(n8555), .A2(n8935), .ZN(n8936) );
  NAND2_X1 U11534 ( .A1(n15350), .A2(n15214), .ZN(n15174) );
  INV_X1 U11535 ( .A(n15140), .ZN(n15177) );
  OR2_X1 U11536 ( .A1(n15339), .A2(n15177), .ZN(n8944) );
  INV_X1 U11537 ( .A(n15134), .ZN(n15132) );
  INV_X1 U11538 ( .A(n15117), .ZN(n8948) );
  NAND2_X1 U11539 ( .A1(n15319), .A2(n8948), .ZN(n8945) );
  OAI211_X1 U11540 ( .C1(n15127), .C2(n15139), .A(n15095), .B(n8945), .ZN(
        n8946) );
  OR2_X1 U11541 ( .A1(n15324), .A2(n15098), .ZN(n15096) );
  NAND2_X1 U11542 ( .A1(n15096), .A2(n8948), .ZN(n8947) );
  NAND2_X1 U11543 ( .A1(n8947), .A2(n15107), .ZN(n8950) );
  OR3_X1 U11544 ( .A1(n15324), .A2(n15098), .A3(n8948), .ZN(n8949) );
  INV_X1 U11545 ( .A(n15076), .ZN(n15083) );
  OR2_X1 U11546 ( .A1(n15090), .A2(n14840), .ZN(n8952) );
  INV_X1 U11547 ( .A(n14839), .ZN(n14766) );
  AND2_X1 U11548 ( .A1(n10073), .A2(n14766), .ZN(n8953) );
  XNOR2_X1 U11549 ( .A(n14986), .B(n8957), .ZN(n8964) );
  NAND2_X1 U11550 ( .A1(n8958), .A2(n8971), .ZN(n8960) );
  NAND2_X1 U11551 ( .A1(n15199), .A2(n15440), .ZN(n8959) );
  INV_X1 U11552 ( .A(n8965), .ZN(n8967) );
  INV_X1 U11553 ( .A(n11500), .ZN(n15563) );
  AND2_X1 U11554 ( .A1(n11497), .A2(n15563), .ZN(n11571) );
  INV_X1 U11555 ( .A(n11576), .ZN(n15570) );
  INV_X1 U11556 ( .A(n15391), .ZN(n11922) );
  NAND2_X1 U11557 ( .A1(n11920), .A2(n11922), .ZN(n11996) );
  INV_X1 U11558 ( .A(n14788), .ZN(n15372) );
  NOR2_X2 U11559 ( .A1(n15235), .A2(n8898), .ZN(n15193) );
  INV_X1 U11560 ( .A(n15339), .ZN(n15159) );
  NOR2_X2 U11561 ( .A1(n15137), .A2(n15324), .ZN(n15113) );
  NOR2_X2 U11562 ( .A1(n15055), .A2(n15030), .ZN(n15029) );
  INV_X1 U11563 ( .A(n10665), .ZN(n8972) );
  NAND2_X1 U11564 ( .A1(n8970), .A2(n8969), .ZN(n10139) );
  AOI21_X1 U11565 ( .B1(n14984), .B2(n8972), .A(n15571), .ZN(n8973) );
  INV_X1 U11566 ( .A(n10139), .ZN(n11019) );
  INV_X1 U11567 ( .A(n8974), .ZN(n8975) );
  NAND2_X1 U11568 ( .A1(n12565), .A2(P1_B_REG_SCAN_IN), .ZN(n8981) );
  MUX2_X1 U11569 ( .A(P1_B_REG_SCAN_IN), .B(n8981), .S(n8980), .Z(n8982) );
  OR2_X1 U11570 ( .A1(n10867), .A2(P1_D_REG_1__SCAN_IN), .ZN(n8984) );
  INV_X1 U11571 ( .A(n10868), .ZN(n15439) );
  NAND2_X1 U11572 ( .A1(n12565), .A2(n15439), .ZN(n8983) );
  NAND2_X1 U11573 ( .A1(n8984), .A2(n8983), .ZN(n10118) );
  NOR2_X1 U11574 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .ZN(
        n12502) );
  NOR4_X1 U11575 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n8987) );
  NOR4_X1 U11576 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n8986) );
  NOR4_X1 U11577 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n8985) );
  AND4_X1 U11578 ( .A1(n12502), .A2(n8987), .A3(n8986), .A4(n8985), .ZN(n8993)
         );
  NOR4_X1 U11579 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n8991) );
  NOR4_X1 U11580 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n8990) );
  NOR4_X1 U11581 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n8989) );
  NOR4_X1 U11582 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n8988) );
  AND4_X1 U11583 ( .A1(n8991), .A2(n8990), .A3(n8989), .A4(n8988), .ZN(n8992)
         );
  AND2_X1 U11584 ( .A1(n8993), .A2(n8992), .ZN(n8994) );
  NAND2_X1 U11585 ( .A1(n8980), .A2(n15439), .ZN(n10875) );
  NOR2_X1 U11586 ( .A1(n10654), .A2(n9000), .ZN(n8996) );
  NAND2_X1 U11587 ( .A1(n9003), .A2(n15599), .ZN(n8999) );
  INV_X1 U11588 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n8997) );
  NAND2_X1 U11589 ( .A1(n8999), .A2(n8998), .ZN(P1_U3556) );
  INV_X1 U11590 ( .A(n9000), .ZN(n10656) );
  NAND2_X1 U11591 ( .A1(n9003), .A2(n15588), .ZN(n9005) );
  OR2_X1 U11592 ( .A1(n15588), .A2(n8769), .ZN(n9004) );
  NAND2_X1 U11593 ( .A1(n9005), .A2(n9004), .ZN(P1_U3524) );
  NOR2_X1 U11594 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_20__SCAN_IN), 
        .ZN(n9008) );
  NAND4_X1 U11595 ( .A1(n9008), .A2(n9007), .A3(n9006), .A4(n9335), .ZN(n9492)
         );
  NAND4_X1 U11596 ( .A1(n9575), .A2(n7971), .A3(n9541), .A4(n9544), .ZN(n9009)
         );
  NOR2_X2 U11597 ( .A1(n9492), .A2(n9009), .ZN(n9547) );
  INV_X1 U11598 ( .A(n9021), .ZN(n12557) );
  INV_X1 U11599 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n9015) );
  NAND2_X1 U11600 ( .A1(n9176), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9025) );
  NAND2_X1 U11601 ( .A1(n12557), .A2(n9020), .ZN(n9041) );
  INV_X1 U11602 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n11325) );
  OR2_X1 U11603 ( .A1(n9041), .A2(n11325), .ZN(n9023) );
  INV_X1 U11604 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n11404) );
  OR2_X1 U11605 ( .A1(n9058), .A2(n11404), .ZN(n9022) );
  XNOR2_X2 U11606 ( .A(n9027), .B(n9026), .ZN(n9503) );
  NAND2_X1 U11607 ( .A1(n9028), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9029) );
  AND2_X1 U11608 ( .A1(n9048), .A2(n9029), .ZN(n10837) );
  NAND2_X1 U11609 ( .A1(n9101), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9030) );
  INV_X1 U11610 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n12452) );
  OR2_X1 U11611 ( .A1(n9089), .A2(n12452), .ZN(n9034) );
  INV_X1 U11612 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11099) );
  OR2_X1 U11613 ( .A1(n9058), .A2(n11099), .ZN(n9032) );
  NAND2_X1 U11614 ( .A1(n6518), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n9031) );
  XNOR2_X1 U11615 ( .A(n9049), .B(n9048), .ZN(n10849) );
  NAND2_X1 U11616 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n9035) );
  NAND2_X1 U11617 ( .A1(n9101), .A2(n10848), .ZN(n9036) );
  INV_X1 U11618 ( .A(n13042), .ZN(n9037) );
  INV_X1 U11619 ( .A(n13042), .ZN(n15860) );
  NAND2_X1 U11620 ( .A1(n15860), .A2(n11661), .ZN(n9038) );
  INV_X1 U11621 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n9040) );
  OR2_X1 U11622 ( .A1(n9089), .A2(n9040), .ZN(n9044) );
  NAND2_X1 U11623 ( .A1(n6518), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9043) );
  INV_X1 U11624 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9619) );
  OR2_X1 U11625 ( .A1(n9041), .A2(n9619), .ZN(n9042) );
  INV_X1 U11626 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15856) );
  OR2_X1 U11627 ( .A1(n9058), .A2(n15856), .ZN(n9045) );
  NAND2_X1 U11628 ( .A1(n10847), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9050) );
  XNOR2_X1 U11629 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n9052) );
  XNOR2_X1 U11630 ( .A(n9066), .B(n9052), .ZN(n10853) );
  OR2_X1 U11631 ( .A1(n9064), .A2(n10853), .ZN(n9054) );
  OR2_X1 U11632 ( .A1(n9069), .A2(SI_2_), .ZN(n9053) );
  INV_X1 U11633 ( .A(n15852), .ZN(n11283) );
  NOR2_X1 U11634 ( .A1(n9055), .A2(n11283), .ZN(n9056) );
  NAND2_X1 U11635 ( .A1(n9466), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9062) );
  OR2_X1 U11636 ( .A1(n9346), .A2(n15910), .ZN(n9061) );
  INV_X1 U11637 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n9057) );
  OR2_X1 U11638 ( .A1(n9089), .A2(n9057), .ZN(n9060) );
  OR2_X1 U11639 ( .A1(n9058), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n9059) );
  NAND2_X1 U11640 ( .A1(n12482), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n9065) );
  NAND2_X1 U11641 ( .A1(n10840), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9067) );
  XNOR2_X1 U11642 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n9068) );
  XNOR2_X1 U11643 ( .A(n9084), .B(n9068), .ZN(n10832) );
  OR2_X1 U11644 ( .A1(n9064), .A2(n10832), .ZN(n9071) );
  OR2_X1 U11645 ( .A1(n9069), .A2(SI_3_), .ZN(n9070) );
  OAI211_X1 U11646 ( .C1(n9605), .C2(n11124), .A(n9071), .B(n9070), .ZN(n15881) );
  NAND2_X1 U11647 ( .A1(n13041), .A2(n15881), .ZN(n12910) );
  NAND2_X1 U11648 ( .A1(n13041), .A2(n7250), .ZN(n9072) );
  NAND2_X1 U11649 ( .A1(n9466), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9081) );
  INV_X1 U11650 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n9073) );
  OR2_X1 U11651 ( .A1(n9346), .A2(n9073), .ZN(n9080) );
  NAND2_X1 U11652 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n9076) );
  AND2_X1 U11653 ( .A1(n9087), .A2(n9076), .ZN(n11632) );
  OR2_X1 U11654 ( .A1(n9058), .A2(n11632), .ZN(n9079) );
  INV_X1 U11655 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n9077) );
  OR2_X1 U11656 ( .A1(n9089), .A2(n9077), .ZN(n9078) );
  NAND2_X1 U11657 ( .A1(n12296), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n9082) );
  XNOR2_X1 U11658 ( .A(n9097), .B(n9095), .ZN(n10830) );
  INV_X1 U11659 ( .A(n15885), .ZN(n11531) );
  NAND2_X1 U11660 ( .A1(n13040), .A2(n11531), .ZN(n9085) );
  NAND2_X1 U11661 ( .A1(n9466), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n9094) );
  INV_X1 U11662 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15913) );
  OR2_X1 U11663 ( .A1(n9346), .A2(n15913), .ZN(n9093) );
  NAND2_X1 U11664 ( .A1(n9087), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n9088) );
  AND2_X1 U11665 ( .A1(n9109), .A2(n9088), .ZN(n11617) );
  OR2_X1 U11666 ( .A1(n9058), .A2(n11617), .ZN(n9092) );
  INV_X1 U11667 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n9090) );
  OR2_X1 U11668 ( .A1(n12847), .A2(n9090), .ZN(n9091) );
  NAND4_X1 U11669 ( .A1(n9094), .A2(n9093), .A3(n9092), .A4(n9091), .ZN(n13039) );
  INV_X1 U11670 ( .A(n9095), .ZN(n9096) );
  NAND2_X1 U11671 ( .A1(n9098), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n9099) );
  XNOR2_X1 U11672 ( .A(n9118), .B(P1_DATAO_REG_5__SCAN_IN), .ZN(n9115) );
  XNOR2_X1 U11673 ( .A(n9117), .B(n9115), .ZN(n10844) );
  OR2_X1 U11674 ( .A1(n9064), .A2(n10844), .ZN(n9106) );
  OR2_X1 U11675 ( .A1(n7381), .A2(SI_5_), .ZN(n9105) );
  NOR2_X1 U11676 ( .A1(n9102), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n9122) );
  OR2_X1 U11677 ( .A1(n9122), .A2(n9015), .ZN(n9103) );
  NAND2_X1 U11678 ( .A1(n9356), .A2(n11202), .ZN(n9104) );
  XNOR2_X1 U11679 ( .A(n13039), .B(n11614), .ZN(n12916) );
  INV_X1 U11680 ( .A(n11614), .ZN(n15892) );
  NAND2_X1 U11681 ( .A1(n11772), .A2(n15892), .ZN(n9108) );
  NAND2_X1 U11682 ( .A1(n9466), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9114) );
  OR2_X1 U11683 ( .A1(n9346), .A2(n15915), .ZN(n9113) );
  NAND2_X1 U11684 ( .A1(n9109), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9110) );
  AND2_X1 U11685 ( .A1(n9128), .A2(n9110), .ZN(n11777) );
  INV_X1 U11686 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n9111) );
  INV_X1 U11687 ( .A(n9115), .ZN(n9116) );
  NAND2_X1 U11688 ( .A1(n9118), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n9119) );
  NAND2_X1 U11689 ( .A1(n10886), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n9120) );
  XNOR2_X1 U11690 ( .A(n9138), .B(n9135), .ZN(n10858) );
  OR2_X1 U11691 ( .A1(n9064), .A2(n10858), .ZN(n9126) );
  INV_X1 U11692 ( .A(SI_6_), .ZN(n10857) );
  OR2_X1 U11693 ( .A1(n7381), .A2(n10857), .ZN(n9125) );
  NAND2_X1 U11694 ( .A1(n9122), .A2(n9121), .ZN(n9220) );
  NAND2_X1 U11695 ( .A1(n9220), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9123) );
  XNOR2_X1 U11696 ( .A(n9123), .B(P3_IR_REG_6__SCAN_IN), .ZN(n9644) );
  NAND2_X1 U11697 ( .A1(n9356), .A2(n9644), .ZN(n9124) );
  INV_X1 U11698 ( .A(n12922), .ZN(n12919) );
  INV_X1 U11699 ( .A(n15896), .ZN(n11774) );
  NAND2_X1 U11700 ( .A1(n13038), .A2(n11774), .ZN(n11845) );
  NAND2_X1 U11701 ( .A1(n11688), .A2(n11845), .ZN(n9145) );
  NAND2_X1 U11702 ( .A1(n9466), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n9134) );
  INV_X1 U11703 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n9648) );
  OR2_X1 U11704 ( .A1(n9346), .A2(n9648), .ZN(n9133) );
  NAND2_X1 U11705 ( .A1(n9128), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9129) );
  AND2_X1 U11706 ( .A1(n9147), .A2(n9129), .ZN(n11844) );
  OR2_X1 U11707 ( .A1(n9058), .A2(n11844), .ZN(n9132) );
  INV_X1 U11708 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n9130) );
  OR2_X1 U11709 ( .A1(n12847), .A2(n9130), .ZN(n9131) );
  INV_X1 U11710 ( .A(n9135), .ZN(n9137) );
  XNOR2_X1 U11711 ( .A(n9155), .B(n9154), .ZN(n10852) );
  NAND2_X1 U11712 ( .A1(n10852), .A2(n7262), .ZN(n9144) );
  OR2_X1 U11713 ( .A1(n7381), .A2(SI_7_), .ZN(n9143) );
  NAND2_X1 U11714 ( .A1(n9157), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9141) );
  INV_X1 U11715 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n9140) );
  XNOR2_X1 U11716 ( .A(n9141), .B(n9140), .ZN(n11297) );
  NAND2_X1 U11717 ( .A1(n9356), .A2(n11297), .ZN(n9142) );
  NAND2_X1 U11718 ( .A1(n13037), .A2(n11815), .ZN(n9146) );
  NAND2_X1 U11719 ( .A1(n9466), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n9153) );
  INV_X1 U11720 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n9656) );
  OR2_X1 U11721 ( .A1(n9346), .A2(n9656), .ZN(n9152) );
  NAND2_X1 U11722 ( .A1(n9147), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n9148) );
  AND2_X1 U11723 ( .A1(n9178), .A2(n9148), .ZN(n12096) );
  OR2_X1 U11724 ( .A1(n9058), .A2(n12096), .ZN(n9151) );
  INV_X1 U11725 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n9149) );
  OR2_X1 U11726 ( .A1(n12847), .A2(n9149), .ZN(n9150) );
  XNOR2_X1 U11727 ( .A(n10912), .B(P2_DATAO_REG_8__SCAN_IN), .ZN(n9156) );
  XNOR2_X1 U11728 ( .A(n9164), .B(n9156), .ZN(n10841) );
  NAND2_X1 U11729 ( .A1(n10841), .A2(n7262), .ZN(n9160) );
  NAND2_X1 U11730 ( .A1(n9166), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9158) );
  XNOR2_X1 U11731 ( .A(n9158), .B(P3_IR_REG_8__SCAN_IN), .ZN(n9657) );
  AOI22_X1 U11732 ( .A1(n12863), .A2(SI_8_), .B1(n9356), .B2(n9657), .ZN(n9159) );
  NAND2_X1 U11733 ( .A1(n9160), .A2(n9159), .ZN(n13498) );
  NAND2_X1 U11734 ( .A1(n11944), .A2(n13498), .ZN(n12932) );
  INV_X1 U11735 ( .A(n13498), .ZN(n9794) );
  NAND2_X1 U11736 ( .A1(n9794), .A2(n13036), .ZN(n12933) );
  NAND2_X1 U11737 ( .A1(n9794), .A2(n11944), .ZN(n9161) );
  NAND2_X1 U11738 ( .A1(n10912), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n9162) );
  XNOR2_X1 U11739 ( .A(n12483), .B(P1_DATAO_REG_9__SCAN_IN), .ZN(n9165) );
  XNOR2_X1 U11740 ( .A(n9186), .B(n9165), .ZN(n10861) );
  NAND2_X1 U11741 ( .A1(n10861), .A2(n7262), .ZN(n9175) );
  INV_X1 U11742 ( .A(n9166), .ZN(n9168) );
  INV_X1 U11743 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n9167) );
  NAND2_X1 U11744 ( .A1(n9168), .A2(n9167), .ZN(n9170) );
  NAND2_X1 U11745 ( .A1(n9170), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9169) );
  MUX2_X1 U11746 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9169), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n9173) );
  INV_X1 U11747 ( .A(n9170), .ZN(n9172) );
  INV_X1 U11748 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9171) );
  NAND2_X1 U11749 ( .A1(n9172), .A2(n9171), .ZN(n9205) );
  NAND2_X1 U11750 ( .A1(n9173), .A2(n9205), .ZN(n11740) );
  INV_X1 U11751 ( .A(SI_9_), .ZN(n10860) );
  AOI22_X1 U11752 ( .A1(n9356), .A2(n11740), .B1(n12863), .B2(n10860), .ZN(
        n9174) );
  NAND2_X1 U11753 ( .A1(n9175), .A2(n9174), .ZN(n11950) );
  NAND2_X1 U11754 ( .A1(n9176), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9183) );
  INV_X1 U11755 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n12462) );
  OR2_X1 U11756 ( .A1(n9346), .A2(n12462), .ZN(n9182) );
  NAND2_X1 U11757 ( .A1(n9178), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n9179) );
  AND2_X1 U11758 ( .A1(n9194), .A2(n9179), .ZN(n11949) );
  OR2_X1 U11759 ( .A1(n9058), .A2(n11949), .ZN(n9181) );
  INV_X1 U11760 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11948) );
  OR2_X1 U11761 ( .A1(n12858), .A2(n11948), .ZN(n9180) );
  NAND4_X1 U11762 ( .A1(n9183), .A2(n9182), .A3(n9181), .A4(n9180), .ZN(n13035) );
  AND2_X1 U11763 ( .A1(n11950), .A2(n12148), .ZN(n9185) );
  NAND2_X1 U11764 ( .A1(n10945), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n9187) );
  NAND2_X1 U11765 ( .A1(n12483), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9189) );
  XNOR2_X1 U11766 ( .A(n9202), .B(n9201), .ZN(n10874) );
  NAND2_X1 U11767 ( .A1(n10874), .A2(n7262), .ZN(n9193) );
  NAND2_X1 U11768 ( .A1(n9205), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9191) );
  INV_X1 U11769 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9190) );
  INV_X1 U11770 ( .A(SI_10_), .ZN(n10873) );
  AOI22_X1 U11771 ( .A1(n10872), .A2(n9356), .B1(n12863), .B2(n10873), .ZN(
        n9192) );
  NAND2_X1 U11772 ( .A1(n12855), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9199) );
  INV_X1 U11773 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n13596) );
  OR2_X1 U11774 ( .A1(n12847), .A2(n13596), .ZN(n9198) );
  NAND2_X1 U11775 ( .A1(n9194), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9195) );
  AND2_X1 U11776 ( .A1(n9210), .A2(n9195), .ZN(n12153) );
  OR2_X1 U11777 ( .A1(n9058), .A2(n12153), .ZN(n9197) );
  INV_X1 U11778 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n12154) );
  OR2_X1 U11779 ( .A1(n12858), .A2(n12154), .ZN(n9196) );
  NAND4_X1 U11780 ( .A1(n9199), .A2(n9198), .A3(n9197), .A4(n9196), .ZN(n13423) );
  NAND2_X1 U11781 ( .A1(n13598), .A2(n13423), .ZN(n12942) );
  NAND2_X1 U11782 ( .A1(n12943), .A2(n12942), .ZN(n12941) );
  INV_X1 U11783 ( .A(n13423), .ZN(n12207) );
  OR2_X1 U11784 ( .A1(n13598), .A2(n12207), .ZN(n9200) );
  NAND2_X1 U11785 ( .A1(n10967), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n9216) );
  NAND2_X1 U11786 ( .A1(n12309), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n9204) );
  XNOR2_X1 U11787 ( .A(n9217), .B(n6694), .ZN(n10902) );
  NAND2_X1 U11788 ( .A1(n10902), .A2(n7262), .ZN(n9209) );
  OAI21_X1 U11789 ( .B1(n9205), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9207) );
  INV_X1 U11790 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n9206) );
  XNOR2_X1 U11791 ( .A(n9207), .B(n9206), .ZN(n10903) );
  AOI22_X1 U11792 ( .A1(n10903), .A2(n9356), .B1(n12863), .B2(n10901), .ZN(
        n9208) );
  NAND2_X1 U11793 ( .A1(n9209), .A2(n9208), .ZN(n12205) );
  NAND2_X1 U11794 ( .A1(n9466), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n9215) );
  INV_X1 U11795 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n13487) );
  OR2_X1 U11796 ( .A1(n9346), .A2(n13487), .ZN(n9214) );
  INV_X1 U11797 ( .A(n6591), .ZN(n9226) );
  NAND2_X1 U11798 ( .A1(n9210), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9211) );
  AND2_X1 U11799 ( .A1(n9226), .A2(n9211), .ZN(n13425) );
  OR2_X1 U11800 ( .A1(n9058), .A2(n13425), .ZN(n9213) );
  INV_X1 U11801 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n13589) );
  OR2_X1 U11802 ( .A1(n12847), .A2(n13589), .ZN(n9212) );
  XNOR2_X1 U11803 ( .A(n11023), .B(P2_DATAO_REG_12__SCAN_IN), .ZN(n9234) );
  XNOR2_X1 U11804 ( .A(n9235), .B(n9234), .ZN(n10916) );
  NAND2_X1 U11805 ( .A1(n10916), .A2(n7262), .ZN(n9224) );
  INV_X1 U11806 ( .A(n9218), .ZN(n9219) );
  OAI21_X1 U11807 ( .B1(n9220), .B2(n9219), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n9222) );
  INV_X1 U11808 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n9221) );
  XNOR2_X1 U11809 ( .A(n9222), .B(n9221), .ZN(n10917) );
  AOI22_X1 U11810 ( .A1(n12863), .A2(n10915), .B1(n9356), .B2(n10917), .ZN(
        n9223) );
  NAND2_X1 U11811 ( .A1(n9466), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n9231) );
  INV_X1 U11812 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n13485) );
  OR2_X1 U11813 ( .A1(n9346), .A2(n13485), .ZN(n9230) );
  NAND2_X1 U11814 ( .A1(n9226), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9227) );
  AND2_X1 U11815 ( .A1(n9264), .A2(n9227), .ZN(n13409) );
  OR2_X1 U11816 ( .A1(n9058), .A2(n13409), .ZN(n9229) );
  INV_X1 U11817 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n13585) );
  OR2_X1 U11818 ( .A1(n12847), .A2(n13585), .ZN(n9228) );
  NAND4_X1 U11819 ( .A1(n9231), .A2(n9230), .A3(n9229), .A4(n9228), .ZN(n13421) );
  NAND2_X1 U11820 ( .A1(n12954), .A2(n12531), .ZN(n9233) );
  NOR2_X1 U11821 ( .A1(n12954), .A2(n12531), .ZN(n9232) );
  NAND2_X1 U11822 ( .A1(n9236), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n9237) );
  XNOR2_X1 U11823 ( .A(n9277), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n9257) );
  NAND2_X1 U11824 ( .A1(n9257), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n9240) );
  NAND2_X1 U11825 ( .A1(n9277), .A2(n11047), .ZN(n9239) );
  NAND2_X1 U11826 ( .A1(n9240), .A2(n9239), .ZN(n9242) );
  NAND2_X1 U11827 ( .A1(n11320), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9272) );
  NAND2_X1 U11828 ( .A1(n11323), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n9273) );
  NAND2_X1 U11829 ( .A1(n9272), .A2(n9273), .ZN(n9241) );
  XNOR2_X1 U11830 ( .A(n9242), .B(n9241), .ZN(n11043) );
  NAND2_X1 U11831 ( .A1(n11043), .A2(n7262), .ZN(n9249) );
  NOR2_X1 U11832 ( .A1(n9260), .A2(n9015), .ZN(n9243) );
  MUX2_X1 U11833 ( .A(n9015), .B(n9243), .S(P3_IR_REG_14__SCAN_IN), .Z(n9246)
         );
  INV_X1 U11834 ( .A(n9493), .ZN(n9245) );
  INV_X1 U11835 ( .A(n13095), .ZN(n9247) );
  AOI22_X1 U11836 ( .A1(n12863), .A2(SI_14_), .B1(n9356), .B2(n9247), .ZN(
        n9248) );
  NAND2_X1 U11837 ( .A1(n9266), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9252) );
  NAND2_X1 U11838 ( .A1(n6543), .A2(n9252), .ZN(n13385) );
  NAND2_X1 U11839 ( .A1(n9497), .A2(n13385), .ZN(n9256) );
  NAND2_X1 U11840 ( .A1(n12855), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9255) );
  INV_X1 U11841 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13573) );
  OR2_X1 U11842 ( .A1(n12847), .A2(n13573), .ZN(n9254) );
  INV_X1 U11843 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13384) );
  OR2_X1 U11844 ( .A1(n12858), .A2(n13384), .ZN(n9253) );
  NAND4_X1 U11845 ( .A1(n9256), .A2(n9255), .A3(n9254), .A4(n9253), .ZN(n13392) );
  NAND2_X1 U11846 ( .A1(n13574), .A2(n12837), .ZN(n12958) );
  XNOR2_X1 U11847 ( .A(n9257), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n11000) );
  NAND2_X1 U11848 ( .A1(n11000), .A2(n7262), .ZN(n9263) );
  NOR2_X1 U11849 ( .A1(n9258), .A2(n9015), .ZN(n9259) );
  MUX2_X1 U11850 ( .A(n9015), .B(n9259), .S(P3_IR_REG_13__SCAN_IN), .Z(n9261)
         );
  OR2_X1 U11851 ( .A1(n9261), .A2(n9260), .ZN(n10998) );
  AOI22_X1 U11852 ( .A1(n12863), .A2(n10999), .B1(n9356), .B2(n10998), .ZN(
        n9262) );
  NAND2_X1 U11853 ( .A1(n9466), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n9270) );
  INV_X1 U11854 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n13480) );
  OR2_X1 U11855 ( .A1(n9346), .A2(n13480), .ZN(n9269) );
  NAND2_X1 U11856 ( .A1(n9264), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9265) );
  AND2_X1 U11857 ( .A1(n9266), .A2(n9265), .ZN(n12242) );
  OR2_X1 U11858 ( .A1(n9058), .A2(n12242), .ZN(n9268) );
  INV_X1 U11859 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n13579) );
  OR2_X1 U11860 ( .A1(n12847), .A2(n13579), .ZN(n9267) );
  NAND2_X1 U11861 ( .A1(n12896), .A2(n13403), .ZN(n13367) );
  INV_X1 U11862 ( .A(n13367), .ZN(n12957) );
  OR2_X1 U11863 ( .A1(n12896), .A2(n13403), .ZN(n12875) );
  NAND2_X1 U11864 ( .A1(n11047), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n9271) );
  NAND2_X1 U11865 ( .A1(n9272), .A2(n9271), .ZN(n9276) );
  NAND3_X1 U11866 ( .A1(n9272), .A2(P2_DATAO_REG_13__SCAN_IN), .A3(n11051), 
        .ZN(n9274) );
  XNOR2_X1 U11867 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n9290) );
  XNOR2_X1 U11868 ( .A(n9291), .B(n9290), .ZN(n11013) );
  NAND2_X1 U11869 ( .A1(n11013), .A2(n7262), .ZN(n9280) );
  NAND2_X1 U11870 ( .A1(n9493), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9278) );
  XNOR2_X1 U11871 ( .A(n9278), .B(P3_IR_REG_15__SCAN_IN), .ZN(n13111) );
  AOI22_X1 U11872 ( .A1(n12863), .A2(SI_15_), .B1(n9356), .B2(n13111), .ZN(
        n9279) );
  INV_X1 U11873 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13567) );
  AOI22_X1 U11874 ( .A1(n9466), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n12855), 
        .B2(P3_REG1_REG_15__SCAN_IN), .ZN(n9284) );
  NAND2_X1 U11875 ( .A1(n6543), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9282) );
  NAND2_X1 U11876 ( .A1(n9294), .A2(n9282), .ZN(n13375) );
  NAND2_X1 U11877 ( .A1(n13375), .A2(n9497), .ZN(n9283) );
  NAND2_X1 U11878 ( .A1(n13568), .A2(n13382), .ZN(n9285) );
  NAND2_X1 U11879 ( .A1(n13574), .A2(n13392), .ZN(n13368) );
  OAI211_X1 U11880 ( .C1(n13369), .C2(n12875), .A(n9285), .B(n13368), .ZN(
        n9286) );
  INV_X1 U11881 ( .A(n9286), .ZN(n9287) );
  NAND2_X1 U11882 ( .A1(n11377), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9292) );
  XNOR2_X1 U11883 ( .A(n11217), .B(P2_DATAO_REG_16__SCAN_IN), .ZN(n9298) );
  XNOR2_X1 U11884 ( .A(n9300), .B(n9298), .ZN(n11052) );
  NAND2_X1 U11885 ( .A1(n6648), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9304) );
  XNOR2_X1 U11886 ( .A(n9304), .B(n9335), .ZN(n13123) );
  OAI22_X1 U11887 ( .A1(n7381), .A2(n11053), .B1(n13123), .B2(n9605), .ZN(
        n9293) );
  INV_X1 U11888 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13561) );
  NAND2_X1 U11889 ( .A1(n9294), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9295) );
  NAND2_X1 U11890 ( .A1(n9323), .A2(n9295), .ZN(n13361) );
  NAND2_X1 U11891 ( .A1(n13361), .A2(n9497), .ZN(n9297) );
  AOI22_X1 U11892 ( .A1(n9466), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n12855), 
        .B2(P3_REG1_REG_16__SCAN_IN), .ZN(n9296) );
  INV_X1 U11893 ( .A(n13373), .ZN(n12774) );
  INV_X1 U11894 ( .A(n9298), .ZN(n9299) );
  NAND2_X1 U11895 ( .A1(n11214), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9301) );
  XNOR2_X1 U11896 ( .A(n7796), .B(P2_DATAO_REG_17__SCAN_IN), .ZN(n9303) );
  XNOR2_X1 U11897 ( .A(n9316), .B(n9303), .ZN(n11065) );
  NAND2_X1 U11898 ( .A1(n11065), .A2(n7262), .ZN(n9308) );
  NAND2_X1 U11899 ( .A1(n9304), .A2(n9335), .ZN(n9305) );
  NAND2_X1 U11900 ( .A1(n9305), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9306) );
  XNOR2_X1 U11901 ( .A(n9306), .B(P3_IR_REG_17__SCAN_IN), .ZN(n13151) );
  AOI22_X1 U11902 ( .A1(n9356), .A2(n13151), .B1(n12863), .B2(SI_17_), .ZN(
        n9307) );
  XNOR2_X1 U11903 ( .A(n9323), .B(P3_REG3_REG_17__SCAN_IN), .ZN(n13352) );
  NAND2_X1 U11904 ( .A1(n13352), .A2(n9497), .ZN(n9313) );
  INV_X1 U11905 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13351) );
  NAND2_X1 U11906 ( .A1(n12855), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9310) );
  NAND2_X1 U11907 ( .A1(n9176), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n9309) );
  OAI211_X1 U11908 ( .C1(n13351), .C2(n12858), .A(n9310), .B(n9309), .ZN(n9311) );
  INV_X1 U11909 ( .A(n9311), .ZN(n9312) );
  XNOR2_X1 U11910 ( .A(n13556), .B(n13358), .ZN(n13348) );
  INV_X1 U11911 ( .A(n13556), .ZN(n12778) );
  NAND2_X1 U11912 ( .A1(n11657), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n9318) );
  INV_X1 U11913 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11656) );
  NAND2_X1 U11914 ( .A1(n11656), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n9317) );
  NAND2_X1 U11915 ( .A1(n9318), .A2(n9317), .ZN(n9350) );
  NAND2_X1 U11916 ( .A1(n11780), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n9320) );
  INV_X1 U11917 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11782) );
  NAND2_X1 U11918 ( .A1(n11782), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n9319) );
  XNOR2_X1 U11919 ( .A(n9369), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n11696) );
  NAND2_X1 U11920 ( .A1(n11696), .A2(n7262), .ZN(n9322) );
  NAND2_X1 U11921 ( .A1(n12863), .A2(SI_20_), .ZN(n9321) );
  INV_X1 U11922 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n9324) );
  NAND2_X1 U11923 ( .A1(n9343), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9325) );
  NAND2_X1 U11924 ( .A1(n9378), .A2(n9325), .ZN(n13311) );
  NAND2_X1 U11925 ( .A1(n13311), .A2(n9497), .ZN(n9330) );
  INV_X1 U11926 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13460) );
  NAND2_X1 U11927 ( .A1(n9466), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n9327) );
  NAND2_X1 U11928 ( .A1(n9176), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n9326) );
  OAI211_X1 U11929 ( .C1(n9346), .C2(n13460), .A(n9327), .B(n9326), .ZN(n9328)
         );
  INV_X1 U11930 ( .A(n9328), .ZN(n9329) );
  NAND2_X1 U11931 ( .A1(n13538), .A2(n13323), .ZN(n12984) );
  OR2_X1 U11932 ( .A1(n9332), .A2(n9331), .ZN(n9333) );
  NAND2_X1 U11933 ( .A1(n9334), .A2(n9333), .ZN(n11362) );
  NAND2_X1 U11934 ( .A1(n11362), .A2(n7262), .ZN(n9340) );
  INV_X1 U11935 ( .A(n9487), .ZN(n9337) );
  NAND2_X1 U11936 ( .A1(n9337), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9338) );
  INV_X1 U11937 ( .A(SI_19_), .ZN(n11363) );
  AOI22_X1 U11938 ( .A1(n13170), .A2(n9356), .B1(n12863), .B2(n11363), .ZN(
        n9339) );
  NAND2_X1 U11939 ( .A1(n9362), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9342) );
  NAND2_X1 U11940 ( .A1(n13327), .A2(n9497), .ZN(n9349) );
  INV_X1 U11941 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13463) );
  NAND2_X1 U11942 ( .A1(n9176), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9345) );
  NAND2_X1 U11943 ( .A1(n9466), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n9344) );
  OAI211_X1 U11944 ( .C1(n9346), .C2(n13463), .A(n9345), .B(n9344), .ZN(n9347)
         );
  INV_X1 U11945 ( .A(n9347), .ZN(n9348) );
  NAND2_X1 U11946 ( .A1(n12735), .A2(n13336), .ZN(n13299) );
  NAND2_X1 U11947 ( .A1(n9351), .A2(n9350), .ZN(n9352) );
  NAND2_X1 U11948 ( .A1(n9353), .A2(n9352), .ZN(n11128) );
  OR2_X1 U11949 ( .A1(n11128), .A2(n9064), .ZN(n9358) );
  NAND2_X1 U11950 ( .A1(n9354), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9355) );
  XNOR2_X1 U11951 ( .A(n9355), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13160) );
  AOI22_X1 U11952 ( .A1(SI_18_), .A2(n12863), .B1(n13160), .B2(n9356), .ZN(
        n9357) );
  INV_X1 U11953 ( .A(n9359), .ZN(n9360) );
  NAND2_X1 U11954 ( .A1(n9360), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9361) );
  NAND2_X1 U11955 ( .A1(n9362), .A2(n9361), .ZN(n13339) );
  NAND2_X1 U11956 ( .A1(n13339), .A2(n9497), .ZN(n9367) );
  INV_X1 U11957 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13549) );
  NAND2_X1 U11958 ( .A1(n12855), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9364) );
  NAND2_X1 U11959 ( .A1(n9466), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9363) );
  OAI211_X1 U11960 ( .C1(n13549), .C2(n12847), .A(n9364), .B(n9363), .ZN(n9365) );
  INV_X1 U11961 ( .A(n9365), .ZN(n9366) );
  AND2_X1 U11962 ( .A1(n12811), .A2(n13322), .ZN(n13319) );
  OR2_X1 U11963 ( .A1(n12735), .A2(n12792), .ZN(n13306) );
  AND2_X1 U11964 ( .A1(n13305), .A2(n13306), .ZN(n9368) );
  NAND2_X1 U11965 ( .A1(n12811), .A2(n13349), .ZN(n13316) );
  NAND2_X1 U11966 ( .A1(n13550), .A2(n13322), .ZN(n12976) );
  NAND2_X1 U11967 ( .A1(n13316), .A2(n12976), .ZN(n13334) );
  NAND2_X1 U11968 ( .A1(n13306), .A2(n13334), .ZN(n13282) );
  NAND2_X1 U11969 ( .A1(n13538), .A2(n13288), .ZN(n13283) );
  INV_X1 U11970 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11783) );
  NAND2_X1 U11971 ( .A1(n11783), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9385) );
  INV_X1 U11972 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12484) );
  NAND2_X1 U11973 ( .A1(n12484), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9373) );
  NAND2_X1 U11974 ( .A1(n9385), .A2(n9373), .ZN(n9374) );
  NAND2_X1 U11975 ( .A1(n9375), .A2(n9374), .ZN(n9376) );
  NAND2_X1 U11976 ( .A1(n12863), .A2(SI_21_), .ZN(n9377) );
  NAND2_X1 U11977 ( .A1(n9378), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9379) );
  NAND2_X1 U11978 ( .A1(n9389), .A2(n9379), .ZN(n13292) );
  INV_X1 U11979 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13531) );
  NAND2_X1 U11980 ( .A1(n9466), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9381) );
  NAND2_X1 U11981 ( .A1(n12855), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n9380) );
  OAI211_X1 U11982 ( .C1(n13531), .C2(n12847), .A(n9381), .B(n9380), .ZN(n9382) );
  AOI21_X1 U11983 ( .B1(n13292), .B2(n9497), .A(n9382), .ZN(n9384) );
  INV_X1 U11984 ( .A(n12989), .ZN(n9525) );
  XNOR2_X1 U11985 ( .A(n11873), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n9398) );
  XNOR2_X1 U11986 ( .A(n9399), .B(n9398), .ZN(n11806) );
  NAND2_X1 U11987 ( .A1(n11806), .A2(n7262), .ZN(n9388) );
  NAND2_X1 U11988 ( .A1(n12863), .A2(SI_22_), .ZN(n9387) );
  NAND2_X1 U11989 ( .A1(n9389), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9390) );
  NAND2_X1 U11990 ( .A1(n9402), .A2(n9390), .ZN(n13277) );
  NAND2_X1 U11991 ( .A1(n13277), .A2(n9497), .ZN(n9395) );
  INV_X1 U11992 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13525) );
  NAND2_X1 U11993 ( .A1(n9466), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n9392) );
  NAND2_X1 U11994 ( .A1(n12855), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n9391) );
  OAI211_X1 U11995 ( .C1(n13525), .C2(n12847), .A(n9392), .B(n9391), .ZN(n9393) );
  INV_X1 U11996 ( .A(n9393), .ZN(n9394) );
  NAND2_X1 U11997 ( .A1(n13526), .A2(n13289), .ZN(n9397) );
  INV_X1 U11998 ( .A(n13526), .ZN(n9396) );
  XNOR2_X1 U11999 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n9409) );
  XNOR2_X1 U12000 ( .A(n9410), .B(n9409), .ZN(n11929) );
  NAND2_X1 U12001 ( .A1(n11929), .A2(n7262), .ZN(n9401) );
  NAND2_X1 U12002 ( .A1(n12863), .A2(SI_23_), .ZN(n9400) );
  NAND2_X1 U12003 ( .A1(n9402), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9403) );
  NAND2_X1 U12004 ( .A1(n9416), .A2(n9403), .ZN(n13264) );
  NAND2_X1 U12005 ( .A1(n13264), .A2(n9497), .ZN(n9408) );
  INV_X1 U12006 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13521) );
  NAND2_X1 U12007 ( .A1(n12855), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n9405) );
  INV_X1 U12008 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12512) );
  OR2_X1 U12009 ( .A1(n12858), .A2(n12512), .ZN(n9404) );
  OAI211_X1 U12010 ( .C1(n13521), .C2(n12847), .A(n9405), .B(n9404), .ZN(n9406) );
  INV_X1 U12011 ( .A(n9406), .ZN(n9407) );
  NAND2_X1 U12012 ( .A1(n12728), .A2(n12801), .ZN(n12994) );
  NAND2_X1 U12013 ( .A1(n12998), .A2(n12994), .ZN(n13263) );
  INV_X1 U12014 ( .A(n12728), .ZN(n13523) );
  INV_X1 U12015 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n12039) );
  INV_X1 U12016 ( .A(n9411), .ZN(n9412) );
  INV_X1 U12017 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12159) );
  NAND2_X1 U12018 ( .A1(n9412), .A2(n12159), .ZN(n9413) );
  INV_X1 U12019 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12161) );
  XNOR2_X1 U12020 ( .A(n9426), .B(n12161), .ZN(n12693) );
  NAND2_X1 U12021 ( .A1(n12693), .A2(n7262), .ZN(n9415) );
  NAND2_X1 U12022 ( .A1(n12863), .A2(SI_24_), .ZN(n9414) );
  INV_X1 U12023 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n12783) );
  NAND2_X1 U12024 ( .A1(n9416), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9417) );
  NAND2_X1 U12025 ( .A1(n9432), .A2(n9417), .ZN(n13252) );
  NAND2_X1 U12026 ( .A1(n13252), .A2(n9497), .ZN(n9423) );
  INV_X1 U12027 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13517) );
  NAND2_X1 U12028 ( .A1(n12855), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9420) );
  INV_X1 U12029 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n9418) );
  OR2_X1 U12030 ( .A1(n12858), .A2(n9418), .ZN(n9419) );
  OAI211_X1 U12031 ( .C1(n13517), .C2(n12847), .A(n9420), .B(n9419), .ZN(n9421) );
  INV_X1 U12032 ( .A(n9421), .ZN(n9422) );
  XNOR2_X1 U12033 ( .A(n9835), .B(n13259), .ZN(n13251) );
  NAND2_X1 U12034 ( .A1(n9835), .A2(n13259), .ZN(n9424) );
  INV_X1 U12035 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12549) );
  XNOR2_X1 U12036 ( .A(n12549), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n9427) );
  XNOR2_X1 U12037 ( .A(n9441), .B(n9427), .ZN(n13617) );
  NAND2_X1 U12038 ( .A1(n13617), .A2(n7262), .ZN(n9429) );
  NAND2_X1 U12039 ( .A1(n12863), .A2(SI_25_), .ZN(n9428) );
  INV_X1 U12040 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9430) );
  NAND2_X1 U12041 ( .A1(n9432), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9433) );
  NAND2_X1 U12042 ( .A1(n9447), .A2(n9433), .ZN(n13238) );
  NAND2_X1 U12043 ( .A1(n13238), .A2(n9497), .ZN(n9439) );
  INV_X1 U12044 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n9436) );
  NAND2_X1 U12045 ( .A1(n9466), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9435) );
  NAND2_X1 U12046 ( .A1(n12855), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9434) );
  OAI211_X1 U12047 ( .C1(n9436), .C2(n12847), .A(n9435), .B(n9434), .ZN(n9437)
         );
  INV_X1 U12048 ( .A(n9437), .ZN(n9438) );
  NAND2_X1 U12049 ( .A1(n13443), .A2(n13249), .ZN(n13008) );
  NAND2_X1 U12050 ( .A1(n13233), .A2(n13232), .ZN(n13231) );
  INV_X1 U12051 ( .A(n13443), .ZN(n13240) );
  NAND2_X1 U12052 ( .A1(n12549), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9440) );
  INV_X1 U12053 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12567) );
  NAND2_X1 U12054 ( .A1(n12567), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9442) );
  INV_X1 U12055 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14672) );
  XNOR2_X1 U12056 ( .A(n14672), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n9444) );
  XNOR2_X1 U12057 ( .A(n9458), .B(n9444), .ZN(n13613) );
  NAND2_X1 U12058 ( .A1(n13613), .A2(n7262), .ZN(n9446) );
  NAND2_X1 U12059 ( .A1(n12863), .A2(SI_26_), .ZN(n9445) );
  INV_X1 U12060 ( .A(n13438), .ZN(n12828) );
  NAND2_X1 U12061 ( .A1(n9447), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9448) );
  NAND2_X1 U12062 ( .A1(n9464), .A2(n9448), .ZN(n13225) );
  NAND2_X1 U12063 ( .A1(n13225), .A2(n9497), .ZN(n9454) );
  INV_X1 U12064 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n9451) );
  NAND2_X1 U12065 ( .A1(n12855), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9450) );
  NAND2_X1 U12066 ( .A1(n9176), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n9449) );
  OAI211_X1 U12067 ( .C1(n9451), .C2(n12858), .A(n9450), .B(n9449), .ZN(n9452)
         );
  INV_X1 U12068 ( .A(n9452), .ZN(n9453) );
  NAND2_X1 U12069 ( .A1(n12828), .A2(n12756), .ZN(n9456) );
  NOR2_X1 U12070 ( .A1(n12828), .A2(n12756), .ZN(n9455) );
  INV_X1 U12071 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15436) );
  AND2_X1 U12072 ( .A1(n15436), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9457) );
  NAND2_X1 U12073 ( .A1(n14672), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9459) );
  XNOR2_X1 U12074 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n9460) );
  XNOR2_X1 U12075 ( .A(n9475), .B(n9460), .ZN(n13608) );
  NAND2_X1 U12076 ( .A1(n13608), .A2(n7262), .ZN(n9462) );
  NAND2_X1 U12077 ( .A1(n12863), .A2(SI_27_), .ZN(n9461) );
  INV_X1 U12078 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9867) );
  NAND2_X1 U12079 ( .A1(n9464), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9465) );
  NAND2_X1 U12080 ( .A1(n9479), .A2(n9465), .ZN(n13208) );
  NAND2_X1 U12081 ( .A1(n13208), .A2(n9497), .ZN(n9472) );
  INV_X1 U12082 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n9469) );
  NAND2_X1 U12083 ( .A1(n12855), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9468) );
  NAND2_X1 U12084 ( .A1(n9466), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9467) );
  OAI211_X1 U12085 ( .C1(n9469), .C2(n12847), .A(n9468), .B(n9467), .ZN(n9470)
         );
  INV_X1 U12086 ( .A(n9470), .ZN(n9471) );
  NOR2_X1 U12087 ( .A1(n13207), .A2(n12823), .ZN(n13014) );
  INV_X1 U12088 ( .A(n13014), .ZN(n9473) );
  NAND2_X1 U12089 ( .A1(n10677), .A2(n13192), .ZN(n9485) );
  INV_X1 U12090 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14670) );
  AND2_X1 U12091 ( .A1(n14670), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9474) );
  XNOR2_X1 U12092 ( .A(n14667), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n9476) );
  NAND2_X1 U12093 ( .A1(n12568), .A2(n7262), .ZN(n9478) );
  NAND2_X1 U12094 ( .A1(n12863), .A2(SI_28_), .ZN(n9477) );
  NAND2_X1 U12095 ( .A1(n9479), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9480) );
  INV_X1 U12096 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n9483) );
  NAND2_X1 U12097 ( .A1(n12855), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9482) );
  NAND2_X1 U12098 ( .A1(n9466), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n9481) );
  OAI211_X1 U12099 ( .C1(n9483), .C2(n12847), .A(n9482), .B(n9481), .ZN(n9484)
         );
  XNOR2_X1 U12100 ( .A(n9485), .B(n13194), .ZN(n9507) );
  NAND2_X1 U12101 ( .A1(n9487), .A2(n9486), .ZN(n9489) );
  NAND2_X1 U12102 ( .A1(n9489), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9491) );
  INV_X1 U12103 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9490) );
  INV_X1 U12104 ( .A(n11699), .ZN(n9571) );
  AND2_X1 U12105 ( .A1(n9778), .A2(n9571), .ZN(n13025) );
  NAND2_X1 U12106 ( .A1(n9495), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9494) );
  MUX2_X1 U12107 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9494), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n9496) );
  INV_X1 U12108 ( .A(n13028), .ZN(n9532) );
  NOR2_X1 U12109 ( .A1(n13170), .A2(n9532), .ZN(n9572) );
  OR2_X2 U12110 ( .A1(n13025), .A2(n9572), .ZN(n15864) );
  INV_X1 U12111 ( .A(n13186), .ZN(n9498) );
  NAND2_X1 U12112 ( .A1(n9498), .A2(n9497), .ZN(n12861) );
  INV_X1 U12113 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n13510) );
  NAND2_X1 U12114 ( .A1(n9466), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9500) );
  NAND2_X1 U12115 ( .A1(n12855), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9499) );
  OAI211_X1 U12116 ( .C1(n13510), .C2(n12847), .A(n9500), .B(n9499), .ZN(n9501) );
  INV_X1 U12117 ( .A(n9501), .ZN(n9502) );
  INV_X1 U12118 ( .A(n9503), .ZN(n9686) );
  NAND2_X1 U12119 ( .A1(n9686), .A2(n13164), .ZN(n9609) );
  INV_X1 U12120 ( .A(n9505), .ZN(n9504) );
  OAI22_X1 U12121 ( .A1(n12868), .A2(n15859), .B1(n12823), .B2(n15861), .ZN(
        n9506) );
  AOI21_X2 U12122 ( .B1(n9507), .B2(n15864), .A(n9506), .ZN(n12699) );
  INV_X1 U12123 ( .A(n12879), .ZN(n9508) );
  NAND2_X1 U12124 ( .A1(n11476), .A2(n9508), .ZN(n9509) );
  NAND2_X1 U12125 ( .A1(n9509), .A2(n12904), .ZN(n11631) );
  INV_X1 U12126 ( .A(n12905), .ZN(n12881) );
  OR2_X1 U12127 ( .A1(n13040), .A2(n15885), .ZN(n12913) );
  NAND2_X1 U12128 ( .A1(n13039), .A2(n15892), .ZN(n9510) );
  NAND2_X1 U12129 ( .A1(n11772), .A2(n11614), .ZN(n9511) );
  NAND2_X1 U12130 ( .A1(n11950), .A2(n13035), .ZN(n12937) );
  OR2_X1 U12131 ( .A1(n11950), .A2(n13035), .ZN(n12936) );
  XNOR2_X1 U12132 ( .A(n12205), .B(n13034), .ZN(n13416) );
  NOR2_X1 U12133 ( .A1(n12205), .A2(n13034), .ZN(n12948) );
  INV_X1 U12134 ( .A(n12948), .ZN(n9512) );
  XNOR2_X1 U12135 ( .A(n12954), .B(n12531), .ZN(n13405) );
  NOR2_X1 U12136 ( .A1(n12954), .A2(n13421), .ZN(n12949) );
  NOR2_X1 U12137 ( .A1(n12896), .A2(n13381), .ZN(n9514) );
  NAND2_X1 U12138 ( .A1(n12896), .A2(n13381), .ZN(n9513) );
  OAI21_X1 U12139 ( .B1(n13388), .B2(n9514), .A(n9513), .ZN(n13364) );
  INV_X1 U12140 ( .A(n12959), .ZN(n9515) );
  INV_X1 U12141 ( .A(n12958), .ZN(n13365) );
  INV_X1 U12142 ( .A(n12961), .ZN(n9516) );
  INV_X1 U12143 ( .A(n13382), .ZN(n12765) );
  AOI21_X1 U12144 ( .B1(n13365), .B2(n9516), .A(n12966), .ZN(n9517) );
  AND2_X1 U12145 ( .A1(n12769), .A2(n13373), .ZN(n12962) );
  INV_X1 U12146 ( .A(n12962), .ZN(n12969) );
  NAND2_X1 U12147 ( .A1(n12969), .A2(n12968), .ZN(n13356) );
  NOR2_X1 U12148 ( .A1(n13556), .A2(n12810), .ZN(n12977) );
  INV_X1 U12149 ( .A(n12977), .ZN(n9518) );
  AND2_X1 U12150 ( .A1(n13316), .A2(n9518), .ZN(n13296) );
  AND2_X1 U12151 ( .A1(n13296), .A2(n13299), .ZN(n9519) );
  AND2_X1 U12152 ( .A1(n13556), .A2(n12810), .ZN(n12972) );
  INV_X1 U12153 ( .A(n12972), .ZN(n13314) );
  NAND2_X1 U12154 ( .A1(n13314), .A2(n13349), .ZN(n9520) );
  AOI22_X1 U12155 ( .A1(n13550), .A2(n9520), .B1(n12972), .B2(n13322), .ZN(
        n9521) );
  AND2_X1 U12156 ( .A1(n12981), .A2(n9521), .ZN(n13297) );
  INV_X1 U12157 ( .A(n13297), .ZN(n9522) );
  NAND2_X1 U12158 ( .A1(n9522), .A2(n13299), .ZN(n9523) );
  NAND2_X1 U12159 ( .A1(n13526), .A2(n12745), .ZN(n12995) );
  NAND2_X1 U12160 ( .A1(n9527), .A2(n12992), .ZN(n13262) );
  INV_X1 U12161 ( .A(n13263), .ZN(n12888) );
  NAND2_X1 U12162 ( .A1(n9835), .A2(n13237), .ZN(n12999) );
  INV_X1 U12163 ( .A(n13008), .ZN(n9529) );
  INV_X1 U12164 ( .A(n13012), .ZN(n9530) );
  NAND2_X1 U12165 ( .A1(n13438), .A2(n12756), .ZN(n13005) );
  NOR2_X1 U12166 ( .A1(n12867), .A2(n7771), .ZN(n9531) );
  OR2_X1 U12167 ( .A1(n9571), .A2(n9778), .ZN(n9533) );
  NAND2_X1 U12168 ( .A1(n9533), .A2(n9532), .ZN(n9536) );
  AOI21_X1 U12169 ( .B1(n11699), .B2(n13028), .A(n13170), .ZN(n9534) );
  OR2_X1 U12170 ( .A1(n9534), .A2(n9778), .ZN(n9535) );
  NAND2_X1 U12171 ( .A1(n9536), .A2(n9535), .ZN(n9859) );
  NAND2_X1 U12172 ( .A1(n9859), .A2(n15901), .ZN(n11083) );
  NAND2_X1 U12173 ( .A1(n11699), .A2(n13170), .ZN(n13022) );
  OR2_X1 U12174 ( .A1(n11083), .A2(n13022), .ZN(n9539) );
  AND2_X1 U12175 ( .A1(n13170), .A2(n13028), .ZN(n9537) );
  AND2_X1 U12176 ( .A1(n13022), .A2(n9537), .ZN(n10687) );
  INV_X1 U12177 ( .A(n10687), .ZN(n9538) );
  NAND2_X1 U12178 ( .A1(n6568), .A2(n15899), .ZN(n9540) );
  XNOR2_X1 U12179 ( .A(n9558), .B(P3_B_REG_SCAN_IN), .ZN(n9546) );
  NAND2_X1 U12180 ( .A1(n9546), .A2(n13620), .ZN(n9554) );
  INV_X1 U12181 ( .A(n9548), .ZN(n9549) );
  OAI21_X1 U12182 ( .B1(n9493), .B2(n9549), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n9550) );
  MUX2_X1 U12183 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9550), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n9552) );
  NAND2_X1 U12184 ( .A1(n9552), .A2(n9551), .ZN(n13616) );
  INV_X1 U12185 ( .A(n13616), .ZN(n9553) );
  OR2_X1 U12186 ( .A1(n9557), .A2(P3_D_REG_1__SCAN_IN), .ZN(n9556) );
  NAND2_X1 U12187 ( .A1(n13620), .A2(n13616), .ZN(n9555) );
  NAND2_X1 U12188 ( .A1(n9558), .A2(n13616), .ZN(n9559) );
  NOR4_X1 U12189 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_6__SCAN_IN), .A4(P3_D_REG_22__SCAN_IN), .ZN(n12508) );
  NOR2_X1 U12190 ( .A1(P3_D_REG_8__SCAN_IN), .A2(P3_D_REG_7__SCAN_IN), .ZN(
        n9562) );
  NOR4_X1 U12191 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_D_REG_25__SCAN_IN), .A3(
        P3_D_REG_20__SCAN_IN), .A4(P3_D_REG_27__SCAN_IN), .ZN(n9561) );
  NOR4_X1 U12192 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), .A3(
        P3_D_REG_17__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n9560) );
  NAND4_X1 U12193 ( .A1(n12508), .A2(n9562), .A3(n9561), .A4(n9560), .ZN(n9568) );
  NOR4_X1 U12194 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_11__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n9566) );
  NOR4_X1 U12195 ( .A1(P3_D_REG_24__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n9565) );
  NOR4_X1 U12196 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_2__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_4__SCAN_IN), .ZN(n9564) );
  NOR4_X1 U12197 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_3__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n9563) );
  NAND4_X1 U12198 ( .A1(n9566), .A2(n9565), .A3(n9564), .A4(n9563), .ZN(n9567)
         );
  NOR2_X1 U12199 ( .A1(n9568), .A2(n9567), .ZN(n9569) );
  INV_X1 U12200 ( .A(n10684), .ZN(n9570) );
  INV_X1 U12201 ( .A(n9778), .ZN(n11753) );
  INV_X1 U12202 ( .A(n9572), .ZN(n9573) );
  NAND3_X1 U12203 ( .A1(n11105), .A2(n11101), .A3(n10684), .ZN(n9870) );
  INV_X1 U12204 ( .A(n9859), .ZN(n9574) );
  OAI22_X1 U12205 ( .A1(n9860), .A2(n9854), .B1(n9870), .B2(n9574), .ZN(n9577)
         );
  NAND2_X1 U12206 ( .A1(n6566), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9576) );
  NAND2_X1 U12207 ( .A1(n9577), .A2(n10683), .ZN(n9580) );
  INV_X1 U12208 ( .A(n9860), .ZN(n9578) );
  NOR2_X1 U12209 ( .A1(n9852), .A2(n13022), .ZN(n9868) );
  AND2_X1 U12210 ( .A1(n9868), .A2(n13006), .ZN(n9864) );
  NAND2_X1 U12211 ( .A1(n9578), .A2(n9864), .ZN(n9579) );
  NOR2_X1 U12212 ( .A1(n15905), .A2(n9483), .ZN(n9582) );
  INV_X1 U12213 ( .A(n13123), .ZN(n9680) );
  INV_X1 U12214 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13360) );
  INV_X1 U12215 ( .A(n9657), .ZN(n11552) );
  INV_X1 U12216 ( .A(n9644), .ZN(n11185) );
  NAND2_X1 U12217 ( .A1(n12295), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9585) );
  AND2_X1 U12218 ( .A1(n9614), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9586) );
  INV_X1 U12219 ( .A(n9586), .ZN(n9587) );
  NAND2_X1 U12220 ( .A1(n11032), .A2(n9587), .ZN(n11132) );
  INV_X1 U12221 ( .A(n11145), .ZN(n10856) );
  NAND2_X1 U12222 ( .A1(n10856), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9588) );
  INV_X1 U12223 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n9590) );
  OR2_X1 U12224 ( .A1(n11158), .A2(n9590), .ZN(n9592) );
  NAND2_X1 U12225 ( .A1(n11158), .A2(n9590), .ZN(n9591) );
  INV_X1 U12226 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n9643) );
  XNOR2_X1 U12227 ( .A(n9644), .B(n9643), .ZN(n11180) );
  INV_X1 U12228 ( .A(n9593), .ZN(n11545) );
  INV_X1 U12229 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n12095) );
  XNOR2_X1 U12230 ( .A(n9657), .B(n12095), .ZN(n11546) );
  AOI21_X1 U12231 ( .B1(n9594), .B2(n9662), .A(n9595), .ZN(n11737) );
  INV_X1 U12232 ( .A(n9595), .ZN(n11889) );
  XNOR2_X1 U12233 ( .A(n10872), .B(P3_REG2_REG_10__SCAN_IN), .ZN(n11890) );
  INV_X1 U12234 ( .A(n10903), .ZN(n12106) );
  INV_X1 U12235 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n13424) );
  INV_X1 U12236 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n9596) );
  XNOR2_X1 U12237 ( .A(n10917), .B(n9596), .ZN(n13045) );
  INV_X1 U12238 ( .A(n10917), .ZN(n13052) );
  INV_X1 U12239 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13394) );
  INV_X1 U12240 ( .A(n13083), .ZN(n9599) );
  NAND2_X1 U12241 ( .A1(n13095), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9674) );
  OAI21_X1 U12242 ( .B1(n13095), .B2(P3_REG2_REG_14__SCAN_IN), .A(n9674), .ZN(
        n13082) );
  INV_X1 U12243 ( .A(n13082), .ZN(n9598) );
  NAND2_X1 U12244 ( .A1(n13084), .A2(n9674), .ZN(n9600) );
  NAND2_X1 U12245 ( .A1(n9600), .A2(n7404), .ZN(n9601) );
  INV_X1 U12246 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13374) );
  INV_X1 U12247 ( .A(n9601), .ZN(n13125) );
  XNOR2_X1 U12248 ( .A(n13123), .B(n13360), .ZN(n13124) );
  INV_X1 U12249 ( .A(n13151), .ZN(n11066) );
  INV_X1 U12250 ( .A(n13160), .ZN(n13175) );
  NAND2_X1 U12251 ( .A1(n13175), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n13158) );
  INV_X1 U12252 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13338) );
  NAND2_X1 U12253 ( .A1(n13160), .A2(n13338), .ZN(n9603) );
  AND2_X1 U12254 ( .A1(n13158), .A2(n9603), .ZN(n9604) );
  NAND2_X1 U12255 ( .A1(n13006), .A2(n9855), .ZN(n9606) );
  NAND2_X1 U12256 ( .A1(n9606), .A2(n9605), .ZN(n9689) );
  INV_X1 U12257 ( .A(n9855), .ZN(n9607) );
  NAND2_X1 U12258 ( .A1(n9607), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13031) );
  NAND2_X1 U12259 ( .A1(n9852), .A2(n13031), .ZN(n9688) );
  INV_X1 U12260 ( .A(n9688), .ZN(n9608) );
  INV_X1 U12261 ( .A(n9687), .ZN(n9611) );
  INV_X1 U12262 ( .A(n9609), .ZN(n9610) );
  AOI21_X1 U12263 ( .B1(n13159), .B2(n9612), .A(n13182), .ZN(n9613) );
  INV_X1 U12264 ( .A(n9613), .ZN(n9694) );
  XNOR2_X1 U12265 ( .A(n13160), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n13176) );
  NAND2_X1 U12266 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n10917), .ZN(n9627) );
  AOI22_X1 U12267 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n10917), .B1(n13052), 
        .B2(n13485), .ZN(n13055) );
  INV_X1 U12268 ( .A(n11158), .ZN(n9640) );
  NAND2_X1 U12269 ( .A1(n12295), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9615) );
  AND2_X1 U12270 ( .A1(n9614), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9616) );
  NAND2_X1 U12271 ( .A1(n11033), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9618) );
  INV_X1 U12272 ( .A(n9616), .ZN(n9617) );
  NAND2_X1 U12273 ( .A1(n9618), .A2(n9617), .ZN(n11138) );
  MUX2_X1 U12274 ( .A(n9619), .B(P3_REG1_REG_2__SCAN_IN), .S(n11145), .Z(
        n11139) );
  NAND2_X1 U12275 ( .A1(n10856), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9620) );
  XNOR2_X1 U12276 ( .A(n9622), .B(n11202), .ZN(n11196) );
  INV_X1 U12277 ( .A(n9622), .ZN(n9623) );
  INV_X1 U12278 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15915) );
  MUX2_X1 U12279 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n15915), .S(n9644), .Z(
        n11177) );
  XNOR2_X1 U12280 ( .A(n9624), .B(n9650), .ZN(n11294) );
  OAI22_X1 U12281 ( .A1(n11294), .A2(n9648), .B1(n9650), .B2(n9624), .ZN(
        n11544) );
  XNOR2_X1 U12282 ( .A(n9657), .B(P3_REG1_REG_8__SCAN_IN), .ZN(n11543) );
  INV_X1 U12283 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n13494) );
  XNOR2_X1 U12284 ( .A(n10872), .B(n13494), .ZN(n11886) );
  OR2_X1 U12285 ( .A1(n9625), .A2(n12106), .ZN(n9626) );
  NAND2_X1 U12286 ( .A1(n13095), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9675) );
  OAI21_X1 U12287 ( .B1(n13095), .B2(P3_REG1_REG_14__SCAN_IN), .A(n9675), .ZN(
        n13080) );
  INV_X1 U12288 ( .A(n13080), .ZN(n9629) );
  INV_X1 U12289 ( .A(n9675), .ZN(n9628) );
  NOR2_X1 U12290 ( .A1(n9630), .A2(n13111), .ZN(n13135) );
  INV_X1 U12291 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13471) );
  XNOR2_X1 U12292 ( .A(n13123), .B(n13471), .ZN(n13133) );
  NAND2_X1 U12293 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n13123), .ZN(n9631) );
  INV_X1 U12294 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13468) );
  NOR2_X2 U12295 ( .A1(n9687), .A2(n13164), .ZN(n13180) );
  MUX2_X1 U12296 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13612), .Z(n9681) );
  INV_X1 U12297 ( .A(n9635), .ZN(n9636) );
  XOR2_X1 U12298 ( .A(n10848), .B(n9635), .Z(n11037) );
  INV_X1 U12299 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11406) );
  MUX2_X1 U12300 ( .A(n11406), .B(n11325), .S(n13612), .Z(n11409) );
  NAND2_X1 U12301 ( .A1(n11409), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11403) );
  NOR2_X1 U12302 ( .A1(n11037), .A2(n11403), .ZN(n11036) );
  AOI21_X1 U12303 ( .B1(n10848), .B2(n9636), .A(n11036), .ZN(n11129) );
  MUX2_X1 U12304 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n13612), .Z(n9637) );
  XOR2_X1 U12305 ( .A(n11145), .B(n9637), .Z(n11130) );
  OAI22_X1 U12306 ( .A1(n11129), .A2(n11130), .B1(n9637), .B2(n10856), .ZN(
        n11113) );
  MUX2_X1 U12307 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n13612), .Z(n9638) );
  XNOR2_X1 U12308 ( .A(n9638), .B(n11124), .ZN(n11114) );
  INV_X1 U12309 ( .A(n9638), .ZN(n9639) );
  AOI22_X1 U12310 ( .A1(n11113), .A2(n11114), .B1(n11124), .B2(n9639), .ZN(
        n11147) );
  MUX2_X1 U12311 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n13612), .Z(n9641) );
  XOR2_X1 U12312 ( .A(n11158), .B(n9641), .Z(n11148) );
  MUX2_X1 U12313 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n13612), .Z(n9642) );
  NOR2_X1 U12314 ( .A1(n9642), .A2(n11202), .ZN(n11191) );
  NAND2_X1 U12315 ( .A1(n9642), .A2(n11202), .ZN(n11192) );
  MUX2_X1 U12316 ( .A(n9643), .B(n15915), .S(n13612), .Z(n9645) );
  NAND2_X1 U12317 ( .A1(n9645), .A2(n9644), .ZN(n11300) );
  INV_X1 U12318 ( .A(n9645), .ZN(n9646) );
  NAND2_X1 U12319 ( .A1(n9646), .A2(n11185), .ZN(n9647) );
  NAND2_X1 U12320 ( .A1(n11300), .A2(n9647), .ZN(n11174) );
  INV_X1 U12321 ( .A(n11300), .ZN(n9655) );
  INV_X1 U12322 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n9649) );
  MUX2_X1 U12323 ( .A(n9649), .B(n9648), .S(n13612), .Z(n9651) );
  NAND2_X1 U12324 ( .A1(n9651), .A2(n9650), .ZN(n11554) );
  INV_X1 U12325 ( .A(n9651), .ZN(n9652) );
  NAND2_X1 U12326 ( .A1(n9652), .A2(n11297), .ZN(n9653) );
  NAND2_X1 U12327 ( .A1(n11554), .A2(n9653), .ZN(n11299) );
  INV_X1 U12328 ( .A(n11299), .ZN(n9654) );
  MUX2_X1 U12329 ( .A(n12095), .B(n9656), .S(n13612), .Z(n9658) );
  NAND2_X1 U12330 ( .A1(n9658), .A2(n9657), .ZN(n9661) );
  INV_X1 U12331 ( .A(n9658), .ZN(n9659) );
  NAND2_X1 U12332 ( .A1(n9659), .A2(n11552), .ZN(n9660) );
  NAND2_X1 U12333 ( .A1(n9661), .A2(n9660), .ZN(n11553) );
  AOI21_X1 U12334 ( .B1(n11555), .B2(n11554), .A(n11553), .ZN(n11745) );
  INV_X1 U12335 ( .A(n9661), .ZN(n11744) );
  MUX2_X1 U12336 ( .A(n11948), .B(n12462), .S(n13612), .Z(n9663) );
  NAND2_X1 U12337 ( .A1(n9662), .A2(n9663), .ZN(n11898) );
  INV_X1 U12338 ( .A(n9663), .ZN(n9664) );
  NAND2_X1 U12339 ( .A1(n9664), .A2(n11740), .ZN(n9665) );
  AND2_X1 U12340 ( .A1(n11898), .A2(n9665), .ZN(n11743) );
  INV_X1 U12341 ( .A(n10872), .ZN(n11896) );
  MUX2_X1 U12342 ( .A(n12154), .B(n13494), .S(n13612), .Z(n9666) );
  NAND2_X1 U12343 ( .A1(n11896), .A2(n9666), .ZN(n9669) );
  INV_X1 U12344 ( .A(n9666), .ZN(n9667) );
  NAND2_X1 U12345 ( .A1(n10872), .A2(n9667), .ZN(n9668) );
  NAND2_X1 U12346 ( .A1(n9669), .A2(n9668), .ZN(n11897) );
  MUX2_X1 U12347 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13612), .Z(n9670) );
  XNOR2_X1 U12348 ( .A(n10903), .B(n9670), .ZN(n12102) );
  NOR2_X1 U12349 ( .A1(n10903), .A2(n9670), .ZN(n13058) );
  MUX2_X1 U12350 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n13612), .Z(n9671) );
  XNOR2_X1 U12351 ( .A(n9671), .B(n10917), .ZN(n13057) );
  NOR3_X1 U12352 ( .A1(n13059), .A2(n13058), .A3(n13057), .ZN(n13071) );
  INV_X1 U12353 ( .A(n9671), .ZN(n9672) );
  NOR2_X1 U12354 ( .A1(n9672), .A2(n13052), .ZN(n13070) );
  MUX2_X1 U12355 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13612), .Z(n9673) );
  XNOR2_X1 U12356 ( .A(n9673), .B(n10998), .ZN(n13069) );
  NOR2_X1 U12357 ( .A1(n9673), .A2(n10998), .ZN(n13088) );
  MUX2_X1 U12358 ( .A(n13080), .B(n13082), .S(n13164), .Z(n13087) );
  MUX2_X1 U12359 ( .A(n9675), .B(n9674), .S(n13164), .Z(n9676) );
  INV_X1 U12360 ( .A(n9677), .ZN(n9678) );
  MUX2_X1 U12361 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n13612), .Z(n13106) );
  NOR2_X1 U12362 ( .A1(n13107), .A2(n13106), .ZN(n13105) );
  MUX2_X1 U12363 ( .A(n13360), .B(n13471), .S(n13612), .Z(n9679) );
  NAND2_X1 U12364 ( .A1(n9680), .A2(n9679), .ZN(n13118) );
  XOR2_X1 U12365 ( .A(n9681), .B(n13151), .Z(n13148) );
  XNOR2_X1 U12366 ( .A(n13161), .B(n13160), .ZN(n9683) );
  MUX2_X1 U12367 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n13612), .Z(n9682) );
  OR2_X1 U12368 ( .A1(n9683), .A2(n9682), .ZN(n13163) );
  NAND2_X1 U12369 ( .A1(n9683), .A2(n9682), .ZN(n9684) );
  AOI21_X1 U12370 ( .B1(n13163), .B2(n9684), .A(n13146), .ZN(n9685) );
  INV_X1 U12371 ( .A(n9685), .ZN(n9693) );
  MUX2_X1 U12372 ( .A(n9687), .B(n13043), .S(n9686), .Z(n13171) );
  NAND2_X1 U12373 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12808)
         );
  NAND2_X1 U12374 ( .A1(n15849), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n9690) );
  OAI211_X1 U12375 ( .C1(n13171), .C2(n13175), .A(n12808), .B(n9690), .ZN(
        n9691) );
  INV_X1 U12376 ( .A(n9691), .ZN(n9692) );
  NAND4_X1 U12377 ( .A1(n9694), .A2(n6623), .A3(n9693), .A4(n9692), .ZN(
        P3_U3200) );
  INV_X1 U12378 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n13143) );
  INV_X1 U12379 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14944) );
  INV_X1 U12380 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9760) );
  AND2_X1 U12381 ( .A1(n9760), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n9713) );
  INV_X1 U12382 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n13104) );
  INV_X1 U12383 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n11623) );
  INV_X1 U12384 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n11603) );
  INV_X1 U12385 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n13050) );
  XOR2_X1 U12386 ( .A(n13050), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n9715) );
  INV_X1 U12387 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n12257) );
  INV_X1 U12388 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14932) );
  INV_X1 U12389 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n9708) );
  XOR2_X1 U12390 ( .A(n9708), .B(P1_ADDR_REG_9__SCAN_IN), .Z(n9717) );
  NAND2_X1 U12391 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n12249), .ZN(n9695) );
  NOR2_X1 U12392 ( .A1(n9698), .A2(n9697), .ZN(n9699) );
  NOR2_X1 U12393 ( .A1(n9701), .A2(n9700), .ZN(n9702) );
  INV_X1 U12394 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10922) );
  NOR2_X1 U12395 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n10932), .ZN(n9704) );
  INV_X1 U12396 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14916) );
  NOR2_X1 U12397 ( .A1(P3_ADDR_REG_8__SCAN_IN), .A2(n9706), .ZN(n9707) );
  NOR2_X1 U12398 ( .A1(n14932), .A2(n9709), .ZN(n9710) );
  INV_X1 U12399 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n12101) );
  AOI22_X1 U12400 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P3_ADDR_REG_11__SCAN_IN), 
        .B1(n12101), .B2(n12257), .ZN(n9749) );
  NAND2_X1 U12401 ( .A1(n9715), .A2(n9714), .ZN(n9711) );
  INV_X1 U12402 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n13068) );
  NAND2_X1 U12403 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n13068), .ZN(n9712) );
  XNOR2_X1 U12404 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(n11623), .ZN(n9753) );
  INV_X1 U12405 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n11879) );
  NOR2_X1 U12406 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n11879), .ZN(n9756) );
  XOR2_X1 U12407 ( .A(n9715), .B(n9714), .Z(n15476) );
  INV_X1 U12408 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n15474) );
  XOR2_X1 U12409 ( .A(n9717), .B(n9716), .Z(n15459) );
  XOR2_X1 U12410 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9718), .Z(n15927) );
  XOR2_X1 U12411 ( .A(n9719), .B(P1_ADDR_REG_3__SCAN_IN), .Z(n15930) );
  XNOR2_X1 U12412 ( .A(n9720), .B(n6670), .ZN(n9725) );
  AOI21_X1 U12413 ( .B1(n11405), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n9721), .ZN(
        n9722) );
  INV_X1 U12414 ( .A(n9722), .ZN(n15924) );
  NAND2_X1 U12415 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15924), .ZN(n15934) );
  INV_X1 U12416 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n15452) );
  NAND2_X1 U12417 ( .A1(n15930), .A2(n15929), .ZN(n9726) );
  INV_X1 U12418 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n15625) );
  NAND2_X1 U12419 ( .A1(n9731), .A2(n9730), .ZN(n9733) );
  INV_X1 U12420 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15922) );
  XOR2_X1 U12421 ( .A(n10932), .B(P3_ADDR_REG_6__SCAN_IN), .Z(n9734) );
  XNOR2_X1 U12422 ( .A(n9735), .B(n9734), .ZN(n15454) );
  NOR2_X1 U12423 ( .A1(n9736), .A2(n7735), .ZN(n9737) );
  INV_X1 U12424 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10957) );
  XOR2_X1 U12425 ( .A(n10957), .B(n9740), .Z(n9741) );
  NAND2_X1 U12426 ( .A1(n9742), .A2(n9741), .ZN(n9743) );
  INV_X1 U12427 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n15663) );
  XNOR2_X1 U12428 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n9745), .ZN(n15464) );
  XOR2_X1 U12429 ( .A(n9749), .B(n9748), .Z(n9750) );
  XOR2_X1 U12430 ( .A(n13068), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n9752) );
  XOR2_X1 U12431 ( .A(n9752), .B(n9751), .Z(n15480) );
  XOR2_X1 U12432 ( .A(n9754), .B(n9753), .Z(n15484) );
  AOI21_X1 U12433 ( .B1(P3_ADDR_REG_15__SCAN_IN), .B2(n11879), .A(n9756), .ZN(
        n9758) );
  XNOR2_X1 U12434 ( .A(n9758), .B(n9757), .ZN(n15488) );
  NAND2_X1 U12435 ( .A1(n15489), .A2(n15488), .ZN(n9759) );
  XNOR2_X1 U12436 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n9760), .ZN(n9761) );
  XNOR2_X1 U12437 ( .A(n9762), .B(n9761), .ZN(n15493) );
  INV_X1 U12438 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n9768) );
  XOR2_X1 U12439 ( .A(n9768), .B(P1_ADDR_REG_18__SCAN_IN), .Z(n9767) );
  NOR2_X1 U12440 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n9763), .ZN(n9766) );
  NOR2_X1 U12441 ( .A1(n13143), .A2(n9764), .ZN(n9765) );
  INV_X1 U12442 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14958) );
  NAND2_X1 U12443 ( .A1(P3_ADDR_REG_18__SCAN_IN), .A2(n14958), .ZN(n9769) );
  AOI22_X1 U12444 ( .A1(n9770), .A2(n9769), .B1(P1_ADDR_REG_18__SCAN_IN), .B2(
        n9768), .ZN(n9771) );
  INV_X1 U12445 ( .A(n9771), .ZN(n9774) );
  XNOR2_X1 U12446 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n9772) );
  XNOR2_X1 U12447 ( .A(n9772), .B(n6983), .ZN(n9773) );
  INV_X1 U12448 ( .A(n13024), .ZN(n9776) );
  NAND2_X1 U12449 ( .A1(n9777), .A2(n9776), .ZN(n9780) );
  OAI21_X1 U12450 ( .B1(n9778), .B2(n13170), .A(n11699), .ZN(n9779) );
  NAND2_X4 U12451 ( .A1(n9780), .A2(n9779), .ZN(n9834) );
  XNOR2_X1 U12452 ( .A(n13207), .B(n9781), .ZN(n12577) );
  NOR2_X1 U12453 ( .A1(n12577), .A2(n13217), .ZN(n12573) );
  AOI21_X1 U12454 ( .B1(n12577), .B2(n13217), .A(n12573), .ZN(n9850) );
  XNOR2_X1 U12455 ( .A(n13556), .B(n12571), .ZN(n9823) );
  XNOR2_X1 U12456 ( .A(n12769), .B(n12571), .ZN(n9821) );
  INV_X1 U12457 ( .A(n9821), .ZN(n9822) );
  XNOR2_X1 U12458 ( .A(n12896), .B(n12571), .ZN(n12239) );
  INV_X1 U12459 ( .A(n12239), .ZN(n9816) );
  XNOR2_X1 U12460 ( .A(n9834), .B(n7250), .ZN(n9785) );
  XNOR2_X1 U12461 ( .A(n9785), .B(n13041), .ZN(n11331) );
  XNOR2_X1 U12462 ( .A(n9834), .B(n11283), .ZN(n9782) );
  NAND2_X1 U12463 ( .A1(n9782), .A2(n11668), .ZN(n11328) );
  AND2_X1 U12464 ( .A1(n11331), .A2(n11328), .ZN(n9784) );
  XNOR2_X1 U12465 ( .A(n9782), .B(n9055), .ZN(n11280) );
  OAI21_X1 U12466 ( .B1(n9834), .B2(n11662), .A(n12897), .ZN(n11094) );
  NAND2_X1 U12467 ( .A1(n11095), .A2(n11094), .ZN(n11093) );
  INV_X1 U12468 ( .A(n11095), .ZN(n9783) );
  NAND2_X1 U12469 ( .A1(n11280), .A2(n11279), .ZN(n11329) );
  INV_X1 U12470 ( .A(n9785), .ZN(n9786) );
  NAND2_X1 U12471 ( .A1(n9786), .A2(n13041), .ZN(n9787) );
  XNOR2_X1 U12472 ( .A(n9834), .B(n11531), .ZN(n9788) );
  INV_X1 U12473 ( .A(n13040), .ZN(n11612) );
  NAND2_X1 U12474 ( .A1(n9788), .A2(n11612), .ZN(n9792) );
  INV_X1 U12475 ( .A(n9788), .ZN(n9789) );
  NAND2_X1 U12476 ( .A1(n9789), .A2(n13040), .ZN(n9790) );
  NAND2_X1 U12477 ( .A1(n9792), .A2(n9790), .ZN(n11525) );
  NAND2_X1 U12478 ( .A1(n11523), .A2(n9792), .ZN(n11607) );
  XNOR2_X1 U12479 ( .A(n9834), .B(n11614), .ZN(n9793) );
  XNOR2_X1 U12480 ( .A(n9793), .B(n13039), .ZN(n11608) );
  XNOR2_X1 U12481 ( .A(n9834), .B(n15896), .ZN(n11767) );
  NAND2_X1 U12482 ( .A1(n9793), .A2(n11772), .ZN(n11765) );
  XNOR2_X1 U12483 ( .A(n9834), .B(n9794), .ZN(n9798) );
  NAND2_X1 U12484 ( .A1(n11766), .A2(n9796), .ZN(n9802) );
  INV_X1 U12485 ( .A(n11955), .ZN(n9797) );
  OAI21_X1 U12486 ( .B1(n11958), .B2(n6954), .A(n9797), .ZN(n9800) );
  NAND2_X1 U12487 ( .A1(n11767), .A2(n13038), .ZN(n11809) );
  OAI21_X1 U12488 ( .B1(n11958), .B2(n11809), .A(n11955), .ZN(n9799) );
  AOI22_X1 U12489 ( .A1(n9800), .A2(n9799), .B1(n9798), .B2(n13036), .ZN(n9801) );
  NAND2_X1 U12490 ( .A1(n9802), .A2(n9801), .ZN(n11819) );
  XNOR2_X1 U12491 ( .A(n9834), .B(n11950), .ZN(n9804) );
  XNOR2_X1 U12492 ( .A(n9804), .B(n13035), .ZN(n11820) );
  INV_X1 U12493 ( .A(n11820), .ZN(n9803) );
  XNOR2_X1 U12494 ( .A(n9834), .B(n13598), .ZN(n9807) );
  XNOR2_X1 U12495 ( .A(n9807), .B(n12207), .ZN(n11856) );
  INV_X1 U12496 ( .A(n9804), .ZN(n9805) );
  NAND2_X1 U12497 ( .A1(n9805), .A2(n12148), .ZN(n11853) );
  AND2_X1 U12498 ( .A1(n11856), .A2(n11853), .ZN(n9806) );
  NAND2_X1 U12499 ( .A1(n9807), .A2(n13423), .ZN(n9808) );
  XNOR2_X1 U12500 ( .A(n12205), .B(n12571), .ZN(n12526) );
  XNOR2_X1 U12501 ( .A(n12954), .B(n9781), .ZN(n12530) );
  NAND2_X1 U12502 ( .A1(n12530), .A2(n12531), .ZN(n12529) );
  INV_X1 U12503 ( .A(n9809), .ZN(n9810) );
  AOI21_X1 U12504 ( .B1(n12526), .B2(n13034), .A(n13421), .ZN(n9812) );
  NAND3_X1 U12505 ( .A1(n12526), .A2(n13421), .A3(n13034), .ZN(n9811) );
  NAND2_X1 U12506 ( .A1(n12241), .A2(n9814), .ZN(n9815) );
  XNOR2_X1 U12507 ( .A(n13574), .B(n12571), .ZN(n9817) );
  XNOR2_X1 U12508 ( .A(n9817), .B(n13392), .ZN(n12540) );
  INV_X1 U12509 ( .A(n9817), .ZN(n9818) );
  XNOR2_X1 U12510 ( .A(n12843), .B(n12571), .ZN(n9819) );
  NOR2_X1 U12511 ( .A1(n9819), .A2(n13382), .ZN(n9820) );
  AOI21_X1 U12512 ( .B1(n9819), .B2(n13382), .A(n9820), .ZN(n12831) );
  INV_X1 U12513 ( .A(n9820), .ZN(n12760) );
  XNOR2_X1 U12514 ( .A(n9821), .B(n13373), .ZN(n12761) );
  XNOR2_X1 U12515 ( .A(n9823), .B(n13358), .ZN(n12771) );
  XNOR2_X1 U12516 ( .A(n12811), .B(n12571), .ZN(n9824) );
  XNOR2_X1 U12517 ( .A(n9824), .B(n13322), .ZN(n12806) );
  XNOR2_X1 U12518 ( .A(n12735), .B(n12571), .ZN(n12731) );
  NOR2_X1 U12519 ( .A1(n12731), .A2(n13336), .ZN(n9826) );
  INV_X1 U12520 ( .A(n12731), .ZN(n9825) );
  XNOR2_X1 U12521 ( .A(n13538), .B(n12571), .ZN(n9827) );
  XNOR2_X1 U12522 ( .A(n9827), .B(n13288), .ZN(n12788) );
  INV_X1 U12523 ( .A(n9827), .ZN(n9828) );
  XNOR2_X1 U12524 ( .A(n13532), .B(n9781), .ZN(n9829) );
  NOR2_X1 U12525 ( .A1(n9829), .A2(n6797), .ZN(n9830) );
  AOI21_X1 U12526 ( .B1(n9829), .B2(n6797), .A(n9830), .ZN(n12742) );
  XNOR2_X1 U12527 ( .A(n13526), .B(n12571), .ZN(n9832) );
  XNOR2_X1 U12528 ( .A(n9835), .B(n9834), .ZN(n9837) );
  NAND2_X1 U12529 ( .A1(n9837), .A2(n13237), .ZN(n9842) );
  XNOR2_X1 U12530 ( .A(n12728), .B(n12571), .ZN(n12722) );
  NAND2_X1 U12531 ( .A1(n12722), .A2(n12801), .ZN(n12749) );
  XNOR2_X1 U12532 ( .A(n13443), .B(n9781), .ZN(n9836) );
  NOR2_X1 U12533 ( .A1(n9836), .A2(n13218), .ZN(n9845) );
  AOI21_X1 U12534 ( .B1(n9836), .B2(n13218), .A(n9845), .ZN(n12751) );
  INV_X1 U12535 ( .A(n9837), .ZN(n9838) );
  NAND2_X1 U12536 ( .A1(n9838), .A2(n13259), .ZN(n9839) );
  NAND2_X1 U12537 ( .A1(n9842), .A2(n9839), .ZN(n12779) );
  INV_X1 U12538 ( .A(n12722), .ZN(n9840) );
  AND2_X1 U12539 ( .A1(n9840), .A2(n13274), .ZN(n9841) );
  INV_X1 U12540 ( .A(n9845), .ZN(n9846) );
  XNOR2_X1 U12541 ( .A(n13438), .B(n9781), .ZN(n9847) );
  NOR2_X1 U12542 ( .A1(n9847), .A2(n13234), .ZN(n9848) );
  AOI21_X1 U12543 ( .B1(n9847), .B2(n13234), .A(n9848), .ZN(n12819) );
  NAND2_X1 U12544 ( .A1(n12818), .A2(n12819), .ZN(n12817) );
  INV_X1 U12545 ( .A(n9848), .ZN(n9849) );
  OAI22_X1 U12546 ( .A1(n9860), .A2(n11083), .B1(n9870), .B2(n9854), .ZN(n9851) );
  NAND2_X1 U12547 ( .A1(n9860), .A2(n13023), .ZN(n9853) );
  INV_X1 U12548 ( .A(n9854), .ZN(n9858) );
  NAND2_X1 U12549 ( .A1(n13006), .A2(n13022), .ZN(n10688) );
  NAND3_X1 U12550 ( .A1(n10688), .A2(n9856), .A3(n9855), .ZN(n9857) );
  AOI21_X1 U12551 ( .B1(n9870), .B2(n9858), .A(n9857), .ZN(n9862) );
  NAND2_X1 U12552 ( .A1(n9860), .A2(n9859), .ZN(n9861) );
  NAND2_X1 U12553 ( .A1(n9862), .A2(n9861), .ZN(n9863) );
  NAND2_X1 U12554 ( .A1(n9863), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9866) );
  NAND2_X1 U12555 ( .A1(n9870), .A2(n9864), .ZN(n9865) );
  NAND2_X1 U12556 ( .A1(n9868), .A2(n13422), .ZN(n13027) );
  OAI22_X1 U12557 ( .A1(n12756), .A2(n12836), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9867), .ZN(n9872) );
  INV_X1 U12558 ( .A(n9868), .ZN(n9869) );
  NOR2_X1 U12559 ( .A1(n13201), .A2(n12822), .ZN(n9871) );
  AOI211_X1 U12560 ( .C1(n13208), .C2(n12839), .A(n9872), .B(n9871), .ZN(n9873) );
  OAI21_X1 U12561 ( .B1(n10700), .B2(n12842), .A(n9873), .ZN(n9874) );
  INV_X1 U12562 ( .A(n9874), .ZN(n9875) );
  NAND2_X1 U12563 ( .A1(n9876), .A2(n9875), .ZN(P3_U3154) );
  INV_X2 U12564 ( .A(n10059), .ZN(n9886) );
  NAND2_X1 U12565 ( .A1(n8898), .A2(n10098), .ZN(n9879) );
  INV_X1 U12566 ( .A(n15228), .ZN(n14843) );
  NAND2_X1 U12567 ( .A1(n14843), .A2(n6513), .ZN(n9878) );
  NAND2_X1 U12568 ( .A1(n9879), .A2(n9878), .ZN(n9880) );
  XNOR2_X1 U12569 ( .A(n9880), .B(n10123), .ZN(n10010) );
  NAND2_X1 U12570 ( .A1(n8898), .A2(n6513), .ZN(n9882) );
  AND2_X2 U12571 ( .A1(n9886), .A2(n15138), .ZN(n9893) );
  NAND2_X1 U12572 ( .A1(n14843), .A2(n9996), .ZN(n9881) );
  NAND2_X1 U12573 ( .A1(n9882), .A2(n9881), .ZN(n14824) );
  NAND2_X1 U12574 ( .A1(n9893), .A2(n14856), .ZN(n9884) );
  INV_X1 U12575 ( .A(n10724), .ZN(n9885) );
  AOI22_X1 U12576 ( .A1(n10108), .A2(n11055), .B1(n9885), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n9883) );
  AND2_X1 U12577 ( .A1(n9884), .A2(n9883), .ZN(n11057) );
  NAND2_X1 U12578 ( .A1(n14856), .A2(n10108), .ZN(n9888) );
  AOI22_X1 U12579 ( .A1(n9886), .A2(n11055), .B1(n9885), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n9887) );
  NAND2_X1 U12580 ( .A1(n9888), .A2(n9887), .ZN(n11056) );
  NAND2_X1 U12581 ( .A1(n11057), .A2(n11056), .ZN(n9891) );
  INV_X1 U12582 ( .A(n11056), .ZN(n9889) );
  OR2_X1 U12583 ( .A1(n15535), .A2(n9953), .ZN(n9894) );
  NAND2_X1 U12584 ( .A1(n9895), .A2(n9894), .ZN(n9896) );
  INV_X1 U12585 ( .A(n9896), .ZN(n9897) );
  NAND2_X1 U12586 ( .A1(n9898), .A2(n9897), .ZN(n9899) );
  NAND2_X1 U12587 ( .A1(n14710), .A2(n9899), .ZN(n11024) );
  OR2_X1 U12588 ( .A1(n8299), .A2(n10059), .ZN(n9900) );
  NAND2_X1 U12589 ( .A1(n9901), .A2(n9900), .ZN(n9902) );
  NAND2_X1 U12590 ( .A1(n9893), .A2(n14855), .ZN(n9904) );
  OR2_X1 U12591 ( .A1(n8299), .A2(n9953), .ZN(n9903) );
  NAND2_X1 U12592 ( .A1(n9904), .A2(n9903), .ZN(n9905) );
  XNOR2_X1 U12593 ( .A(n9907), .B(n9905), .ZN(n11025) );
  INV_X1 U12594 ( .A(n9905), .ZN(n9906) );
  NAND2_X1 U12595 ( .A1(n9907), .A2(n9906), .ZN(n9908) );
  NAND2_X1 U12596 ( .A1(n14854), .A2(n10108), .ZN(n9910) );
  OR2_X1 U12597 ( .A1(n15502), .A2(n10059), .ZN(n9909) );
  NAND2_X1 U12598 ( .A1(n9910), .A2(n9909), .ZN(n9911) );
  XNOR2_X1 U12599 ( .A(n9911), .B(n10123), .ZN(n9914) );
  NAND2_X1 U12600 ( .A1(n9893), .A2(n14854), .ZN(n9913) );
  OR2_X1 U12601 ( .A1(n15502), .A2(n9953), .ZN(n9912) );
  NAND2_X1 U12602 ( .A1(n9913), .A2(n9912), .ZN(n9915) );
  NAND2_X1 U12603 ( .A1(n9914), .A2(n9915), .ZN(n9920) );
  INV_X1 U12604 ( .A(n9914), .ZN(n9917) );
  INV_X1 U12605 ( .A(n9915), .ZN(n9916) );
  NAND2_X1 U12606 ( .A1(n9917), .A2(n9916), .ZN(n9918) );
  NAND2_X1 U12607 ( .A1(n9920), .A2(n9918), .ZN(n15497) );
  NAND2_X1 U12608 ( .A1(n15505), .A2(n9920), .ZN(n9924) );
  INV_X2 U12609 ( .A(n9893), .ZN(n10091) );
  NAND2_X1 U12610 ( .A1(n15554), .A2(n6513), .ZN(n9921) );
  OAI21_X1 U12611 ( .B1(n11489), .B2(n10091), .A(n9921), .ZN(n9925) );
  NAND2_X1 U12612 ( .A1(n15554), .A2(n9886), .ZN(n9922) );
  OAI21_X1 U12613 ( .B1(n11489), .B2(n9953), .A(n9922), .ZN(n9923) );
  XNOR2_X1 U12614 ( .A(n9923), .B(n10111), .ZN(n11346) );
  INV_X1 U12615 ( .A(n9925), .ZN(n9926) );
  NAND2_X1 U12616 ( .A1(n11500), .A2(n9886), .ZN(n9928) );
  NAND2_X1 U12617 ( .A1(n14852), .A2(n10108), .ZN(n9927) );
  NAND2_X1 U12618 ( .A1(n9928), .A2(n9927), .ZN(n9929) );
  XNOR2_X1 U12619 ( .A(n9929), .B(n10111), .ZN(n11354) );
  NAND2_X1 U12620 ( .A1(n11500), .A2(n10108), .ZN(n9931) );
  NAND2_X1 U12621 ( .A1(n14852), .A2(n9893), .ZN(n9930) );
  AND2_X1 U12622 ( .A1(n9931), .A2(n9930), .ZN(n11353) );
  AND2_X1 U12623 ( .A1(n11354), .A2(n11353), .ZN(n9932) );
  NAND2_X1 U12624 ( .A1(n11576), .A2(n9886), .ZN(n9934) );
  NAND2_X1 U12625 ( .A1(n14851), .A2(n10108), .ZN(n9933) );
  NAND2_X1 U12626 ( .A1(n9934), .A2(n9933), .ZN(n9935) );
  XNOR2_X1 U12627 ( .A(n9935), .B(n10123), .ZN(n9938) );
  NAND2_X1 U12628 ( .A1(n11576), .A2(n10108), .ZN(n9937) );
  NAND2_X1 U12629 ( .A1(n14851), .A2(n9893), .ZN(n9936) );
  NAND2_X1 U12630 ( .A1(n9937), .A2(n9936), .ZN(n9939) );
  AND2_X1 U12631 ( .A1(n9938), .A2(n9939), .ZN(n11513) );
  INV_X1 U12632 ( .A(n11513), .ZN(n9942) );
  INV_X1 U12633 ( .A(n9938), .ZN(n9941) );
  INV_X1 U12634 ( .A(n9939), .ZN(n9940) );
  NAND2_X1 U12635 ( .A1(n11700), .A2(n9886), .ZN(n9944) );
  NAND2_X1 U12636 ( .A1(n14849), .A2(n10108), .ZN(n9943) );
  NAND2_X1 U12637 ( .A1(n9944), .A2(n9943), .ZN(n9945) );
  XNOR2_X1 U12638 ( .A(n9945), .B(n10123), .ZN(n9949) );
  NOR2_X1 U12639 ( .A1(n11677), .A2(n10091), .ZN(n9946) );
  AOI21_X1 U12640 ( .B1(n11700), .B2(n6513), .A(n9946), .ZN(n9947) );
  XNOR2_X1 U12641 ( .A(n9949), .B(n9947), .ZN(n11702) );
  INV_X1 U12642 ( .A(n9947), .ZN(n9948) );
  NAND2_X1 U12643 ( .A1(n15581), .A2(n10098), .ZN(n9951) );
  NAND2_X1 U12644 ( .A1(n14848), .A2(n6513), .ZN(n9950) );
  NAND2_X1 U12645 ( .A1(n9951), .A2(n9950), .ZN(n9952) );
  XNOR2_X1 U12646 ( .A(n9952), .B(n10111), .ZN(n9957) );
  NOR2_X1 U12647 ( .A1(n11832), .A2(n10091), .ZN(n9954) );
  AOI21_X1 U12648 ( .B1(n15581), .B2(n6513), .A(n9954), .ZN(n9956) );
  XNOR2_X1 U12649 ( .A(n9957), .B(n9956), .ZN(n11865) );
  INV_X1 U12650 ( .A(n11865), .ZN(n9955) );
  NAND2_X1 U12651 ( .A1(n9957), .A2(n9956), .ZN(n9958) );
  NAND2_X1 U12652 ( .A1(n15391), .A2(n9886), .ZN(n9960) );
  NAND2_X1 U12653 ( .A1(n14846), .A2(n6513), .ZN(n9959) );
  NAND2_X1 U12654 ( .A1(n9960), .A2(n9959), .ZN(n9961) );
  XNOR2_X1 U12655 ( .A(n9961), .B(n10123), .ZN(n12179) );
  NOR2_X1 U12656 ( .A1(n12169), .A2(n10091), .ZN(n9962) );
  AOI21_X1 U12657 ( .B1(n15391), .B2(n6513), .A(n9962), .ZN(n12178) );
  INV_X1 U12658 ( .A(n12178), .ZN(n9968) );
  NAND2_X1 U12659 ( .A1(n15396), .A2(n6513), .ZN(n9964) );
  NAND2_X1 U12660 ( .A1(n14847), .A2(n9996), .ZN(n9963) );
  INV_X1 U12661 ( .A(n12175), .ZN(n12060) );
  NAND2_X1 U12662 ( .A1(n15396), .A2(n9886), .ZN(n9966) );
  NAND2_X1 U12663 ( .A1(n14847), .A2(n6513), .ZN(n9965) );
  NAND2_X1 U12664 ( .A1(n9966), .A2(n9965), .ZN(n9967) );
  XNOR2_X1 U12665 ( .A(n9967), .B(n10111), .ZN(n12176) );
  INV_X1 U12666 ( .A(n12176), .ZN(n12061) );
  OAI22_X1 U12667 ( .A1(n12179), .A2(n9968), .B1(n12060), .B2(n12061), .ZN(
        n9972) );
  OAI21_X1 U12668 ( .B1(n12176), .B2(n12175), .A(n12178), .ZN(n9970) );
  AND2_X1 U12669 ( .A1(n9968), .A2(n12060), .ZN(n9969) );
  AOI22_X1 U12670 ( .A1(n9970), .A2(n12179), .B1(n9969), .B2(n12061), .ZN(
        n9971) );
  NAND2_X1 U12671 ( .A1(n15384), .A2(n9886), .ZN(n9974) );
  NAND2_X1 U12672 ( .A1(n14845), .A2(n6513), .ZN(n9973) );
  NAND2_X1 U12673 ( .A1(n9974), .A2(n9973), .ZN(n9975) );
  XNOR2_X1 U12674 ( .A(n9975), .B(n10111), .ZN(n9977) );
  NOR2_X1 U12675 ( .A1(n14729), .A2(n10091), .ZN(n9976) );
  AOI21_X1 U12676 ( .B1(n15384), .B2(n6513), .A(n9976), .ZN(n9978) );
  NAND2_X1 U12677 ( .A1(n9977), .A2(n9978), .ZN(n9983) );
  INV_X1 U12678 ( .A(n9977), .ZN(n9980) );
  INV_X1 U12679 ( .A(n9978), .ZN(n9979) );
  NAND2_X1 U12680 ( .A1(n9980), .A2(n9979), .ZN(n9981) );
  NAND2_X1 U12681 ( .A1(n9983), .A2(n9981), .ZN(n12166) );
  INV_X1 U12682 ( .A(n12166), .ZN(n9982) );
  NAND2_X1 U12683 ( .A1(n8965), .A2(n10098), .ZN(n9985) );
  NAND2_X1 U12684 ( .A1(n15255), .A2(n6513), .ZN(n9984) );
  NAND2_X1 U12685 ( .A1(n9985), .A2(n9984), .ZN(n9986) );
  XNOR2_X1 U12686 ( .A(n9986), .B(n10123), .ZN(n14683) );
  NAND2_X1 U12687 ( .A1(n8965), .A2(n6513), .ZN(n9988) );
  NAND2_X1 U12688 ( .A1(n9996), .A2(n15255), .ZN(n9987) );
  NAND2_X1 U12689 ( .A1(n9988), .A2(n9987), .ZN(n10003) );
  NAND2_X1 U12690 ( .A1(n14788), .A2(n9886), .ZN(n9990) );
  NAND2_X1 U12691 ( .A1(n14844), .A2(n6513), .ZN(n9989) );
  NAND2_X1 U12692 ( .A1(n9990), .A2(n9989), .ZN(n9991) );
  XNOR2_X1 U12693 ( .A(n9991), .B(n10123), .ZN(n14680) );
  NAND2_X1 U12694 ( .A1(n14788), .A2(n10108), .ZN(n9993) );
  NAND2_X1 U12695 ( .A1(n14844), .A2(n9996), .ZN(n9992) );
  NAND2_X1 U12696 ( .A1(n9993), .A2(n9992), .ZN(n14678) );
  NAND2_X1 U12697 ( .A1(n14680), .A2(n14678), .ZN(n14681) );
  NAND2_X1 U12698 ( .A1(n15258), .A2(n6513), .ZN(n9994) );
  NAND2_X1 U12699 ( .A1(n14724), .A2(n10108), .ZN(n9998) );
  NAND2_X1 U12700 ( .A1(n15258), .A2(n9996), .ZN(n9997) );
  NAND2_X1 U12701 ( .A1(n9998), .A2(n9997), .ZN(n10002) );
  NAND2_X1 U12702 ( .A1(n14677), .A2(n10002), .ZN(n9999) );
  INV_X1 U12703 ( .A(n14683), .ZN(n10008) );
  INV_X1 U12704 ( .A(n10002), .ZN(n14676) );
  INV_X1 U12705 ( .A(n14680), .ZN(n10001) );
  OR3_X1 U12706 ( .A1(n14677), .A2(n14678), .A3(n10002), .ZN(n10004) );
  INV_X1 U12707 ( .A(n10003), .ZN(n14682) );
  NAND2_X1 U12708 ( .A1(n10005), .A2(n10004), .ZN(n10006) );
  INV_X1 U12709 ( .A(n10010), .ZN(n14744) );
  INV_X1 U12710 ( .A(n14824), .ZN(n10018) );
  NAND2_X1 U12711 ( .A1(n15350), .A2(n10098), .ZN(n10012) );
  NAND2_X1 U12712 ( .A1(n14842), .A2(n6513), .ZN(n10011) );
  NAND2_X1 U12713 ( .A1(n10012), .A2(n10011), .ZN(n10013) );
  XNOR2_X1 U12714 ( .A(n10013), .B(n10123), .ZN(n10017) );
  NAND2_X1 U12715 ( .A1(n15350), .A2(n10108), .ZN(n10015) );
  NAND2_X1 U12716 ( .A1(n14842), .A2(n9996), .ZN(n10014) );
  NAND2_X1 U12717 ( .A1(n10015), .A2(n10014), .ZN(n10016) );
  NAND2_X1 U12718 ( .A1(n15342), .A2(n10098), .ZN(n10022) );
  NAND2_X1 U12719 ( .A1(n14841), .A2(n10108), .ZN(n10021) );
  NAND2_X1 U12720 ( .A1(n10022), .A2(n10021), .ZN(n10023) );
  XNOR2_X1 U12721 ( .A(n10023), .B(n10111), .ZN(n10025) );
  AND2_X1 U12722 ( .A1(n14841), .A2(n9996), .ZN(n10024) );
  AOI21_X1 U12723 ( .B1(n15342), .B2(n6513), .A(n10024), .ZN(n10026) );
  NAND2_X1 U12724 ( .A1(n10025), .A2(n10026), .ZN(n10030) );
  INV_X1 U12725 ( .A(n10025), .ZN(n10028) );
  INV_X1 U12726 ( .A(n10026), .ZN(n10027) );
  NAND2_X1 U12727 ( .A1(n10028), .A2(n10027), .ZN(n10029) );
  NAND2_X1 U12728 ( .A1(n10030), .A2(n10029), .ZN(n14754) );
  INV_X1 U12729 ( .A(n10030), .ZN(n10031) );
  NAND2_X1 U12730 ( .A1(n15339), .A2(n10098), .ZN(n10033) );
  NAND2_X1 U12731 ( .A1(n15140), .A2(n6513), .ZN(n10032) );
  NAND2_X1 U12732 ( .A1(n10033), .A2(n10032), .ZN(n10034) );
  XNOR2_X1 U12733 ( .A(n10034), .B(n10123), .ZN(n10035) );
  OAI22_X1 U12734 ( .A1(n15159), .A2(n9953), .B1(n15177), .B2(n10091), .ZN(
        n10036) );
  XNOR2_X1 U12735 ( .A(n10035), .B(n10036), .ZN(n14803) );
  INV_X1 U12736 ( .A(n10035), .ZN(n10038) );
  INV_X1 U12737 ( .A(n10036), .ZN(n10037) );
  NAND2_X1 U12738 ( .A1(n15330), .A2(n10098), .ZN(n10040) );
  NAND2_X1 U12739 ( .A1(n15116), .A2(n10108), .ZN(n10039) );
  NAND2_X1 U12740 ( .A1(n10040), .A2(n10039), .ZN(n10041) );
  XNOR2_X1 U12741 ( .A(n10041), .B(n10123), .ZN(n10043) );
  AND2_X1 U12742 ( .A1(n15116), .A2(n9996), .ZN(n10042) );
  AOI21_X1 U12743 ( .B1(n15330), .B2(n6513), .A(n10042), .ZN(n10044) );
  XNOR2_X1 U12744 ( .A(n10043), .B(n10044), .ZN(n14700) );
  INV_X1 U12745 ( .A(n10043), .ZN(n10045) );
  OAI22_X1 U12746 ( .A1(n15127), .A2(n9953), .B1(n15098), .B2(n10091), .ZN(
        n10049) );
  NAND2_X1 U12747 ( .A1(n15324), .A2(n10098), .ZN(n10047) );
  NAND2_X1 U12748 ( .A1(n15139), .A2(n6513), .ZN(n10046) );
  NAND2_X1 U12749 ( .A1(n10047), .A2(n10046), .ZN(n10048) );
  XNOR2_X1 U12750 ( .A(n10048), .B(n10123), .ZN(n10050) );
  XOR2_X1 U12751 ( .A(n10049), .B(n10050), .Z(n14771) );
  NAND2_X1 U12752 ( .A1(n15319), .A2(n10098), .ZN(n10052) );
  NAND2_X1 U12753 ( .A1(n15117), .A2(n6513), .ZN(n10051) );
  NAND2_X1 U12754 ( .A1(n10052), .A2(n10051), .ZN(n10053) );
  XNOR2_X1 U12755 ( .A(n10053), .B(n10123), .ZN(n10057) );
  NAND2_X1 U12756 ( .A1(n15319), .A2(n6513), .ZN(n10055) );
  NAND2_X1 U12757 ( .A1(n15117), .A2(n9996), .ZN(n10054) );
  NAND2_X1 U12758 ( .A1(n10055), .A2(n10054), .ZN(n10056) );
  NOR2_X1 U12759 ( .A1(n10057), .A2(n10056), .ZN(n10058) );
  AOI21_X1 U12760 ( .B1(n10057), .B2(n10056), .A(n10058), .ZN(n14717) );
  INV_X1 U12761 ( .A(n10058), .ZN(n14793) );
  OAI22_X1 U12762 ( .A1(n15090), .A2(n10059), .B1(n15099), .B2(n9953), .ZN(
        n10060) );
  XNOR2_X1 U12763 ( .A(n10060), .B(n10111), .ZN(n10063) );
  OR2_X1 U12764 ( .A1(n15090), .A2(n9953), .ZN(n10062) );
  NAND2_X1 U12765 ( .A1(n14840), .A2(n9996), .ZN(n10061) );
  AND2_X1 U12766 ( .A1(n10062), .A2(n10061), .ZN(n10064) );
  NAND2_X1 U12767 ( .A1(n10063), .A2(n10064), .ZN(n10068) );
  INV_X1 U12768 ( .A(n10063), .ZN(n10066) );
  INV_X1 U12769 ( .A(n10064), .ZN(n10065) );
  NAND2_X1 U12770 ( .A1(n10066), .A2(n10065), .ZN(n10067) );
  NAND2_X1 U12771 ( .A1(n10068), .A2(n10067), .ZN(n14792) );
  INV_X1 U12772 ( .A(n10068), .ZN(n14692) );
  NAND2_X1 U12773 ( .A1(n10073), .A2(n10098), .ZN(n10070) );
  NAND2_X1 U12774 ( .A1(n14839), .A2(n6513), .ZN(n10069) );
  NAND2_X1 U12775 ( .A1(n10070), .A2(n10069), .ZN(n10071) );
  XNOR2_X1 U12776 ( .A(n10071), .B(n10111), .ZN(n10074) );
  AND2_X1 U12777 ( .A1(n14839), .A2(n9893), .ZN(n10072) );
  AOI21_X1 U12778 ( .B1(n10073), .B2(n6513), .A(n10072), .ZN(n10075) );
  NAND2_X1 U12779 ( .A1(n10074), .A2(n10075), .ZN(n14762) );
  INV_X1 U12780 ( .A(n10074), .ZN(n10077) );
  INV_X1 U12781 ( .A(n10075), .ZN(n10076) );
  NAND2_X1 U12782 ( .A1(n10077), .A2(n10076), .ZN(n10078) );
  AND2_X1 U12783 ( .A1(n14762), .A2(n10078), .ZN(n14691) );
  NAND2_X1 U12784 ( .A1(n15031), .A2(n6513), .ZN(n10079) );
  XNOR2_X1 U12785 ( .A(n10080), .B(n10111), .ZN(n10082) );
  AND2_X1 U12786 ( .A1(n15031), .A2(n9893), .ZN(n10081) );
  AOI21_X1 U12787 ( .B1(n15053), .B2(n6513), .A(n10081), .ZN(n10083) );
  NAND2_X1 U12788 ( .A1(n10082), .A2(n10083), .ZN(n10087) );
  INV_X1 U12789 ( .A(n10082), .ZN(n10085) );
  INV_X1 U12790 ( .A(n10083), .ZN(n10084) );
  NAND2_X1 U12791 ( .A1(n10085), .A2(n10084), .ZN(n10086) );
  INV_X1 U12792 ( .A(n10087), .ZN(n14736) );
  NAND2_X1 U12793 ( .A1(n15030), .A2(n9886), .ZN(n10089) );
  NAND2_X1 U12794 ( .A1(n14838), .A2(n6513), .ZN(n10088) );
  NAND2_X1 U12795 ( .A1(n10089), .A2(n10088), .ZN(n10090) );
  XNOR2_X1 U12796 ( .A(n10090), .B(n10111), .ZN(n10093) );
  NOR2_X1 U12797 ( .A1(n14815), .A2(n10091), .ZN(n10092) );
  AOI21_X1 U12798 ( .B1(n15030), .B2(n6513), .A(n10092), .ZN(n10094) );
  INV_X1 U12799 ( .A(n10093), .ZN(n10096) );
  INV_X1 U12800 ( .A(n10094), .ZN(n10095) );
  NAND2_X1 U12801 ( .A1(n15289), .A2(n10098), .ZN(n10100) );
  NAND2_X1 U12802 ( .A1(n15032), .A2(n6513), .ZN(n10099) );
  NAND2_X1 U12803 ( .A1(n10100), .A2(n10099), .ZN(n10101) );
  XNOR2_X1 U12804 ( .A(n10101), .B(n10123), .ZN(n10105) );
  NAND2_X1 U12805 ( .A1(n15289), .A2(n6513), .ZN(n10103) );
  NAND2_X1 U12806 ( .A1(n15032), .A2(n9996), .ZN(n10102) );
  NAND2_X1 U12807 ( .A1(n10103), .A2(n10102), .ZN(n10104) );
  NOR2_X1 U12808 ( .A1(n10105), .A2(n10104), .ZN(n10106) );
  AOI21_X1 U12809 ( .B1(n10105), .B2(n10104), .A(n10106), .ZN(n14812) );
  INV_X1 U12810 ( .A(n10106), .ZN(n10107) );
  NAND2_X1 U12811 ( .A1(n15284), .A2(n9886), .ZN(n10110) );
  NAND2_X1 U12812 ( .A1(n14837), .A2(n10108), .ZN(n10109) );
  NAND2_X1 U12813 ( .A1(n10110), .A2(n10109), .ZN(n10112) );
  XNOR2_X1 U12814 ( .A(n10112), .B(n10111), .ZN(n10115) );
  INV_X1 U12815 ( .A(n10115), .ZN(n10117) );
  AND2_X1 U12816 ( .A1(n14837), .A2(n9996), .ZN(n10113) );
  AOI21_X1 U12817 ( .B1(n15284), .B2(n6513), .A(n10113), .ZN(n10114) );
  INV_X1 U12818 ( .A(n10114), .ZN(n10116) );
  AOI21_X1 U12819 ( .B1(n10117), .B2(n10116), .A(n10130), .ZN(n10150) );
  NAND2_X1 U12820 ( .A1(n10149), .A2(n10150), .ZN(n10148) );
  INV_X1 U12821 ( .A(n10148), .ZN(n10127) );
  INV_X1 U12822 ( .A(n10654), .ZN(n10119) );
  INV_X1 U12823 ( .A(n10118), .ZN(n10657) );
  NAND3_X1 U12824 ( .A1(n10119), .A2(n10657), .A3(n10655), .ZN(n10132) );
  OR2_X1 U12825 ( .A1(n15580), .A2(n10758), .ZN(n10120) );
  NAND2_X1 U12826 ( .A1(n14984), .A2(n6513), .ZN(n10122) );
  NAND2_X1 U12827 ( .A1(n14982), .A2(n9996), .ZN(n10121) );
  NAND2_X1 U12828 ( .A1(n10122), .A2(n10121), .ZN(n10124) );
  XNOR2_X1 U12829 ( .A(n10124), .B(n10123), .ZN(n10126) );
  AOI22_X1 U12830 ( .A1(n14984), .A2(n9886), .B1(n6513), .B2(n14982), .ZN(
        n10125) );
  XNOR2_X1 U12831 ( .A(n10126), .B(n10125), .ZN(n10131) );
  INV_X1 U12832 ( .A(n10131), .ZN(n10129) );
  INV_X1 U12833 ( .A(n10130), .ZN(n10128) );
  NAND3_X1 U12834 ( .A1(n10131), .A2(n10130), .A3(n14813), .ZN(n10145) );
  NAND2_X1 U12835 ( .A1(n10132), .A2(n10140), .ZN(n10134) );
  NAND2_X1 U12836 ( .A1(n10134), .A2(n10133), .ZN(n11029) );
  INV_X1 U12837 ( .A(n15508), .ZN(n14829) );
  INV_X1 U12838 ( .A(n10135), .ZN(n10136) );
  NAND2_X1 U12839 ( .A1(n15500), .A2(n15257), .ZN(n14825) );
  AOI22_X1 U12840 ( .A1(n14835), .A2(n14773), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10137) );
  OAI21_X1 U12841 ( .B1(n14816), .B2(n14825), .A(n10137), .ZN(n10143) );
  INV_X1 U12842 ( .A(n10138), .ZN(n10141) );
  NOR2_X1 U12843 ( .A1(n10139), .A2(n11828), .ZN(n10666) );
  AOI21_X2 U12844 ( .B1(n10141), .B2(n10666), .A(n15513), .ZN(n15503) );
  NOR2_X1 U12845 ( .A1(n14983), .A2(n15503), .ZN(n10142) );
  AOI211_X1 U12846 ( .C1(n12685), .C2(n14829), .A(n10143), .B(n10142), .ZN(
        n10144) );
  NAND2_X1 U12847 ( .A1(n10145), .A2(n10144), .ZN(n10146) );
  AOI21_X1 U12848 ( .B1(n10148), .B2(n8081), .A(n10146), .ZN(n10147) );
  NAND2_X1 U12849 ( .A1(n14982), .A2(n15256), .ZN(n10152) );
  NAND2_X1 U12850 ( .A1(n15032), .A2(n15257), .ZN(n10151) );
  NAND2_X1 U12851 ( .A1(n10152), .A2(n10151), .ZN(n10661) );
  OAI22_X1 U12852 ( .A1(n10668), .A2(n15508), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10153), .ZN(n10154) );
  AOI21_X1 U12853 ( .B1(n10661), .B2(n15500), .A(n10154), .ZN(n10155) );
  NAND2_X1 U12854 ( .A1(n10158), .A2(n10157), .ZN(P1_U3214) );
  NOR2_X1 U12855 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .ZN(n10159) );
  INV_X1 U12856 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10164) );
  INV_X1 U12857 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12559) );
  OR2_X1 U12858 ( .A1(n10185), .A2(n12559), .ZN(n10169) );
  NAND2_X1 U12859 ( .A1(n11779), .A2(n10301), .ZN(n10176) );
  INV_X1 U12860 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U12861 ( .A1(n10275), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n14176), 
        .B2(n10274), .ZN(n10175) );
  NAND2_X1 U12862 ( .A1(n10878), .A2(SI_0_), .ZN(n10179) );
  NAND2_X1 U12863 ( .A1(n10179), .A2(n10178), .ZN(n10181) );
  AND2_X1 U12864 ( .A1(n10180), .A2(n10181), .ZN(n14675) );
  MUX2_X1 U12865 ( .A(P2_IR_REG_0__SCAN_IN), .B(n14675), .S(n10184), .Z(n11400) );
  OR2_X1 U12866 ( .A1(n10184), .A2(n15609), .ZN(n10187) );
  OR2_X1 U12867 ( .A1(n10185), .A2(n10840), .ZN(n10186) );
  NAND2_X1 U12868 ( .A1(n10190), .A2(n10189), .ZN(n10223) );
  NAND2_X1 U12869 ( .A1(n10223), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10192) );
  INV_X1 U12870 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n10191) );
  XNOR2_X1 U12871 ( .A(n10192), .B(n10191), .ZN(n14117) );
  OR2_X1 U12872 ( .A1(n10184), .A2(n14117), .ZN(n10194) );
  OR2_X1 U12873 ( .A1(n10185), .A2(n10839), .ZN(n10193) );
  AND3_X2 U12874 ( .A1(n10195), .A2(n10194), .A3(n10193), .ZN(n11905) );
  NAND2_X1 U12875 ( .A1(n10859), .A2(n10251), .ZN(n10197) );
  NAND2_X1 U12876 ( .A1(n10199), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10196) );
  XNOR2_X1 U12877 ( .A(n10196), .B(P2_IR_REG_4__SCAN_IN), .ZN(n11253) );
  NAND2_X1 U12878 ( .A1(n10863), .A2(n10251), .ZN(n10206) );
  INV_X1 U12879 ( .A(n10199), .ZN(n10201) );
  INV_X1 U12880 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n10200) );
  NAND2_X1 U12881 ( .A1(n10201), .A2(n10200), .ZN(n10203) );
  NAND2_X1 U12882 ( .A1(n10203), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10202) );
  MUX2_X1 U12883 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10202), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n10204) );
  AOI22_X1 U12884 ( .A1(n10275), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n10274), 
        .B2(n11255), .ZN(n10205) );
  NAND2_X1 U12885 ( .A1(n10206), .A2(n10205), .ZN(n15813) );
  NAND2_X1 U12886 ( .A1(n10882), .A2(n10251), .ZN(n10213) );
  NAND2_X1 U12887 ( .A1(n10208), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10207) );
  MUX2_X1 U12888 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10207), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n10211) );
  INV_X1 U12889 ( .A(n10208), .ZN(n10210) );
  INV_X1 U12890 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n10209) );
  NAND2_X1 U12891 ( .A1(n10210), .A2(n10209), .ZN(n10217) );
  NAND2_X1 U12892 ( .A1(n10211), .A2(n10217), .ZN(n15646) );
  INV_X1 U12893 ( .A(n15646), .ZN(n11257) );
  AOI22_X1 U12894 ( .A1(n10275), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n10274), 
        .B2(n11257), .ZN(n10212) );
  NAND2_X1 U12895 ( .A1(n10213), .A2(n10212), .ZN(n15764) );
  INV_X1 U12896 ( .A(n15764), .ZN(n15824) );
  NAND2_X1 U12897 ( .A1(n10904), .A2(n10251), .ZN(n10216) );
  NAND2_X1 U12898 ( .A1(n10217), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10214) );
  XNOR2_X1 U12899 ( .A(n10214), .B(P2_IR_REG_7__SCAN_IN), .ZN(n11259) );
  AOI22_X1 U12900 ( .A1(n10275), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n10274), 
        .B2(n11259), .ZN(n10215) );
  NAND2_X1 U12901 ( .A1(n10911), .A2(n10251), .ZN(n10220) );
  OAI21_X1 U12902 ( .B1(n10217), .B2(P2_IR_REG_7__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n10218) );
  XNOR2_X1 U12903 ( .A(n10218), .B(P2_IR_REG_8__SCAN_IN), .ZN(n11262) );
  AOI22_X1 U12904 ( .A1(n10275), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n10274), 
        .B2(n11262), .ZN(n10219) );
  INV_X1 U12905 ( .A(n10223), .ZN(n10225) );
  NAND2_X1 U12906 ( .A1(n10225), .A2(n10224), .ZN(n10227) );
  NAND2_X1 U12907 ( .A1(n10227), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10226) );
  MUX2_X1 U12908 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10226), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n10228) );
  AOI22_X1 U12909 ( .A1(n10275), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n10274), 
        .B2(n11263), .ZN(n10229) );
  NAND2_X1 U12910 ( .A1(n10949), .A2(n10251), .ZN(n10235) );
  NAND2_X1 U12911 ( .A1(n10230), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10231) );
  MUX2_X1 U12912 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10231), .S(
        P2_IR_REG_10__SCAN_IN), .Z(n10233) );
  NAND2_X1 U12913 ( .A1(n10233), .A2(n10239), .ZN(n11232) );
  AOI22_X1 U12914 ( .A1(n10275), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n10274), 
        .B2(n15690), .ZN(n10234) );
  NAND2_X1 U12915 ( .A1(n10966), .A2(n10251), .ZN(n10238) );
  NAND2_X1 U12916 ( .A1(n10239), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10236) );
  XNOR2_X1 U12917 ( .A(n10236), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U12918 ( .A1(n10275), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n10274), 
        .B2(n11644), .ZN(n10237) );
  NAND2_X1 U12919 ( .A1(n11001), .A2(n10251), .ZN(n10242) );
  OR2_X1 U12920 ( .A1(n10239), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n10243) );
  NAND2_X1 U12921 ( .A1(n10243), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10240) );
  XNOR2_X1 U12922 ( .A(n10240), .B(P2_IR_REG_12__SCAN_IN), .ZN(n15701) );
  AOI22_X1 U12923 ( .A1(n10275), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n10274), 
        .B2(n15701), .ZN(n10241) );
  AND2_X2 U12924 ( .A1(n14457), .A2(n14458), .ZN(n14460) );
  NAND2_X1 U12925 ( .A1(n11046), .A2(n10251), .ZN(n10250) );
  INV_X1 U12926 ( .A(n10243), .ZN(n10245) );
  INV_X1 U12927 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n10244) );
  NAND2_X1 U12928 ( .A1(n10245), .A2(n10244), .ZN(n10247) );
  NAND2_X1 U12929 ( .A1(n10247), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10246) );
  MUX2_X1 U12930 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10246), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n10248) );
  AOI22_X1 U12931 ( .A1(n10275), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n10274), 
        .B2(n14149), .ZN(n10249) );
  NAND2_X1 U12932 ( .A1(n14460), .A2(n14645), .ZN(n14413) );
  NAND2_X1 U12933 ( .A1(n10253), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10252) );
  MUX2_X1 U12934 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10252), .S(
        P2_IR_REG_14__SCAN_IN), .Z(n10256) );
  INV_X1 U12935 ( .A(n10253), .ZN(n10255) );
  INV_X1 U12936 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n10254) );
  NAND2_X1 U12937 ( .A1(n10255), .A2(n10254), .ZN(n10263) );
  NAND2_X1 U12938 ( .A1(n10256), .A2(n10263), .ZN(n14152) );
  AOI22_X1 U12939 ( .A1(n10275), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n10274), 
        .B2(n15713), .ZN(n10257) );
  NAND2_X1 U12940 ( .A1(n10259), .A2(n10301), .ZN(n10262) );
  NAND2_X1 U12941 ( .A1(n10263), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10260) );
  XNOR2_X1 U12942 ( .A(n10260), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14155) );
  AOI22_X1 U12943 ( .A1(n10275), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n10274), 
        .B2(n14155), .ZN(n10261) );
  OAI21_X1 U12944 ( .B1(n10263), .B2(P2_IR_REG_15__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n10264) );
  XNOR2_X1 U12945 ( .A(n10264), .B(P2_IR_REG_16__SCAN_IN), .ZN(n15738) );
  AOI22_X1 U12946 ( .A1(n10275), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n15738), 
        .B2(n10274), .ZN(n10265) );
  NAND2_X1 U12947 ( .A1(n11446), .A2(n10301), .ZN(n10272) );
  NAND2_X1 U12948 ( .A1(n10266), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10268) );
  MUX2_X1 U12949 ( .A(n10268), .B(P2_IR_REG_31__SCAN_IN), .S(n10267), .Z(
        n10270) );
  NAND2_X1 U12950 ( .A1(n10270), .A2(n10269), .ZN(n14159) );
  INV_X1 U12951 ( .A(n14159), .ZN(n14167) );
  AOI22_X1 U12952 ( .A1(n10275), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n10274), 
        .B2(n14167), .ZN(n10271) );
  NAND2_X1 U12953 ( .A1(n10269), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10273) );
  XNOR2_X1 U12954 ( .A(n10273), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14170) );
  AOI22_X1 U12955 ( .A1(n10275), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n10274), 
        .B2(n14170), .ZN(n10276) );
  NAND2_X1 U12956 ( .A1(n11827), .A2(n10301), .ZN(n10279) );
  OR2_X1 U12957 ( .A1(n10185), .A2(n12359), .ZN(n10278) );
  OR2_X1 U12958 ( .A1(n10185), .A2(n12484), .ZN(n10280) );
  OR2_X2 U12959 ( .A1(n6563), .A2(n14539), .ZN(n14294) );
  NAND2_X1 U12960 ( .A1(n10283), .A2(n10282), .ZN(n10284) );
  OR2_X1 U12961 ( .A1(n6519), .A2(n11873), .ZN(n10286) );
  NAND2_X1 U12962 ( .A1(n12036), .A2(n10301), .ZN(n10288) );
  OR2_X1 U12963 ( .A1(n10185), .A2(n12039), .ZN(n10287) );
  OR2_X1 U12964 ( .A1(n10185), .A2(n12159), .ZN(n10289) );
  NAND2_X1 U12965 ( .A1(n12547), .A2(n10301), .ZN(n10291) );
  OR2_X1 U12966 ( .A1(n10185), .A2(n12549), .ZN(n10290) );
  OR2_X1 U12967 ( .A1(n10185), .A2(n14672), .ZN(n10293) );
  NAND2_X1 U12968 ( .A1(n14668), .A2(n10301), .ZN(n10296) );
  OR2_X1 U12969 ( .A1(n6519), .A2(n14670), .ZN(n10295) );
  NAND2_X1 U12970 ( .A1(n10297), .A2(n10301), .ZN(n10299) );
  OR2_X1 U12971 ( .A1(n10185), .A2(n14667), .ZN(n10298) );
  OR2_X1 U12972 ( .A1(n6519), .A2(n12697), .ZN(n10300) );
  INV_X1 U12973 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n14658) );
  OR2_X1 U12974 ( .A1(n6519), .A2(n14658), .ZN(n13981) );
  XNOR2_X2 U12975 ( .A(n10303), .B(P2_IR_REG_22__SCAN_IN), .ZN(n10315) );
  INV_X1 U12976 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n10304) );
  OAI21_X1 U12977 ( .B1(n10305), .B2(n10304), .A(P2_IR_REG_21__SCAN_IN), .ZN(
        n10308) );
  XNOR2_X2 U12978 ( .A(n10312), .B(n10311), .ZN(n14075) );
  NAND2_X1 U12979 ( .A1(n10313), .A2(n15767), .ZN(n12564) );
  NAND2_X1 U12980 ( .A1(n10315), .A2(n14066), .ZN(n10810) );
  INV_X1 U12981 ( .A(P2_B_REG_SCAN_IN), .ZN(n12479) );
  OR2_X1 U12982 ( .A1(n14669), .A2(n12479), .ZN(n10317) );
  NAND2_X1 U12983 ( .A1(n14449), .A2(n10317), .ZN(n14194) );
  NAND2_X1 U12984 ( .A1(n13968), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n10324) );
  NAND2_X1 U12985 ( .A1(n7281), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n10323) );
  NAND2_X1 U12986 ( .A1(n10373), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n10322) );
  NAND3_X1 U12987 ( .A1(n10324), .A2(n10323), .A3(n10322), .ZN(n14085) );
  INV_X1 U12988 ( .A(n14085), .ZN(n14023) );
  OR2_X1 U12989 ( .A1(n14194), .A2(n14023), .ZN(n14490) );
  NOR4_X1 U12990 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n10328) );
  NOR4_X1 U12991 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n10327) );
  NOR4_X1 U12992 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n10326) );
  NOR4_X1 U12993 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n10325) );
  NAND4_X1 U12994 ( .A1(n10328), .A2(n10327), .A3(n10326), .A4(n10325), .ZN(
        n10349) );
  NOR2_X1 U12995 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .ZN(
        n10332) );
  NOR4_X1 U12996 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n10331) );
  NOR4_X1 U12997 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n10330) );
  NOR4_X1 U12998 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n10329) );
  NAND4_X1 U12999 ( .A1(n10332), .A2(n10331), .A3(n10330), .A4(n10329), .ZN(
        n10348) );
  OAI21_X1 U13000 ( .B1(n10269), .B2(n10333), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n10334) );
  MUX2_X1 U13001 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10334), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n10336) );
  NAND2_X1 U13002 ( .A1(n10336), .A2(n10335), .ZN(n12548) );
  XNOR2_X1 U13003 ( .A(n12160), .B(P2_B_REG_SCAN_IN), .ZN(n10342) );
  NAND2_X1 U13004 ( .A1(n12548), .A2(n10342), .ZN(n10347) );
  NAND2_X1 U13005 ( .A1(n10335), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10343) );
  MUX2_X1 U13006 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10343), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n10345) );
  NAND2_X1 U13007 ( .A1(n10345), .A2(n10344), .ZN(n14674) );
  INV_X1 U13008 ( .A(n14674), .ZN(n10346) );
  INV_X1 U13009 ( .A(n10725), .ZN(n10808) );
  OAI211_X1 U13010 ( .C1(n10810), .C2(n14070), .A(n12037), .B(n10808), .ZN(
        n10817) );
  NAND2_X1 U13011 ( .A1(n11209), .A2(n11791), .ZN(n10823) );
  INV_X1 U13012 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15794) );
  NAND2_X1 U13013 ( .A1(n15784), .A2(n15794), .ZN(n10353) );
  NAND2_X1 U13014 ( .A1(n12548), .A2(n14674), .ZN(n10352) );
  NAND2_X1 U13015 ( .A1(n10353), .A2(n10352), .ZN(n15795) );
  NAND2_X1 U13016 ( .A1(n10823), .A2(n15795), .ZN(n10354) );
  NOR2_X1 U13017 ( .A1(n11273), .A2(n10354), .ZN(n10355) );
  NAND2_X1 U13018 ( .A1(n12160), .A2(n14674), .ZN(n10357) );
  INV_X1 U13019 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15791) );
  NAND2_X1 U13020 ( .A1(n15784), .A2(n15791), .ZN(n10356) );
  INV_X1 U13021 ( .A(n15792), .ZN(n10358) );
  INV_X1 U13022 ( .A(n14070), .ZN(n13966) );
  INV_X1 U13023 ( .A(n10404), .ZN(n10361) );
  INV_X1 U13024 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10495) );
  INV_X1 U13025 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10508) );
  INV_X1 U13026 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10520) );
  INV_X1 U13027 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10364) );
  NAND2_X1 U13028 ( .A1(n10523), .A2(n10364), .ZN(n10365) );
  AND2_X1 U13029 ( .A1(n10529), .A2(n10365), .ZN(n14313) );
  NAND2_X1 U13030 ( .A1(n14313), .A2(n10720), .ZN(n10372) );
  INV_X1 U13031 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n10369) );
  NAND2_X1 U13032 ( .A1(n10373), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n10368) );
  NAND2_X1 U13033 ( .A1(n13968), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n10367) );
  OAI211_X1 U13034 ( .C1(n10369), .C2(n6522), .A(n10368), .B(n10367), .ZN(
        n10370) );
  INV_X1 U13035 ( .A(n10370), .ZN(n10371) );
  INV_X1 U13036 ( .A(n14544), .ZN(n14316) );
  NAND2_X1 U13037 ( .A1(n6521), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10374) );
  NAND2_X1 U13038 ( .A1(n6512), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10377) );
  NAND2_X1 U13039 ( .A1(n10373), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n10376) );
  AND2_X1 U13040 ( .A1(n10586), .A2(n11400), .ZN(n11338) );
  NAND2_X1 U13041 ( .A1(n11972), .A2(n11338), .ZN(n10388) );
  INV_X1 U13042 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10380) );
  OR2_X1 U13043 ( .A1(n10643), .A2(n10380), .ZN(n10385) );
  NAND2_X1 U13044 ( .A1(n13969), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10383) );
  INV_X1 U13045 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15804) );
  NAND2_X1 U13046 ( .A1(n11275), .A2(n15800), .ZN(n10386) );
  NAND2_X1 U13047 ( .A1(n10389), .A2(n13813), .ZN(n10589) );
  NAND2_X1 U13048 ( .A1(n10389), .A2(n15800), .ZN(n10390) );
  NAND2_X1 U13049 ( .A1(n13968), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10395) );
  INV_X1 U13050 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10391) );
  NAND2_X1 U13051 ( .A1(n10720), .A2(n10391), .ZN(n10394) );
  NAND2_X1 U13052 ( .A1(n13969), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10393) );
  NAND2_X1 U13053 ( .A1(n10373), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n10392) );
  XNOR2_X1 U13054 ( .A(n14101), .B(n11905), .ZN(n11370) );
  INV_X1 U13055 ( .A(n14101), .ZN(n11462) );
  NAND2_X1 U13056 ( .A1(n11462), .A2(n11905), .ZN(n10396) );
  NAND2_X1 U13057 ( .A1(n11369), .A2(n10396), .ZN(n12009) );
  NAND2_X1 U13058 ( .A1(n13968), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10401) );
  OAI21_X1 U13059 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n10404), .ZN(n10397) );
  INV_X1 U13060 ( .A(n10397), .ZN(n12014) );
  NAND2_X1 U13061 ( .A1(n10720), .A2(n12014), .ZN(n10400) );
  NAND2_X1 U13062 ( .A1(n13969), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10399) );
  NAND2_X1 U13063 ( .A1(n10373), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n10398) );
  NAND4_X1 U13064 ( .A1(n10401), .A2(n10400), .A3(n10399), .A4(n10398), .ZN(
        n14100) );
  XNOR2_X1 U13065 ( .A(n14100), .B(n15806), .ZN(n12008) );
  NAND2_X1 U13066 ( .A1(n12009), .A2(n12008), .ZN(n12011) );
  INV_X1 U13067 ( .A(n14100), .ZN(n13842) );
  NAND2_X1 U13068 ( .A1(n13842), .A2(n15806), .ZN(n10402) );
  NAND2_X1 U13069 ( .A1(n12011), .A2(n10402), .ZN(n11784) );
  NAND2_X1 U13070 ( .A1(n13968), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10409) );
  INV_X1 U13071 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10403) );
  NAND2_X1 U13072 ( .A1(n10404), .A2(n10403), .ZN(n10405) );
  AND2_X1 U13073 ( .A1(n10414), .A2(n10405), .ZN(n11801) );
  NAND2_X1 U13074 ( .A1(n10720), .A2(n11801), .ZN(n10408) );
  NAND2_X1 U13075 ( .A1(n13970), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n10407) );
  NAND2_X1 U13076 ( .A1(n7281), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10406) );
  NAND4_X1 U13077 ( .A1(n10409), .A2(n10408), .A3(n10407), .A4(n10406), .ZN(
        n14099) );
  NAND2_X1 U13078 ( .A1(n15813), .A2(n14099), .ZN(n10410) );
  NAND2_X1 U13079 ( .A1(n11784), .A2(n10410), .ZN(n10412) );
  INV_X1 U13080 ( .A(n14099), .ZN(n13849) );
  INV_X1 U13081 ( .A(n15813), .ZN(n13850) );
  NAND2_X1 U13082 ( .A1(n13849), .A2(n13850), .ZN(n10411) );
  NAND2_X1 U13083 ( .A1(n13970), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n10419) );
  NAND2_X1 U13084 ( .A1(n13968), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10418) );
  INV_X1 U13085 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10413) );
  NAND2_X1 U13086 ( .A1(n10414), .A2(n10413), .ZN(n10415) );
  AND2_X1 U13087 ( .A1(n10422), .A2(n10415), .ZN(n15761) );
  NAND2_X1 U13088 ( .A1(n10720), .A2(n15761), .ZN(n10417) );
  NAND2_X1 U13089 ( .A1(n7281), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10416) );
  NAND2_X1 U13090 ( .A1(n15766), .A2(n15765), .ZN(n10421) );
  INV_X1 U13091 ( .A(n13855), .ZN(n14098) );
  OR2_X1 U13092 ( .A1(n15764), .A2(n14098), .ZN(n10420) );
  NAND2_X1 U13093 ( .A1(n10421), .A2(n10420), .ZN(n11935) );
  NAND2_X1 U13094 ( .A1(n13968), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10427) );
  NAND2_X1 U13095 ( .A1(n10373), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n10426) );
  NAND2_X1 U13096 ( .A1(n10422), .A2(n12308), .ZN(n10423) );
  AND2_X1 U13097 ( .A1(n10431), .A2(n10423), .ZN(n11937) );
  NAND2_X1 U13098 ( .A1(n10720), .A2(n11937), .ZN(n10425) );
  NAND2_X1 U13099 ( .A1(n7281), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10424) );
  INV_X1 U13100 ( .A(n13859), .ZN(n14097) );
  OR2_X1 U13101 ( .A1(n13858), .A2(n14097), .ZN(n10428) );
  NAND2_X1 U13102 ( .A1(n13968), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10436) );
  NAND2_X1 U13103 ( .A1(n10431), .A2(n10430), .ZN(n10432) );
  NAND2_X1 U13104 ( .A1(n10720), .A2(n8087), .ZN(n10435) );
  NAND2_X1 U13105 ( .A1(n13970), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n10434) );
  NAND2_X1 U13106 ( .A1(n7281), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10433) );
  NAND4_X1 U13107 ( .A1(n10436), .A2(n10435), .A3(n10434), .A4(n10433), .ZN(
        n14096) );
  NAND2_X1 U13108 ( .A1(n13970), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n10443) );
  NAND2_X1 U13109 ( .A1(n13968), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n10442) );
  NAND2_X1 U13110 ( .A1(n10438), .A2(n10437), .ZN(n10439) );
  AND2_X1 U13111 ( .A1(n10447), .A2(n10439), .ZN(n12591) );
  NAND2_X1 U13112 ( .A1(n10720), .A2(n12591), .ZN(n10441) );
  NAND2_X1 U13113 ( .A1(n7281), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10440) );
  OR2_X1 U13114 ( .A1(n14044), .A2(n10597), .ZN(n10444) );
  NAND2_X1 U13115 ( .A1(n13870), .A2(n8009), .ZN(n10445) );
  NAND2_X1 U13116 ( .A1(n7205), .A2(n14096), .ZN(n12070) );
  NAND2_X1 U13117 ( .A1(n13968), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10452) );
  INV_X1 U13118 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10446) );
  NAND2_X1 U13119 ( .A1(n10447), .A2(n10446), .ZN(n10448) );
  AND2_X1 U13120 ( .A1(n10457), .A2(n10448), .ZN(n12230) );
  NAND2_X1 U13121 ( .A1(n10720), .A2(n12230), .ZN(n10451) );
  NAND2_X1 U13122 ( .A1(n13970), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n10450) );
  NAND2_X1 U13123 ( .A1(n7281), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10449) );
  NAND4_X1 U13124 ( .A1(n10452), .A2(n10451), .A3(n10450), .A4(n10449), .ZN(
        n14095) );
  INV_X1 U13125 ( .A(n14047), .ZN(n10453) );
  AND2_X1 U13126 ( .A1(n12026), .A2(n10453), .ZN(n10454) );
  OR2_X1 U13127 ( .A1(n14605), .A2(n14095), .ZN(n10455) );
  NAND2_X1 U13128 ( .A1(n13968), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10462) );
  NAND2_X1 U13129 ( .A1(n10457), .A2(n10456), .ZN(n10458) );
  AND2_X1 U13130 ( .A1(n10466), .A2(n10458), .ZN(n14484) );
  NAND2_X1 U13131 ( .A1(n10720), .A2(n14484), .ZN(n10461) );
  NAND2_X1 U13132 ( .A1(n7281), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10460) );
  NAND2_X1 U13133 ( .A1(n13970), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n10459) );
  NAND4_X1 U13134 ( .A1(n10462), .A2(n10461), .A3(n10460), .A4(n10459), .ZN(
        n14450) );
  XNOR2_X1 U13135 ( .A(n14483), .B(n14450), .ZN(n14470) );
  NAND2_X1 U13136 ( .A1(n14483), .A2(n14450), .ZN(n10464) );
  NAND2_X1 U13137 ( .A1(n13968), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10471) );
  INV_X1 U13138 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10465) );
  NAND2_X1 U13139 ( .A1(n10466), .A2(n10465), .ZN(n10467) );
  AND2_X1 U13140 ( .A1(n10475), .A2(n10467), .ZN(n13680) );
  NAND2_X1 U13141 ( .A1(n10720), .A2(n13680), .ZN(n10470) );
  NAND2_X1 U13142 ( .A1(n13970), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n10469) );
  NAND2_X1 U13143 ( .A1(n7281), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n10468) );
  NAND4_X1 U13144 ( .A1(n10471), .A2(n10470), .A3(n10469), .A4(n10468), .ZN(
        n14094) );
  OR2_X1 U13145 ( .A1(n14588), .A2(n14094), .ZN(n10472) );
  NAND2_X1 U13146 ( .A1(n14440), .A2(n10472), .ZN(n10474) );
  NAND2_X1 U13147 ( .A1(n14588), .A2(n14094), .ZN(n10473) );
  NAND2_X1 U13148 ( .A1(n10474), .A2(n10473), .ZN(n14428) );
  NAND2_X1 U13149 ( .A1(n13968), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10480) );
  NAND2_X1 U13150 ( .A1(n10475), .A2(n13741), .ZN(n10476) );
  AND2_X1 U13151 ( .A1(n10483), .A2(n10476), .ZN(n14433) );
  NAND2_X1 U13152 ( .A1(n10720), .A2(n14433), .ZN(n10479) );
  NAND2_X1 U13153 ( .A1(n13970), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n10478) );
  NAND2_X1 U13154 ( .A1(n7281), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10477) );
  NAND4_X1 U13155 ( .A1(n10480), .A2(n10479), .A3(n10478), .A4(n10477), .ZN(
        n14448) );
  AND2_X1 U13156 ( .A1(n14432), .A2(n14448), .ZN(n10481) );
  NAND2_X1 U13157 ( .A1(n6512), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n10488) );
  NAND2_X1 U13158 ( .A1(n10483), .A2(n10482), .ZN(n10484) );
  AND2_X1 U13159 ( .A1(n10491), .A2(n10484), .ZN(n14415) );
  NAND2_X1 U13160 ( .A1(n10720), .A2(n14415), .ZN(n10487) );
  NAND2_X1 U13161 ( .A1(n13970), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n10486) );
  NAND2_X1 U13162 ( .A1(n7281), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n10485) );
  NAND4_X1 U13163 ( .A1(n10488), .A2(n10487), .A3(n10486), .A4(n10485), .ZN(
        n14397) );
  NOR2_X1 U13164 ( .A1(n14580), .A2(n14397), .ZN(n14034) );
  INV_X1 U13165 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n14389) );
  NAND2_X1 U13166 ( .A1(n13970), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n10490) );
  NAND2_X1 U13167 ( .A1(n6512), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n10489) );
  AND2_X1 U13168 ( .A1(n10490), .A2(n10489), .ZN(n10494) );
  NAND2_X1 U13169 ( .A1(n10491), .A2(n6971), .ZN(n10492) );
  NAND2_X1 U13170 ( .A1(n10496), .A2(n10492), .ZN(n14388) );
  OR2_X1 U13171 ( .A1(n14388), .A2(n7879), .ZN(n10493) );
  OAI211_X1 U13172 ( .C1(n6522), .C2(n14389), .A(n10494), .B(n10493), .ZN(
        n14093) );
  XNOR2_X1 U13173 ( .A(n14393), .B(n14093), .ZN(n14394) );
  NAND2_X1 U13174 ( .A1(n10496), .A2(n10495), .ZN(n10497) );
  NAND2_X1 U13175 ( .A1(n10500), .A2(n10497), .ZN(n14379) );
  AOI22_X1 U13176 ( .A1(n7281), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n13968), 
        .B2(P2_REG1_REG_16__SCAN_IN), .ZN(n10499) );
  NAND2_X1 U13177 ( .A1(n13970), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n10498) );
  OAI211_X1 U13178 ( .C1(n14379), .C2(n7879), .A(n10499), .B(n10498), .ZN(
        n14398) );
  AND2_X1 U13179 ( .A1(n14568), .A2(n14398), .ZN(n14356) );
  NAND2_X1 U13180 ( .A1(n10500), .A2(n6972), .ZN(n10501) );
  NAND2_X1 U13181 ( .A1(n10509), .A2(n10501), .ZN(n14365) );
  OR2_X1 U13182 ( .A1(n14365), .A2(n7879), .ZN(n10504) );
  AOI22_X1 U13183 ( .A1(n13970), .A2(P2_REG0_REG_17__SCAN_IN), .B1(n13968), 
        .B2(P2_REG1_REG_17__SCAN_IN), .ZN(n10503) );
  NAND2_X1 U13184 ( .A1(n7281), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n10502) );
  XNOR2_X1 U13185 ( .A(n14364), .B(n14376), .ZN(n14051) );
  OR2_X1 U13186 ( .A1(n14393), .A2(n14093), .ZN(n14355) );
  OAI22_X1 U13187 ( .A1(n14355), .A2(n14356), .B1(n14398), .B2(n14568), .ZN(
        n10505) );
  INV_X1 U13188 ( .A(n10505), .ZN(n10506) );
  NAND2_X1 U13189 ( .A1(n14364), .A2(n14339), .ZN(n10507) );
  NAND2_X1 U13190 ( .A1(n10509), .A2(n10508), .ZN(n10510) );
  NAND2_X1 U13191 ( .A1(n10521), .A2(n10510), .ZN(n14344) );
  OR2_X1 U13192 ( .A1(n14344), .A2(n7879), .ZN(n10515) );
  INV_X1 U13193 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n14345) );
  NAND2_X1 U13194 ( .A1(n13970), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n10512) );
  NAND2_X1 U13195 ( .A1(n6512), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n10511) );
  OAI211_X1 U13196 ( .C1(n14345), .C2(n6522), .A(n10512), .B(n10511), .ZN(
        n10513) );
  INV_X1 U13197 ( .A(n10513), .ZN(n10514) );
  NAND2_X1 U13198 ( .A1(n10515), .A2(n10514), .ZN(n14092) );
  NAND2_X1 U13199 ( .A1(n10521), .A2(n10520), .ZN(n10522) );
  NAND2_X1 U13200 ( .A1(n10523), .A2(n10522), .ZN(n14326) );
  INV_X1 U13201 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n14327) );
  NAND2_X1 U13202 ( .A1(n13968), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n10525) );
  NAND2_X1 U13203 ( .A1(n10373), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n10524) );
  OAI211_X1 U13204 ( .C1(n14327), .C2(n6522), .A(n10525), .B(n10524), .ZN(
        n10526) );
  INV_X1 U13205 ( .A(n10526), .ZN(n10527) );
  OAI21_X1 U13206 ( .B1(n14326), .B2(n7879), .A(n10527), .ZN(n14340) );
  NAND2_X1 U13207 ( .A1(n14329), .A2(n14340), .ZN(n10528) );
  INV_X1 U13208 ( .A(n14340), .ZN(n13907) );
  XNOR2_X1 U13209 ( .A(n14544), .B(n13909), .ZN(n14309) );
  INV_X1 U13210 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13672) );
  NAND2_X1 U13211 ( .A1(n10529), .A2(n13672), .ZN(n10530) );
  NAND2_X1 U13212 ( .A1(n10538), .A2(n10530), .ZN(n14296) );
  OR2_X1 U13213 ( .A1(n14296), .A2(n7879), .ZN(n10536) );
  INV_X1 U13214 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n10533) );
  NAND2_X1 U13215 ( .A1(n10373), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n10532) );
  NAND2_X1 U13216 ( .A1(n6512), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n10531) );
  OAI211_X1 U13217 ( .C1(n10533), .C2(n6522), .A(n10532), .B(n10531), .ZN(
        n10534) );
  INV_X1 U13218 ( .A(n10534), .ZN(n10535) );
  NAND2_X1 U13219 ( .A1(n10536), .A2(n10535), .ZN(n14091) );
  AND2_X1 U13220 ( .A1(n14539), .A2(n14091), .ZN(n14032) );
  OR2_X1 U13221 ( .A1(n14539), .A2(n14091), .ZN(n14031) );
  INV_X1 U13222 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10537) );
  NAND2_X1 U13223 ( .A1(n10538), .A2(n10537), .ZN(n10539) );
  AND2_X1 U13224 ( .A1(n10546), .A2(n10539), .ZN(n14285) );
  NAND2_X1 U13225 ( .A1(n14285), .A2(n10720), .ZN(n10545) );
  INV_X1 U13226 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n10542) );
  NAND2_X1 U13227 ( .A1(n6512), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n10541) );
  NAND2_X1 U13228 ( .A1(n13970), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n10540) );
  OAI211_X1 U13229 ( .C1(n10542), .C2(n6522), .A(n10541), .B(n10540), .ZN(
        n10543) );
  INV_X1 U13230 ( .A(n10543), .ZN(n10544) );
  XNOR2_X1 U13231 ( .A(n14284), .B(n14263), .ZN(n14282) );
  INV_X1 U13232 ( .A(n14263), .ZN(n13671) );
  INV_X1 U13233 ( .A(n14284), .ZN(n14626) );
  INV_X1 U13234 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n12504) );
  NAND2_X1 U13235 ( .A1(n10546), .A2(n12504), .ZN(n10547) );
  NAND2_X1 U13236 ( .A1(n10563), .A2(n10547), .ZN(n14261) );
  INV_X1 U13237 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n14272) );
  NAND2_X1 U13238 ( .A1(n13970), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n10549) );
  NAND2_X1 U13239 ( .A1(n13968), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n10548) );
  OAI211_X1 U13240 ( .C1(n14272), .C2(n6522), .A(n10549), .B(n10548), .ZN(
        n10550) );
  INV_X1 U13241 ( .A(n10550), .ZN(n10551) );
  AND2_X1 U13242 ( .A1(n14528), .A2(n14090), .ZN(n14029) );
  NOR2_X1 U13243 ( .A1(n14528), .A2(n14090), .ZN(n14030) );
  XNOR2_X1 U13244 ( .A(n10563), .B(P2_REG3_REG_24__SCAN_IN), .ZN(n14254) );
  NAND2_X1 U13245 ( .A1(n14254), .A2(n10720), .ZN(n10558) );
  INV_X1 U13246 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n10555) );
  NAND2_X1 U13247 ( .A1(n10373), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n10554) );
  NAND2_X1 U13248 ( .A1(n13968), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n10553) );
  OAI211_X1 U13249 ( .C1(n10555), .C2(n6522), .A(n10554), .B(n10553), .ZN(
        n10556) );
  INV_X1 U13250 ( .A(n10556), .ZN(n10557) );
  XNOR2_X1 U13251 ( .A(n14522), .B(n14262), .ZN(n14249) );
  NAND2_X1 U13252 ( .A1(n14522), .A2(n10559), .ZN(n10560) );
  INV_X1 U13253 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13719) );
  INV_X1 U13254 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10561) );
  OAI21_X1 U13255 ( .B1(n10563), .B2(n13719), .A(n10561), .ZN(n10564) );
  NAND2_X1 U13256 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n10562) );
  NAND2_X1 U13257 ( .A1(n14232), .A2(n10720), .ZN(n10570) );
  INV_X1 U13258 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n10567) );
  NAND2_X1 U13259 ( .A1(n10373), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n10566) );
  NAND2_X1 U13260 ( .A1(n13968), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n10565) );
  OAI211_X1 U13261 ( .C1(n10567), .C2(n6522), .A(n10566), .B(n10565), .ZN(
        n10568) );
  INV_X1 U13262 ( .A(n10568), .ZN(n10569) );
  NAND2_X1 U13263 ( .A1(n14234), .A2(n13718), .ZN(n10571) );
  INV_X1 U13264 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13790) );
  NAND2_X1 U13265 ( .A1(n10573), .A2(n13790), .ZN(n10574) );
  INV_X1 U13266 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n14218) );
  NAND2_X1 U13267 ( .A1(n13970), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n10576) );
  NAND2_X1 U13268 ( .A1(n6512), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n10575) );
  OAI211_X1 U13269 ( .C1(n14218), .C2(n6522), .A(n10576), .B(n10575), .ZN(
        n10577) );
  INV_X1 U13270 ( .A(n10577), .ZN(n10578) );
  XNOR2_X1 U13271 ( .A(n10639), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n14209) );
  INV_X1 U13272 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n10582) );
  NAND2_X1 U13273 ( .A1(n13970), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n10581) );
  NAND2_X1 U13274 ( .A1(n6512), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n10580) );
  OAI211_X1 U13275 ( .C1(n10582), .C2(n6522), .A(n10581), .B(n10580), .ZN(
        n10583) );
  NAND2_X1 U13276 ( .A1(n13992), .A2(n13993), .ZN(n10711) );
  OR2_X1 U13277 ( .A1(n13992), .A2(n13993), .ZN(n10584) );
  XNOR2_X1 U13278 ( .A(n10709), .B(n14058), .ZN(n14214) );
  NAND2_X2 U13279 ( .A1(n14066), .A2(n14075), .ZN(n14068) );
  XNOR2_X1 U13280 ( .A(n14068), .B(n10315), .ZN(n10585) );
  INV_X1 U13281 ( .A(n11400), .ZN(n13820) );
  NOR2_X1 U13282 ( .A1(n13819), .A2(n13820), .ZN(n11339) );
  NAND2_X1 U13283 ( .A1(n13816), .A2(n10379), .ZN(n11965) );
  INV_X1 U13284 ( .A(n10587), .ZN(n14036) );
  NAND2_X1 U13285 ( .A1(n10588), .A2(n14036), .ZN(n11968) );
  NAND2_X1 U13286 ( .A1(n11968), .A2(n10589), .ZN(n11372) );
  INV_X1 U13287 ( .A(n11370), .ZN(n14037) );
  NAND2_X1 U13288 ( .A1(n11372), .A2(n14037), .ZN(n11371) );
  NAND2_X1 U13289 ( .A1(n11462), .A2(n7648), .ZN(n10590) );
  NAND2_X1 U13290 ( .A1(n11371), .A2(n10590), .ZN(n12017) );
  INV_X1 U13291 ( .A(n12008), .ZN(n14038) );
  NAND2_X1 U13292 ( .A1(n13842), .A2(n13843), .ZN(n10591) );
  AND2_X1 U13293 ( .A1(n13849), .A2(n15813), .ZN(n11786) );
  NAND2_X1 U13294 ( .A1(n13850), .A2(n14099), .ZN(n11785) );
  NAND2_X1 U13295 ( .A1(n15764), .A2(n13855), .ZN(n10593) );
  AND2_X1 U13296 ( .A1(n13858), .A2(n13859), .ZN(n10594) );
  INV_X1 U13297 ( .A(n14096), .ZN(n13865) );
  OR2_X1 U13298 ( .A1(n7205), .A2(n13865), .ZN(n10595) );
  NAND2_X1 U13299 ( .A1(n10596), .A2(n10595), .ZN(n12075) );
  NAND2_X1 U13300 ( .A1(n12075), .A2(n10597), .ZN(n10599) );
  OR2_X1 U13301 ( .A1(n13870), .A2(n13868), .ZN(n10598) );
  INV_X1 U13302 ( .A(n14095), .ZN(n14473) );
  OR2_X1 U13303 ( .A1(n14605), .A2(n14473), .ZN(n10600) );
  XNOR2_X1 U13304 ( .A(n14432), .B(n14448), .ZN(n14429) );
  INV_X1 U13305 ( .A(n14450), .ZN(n13878) );
  NAND2_X1 U13306 ( .A1(n14483), .A2(n13878), .ZN(n14422) );
  NAND2_X1 U13307 ( .A1(n14422), .A2(n14094), .ZN(n10602) );
  NOR2_X1 U13308 ( .A1(n14450), .A2(n14094), .ZN(n10601) );
  AOI22_X1 U13309 ( .A1(n14588), .A2(n10602), .B1(n10601), .B2(n14483), .ZN(
        n10603) );
  AND2_X1 U13310 ( .A1(n14429), .A2(n10603), .ZN(n10604) );
  INV_X1 U13311 ( .A(n14580), .ZN(n14418) );
  INV_X1 U13312 ( .A(n14448), .ZN(n14411) );
  NOR2_X1 U13313 ( .A1(n14432), .A2(n14411), .ZN(n14406) );
  AOI21_X1 U13314 ( .B1(n14418), .B2(n14397), .A(n14406), .ZN(n10606) );
  INV_X1 U13315 ( .A(n10604), .ZN(n14404) );
  OR2_X1 U13316 ( .A1(n14588), .A2(n14475), .ZN(n14423) );
  OR2_X1 U13317 ( .A1(n14483), .A2(n13878), .ZN(n10605) );
  AND2_X1 U13318 ( .A1(n14423), .A2(n10605), .ZN(n14405) );
  INV_X1 U13319 ( .A(n14397), .ZN(n14427) );
  NAND2_X1 U13320 ( .A1(n14580), .A2(n14427), .ZN(n10609) );
  INV_X1 U13321 ( .A(n14093), .ZN(n14412) );
  AND2_X1 U13322 ( .A1(n14393), .A2(n14412), .ZN(n10611) );
  XNOR2_X1 U13323 ( .A(n14568), .B(n14398), .ZN(n14374) );
  INV_X1 U13324 ( .A(n14398), .ZN(n14361) );
  OR2_X1 U13325 ( .A1(n14568), .A2(n14361), .ZN(n10612) );
  INV_X1 U13326 ( .A(n14051), .ZN(n14359) );
  OR2_X1 U13327 ( .A1(n14364), .A2(n14376), .ZN(n10613) );
  NAND2_X1 U13328 ( .A1(n14351), .A2(n10517), .ZN(n10614) );
  OR2_X1 U13329 ( .A1(n14351), .A2(n10517), .ZN(n10615) );
  NAND2_X1 U13330 ( .A1(n14329), .A2(n13907), .ZN(n10616) );
  NAND2_X1 U13331 ( .A1(n14320), .A2(n10616), .ZN(n10618) );
  OR2_X1 U13332 ( .A1(n14329), .A2(n13907), .ZN(n10617) );
  NOR2_X1 U13333 ( .A1(n14544), .A2(n13909), .ZN(n10619) );
  NAND2_X1 U13334 ( .A1(n14544), .A2(n13909), .ZN(n10620) );
  INV_X1 U13335 ( .A(n14091), .ZN(n13729) );
  AND2_X1 U13336 ( .A1(n14539), .A2(n13729), .ZN(n10621) );
  NAND2_X1 U13337 ( .A1(n14528), .A2(n13717), .ZN(n14242) );
  NAND2_X1 U13338 ( .A1(n14522), .A2(n14262), .ZN(n10622) );
  AND2_X1 U13339 ( .A1(n14242), .A2(n10622), .ZN(n10627) );
  INV_X1 U13340 ( .A(n10622), .ZN(n10623) );
  INV_X1 U13341 ( .A(n14249), .ZN(n14244) );
  XNOR2_X1 U13342 ( .A(n14234), .B(n13718), .ZN(n14235) );
  AND2_X1 U13343 ( .A1(n14517), .A2(n13718), .ZN(n10625) );
  INV_X1 U13344 ( .A(n10629), .ZN(n10626) );
  AOI21_X1 U13345 ( .B1(n14234), .B2(n14089), .A(n14088), .ZN(n10632) );
  NAND2_X1 U13346 ( .A1(n14088), .A2(n14089), .ZN(n10631) );
  OAI22_X1 U13347 ( .A1(n10632), .A2(n14217), .B1(n14517), .B2(n10631), .ZN(
        n10633) );
  NOR2_X1 U13348 ( .A1(n14058), .A2(n10633), .ZN(n10634) );
  NAND2_X1 U13349 ( .A1(n10315), .A2(n14176), .ZN(n10636) );
  INV_X1 U13350 ( .A(n14075), .ZN(n14065) );
  NAND2_X1 U13351 ( .A1(n14066), .A2(n14065), .ZN(n10635) );
  INV_X1 U13352 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13628) );
  INV_X1 U13353 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10637) );
  OAI21_X1 U13354 ( .B1(n10639), .B2(n13628), .A(n10637), .ZN(n10640) );
  NAND2_X1 U13355 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n10638) );
  NAND2_X1 U13356 ( .A1(n14203), .A2(n10720), .ZN(n10647) );
  INV_X1 U13357 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n10644) );
  NAND2_X1 U13358 ( .A1(n13970), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n10642) );
  NAND2_X1 U13359 ( .A1(n7281), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n10641) );
  OAI211_X1 U13360 ( .C1(n10644), .C2(n10643), .A(n10642), .B(n10641), .ZN(
        n10645) );
  INV_X1 U13361 ( .A(n10645), .ZN(n10646) );
  INV_X1 U13362 ( .A(n10314), .ZN(n10648) );
  OAI22_X1 U13363 ( .A1(n14196), .A2(n14474), .B1(n10649), .B2(n14472), .ZN(
        n13631) );
  INV_X1 U13364 ( .A(n10651), .ZN(n14215) );
  INV_X1 U13365 ( .A(n10722), .ZN(n10652) );
  OAI211_X1 U13366 ( .C1(n14511), .C2(n14215), .A(n10652), .B(n15767), .ZN(
        n14208) );
  OAI211_X1 U13367 ( .C1(n14214), .C2(n15817), .A(n14211), .B(n14208), .ZN(
        n14510) );
  NAND4_X1 U13368 ( .A1(n10657), .A2(n10656), .A3(n10655), .A4(n10654), .ZN(
        n11390) );
  NOR2_X1 U13369 ( .A1(n15262), .A2(n10658), .ZN(n15521) );
  AOI21_X1 U13370 ( .B1(n15552), .B2(n15232), .A(n15521), .ZN(n15169) );
  NOR2_X1 U13371 ( .A1(n15287), .A2(n15169), .ZN(n10674) );
  XNOR2_X1 U13372 ( .A(n10660), .B(n10659), .ZN(n10662) );
  NAND2_X1 U13373 ( .A1(n15284), .A2(n15015), .ZN(n10663) );
  NAND2_X1 U13374 ( .A1(n10663), .A2(n15555), .ZN(n10664) );
  NOR2_X1 U13375 ( .A1(n10665), .A2(n10664), .ZN(n15283) );
  OR2_X1 U13376 ( .A1(n11390), .A2(n15199), .ZN(n15067) );
  INV_X1 U13377 ( .A(n15067), .ZN(n15254) );
  INV_X1 U13378 ( .A(n10666), .ZN(n10667) );
  OR2_X2 U13379 ( .A1(n15262), .A2(n10667), .ZN(n15517) );
  INV_X1 U13380 ( .A(n10668), .ZN(n10669) );
  AOI22_X1 U13381 ( .A1(n10669), .A2(n15513), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n15262), .ZN(n10670) );
  OAI21_X1 U13382 ( .B1(n7840), .B2(n15517), .A(n10670), .ZN(n10671) );
  AOI21_X1 U13383 ( .B1(n15283), .B2(n15254), .A(n10671), .ZN(n10672) );
  INV_X1 U13384 ( .A(n12867), .ZN(n10676) );
  INV_X1 U13385 ( .A(n10679), .ZN(n10682) );
  OAI21_X1 U13386 ( .B1(n13199), .B2(n12890), .A(n10677), .ZN(n10678) );
  INV_X1 U13387 ( .A(n15866), .ZN(n12150) );
  OAI22_X1 U13388 ( .A1(n13201), .A2(n15859), .B1(n12756), .B2(n15861), .ZN(
        n10680) );
  INV_X1 U13389 ( .A(n10680), .ZN(n10681) );
  OAI21_X1 U13390 ( .B1(n10682), .B2(n15886), .A(n13214), .ZN(n10697) );
  AND2_X1 U13391 ( .A1(n10684), .A2(n10683), .ZN(n10685) );
  NAND2_X1 U13392 ( .A1(n11104), .A2(n10688), .ZN(n11102) );
  INV_X1 U13393 ( .A(n11104), .ZN(n10689) );
  OAI211_X1 U13394 ( .C1(n15901), .C2(n13023), .A(n9777), .B(n10689), .ZN(
        n10690) );
  OAI21_X1 U13395 ( .B1(n11102), .B2(n11105), .A(n10690), .ZN(n10691) );
  OR2_X1 U13396 ( .A1(n10697), .A2(n10706), .ZN(n10694) );
  INV_X1 U13397 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n10692) );
  NAND2_X1 U13398 ( .A1(n10706), .A2(n10692), .ZN(n10693) );
  NAND2_X1 U13399 ( .A1(n10694), .A2(n10693), .ZN(n10696) );
  NAND2_X1 U13400 ( .A1(n10696), .A2(n10695), .ZN(P3_U3486) );
  OR2_X1 U13401 ( .A1(n10697), .A2(n15906), .ZN(n10699) );
  OR2_X1 U13402 ( .A1(n15905), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n10698) );
  NAND2_X1 U13403 ( .A1(n10699), .A2(n10698), .ZN(n10703) );
  NAND2_X1 U13404 ( .A1(n10703), .A2(n10702), .ZN(P3_U3454) );
  INV_X1 U13405 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n10704) );
  NAND2_X1 U13406 ( .A1(n10706), .A2(n10704), .ZN(n10705) );
  NAND2_X1 U13407 ( .A1(n10708), .A2(n8082), .ZN(P3_U3487) );
  NAND2_X1 U13408 ( .A1(n14184), .A2(n14196), .ZN(n10710) );
  XNOR2_X1 U13409 ( .A(n14182), .B(n14496), .ZN(n14201) );
  NAND2_X1 U13410 ( .A1(n10714), .A2(n10711), .ZN(n10715) );
  INV_X1 U13411 ( .A(n10711), .ZN(n10712) );
  NOR2_X1 U13412 ( .A1(n14496), .A2(n10712), .ZN(n10713) );
  INV_X1 U13413 ( .A(n10716), .ZN(n14188) );
  INV_X1 U13414 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n12511) );
  NAND2_X1 U13415 ( .A1(n6512), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n10718) );
  NAND2_X1 U13416 ( .A1(n7281), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n10717) );
  OAI211_X1 U13417 ( .C1(n10381), .C2(n12511), .A(n10718), .B(n10717), .ZN(
        n10719) );
  OAI22_X1 U13418 ( .A1(n13993), .A2(n14472), .B1(n14059), .B2(n14474), .ZN(
        n12673) );
  OAI211_X1 U13419 ( .C1(n14205), .C2(n10722), .A(n11714), .B(n14187), .ZN(
        n14202) );
  INV_X1 U13420 ( .A(n10876), .ZN(n10869) );
  AND2_X1 U13421 ( .A1(n12037), .A2(n10725), .ZN(n11237) );
  INV_X1 U13422 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n15589) );
  MUX2_X1 U13423 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n15589), .S(n14859), .Z(
        n14862) );
  AND2_X1 U13424 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14861) );
  NAND2_X1 U13425 ( .A1(n14862), .A2(n14861), .ZN(n14860) );
  NAND2_X1 U13426 ( .A1(n14859), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10726) );
  NAND2_X1 U13427 ( .A1(n14860), .A2(n10726), .ZN(n14884) );
  INV_X1 U13428 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n15591) );
  MUX2_X1 U13429 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n15591), .S(n14879), .Z(
        n14885) );
  NAND2_X1 U13430 ( .A1(n14884), .A2(n14885), .ZN(n14883) );
  NAND2_X1 U13431 ( .A1(n14879), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n10727) );
  NAND2_X1 U13432 ( .A1(n14883), .A2(n10727), .ZN(n14897) );
  INV_X1 U13433 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n11089) );
  MUX2_X1 U13434 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n11089), .S(n14892), .Z(
        n14898) );
  NAND2_X1 U13435 ( .A1(n14897), .A2(n14898), .ZN(n14896) );
  NAND2_X1 U13436 ( .A1(n14892), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10728) );
  NAND2_X1 U13437 ( .A1(n14896), .A2(n10728), .ZN(n14906) );
  INV_X1 U13438 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n15593) );
  MUX2_X1 U13439 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n15593), .S(n14904), .Z(
        n14907) );
  NAND2_X1 U13440 ( .A1(n14906), .A2(n14907), .ZN(n14905) );
  NAND2_X1 U13441 ( .A1(n14904), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10729) );
  NAND2_X1 U13442 ( .A1(n14905), .A2(n10729), .ZN(n10920) );
  XNOR2_X1 U13443 ( .A(n10924), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n10921) );
  OR2_X1 U13444 ( .A1(n10924), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n10730) );
  NAND2_X1 U13445 ( .A1(n10918), .A2(n10730), .ZN(n10935) );
  INV_X1 U13446 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10731) );
  MUX2_X1 U13447 ( .A(n10731), .B(P1_REG1_REG_6__SCAN_IN), .S(n10939), .Z(
        n10936) );
  NAND2_X1 U13448 ( .A1(n10939), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10732) );
  NAND2_X1 U13449 ( .A1(n10933), .A2(n10732), .ZN(n14920) );
  INV_X1 U13450 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n11592) );
  MUX2_X1 U13451 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n11592), .S(n14918), .Z(
        n14921) );
  NAND2_X1 U13452 ( .A1(n14920), .A2(n14921), .ZN(n14919) );
  NAND2_X1 U13453 ( .A1(n14918), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10733) );
  NAND2_X1 U13454 ( .A1(n14919), .A2(n10733), .ZN(n10954) );
  MUX2_X1 U13455 ( .A(n8352), .B(P1_REG1_REG_8__SCAN_IN), .S(n10959), .Z(
        n10955) );
  OR2_X1 U13456 ( .A1(n10959), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10734) );
  XNOR2_X1 U13457 ( .A(n11006), .B(n10735), .ZN(n11004) );
  NOR2_X1 U13458 ( .A1(n11006), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n10736) );
  AOI21_X1 U13459 ( .B1(n11003), .B2(n11004), .A(n10736), .ZN(n14930) );
  INV_X1 U13460 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10737) );
  XNOR2_X1 U13461 ( .A(n14934), .B(n10737), .ZN(n14929) );
  NAND2_X1 U13462 ( .A1(n14930), .A2(n14929), .ZN(n14928) );
  NAND2_X1 U13463 ( .A1(n14934), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10738) );
  NAND2_X1 U13464 ( .A1(n14928), .A2(n10738), .ZN(n11163) );
  XNOR2_X1 U13465 ( .A(n11166), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n11164) );
  OR2_X1 U13466 ( .A1(n11166), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10739) );
  NAND2_X1 U13467 ( .A1(n11161), .A2(n10739), .ZN(n11307) );
  INV_X1 U13468 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10740) );
  XNOR2_X1 U13469 ( .A(n11316), .B(n10740), .ZN(n11308) );
  NAND2_X1 U13470 ( .A1(n11307), .A2(n11308), .ZN(n10742) );
  OR2_X1 U13471 ( .A1(n11316), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10741) );
  NAND2_X1 U13472 ( .A1(n10742), .A2(n10741), .ZN(n11595) );
  XNOR2_X1 U13473 ( .A(n11601), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n11596) );
  NAND2_X1 U13474 ( .A1(n11601), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n10743) );
  INV_X1 U13475 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10744) );
  XNOR2_X1 U13476 ( .A(n11621), .B(n10744), .ZN(n11620) );
  NAND2_X1 U13477 ( .A1(n11619), .A2(n11620), .ZN(n11618) );
  OR2_X1 U13478 ( .A1(n11621), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n10745) );
  NAND2_X1 U13479 ( .A1(n11618), .A2(n10745), .ZN(n10746) );
  XNOR2_X1 U13480 ( .A(n10746), .B(n11881), .ZN(n11877) );
  INV_X1 U13481 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n11876) );
  NAND2_X1 U13482 ( .A1(n11877), .A2(n11876), .ZN(n10748) );
  INV_X1 U13483 ( .A(n11881), .ZN(n11378) );
  NAND2_X1 U13484 ( .A1(n10746), .A2(n11378), .ZN(n10747) );
  NAND2_X1 U13485 ( .A1(n10748), .A2(n10747), .ZN(n12216) );
  XNOR2_X1 U13486 ( .A(n11212), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n12217) );
  NAND2_X1 U13487 ( .A1(n11212), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n10749) );
  NAND2_X1 U13488 ( .A1(n12213), .A2(n10749), .ZN(n14943) );
  XNOR2_X1 U13489 ( .A(n11448), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n14942) );
  NAND2_X1 U13490 ( .A1(n14943), .A2(n14942), .ZN(n14941) );
  NAND2_X1 U13491 ( .A1(n14947), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n10750) );
  NAND2_X1 U13492 ( .A1(n14941), .A2(n10750), .ZN(n10751) );
  NAND2_X1 U13493 ( .A1(n10751), .A2(n14961), .ZN(n10753) );
  AND2_X1 U13494 ( .A1(n10752), .A2(n10753), .ZN(n14956) );
  NAND2_X1 U13495 ( .A1(n14956), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n14955) );
  NAND2_X1 U13496 ( .A1(n14955), .A2(n10753), .ZN(n10754) );
  XNOR2_X1 U13497 ( .A(n10754), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n10791) );
  NAND2_X1 U13498 ( .A1(n10865), .A2(n10755), .ZN(n10796) );
  AOI21_X1 U13499 ( .B1(n10758), .B2(n10757), .A(n10756), .ZN(n10794) );
  NAND2_X1 U13500 ( .A1(n10796), .A2(n10794), .ZN(n10887) );
  INV_X1 U13501 ( .A(n15433), .ZN(n14971) );
  NAND2_X1 U13502 ( .A1(n10791), .A2(n14954), .ZN(n10789) );
  INV_X1 U13503 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n11435) );
  MUX2_X1 U13504 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n11435), .S(n14859), .Z(
        n14864) );
  AND2_X1 U13505 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14868) );
  NAND2_X1 U13506 ( .A1(n14864), .A2(n14868), .ZN(n14863) );
  NAND2_X1 U13507 ( .A1(n14859), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10759) );
  NAND2_X1 U13508 ( .A1(n14863), .A2(n10759), .ZN(n14881) );
  INV_X1 U13509 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n11506) );
  MUX2_X1 U13510 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n11506), .S(n14879), .Z(
        n14882) );
  NAND2_X1 U13511 ( .A1(n14881), .A2(n14882), .ZN(n14880) );
  NAND2_X1 U13512 ( .A1(n14879), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n10760) );
  NAND2_X1 U13513 ( .A1(n14880), .A2(n10760), .ZN(n14894) );
  INV_X1 U13514 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10761) );
  MUX2_X1 U13515 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10761), .S(n14892), .Z(
        n14895) );
  NAND2_X1 U13516 ( .A1(n14894), .A2(n14895), .ZN(n14893) );
  NAND2_X1 U13517 ( .A1(n14892), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n10762) );
  NAND2_X1 U13518 ( .A1(n14893), .A2(n10762), .ZN(n14909) );
  MUX2_X1 U13519 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n11389), .S(n14904), .Z(
        n14910) );
  NAND2_X1 U13520 ( .A1(n14909), .A2(n14910), .ZN(n14908) );
  NAND2_X1 U13521 ( .A1(n14904), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10763) );
  NAND2_X1 U13522 ( .A1(n14908), .A2(n10763), .ZN(n10926) );
  XNOR2_X1 U13523 ( .A(n10924), .B(n11495), .ZN(n10927) );
  NAND2_X1 U13524 ( .A1(n10926), .A2(n10927), .ZN(n10925) );
  NAND2_X1 U13525 ( .A1(n10924), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10764) );
  NAND2_X1 U13526 ( .A1(n10925), .A2(n10764), .ZN(n10941) );
  XNOR2_X1 U13527 ( .A(n10939), .B(n11574), .ZN(n10942) );
  NAND2_X1 U13528 ( .A1(n10941), .A2(n10942), .ZN(n10940) );
  NAND2_X1 U13529 ( .A1(n10939), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10765) );
  NAND2_X1 U13530 ( .A1(n10940), .A2(n10765), .ZN(n14923) );
  MUX2_X1 U13531 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n8334), .S(n14918), .Z(
        n14924) );
  NAND2_X1 U13532 ( .A1(n14923), .A2(n14924), .ZN(n14922) );
  NAND2_X1 U13533 ( .A1(n14918), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10766) );
  NAND2_X1 U13534 ( .A1(n14922), .A2(n10766), .ZN(n10962) );
  INV_X1 U13535 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11681) );
  XNOR2_X1 U13536 ( .A(n10959), .B(n11681), .ZN(n10961) );
  NAND2_X1 U13537 ( .A1(n10962), .A2(n10961), .ZN(n10960) );
  NAND2_X1 U13538 ( .A1(n10959), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10767) );
  NAND2_X1 U13539 ( .A1(n10960), .A2(n10767), .ZN(n11009) );
  INV_X1 U13540 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10768) );
  MUX2_X1 U13541 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10768), .S(n11006), .Z(
        n11008) );
  NAND2_X1 U13542 ( .A1(n11009), .A2(n11008), .ZN(n11007) );
  NAND2_X1 U13543 ( .A1(n11006), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10769) );
  NAND2_X1 U13544 ( .A1(n11007), .A2(n10769), .ZN(n14937) );
  XNOR2_X1 U13545 ( .A(n14934), .B(n11923), .ZN(n14936) );
  NAND2_X1 U13546 ( .A1(n14937), .A2(n14936), .ZN(n14935) );
  NAND2_X1 U13547 ( .A1(n14934), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10770) );
  NAND2_X1 U13548 ( .A1(n14935), .A2(n10770), .ZN(n11169) );
  XNOR2_X1 U13549 ( .A(n11166), .B(n10771), .ZN(n11168) );
  NAND2_X1 U13550 ( .A1(n11169), .A2(n11168), .ZN(n11167) );
  NAND2_X1 U13551 ( .A1(n11166), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10772) );
  NAND2_X1 U13552 ( .A1(n11167), .A2(n10772), .ZN(n11311) );
  MUX2_X1 U13553 ( .A(n12198), .B(P1_REG2_REG_12__SCAN_IN), .S(n11316), .Z(
        n11310) );
  OR2_X1 U13554 ( .A1(n11316), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10773) );
  NAND2_X1 U13555 ( .A1(n11313), .A2(n10773), .ZN(n11599) );
  XNOR2_X1 U13556 ( .A(n11601), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n11600) );
  NAND2_X1 U13557 ( .A1(n11601), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n10774) );
  NAND2_X1 U13558 ( .A1(n11597), .A2(n10774), .ZN(n11628) );
  INV_X1 U13559 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10775) );
  MUX2_X1 U13560 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n10775), .S(n11621), .Z(
        n11627) );
  NAND2_X1 U13561 ( .A1(n11628), .A2(n11627), .ZN(n11626) );
  NAND2_X1 U13562 ( .A1(n11621), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n10776) );
  NAND2_X1 U13563 ( .A1(n11626), .A2(n10776), .ZN(n10777) );
  XNOR2_X1 U13564 ( .A(n10777), .B(n11378), .ZN(n11874) );
  INV_X1 U13565 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11875) );
  NAND2_X1 U13566 ( .A1(n11874), .A2(n11875), .ZN(n10779) );
  OR2_X1 U13567 ( .A1(n10777), .A2(n11881), .ZN(n10778) );
  NAND2_X1 U13568 ( .A1(n10779), .A2(n10778), .ZN(n12221) );
  XNOR2_X1 U13569 ( .A(n11212), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n12222) );
  NAND2_X1 U13570 ( .A1(n11212), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n10780) );
  NAND2_X1 U13571 ( .A1(n12218), .A2(n10780), .ZN(n14950) );
  INV_X1 U13572 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n12520) );
  MUX2_X1 U13573 ( .A(n12520), .B(P1_REG2_REG_17__SCAN_IN), .S(n11448), .Z(
        n14949) );
  NAND2_X1 U13574 ( .A1(n14950), .A2(n14949), .ZN(n14948) );
  NAND2_X1 U13575 ( .A1(n14947), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n10781) );
  NAND2_X1 U13576 ( .A1(n14948), .A2(n10781), .ZN(n10782) );
  NAND2_X1 U13577 ( .A1(n10782), .A2(n14961), .ZN(n10785) );
  OR2_X1 U13578 ( .A1(n10782), .A2(n14961), .ZN(n10783) );
  NAND2_X1 U13579 ( .A1(n10785), .A2(n10783), .ZN(n14963) );
  INV_X1 U13580 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10784) );
  OR2_X1 U13581 ( .A1(n14963), .A2(n10784), .ZN(n14964) );
  NAND2_X1 U13582 ( .A1(n14964), .A2(n10785), .ZN(n10786) );
  XNOR2_X1 U13583 ( .A(n10786), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n10790) );
  NAND2_X1 U13584 ( .A1(n10888), .A2(n14971), .ZN(n10787) );
  OR2_X1 U13585 ( .A1(n10887), .A2(n10787), .ZN(n12220) );
  NAND2_X1 U13586 ( .A1(n10790), .A2(n14965), .ZN(n10788) );
  OR2_X1 U13587 ( .A1(n10887), .A2(n10888), .ZN(n12225) );
  NAND3_X1 U13588 ( .A1(n10789), .A2(n10788), .A3(n12225), .ZN(n10793) );
  OAI22_X1 U13589 ( .A1(n10791), .A2(n12215), .B1(n10790), .B2(n12220), .ZN(
        n10792) );
  AND2_X1 U13590 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14704) );
  INV_X1 U13591 ( .A(n10794), .ZN(n10795) );
  NAND2_X1 U13592 ( .A1(n10796), .A2(n10795), .ZN(n14959) );
  NOR2_X1 U13593 ( .A1(n14959), .A2(n8117), .ZN(n10797) );
  XNOR2_X1 U13594 ( .A(n11420), .B(n15800), .ZN(n13757) );
  NAND2_X1 U13595 ( .A1(n11338), .A2(n14311), .ZN(n11398) );
  NAND2_X1 U13596 ( .A1(n10801), .A2(n13757), .ZN(n10803) );
  INV_X1 U13597 ( .A(n13762), .ZN(n11270) );
  XNOR2_X1 U13598 ( .A(n7648), .B(n11420), .ZN(n11460) );
  AND2_X1 U13599 ( .A1(n14311), .A2(n14101), .ZN(n10804) );
  NAND2_X1 U13600 ( .A1(n11460), .A2(n10804), .ZN(n11416) );
  NAND2_X1 U13601 ( .A1(n11416), .A2(n10805), .ZN(n10815) );
  INV_X1 U13602 ( .A(n15795), .ZN(n10807) );
  NAND2_X1 U13603 ( .A1(n10807), .A2(n10806), .ZN(n11787) );
  INV_X1 U13604 ( .A(n15812), .ZN(n15831) );
  NAND3_X1 U13605 ( .A1(n15831), .A2(n15796), .A3(n10810), .ZN(n10811) );
  OR2_X2 U13606 ( .A1(n10822), .A2(n10811), .ZN(n13796) );
  INV_X1 U13607 ( .A(n11457), .ZN(n10814) );
  NAND2_X1 U13608 ( .A1(n10822), .A2(n10823), .ZN(n11274) );
  INV_X1 U13609 ( .A(n10817), .ZN(n10818) );
  NAND2_X1 U13610 ( .A1(n11274), .A2(n10818), .ZN(n10819) );
  NOR2_X1 U13611 ( .A1(n13804), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n10828) );
  NAND2_X1 U13612 ( .A1(n15796), .A2(n14070), .ZN(n10820) );
  OAI22_X1 U13613 ( .A1(n10389), .A2(n13805), .B1(n13803), .B2(n13842), .ZN(
        n10827) );
  AND2_X1 U13614 ( .A1(n11209), .A2(n14065), .ZN(n11800) );
  NAND2_X1 U13615 ( .A1(n11800), .A2(n15796), .ZN(n10821) );
  OR2_X1 U13616 ( .A1(n10822), .A2(n10821), .ZN(n10825) );
  OAI22_X1 U13617 ( .A1(n13733), .A2(n11905), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10391), .ZN(n10826) );
  OR4_X1 U13618 ( .A1(n10829), .A2(n10828), .A3(n10827), .A4(n10826), .ZN(
        P2_U3190) );
  NAND2_X1 U13619 ( .A1(n10879), .A2(P3_U3151), .ZN(n13611) );
  INV_X1 U13620 ( .A(n13611), .ZN(n11928) );
  AND2_X1 U13621 ( .A1(n10878), .A2(P3_U3151), .ZN(n13605) );
  AOI222_X1 U13622 ( .A1(n10830), .A2(n11928), .B1(SI_4_), .B2(n13605), .C1(
        n11158), .C2(P3_STATE_REG_SCAN_IN), .ZN(n10831) );
  INV_X1 U13623 ( .A(n10831), .ZN(P3_U3291) );
  INV_X2 U13624 ( .A(n13605), .ZN(n13618) );
  INV_X1 U13625 ( .A(SI_3_), .ZN(n10835) );
  INV_X1 U13626 ( .A(n10832), .ZN(n10834) );
  OAI222_X1 U13627 ( .A1(n13618), .A2(n10835), .B1(n13611), .B2(n10834), .C1(
        P3_U3151), .C2(n10833), .ZN(P3_U3292) );
  OAI222_X1 U13628 ( .A1(n12295), .A2(P3_U3151), .B1(n13611), .B2(n10837), 
        .C1(n10836), .C2(n13618), .ZN(P3_U3295) );
  NAND2_X1 U13629 ( .A1(n10878), .A2(P2_U3088), .ZN(n14663) );
  INV_X1 U13630 ( .A(n14663), .ZN(n14664) );
  INV_X1 U13631 ( .A(n14664), .ZN(n14673) );
  INV_X1 U13632 ( .A(n10838), .ZN(n10899) );
  OAI222_X1 U13633 ( .A1(n14671), .A2(n10839), .B1(n14673), .B2(n10899), .C1(
        n11242), .C2(n14117), .ZN(P2_U3324) );
  OAI222_X1 U13634 ( .A1(n14671), .A2(n10840), .B1(n14673), .B2(n10881), .C1(
        P2_U3088), .C2(n15609), .ZN(P2_U3325) );
  INV_X1 U13635 ( .A(n10841), .ZN(n10843) );
  INV_X1 U13636 ( .A(SI_8_), .ZN(n10842) );
  OAI222_X1 U13637 ( .A1(n13622), .A2(n10843), .B1(n13618), .B2(n10842), .C1(
        n11552), .C2(P3_U3151), .ZN(P3_U3287) );
  INV_X1 U13638 ( .A(n10844), .ZN(n10846) );
  INV_X1 U13639 ( .A(SI_5_), .ZN(n10845) );
  OAI222_X1 U13640 ( .A1(n13622), .A2(n10846), .B1(n13618), .B2(n10845), .C1(
        n11202), .C2(P3_U3151), .ZN(P3_U3290) );
  OAI222_X1 U13641 ( .A1(n14105), .A2(n11242), .B1(n14663), .B2(n10907), .C1(
        n10847), .C2(n14671), .ZN(P2_U3326) );
  INV_X1 U13642 ( .A(n10848), .ZN(n11042) );
  OAI222_X1 U13643 ( .A1(P3_U3151), .A2(n11042), .B1(n13618), .B2(n10850), 
        .C1(n13622), .C2(n10849), .ZN(P3_U3294) );
  INV_X1 U13644 ( .A(SI_7_), .ZN(n10851) );
  OAI222_X1 U13645 ( .A1(n11297), .A2(P3_U3151), .B1(n13622), .B2(n10852), 
        .C1(n10851), .C2(n13618), .ZN(P3_U3288) );
  INV_X1 U13646 ( .A(n10853), .ZN(n10855) );
  OAI222_X1 U13647 ( .A1(n10856), .A2(P3_U3151), .B1(n13622), .B2(n10855), 
        .C1(n10854), .C2(n13618), .ZN(P3_U3293) );
  OAI222_X1 U13648 ( .A1(n11185), .A2(P3_U3151), .B1(n13622), .B2(n10858), 
        .C1(n10857), .C2(n13618), .ZN(P3_U3289) );
  INV_X1 U13649 ( .A(n10859), .ZN(n10895) );
  INV_X1 U13650 ( .A(n11253), .ZN(n15621) );
  OAI222_X1 U13651 ( .A1(n14671), .A2(n7693), .B1(n14673), .B2(n10895), .C1(
        n11242), .C2(n15621), .ZN(P2_U3323) );
  OAI222_X1 U13652 ( .A1(n11740), .A2(P3_U3151), .B1(n13622), .B2(n10861), 
        .C1(n10860), .C2(n13618), .ZN(P3_U3286) );
  NAND2_X1 U13653 ( .A1(n14836), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n10862) );
  OAI21_X1 U13654 ( .B1(n15008), .B2(n14836), .A(n10862), .ZN(P1_U3590) );
  INV_X1 U13655 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10864) );
  INV_X1 U13656 ( .A(n10863), .ZN(n10897) );
  INV_X1 U13657 ( .A(n11255), .ZN(n15634) );
  OAI222_X1 U13658 ( .A1(n14671), .A2(n10864), .B1(n14673), .B2(n10897), .C1(
        n6510), .C2(n15634), .ZN(P2_U3322) );
  INV_X1 U13659 ( .A(n10865), .ZN(n10866) );
  INV_X1 U13660 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10871) );
  NOR3_X1 U13661 ( .A1(n8979), .A2(n10869), .A3(n10868), .ZN(n10870) );
  AOI21_X1 U13662 ( .B1(n15531), .B2(n10871), .A(n10870), .ZN(P1_U3446) );
  OAI222_X1 U13663 ( .A1(n13622), .A2(n10874), .B1(n13618), .B2(n10873), .C1(
        n10872), .C2(P3_U3151), .ZN(P3_U3285) );
  INV_X1 U13664 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n12509) );
  INV_X1 U13665 ( .A(n10875), .ZN(n10877) );
  AOI22_X1 U13666 ( .A1(n15531), .A2(n12509), .B1(n10877), .B2(n10876), .ZN(
        P1_U3445) );
  NAND2_X1 U13667 ( .A1(n10878), .A2(P1_U3086), .ZN(n15435) );
  INV_X1 U13668 ( .A(n14879), .ZN(n10880) );
  OAI222_X1 U13669 ( .A1(n15435), .A2(n12482), .B1(n15438), .B2(n10881), .C1(
        P1_U3086), .C2(n10880), .ZN(P1_U3353) );
  INV_X1 U13670 ( .A(n14959), .ZN(n12223) );
  NOR2_X1 U13671 ( .A1(n12223), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U13672 ( .A(n10882), .ZN(n10885) );
  OAI222_X1 U13673 ( .A1(n14671), .A2(n10883), .B1(n14673), .B2(n10885), .C1(
        P2_U3088), .C2(n15646), .ZN(P2_U3321) );
  INV_X1 U13674 ( .A(n10939), .ZN(n10884) );
  OAI222_X1 U13675 ( .A1(n15435), .A2(n10886), .B1(n15438), .B2(n10885), .C1(
        P1_U3086), .C2(n10884), .ZN(P1_U3349) );
  INV_X1 U13676 ( .A(n10887), .ZN(n10892) );
  INV_X1 U13677 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10889) );
  OAI21_X1 U13678 ( .B1(n15433), .B2(P1_REG2_REG_0__SCAN_IN), .A(n10888), .ZN(
        n14872) );
  AOI21_X1 U13679 ( .B1(n15433), .B2(n10889), .A(n14872), .ZN(n10890) );
  INV_X1 U13680 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14871) );
  XNOR2_X1 U13681 ( .A(n10890), .B(n14871), .ZN(n10891) );
  AOI22_X1 U13682 ( .A1(n10892), .A2(n10891), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10893) );
  OAI21_X1 U13683 ( .B1(n14959), .B2(n7320), .A(n10893), .ZN(P1_U3243) );
  INV_X1 U13684 ( .A(n15435), .ZN(n15424) );
  AOI22_X1 U13685 ( .A1(n14904), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n15424), .ZN(n10894) );
  OAI21_X1 U13686 ( .B1(n10895), .B2(n15438), .A(n10894), .ZN(P1_U3351) );
  AOI22_X1 U13687 ( .A1(n10924), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n15424), .ZN(n10896) );
  OAI21_X1 U13688 ( .B1(n10897), .B2(n15438), .A(n10896), .ZN(P1_U3350) );
  INV_X1 U13689 ( .A(n14892), .ZN(n10898) );
  OAI222_X1 U13690 ( .A1(n15435), .A2(n12296), .B1(n15438), .B2(n10899), .C1(
        P1_U3086), .C2(n10898), .ZN(P1_U3352) );
  NAND2_X1 U13691 ( .A1(n10972), .A2(P3_D_REG_1__SCAN_IN), .ZN(n10900) );
  OAI21_X1 U13692 ( .B1(n11105), .B2(n10972), .A(n10900), .ZN(P3_U3377) );
  OAI222_X1 U13693 ( .A1(n10903), .A2(P3_U3151), .B1(n13622), .B2(n10902), 
        .C1(n10901), .C2(n13618), .ZN(P3_U3284) );
  INV_X1 U13694 ( .A(n10904), .ZN(n10909) );
  AOI22_X1 U13695 ( .A1(n14918), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n15424), .ZN(n10905) );
  OAI21_X1 U13696 ( .B1(n10909), .B2(n15438), .A(n10905), .ZN(P1_U3348) );
  INV_X1 U13697 ( .A(n14859), .ZN(n10908) );
  OAI222_X1 U13698 ( .A1(n10908), .A2(P1_U3086), .B1(n15438), .B2(n10907), 
        .C1(n10906), .C2(n15435), .ZN(P1_U3354) );
  INV_X1 U13699 ( .A(n11259), .ZN(n14129) );
  OAI222_X1 U13700 ( .A1(n14671), .A2(n10910), .B1(n14673), .B2(n10909), .C1(
        n6510), .C2(n14129), .ZN(P2_U3320) );
  INV_X1 U13701 ( .A(n10911), .ZN(n10914) );
  INV_X1 U13702 ( .A(n11262), .ZN(n15659) );
  OAI222_X1 U13703 ( .A1(n14671), .A2(n10912), .B1(n14673), .B2(n10914), .C1(
        P2_U3088), .C2(n15659), .ZN(P2_U3319) );
  INV_X1 U13704 ( .A(n10959), .ZN(n10913) );
  OAI222_X1 U13705 ( .A1(n15435), .A2(n8144), .B1(n15438), .B2(n10914), .C1(
        P1_U3086), .C2(n10913), .ZN(P1_U3347) );
  OAI222_X1 U13706 ( .A1(n10917), .A2(P3_U3151), .B1(n13622), .B2(n10916), 
        .C1(n10915), .C2(n13618), .ZN(P3_U3283) );
  INV_X1 U13707 ( .A(n10918), .ZN(n10919) );
  AOI21_X1 U13708 ( .B1(n10921), .B2(n10920), .A(n10919), .ZN(n10930) );
  NAND2_X1 U13709 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n11357) );
  OAI21_X1 U13710 ( .B1(n14959), .B2(n10922), .A(n11357), .ZN(n10923) );
  AOI21_X1 U13711 ( .B1(n14962), .B2(n10924), .A(n10923), .ZN(n10929) );
  OAI211_X1 U13712 ( .C1(n10927), .C2(n10926), .A(n14965), .B(n10925), .ZN(
        n10928) );
  OAI211_X1 U13713 ( .C1(n10930), .C2(n12215), .A(n10929), .B(n10928), .ZN(
        P1_U3248) );
  NAND2_X1 U13714 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n10931) );
  OAI21_X1 U13715 ( .B1(n14959), .B2(n10932), .A(n10931), .ZN(n10938) );
  INV_X1 U13716 ( .A(n10933), .ZN(n10934) );
  AOI211_X1 U13717 ( .C1(n10936), .C2(n10935), .A(n10934), .B(n12215), .ZN(
        n10937) );
  AOI211_X1 U13718 ( .C1(n14962), .C2(n10939), .A(n10938), .B(n10937), .ZN(
        n10944) );
  OAI211_X1 U13719 ( .C1(n10942), .C2(n10941), .A(n14965), .B(n10940), .ZN(
        n10943) );
  NAND2_X1 U13720 ( .A1(n10944), .A2(n10943), .ZN(P1_U3249) );
  INV_X1 U13721 ( .A(n10222), .ZN(n10947) );
  INV_X1 U13722 ( .A(n11263), .ZN(n15676) );
  OAI222_X1 U13723 ( .A1(n14671), .A2(n10945), .B1(n14673), .B2(n10947), .C1(
        n6510), .C2(n15676), .ZN(P2_U3318) );
  INV_X1 U13724 ( .A(n11006), .ZN(n10946) );
  OAI222_X1 U13725 ( .A1(n15435), .A2(n12483), .B1(n15438), .B2(n10947), .C1(
        P1_U3086), .C2(n10946), .ZN(P1_U3346) );
  NAND2_X1 U13726 ( .A1(n13819), .A2(P2_U3947), .ZN(n10948) );
  OAI21_X1 U13727 ( .B1(n9028), .B2(P2_U3947), .A(n10948), .ZN(P2_U3531) );
  INV_X1 U13728 ( .A(n10949), .ZN(n10970) );
  AOI22_X1 U13729 ( .A1(n14934), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n15424), .ZN(n10950) );
  OAI21_X1 U13730 ( .B1(n10970), .B2(n15438), .A(n10950), .ZN(P1_U3345) );
  INV_X1 U13731 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n12418) );
  NAND2_X1 U13732 ( .A1(P3_U3897), .A2(n9055), .ZN(n10951) );
  OAI21_X1 U13733 ( .B1(P3_U3897), .B2(n12418), .A(n10951), .ZN(P3_U3493) );
  INV_X1 U13734 ( .A(n10952), .ZN(n10953) );
  AOI21_X1 U13735 ( .B1(n10955), .B2(n10954), .A(n10953), .ZN(n10965) );
  NAND2_X1 U13736 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n10956) );
  OAI21_X1 U13737 ( .B1(n14959), .B2(n10957), .A(n10956), .ZN(n10958) );
  AOI21_X1 U13738 ( .B1(n14962), .B2(n10959), .A(n10958), .ZN(n10964) );
  OAI211_X1 U13739 ( .C1(n10962), .C2(n10961), .A(n10960), .B(n14965), .ZN(
        n10963) );
  OAI211_X1 U13740 ( .C1(n10965), .C2(n12215), .A(n10964), .B(n10963), .ZN(
        P1_U3251) );
  INV_X1 U13741 ( .A(n10966), .ZN(n10969) );
  INV_X1 U13742 ( .A(n11644), .ZN(n11247) );
  OAI222_X1 U13743 ( .A1(n14671), .A2(n10967), .B1(n14663), .B2(n10969), .C1(
        P2_U3088), .C2(n11247), .ZN(P2_U3316) );
  INV_X1 U13744 ( .A(n11166), .ZN(n10968) );
  OAI222_X1 U13745 ( .A1(n15435), .A2(n12309), .B1(n15438), .B2(n10969), .C1(
        P1_U3086), .C2(n10968), .ZN(P1_U3344) );
  INV_X1 U13746 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10971) );
  OAI222_X1 U13747 ( .A1(n14671), .A2(n10971), .B1(n14663), .B2(n10970), .C1(
        n6510), .C2(n11232), .ZN(P2_U3317) );
  INV_X1 U13748 ( .A(n9557), .ZN(n10973) );
  INV_X1 U13749 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10974) );
  NOR2_X1 U13750 ( .A1(n10993), .A2(n10974), .ZN(P3_U3262) );
  CLKBUF_X1 U13751 ( .A(n10975), .Z(n10993) );
  INV_X1 U13752 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10976) );
  NOR2_X1 U13753 ( .A1(n10993), .A2(n10976), .ZN(P3_U3263) );
  INV_X1 U13754 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10977) );
  NOR2_X1 U13755 ( .A1(n10975), .A2(n10977), .ZN(P3_U3241) );
  INV_X1 U13756 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10978) );
  NOR2_X1 U13757 ( .A1(n10975), .A2(n10978), .ZN(P3_U3239) );
  INV_X1 U13758 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10979) );
  NOR2_X1 U13759 ( .A1(n10975), .A2(n10979), .ZN(P3_U3238) );
  INV_X1 U13760 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10980) );
  NOR2_X1 U13761 ( .A1(n10975), .A2(n10980), .ZN(P3_U3237) );
  INV_X1 U13762 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10981) );
  NOR2_X1 U13763 ( .A1(n10975), .A2(n10981), .ZN(P3_U3236) );
  INV_X1 U13764 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10982) );
  NOR2_X1 U13765 ( .A1(n10975), .A2(n10982), .ZN(P3_U3235) );
  INV_X1 U13766 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n12481) );
  NOR2_X1 U13767 ( .A1(n10975), .A2(n12481), .ZN(P3_U3234) );
  INV_X1 U13768 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10983) );
  NOR2_X1 U13769 ( .A1(n10993), .A2(n10983), .ZN(P3_U3261) );
  INV_X1 U13770 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10984) );
  NOR2_X1 U13771 ( .A1(n10975), .A2(n10984), .ZN(P3_U3260) );
  INV_X1 U13772 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n12347) );
  NOR2_X1 U13773 ( .A1(n10993), .A2(n12347), .ZN(P3_U3259) );
  INV_X1 U13774 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10985) );
  NOR2_X1 U13775 ( .A1(n10975), .A2(n10985), .ZN(P3_U3258) );
  INV_X1 U13776 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10986) );
  NOR2_X1 U13777 ( .A1(n10993), .A2(n10986), .ZN(P3_U3257) );
  INV_X1 U13778 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10987) );
  NOR2_X1 U13779 ( .A1(n10993), .A2(n10987), .ZN(P3_U3256) );
  INV_X1 U13780 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10988) );
  NOR2_X1 U13781 ( .A1(n10993), .A2(n10988), .ZN(P3_U3255) );
  INV_X1 U13782 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10989) );
  NOR2_X1 U13783 ( .A1(n10993), .A2(n10989), .ZN(P3_U3254) );
  INV_X1 U13784 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n12426) );
  NOR2_X1 U13785 ( .A1(n10993), .A2(n12426), .ZN(P3_U3253) );
  INV_X1 U13786 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10990) );
  NOR2_X1 U13787 ( .A1(n10993), .A2(n10990), .ZN(P3_U3252) );
  INV_X1 U13788 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n12420) );
  NOR2_X1 U13789 ( .A1(n10993), .A2(n12420), .ZN(P3_U3251) );
  INV_X1 U13790 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n12354) );
  NOR2_X1 U13791 ( .A1(n10993), .A2(n12354), .ZN(P3_U3250) );
  INV_X1 U13792 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10991) );
  NOR2_X1 U13793 ( .A1(n10993), .A2(n10991), .ZN(P3_U3249) );
  INV_X1 U13794 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n12344) );
  NOR2_X1 U13795 ( .A1(n10993), .A2(n12344), .ZN(P3_U3248) );
  INV_X1 U13796 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10992) );
  NOR2_X1 U13797 ( .A1(n10993), .A2(n10992), .ZN(P3_U3247) );
  INV_X1 U13798 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n12288) );
  NOR2_X1 U13799 ( .A1(n10993), .A2(n12288), .ZN(P3_U3246) );
  INV_X1 U13800 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10994) );
  NOR2_X1 U13801 ( .A1(n10975), .A2(n10994), .ZN(P3_U3245) );
  INV_X1 U13802 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10995) );
  NOR2_X1 U13803 ( .A1(n10975), .A2(n10995), .ZN(P3_U3244) );
  INV_X1 U13804 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n12282) );
  NOR2_X1 U13805 ( .A1(n10993), .A2(n12282), .ZN(P3_U3243) );
  INV_X1 U13806 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10996) );
  NOR2_X1 U13807 ( .A1(n10993), .A2(n10996), .ZN(P3_U3242) );
  INV_X1 U13808 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10997) );
  NOR2_X1 U13809 ( .A1(n10993), .A2(n10997), .ZN(P3_U3240) );
  OAI222_X1 U13810 ( .A1(n13611), .A2(n11000), .B1(n13618), .B2(n10999), .C1(
        n10998), .C2(P3_U3151), .ZN(P3_U3282) );
  INV_X1 U13811 ( .A(n11001), .ZN(n11022) );
  AOI22_X1 U13812 ( .A1(n11316), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n15424), .ZN(n11002) );
  OAI21_X1 U13813 ( .B1(n11022), .B2(n15438), .A(n11002), .ZN(P1_U3343) );
  XOR2_X1 U13814 ( .A(n11004), .B(n11003), .Z(n11012) );
  NAND2_X1 U13815 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n12063) );
  OAI21_X1 U13816 ( .B1(n14959), .B2(n6813), .A(n12063), .ZN(n11005) );
  AOI21_X1 U13817 ( .B1(n14962), .B2(n11006), .A(n11005), .ZN(n11011) );
  OAI211_X1 U13818 ( .C1(n11009), .C2(n11008), .A(n11007), .B(n14965), .ZN(
        n11010) );
  OAI211_X1 U13819 ( .C1(n11012), .C2(n12215), .A(n11011), .B(n11010), .ZN(
        P1_U3252) );
  INV_X1 U13820 ( .A(n11013), .ZN(n11015) );
  OAI222_X1 U13821 ( .A1(n7404), .A2(P3_U3151), .B1(n13611), .B2(n11015), .C1(
        n11014), .C2(n13618), .ZN(P3_U3280) );
  INV_X1 U13822 ( .A(n11450), .ZN(n11018) );
  INV_X1 U13823 ( .A(n11453), .ZN(n11016) );
  AOI21_X1 U13824 ( .B1(n15360), .B2(n15560), .A(n11016), .ZN(n11017) );
  AOI211_X1 U13825 ( .C1(n11019), .C2(n11055), .A(n11018), .B(n11017), .ZN(
        n15533) );
  NAND2_X1 U13826 ( .A1(n15597), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n11020) );
  OAI21_X1 U13827 ( .B1(n15533), .B2(n15597), .A(n11020), .ZN(P1_U3528) );
  INV_X1 U13828 ( .A(n15701), .ZN(n11021) );
  OAI222_X1 U13829 ( .A1(n14671), .A2(n11023), .B1(n14663), .B2(n11022), .C1(
        n11021), .C2(P2_U3088), .ZN(P2_U3315) );
  XNOR2_X1 U13830 ( .A(n11024), .B(n11025), .ZN(n11026) );
  NAND2_X1 U13831 ( .A1(n11026), .A2(n14813), .ZN(n11031) );
  NAND2_X1 U13832 ( .A1(n14854), .A2(n15256), .ZN(n11027) );
  NAND2_X1 U13833 ( .A1(n11028), .A2(n11027), .ZN(n15541) );
  OR2_X1 U13834 ( .A1(n11029), .A2(P1_U3086), .ZN(n14708) );
  AOI22_X1 U13835 ( .A1(n15500), .A2(n15541), .B1(n14708), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n11030) );
  OAI211_X1 U13836 ( .C1(n8299), .C2(n15503), .A(n11031), .B(n11030), .ZN(
        P1_U3237) );
  XNOR2_X1 U13837 ( .A(n11033), .B(P3_REG1_REG_1__SCAN_IN), .ZN(n11034) );
  AOI22_X1 U13838 ( .A1(n13097), .A2(n11035), .B1(n13180), .B2(n11034), .ZN(
        n11041) );
  AOI21_X1 U13839 ( .B1(n11037), .B2(n11403), .A(n11036), .ZN(n11038) );
  OAI22_X1 U13840 ( .A1(n13146), .A2(n11038), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11099), .ZN(n11039) );
  AOI21_X1 U13841 ( .B1(n15849), .B2(P3_ADDR_REG_1__SCAN_IN), .A(n11039), .ZN(
        n11040) );
  OAI211_X1 U13842 ( .C1(n11042), .C2(n13171), .A(n11041), .B(n11040), .ZN(
        P3_U3183) );
  INV_X1 U13843 ( .A(n11043), .ZN(n11045) );
  OAI222_X1 U13844 ( .A1(n13095), .A2(P3_U3151), .B1(n13611), .B2(n11045), 
        .C1(n11044), .C2(n13618), .ZN(P3_U3281) );
  INV_X1 U13845 ( .A(n11601), .ZN(n11048) );
  INV_X1 U13846 ( .A(n11046), .ZN(n11050) );
  OAI222_X1 U13847 ( .A1(P1_U3086), .A2(n11048), .B1(n15438), .B2(n11050), 
        .C1(n11047), .C2(n15435), .ZN(P1_U3342) );
  INV_X1 U13848 ( .A(n14149), .ZN(n11049) );
  OAI222_X1 U13849 ( .A1(n14671), .A2(n11051), .B1(n14663), .B2(n11050), .C1(
        n11049), .C2(n6510), .ZN(P2_U3314) );
  INV_X1 U13850 ( .A(n11052), .ZN(n11054) );
  OAI222_X1 U13851 ( .A1(n13611), .A2(n11054), .B1(n13618), .B2(n11053), .C1(
        n13123), .C2(P3_U3151), .ZN(P3_U3279) );
  XNOR2_X1 U13852 ( .A(n11057), .B(n11056), .ZN(n14870) );
  AOI22_X1 U13853 ( .A1(n14813), .A2(n14870), .B1(n14708), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n11058) );
  NAND2_X1 U13854 ( .A1(n11059), .A2(n11058), .ZN(P1_U3232) );
  NOR2_X1 U13855 ( .A1(n12839), .A2(P3_U3151), .ZN(n11286) );
  NAND2_X1 U13856 ( .A1(n13044), .A2(n11327), .ZN(n12899) );
  INV_X1 U13857 ( .A(n12899), .ZN(n11061) );
  INV_X1 U13858 ( .A(n12897), .ZN(n11060) );
  NOR2_X1 U13859 ( .A1(n11061), .A2(n11060), .ZN(n12877) );
  INV_X1 U13860 ( .A(n12877), .ZN(n11063) );
  OAI22_X1 U13861 ( .A1(n12842), .A2(n11327), .B1(n15860), .B2(n12822), .ZN(
        n11062) );
  AOI21_X1 U13862 ( .B1(n12832), .B2(n11063), .A(n11062), .ZN(n11064) );
  OAI21_X1 U13863 ( .B1(n11286), .B2(n11404), .A(n11064), .ZN(P3_U3172) );
  INV_X1 U13864 ( .A(n11065), .ZN(n11068) );
  OAI222_X1 U13865 ( .A1(n13611), .A2(n11068), .B1(n13618), .B2(n11067), .C1(
        n11066), .C2(P3_U3151), .ZN(P3_U3278) );
  INV_X1 U13866 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n11082) );
  XNOR2_X1 U13867 ( .A(n11069), .B(n11070), .ZN(n11468) );
  NAND2_X1 U13868 ( .A1(n11468), .A2(n15552), .ZN(n11077) );
  OAI21_X1 U13869 ( .B1(n11073), .B2(n11072), .A(n11071), .ZN(n11075) );
  NAND2_X1 U13870 ( .A1(n14855), .A2(n15257), .ZN(n11074) );
  OAI21_X1 U13871 ( .B1(n11489), .B2(n15227), .A(n11074), .ZN(n15499) );
  AOI21_X1 U13872 ( .B1(n11075), .B2(n15545), .A(n15499), .ZN(n11076) );
  AND2_X1 U13873 ( .A1(n11077), .A2(n11076), .ZN(n11469) );
  INV_X1 U13874 ( .A(n15548), .ZN(n15574) );
  NAND2_X1 U13875 ( .A1(n11504), .A2(n11472), .ZN(n11078) );
  NAND2_X1 U13876 ( .A1(n11391), .A2(n11078), .ZN(n11470) );
  OAI22_X1 U13877 ( .A1(n11470), .A2(n15571), .B1(n15502), .B2(n15569), .ZN(
        n11079) );
  AOI21_X1 U13878 ( .B1(n11468), .B2(n15574), .A(n11079), .ZN(n11080) );
  NAND2_X1 U13879 ( .A1(n11469), .A2(n11080), .ZN(n11087) );
  NAND2_X1 U13880 ( .A1(n11087), .A2(n15588), .ZN(n11081) );
  OAI21_X1 U13881 ( .B1(n15588), .B2(n11082), .A(n11081), .ZN(P1_U3468) );
  AOI21_X1 U13882 ( .B1(n13401), .B2(n11083), .A(n12877), .ZN(n11084) );
  AOI21_X1 U13883 ( .B1(n13420), .B2(n13042), .A(n11084), .ZN(n11324) );
  INV_X1 U13884 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11085) );
  MUX2_X1 U13885 ( .A(n11324), .B(n11085), .S(n15906), .Z(n11086) );
  OAI21_X1 U13886 ( .B1(n11327), .B2(n13599), .A(n11086), .ZN(P3_U3390) );
  NAND2_X1 U13887 ( .A1(n11087), .A2(n15599), .ZN(n11088) );
  OAI21_X1 U13888 ( .B1(n15599), .B2(n11089), .A(n11088), .ZN(P1_U3531) );
  INV_X1 U13889 ( .A(n13044), .ZN(n11090) );
  OAI22_X1 U13890 ( .A1(n11090), .A2(n12836), .B1(n12822), .B2(n11668), .ZN(
        n11091) );
  AOI21_X1 U13891 ( .B1(n12803), .B2(n11092), .A(n11091), .ZN(n11098) );
  OAI21_X1 U13892 ( .B1(n11095), .B2(n11094), .A(n11093), .ZN(n11096) );
  NAND2_X1 U13893 ( .A1(n11096), .A2(n12832), .ZN(n11097) );
  OAI211_X1 U13894 ( .C1(n11286), .C2(n11099), .A(n11098), .B(n11097), .ZN(
        P3_U3162) );
  NAND2_X1 U13895 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n14103), .ZN(n11100) );
  OAI21_X1 U13896 ( .B1(n13909), .B2(n14103), .A(n11100), .ZN(P2_U3551) );
  OR2_X1 U13897 ( .A1(n11102), .A2(n11101), .ZN(n11103) );
  OAI21_X1 U13898 ( .B1(n11105), .B2(n11104), .A(n11103), .ZN(n11108) );
  NAND2_X1 U13899 ( .A1(n11110), .A2(n11108), .ZN(n11107) );
  MUX2_X1 U13900 ( .A(n11324), .B(n11406), .S(n15873), .Z(n11112) );
  NOR2_X1 U13901 ( .A1(n15901), .A2(n15853), .ZN(n11109) );
  AOI22_X1 U13902 ( .A1(n13428), .A2(n11662), .B1(n13427), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n11111) );
  NAND2_X1 U13903 ( .A1(n11112), .A2(n11111), .ZN(P3_U3233) );
  XOR2_X1 U13904 ( .A(n11114), .B(n11113), .Z(n11126) );
  OAI21_X1 U13905 ( .B1(P3_REG2_REG_3__SCAN_IN), .B2(n11116), .A(n11115), .ZN(
        n11117) );
  INV_X1 U13906 ( .A(n11117), .ZN(n11122) );
  XNOR2_X1 U13907 ( .A(n11118), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n11119) );
  NAND2_X1 U13908 ( .A1(n13180), .A2(n11119), .ZN(n11121) );
  NOR2_X1 U13909 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9075), .ZN(n11333) );
  AOI21_X1 U13910 ( .B1(n15849), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n11333), .ZN(
        n11120) );
  OAI211_X1 U13911 ( .C1(n11122), .C2(n13182), .A(n11121), .B(n11120), .ZN(
        n11123) );
  AOI21_X1 U13912 ( .B1(n13152), .B2(n11124), .A(n11123), .ZN(n11125) );
  OAI21_X1 U13913 ( .B1(n11126), .B2(n13146), .A(n11125), .ZN(P3_U3185) );
  OAI222_X1 U13914 ( .A1(n13611), .A2(n11128), .B1(n13618), .B2(n11127), .C1(
        n13175), .C2(P3_U3151), .ZN(P3_U3277) );
  XOR2_X1 U13915 ( .A(n11130), .B(n11129), .Z(n11143) );
  OAI21_X1 U13916 ( .B1(n11133), .B2(n11132), .A(n11131), .ZN(n11136) );
  NAND2_X1 U13917 ( .A1(n15849), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n11134) );
  OAI21_X1 U13918 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n15856), .A(n11134), .ZN(
        n11135) );
  AOI21_X1 U13919 ( .B1(n13097), .B2(n11136), .A(n11135), .ZN(n11142) );
  OAI21_X1 U13920 ( .B1(n11139), .B2(n11138), .A(n11137), .ZN(n11140) );
  NAND2_X1 U13921 ( .A1(n13180), .A2(n11140), .ZN(n11141) );
  OAI211_X1 U13922 ( .C1(n11143), .C2(n13146), .A(n11142), .B(n11141), .ZN(
        n11144) );
  AOI21_X1 U13923 ( .B1(n11145), .B2(n13152), .A(n11144), .ZN(n11146) );
  INV_X1 U13924 ( .A(n11146), .ZN(P3_U3184) );
  XOR2_X1 U13925 ( .A(n11148), .B(n11147), .Z(n11160) );
  AOI21_X1 U13926 ( .B1(n11150), .B2(n11149), .A(n6723), .ZN(n11156) );
  AND2_X1 U13927 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n11527) );
  AOI21_X1 U13928 ( .B1(n15849), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n11527), .ZN(
        n11155) );
  NAND2_X1 U13929 ( .A1(n13097), .A2(n11153), .ZN(n11154) );
  OAI211_X1 U13930 ( .C1(n13101), .C2(n11156), .A(n11155), .B(n11154), .ZN(
        n11157) );
  AOI21_X1 U13931 ( .B1(n11158), .B2(n13152), .A(n11157), .ZN(n11159) );
  OAI21_X1 U13932 ( .B1(n11160), .B2(n13146), .A(n11159), .ZN(P3_U3186) );
  INV_X1 U13933 ( .A(n11161), .ZN(n11162) );
  AOI21_X1 U13934 ( .B1(n11164), .B2(n11163), .A(n11162), .ZN(n11172) );
  NAND2_X1 U13935 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n12167)
         );
  OAI21_X1 U13936 ( .B1(n14959), .B2(n12257), .A(n12167), .ZN(n11165) );
  AOI21_X1 U13937 ( .B1(n14962), .B2(n11166), .A(n11165), .ZN(n11171) );
  OAI211_X1 U13938 ( .C1(n11169), .C2(n11168), .A(n11167), .B(n14965), .ZN(
        n11170) );
  OAI211_X1 U13939 ( .C1(n11172), .C2(n12215), .A(n11171), .B(n11170), .ZN(
        P1_U3254) );
  AOI21_X1 U13940 ( .B1(n11174), .B2(n11173), .A(n11298), .ZN(n11190) );
  AOI21_X1 U13941 ( .B1(n11177), .B2(n11176), .A(n11175), .ZN(n11178) );
  NOR2_X1 U13942 ( .A1(n11178), .A2(n13101), .ZN(n11188) );
  NAND3_X1 U13943 ( .A1(n11197), .A2(n11180), .A3(n11179), .ZN(n11181) );
  AOI21_X1 U13944 ( .B1(n11182), .B2(n11181), .A(n13182), .ZN(n11187) );
  NAND2_X1 U13945 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n11770) );
  INV_X1 U13946 ( .A(n11770), .ZN(n11183) );
  AOI21_X1 U13947 ( .B1(n15849), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n11183), .ZN(
        n11184) );
  OAI21_X1 U13948 ( .B1(n13171), .B2(n11185), .A(n11184), .ZN(n11186) );
  NOR3_X1 U13949 ( .A1(n11188), .A2(n11187), .A3(n11186), .ZN(n11189) );
  OAI21_X1 U13950 ( .B1(n11190), .B2(n13146), .A(n11189), .ZN(P3_U3188) );
  INV_X1 U13951 ( .A(n11191), .ZN(n11193) );
  NAND2_X1 U13952 ( .A1(n11193), .A2(n11192), .ZN(n11194) );
  XNOR2_X1 U13953 ( .A(n11195), .B(n11194), .ZN(n11207) );
  XNOR2_X1 U13954 ( .A(n11196), .B(P3_REG1_REG_5__SCAN_IN), .ZN(n11205) );
  OAI21_X1 U13955 ( .B1(P3_REG2_REG_5__SCAN_IN), .B2(n11198), .A(n11197), .ZN(
        n11199) );
  INV_X1 U13956 ( .A(n11199), .ZN(n11201) );
  AND2_X1 U13957 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n11610) );
  AOI21_X1 U13958 ( .B1(n15849), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11610), .ZN(
        n11200) );
  OAI21_X1 U13959 ( .B1(n13182), .B2(n11201), .A(n11200), .ZN(n11204) );
  NOR2_X1 U13960 ( .A1(n13171), .A2(n11202), .ZN(n11203) );
  AOI211_X1 U13961 ( .C1(n13180), .C2(n11205), .A(n11204), .B(n11203), .ZN(
        n11206) );
  OAI21_X1 U13962 ( .B1(n11207), .B2(n13146), .A(n11206), .ZN(P3_U3187) );
  XNOR2_X1 U13963 ( .A(n13819), .B(n11400), .ZN(n15774) );
  AND2_X1 U13964 ( .A1(n14479), .A2(n14425), .ZN(n11208) );
  OAI22_X1 U13965 ( .A1(n15774), .A2(n11208), .B1(n13816), .B2(n14474), .ZN(
        n15777) );
  NAND2_X1 U13966 ( .A1(n11209), .A2(n11400), .ZN(n15775) );
  OAI21_X1 U13967 ( .B1(n15774), .B2(n13811), .A(n15775), .ZN(n11210) );
  NOR2_X1 U13968 ( .A1(n15777), .A2(n11210), .ZN(n15798) );
  NAND2_X1 U13969 ( .A1(n7285), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n11211) );
  OAI21_X1 U13970 ( .B1(n7285), .B2(n15798), .A(n11211), .ZN(P2_U3499) );
  INV_X1 U13971 ( .A(n11212), .ZN(n12226) );
  INV_X1 U13972 ( .A(n11213), .ZN(n11216) );
  OAI222_X1 U13973 ( .A1(P1_U3086), .A2(n12226), .B1(n15438), .B2(n11216), 
        .C1(n11214), .C2(n15435), .ZN(P1_U3339) );
  INV_X1 U13974 ( .A(n15738), .ZN(n11215) );
  OAI222_X1 U13975 ( .A1(n14671), .A2(n11217), .B1(n14663), .B2(n11216), .C1(
        n11215), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U13976 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n12315) );
  MUX2_X1 U13977 ( .A(n12315), .B(P2_REG2_REG_11__SCAN_IN), .S(n11644), .Z(
        n11236) );
  INV_X1 U13978 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n11218) );
  MUX2_X1 U13979 ( .A(n11218), .B(P2_REG2_REG_1__SCAN_IN), .S(n14105), .Z(
        n14112) );
  AND2_X1 U13980 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n14111) );
  NAND2_X1 U13981 ( .A1(n14112), .A2(n14111), .ZN(n14110) );
  INV_X1 U13982 ( .A(n14105), .ZN(n11249) );
  NAND2_X1 U13983 ( .A1(n11249), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n11219) );
  NAND2_X1 U13984 ( .A1(n14110), .A2(n11219), .ZN(n15605) );
  INV_X1 U13985 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n11980) );
  MUX2_X1 U13986 ( .A(n11980), .B(P2_REG2_REG_2__SCAN_IN), .S(n15609), .Z(
        n15606) );
  NAND2_X1 U13987 ( .A1(n15605), .A2(n15606), .ZN(n15604) );
  OR2_X1 U13988 ( .A1(n15609), .A2(n11980), .ZN(n11220) );
  NAND2_X1 U13989 ( .A1(n15604), .A2(n11220), .ZN(n14120) );
  INV_X1 U13990 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n12417) );
  MUX2_X1 U13991 ( .A(n12417), .B(P2_REG2_REG_3__SCAN_IN), .S(n14117), .Z(
        n14121) );
  NAND2_X1 U13992 ( .A1(n14120), .A2(n14121), .ZN(n14119) );
  OR2_X1 U13993 ( .A1(n14117), .A2(n12417), .ZN(n11221) );
  NAND2_X1 U13994 ( .A1(n14119), .A2(n11221), .ZN(n15617) );
  INV_X1 U13995 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n12325) );
  MUX2_X1 U13996 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n12325), .S(n11253), .Z(
        n15618) );
  NAND2_X1 U13997 ( .A1(n15617), .A2(n15618), .ZN(n15616) );
  NAND2_X1 U13998 ( .A1(n11253), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n11222) );
  NAND2_X1 U13999 ( .A1(n15616), .A2(n11222), .ZN(n15630) );
  INV_X1 U14000 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11223) );
  MUX2_X1 U14001 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11223), .S(n11255), .Z(
        n15631) );
  NAND2_X1 U14002 ( .A1(n15630), .A2(n15631), .ZN(n15629) );
  NAND2_X1 U14003 ( .A1(n11255), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n11224) );
  NAND2_X1 U14004 ( .A1(n15629), .A2(n11224), .ZN(n15642) );
  XNOR2_X1 U14005 ( .A(n15646), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n15643) );
  NAND2_X1 U14006 ( .A1(n15642), .A2(n15643), .ZN(n15641) );
  NAND2_X1 U14007 ( .A1(n11257), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n11225) );
  NAND2_X1 U14008 ( .A1(n15641), .A2(n11225), .ZN(n14135) );
  INV_X1 U14009 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11226) );
  XNOR2_X1 U14010 ( .A(n11259), .B(n11226), .ZN(n14136) );
  NAND2_X1 U14011 ( .A1(n14135), .A2(n14136), .ZN(n14134) );
  NAND2_X1 U14012 ( .A1(n11259), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n11227) );
  NAND2_X1 U14013 ( .A1(n14134), .A2(n11227), .ZN(n15655) );
  INV_X1 U14014 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11228) );
  XNOR2_X1 U14015 ( .A(n11262), .B(n11228), .ZN(n15656) );
  NAND2_X1 U14016 ( .A1(n15655), .A2(n15656), .ZN(n15654) );
  NAND2_X1 U14017 ( .A1(n11262), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n11229) );
  NAND2_X1 U14018 ( .A1(n15654), .A2(n11229), .ZN(n15670) );
  MUX2_X1 U14019 ( .A(n12080), .B(P2_REG2_REG_9__SCAN_IN), .S(n11263), .Z(
        n15669) );
  INV_X1 U14020 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n12080) );
  NAND2_X1 U14021 ( .A1(n15676), .A2(n12080), .ZN(n11230) );
  NAND2_X1 U14022 ( .A1(n15672), .A2(n11230), .ZN(n15683) );
  INV_X1 U14023 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11231) );
  XNOR2_X1 U14024 ( .A(n11232), .B(n11231), .ZN(n15684) );
  NAND2_X1 U14025 ( .A1(n15690), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n11233) );
  NAND2_X1 U14026 ( .A1(n15680), .A2(n11233), .ZN(n11235) );
  INV_X1 U14027 ( .A(n11646), .ZN(n11234) );
  AOI21_X1 U14028 ( .B1(n11236), .B2(n11235), .A(n11234), .ZN(n11269) );
  INV_X1 U14029 ( .A(n11237), .ZN(n11241) );
  NAND2_X1 U14030 ( .A1(n11238), .A2(n12037), .ZN(n11239) );
  NAND2_X1 U14031 ( .A1(n11239), .A2(n10184), .ZN(n11240) );
  INV_X1 U14032 ( .A(n11244), .ZN(n11246) );
  OR2_X1 U14033 ( .A1(n10314), .A2(n11242), .ZN(n14665) );
  INV_X1 U14034 ( .A(n14665), .ZN(n11243) );
  AND2_X1 U14035 ( .A1(n11246), .A2(n11243), .ZN(n11264) );
  INV_X1 U14036 ( .A(n14669), .ZN(n14071) );
  INV_X1 U14037 ( .A(n15752), .ZN(n15682) );
  AND2_X1 U14038 ( .A1(n11244), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15600) );
  AND2_X1 U14039 ( .A1(n10314), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11245) );
  NAND2_X1 U14040 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n12137)
         );
  OAI21_X1 U14041 ( .B1(n15749), .B2(n11247), .A(n12137), .ZN(n11267) );
  INV_X1 U14042 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n11248) );
  MUX2_X1 U14043 ( .A(n11248), .B(P2_REG1_REG_1__SCAN_IN), .S(n14105), .Z(
        n14109) );
  AND2_X1 U14044 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n14108) );
  NAND2_X1 U14045 ( .A1(n14109), .A2(n14108), .ZN(n14107) );
  NAND2_X1 U14046 ( .A1(n11249), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n11250) );
  NAND2_X1 U14047 ( .A1(n14107), .A2(n11250), .ZN(n15602) );
  MUX2_X1 U14048 ( .A(n10380), .B(P2_REG1_REG_2__SCAN_IN), .S(n15609), .Z(
        n15603) );
  NAND2_X1 U14049 ( .A1(n15602), .A2(n15603), .ZN(n15601) );
  OR2_X1 U14050 ( .A1(n15609), .A2(n10380), .ZN(n11251) );
  NAND2_X1 U14051 ( .A1(n15601), .A2(n11251), .ZN(n14123) );
  INV_X1 U14052 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n12431) );
  MUX2_X1 U14053 ( .A(n12431), .B(P2_REG1_REG_3__SCAN_IN), .S(n14117), .Z(
        n14124) );
  NAND2_X1 U14054 ( .A1(n14123), .A2(n14124), .ZN(n14122) );
  OR2_X1 U14055 ( .A1(n14117), .A2(n12431), .ZN(n11252) );
  INV_X1 U14056 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n15840) );
  MUX2_X1 U14057 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n15840), .S(n11253), .Z(
        n15615) );
  NAND2_X1 U14058 ( .A1(n11253), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n11254) );
  INV_X1 U14059 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n15842) );
  MUX2_X1 U14060 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n15842), .S(n11255), .Z(
        n15628) );
  NAND2_X1 U14061 ( .A1(n11255), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n11256) );
  NAND2_X1 U14062 ( .A1(n15626), .A2(n11256), .ZN(n15639) );
  INV_X1 U14063 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n15844) );
  MUX2_X1 U14064 ( .A(n15844), .B(P2_REG1_REG_6__SCAN_IN), .S(n15646), .Z(
        n15640) );
  NAND2_X1 U14065 ( .A1(n15639), .A2(n15640), .ZN(n15638) );
  NAND2_X1 U14066 ( .A1(n11257), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n11258) );
  NAND2_X1 U14067 ( .A1(n15638), .A2(n11258), .ZN(n14132) );
  INV_X1 U14068 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n15846) );
  MUX2_X1 U14069 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n15846), .S(n11259), .Z(
        n14133) );
  NAND2_X1 U14070 ( .A1(n14132), .A2(n14133), .ZN(n14131) );
  NAND2_X1 U14071 ( .A1(n11259), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n11260) );
  INV_X1 U14072 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n11261) );
  XNOR2_X1 U14073 ( .A(n11262), .B(n11261), .ZN(n15653) );
  XNOR2_X1 U14074 ( .A(n11263), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n15664) );
  XNOR2_X1 U14075 ( .A(n15690), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n15687) );
  XNOR2_X1 U14076 ( .A(n11644), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n11265) );
  NAND2_X1 U14077 ( .A1(n11264), .A2(n14669), .ZN(n15733) );
  AOI211_X1 U14078 ( .C1(n6527), .C2(n11265), .A(n15733), .B(n11641), .ZN(
        n11266) );
  AOI211_X1 U14079 ( .C1(n15600), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n11267), 
        .B(n11266), .ZN(n11268) );
  OAI21_X1 U14080 ( .B1(n11269), .B2(n15682), .A(n11268), .ZN(P2_U3225) );
  XNOR2_X1 U14081 ( .A(n13761), .B(n11270), .ZN(n11272) );
  NOR2_X1 U14082 ( .A1(n11272), .A2(n11271), .ZN(n13767) );
  AOI21_X1 U14083 ( .B1(n11272), .B2(n11271), .A(n13767), .ZN(n11278) );
  INV_X1 U14084 ( .A(n11273), .ZN(n11789) );
  NAND2_X1 U14085 ( .A1(n11274), .A2(n11789), .ZN(n13768) );
  AOI22_X1 U14086 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(n13768), .B1(n13808), 
        .B2(n10379), .ZN(n11277) );
  AOI22_X1 U14087 ( .A1(n13770), .A2(n13819), .B1(n13769), .B2(n14102), .ZN(
        n11276) );
  OAI211_X1 U14088 ( .C1(n11278), .C2(n13796), .A(n11277), .B(n11276), .ZN(
        P2_U3194) );
  OAI21_X1 U14089 ( .B1(n11280), .B2(n11279), .A(n11329), .ZN(n11281) );
  NAND2_X1 U14090 ( .A1(n11281), .A2(n12832), .ZN(n11285) );
  OAI22_X1 U14091 ( .A1(n15860), .A2(n12836), .B1(n12822), .B2(n7251), .ZN(
        n11282) );
  AOI21_X1 U14092 ( .B1(n11283), .B2(n12803), .A(n11282), .ZN(n11284) );
  OAI211_X1 U14093 ( .C1(n11286), .C2(n15856), .A(n11285), .B(n11284), .ZN(
        P3_U3177) );
  INV_X1 U14094 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n11287) );
  NAND2_X1 U14095 ( .A1(n15752), .A2(n11287), .ZN(n11288) );
  OAI211_X1 U14096 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n15733), .A(n11288), .B(
        n15749), .ZN(n11289) );
  INV_X1 U14097 ( .A(n11289), .ZN(n11291) );
  AOI22_X1 U14098 ( .A1(n15744), .A2(P2_REG1_REG_0__SCAN_IN), .B1(n15752), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n11290) );
  MUX2_X1 U14099 ( .A(n11291), .B(n11290), .S(n10164), .Z(n11293) );
  AOI22_X1 U14100 ( .A1(n15600), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n11292) );
  NAND2_X1 U14101 ( .A1(n11293), .A2(n11292), .ZN(P2_U3214) );
  XNOR2_X1 U14102 ( .A(n11294), .B(P3_REG1_REG_7__SCAN_IN), .ZN(n11306) );
  OAI21_X1 U14103 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(n11295), .A(n11547), .ZN(
        n11304) );
  AND2_X1 U14104 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11811) );
  AOI21_X1 U14105 ( .B1(n15849), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11811), .ZN(
        n11296) );
  OAI21_X1 U14106 ( .B1(n13171), .B2(n11297), .A(n11296), .ZN(n11303) );
  NAND3_X1 U14107 ( .A1(n7432), .A2(n11300), .A3(n11299), .ZN(n11301) );
  AOI21_X1 U14108 ( .B1(n11555), .B2(n11301), .A(n13146), .ZN(n11302) );
  AOI211_X1 U14109 ( .C1(n13097), .C2(n11304), .A(n11303), .B(n11302), .ZN(
        n11305) );
  OAI21_X1 U14110 ( .B1(n11306), .B2(n13101), .A(n11305), .ZN(P3_U3189) );
  XOR2_X1 U14111 ( .A(n11308), .B(n11307), .Z(n11318) );
  AND2_X1 U14112 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n14731) );
  INV_X1 U14113 ( .A(n14731), .ZN(n11309) );
  OAI21_X1 U14114 ( .B1(n14959), .B2(n7568), .A(n11309), .ZN(n11315) );
  NAND2_X1 U14115 ( .A1(n11311), .A2(n11310), .ZN(n11312) );
  AOI21_X1 U14116 ( .B1(n11313), .B2(n11312), .A(n12220), .ZN(n11314) );
  AOI211_X1 U14117 ( .C1(n14962), .C2(n11316), .A(n11315), .B(n11314), .ZN(
        n11317) );
  OAI21_X1 U14118 ( .B1(n12215), .B2(n11318), .A(n11317), .ZN(P1_U3255) );
  INV_X1 U14119 ( .A(n11621), .ZN(n11321) );
  INV_X1 U14120 ( .A(n11319), .ZN(n11322) );
  OAI222_X1 U14121 ( .A1(P1_U3086), .A2(n11321), .B1(n15438), .B2(n11322), 
        .C1(n11320), .C2(n15435), .ZN(P1_U3341) );
  OAI222_X1 U14122 ( .A1(n14671), .A2(n11323), .B1(n14663), .B2(n11322), .C1(
        n14152), .C2(n6510), .ZN(P2_U3313) );
  MUX2_X1 U14123 ( .A(n11325), .B(n11324), .S(n15918), .Z(n11326) );
  OAI21_X1 U14124 ( .B1(n11327), .B2(n13496), .A(n11326), .ZN(P3_U3459) );
  INV_X1 U14125 ( .A(n12839), .ZN(n12536) );
  AND2_X1 U14126 ( .A1(n11329), .A2(n11328), .ZN(n11332) );
  OAI211_X1 U14127 ( .C1(n11332), .C2(n11331), .A(n12832), .B(n11330), .ZN(
        n11337) );
  AOI21_X1 U14128 ( .B1(n12834), .B2(n13040), .A(n11333), .ZN(n11334) );
  OAI21_X1 U14129 ( .B1(n11668), .B2(n12836), .A(n11334), .ZN(n11335) );
  AOI21_X1 U14130 ( .B1(n7250), .B2(n12803), .A(n11335), .ZN(n11336) );
  OAI211_X1 U14131 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12536), .A(n11337), .B(
        n11336), .ZN(P3_U3158) );
  NOR2_X1 U14132 ( .A1(n14035), .A2(n11338), .ZN(n11975) );
  AOI21_X1 U14133 ( .B1(n11338), .B2(n14035), .A(n11975), .ZN(n12040) );
  AOI22_X1 U14134 ( .A1(n14102), .A2(n14449), .B1(n14451), .B2(n13819), .ZN(
        n11342) );
  OAI21_X1 U14135 ( .B1(n11339), .B2(n14035), .A(n11966), .ZN(n11340) );
  NAND2_X1 U14136 ( .A1(n11340), .A2(n15759), .ZN(n11341) );
  OAI211_X1 U14137 ( .C1(n12040), .C2(n14479), .A(n11342), .B(n11341), .ZN(
        n12043) );
  OAI211_X1 U14138 ( .C1(n11364), .C2(n13820), .A(n15767), .B(n11976), .ZN(
        n12042) );
  OAI21_X1 U14139 ( .B1(n12040), .B2(n13811), .A(n12042), .ZN(n11343) );
  NOR2_X1 U14140 ( .A1(n12043), .A2(n11343), .ZN(n11367) );
  INV_X1 U14141 ( .A(n14602), .ZN(n12142) );
  AOI22_X1 U14142 ( .A1(n12142), .A2(n10379), .B1(n7285), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n11344) );
  OAI21_X1 U14143 ( .B1(n11367), .B2(n7285), .A(n11344), .ZN(P2_U3500) );
  NAND2_X1 U14144 ( .A1(n6556), .A2(n11345), .ZN(n11347) );
  XNOR2_X1 U14145 ( .A(n11347), .B(n11346), .ZN(n11352) );
  NAND2_X1 U14146 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14902) );
  OAI21_X1 U14147 ( .B1(n15503), .B2(n11393), .A(n14902), .ZN(n11350) );
  OAI22_X1 U14148 ( .A1(n14825), .A2(n11348), .B1(n11392), .B2(n15508), .ZN(
        n11349) );
  AOI211_X1 U14149 ( .C1(n14773), .C2(n14852), .A(n11350), .B(n11349), .ZN(
        n11351) );
  OAI21_X1 U14150 ( .B1(n11352), .B2(n15496), .A(n11351), .ZN(P1_U3230) );
  XNOR2_X1 U14151 ( .A(n11354), .B(n11353), .ZN(n11355) );
  XNOR2_X1 U14152 ( .A(n11356), .B(n11355), .ZN(n11361) );
  INV_X1 U14153 ( .A(n14825), .ZN(n14707) );
  OAI21_X1 U14154 ( .B1(n15508), .B2(n11494), .A(n11357), .ZN(n11359) );
  OAI22_X1 U14155 ( .A1(n14826), .A2(n11703), .B1(n15563), .B2(n15503), .ZN(
        n11358) );
  AOI211_X1 U14156 ( .C1(n14707), .C2(n14853), .A(n11359), .B(n11358), .ZN(
        n11360) );
  OAI21_X1 U14157 ( .B1(n11361), .B2(n15496), .A(n11360), .ZN(P1_U3227) );
  OAI222_X1 U14158 ( .A1(n13170), .A2(P3_U3151), .B1(n13618), .B2(n11363), 
        .C1(n13622), .C2(n11362), .ZN(P3_U3276) );
  OAI22_X1 U14159 ( .A1(n14652), .A2(n11364), .B1(n15838), .B2(n7881), .ZN(
        n11365) );
  INV_X1 U14160 ( .A(n11365), .ZN(n11366) );
  OAI21_X1 U14161 ( .B1(n11367), .B2(n7304), .A(n11366), .ZN(P2_U3433) );
  OAI21_X1 U14162 ( .B1(n11368), .B2(n11370), .A(n11369), .ZN(n11911) );
  INV_X1 U14163 ( .A(n11911), .ZN(n11374) );
  OAI21_X1 U14164 ( .B1(n11372), .B2(n14037), .A(n11371), .ZN(n11373) );
  AOI222_X1 U14165 ( .A1(n15759), .A2(n11373), .B1(n14100), .B2(n14449), .C1(
        n14102), .C2(n14451), .ZN(n11907) );
  OAI211_X1 U14166 ( .C1(n11977), .C2(n11905), .A(n11714), .B(n12012), .ZN(
        n11906) );
  OAI211_X1 U14167 ( .C1(n15817), .C2(n11374), .A(n11907), .B(n11906), .ZN(
        n11382) );
  INV_X1 U14168 ( .A(n11382), .ZN(n11376) );
  AOI22_X1 U14169 ( .A1(n12142), .A2(n7648), .B1(n7285), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n11375) );
  OAI21_X1 U14170 ( .B1(n11376), .B2(n7285), .A(n11375), .ZN(P2_U3502) );
  INV_X1 U14171 ( .A(n10259), .ZN(n11379) );
  OAI222_X1 U14172 ( .A1(P1_U3086), .A2(n11378), .B1(n15438), .B2(n11379), 
        .C1(n11377), .C2(n15435), .ZN(P1_U3340) );
  INV_X1 U14173 ( .A(n14155), .ZN(n15723) );
  OAI222_X1 U14174 ( .A1(n14671), .A2(n12274), .B1(n14663), .B2(n11379), .C1(
        n15723), .C2(n6510), .ZN(P2_U3312) );
  INV_X1 U14175 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n11380) );
  OAI22_X1 U14176 ( .A1(n14652), .A2(n11905), .B1(n15838), .B2(n11380), .ZN(
        n11381) );
  AOI21_X1 U14177 ( .B1(n11382), .B2(n15838), .A(n11381), .ZN(n11383) );
  INV_X1 U14178 ( .A(n11383), .ZN(P2_U3439) );
  XNOR2_X1 U14179 ( .A(n11385), .B(n6515), .ZN(n15559) );
  OAI21_X1 U14180 ( .B1(n11387), .B2(n6515), .A(n11386), .ZN(n11388) );
  AOI222_X1 U14181 ( .A1(n15545), .A2(n11388), .B1(n14852), .B2(n15256), .C1(
        n14854), .C2(n15257), .ZN(n15558) );
  MUX2_X1 U14182 ( .A(n11389), .B(n15558), .S(n15232), .Z(n11396) );
  OR2_X1 U14183 ( .A1(n11390), .A2(n15138), .ZN(n15236) );
  INV_X1 U14184 ( .A(n15236), .ZN(n15520) );
  AOI21_X1 U14185 ( .B1(n15554), .B2(n11391), .A(n11497), .ZN(n15556) );
  OAI22_X1 U14186 ( .A1(n15517), .A2(n11393), .B1(n15259), .B2(n11392), .ZN(
        n11394) );
  AOI21_X1 U14187 ( .B1(n15520), .B2(n15556), .A(n11394), .ZN(n11395) );
  OAI211_X1 U14188 ( .C1(n15267), .C2(n15559), .A(n11396), .B(n11395), .ZN(
        P1_U3289) );
  NOR2_X1 U14189 ( .A1(n13796), .A2(n15767), .ZN(n13799) );
  INV_X1 U14190 ( .A(n13799), .ZN(n13758) );
  INV_X1 U14191 ( .A(n13819), .ZN(n11397) );
  OAI22_X1 U14192 ( .A1(n13758), .A2(n11397), .B1(n13820), .B2(n13796), .ZN(
        n11399) );
  NAND2_X1 U14193 ( .A1(n11399), .A2(n11398), .ZN(n11402) );
  AOI22_X1 U14194 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(n13768), .B1(n13808), 
        .B2(n11400), .ZN(n11401) );
  OAI211_X1 U14195 ( .C1(n13816), .C2(n13803), .A(n11402), .B(n11401), .ZN(
        P2_U3204) );
  INV_X1 U14196 ( .A(n11403), .ZN(n11414) );
  NAND3_X1 U14197 ( .A1(n13101), .A2(n13182), .A3(n13146), .ZN(n11413) );
  OAI22_X1 U14198 ( .A1(n13144), .A2(n11405), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11404), .ZN(n11412) );
  NAND2_X1 U14199 ( .A1(n13180), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n11408) );
  OR2_X1 U14200 ( .A1(n13182), .A2(n11406), .ZN(n11407) );
  OAI211_X1 U14201 ( .C1(n13146), .C2(n11409), .A(n11408), .B(n11407), .ZN(
        n11410) );
  MUX2_X1 U14202 ( .A(n13152), .B(n11410), .S(n12295), .Z(n11411) );
  AOI211_X1 U14203 ( .C1(n11414), .C2(n11413), .A(n11412), .B(n11411), .ZN(
        n11415) );
  INV_X1 U14204 ( .A(n11415), .ZN(P3_U3182) );
  NAND2_X1 U14205 ( .A1(n14311), .A2(n14100), .ZN(n11418) );
  INV_X1 U14206 ( .A(n11417), .ZN(n11429) );
  NAND2_X1 U14207 ( .A1(n11429), .A2(n11418), .ZN(n11419) );
  XNOR2_X1 U14208 ( .A(n12669), .B(n15813), .ZN(n11708) );
  NAND2_X1 U14209 ( .A1(n14311), .A2(n14099), .ZN(n11709) );
  XNOR2_X1 U14210 ( .A(n11708), .B(n11709), .ZN(n11427) );
  OR2_X1 U14211 ( .A1(n13855), .A2(n14474), .ZN(n11423) );
  NAND2_X1 U14212 ( .A1(n14451), .A2(n14100), .ZN(n11422) );
  NAND2_X1 U14213 ( .A1(n11423), .A2(n11422), .ZN(n11795) );
  AOI22_X1 U14214 ( .A1(n13730), .A2(n11795), .B1(P2_REG3_REG_5__SCAN_IN), 
        .B2(n6510), .ZN(n11425) );
  NAND2_X1 U14215 ( .A1(n13750), .A2(n11801), .ZN(n11424) );
  OAI211_X1 U14216 ( .C1(n13850), .C2(n13733), .A(n11425), .B(n11424), .ZN(
        n11426) );
  INV_X1 U14217 ( .A(n11426), .ZN(n11433) );
  INV_X1 U14218 ( .A(n11427), .ZN(n11431) );
  NAND2_X1 U14219 ( .A1(n13799), .A2(n14100), .ZN(n11428) );
  OAI21_X1 U14220 ( .B1(n11429), .B2(n13796), .A(n11428), .ZN(n11430) );
  NAND3_X1 U14221 ( .A1(n11456), .A2(n11431), .A3(n11430), .ZN(n11432) );
  OAI211_X1 U14222 ( .C1(n11712), .C2(n13796), .A(n11433), .B(n11432), .ZN(
        P2_U3199) );
  XOR2_X1 U14223 ( .A(n11439), .B(n11434), .Z(n15534) );
  INV_X1 U14224 ( .A(n15521), .ZN(n12204) );
  NOR2_X1 U14225 ( .A1(n15535), .A2(n8966), .ZN(n11436) );
  OR2_X1 U14226 ( .A1(n11436), .A2(n11505), .ZN(n15536) );
  INV_X1 U14227 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n14857) );
  OAI22_X1 U14228 ( .A1(n15236), .A2(n15536), .B1(n14857), .B2(n15259), .ZN(
        n11438) );
  NOR2_X1 U14229 ( .A1(n15517), .A2(n15535), .ZN(n11437) );
  AOI211_X1 U14230 ( .C1(n15262), .C2(P1_REG2_REG_1__SCAN_IN), .A(n11438), .B(
        n11437), .ZN(n11445) );
  AOI22_X1 U14231 ( .A1(n15256), .A2(n14855), .B1(n14856), .B2(n15257), .ZN(
        n11443) );
  MUX2_X1 U14232 ( .A(n11440), .B(n11439), .S(n14856), .Z(n11441) );
  NAND2_X1 U14233 ( .A1(n11441), .A2(n15545), .ZN(n11442) );
  OAI211_X1 U14234 ( .C1(n15534), .C2(n11493), .A(n11443), .B(n11442), .ZN(
        n15537) );
  NAND2_X1 U14235 ( .A1(n15537), .A2(n15232), .ZN(n11444) );
  OAI211_X1 U14236 ( .C1(n15534), .C2(n12204), .A(n11445), .B(n11444), .ZN(
        P1_U3292) );
  INV_X1 U14237 ( .A(n11446), .ZN(n11447) );
  OAI222_X1 U14238 ( .A1(n14671), .A2(n7796), .B1(n14663), .B2(n11447), .C1(
        n14159), .C2(P2_U3088), .ZN(P2_U3310) );
  OAI222_X1 U14239 ( .A1(P1_U3086), .A2(n11448), .B1(n15438), .B2(n11447), 
        .C1(n12251), .C2(n15435), .ZN(P1_U3338) );
  INV_X1 U14240 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11449) );
  OAI22_X1 U14241 ( .A1(n15262), .A2(n11450), .B1(n11449), .B2(n15259), .ZN(
        n11452) );
  AOI21_X1 U14242 ( .B1(n15517), .B2(n15236), .A(n8966), .ZN(n11451) );
  AOI211_X1 U14243 ( .C1(n15262), .C2(P1_REG2_REG_0__SCAN_IN), .A(n11452), .B(
        n11451), .ZN(n11455) );
  OR2_X1 U14244 ( .A1(n15262), .A2(n15360), .ZN(n15245) );
  OAI21_X1 U14245 ( .B1(n7490), .B2(n15242), .A(n11453), .ZN(n11454) );
  NAND2_X1 U14246 ( .A1(n11455), .A2(n11454), .ZN(P1_U3293) );
  OAI21_X1 U14247 ( .B1(n11457), .B2(n11459), .A(n11456), .ZN(n11466) );
  AOI22_X1 U14248 ( .A1(n13769), .A2(n14099), .B1(n13750), .B2(n12014), .ZN(
        n11458) );
  NAND2_X1 U14249 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(n6510), .ZN(n15623) );
  OAI211_X1 U14250 ( .C1(n15806), .C2(n13733), .A(n11458), .B(n15623), .ZN(
        n11465) );
  INV_X1 U14251 ( .A(n11459), .ZN(n11461) );
  NAND3_X1 U14252 ( .A1(n11461), .A2(n13799), .A3(n11460), .ZN(n11463) );
  AOI21_X1 U14253 ( .B1(n11463), .B2(n13805), .A(n11462), .ZN(n11464) );
  AOI211_X1 U14254 ( .C1(n13798), .C2(n11466), .A(n11465), .B(n11464), .ZN(
        n11467) );
  INV_X1 U14255 ( .A(n11467), .ZN(P2_U3202) );
  INV_X1 U14256 ( .A(n11468), .ZN(n11475) );
  MUX2_X1 U14257 ( .A(n10761), .B(n11469), .S(n15232), .Z(n11474) );
  INV_X1 U14258 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n12475) );
  OAI22_X1 U14259 ( .A1(n15236), .A2(n11470), .B1(n15259), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n11471) );
  AOI21_X1 U14260 ( .B1(n15239), .B2(n11472), .A(n11471), .ZN(n11473) );
  OAI211_X1 U14261 ( .C1(n11475), .C2(n12204), .A(n11474), .B(n11473), .ZN(
        P1_U3290) );
  XNOR2_X1 U14262 ( .A(n11476), .B(n12879), .ZN(n15882) );
  NAND2_X1 U14263 ( .A1(n15853), .A2(n9778), .ZN(n15850) );
  NOR2_X1 U14264 ( .A1(n15873), .A2(n15850), .ZN(n13212) );
  INV_X1 U14265 ( .A(n13212), .ZN(n11485) );
  INV_X1 U14266 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11482) );
  AOI22_X1 U14267 ( .A1(n13420), .A2(n13040), .B1(n13422), .B2(n9055), .ZN(
        n11480) );
  OAI211_X1 U14268 ( .C1(n11478), .C2(n12879), .A(n11477), .B(n15864), .ZN(
        n11479) );
  OAI211_X1 U14269 ( .C1(n15882), .C2(n15866), .A(n11480), .B(n11479), .ZN(
        n15884) );
  INV_X1 U14270 ( .A(n15884), .ZN(n11481) );
  MUX2_X1 U14271 ( .A(n11482), .B(n11481), .S(n15870), .Z(n11484) );
  AOI22_X1 U14272 ( .A1(n13428), .A2(n7250), .B1(n13427), .B2(n9075), .ZN(
        n11483) );
  OAI211_X1 U14273 ( .C1(n15882), .C2(n11485), .A(n11484), .B(n11483), .ZN(
        P3_U3230) );
  XNOR2_X1 U14274 ( .A(n11486), .B(n11487), .ZN(n15562) );
  XNOR2_X1 U14275 ( .A(n11488), .B(n11487), .ZN(n11491) );
  OAI22_X1 U14276 ( .A1(n11703), .A2(n15227), .B1(n11489), .B2(n15225), .ZN(
        n11490) );
  AOI21_X1 U14277 ( .B1(n11491), .B2(n15545), .A(n11490), .ZN(n11492) );
  OAI21_X1 U14278 ( .B1(n15562), .B2(n11493), .A(n11492), .ZN(n15565) );
  NAND2_X1 U14279 ( .A1(n15565), .A2(n15232), .ZN(n11502) );
  OAI22_X1 U14280 ( .A1(n15232), .A2(n11495), .B1(n11494), .B2(n15259), .ZN(
        n11499) );
  INV_X1 U14281 ( .A(n11571), .ZN(n11496) );
  OAI21_X1 U14282 ( .B1(n15563), .B2(n11497), .A(n11496), .ZN(n15564) );
  NOR2_X1 U14283 ( .A1(n15564), .A2(n15236), .ZN(n11498) );
  AOI211_X1 U14284 ( .C1(n15239), .C2(n11500), .A(n11499), .B(n11498), .ZN(
        n11501) );
  OAI211_X1 U14285 ( .C1(n15562), .C2(n12204), .A(n11502), .B(n11501), .ZN(
        P1_U3288) );
  XNOR2_X1 U14286 ( .A(n11503), .B(n11509), .ZN(n15549) );
  OAI211_X1 U14287 ( .C1(n11505), .C2(n8299), .A(n11504), .B(n15555), .ZN(
        n15543) );
  INV_X1 U14288 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14876) );
  OAI22_X1 U14289 ( .A1(n15067), .A2(n15543), .B1(n14876), .B2(n15259), .ZN(
        n11508) );
  NOR2_X1 U14290 ( .A1(n15232), .A2(n11506), .ZN(n11507) );
  AOI211_X1 U14291 ( .C1(n15232), .C2(n15541), .A(n11508), .B(n11507), .ZN(
        n11512) );
  AOI22_X1 U14292 ( .A1(n7490), .A2(n15546), .B1(n15239), .B2(n6516), .ZN(
        n11511) );
  OAI211_X1 U14293 ( .C1(n15169), .C2(n15549), .A(n11512), .B(n11511), .ZN(
        P1_U3291) );
  NOR2_X1 U14294 ( .A1(n8083), .A2(n11513), .ZN(n11514) );
  XNOR2_X1 U14295 ( .A(n11515), .B(n11514), .ZN(n11520) );
  OAI22_X1 U14296 ( .A1(n15508), .A2(n11573), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11516), .ZN(n11518) );
  OAI22_X1 U14297 ( .A1(n14826), .A2(n11677), .B1(n11564), .B2(n14825), .ZN(
        n11517) );
  AOI211_X1 U14298 ( .C1(n11576), .C2(n14830), .A(n11518), .B(n11517), .ZN(
        n11519) );
  OAI21_X1 U14299 ( .B1(n11520), .B2(n15496), .A(n11519), .ZN(P1_U3239) );
  INV_X1 U14300 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n12259) );
  NAND2_X1 U14301 ( .A1(n13274), .A2(P3_U3897), .ZN(n11521) );
  OAI21_X1 U14302 ( .B1(P3_U3897), .B2(n12259), .A(n11521), .ZN(P3_U3514) );
  INV_X1 U14303 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n12336) );
  NAND2_X1 U14304 ( .A1(n13259), .A2(P3_U3897), .ZN(n11522) );
  OAI21_X1 U14305 ( .B1(P3_U3897), .B2(n12336), .A(n11522), .ZN(P3_U3515) );
  INV_X1 U14306 ( .A(n11523), .ZN(n11524) );
  AOI21_X1 U14307 ( .B1(n11526), .B2(n11525), .A(n11524), .ZN(n11533) );
  AOI21_X1 U14308 ( .B1(n12834), .B2(n13039), .A(n11527), .ZN(n11528) );
  OAI21_X1 U14309 ( .B1(n7251), .B2(n12836), .A(n11528), .ZN(n11530) );
  NOR2_X1 U14310 ( .A1(n12536), .A2(n11632), .ZN(n11529) );
  AOI211_X1 U14311 ( .C1(n12803), .C2(n11531), .A(n11530), .B(n11529), .ZN(
        n11532) );
  OAI21_X1 U14312 ( .B1(n11533), .B2(n12815), .A(n11532), .ZN(P3_U3170) );
  NAND2_X1 U14313 ( .A1(n15866), .A2(n15850), .ZN(n11534) );
  XOR2_X1 U14314 ( .A(n12916), .B(n11535), .Z(n15890) );
  INV_X1 U14315 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11539) );
  OAI21_X1 U14316 ( .B1(n11537), .B2(n9107), .A(n7321), .ZN(n11538) );
  AOI222_X1 U14317 ( .A1(n15864), .A2(n11538), .B1(n13038), .B2(n13420), .C1(
        n13040), .C2(n13422), .ZN(n15891) );
  MUX2_X1 U14318 ( .A(n11539), .B(n15891), .S(n15870), .Z(n11542) );
  INV_X1 U14319 ( .A(n11617), .ZN(n11540) );
  AOI22_X1 U14320 ( .A1(n13428), .A2(n11614), .B1(n13427), .B2(n11540), .ZN(
        n11541) );
  OAI211_X1 U14321 ( .C1(n13431), .C2(n15890), .A(n11542), .B(n11541), .ZN(
        P3_U3228) );
  XNOR2_X1 U14322 ( .A(n11544), .B(n11543), .ZN(n11560) );
  AND3_X1 U14323 ( .A1(n11547), .A2(n11546), .A3(n11545), .ZN(n11548) );
  OAI21_X1 U14324 ( .B1(n11549), .B2(n11548), .A(n13097), .ZN(n11551) );
  NOR2_X1 U14325 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7390), .ZN(n11959) );
  AOI21_X1 U14326 ( .B1(n15849), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11959), .ZN(
        n11550) );
  OAI211_X1 U14327 ( .C1(n13171), .C2(n11552), .A(n11551), .B(n11550), .ZN(
        n11559) );
  INV_X1 U14328 ( .A(n11745), .ZN(n11557) );
  NAND3_X1 U14329 ( .A1(n11555), .A2(n11554), .A3(n11553), .ZN(n11556) );
  AOI21_X1 U14330 ( .B1(n11557), .B2(n11556), .A(n13146), .ZN(n11558) );
  AOI211_X1 U14331 ( .C1(n13180), .C2(n11560), .A(n11559), .B(n11558), .ZN(
        n11561) );
  INV_X1 U14332 ( .A(n11561), .ZN(P3_U3190) );
  XNOR2_X1 U14333 ( .A(n11562), .B(n11563), .ZN(n11566) );
  OAI22_X1 U14334 ( .A1(n11677), .A2(n15227), .B1(n11564), .B2(n15225), .ZN(
        n11565) );
  AOI21_X1 U14335 ( .B1(n11566), .B2(n15545), .A(n11565), .ZN(n11570) );
  XNOR2_X1 U14336 ( .A(n11567), .B(n11568), .ZN(n15575) );
  NAND2_X1 U14337 ( .A1(n15575), .A2(n15552), .ZN(n11569) );
  AND2_X1 U14338 ( .A1(n11570), .A2(n11569), .ZN(n15577) );
  OR2_X1 U14339 ( .A1(n11571), .A2(n15570), .ZN(n11572) );
  NAND2_X1 U14340 ( .A1(n11587), .A2(n11572), .ZN(n15572) );
  OAI22_X1 U14341 ( .A1(n15232), .A2(n11574), .B1(n11573), .B2(n15259), .ZN(
        n11575) );
  AOI21_X1 U14342 ( .B1(n15239), .B2(n11576), .A(n11575), .ZN(n11577) );
  OAI21_X1 U14343 ( .B1(n15236), .B2(n15572), .A(n11577), .ZN(n11578) );
  AOI21_X1 U14344 ( .B1(n15575), .B2(n15521), .A(n11578), .ZN(n11579) );
  OAI21_X1 U14345 ( .B1(n15577), .B2(n15262), .A(n11579), .ZN(P1_U3287) );
  XOR2_X1 U14346 ( .A(n11580), .B(n11581), .Z(n15509) );
  AOI21_X1 U14347 ( .B1(n11582), .B2(n11581), .A(n15360), .ZN(n11585) );
  OAI22_X1 U14348 ( .A1(n11832), .A2(n15227), .B1(n11703), .B2(n15225), .ZN(
        n11583) );
  AOI21_X1 U14349 ( .B1(n11585), .B2(n11584), .A(n11583), .ZN(n15510) );
  AOI21_X1 U14350 ( .B1(n11700), .B2(n11587), .A(n11586), .ZN(n15519) );
  AOI22_X1 U14351 ( .A1(n15519), .A2(n15555), .B1(n15580), .B2(n11700), .ZN(
        n11588) );
  OAI211_X1 U14352 ( .C1(n15509), .C2(n15560), .A(n15510), .B(n11588), .ZN(
        n11590) );
  NAND2_X1 U14353 ( .A1(n11590), .A2(n15588), .ZN(n11589) );
  OAI21_X1 U14354 ( .B1(n15588), .B2(n8337), .A(n11589), .ZN(P1_U3480) );
  NAND2_X1 U14355 ( .A1(n11590), .A2(n15599), .ZN(n11591) );
  OAI21_X1 U14356 ( .B1(n15599), .B2(n11592), .A(n11591), .ZN(P1_U3535) );
  INV_X1 U14357 ( .A(n11593), .ZN(n11594) );
  AOI211_X1 U14358 ( .C1(n11596), .C2(n11595), .A(n12215), .B(n11594), .ZN(
        n11606) );
  INV_X1 U14359 ( .A(n11597), .ZN(n11598) );
  AOI211_X1 U14360 ( .C1(n11600), .C2(n11599), .A(n12220), .B(n11598), .ZN(
        n11605) );
  NAND2_X1 U14361 ( .A1(n14962), .A2(n11601), .ZN(n11602) );
  NAND2_X1 U14362 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n14784)
         );
  OAI211_X1 U14363 ( .C1(n11603), .C2(n14959), .A(n11602), .B(n14784), .ZN(
        n11604) );
  OR3_X1 U14364 ( .A1(n11606), .A2(n11605), .A3(n11604), .ZN(P1_U3256) );
  OAI21_X1 U14365 ( .B1(n11608), .B2(n11607), .A(n11766), .ZN(n11609) );
  NAND2_X1 U14366 ( .A1(n11609), .A2(n12832), .ZN(n11616) );
  AOI21_X1 U14367 ( .B1(n12834), .B2(n13038), .A(n11610), .ZN(n11611) );
  OAI21_X1 U14368 ( .B1(n11612), .B2(n12836), .A(n11611), .ZN(n11613) );
  AOI21_X1 U14369 ( .B1(n11614), .B2(n12803), .A(n11613), .ZN(n11615) );
  OAI211_X1 U14370 ( .C1(n11617), .C2(n12536), .A(n11616), .B(n11615), .ZN(
        P3_U3167) );
  OAI21_X1 U14371 ( .B1(n11620), .B2(n11619), .A(n11618), .ZN(n11625) );
  NAND2_X1 U14372 ( .A1(n11621), .A2(n14962), .ZN(n11622) );
  NAND2_X1 U14373 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n14686)
         );
  OAI211_X1 U14374 ( .C1(n11623), .C2(n14959), .A(n11622), .B(n14686), .ZN(
        n11624) );
  AOI21_X1 U14375 ( .B1(n11625), .B2(n14954), .A(n11624), .ZN(n11630) );
  OAI211_X1 U14376 ( .C1(n11628), .C2(n11627), .A(n11626), .B(n14965), .ZN(
        n11629) );
  NAND2_X1 U14377 ( .A1(n11630), .A2(n11629), .ZN(P1_U3257) );
  XNOR2_X1 U14378 ( .A(n11631), .B(n12905), .ZN(n15887) );
  INV_X1 U14379 ( .A(n15887), .ZN(n11639) );
  OAI22_X1 U14380 ( .A1(n13266), .A2(n15885), .B1(n11632), .B2(n15855), .ZN(
        n11638) );
  AOI22_X1 U14381 ( .A1(n13420), .A2(n13039), .B1(n13422), .B2(n13041), .ZN(
        n11636) );
  OAI211_X1 U14382 ( .C1(n11634), .C2(n12905), .A(n11633), .B(n15864), .ZN(
        n11635) );
  OAI211_X1 U14383 ( .C1(n15887), .C2(n15866), .A(n11636), .B(n11635), .ZN(
        n15889) );
  MUX2_X1 U14384 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n15889), .S(n15870), .Z(
        n11637) );
  AOI211_X1 U14385 ( .C1(n11639), .C2(n13212), .A(n11638), .B(n11637), .ZN(
        n11640) );
  INV_X1 U14386 ( .A(n11640), .ZN(P3_U3229) );
  XNOR2_X1 U14387 ( .A(n14149), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n11643) );
  XOR2_X1 U14388 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n15701), .Z(n15699) );
  OAI21_X1 U14389 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n15701), .A(n15697), 
        .ZN(n11642) );
  NOR2_X1 U14390 ( .A1(n11642), .A2(n11643), .ZN(n14140) );
  AOI211_X1 U14391 ( .C1(n11643), .C2(n11642), .A(n15733), .B(n14140), .ZN(
        n11655) );
  OR2_X1 U14392 ( .A1(n11644), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n11645) );
  NAND2_X1 U14393 ( .A1(n11646), .A2(n11645), .ZN(n15695) );
  INV_X1 U14394 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n14456) );
  MUX2_X1 U14395 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n14456), .S(n15701), .Z(
        n15696) );
  NAND2_X1 U14396 ( .A1(n15695), .A2(n15696), .ZN(n15694) );
  OR2_X1 U14397 ( .A1(n15701), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n11647) );
  INV_X1 U14398 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11648) );
  XNOR2_X1 U14399 ( .A(n14149), .B(n11648), .ZN(n11649) );
  NAND2_X1 U14400 ( .A1(n11650), .A2(n11649), .ZN(n14151) );
  OAI211_X1 U14401 ( .C1(n11650), .C2(n11649), .A(n14151), .B(n15752), .ZN(
        n11653) );
  INV_X1 U14402 ( .A(n15749), .ZN(n15739) );
  AND2_X1 U14403 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n11651) );
  AOI21_X1 U14404 ( .B1(n15739), .B2(n14149), .A(n11651), .ZN(n11652) );
  OAI211_X1 U14405 ( .C1(n7734), .C2(n15755), .A(n11653), .B(n11652), .ZN(
        n11654) );
  OR2_X1 U14406 ( .A1(n11655), .A2(n11654), .ZN(P2_U3227) );
  INV_X1 U14407 ( .A(n14170), .ZN(n15748) );
  OAI222_X1 U14408 ( .A1(n14671), .A2(n11656), .B1(n14663), .B2(n11658), .C1(
        n15748), .C2(n11242), .ZN(P2_U3309) );
  INV_X1 U14409 ( .A(n14961), .ZN(n11659) );
  OAI222_X1 U14410 ( .A1(P1_U3086), .A2(n11659), .B1(n15438), .B2(n11658), 
        .C1(n11657), .C2(n15435), .ZN(P1_U3337) );
  XNOR2_X1 U14411 ( .A(n11660), .B(n12897), .ZN(n15876) );
  AOI22_X1 U14412 ( .A1(n13411), .A2(n15876), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n13427), .ZN(n11671) );
  NOR2_X1 U14413 ( .A1(n15901), .A2(n11661), .ZN(n15875) );
  NAND2_X1 U14414 ( .A1(n15864), .A2(n11662), .ZN(n11663) );
  OAI21_X1 U14415 ( .B1(n11663), .B2(n11660), .A(n15861), .ZN(n11664) );
  NAND2_X1 U14416 ( .A1(n11664), .A2(n13044), .ZN(n11667) );
  NAND3_X1 U14417 ( .A1(n11660), .A2(n15864), .A3(n11665), .ZN(n11666) );
  OAI211_X1 U14418 ( .C1(n11668), .C2(n15859), .A(n11667), .B(n11666), .ZN(
        n15874) );
  AOI21_X1 U14419 ( .B1(n15875), .B2(n13023), .A(n15874), .ZN(n11669) );
  MUX2_X1 U14420 ( .A(n11669), .B(n7400), .S(n15873), .Z(n11670) );
  NAND2_X1 U14421 ( .A1(n11671), .A2(n11670), .ZN(P3_U3232) );
  XNOR2_X1 U14422 ( .A(n11672), .B(n11673), .ZN(n15579) );
  INV_X1 U14423 ( .A(n15579), .ZN(n11686) );
  OAI211_X1 U14424 ( .C1(n11676), .C2(n11675), .A(n11674), .B(n15545), .ZN(
        n11679) );
  OAI22_X1 U14425 ( .A1(n11677), .A2(n15225), .B1(n12183), .B2(n15227), .ZN(
        n11866) );
  INV_X1 U14426 ( .A(n11866), .ZN(n11678) );
  NAND2_X1 U14427 ( .A1(n11679), .A2(n11678), .ZN(n15586) );
  AOI21_X1 U14428 ( .B1(n7857), .B2(n15581), .A(n15571), .ZN(n11680) );
  NAND2_X1 U14429 ( .A1(n11680), .A2(n11834), .ZN(n15583) );
  OAI22_X1 U14430 ( .A1(n15232), .A2(n11681), .B1(n11868), .B2(n15259), .ZN(
        n11682) );
  AOI21_X1 U14431 ( .B1(n15239), .B2(n15581), .A(n11682), .ZN(n11683) );
  OAI21_X1 U14432 ( .B1(n15583), .B2(n15067), .A(n11683), .ZN(n11684) );
  AOI21_X1 U14433 ( .B1(n15586), .B2(n15232), .A(n11684), .ZN(n11685) );
  OAI21_X1 U14434 ( .B1(n11686), .B2(n15267), .A(n11685), .ZN(P1_U3285) );
  AOI21_X1 U14435 ( .B1(n11687), .B2(n12918), .A(n13401), .ZN(n11691) );
  OAI22_X1 U14436 ( .A1(n15861), .A2(n11772), .B1(n6954), .B2(n15859), .ZN(
        n11690) );
  AOI21_X1 U14437 ( .B1(n11691), .B2(n11689), .A(n11690), .ZN(n15895) );
  XNOR2_X1 U14438 ( .A(n11692), .B(n12918), .ZN(n15898) );
  NOR2_X1 U14439 ( .A1(n15870), .A2(n9643), .ZN(n11694) );
  OAI22_X1 U14440 ( .A1(n13266), .A2(n15896), .B1(n11777), .B2(n15855), .ZN(
        n11693) );
  AOI211_X1 U14441 ( .C1(n15898), .C2(n13411), .A(n11694), .B(n11693), .ZN(
        n11695) );
  OAI21_X1 U14442 ( .B1(n15895), .B2(n15873), .A(n11695), .ZN(P3_U3227) );
  INV_X1 U14443 ( .A(n11696), .ZN(n11697) );
  OAI222_X1 U14444 ( .A1(n11699), .A2(P3_U3151), .B1(n13618), .B2(n11698), 
        .C1(n13622), .C2(n11697), .ZN(P3_U3275) );
  INV_X1 U14445 ( .A(n11700), .ZN(n15516) );
  OAI211_X1 U14446 ( .C1(n6715), .C2(n11702), .A(n11701), .B(n14813), .ZN(
        n11707) );
  NOR2_X1 U14447 ( .A1(n15508), .A2(n15512), .ZN(n11705) );
  OAI22_X1 U14448 ( .A1(n14826), .A2(n11832), .B1(n11703), .B2(n14825), .ZN(
        n11704) );
  AOI211_X1 U14449 ( .C1(P1_REG3_REG_7__SCAN_IN), .C2(P1_U3086), .A(n11705), 
        .B(n11704), .ZN(n11706) );
  OAI211_X1 U14450 ( .C1(n15516), .C2(n15503), .A(n11707), .B(n11706), .ZN(
        P1_U3213) );
  INV_X1 U14451 ( .A(n11708), .ZN(n11710) );
  NAND2_X1 U14452 ( .A1(n11710), .A2(n11709), .ZN(n11711) );
  INV_X2 U14453 ( .A(n11713), .ZN(n12669) );
  XNOR2_X1 U14454 ( .A(n15764), .B(n12669), .ZN(n11723) );
  NOR2_X1 U14455 ( .A1(n13855), .A2(n11714), .ZN(n11715) );
  NAND2_X1 U14456 ( .A1(n11723), .A2(n11715), .ZN(n11725) );
  OR2_X1 U14457 ( .A1(n11723), .A2(n11715), .ZN(n11716) );
  NAND2_X1 U14458 ( .A1(n11725), .A2(n11716), .ZN(n11761) );
  XNOR2_X1 U14459 ( .A(n13858), .B(n12669), .ZN(n11718) );
  NOR2_X1 U14460 ( .A1(n13859), .A2(n15767), .ZN(n11719) );
  NAND2_X1 U14461 ( .A1(n11718), .A2(n11719), .ZN(n12118) );
  INV_X1 U14462 ( .A(n11718), .ZN(n12713) );
  INV_X1 U14463 ( .A(n11719), .ZN(n11720) );
  NAND2_X1 U14464 ( .A1(n12713), .A2(n11720), .ZN(n11721) );
  AND2_X1 U14465 ( .A1(n12118), .A2(n11721), .ZN(n11726) );
  INV_X1 U14466 ( .A(n11726), .ZN(n11722) );
  AOI21_X1 U14467 ( .B1(n11758), .B2(n11722), .A(n13796), .ZN(n11729) );
  INV_X1 U14468 ( .A(n11723), .ZN(n11724) );
  NOR3_X1 U14469 ( .A1(n13758), .A2(n13855), .A3(n11724), .ZN(n11728) );
  OAI21_X1 U14470 ( .B1(n11729), .B2(n11728), .A(n12712), .ZN(n11735) );
  OR2_X1 U14471 ( .A1(n13855), .A2(n14472), .ZN(n11731) );
  NAND2_X1 U14472 ( .A1(n14449), .A2(n14096), .ZN(n11730) );
  NAND2_X1 U14473 ( .A1(n11731), .A2(n11730), .ZN(n11932) );
  INV_X1 U14474 ( .A(n11932), .ZN(n11732) );
  OAI22_X1 U14475 ( .A1(n13789), .A2(n11732), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12308), .ZN(n11733) );
  AOI21_X1 U14476 ( .B1(n11937), .B2(n13750), .A(n11733), .ZN(n11734) );
  OAI211_X1 U14477 ( .C1(n7911), .C2(n13733), .A(n11735), .B(n11734), .ZN(
        P2_U3185) );
  XNOR2_X1 U14478 ( .A(n11736), .B(P3_REG1_REG_9__SCAN_IN), .ZN(n11750) );
  OAI21_X1 U14479 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n11737), .A(n11891), .ZN(
        n11742) );
  NAND2_X1 U14480 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n11821) );
  INV_X1 U14481 ( .A(n11821), .ZN(n11738) );
  AOI21_X1 U14482 ( .B1(n15849), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11738), .ZN(
        n11739) );
  OAI21_X1 U14483 ( .B1(n13171), .B2(n11740), .A(n11739), .ZN(n11741) );
  AOI21_X1 U14484 ( .B1(n11742), .B2(n13097), .A(n11741), .ZN(n11749) );
  INV_X1 U14485 ( .A(n11899), .ZN(n11747) );
  NOR3_X1 U14486 ( .A1(n11745), .A2(n11744), .A3(n11743), .ZN(n11746) );
  OAI21_X1 U14487 ( .B1(n11747), .B2(n11746), .A(n13173), .ZN(n11748) );
  OAI211_X1 U14488 ( .C1(n11750), .C2(n13101), .A(n11749), .B(n11748), .ZN(
        P3_U3191) );
  INV_X1 U14489 ( .A(SI_21_), .ZN(n11752) );
  OAI222_X1 U14490 ( .A1(P3_U3151), .A2(n11753), .B1(n13618), .B2(n11752), 
        .C1(n13622), .C2(n11751), .ZN(P3_U3274) );
  INV_X1 U14491 ( .A(n15761), .ZN(n11757) );
  OR2_X1 U14492 ( .A1(n13859), .A2(n14474), .ZN(n11755) );
  NAND2_X1 U14493 ( .A1(n14451), .A2(n14099), .ZN(n11754) );
  NAND2_X1 U14494 ( .A1(n11755), .A2(n11754), .ZN(n15758) );
  AOI22_X1 U14495 ( .A1(n13730), .A2(n15758), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11756) );
  OAI21_X1 U14496 ( .B1(n13804), .B2(n11757), .A(n11756), .ZN(n11763) );
  INV_X1 U14497 ( .A(n11758), .ZN(n11759) );
  AOI211_X1 U14498 ( .C1(n11761), .C2(n11760), .A(n13796), .B(n11759), .ZN(
        n11762) );
  AOI211_X1 U14499 ( .C1(n15764), .C2(n13808), .A(n11763), .B(n11762), .ZN(
        n11764) );
  INV_X1 U14500 ( .A(n11764), .ZN(P2_U3211) );
  AND2_X1 U14501 ( .A1(n11766), .A2(n11765), .ZN(n11769) );
  XOR2_X1 U14502 ( .A(n13038), .B(n11767), .Z(n11768) );
  NAND2_X1 U14503 ( .A1(n11769), .A2(n11768), .ZN(n11810) );
  OAI211_X1 U14504 ( .C1(n11769), .C2(n11768), .A(n11810), .B(n12832), .ZN(
        n11776) );
  NAND2_X1 U14505 ( .A1(n12834), .A2(n13037), .ZN(n11771) );
  OAI211_X1 U14506 ( .C1(n11772), .C2(n12836), .A(n11771), .B(n11770), .ZN(
        n11773) );
  AOI21_X1 U14507 ( .B1(n12803), .B2(n11774), .A(n11773), .ZN(n11775) );
  OAI211_X1 U14508 ( .C1(n11777), .C2(n12536), .A(n11776), .B(n11775), .ZN(
        P3_U3179) );
  NAND2_X1 U14509 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n14103), .ZN(n11778) );
  OAI21_X1 U14510 ( .B1(n14059), .B2(n14103), .A(n11778), .ZN(P2_U3560) );
  INV_X1 U14511 ( .A(n11779), .ZN(n11781) );
  OAI222_X1 U14512 ( .A1(n15435), .A2(n11780), .B1(n15438), .B2(n11781), .C1(
        P1_U3086), .C2(n15163), .ZN(P1_U3336) );
  OAI222_X1 U14513 ( .A1(n14671), .A2(n11782), .B1(n14673), .B2(n11781), .C1(
        n14076), .C2(n11242), .ZN(P2_U3308) );
  OAI222_X1 U14514 ( .A1(n15435), .A2(n11783), .B1(n15438), .B2(n11913), .C1(
        n8970), .C2(P1_U3086), .ZN(P1_U3334) );
  NOR2_X1 U14515 ( .A1(n7909), .A2(n11786), .ZN(n14039) );
  XNOR2_X1 U14516 ( .A(n11784), .B(n14039), .ZN(n15818) );
  INV_X1 U14517 ( .A(n11787), .ZN(n11788) );
  NAND3_X1 U14518 ( .A1(n11789), .A2(n15792), .A3(n11788), .ZN(n11790) );
  INV_X1 U14519 ( .A(n15780), .ZN(n11792) );
  NAND2_X1 U14520 ( .A1(n14479), .A2(n11792), .ZN(n11793) );
  XNOR2_X1 U14521 ( .A(n11794), .B(n14039), .ZN(n11796) );
  AOI21_X1 U14522 ( .B1(n11796), .B2(n15759), .A(n11795), .ZN(n15821) );
  MUX2_X1 U14523 ( .A(n11223), .B(n15821), .S(n15781), .Z(n11805) );
  NAND2_X1 U14524 ( .A1(n12013), .A2(n15813), .ZN(n11798) );
  NAND2_X1 U14525 ( .A1(n11798), .A2(n15767), .ZN(n11799) );
  NOR2_X1 U14526 ( .A1(n11797), .A2(n11799), .ZN(n15814) );
  INV_X1 U14527 ( .A(n11801), .ZN(n11802) );
  OAI22_X1 U14528 ( .A1(n14436), .A2(n13850), .B1(n15776), .B2(n11802), .ZN(
        n11803) );
  AOI21_X1 U14529 ( .B1(n15770), .B2(n15814), .A(n11803), .ZN(n11804) );
  OAI211_X1 U14530 ( .C1(n15818), .C2(n14421), .A(n11805), .B(n11804), .ZN(
        P2_U3260) );
  INV_X1 U14531 ( .A(n11806), .ZN(n11808) );
  OAI22_X1 U14532 ( .A1(n13028), .A2(P3_U3151), .B1(SI_22_), .B2(n13618), .ZN(
        n11807) );
  AOI21_X1 U14533 ( .B1(n11808), .B2(n11928), .A(n11807), .ZN(P3_U3273) );
  NAND2_X1 U14534 ( .A1(n11810), .A2(n11809), .ZN(n11956) );
  XNOR2_X1 U14535 ( .A(n11956), .B(n11955), .ZN(n11817) );
  AOI21_X1 U14536 ( .B1(n12834), .B2(n13036), .A(n11811), .ZN(n11812) );
  OAI21_X1 U14537 ( .B1(n6952), .B2(n12836), .A(n11812), .ZN(n11814) );
  NOR2_X1 U14538 ( .A1(n12536), .A2(n11844), .ZN(n11813) );
  AOI211_X1 U14539 ( .C1(n12803), .C2(n11815), .A(n11814), .B(n11813), .ZN(
        n11816) );
  OAI21_X1 U14540 ( .B1(n11817), .B2(n12815), .A(n11816), .ZN(P3_U3153) );
  INV_X1 U14541 ( .A(n11854), .ZN(n11818) );
  AOI21_X1 U14542 ( .B1(n11820), .B2(n11819), .A(n11818), .ZN(n11826) );
  INV_X1 U14543 ( .A(n11950), .ZN(n11989) );
  NAND2_X1 U14544 ( .A1(n12834), .A2(n13423), .ZN(n11822) );
  OAI211_X1 U14545 ( .C1(n11944), .C2(n12836), .A(n11822), .B(n11821), .ZN(
        n11824) );
  NOR2_X1 U14546 ( .A1(n12536), .A2(n11949), .ZN(n11823) );
  AOI211_X1 U14547 ( .C1(n12803), .C2(n11989), .A(n11824), .B(n11823), .ZN(
        n11825) );
  OAI21_X1 U14548 ( .B1(n11826), .B2(n12815), .A(n11825), .ZN(P3_U3171) );
  INV_X1 U14549 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11829) );
  INV_X1 U14550 ( .A(n11827), .ZN(n11916) );
  OAI222_X1 U14551 ( .A1(n15435), .A2(n11829), .B1(n15438), .B2(n11916), .C1(
        n11828), .C2(P1_U3086), .ZN(P1_U3335) );
  OAI21_X1 U14552 ( .B1(n11831), .B2(n6959), .A(n11830), .ZN(n11833) );
  OAI22_X1 U14553 ( .A1(n12169), .A2(n15227), .B1(n11832), .B2(n15225), .ZN(
        n12062) );
  AOI21_X1 U14554 ( .B1(n11833), .B2(n15545), .A(n12062), .ZN(n15398) );
  AOI211_X1 U14555 ( .C1(n15396), .C2(n11834), .A(n15571), .B(n11920), .ZN(
        n15395) );
  INV_X1 U14556 ( .A(n12065), .ZN(n11835) );
  AOI22_X1 U14557 ( .A1(n15262), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n11835), 
        .B2(n15513), .ZN(n11836) );
  OAI21_X1 U14558 ( .B1(n11837), .B2(n15517), .A(n11836), .ZN(n11841) );
  XOR2_X1 U14559 ( .A(n11838), .B(n11839), .Z(n15399) );
  NOR2_X1 U14560 ( .A1(n15399), .A2(n15169), .ZN(n11840) );
  AOI211_X1 U14561 ( .C1(n15395), .C2(n15254), .A(n11841), .B(n11840), .ZN(
        n11842) );
  OAI21_X1 U14562 ( .B1(n15262), .B2(n15398), .A(n11842), .ZN(P1_U3284) );
  XNOR2_X1 U14563 ( .A(n11843), .B(n12884), .ZN(n15900) );
  OAI22_X1 U14564 ( .A1(n13266), .A2(n6956), .B1(n11844), .B2(n15855), .ZN(
        n11851) );
  NAND3_X1 U14565 ( .A1(n11689), .A2(n12924), .A3(n11845), .ZN(n11846) );
  NAND3_X1 U14566 ( .A1(n7324), .A2(n15864), .A3(n11846), .ZN(n11849) );
  AOI22_X1 U14567 ( .A1(n13420), .A2(n13036), .B1(n13422), .B2(n13038), .ZN(
        n11848) );
  NAND2_X1 U14568 ( .A1(n11849), .A2(n11848), .ZN(n15904) );
  MUX2_X1 U14569 ( .A(n15904), .B(P3_REG2_REG_7__SCAN_IN), .S(n15873), .Z(
        n11850) );
  AOI211_X1 U14570 ( .C1(n13411), .C2(n15900), .A(n11851), .B(n11850), .ZN(
        n11852) );
  INV_X1 U14571 ( .A(n11852), .ZN(P3_U3226) );
  AND2_X1 U14572 ( .A1(n11854), .A2(n11853), .ZN(n11857) );
  OAI211_X1 U14573 ( .C1(n11857), .C2(n11856), .A(n12832), .B(n11855), .ZN(
        n11861) );
  NAND2_X1 U14574 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n11887)
         );
  OAI21_X1 U14575 ( .B1(n12836), .B2(n12148), .A(n11887), .ZN(n11859) );
  NOR2_X1 U14576 ( .A1(n12842), .A2(n13598), .ZN(n11858) );
  AOI211_X1 U14577 ( .C1(n12834), .C2(n13034), .A(n11859), .B(n11858), .ZN(
        n11860) );
  OAI211_X1 U14578 ( .C1(n12153), .C2(n12536), .A(n11861), .B(n11860), .ZN(
        P3_U3157) );
  INV_X1 U14579 ( .A(n11862), .ZN(n11863) );
  AOI21_X1 U14580 ( .B1(n11865), .B2(n11864), .A(n11863), .ZN(n11871) );
  AOI22_X1 U14581 ( .A1(n15500), .A2(n11866), .B1(P1_REG3_REG_8__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11867) );
  OAI21_X1 U14582 ( .B1(n11868), .B2(n15508), .A(n11867), .ZN(n11869) );
  AOI21_X1 U14583 ( .B1(n15581), .B2(n14830), .A(n11869), .ZN(n11870) );
  OAI21_X1 U14584 ( .B1(n11871), .B2(n15496), .A(n11870), .ZN(P1_U3221) );
  OAI222_X1 U14585 ( .A1(n14671), .A2(n11873), .B1(n6510), .B2(n13812), .C1(
        n14673), .C2(n11872), .ZN(P2_U3305) );
  XOR2_X1 U14586 ( .A(n11875), .B(n11874), .Z(n11884) );
  XNOR2_X1 U14587 ( .A(n11877), .B(n11876), .ZN(n11878) );
  NAND2_X1 U14588 ( .A1(n11878), .A2(n14954), .ZN(n11883) );
  AND2_X1 U14589 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14828) );
  NOR2_X1 U14590 ( .A1(n14959), .A2(n11879), .ZN(n11880) );
  AOI211_X1 U14591 ( .C1(n14962), .C2(n11881), .A(n14828), .B(n11880), .ZN(
        n11882) );
  OAI211_X1 U14592 ( .C1(n11884), .C2(n12220), .A(n11883), .B(n11882), .ZN(
        P1_U3258) );
  XOR2_X1 U14593 ( .A(n11885), .B(n11886), .Z(n11904) );
  NAND2_X1 U14594 ( .A1(n15849), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n11888) );
  NAND2_X1 U14595 ( .A1(n11888), .A2(n11887), .ZN(n11895) );
  NAND3_X1 U14596 ( .A1(n11891), .A2(n11890), .A3(n11889), .ZN(n11892) );
  AOI21_X1 U14597 ( .B1(n11893), .B2(n11892), .A(n13182), .ZN(n11894) );
  AOI211_X1 U14598 ( .C1(n13152), .C2(n11896), .A(n11895), .B(n11894), .ZN(
        n11903) );
  AND3_X1 U14599 ( .A1(n11899), .A2(n11898), .A3(n11897), .ZN(n11900) );
  OAI21_X1 U14600 ( .B1(n11901), .B2(n11900), .A(n13173), .ZN(n11902) );
  OAI211_X1 U14601 ( .C1(n11904), .C2(n13101), .A(n11903), .B(n11902), .ZN(
        P3_U3192) );
  OAI22_X1 U14602 ( .A1(n14461), .A2(n11906), .B1(n11905), .B2(n14436), .ZN(
        n11910) );
  OAI21_X1 U14603 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n15776), .A(n11907), .ZN(
        n11908) );
  MUX2_X1 U14604 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11908), .S(n15781), .Z(
        n11909) );
  AOI211_X1 U14605 ( .C1(n15771), .C2(n11911), .A(n11910), .B(n11909), .ZN(
        n11912) );
  INV_X1 U14606 ( .A(n11912), .ZN(P2_U3262) );
  OAI222_X1 U14607 ( .A1(n14671), .A2(n12484), .B1(n11242), .B2(n14077), .C1(
        n14673), .C2(n11913), .ZN(P2_U3306) );
  INV_X1 U14608 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n12272) );
  INV_X1 U14609 ( .A(n12868), .ZN(n11914) );
  NAND2_X1 U14610 ( .A1(n11914), .A2(P3_U3897), .ZN(n11915) );
  OAI21_X1 U14611 ( .B1(P3_U3897), .B2(n12272), .A(n11915), .ZN(P3_U3520) );
  OAI222_X1 U14612 ( .A1(n14671), .A2(n12359), .B1(P2_U3088), .B2(n14075), 
        .C1(n14673), .C2(n11916), .ZN(P2_U3307) );
  XNOR2_X1 U14613 ( .A(n11917), .B(n8049), .ZN(n15394) );
  OAI211_X1 U14614 ( .C1(n6709), .C2(n8049), .A(n15545), .B(n11918), .ZN(
        n15393) );
  INV_X1 U14615 ( .A(n15393), .ZN(n11919) );
  NOR2_X1 U14616 ( .A1(n12183), .A2(n15225), .ZN(n15390) );
  OAI21_X1 U14617 ( .B1(n11919), .B2(n15390), .A(n15232), .ZN(n11927) );
  OAI211_X1 U14618 ( .C1(n11920), .C2(n11922), .A(n11996), .B(n15555), .ZN(
        n11921) );
  OAI21_X1 U14619 ( .B1(n14729), .B2(n15227), .A(n11921), .ZN(n15389) );
  NOR2_X1 U14620 ( .A1(n11922), .A2(n15517), .ZN(n11925) );
  OAI22_X1 U14621 ( .A1(n15232), .A2(n11923), .B1(n12182), .B2(n15259), .ZN(
        n11924) );
  AOI211_X1 U14622 ( .C1(n15389), .C2(n15254), .A(n11925), .B(n11924), .ZN(
        n11926) );
  OAI211_X1 U14623 ( .C1(n15394), .C2(n15267), .A(n11927), .B(n11926), .ZN(
        P1_U3283) );
  INV_X1 U14624 ( .A(SI_23_), .ZN(n12451) );
  NAND2_X1 U14625 ( .A1(n11929), .A2(n11928), .ZN(n11930) );
  OAI211_X1 U14626 ( .C1(n12451), .C2(n13618), .A(n11930), .B(n13031), .ZN(
        P3_U3272) );
  INV_X1 U14627 ( .A(n11934), .ZN(n14042) );
  XNOR2_X1 U14628 ( .A(n11931), .B(n14042), .ZN(n11933) );
  AOI21_X1 U14629 ( .B1(n11933), .B2(n15759), .A(n11932), .ZN(n15832) );
  XNOR2_X1 U14630 ( .A(n11935), .B(n11934), .ZN(n15836) );
  OAI211_X1 U14631 ( .C1(n11936), .C2(n7911), .A(n15767), .B(n12054), .ZN(
        n15830) );
  AOI22_X1 U14632 ( .A1(n15783), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n11937), 
        .B2(n15762), .ZN(n11939) );
  NAND2_X1 U14633 ( .A1(n15763), .A2(n13858), .ZN(n11938) );
  OAI211_X1 U14634 ( .C1(n15830), .C2(n14461), .A(n11939), .B(n11938), .ZN(
        n11940) );
  AOI21_X1 U14635 ( .B1(n15836), .B2(n15771), .A(n11940), .ZN(n11941) );
  OAI21_X1 U14636 ( .B1(n15832), .B2(n15783), .A(n11941), .ZN(P2_U3258) );
  AND2_X1 U14637 ( .A1(n12936), .A2(n12937), .ZN(n12935) );
  XNOR2_X1 U14638 ( .A(n11942), .B(n12935), .ZN(n11947) );
  XNOR2_X1 U14639 ( .A(n11943), .B(n12935), .ZN(n11987) );
  OAI22_X1 U14640 ( .A1(n15861), .A2(n11944), .B1(n12207), .B2(n15859), .ZN(
        n11945) );
  AOI21_X1 U14641 ( .B1(n11987), .B2(n12150), .A(n11945), .ZN(n11946) );
  OAI21_X1 U14642 ( .B1(n11947), .B2(n13401), .A(n11946), .ZN(n11986) );
  INV_X1 U14643 ( .A(n11986), .ZN(n11954) );
  NOR2_X1 U14644 ( .A1(n15870), .A2(n11948), .ZN(n11952) );
  OAI22_X1 U14645 ( .A1(n13266), .A2(n11950), .B1(n11949), .B2(n15855), .ZN(
        n11951) );
  AOI211_X1 U14646 ( .C1(n11987), .C2(n13212), .A(n11952), .B(n11951), .ZN(
        n11953) );
  OAI21_X1 U14647 ( .B1(n11954), .B2(n15873), .A(n11953), .ZN(P3_U3224) );
  MUX2_X1 U14648 ( .A(n13037), .B(n11956), .S(n11955), .Z(n11957) );
  XOR2_X1 U14649 ( .A(n11958), .B(n11957), .Z(n11964) );
  AOI21_X1 U14650 ( .B1(n12834), .B2(n13035), .A(n11959), .ZN(n11960) );
  OAI21_X1 U14651 ( .B1(n6954), .B2(n12836), .A(n11960), .ZN(n11962) );
  NOR2_X1 U14652 ( .A1(n12536), .A2(n12096), .ZN(n11961) );
  AOI211_X1 U14653 ( .C1(n12803), .C2(n13498), .A(n11962), .B(n11961), .ZN(
        n11963) );
  OAI21_X1 U14654 ( .B1(n11964), .B2(n12815), .A(n11963), .ZN(P3_U3161) );
  NAND3_X1 U14655 ( .A1(n11966), .A2(n10587), .A3(n11965), .ZN(n11967) );
  NAND2_X1 U14656 ( .A1(n11968), .A2(n11967), .ZN(n11969) );
  NAND2_X1 U14657 ( .A1(n11969), .A2(n15759), .ZN(n11971) );
  AOI22_X1 U14658 ( .A1(n14104), .A2(n14451), .B1(n14449), .B2(n14101), .ZN(
        n11970) );
  NAND2_X1 U14659 ( .A1(n11971), .A2(n11970), .ZN(n15801) );
  INV_X1 U14660 ( .A(n15801), .ZN(n11985) );
  NAND2_X1 U14661 ( .A1(n14036), .A2(n11972), .ZN(n11974) );
  OAI21_X1 U14662 ( .B1(n11975), .B2(n11974), .A(n11973), .ZN(n15803) );
  INV_X1 U14663 ( .A(n11976), .ZN(n11979) );
  INV_X1 U14664 ( .A(n11977), .ZN(n11978) );
  OAI211_X1 U14665 ( .C1(n15800), .C2(n11979), .A(n11978), .B(n11714), .ZN(
        n15799) );
  OAI22_X1 U14666 ( .A1(n15781), .A2(n11980), .B1(n7274), .B2(n15776), .ZN(
        n11981) );
  AOI21_X1 U14667 ( .B1(n15763), .B2(n13813), .A(n11981), .ZN(n11982) );
  OAI21_X1 U14668 ( .B1(n14461), .B2(n15799), .A(n11982), .ZN(n11983) );
  AOI21_X1 U14669 ( .B1(n15771), .B2(n15803), .A(n11983), .ZN(n11984) );
  OAI21_X1 U14670 ( .B1(n15783), .B2(n11985), .A(n11984), .ZN(P2_U3263) );
  INV_X1 U14671 ( .A(n15886), .ZN(n15879) );
  AOI21_X1 U14672 ( .B1(n15879), .B2(n11987), .A(n11986), .ZN(n11991) );
  AOI22_X1 U14673 ( .A1(n10701), .A2(n11989), .B1(P3_REG0_REG_9__SCAN_IN), 
        .B2(n15906), .ZN(n11988) );
  OAI21_X1 U14674 ( .B1(n11991), .B2(n15906), .A(n11988), .ZN(P3_U3417) );
  AOI22_X1 U14675 ( .A1(n13488), .A2(n11989), .B1(P3_REG1_REG_9__SCAN_IN), 
        .B2(n10706), .ZN(n11990) );
  OAI21_X1 U14676 ( .B1(n11991), .B2(n10706), .A(n11990), .ZN(P3_U3468) );
  OAI211_X1 U14677 ( .C1(n11993), .C2(n12001), .A(n11992), .B(n15545), .ZN(
        n11995) );
  AOI22_X1 U14678 ( .A1(n15256), .A2(n15258), .B1(n14846), .B2(n15257), .ZN(
        n11994) );
  NAND2_X1 U14679 ( .A1(n11996), .A2(n15384), .ZN(n11997) );
  AND2_X1 U14680 ( .A1(n6702), .A2(n11997), .ZN(n15385) );
  INV_X1 U14681 ( .A(n12168), .ZN(n11998) );
  AOI22_X1 U14682 ( .A1(n15262), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n11998), 
        .B2(n15513), .ZN(n11999) );
  OAI21_X1 U14683 ( .B1(n7846), .B2(n15517), .A(n11999), .ZN(n12003) );
  XNOR2_X1 U14684 ( .A(n12000), .B(n12001), .ZN(n15388) );
  NOR2_X1 U14685 ( .A1(n15388), .A2(n15267), .ZN(n12002) );
  AOI211_X1 U14686 ( .C1(n15385), .C2(n15520), .A(n12003), .B(n12002), .ZN(
        n12004) );
  OAI21_X1 U14687 ( .B1(n15262), .B2(n15387), .A(n12004), .ZN(P1_U3282) );
  INV_X1 U14688 ( .A(n12036), .ZN(n12007) );
  AOI21_X1 U14689 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n15424), .A(n12005), 
        .ZN(n12006) );
  OAI21_X1 U14690 ( .B1(n12007), .B2(n15438), .A(n12006), .ZN(P1_U3332) );
  AND2_X1 U14691 ( .A1(n15781), .A2(n15780), .ZN(n12056) );
  OR2_X1 U14692 ( .A1(n12009), .A2(n12008), .ZN(n12010) );
  AND2_X1 U14693 ( .A1(n12011), .A2(n12010), .ZN(n12021) );
  INV_X1 U14694 ( .A(n12021), .ZN(n15809) );
  OAI211_X1 U14695 ( .C1(n10198), .C2(n15806), .A(n15767), .B(n12013), .ZN(
        n15805) );
  AOI22_X1 U14696 ( .A1(n15763), .A2(n13843), .B1(n12014), .B2(n15762), .ZN(
        n12015) );
  OAI21_X1 U14697 ( .B1(n14461), .B2(n15805), .A(n12015), .ZN(n12023) );
  OAI21_X1 U14698 ( .B1(n12017), .B2(n14038), .A(n12016), .ZN(n12018) );
  NAND2_X1 U14699 ( .A1(n12018), .A2(n15759), .ZN(n12020) );
  AOI22_X1 U14700 ( .A1(n14449), .A2(n14099), .B1(n14451), .B2(n14101), .ZN(
        n12019) );
  OAI211_X1 U14701 ( .C1(n12021), .C2(n14479), .A(n12020), .B(n12019), .ZN(
        n15807) );
  MUX2_X1 U14702 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n15807), .S(n15781), .Z(
        n12022) );
  AOI211_X1 U14703 ( .C1(n12056), .C2(n15809), .A(n12023), .B(n12022), .ZN(
        n12024) );
  INV_X1 U14704 ( .A(n12024), .ZN(P2_U3261) );
  INV_X1 U14705 ( .A(n14479), .ZN(n14446) );
  NAND2_X1 U14706 ( .A1(n12025), .A2(n12026), .ZN(n12027) );
  XNOR2_X1 U14707 ( .A(n14047), .B(n12027), .ZN(n14603) );
  XNOR2_X1 U14708 ( .A(n14047), .B(n12028), .ZN(n12030) );
  AOI22_X1 U14709 ( .A1(n8009), .A2(n14451), .B1(n14450), .B2(n14449), .ZN(
        n12029) );
  OAI21_X1 U14710 ( .B1(n12030), .B2(n14425), .A(n12029), .ZN(n12031) );
  AOI21_X1 U14711 ( .B1(n14446), .B2(n14603), .A(n12031), .ZN(n14607) );
  AOI211_X1 U14712 ( .C1(n14605), .C2(n12083), .A(n14481), .B(n14480), .ZN(
        n14604) );
  NAND2_X1 U14713 ( .A1(n14604), .A2(n15770), .ZN(n12033) );
  AOI22_X1 U14714 ( .A1(n15783), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n12230), 
        .B2(n15762), .ZN(n12032) );
  OAI211_X1 U14715 ( .C1(n7655), .C2(n14436), .A(n12033), .B(n12032), .ZN(
        n12034) );
  AOI21_X1 U14716 ( .B1(n14603), .B2(n12056), .A(n12034), .ZN(n12035) );
  OAI21_X1 U14717 ( .B1(n14607), .B2(n15783), .A(n12035), .ZN(P2_U3255) );
  NAND2_X1 U14718 ( .A1(n12036), .A2(n14664), .ZN(n12038) );
  OR2_X1 U14719 ( .A1(n12037), .A2(n6510), .ZN(n14073) );
  OAI211_X1 U14720 ( .C1(n12039), .C2(n14671), .A(n12038), .B(n14073), .ZN(
        P2_U3304) );
  INV_X1 U14721 ( .A(n12040), .ZN(n12046) );
  AOI22_X1 U14722 ( .A1(n15763), .A2(n10379), .B1(n15762), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n12041) );
  OAI21_X1 U14723 ( .B1(n14461), .B2(n12042), .A(n12041), .ZN(n12045) );
  MUX2_X1 U14724 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n12043), .S(n15781), .Z(
        n12044) );
  AOI211_X1 U14725 ( .C1(n12056), .C2(n12046), .A(n12045), .B(n12044), .ZN(
        n12047) );
  INV_X1 U14726 ( .A(n12047), .ZN(P2_U3264) );
  XOR2_X1 U14727 ( .A(n12048), .B(n14044), .Z(n12052) );
  OAI22_X1 U14728 ( .A1(n13859), .A2(n14472), .B1(n13868), .B2(n14474), .ZN(
        n12051) );
  XNOR2_X1 U14729 ( .A(n12049), .B(n14044), .ZN(n14612) );
  NOR2_X1 U14730 ( .A1(n14612), .A2(n14479), .ZN(n12050) );
  AOI211_X1 U14731 ( .C1(n12052), .C2(n15759), .A(n12051), .B(n12050), .ZN(
        n14611) );
  INV_X1 U14732 ( .A(n12081), .ZN(n12053) );
  AOI211_X1 U14733 ( .C1(n7205), .C2(n12054), .A(n14481), .B(n12053), .ZN(
        n14609) );
  AOI22_X1 U14734 ( .A1(n15783), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n8087), .B2(
        n15762), .ZN(n12055) );
  OAI21_X1 U14735 ( .B1(n10221), .B2(n14436), .A(n12055), .ZN(n12058) );
  NOR2_X1 U14736 ( .A1(n14612), .A2(n14489), .ZN(n12057) );
  AOI211_X1 U14737 ( .C1(n14609), .C2(n15770), .A(n12058), .B(n12057), .ZN(
        n12059) );
  OAI21_X1 U14738 ( .B1(n14611), .B2(n15783), .A(n12059), .ZN(P2_U3257) );
  XNOR2_X1 U14739 ( .A(n12174), .B(n12060), .ZN(n12177) );
  XNOR2_X1 U14740 ( .A(n12177), .B(n12061), .ZN(n12068) );
  NAND2_X1 U14741 ( .A1(n15500), .A2(n12062), .ZN(n12064) );
  OAI211_X1 U14742 ( .C1(n15508), .C2(n12065), .A(n12064), .B(n12063), .ZN(
        n12066) );
  AOI21_X1 U14743 ( .B1(n15396), .B2(n14830), .A(n12066), .ZN(n12067) );
  OAI21_X1 U14744 ( .B1(n12068), .B2(n15496), .A(n12067), .ZN(P1_U3231) );
  AND2_X1 U14745 ( .A1(n12025), .A2(n12069), .ZN(n12074) );
  OR2_X1 U14746 ( .A1(n12049), .A2(n14044), .ZN(n12071) );
  NAND2_X1 U14747 ( .A1(n12071), .A2(n12070), .ZN(n12072) );
  OR2_X1 U14748 ( .A1(n12072), .A2(n14046), .ZN(n12073) );
  NAND2_X1 U14749 ( .A1(n12074), .A2(n12073), .ZN(n12113) );
  XNOR2_X1 U14750 ( .A(n12075), .B(n14046), .ZN(n12076) );
  NAND2_X1 U14751 ( .A1(n12076), .A2(n15759), .ZN(n12078) );
  AOI22_X1 U14752 ( .A1(n14451), .A2(n14096), .B1(n14449), .B2(n14095), .ZN(
        n12077) );
  OAI211_X1 U14753 ( .C1(n14479), .C2(n12113), .A(n12078), .B(n12077), .ZN(
        n12114) );
  INV_X1 U14754 ( .A(n12114), .ZN(n12079) );
  MUX2_X1 U14755 ( .A(n12080), .B(n12079), .S(n15781), .Z(n12087) );
  AOI21_X1 U14756 ( .B1(n12081), .B2(n13870), .A(n14481), .ZN(n12082) );
  AND2_X1 U14757 ( .A1(n12083), .A2(n12082), .ZN(n12115) );
  INV_X1 U14758 ( .A(n13870), .ZN(n13869) );
  INV_X1 U14759 ( .A(n12591), .ZN(n12084) );
  OAI22_X1 U14760 ( .A1(n13869), .A2(n14436), .B1(n12084), .B2(n15776), .ZN(
        n12085) );
  AOI21_X1 U14761 ( .B1(n12115), .B2(n15770), .A(n12085), .ZN(n12086) );
  OAI211_X1 U14762 ( .C1(n12113), .C2(n14489), .A(n12087), .B(n12086), .ZN(
        P2_U3256) );
  NOR2_X1 U14763 ( .A1(n15873), .A2(n15866), .ZN(n12088) );
  OR2_X1 U14764 ( .A1(n13212), .A2(n12088), .ZN(n13268) );
  INV_X1 U14765 ( .A(n13268), .ZN(n13243) );
  XOR2_X1 U14766 ( .A(n12089), .B(n12930), .Z(n13501) );
  INV_X1 U14767 ( .A(n12090), .ZN(n12091) );
  AOI21_X1 U14768 ( .B1(n12930), .B2(n12092), .A(n12091), .ZN(n12093) );
  OAI222_X1 U14769 ( .A1(n15859), .A2(n12148), .B1(n15861), .B2(n6954), .C1(
        n13401), .C2(n12093), .ZN(n13497) );
  INV_X1 U14770 ( .A(n13497), .ZN(n12094) );
  MUX2_X1 U14771 ( .A(n12095), .B(n12094), .S(n15870), .Z(n12099) );
  INV_X1 U14772 ( .A(n12096), .ZN(n12097) );
  AOI22_X1 U14773 ( .A1(n13428), .A2(n13498), .B1(n13427), .B2(n12097), .ZN(
        n12098) );
  OAI211_X1 U14774 ( .C1(n13243), .C2(n13501), .A(n12099), .B(n12098), .ZN(
        P3_U3225) );
  AOI21_X1 U14775 ( .B1(n13424), .B2(n12100), .A(n13046), .ZN(n12112) );
  NAND2_X1 U14776 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n12206)
         );
  OAI21_X1 U14777 ( .B1(n13144), .B2(n12101), .A(n12206), .ZN(n12105) );
  AOI21_X1 U14778 ( .B1(n6703), .B2(n12102), .A(n13059), .ZN(n12103) );
  NOR2_X1 U14779 ( .A1(n12103), .A2(n13146), .ZN(n12104) );
  AOI211_X1 U14780 ( .C1(n13152), .C2(n12106), .A(n12105), .B(n12104), .ZN(
        n12111) );
  OAI21_X1 U14781 ( .B1(n12108), .B2(P3_REG1_REG_11__SCAN_IN), .A(n12107), 
        .ZN(n12109) );
  NAND2_X1 U14782 ( .A1(n12109), .A2(n13180), .ZN(n12110) );
  OAI211_X1 U14783 ( .C1(n12112), .C2(n13182), .A(n12111), .B(n12110), .ZN(
        P3_U3193) );
  INV_X1 U14784 ( .A(n12113), .ZN(n12116) );
  INV_X1 U14785 ( .A(n13811), .ZN(n15810) );
  AOI211_X1 U14786 ( .C1(n12116), .C2(n15810), .A(n12115), .B(n12114), .ZN(
        n12145) );
  AOI22_X1 U14787 ( .A1(n7368), .A2(n13870), .B1(P2_REG0_REG_9__SCAN_IN), .B2(
        n7304), .ZN(n12117) );
  OAI21_X1 U14788 ( .B1(n12145), .B2(n7304), .A(n12117), .ZN(P2_U3457) );
  NAND2_X1 U14789 ( .A1(n14311), .A2(n14096), .ZN(n12120) );
  XNOR2_X1 U14790 ( .A(n12586), .B(n12120), .ZN(n12716) );
  INV_X1 U14791 ( .A(n12586), .ZN(n12121) );
  XNOR2_X1 U14792 ( .A(n13870), .B(n11713), .ZN(n12124) );
  NOR2_X1 U14793 ( .A1(n13868), .A2(n15767), .ZN(n12122) );
  XNOR2_X1 U14794 ( .A(n12124), .B(n12122), .ZN(n12585) );
  INV_X1 U14795 ( .A(n12122), .ZN(n12123) );
  XNOR2_X1 U14796 ( .A(n14605), .B(n11713), .ZN(n12127) );
  NAND2_X1 U14797 ( .A1(n14481), .A2(n14095), .ZN(n12128) );
  XNOR2_X1 U14798 ( .A(n12127), .B(n12128), .ZN(n12235) );
  INV_X1 U14799 ( .A(n12127), .ZN(n12130) );
  INV_X1 U14800 ( .A(n12128), .ZN(n12129) );
  NAND2_X1 U14801 ( .A1(n12130), .A2(n12129), .ZN(n12131) );
  XNOR2_X1 U14802 ( .A(n14483), .B(n12669), .ZN(n12135) );
  INV_X1 U14803 ( .A(n12135), .ZN(n12133) );
  AND2_X1 U14804 ( .A1(n14481), .A2(n14450), .ZN(n12134) );
  INV_X1 U14805 ( .A(n12134), .ZN(n12132) );
  NAND2_X1 U14806 ( .A1(n12133), .A2(n12132), .ZN(n12600) );
  NAND2_X1 U14807 ( .A1(n12135), .A2(n12134), .ZN(n12598) );
  NAND2_X1 U14808 ( .A1(n12600), .A2(n12598), .ZN(n12136) );
  XNOR2_X1 U14809 ( .A(n12599), .B(n12136), .ZN(n12141) );
  AOI22_X1 U14810 ( .A1(n13770), .A2(n14095), .B1(n13750), .B2(n14484), .ZN(
        n12138) );
  OAI211_X1 U14811 ( .C1(n14475), .C2(n13803), .A(n12138), .B(n12137), .ZN(
        n12139) );
  AOI21_X1 U14812 ( .B1(n14483), .B2(n13808), .A(n12139), .ZN(n12140) );
  OAI21_X1 U14813 ( .B1(n12141), .B2(n13796), .A(n12140), .ZN(P2_U3208) );
  NAND2_X1 U14814 ( .A1(n7285), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n12144) );
  NAND2_X1 U14815 ( .A1(n12142), .A2(n13870), .ZN(n12143) );
  OAI211_X1 U14816 ( .C1(n12145), .C2(n7285), .A(n12144), .B(n12143), .ZN(
        P2_U3508) );
  XNOR2_X1 U14817 ( .A(n12146), .B(n12941), .ZN(n12152) );
  XOR2_X1 U14818 ( .A(n12147), .B(n12941), .Z(n13493) );
  OAI22_X1 U14819 ( .A1(n15861), .A2(n12148), .B1(n13402), .B2(n15859), .ZN(
        n12149) );
  AOI21_X1 U14820 ( .B1(n13493), .B2(n12150), .A(n12149), .ZN(n12151) );
  OAI21_X1 U14821 ( .B1(n13401), .B2(n12152), .A(n12151), .ZN(n13492) );
  INV_X1 U14822 ( .A(n13492), .ZN(n12158) );
  NOR2_X1 U14823 ( .A1(n13266), .A2(n13598), .ZN(n12156) );
  OAI22_X1 U14824 ( .A1(n15870), .A2(n12154), .B1(n12153), .B2(n15855), .ZN(
        n12155) );
  AOI211_X1 U14825 ( .C1(n13493), .C2(n13212), .A(n12156), .B(n12155), .ZN(
        n12157) );
  OAI21_X1 U14826 ( .B1(n12158), .B2(n15873), .A(n12157), .ZN(P3_U3223) );
  OAI222_X1 U14827 ( .A1(P2_U3088), .A2(n12160), .B1(n14673), .B2(n12162), 
        .C1(n12159), .C2(n14671), .ZN(P2_U3303) );
  OAI222_X1 U14828 ( .A1(n8980), .A2(P1_U3086), .B1(n15438), .B2(n12162), .C1(
        n12161), .C2(n15435), .ZN(P1_U3331) );
  INV_X1 U14829 ( .A(n12163), .ZN(n12164) );
  AOI21_X1 U14830 ( .B1(n12166), .B2(n12165), .A(n12164), .ZN(n12173) );
  OAI21_X1 U14831 ( .B1(n15508), .B2(n12168), .A(n12167), .ZN(n12171) );
  OAI22_X1 U14832 ( .A1(n14826), .A2(n14785), .B1(n12169), .B2(n14825), .ZN(
        n12170) );
  AOI211_X1 U14833 ( .C1(n15384), .C2(n14830), .A(n12171), .B(n12170), .ZN(
        n12172) );
  OAI21_X1 U14834 ( .B1(n12173), .B2(n15496), .A(n12172), .ZN(P1_U3236) );
  AOI22_X1 U14835 ( .A1(n12177), .A2(n12176), .B1(n12175), .B2(n12174), .ZN(
        n12181) );
  XNOR2_X1 U14836 ( .A(n12179), .B(n12178), .ZN(n12180) );
  XNOR2_X1 U14837 ( .A(n12181), .B(n12180), .ZN(n12187) );
  NAND2_X1 U14838 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n14931)
         );
  OAI21_X1 U14839 ( .B1(n15508), .B2(n12182), .A(n14931), .ZN(n12185) );
  OAI22_X1 U14840 ( .A1(n14826), .A2(n14729), .B1(n12183), .B2(n14825), .ZN(
        n12184) );
  AOI211_X1 U14841 ( .C1(n15391), .C2(n14830), .A(n12185), .B(n12184), .ZN(
        n12186) );
  OAI21_X1 U14842 ( .B1(n12187), .B2(n15496), .A(n12186), .ZN(P1_U3217) );
  XNOR2_X1 U14843 ( .A(n12188), .B(n12189), .ZN(n12194) );
  INV_X1 U14844 ( .A(n12194), .ZN(n15381) );
  OAI211_X1 U14845 ( .C1(n12192), .C2(n12191), .A(n12190), .B(n15545), .ZN(
        n12197) );
  OAI22_X1 U14846 ( .A1(n15226), .A2(n15227), .B1(n14729), .B2(n15225), .ZN(
        n12193) );
  INV_X1 U14847 ( .A(n12193), .ZN(n12196) );
  NAND2_X1 U14848 ( .A1(n12194), .A2(n15552), .ZN(n12195) );
  NAND3_X1 U14849 ( .A1(n12197), .A2(n12196), .A3(n12195), .ZN(n15383) );
  NAND2_X1 U14850 ( .A1(n15383), .A2(n15232), .ZN(n12203) );
  OAI22_X1 U14851 ( .A1(n15232), .A2(n12198), .B1(n14728), .B2(n15259), .ZN(
        n12201) );
  AND2_X1 U14852 ( .A1(n6702), .A2(n14724), .ZN(n12199) );
  OR2_X1 U14853 ( .A1(n12199), .A2(n15251), .ZN(n15378) );
  NOR2_X1 U14854 ( .A1(n15378), .A2(n15236), .ZN(n12200) );
  AOI211_X1 U14855 ( .C1(n15239), .C2(n14724), .A(n12201), .B(n12200), .ZN(
        n12202) );
  OAI211_X1 U14856 ( .C1(n15381), .C2(n12204), .A(n12203), .B(n12202), .ZN(
        P1_U3281) );
  XOR2_X1 U14857 ( .A(n12527), .B(n12526), .Z(n12528) );
  XNOR2_X1 U14858 ( .A(n12528), .B(n13034), .ZN(n12212) );
  INV_X1 U14859 ( .A(n12205), .ZN(n13590) );
  OAI21_X1 U14860 ( .B1(n12836), .B2(n12207), .A(n12206), .ZN(n12208) );
  AOI21_X1 U14861 ( .B1(n12834), .B2(n13421), .A(n12208), .ZN(n12209) );
  OAI21_X1 U14862 ( .B1(n12536), .B2(n13425), .A(n12209), .ZN(n12210) );
  AOI21_X1 U14863 ( .B1(n13590), .B2(n12803), .A(n12210), .ZN(n12211) );
  OAI21_X1 U14864 ( .B1(n12212), .B2(n12815), .A(n12211), .ZN(P3_U3176) );
  INV_X1 U14865 ( .A(n12213), .ZN(n12214) );
  AOI211_X1 U14866 ( .C1(n12217), .C2(n12216), .A(n12215), .B(n12214), .ZN(
        n12229) );
  INV_X1 U14867 ( .A(n12218), .ZN(n12219) );
  AOI211_X1 U14868 ( .C1(n12222), .C2(n12221), .A(n12220), .B(n12219), .ZN(
        n12228) );
  AND2_X1 U14869 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14751) );
  AOI21_X1 U14870 ( .B1(n12223), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n14751), 
        .ZN(n12224) );
  OAI21_X1 U14871 ( .B1(n12226), .B2(n12225), .A(n12224), .ZN(n12227) );
  OR3_X1 U14872 ( .A1(n12229), .A2(n12228), .A3(n12227), .ZN(P1_U3259) );
  AOI22_X1 U14873 ( .A1(n13769), .A2(n14450), .B1(n13750), .B2(n12230), .ZN(
        n12231) );
  NAND2_X1 U14874 ( .A1(n6510), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n15691) );
  OAI211_X1 U14875 ( .C1(n13868), .C2(n13805), .A(n12231), .B(n15691), .ZN(
        n12237) );
  INV_X1 U14876 ( .A(n12232), .ZN(n12233) );
  AOI211_X1 U14877 ( .C1(n12235), .C2(n12234), .A(n13796), .B(n12233), .ZN(
        n12236) );
  AOI211_X1 U14878 ( .C1(n14605), .C2(n13808), .A(n12237), .B(n12236), .ZN(
        n12238) );
  INV_X1 U14879 ( .A(n12238), .ZN(P2_U3189) );
  XNOR2_X1 U14880 ( .A(n12239), .B(n13381), .ZN(n12240) );
  XNOR2_X1 U14881 ( .A(n12241), .B(n12240), .ZN(n12247) );
  INV_X1 U14882 ( .A(n12242), .ZN(n13395) );
  NAND2_X1 U14883 ( .A1(n12834), .A2(n13392), .ZN(n12243) );
  NAND2_X1 U14884 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n13067)
         );
  OAI211_X1 U14885 ( .C1(n12531), .C2(n12836), .A(n12243), .B(n13067), .ZN(
        n12244) );
  AOI21_X1 U14886 ( .B1(n13395), .B2(n12839), .A(n12244), .ZN(n12245) );
  OAI21_X1 U14887 ( .B1(n12896), .B2(n12842), .A(n12245), .ZN(n12246) );
  AOI21_X1 U14888 ( .B1(n12247), .B2(n12832), .A(n12246), .ZN(n12525) );
  AOI22_X1 U14889 ( .A1(n12249), .A2(keyinput30), .B1(n12451), .B2(keyinput43), 
        .ZN(n12248) );
  OAI221_X1 U14890 ( .B1(n12249), .B2(keyinput30), .C1(n12451), .C2(keyinput43), .A(n12248), .ZN(n12254) );
  AOI22_X1 U14891 ( .A1(n15591), .A2(keyinput113), .B1(n12251), .B2(
        keyinput101), .ZN(n12250) );
  OAI221_X1 U14892 ( .B1(n15591), .B2(keyinput113), .C1(n12251), .C2(
        keyinput101), .A(n12250), .ZN(n12253) );
  INV_X1 U14893 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n15785) );
  XNOR2_X1 U14894 ( .A(n15785), .B(keyinput69), .ZN(n12252) );
  OR3_X1 U14895 ( .A1(n12254), .A2(n12253), .A3(n12252), .ZN(n12263) );
  AOI22_X1 U14896 ( .A1(n12257), .A2(keyinput125), .B1(n12256), .B2(
        keyinput115), .ZN(n12255) );
  OAI221_X1 U14897 ( .B1(n12257), .B2(keyinput125), .C1(n12256), .C2(
        keyinput115), .A(n12255), .ZN(n12262) );
  AOI22_X1 U14898 ( .A1(n12259), .A2(keyinput32), .B1(n9451), .B2(keyinput93), 
        .ZN(n12258) );
  OAI221_X1 U14899 ( .B1(n12259), .B2(keyinput32), .C1(n9451), .C2(keyinput93), 
        .A(n12258), .ZN(n12261) );
  INV_X1 U14900 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n15529) );
  XNOR2_X1 U14901 ( .A(n15529), .B(keyinput21), .ZN(n12260) );
  OR4_X1 U14902 ( .A1(n12263), .A2(n12262), .A3(n12261), .A4(n12260), .ZN(
        n12412) );
  INV_X1 U14903 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U14904 ( .A1(n9418), .A2(keyinput67), .B1(keyinput40), .B2(n12265), 
        .ZN(n12264) );
  OAI221_X1 U14905 ( .B1(n9418), .B2(keyinput67), .C1(n12265), .C2(keyinput40), 
        .A(n12264), .ZN(n12270) );
  INV_X1 U14906 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n12821) );
  AOI22_X1 U14907 ( .A1(n12462), .A2(keyinput28), .B1(n12821), .B2(keyinput59), 
        .ZN(n12266) );
  OAI221_X1 U14908 ( .B1(n12462), .B2(keyinput28), .C1(n12821), .C2(keyinput59), .A(n12266), .ZN(n12269) );
  INV_X1 U14909 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n15429) );
  AOI22_X1 U14910 ( .A1(n15429), .A2(keyinput76), .B1(n12504), .B2(keyinput54), 
        .ZN(n12267) );
  OAI221_X1 U14911 ( .B1(n15429), .B2(keyinput76), .C1(n12504), .C2(keyinput54), .A(n12267), .ZN(n12268) );
  NOR3_X1 U14912 ( .A1(n12270), .A2(n12269), .A3(n12268), .ZN(n12294) );
  AOI22_X1 U14913 ( .A1(n10731), .A2(keyinput122), .B1(keyinput123), .B2(
        n12272), .ZN(n12271) );
  OAI221_X1 U14914 ( .B1(n10731), .B2(keyinput122), .C1(n12272), .C2(
        keyinput123), .A(n12271), .ZN(n12278) );
  AOI22_X1 U14915 ( .A1(n6971), .A2(keyinput37), .B1(n12274), .B2(keyinput78), 
        .ZN(n12273) );
  OAI221_X1 U14916 ( .B1(n6971), .B2(keyinput37), .C1(n12274), .C2(keyinput78), 
        .A(n12273), .ZN(n12277) );
  AOI22_X1 U14917 ( .A1(n12511), .A2(keyinput41), .B1(n12512), .B2(keyinput110), .ZN(n12275) );
  OAI221_X1 U14918 ( .B1(n12511), .B2(keyinput41), .C1(n12512), .C2(
        keyinput110), .A(n12275), .ZN(n12276) );
  NOR3_X1 U14919 ( .A1(n12278), .A2(n12277), .A3(n12276), .ZN(n12293) );
  AOI22_X1 U14920 ( .A1(n12280), .A2(keyinput116), .B1(n12452), .B2(keyinput23), .ZN(n12279) );
  OAI221_X1 U14921 ( .B1(n12280), .B2(keyinput116), .C1(n12452), .C2(
        keyinput23), .A(n12279), .ZN(n12284) );
  INV_X1 U14922 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U14923 ( .A1(n12455), .A2(keyinput48), .B1(n12282), .B2(keyinput4), 
        .ZN(n12281) );
  OAI221_X1 U14924 ( .B1(n12455), .B2(keyinput48), .C1(n12282), .C2(keyinput4), 
        .A(n12281), .ZN(n12283) );
  NOR2_X1 U14925 ( .A1(n12284), .A2(n12283), .ZN(n12292) );
  INV_X1 U14926 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15811) );
  INV_X1 U14927 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n12286) );
  AOI22_X1 U14928 ( .A1(n15811), .A2(keyinput35), .B1(keyinput8), .B2(n12286), 
        .ZN(n12285) );
  OAI221_X1 U14929 ( .B1(n15811), .B2(keyinput35), .C1(n12286), .C2(keyinput8), 
        .A(n12285), .ZN(n12290) );
  INV_X1 U14930 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n12510) );
  AOI22_X1 U14931 ( .A1(n12510), .A2(keyinput126), .B1(n12288), .B2(keyinput94), .ZN(n12287) );
  OAI221_X1 U14932 ( .B1(n12510), .B2(keyinput126), .C1(n12288), .C2(
        keyinput94), .A(n12287), .ZN(n12289) );
  NOR2_X1 U14933 ( .A1(n12290), .A2(n12289), .ZN(n12291) );
  NAND4_X1 U14934 ( .A1(n12294), .A2(n12293), .A3(n12292), .A4(n12291), .ZN(
        n12411) );
  XOR2_X1 U14935 ( .A(P2_IR_REG_5__SCAN_IN), .B(keyinput102), .Z(n12300) );
  XNOR2_X1 U14936 ( .A(n12483), .B(keyinput75), .ZN(n12299) );
  XNOR2_X1 U14937 ( .A(n12295), .B(keyinput86), .ZN(n12298) );
  XNOR2_X1 U14938 ( .A(n12296), .B(keyinput66), .ZN(n12297) );
  NOR4_X1 U14939 ( .A1(n12300), .A2(n12299), .A3(n12298), .A4(n12297), .ZN(
        n12323) );
  XOR2_X1 U14940 ( .A(P3_IR_REG_1__SCAN_IN), .B(keyinput65), .Z(n12307) );
  XNOR2_X1 U14941 ( .A(n12301), .B(keyinput53), .ZN(n12306) );
  XNOR2_X1 U14942 ( .A(n12302), .B(keyinput62), .ZN(n12305) );
  XNOR2_X1 U14943 ( .A(n12303), .B(keyinput73), .ZN(n12304) );
  NOR4_X1 U14944 ( .A1(n12307), .A2(n12306), .A3(n12305), .A4(n12304), .ZN(
        n12322) );
  XNOR2_X1 U14945 ( .A(n12489), .B(keyinput20), .ZN(n12313) );
  XNOR2_X1 U14946 ( .A(n12308), .B(keyinput44), .ZN(n12312) );
  XNOR2_X1 U14947 ( .A(n12309), .B(keyinput14), .ZN(n12311) );
  XNOR2_X1 U14948 ( .A(keyinput107), .B(n8353), .ZN(n12310) );
  NOR4_X1 U14949 ( .A1(n12313), .A2(n12312), .A3(n12311), .A4(n12310), .ZN(
        n12321) );
  INV_X1 U14950 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n12314) );
  XNOR2_X1 U14951 ( .A(keyinput108), .B(n12314), .ZN(n12319) );
  XNOR2_X1 U14952 ( .A(keyinput91), .B(n12315), .ZN(n12318) );
  XNOR2_X1 U14953 ( .A(keyinput71), .B(n10380), .ZN(n12317) );
  XNOR2_X1 U14954 ( .A(keyinput82), .B(n15840), .ZN(n12316) );
  NOR4_X1 U14955 ( .A1(n12319), .A2(n12318), .A3(n12317), .A4(n12316), .ZN(
        n12320) );
  NAND4_X1 U14956 ( .A1(n12323), .A2(n12322), .A3(n12321), .A4(n12320), .ZN(
        n12333) );
  AOI22_X1 U14957 ( .A1(n9723), .A2(keyinput112), .B1(n12570), .B2(keyinput80), 
        .ZN(n12324) );
  OAI221_X1 U14958 ( .B1(n9723), .B2(keyinput112), .C1(n12570), .C2(keyinput80), .A(n12324), .ZN(n12332) );
  INV_X1 U14959 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15705) );
  XNOR2_X1 U14960 ( .A(n15705), .B(keyinput57), .ZN(n12331) );
  INV_X1 U14961 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n15786) );
  XOR2_X1 U14962 ( .A(n15786), .B(keyinput55), .Z(n12329) );
  XOR2_X1 U14963 ( .A(n12325), .B(keyinput33), .Z(n12328) );
  XOR2_X1 U14964 ( .A(n12475), .B(keyinput1), .Z(n12327) );
  XOR2_X1 U14965 ( .A(n10391), .B(keyinput15), .Z(n12326) );
  NAND4_X1 U14966 ( .A1(n12329), .A2(n12328), .A3(n12327), .A4(n12326), .ZN(
        n12330) );
  NOR4_X1 U14967 ( .A1(n12333), .A2(n12332), .A3(n12331), .A4(n12330), .ZN(
        n12409) );
  INV_X1 U14968 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n15788) );
  AOI22_X1 U14969 ( .A1(n15788), .A2(keyinput109), .B1(keyinput120), .B2(
        n12335), .ZN(n12334) );
  OAI221_X1 U14970 ( .B1(n15788), .B2(keyinput109), .C1(n12335), .C2(
        keyinput120), .A(n12334), .ZN(n12338) );
  XNOR2_X1 U14971 ( .A(n12336), .B(keyinput27), .ZN(n12337) );
  NOR2_X1 U14972 ( .A1(n12338), .A2(n12337), .ZN(n12352) );
  INV_X1 U14973 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n15528) );
  AOI22_X1 U14974 ( .A1(n15528), .A2(keyinput92), .B1(n12484), .B2(keyinput121), .ZN(n12339) );
  OAI221_X1 U14975 ( .B1(n15528), .B2(keyinput92), .C1(n12484), .C2(
        keyinput121), .A(n12339), .ZN(n12342) );
  AOI22_X1 U14976 ( .A1(n13521), .A2(keyinput95), .B1(keyinput99), .B2(n7506), 
        .ZN(n12340) );
  OAI221_X1 U14977 ( .B1(n13521), .B2(keyinput95), .C1(n7506), .C2(keyinput99), 
        .A(n12340), .ZN(n12341) );
  NOR2_X1 U14978 ( .A1(n12342), .A2(n12341), .ZN(n12351) );
  AOI22_X1 U14979 ( .A1(n12344), .A2(keyinput31), .B1(keyinput11), .B2(n12509), 
        .ZN(n12343) );
  OAI221_X1 U14980 ( .B1(n12344), .B2(keyinput31), .C1(n12509), .C2(keyinput11), .A(n12343), .ZN(n12349) );
  AOI22_X1 U14981 ( .A1(n12347), .A2(keyinput74), .B1(keyinput87), .B2(n12346), 
        .ZN(n12345) );
  OAI221_X1 U14982 ( .B1(n12347), .B2(keyinput74), .C1(n12346), .C2(keyinput87), .A(n12345), .ZN(n12348) );
  NOR2_X1 U14983 ( .A1(n12349), .A2(n12348), .ZN(n12350) );
  NAND3_X1 U14984 ( .A1(n12352), .A2(n12351), .A3(n12350), .ZN(n12368) );
  AOI22_X1 U14985 ( .A1(n12481), .A2(keyinput100), .B1(keyinput39), .B2(n12354), .ZN(n12353) );
  OAI221_X1 U14986 ( .B1(n12481), .B2(keyinput100), .C1(n12354), .C2(
        keyinput39), .A(n12353), .ZN(n12367) );
  INV_X1 U14987 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n15527) );
  AOI22_X1 U14988 ( .A1(n12479), .A2(keyinput117), .B1(keyinput81), .B2(n15527), .ZN(n12355) );
  OAI221_X1 U14989 ( .B1(n12479), .B2(keyinput117), .C1(n15527), .C2(
        keyinput81), .A(n12355), .ZN(n12366) );
  INV_X1 U14990 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n15787) );
  INV_X1 U14991 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n15553) );
  AOI22_X1 U14992 ( .A1(n15787), .A2(keyinput45), .B1(keyinput29), .B2(n15553), 
        .ZN(n12356) );
  OAI221_X1 U14993 ( .B1(n15787), .B2(keyinput45), .C1(n15553), .C2(keyinput29), .A(n12356), .ZN(n12364) );
  AOI22_X1 U14994 ( .A1(n12359), .A2(keyinput104), .B1(keyinput5), .B2(n12358), 
        .ZN(n12357) );
  OAI221_X1 U14995 ( .B1(n12359), .B2(keyinput104), .C1(n12358), .C2(keyinput5), .A(n12357), .ZN(n12363) );
  INV_X1 U14996 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U14997 ( .A1(n14672), .A2(keyinput98), .B1(keyinput7), .B2(n12361), 
        .ZN(n12360) );
  OAI221_X1 U14998 ( .B1(n14672), .B2(keyinput98), .C1(n12361), .C2(keyinput7), 
        .A(n12360), .ZN(n12362) );
  OR3_X1 U14999 ( .A1(n12364), .A2(n12363), .A3(n12362), .ZN(n12365) );
  NOR4_X1 U15000 ( .A1(n12368), .A2(n12367), .A3(n12366), .A4(n12365), .ZN(
        n12408) );
  INV_X1 U15001 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15910) );
  AOI22_X1 U15002 ( .A1(n15910), .A2(keyinput61), .B1(keyinput106), .B2(n12468), .ZN(n12369) );
  OAI221_X1 U15003 ( .B1(n15910), .B2(keyinput61), .C1(n12468), .C2(
        keyinput106), .A(n12369), .ZN(n12385) );
  AOI22_X1 U15004 ( .A1(n14916), .A2(keyinput124), .B1(n12520), .B2(
        keyinput119), .ZN(n12373) );
  XNOR2_X1 U15005 ( .A(SI_7_), .B(keyinput85), .ZN(n12372) );
  XNOR2_X1 U15006 ( .A(SI_5_), .B(keyinput68), .ZN(n12371) );
  XNOR2_X1 U15007 ( .A(SI_1_), .B(keyinput84), .ZN(n12370) );
  NAND4_X1 U15008 ( .A1(n12373), .A2(n12372), .A3(n12371), .A4(n12370), .ZN(
        n12384) );
  XNOR2_X1 U15009 ( .A(SI_3_), .B(keyinput72), .ZN(n12377) );
  XNOR2_X1 U15010 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput12), .ZN(n12376) );
  XNOR2_X1 U15011 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput9), .ZN(n12375) );
  XNOR2_X1 U15012 ( .A(P1_REG0_REG_12__SCAN_IN), .B(keyinput10), .ZN(n12374)
         );
  NAND4_X1 U15013 ( .A1(n12377), .A2(n12376), .A3(n12375), .A4(n12374), .ZN(
        n12383) );
  XNOR2_X1 U15014 ( .A(P2_IR_REG_0__SCAN_IN), .B(keyinput24), .ZN(n12381) );
  XNOR2_X1 U15015 ( .A(P1_REG1_REG_26__SCAN_IN), .B(keyinput2), .ZN(n12380) );
  XNOR2_X1 U15016 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput25), .ZN(n12379) );
  XNOR2_X1 U15017 ( .A(P2_IR_REG_17__SCAN_IN), .B(keyinput6), .ZN(n12378) );
  NAND4_X1 U15018 ( .A1(n12381), .A2(n12380), .A3(n12379), .A4(n12378), .ZN(
        n12382) );
  NOR4_X1 U15019 ( .A1(n12385), .A2(n12384), .A3(n12383), .A4(n12382), .ZN(
        n12407) );
  XNOR2_X1 U15020 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput83), .ZN(n12389) );
  XNOR2_X1 U15021 ( .A(P2_IR_REG_27__SCAN_IN), .B(keyinput34), .ZN(n12388) );
  XNOR2_X1 U15022 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput56), .ZN(n12387) );
  XNOR2_X1 U15023 ( .A(P2_IR_REG_30__SCAN_IN), .B(keyinput46), .ZN(n12386) );
  NAND4_X1 U15024 ( .A1(n12389), .A2(n12388), .A3(n12387), .A4(n12386), .ZN(
        n12405) );
  XNOR2_X1 U15025 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput63), .ZN(n12393)
         );
  XNOR2_X1 U15026 ( .A(P2_REG0_REG_17__SCAN_IN), .B(keyinput90), .ZN(n12392)
         );
  XNOR2_X1 U15027 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput58), .ZN(n12391)
         );
  XNOR2_X1 U15028 ( .A(P3_IR_REG_27__SCAN_IN), .B(keyinput16), .ZN(n12390) );
  NAND4_X1 U15029 ( .A1(n12393), .A2(n12392), .A3(n12391), .A4(n12390), .ZN(
        n12404) );
  XNOR2_X1 U15030 ( .A(P3_IR_REG_17__SCAN_IN), .B(keyinput22), .ZN(n12397) );
  XNOR2_X1 U15031 ( .A(P3_REG0_REG_24__SCAN_IN), .B(keyinput49), .ZN(n12396)
         );
  XNOR2_X1 U15032 ( .A(P3_REG0_REG_10__SCAN_IN), .B(keyinput70), .ZN(n12395)
         );
  XNOR2_X1 U15033 ( .A(P3_REG1_REG_30__SCAN_IN), .B(keyinput77), .ZN(n12394)
         );
  NAND4_X1 U15034 ( .A1(n12397), .A2(n12396), .A3(n12395), .A4(n12394), .ZN(
        n12403) );
  XNOR2_X1 U15035 ( .A(P1_REG0_REG_10__SCAN_IN), .B(keyinput114), .ZN(n12401)
         );
  XNOR2_X1 U15036 ( .A(P3_IR_REG_15__SCAN_IN), .B(keyinput118), .ZN(n12400) );
  XNOR2_X1 U15037 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput105), .ZN(n12399)
         );
  XNOR2_X1 U15038 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(keyinput111), .ZN(n12398)
         );
  NAND4_X1 U15039 ( .A1(n12401), .A2(n12400), .A3(n12399), .A4(n12398), .ZN(
        n12402) );
  NOR4_X1 U15040 ( .A1(n12405), .A2(n12404), .A3(n12403), .A4(n12402), .ZN(
        n12406) );
  NAND4_X1 U15041 ( .A1(n12409), .A2(n12408), .A3(n12407), .A4(n12406), .ZN(
        n12410) );
  NOR3_X1 U15042 ( .A1(n12412), .A2(n12411), .A3(n12410), .ZN(n12449) );
  AOI22_X1 U15043 ( .A1(n9075), .A2(keyinput26), .B1(keyinput60), .B2(n12559), 
        .ZN(n12413) );
  OAI221_X1 U15044 ( .B1(n9075), .B2(keyinput26), .C1(n12559), .C2(keyinput60), 
        .A(n12413), .ZN(n12424) );
  INV_X1 U15045 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15526) );
  AOI22_X1 U15046 ( .A1(n15526), .A2(keyinput96), .B1(keyinput18), .B2(n12415), 
        .ZN(n12414) );
  OAI221_X1 U15047 ( .B1(n15526), .B2(keyinput96), .C1(n12415), .C2(keyinput18), .A(n12414), .ZN(n12423) );
  AOI22_X1 U15048 ( .A1(n12418), .A2(keyinput89), .B1(n12417), .B2(keyinput38), 
        .ZN(n12416) );
  OAI221_X1 U15049 ( .B1(n12418), .B2(keyinput89), .C1(n12417), .C2(keyinput38), .A(n12416), .ZN(n12422) );
  INV_X1 U15050 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n13188) );
  AOI22_X1 U15051 ( .A1(n12420), .A2(keyinput64), .B1(keyinput13), .B2(n13188), 
        .ZN(n12419) );
  OAI221_X1 U15052 ( .B1(n12420), .B2(keyinput64), .C1(n13188), .C2(keyinput13), .A(n12419), .ZN(n12421) );
  NOR4_X1 U15053 ( .A1(n12424), .A2(n12423), .A3(n12422), .A4(n12421), .ZN(
        n12448) );
  NAND2_X1 U15054 ( .A1(n12426), .A2(keyinput42), .ZN(n12425) );
  OAI221_X1 U15055 ( .B1(n14916), .B2(keyinput124), .C1(n12426), .C2(
        keyinput42), .A(n12425), .ZN(n12435) );
  AOI22_X1 U15056 ( .A1(n13463), .A2(keyinput79), .B1(keyinput103), .B2(n12080), .ZN(n12427) );
  OAI221_X1 U15057 ( .B1(n13463), .B2(keyinput79), .C1(n12080), .C2(
        keyinput103), .A(n12427), .ZN(n12434) );
  INV_X1 U15058 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n12429) );
  AOI22_X1 U15059 ( .A1(n12429), .A2(keyinput36), .B1(n8622), .B2(keyinput3), 
        .ZN(n12428) );
  OAI221_X1 U15060 ( .B1(n12429), .B2(keyinput36), .C1(n8622), .C2(keyinput3), 
        .A(n12428), .ZN(n12433) );
  INV_X1 U15061 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n15693) );
  AOI22_X1 U15062 ( .A1(n15693), .A2(keyinput52), .B1(n12431), .B2(keyinput19), 
        .ZN(n12430) );
  OAI221_X1 U15063 ( .B1(n15693), .B2(keyinput52), .C1(n12431), .C2(keyinput19), .A(n12430), .ZN(n12432) );
  NOR4_X1 U15064 ( .A1(n12435), .A2(n12434), .A3(n12433), .A4(n12432), .ZN(
        n12447) );
  AOI22_X1 U15065 ( .A1(n10555), .A2(keyinput17), .B1(n13351), .B2(keyinput127), .ZN(n12436) );
  OAI221_X1 U15066 ( .B1(n10555), .B2(keyinput17), .C1(n13351), .C2(
        keyinput127), .A(n12436), .ZN(n12445) );
  INV_X1 U15067 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n12467) );
  AOI22_X1 U15068 ( .A1(n12467), .A2(keyinput0), .B1(keyinput88), .B2(n12438), 
        .ZN(n12437) );
  OAI221_X1 U15069 ( .B1(n12467), .B2(keyinput0), .C1(n12438), .C2(keyinput88), 
        .A(n12437), .ZN(n12444) );
  AOI22_X1 U15070 ( .A1(n13460), .A2(keyinput47), .B1(keyinput50), .B2(n13143), 
        .ZN(n12439) );
  OAI221_X1 U15071 ( .B1(n13460), .B2(keyinput47), .C1(n13143), .C2(keyinput50), .A(n12439), .ZN(n12443) );
  AOI22_X1 U15072 ( .A1(n12441), .A2(keyinput97), .B1(keyinput51), .B2(n12476), 
        .ZN(n12440) );
  OAI221_X1 U15073 ( .B1(n12441), .B2(keyinput97), .C1(n12476), .C2(keyinput51), .A(n12440), .ZN(n12442) );
  NOR4_X1 U15074 ( .A1(n12445), .A2(n12444), .A3(n12443), .A4(n12442), .ZN(
        n12446) );
  NAND4_X1 U15075 ( .A1(n12449), .A2(n12448), .A3(n12447), .A4(n12446), .ZN(
        n12523) );
  NAND4_X1 U15076 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_REG1_REG_4__SCAN_IN), 
        .A3(P3_REG2_REG_31__SCAN_IN), .A4(P3_DATAO_REG_2__SCAN_IN), .ZN(n12450) );
  NOR3_X1 U15077 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n12451), .A3(n12450), 
        .ZN(n12464) );
  NAND4_X1 U15078 ( .A1(SI_1_), .A2(SI_3_), .A3(SI_5_), .A4(SI_7_), .ZN(n12453) );
  OR3_X1 U15079 ( .A1(n12453), .A2(P3_REG1_REG_3__SCAN_IN), .A3(n12452), .ZN(
        n12461) );
  NOR4_X1 U15080 ( .A1(P3_REG1_REG_30__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), 
        .A3(n8622), .A4(n15705), .ZN(n12459) );
  NOR4_X1 U15081 ( .A1(P3_REG1_REG_19__SCAN_IN), .A2(P2_REG2_REG_9__SCAN_IN), 
        .A3(P2_REG1_REG_3__SCAN_IN), .A4(P2_ADDR_REG_10__SCAN_IN), .ZN(n12458)
         );
  NOR4_X1 U15082 ( .A1(P3_REG2_REG_24__SCAN_IN), .A2(P3_REG2_REG_30__SCAN_IN), 
        .A3(P2_IR_REG_9__SCAN_IN), .A4(n12454), .ZN(n12457) );
  NOR4_X1 U15083 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(P2_REG2_REG_4__SCAN_IN), 
        .A3(P1_REG1_REG_26__SCAN_IN), .A4(n12455), .ZN(n12456) );
  NAND4_X1 U15084 ( .A1(n12459), .A2(n12458), .A3(n12457), .A4(n12456), .ZN(
        n12460) );
  NOR4_X1 U15085 ( .A1(P3_REG0_REG_10__SCAN_IN), .A2(n12462), .A3(n12461), 
        .A4(n12460), .ZN(n12463) );
  NAND4_X1 U15086 ( .A1(P3_REG0_REG_23__SCAN_IN), .A2(P2_REG2_REG_3__SCAN_IN), 
        .A3(n12464), .A4(n12463), .ZN(n12519) );
  NOR2_X1 U15087 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), 
        .ZN(n12466) );
  NOR4_X1 U15088 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(P3_ADDR_REG_1__SCAN_IN), 
        .A3(n12559), .A4(n9723), .ZN(n12465) );
  NAND4_X1 U15089 ( .A1(n12466), .A2(P2_ADDR_REG_3__SCAN_IN), .A3(
        P3_ADDR_REG_3__SCAN_IN), .A4(n12465), .ZN(n12474) );
  NOR4_X1 U15090 ( .A1(P3_REG1_REG_20__SCAN_IN), .A2(P1_REG2_REG_13__SCAN_IN), 
        .A3(P3_ADDR_REG_17__SCAN_IN), .A4(n10380), .ZN(n12472) );
  NOR4_X1 U15091 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P3_REG2_REG_17__SCAN_IN), 
        .A3(n12467), .A4(n10555), .ZN(n12471) );
  NOR4_X1 U15092 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .A3(P1_IR_REG_26__SCAN_IN), .A4(n12468), .ZN(n12470) );
  NOR4_X1 U15093 ( .A1(SI_28_), .A2(P2_IR_REG_27__SCAN_IN), .A3(
        P2_REG3_REG_3__SCAN_IN), .A4(P2_REG2_REG_11__SCAN_IN), .ZN(n12469) );
  NAND4_X1 U15094 ( .A1(n12472), .A2(n12471), .A3(n12470), .A4(n12469), .ZN(
        n12473) );
  NOR2_X1 U15095 ( .A1(n12474), .A2(n12473), .ZN(n12503) );
  NAND4_X1 U15096 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), 
        .A3(n13517), .A4(n12475), .ZN(n12478) );
  NAND4_X1 U15097 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), 
        .A3(P3_REG3_REG_3__SCAN_IN), .A4(n12476), .ZN(n12477) );
  NOR2_X1 U15098 ( .A1(n12478), .A2(n12477), .ZN(n12501) );
  NOR4_X1 U15099 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_21__SCAN_IN), 
        .A3(P1_REG0_REG_14__SCAN_IN), .A4(P3_DATAO_REG_24__SCAN_IN), .ZN(
        n12480) );
  NAND3_X1 U15100 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n12480), .A3(n12479), .ZN(
        n12499) );
  AND4_X1 U15101 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_17__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(n12481), .ZN(n12497) );
  NAND4_X1 U15102 ( .A1(n12483), .A2(n12482), .A3(n14670), .A4(
        P2_REG3_REG_7__SCAN_IN), .ZN(n12488) );
  INV_X1 U15103 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n12486) );
  NOR4_X1 U15104 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(P1_REG1_REG_2__SCAN_IN), 
        .A3(n12484), .A4(n13790), .ZN(n12485) );
  NAND4_X1 U15105 ( .A1(n15786), .A2(n12486), .A3(n12485), .A4(
        P1_REG0_REG_2__SCAN_IN), .ZN(n12487) );
  NOR2_X1 U15106 ( .A1(n12488), .A2(n12487), .ZN(n12496) );
  NAND4_X1 U15107 ( .A1(n12489), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P1_DATAO_REG_26__SCAN_IN), .A4(P3_IR_REG_15__SCAN_IN), .ZN(n12491) );
  NAND4_X1 U15108 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(P2_DATAO_REG_11__SCAN_IN), .A3(P3_REG3_REG_26__SCAN_IN), .A4(P3_IR_REG_0__SCAN_IN), .ZN(n12490) );
  NOR2_X1 U15109 ( .A1(n12491), .A2(n12490), .ZN(n12495) );
  NAND4_X1 U15110 ( .A1(n14916), .A2(n15787), .A3(P1_REG0_REG_10__SCAN_IN), 
        .A4(P1_REG0_REG_15__SCAN_IN), .ZN(n12493) );
  NAND4_X1 U15111 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .A3(P1_REG3_REG_7__SCAN_IN), .A4(P3_REG3_REG_19__SCAN_IN), .ZN(n12492)
         );
  NOR2_X1 U15112 ( .A1(n12493), .A2(n12492), .ZN(n12494) );
  NAND4_X1 U15113 ( .A1(n12497), .A2(n12496), .A3(n12495), .A4(n12494), .ZN(
        n12498) );
  NOR2_X1 U15114 ( .A1(n12499), .A2(n12498), .ZN(n12500) );
  AND4_X1 U15115 ( .A1(n12503), .A2(n12502), .A3(n12501), .A4(n12500), .ZN(
        n12507) );
  NOR4_X1 U15116 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), 
        .A3(P3_DATAO_REG_0__SCAN_IN), .A4(n15811), .ZN(n12506) );
  NOR4_X1 U15117 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(P1_REG1_REG_6__SCAN_IN), 
        .A3(P3_DATAO_REG_29__SCAN_IN), .A4(n12504), .ZN(n12505) );
  NAND3_X1 U15118 ( .A1(n12507), .A2(n12506), .A3(n12505), .ZN(n12518) );
  INV_X1 U15119 ( .A(n12508), .ZN(n12517) );
  NOR4_X1 U15120 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(n12510), .A3(n12509), .A4(
        n8353), .ZN(n12515) );
  NOR4_X1 U15121 ( .A1(P3_REG2_REG_26__SCAN_IN), .A2(P3_DATAO_REG_23__SCAN_IN), 
        .A3(n12512), .A4(n12511), .ZN(n12514) );
  INV_X1 U15122 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n14637) );
  NOR4_X1 U15123 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(P1_REG2_REG_30__SCAN_IN), 
        .A3(P1_ADDR_REG_11__SCAN_IN), .A4(n14637), .ZN(n12513) );
  NAND3_X1 U15124 ( .A1(n12515), .A2(n12514), .A3(n12513), .ZN(n12516) );
  OR4_X1 U15125 ( .A1(n12519), .A2(n12518), .A3(n12517), .A4(n12516), .ZN(
        n12521) );
  AOI21_X1 U15126 ( .B1(n12521), .B2(keyinput119), .A(n12520), .ZN(n12522) );
  NOR2_X1 U15127 ( .A1(n12523), .A2(n12522), .ZN(n12524) );
  XNOR2_X1 U15128 ( .A(n12525), .B(n12524), .ZN(P3_U3174) );
  AOI22_X1 U15129 ( .A1(n12528), .A2(n13034), .B1(n12527), .B2(n12526), .ZN(
        n12533) );
  OAI21_X1 U15130 ( .B1(n12531), .B2(n12530), .A(n12529), .ZN(n12532) );
  XNOR2_X1 U15131 ( .A(n12533), .B(n12532), .ZN(n12539) );
  INV_X1 U15132 ( .A(n12954), .ZN(n13484) );
  INV_X1 U15133 ( .A(n12836), .ZN(n12798) );
  NAND2_X1 U15134 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n13049)
         );
  OAI21_X1 U15135 ( .B1(n12822), .B2(n13403), .A(n13049), .ZN(n12534) );
  AOI21_X1 U15136 ( .B1(n12798), .B2(n13034), .A(n12534), .ZN(n12535) );
  OAI21_X1 U15137 ( .B1(n12536), .B2(n13409), .A(n12535), .ZN(n12537) );
  AOI21_X1 U15138 ( .B1(n13484), .B2(n12803), .A(n12537), .ZN(n12538) );
  OAI21_X1 U15139 ( .B1(n12539), .B2(n12815), .A(n12538), .ZN(P3_U3164) );
  XNOR2_X1 U15140 ( .A(n12541), .B(n12540), .ZN(n12546) );
  NAND2_X1 U15141 ( .A1(n12839), .A2(n13385), .ZN(n12543) );
  AND2_X1 U15142 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n13092) );
  AOI21_X1 U15143 ( .B1(n12834), .B2(n13382), .A(n13092), .ZN(n12542) );
  OAI211_X1 U15144 ( .C1(n13403), .C2(n12836), .A(n12543), .B(n12542), .ZN(
        n12544) );
  AOI21_X1 U15145 ( .B1(n13574), .B2(n12803), .A(n12544), .ZN(n12545) );
  OAI21_X1 U15146 ( .B1(n12546), .B2(n12815), .A(n12545), .ZN(P3_U3155) );
  INV_X1 U15147 ( .A(n12547), .ZN(n12566) );
  OAI222_X1 U15148 ( .A1(n14671), .A2(n12549), .B1(n14673), .B2(n12566), .C1(
        P2_U3088), .C2(n12548), .ZN(P2_U3302) );
  AND2_X1 U15149 ( .A1(n12684), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12551) );
  NAND2_X1 U15150 ( .A1(n14667), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12550) );
  XNOR2_X1 U15151 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n12705) );
  INV_X1 U15152 ( .A(n12705), .ZN(n12553) );
  NAND2_X1 U15153 ( .A1(n12559), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12848) );
  NAND2_X1 U15154 ( .A1(n15429), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12554) );
  NAND2_X1 U15155 ( .A1(n12848), .A2(n12554), .ZN(n12849) );
  XNOR2_X1 U15156 ( .A(n12850), .B(n12849), .ZN(n12844) );
  INV_X1 U15157 ( .A(n12844), .ZN(n12556) );
  OAI222_X1 U15158 ( .A1(n12557), .A2(P3_U3151), .B1(n13611), .B2(n12556), 
        .C1(n12555), .C2(n13618), .ZN(P3_U3265) );
  INV_X1 U15159 ( .A(n12558), .ZN(n15428) );
  OAI222_X1 U15160 ( .A1(n14673), .A2(n15428), .B1(n11242), .B2(n12560), .C1(
        n12559), .C2(n14671), .ZN(P2_U3297) );
  NOR2_X1 U15161 ( .A1(n15783), .A2(n14490), .ZN(n14180) );
  NOR2_X1 U15162 ( .A1(n12561), .A2(n14436), .ZN(n12562) );
  AOI211_X1 U15163 ( .C1(n15783), .C2(P2_REG2_REG_31__SCAN_IN), .A(n14180), 
        .B(n12562), .ZN(n12563) );
  OAI21_X1 U15164 ( .B1(n12564), .B2(n14461), .A(n12563), .ZN(P2_U3234) );
  OAI222_X1 U15165 ( .A1(n15435), .A2(n12567), .B1(n15438), .B2(n12566), .C1(
        n12565), .C2(P1_U3086), .ZN(P1_U3330) );
  INV_X1 U15166 ( .A(n12568), .ZN(n12569) );
  OAI222_X1 U15167 ( .A1(n9503), .A2(P3_U3151), .B1(n13618), .B2(n12570), .C1(
        n13622), .C2(n12569), .ZN(P3_U3267) );
  XNOR2_X1 U15168 ( .A(n13194), .B(n12571), .ZN(n12578) );
  INV_X1 U15169 ( .A(n12578), .ZN(n12572) );
  NAND2_X1 U15170 ( .A1(n12572), .A2(n12832), .ZN(n12584) );
  INV_X1 U15171 ( .A(n12573), .ZN(n12574) );
  NAND4_X1 U15172 ( .A1(n12583), .A2(n12832), .A3(n12574), .A4(n12578), .ZN(
        n12582) );
  AOI22_X1 U15173 ( .A1(n12700), .A2(n12839), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12576) );
  NAND2_X1 U15174 ( .A1(n13217), .A2(n12798), .ZN(n12575) );
  OAI211_X1 U15175 ( .C1(n12868), .C2(n12822), .A(n12576), .B(n12575), .ZN(
        n12580) );
  NOR4_X1 U15176 ( .A1(n12578), .A2(n12577), .A3(n12815), .A4(n13217), .ZN(
        n12579) );
  AOI211_X1 U15177 ( .C1(n12803), .C2(n13196), .A(n12580), .B(n12579), .ZN(
        n12581) );
  OAI211_X1 U15178 ( .C1(n12584), .C2(n12583), .A(n12582), .B(n12581), .ZN(
        P3_U3160) );
  INV_X1 U15179 ( .A(n12585), .ZN(n12589) );
  NAND2_X1 U15180 ( .A1(n12586), .A2(n13798), .ZN(n12587) );
  OAI21_X1 U15181 ( .B1(n13865), .B2(n13758), .A(n12587), .ZN(n12588) );
  NAND3_X1 U15182 ( .A1(n12721), .A2(n12589), .A3(n12588), .ZN(n12595) );
  NAND2_X1 U15183 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n15678) );
  INV_X1 U15184 ( .A(n15678), .ZN(n12590) );
  AOI21_X1 U15185 ( .B1(n13769), .B2(n14095), .A(n12590), .ZN(n12594) );
  AOI22_X1 U15186 ( .A1(n13770), .A2(n14096), .B1(n13750), .B2(n12591), .ZN(
        n12593) );
  NAND2_X1 U15187 ( .A1(n13870), .A2(n13808), .ZN(n12592) );
  AND4_X1 U15188 ( .A1(n12595), .A2(n12594), .A3(n12593), .A4(n12592), .ZN(
        n12596) );
  OAI21_X1 U15189 ( .B1(n12597), .B2(n13796), .A(n12596), .ZN(P2_U3203) );
  NAND2_X1 U15190 ( .A1(n14088), .A2(n14481), .ZN(n12664) );
  XNOR2_X1 U15191 ( .A(n14217), .B(n12669), .ZN(n12666) );
  XNOR2_X1 U15192 ( .A(n14588), .B(n11713), .ZN(n12601) );
  NAND2_X1 U15193 ( .A1(n14481), .A2(n14094), .ZN(n12602) );
  NAND2_X1 U15194 ( .A1(n12601), .A2(n12602), .ZN(n12606) );
  INV_X1 U15195 ( .A(n12601), .ZN(n12604) );
  INV_X1 U15196 ( .A(n12602), .ZN(n12603) );
  NAND2_X1 U15197 ( .A1(n12604), .A2(n12603), .ZN(n12605) );
  AND2_X1 U15198 ( .A1(n12606), .A2(n12605), .ZN(n13678) );
  INV_X1 U15199 ( .A(n13740), .ZN(n12608) );
  XNOR2_X1 U15200 ( .A(n14432), .B(n11713), .ZN(n12609) );
  NAND2_X1 U15201 ( .A1(n14481), .A2(n14448), .ZN(n12610) );
  XNOR2_X1 U15202 ( .A(n12609), .B(n12610), .ZN(n13739) );
  INV_X1 U15203 ( .A(n13739), .ZN(n12607) );
  INV_X1 U15204 ( .A(n12609), .ZN(n12612) );
  INV_X1 U15205 ( .A(n12610), .ZN(n12611) );
  NAND2_X1 U15206 ( .A1(n12612), .A2(n12611), .ZN(n13633) );
  NAND2_X1 U15207 ( .A1(n14481), .A2(n14397), .ZN(n12614) );
  NAND2_X1 U15208 ( .A1(n12613), .A2(n12614), .ZN(n12619) );
  INV_X1 U15209 ( .A(n12613), .ZN(n12616) );
  INV_X1 U15210 ( .A(n12614), .ZN(n12615) );
  NAND2_X1 U15211 ( .A1(n12616), .A2(n12615), .ZN(n12617) );
  AND2_X1 U15212 ( .A1(n14481), .A2(n14093), .ZN(n12623) );
  XNOR2_X1 U15213 ( .A(n14393), .B(n12669), .ZN(n12621) );
  XNOR2_X1 U15214 ( .A(n14568), .B(n12669), .ZN(n12624) );
  AND2_X1 U15215 ( .A1(n14398), .A2(n14481), .ZN(n12625) );
  AND2_X1 U15216 ( .A1(n12624), .A2(n12625), .ZN(n12622) );
  INV_X1 U15217 ( .A(n12621), .ZN(n13699) );
  INV_X1 U15218 ( .A(n12622), .ZN(n13697) );
  INV_X1 U15219 ( .A(n12623), .ZN(n13797) );
  INV_X1 U15220 ( .A(n12624), .ZN(n12627) );
  INV_X1 U15221 ( .A(n12625), .ZN(n12626) );
  NAND2_X1 U15222 ( .A1(n12627), .A2(n12626), .ZN(n13696) );
  XNOR2_X1 U15223 ( .A(n14364), .B(n11713), .ZN(n12629) );
  NAND2_X1 U15224 ( .A1(n14339), .A2(n14481), .ZN(n12630) );
  NAND2_X1 U15225 ( .A1(n12629), .A2(n12630), .ZN(n12634) );
  INV_X1 U15226 ( .A(n12629), .ZN(n12632) );
  INV_X1 U15227 ( .A(n12630), .ZN(n12631) );
  NAND2_X1 U15228 ( .A1(n12632), .A2(n12631), .ZN(n12633) );
  AND2_X1 U15229 ( .A1(n12634), .A2(n12633), .ZN(n13708) );
  XNOR2_X1 U15230 ( .A(n14351), .B(n11713), .ZN(n12635) );
  NAND2_X1 U15231 ( .A1(n14092), .A2(n14481), .ZN(n12636) );
  XNOR2_X1 U15232 ( .A(n12635), .B(n12636), .ZN(n13775) );
  INV_X1 U15233 ( .A(n12635), .ZN(n12638) );
  INV_X1 U15234 ( .A(n12636), .ZN(n12637) );
  NAND2_X1 U15235 ( .A1(n12638), .A2(n12637), .ZN(n12639) );
  NAND2_X1 U15236 ( .A1(n14091), .A2(n14481), .ZN(n12646) );
  XNOR2_X1 U15237 ( .A(n12648), .B(n12646), .ZN(n13669) );
  XNOR2_X1 U15238 ( .A(n14544), .B(n11713), .ZN(n13662) );
  OR2_X1 U15239 ( .A1(n13909), .A2(n15767), .ZN(n13661) );
  NAND2_X1 U15240 ( .A1(n13662), .A2(n13661), .ZN(n13666) );
  NAND2_X1 U15241 ( .A1(n14340), .A2(n14481), .ZN(n13663) );
  NAND2_X1 U15242 ( .A1(n13726), .A2(n13663), .ZN(n12640) );
  AND3_X1 U15243 ( .A1(n13666), .A2(n13669), .A3(n12640), .ZN(n12645) );
  INV_X1 U15244 ( .A(n13663), .ZN(n13655) );
  INV_X1 U15245 ( .A(n13726), .ZN(n13665) );
  INV_X1 U15246 ( .A(n13662), .ZN(n12642) );
  INV_X1 U15247 ( .A(n13661), .ZN(n12641) );
  NAND2_X1 U15248 ( .A1(n12642), .A2(n12641), .ZN(n12643) );
  INV_X1 U15249 ( .A(n12646), .ZN(n12647) );
  NAND2_X1 U15250 ( .A1(n12648), .A2(n12647), .ZN(n12649) );
  XNOR2_X1 U15251 ( .A(n14284), .B(n12669), .ZN(n12652) );
  XNOR2_X1 U15252 ( .A(n14528), .B(n11713), .ZN(n12654) );
  NAND2_X1 U15253 ( .A1(n12654), .A2(n13717), .ZN(n12651) );
  NAND2_X1 U15254 ( .A1(n14263), .A2(n14481), .ZN(n13644) );
  INV_X1 U15255 ( .A(n13644), .ZN(n12650) );
  NAND2_X1 U15256 ( .A1(n12651), .A2(n12650), .ZN(n12657) );
  NAND2_X1 U15257 ( .A1(n14090), .A2(n14481), .ZN(n13649) );
  INV_X1 U15258 ( .A(n12654), .ZN(n13646) );
  INV_X1 U15259 ( .A(n13649), .ZN(n12655) );
  XNOR2_X1 U15260 ( .A(n14522), .B(n12669), .ZN(n13685) );
  NOR2_X1 U15261 ( .A1(n14262), .A2(n15767), .ZN(n12658) );
  NAND2_X1 U15262 ( .A1(n13685), .A2(n12658), .ZN(n12659) );
  OAI21_X1 U15263 ( .B1(n13685), .B2(n12658), .A(n12659), .ZN(n13714) );
  XNOR2_X1 U15264 ( .A(n14234), .B(n11713), .ZN(n13781) );
  NOR2_X1 U15265 ( .A1(n13718), .A2(n15767), .ZN(n12660) );
  NAND2_X1 U15266 ( .A1(n13781), .A2(n12660), .ZN(n12665) );
  INV_X1 U15267 ( .A(n13781), .ZN(n12662) );
  INV_X1 U15268 ( .A(n12660), .ZN(n12661) );
  NAND2_X1 U15269 ( .A1(n12662), .A2(n12661), .ZN(n12663) );
  AND2_X1 U15270 ( .A1(n12665), .A2(n12663), .ZN(n13686) );
  XNOR2_X1 U15271 ( .A(n12666), .B(n12664), .ZN(n13784) );
  XNOR2_X1 U15272 ( .A(n13992), .B(n12669), .ZN(n12668) );
  NOR2_X1 U15273 ( .A1(n13993), .A2(n15767), .ZN(n12667) );
  NAND2_X1 U15274 ( .A1(n12668), .A2(n12667), .ZN(n12676) );
  OAI21_X1 U15275 ( .B1(n12668), .B2(n12667), .A(n12676), .ZN(n13624) );
  NOR2_X1 U15276 ( .A1(n14196), .A2(n15767), .ZN(n12670) );
  XNOR2_X1 U15277 ( .A(n12670), .B(n12669), .ZN(n12671) );
  XNOR2_X1 U15278 ( .A(n14184), .B(n12671), .ZN(n12672) );
  INV_X1 U15279 ( .A(n12672), .ZN(n12677) );
  NAND3_X1 U15280 ( .A1(n12677), .A2(n13798), .A3(n12676), .ZN(n12682) );
  INV_X1 U15281 ( .A(n12673), .ZN(n12675) );
  AOI22_X1 U15282 ( .A1(n14203), .A2(n13750), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12674) );
  OAI21_X1 U15283 ( .B1(n12675), .B2(n13789), .A(n12674), .ZN(n12679) );
  NOR3_X1 U15284 ( .A1(n12677), .A2(n12676), .A3(n13796), .ZN(n12678) );
  AOI211_X1 U15285 ( .C1(n14184), .C2(n13808), .A(n12679), .B(n12678), .ZN(
        n12680) );
  OAI211_X1 U15286 ( .C1(n13623), .C2(n12682), .A(n12681), .B(n12680), .ZN(
        P2_U3192) );
  INV_X1 U15287 ( .A(n10297), .ZN(n12683) );
  OAI222_X1 U15288 ( .A1(n15435), .A2(n12684), .B1(n15438), .B2(n12683), .C1(
        P1_U3086), .C2(n14874), .ZN(P1_U3327) );
  AOI22_X1 U15289 ( .A1(n12685), .A2(n15513), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n15262), .ZN(n12686) );
  OAI21_X1 U15290 ( .B1(n14983), .B2(n15517), .A(n12686), .ZN(n12687) );
  AOI21_X1 U15291 ( .B1(n8090), .B2(n15254), .A(n12687), .ZN(n12691) );
  NAND3_X1 U15292 ( .A1(n12689), .A2(n15242), .A3(n12688), .ZN(n12690) );
  OAI211_X1 U15293 ( .C1(n12692), .C2(n15262), .A(n12691), .B(n12690), .ZN(
        P1_U3265) );
  INV_X1 U15294 ( .A(n12693), .ZN(n12695) );
  INV_X1 U15295 ( .A(SI_24_), .ZN(n12694) );
  OAI222_X1 U15296 ( .A1(P3_U3151), .A2(n9558), .B1(n13611), .B2(n12695), .C1(
        n12694), .C2(n13618), .ZN(P3_U3271) );
  INV_X1 U15297 ( .A(n12696), .ZN(n15430) );
  OAI222_X1 U15298 ( .A1(n14673), .A2(n15430), .B1(n6510), .B2(n12698), .C1(
        n12697), .C2(n14671), .ZN(P2_U3298) );
  AOI22_X1 U15299 ( .A1(n12700), .A2(n13427), .B1(n15873), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12701) );
  OAI21_X1 U15300 ( .B1(n12702), .B2(n13266), .A(n12701), .ZN(n12703) );
  AOI21_X1 U15301 ( .B1(n6568), .B2(n13411), .A(n12703), .ZN(n12704) );
  OAI21_X1 U15302 ( .B1(n12699), .B2(n15873), .A(n12704), .ZN(P3_U3205) );
  XNOR2_X1 U15303 ( .A(n12706), .B(n12705), .ZN(n12862) );
  INV_X1 U15304 ( .A(n12862), .ZN(n12707) );
  OAI222_X1 U15305 ( .A1(n13618), .A2(n12708), .B1(n13611), .B2(n12707), .C1(
        P3_U3151), .C2(n9019), .ZN(P3_U3266) );
  NAND2_X1 U15306 ( .A1(n13769), .A2(n8009), .ZN(n12711) );
  NAND2_X1 U15307 ( .A1(n13770), .A2(n14097), .ZN(n12710) );
  NAND2_X1 U15308 ( .A1(n13750), .A2(n8087), .ZN(n12709) );
  NAND2_X1 U15309 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(n6510), .ZN(n15661) );
  NAND4_X1 U15310 ( .A1(n12711), .A2(n12710), .A3(n12709), .A4(n15661), .ZN(
        n12719) );
  INV_X1 U15311 ( .A(n12712), .ZN(n12715) );
  NOR3_X1 U15312 ( .A1(n13758), .A2(n12713), .A3(n13859), .ZN(n12714) );
  AOI21_X1 U15313 ( .B1(n12715), .B2(n13798), .A(n12714), .ZN(n12717) );
  NOR2_X1 U15314 ( .A1(n12717), .A2(n12716), .ZN(n12718) );
  AOI211_X1 U15315 ( .C1(n7205), .C2(n13808), .A(n12719), .B(n12718), .ZN(
        n12720) );
  OAI21_X1 U15316 ( .B1(n12721), .B2(n13796), .A(n12720), .ZN(P2_U3193) );
  INV_X1 U15317 ( .A(n12750), .ZN(n12723) );
  AOI21_X1 U15318 ( .B1(n13274), .B2(n12724), .A(n12781), .ZN(n12730) );
  AOI22_X1 U15319 ( .A1(n13289), .A2(n12798), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12726) );
  NAND2_X1 U15320 ( .A1(n13264), .A2(n12839), .ZN(n12725) );
  OAI211_X1 U15321 ( .C1(n13237), .C2(n12822), .A(n12726), .B(n12725), .ZN(
        n12727) );
  AOI21_X1 U15322 ( .B1(n12728), .B2(n12803), .A(n12727), .ZN(n12729) );
  OAI21_X1 U15323 ( .B1(n12730), .B2(n12815), .A(n12729), .ZN(P3_U3156) );
  XNOR2_X1 U15324 ( .A(n12731), .B(n13336), .ZN(n12732) );
  XNOR2_X1 U15325 ( .A(n12733), .B(n12732), .ZN(n12739) );
  NAND2_X1 U15326 ( .A1(n12798), .A2(n13349), .ZN(n12734) );
  NAND2_X1 U15327 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13169)
         );
  OAI211_X1 U15328 ( .C1(n13323), .C2(n12822), .A(n12734), .B(n13169), .ZN(
        n12737) );
  NOR2_X1 U15329 ( .A1(n12735), .A2(n12842), .ZN(n12736) );
  AOI211_X1 U15330 ( .C1(n13327), .C2(n12839), .A(n12737), .B(n12736), .ZN(
        n12738) );
  OAI21_X1 U15331 ( .B1(n12739), .B2(n12815), .A(n12738), .ZN(P3_U3159) );
  OAI21_X1 U15332 ( .B1(n12742), .B2(n12741), .A(n12740), .ZN(n12743) );
  NAND2_X1 U15333 ( .A1(n12743), .A2(n12832), .ZN(n12748) );
  AOI22_X1 U15334 ( .A1(n13288), .A2(n12798), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12744) );
  OAI21_X1 U15335 ( .B1(n12745), .B2(n12822), .A(n12744), .ZN(n12746) );
  AOI21_X1 U15336 ( .B1(n13292), .B2(n12839), .A(n12746), .ZN(n12747) );
  OAI211_X1 U15337 ( .C1(n6798), .C2(n12842), .A(n12748), .B(n12747), .ZN(
        P3_U3163) );
  AOI21_X1 U15338 ( .B1(n12750), .B2(n12749), .A(n6530), .ZN(n12782) );
  NOR3_X1 U15339 ( .A1(n12782), .A2(n7967), .A3(n12751), .ZN(n12754) );
  INV_X1 U15340 ( .A(n12752), .ZN(n12753) );
  OAI21_X1 U15341 ( .B1(n12754), .B2(n12753), .A(n12832), .ZN(n12759) );
  AOI22_X1 U15342 ( .A1(n13259), .A2(n12798), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12755) );
  OAI21_X1 U15343 ( .B1(n12756), .B2(n12822), .A(n12755), .ZN(n12757) );
  AOI21_X1 U15344 ( .B1(n13238), .B2(n12839), .A(n12757), .ZN(n12758) );
  OAI211_X1 U15345 ( .C1(n13240), .C2(n12842), .A(n12759), .B(n12758), .ZN(
        P3_U3165) );
  AND3_X1 U15346 ( .A1(n12829), .A2(n12761), .A3(n12760), .ZN(n12762) );
  OAI21_X1 U15347 ( .B1(n12763), .B2(n12762), .A(n12832), .ZN(n12768) );
  NAND2_X1 U15348 ( .A1(n12834), .A2(n13358), .ZN(n12764) );
  NAND2_X1 U15349 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13122)
         );
  OAI211_X1 U15350 ( .C1(n12765), .C2(n12836), .A(n12764), .B(n13122), .ZN(
        n12766) );
  AOI21_X1 U15351 ( .B1(n13361), .B2(n12839), .A(n12766), .ZN(n12767) );
  OAI211_X1 U15352 ( .C1(n12769), .C2(n12842), .A(n12768), .B(n12767), .ZN(
        P3_U3166) );
  OAI211_X1 U15353 ( .C1(n12772), .C2(n12771), .A(n12770), .B(n12832), .ZN(
        n12777) );
  NAND2_X1 U15354 ( .A1(n12834), .A2(n13349), .ZN(n12773) );
  NAND2_X1 U15355 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13142)
         );
  OAI211_X1 U15356 ( .C1(n12774), .C2(n12836), .A(n12773), .B(n13142), .ZN(
        n12775) );
  AOI21_X1 U15357 ( .B1(n13352), .B2(n12839), .A(n12775), .ZN(n12776) );
  OAI211_X1 U15358 ( .C1(n12778), .C2(n12842), .A(n12777), .B(n12776), .ZN(
        P3_U3168) );
  OAI22_X1 U15359 ( .A1(n12801), .A2(n12836), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12783), .ZN(n12785) );
  NOR2_X1 U15360 ( .A1(n13249), .A2(n12822), .ZN(n12784) );
  AOI211_X1 U15361 ( .C1(n13252), .C2(n12839), .A(n12785), .B(n12784), .ZN(
        n12786) );
  OAI211_X1 U15362 ( .C1(n13519), .C2(n12842), .A(n12787), .B(n12786), .ZN(
        P3_U3169) );
  XNOR2_X1 U15363 ( .A(n12789), .B(n12788), .ZN(n12795) );
  AOI22_X1 U15364 ( .A1(n6797), .A2(n12834), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12791) );
  NAND2_X1 U15365 ( .A1(n12839), .A2(n13311), .ZN(n12790) );
  OAI211_X1 U15366 ( .C1(n12792), .C2(n12836), .A(n12791), .B(n12790), .ZN(
        n12793) );
  AOI21_X1 U15367 ( .B1(n13538), .B2(n12803), .A(n12793), .ZN(n12794) );
  OAI21_X1 U15368 ( .B1(n12795), .B2(n12815), .A(n12794), .ZN(P3_U3173) );
  AOI21_X1 U15369 ( .B1(n13289), .B2(n12797), .A(n12796), .ZN(n12805) );
  AOI22_X1 U15370 ( .A1(n6797), .A2(n12798), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12800) );
  NAND2_X1 U15371 ( .A1(n13277), .A2(n12839), .ZN(n12799) );
  OAI211_X1 U15372 ( .C1(n12801), .C2(n12822), .A(n12800), .B(n12799), .ZN(
        n12802) );
  AOI21_X1 U15373 ( .B1(n13526), .B2(n12803), .A(n12802), .ZN(n12804) );
  OAI21_X1 U15374 ( .B1(n12805), .B2(n12815), .A(n12804), .ZN(P3_U3175) );
  XNOR2_X1 U15375 ( .A(n12807), .B(n12806), .ZN(n12816) );
  NAND2_X1 U15376 ( .A1(n12834), .A2(n13336), .ZN(n12809) );
  OAI211_X1 U15377 ( .C1(n12810), .C2(n12836), .A(n12809), .B(n12808), .ZN(
        n12813) );
  NOR2_X1 U15378 ( .A1(n12811), .A2(n12842), .ZN(n12812) );
  AOI211_X1 U15379 ( .C1(n13339), .C2(n12839), .A(n12813), .B(n12812), .ZN(
        n12814) );
  OAI21_X1 U15380 ( .B1(n12816), .B2(n12815), .A(n12814), .ZN(P3_U3178) );
  OAI21_X1 U15381 ( .B1(n12819), .B2(n12818), .A(n12817), .ZN(n12820) );
  NAND2_X1 U15382 ( .A1(n12820), .A2(n12832), .ZN(n12827) );
  OAI22_X1 U15383 ( .A1(n13249), .A2(n12836), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12821), .ZN(n12825) );
  NOR2_X1 U15384 ( .A1(n12823), .A2(n12822), .ZN(n12824) );
  AOI211_X1 U15385 ( .C1(n13225), .C2(n12839), .A(n12825), .B(n12824), .ZN(
        n12826) );
  OAI211_X1 U15386 ( .C1(n12828), .C2(n12842), .A(n12827), .B(n12826), .ZN(
        P3_U3180) );
  OAI21_X1 U15387 ( .B1(n12831), .B2(n12830), .A(n12829), .ZN(n12833) );
  NAND2_X1 U15388 ( .A1(n12833), .A2(n12832), .ZN(n12841) );
  NAND2_X1 U15389 ( .A1(n12834), .A2(n13373), .ZN(n12835) );
  NAND2_X1 U15390 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n13103)
         );
  OAI211_X1 U15391 ( .C1(n12837), .C2(n12836), .A(n12835), .B(n13103), .ZN(
        n12838) );
  AOI21_X1 U15392 ( .B1(n13375), .B2(n12839), .A(n12838), .ZN(n12840) );
  OAI211_X1 U15393 ( .C1(n12843), .C2(n12842), .A(n12841), .B(n12840), .ZN(
        P3_U3181) );
  INV_X1 U15394 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n12846) );
  AOI22_X1 U15395 ( .A1(n9466), .A2(P3_REG2_REG_30__SCAN_IN), .B1(n12855), 
        .B2(P3_REG1_REG_30__SCAN_IN), .ZN(n12845) );
  OAI211_X1 U15396 ( .C1(n12847), .C2(n12846), .A(n12861), .B(n12845), .ZN(
        n13033) );
  XNOR2_X1 U15397 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12851) );
  XNOR2_X1 U15398 ( .A(n12852), .B(n12851), .ZN(n13602) );
  NAND2_X1 U15399 ( .A1(n13602), .A2(n7262), .ZN(n12854) );
  NAND2_X1 U15400 ( .A1(n12863), .A2(SI_31_), .ZN(n12853) );
  NAND2_X1 U15401 ( .A1(n9176), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12857) );
  NAND2_X1 U15402 ( .A1(n12855), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12856) );
  OAI211_X1 U15403 ( .C1(n12858), .C2(n13188), .A(n12857), .B(n12856), .ZN(
        n12859) );
  INV_X1 U15404 ( .A(n12859), .ZN(n12860) );
  OR2_X1 U15405 ( .A1(n13183), .A2(n13185), .ZN(n13019) );
  OAI21_X1 U15406 ( .B1(n13507), .B2(n13033), .A(n13019), .ZN(n12872) );
  NAND2_X1 U15407 ( .A1(n12862), .A2(n7262), .ZN(n12865) );
  NAND2_X1 U15408 ( .A1(n12863), .A2(SI_29_), .ZN(n12864) );
  NOR2_X1 U15409 ( .A1(n12872), .A2(n12873), .ZN(n13020) );
  INV_X1 U15410 ( .A(n13020), .ZN(n12870) );
  INV_X1 U15411 ( .A(n13185), .ZN(n13032) );
  NAND2_X1 U15412 ( .A1(n13013), .A2(n13010), .ZN(n13017) );
  OAI21_X1 U15413 ( .B1(n12867), .B2(n13017), .A(n12866), .ZN(n13191) );
  INV_X1 U15414 ( .A(n13507), .ZN(n12869) );
  INV_X1 U15415 ( .A(n13033), .ZN(n13203) );
  OAI22_X1 U15416 ( .A1(n12869), .A2(n13203), .B1(n13504), .B2(n13032), .ZN(
        n13018) );
  INV_X1 U15417 ( .A(n13018), .ZN(n12893) );
  XNOR2_X1 U15418 ( .A(n12871), .B(n12895), .ZN(n13026) );
  INV_X1 U15419 ( .A(n12872), .ZN(n12892) );
  INV_X1 U15420 ( .A(n12873), .ZN(n12874) );
  NAND2_X1 U15421 ( .A1(n12992), .A2(n12995), .ZN(n13273) );
  INV_X1 U15422 ( .A(n13307), .ZN(n13300) );
  NAND2_X1 U15423 ( .A1(n12875), .A2(n13367), .ZN(n12955) );
  NOR2_X1 U15424 ( .A1(n12961), .A2(n12966), .ZN(n13370) );
  NAND2_X1 U15425 ( .A1(n12877), .A2(n12876), .ZN(n12880) );
  NAND4_X1 U15426 ( .A1(n12882), .A2(n12930), .A3(n12881), .A4(n12916), .ZN(
        n12885) );
  INV_X1 U15427 ( .A(n12935), .ZN(n12883) );
  NOR4_X1 U15428 ( .A1(n12885), .A2(n12884), .A3(n12941), .A4(n12883), .ZN(
        n12886) );
  NAND4_X1 U15429 ( .A1(n13002), .A2(n12888), .A3(n12887), .A4(n13251), .ZN(
        n12889) );
  NOR4_X1 U15430 ( .A1(n13194), .A2(n12890), .A3(n13224), .A4(n12889), .ZN(
        n12891) );
  NAND4_X1 U15431 ( .A1(n12893), .A2(n12892), .A3(n13200), .A4(n12891), .ZN(
        n12894) );
  INV_X1 U15432 ( .A(n12896), .ZN(n13580) );
  MUX2_X1 U15433 ( .A(n13381), .B(n13580), .S(n13011), .Z(n12956) );
  AOI21_X1 U15434 ( .B1(n9778), .B2(n12899), .A(n12902), .ZN(n12898) );
  OAI22_X1 U15435 ( .A1(n12898), .A2(n13006), .B1(n9778), .B2(n12897), .ZN(
        n12901) );
  AOI21_X1 U15436 ( .B1(n12904), .B2(n12903), .A(n13006), .ZN(n12907) );
  OAI211_X1 U15437 ( .C1(n12908), .C2(n12907), .A(n12912), .B(n12910), .ZN(
        n12917) );
  NAND2_X1 U15438 ( .A1(n12910), .A2(n12909), .ZN(n12911) );
  AOI22_X1 U15439 ( .A1(n12912), .A2(n12911), .B1(n13040), .B2(n15885), .ZN(
        n12914) );
  MUX2_X1 U15440 ( .A(n12914), .B(n12913), .S(n13011), .Z(n12915) );
  AND3_X1 U15441 ( .A1(n12917), .A2(n12916), .A3(n12915), .ZN(n12926) );
  NAND2_X1 U15442 ( .A1(n12918), .A2(n13039), .ZN(n12921) );
  NAND2_X1 U15443 ( .A1(n12919), .A2(n13006), .ZN(n12920) );
  MUX2_X1 U15444 ( .A(n12921), .B(n12920), .S(n15892), .Z(n12925) );
  NAND2_X1 U15445 ( .A1(n13037), .A2(n6956), .ZN(n12927) );
  MUX2_X1 U15446 ( .A(n12928), .B(n12927), .S(n13011), .Z(n12929) );
  MUX2_X1 U15447 ( .A(n12933), .B(n12932), .S(n13011), .Z(n12934) );
  INV_X1 U15448 ( .A(n12936), .ZN(n12939) );
  INV_X1 U15449 ( .A(n12937), .ZN(n12938) );
  MUX2_X1 U15450 ( .A(n12939), .B(n12938), .S(n13011), .Z(n12940) );
  NOR2_X1 U15451 ( .A1(n12941), .A2(n12940), .ZN(n12947) );
  INV_X1 U15452 ( .A(n12942), .ZN(n12945) );
  INV_X1 U15453 ( .A(n12943), .ZN(n12944) );
  MUX2_X1 U15454 ( .A(n12945), .B(n12944), .S(n13011), .Z(n12946) );
  OAI21_X1 U15455 ( .B1(n12949), .B2(n12948), .A(n13011), .ZN(n12950) );
  NAND2_X1 U15456 ( .A1(n12954), .A2(n13421), .ZN(n12952) );
  OAI21_X1 U15457 ( .B1(n13402), .B2(n13590), .A(n12952), .ZN(n12951) );
  MUX2_X1 U15458 ( .A(n12959), .B(n12958), .S(n13011), .Z(n12960) );
  OAI21_X1 U15459 ( .B1(n12962), .B2(n12961), .A(n13011), .ZN(n12964) );
  AOI21_X1 U15460 ( .B1(n12965), .B2(n12964), .A(n12963), .ZN(n12971) );
  INV_X1 U15461 ( .A(n12966), .ZN(n12967) );
  AOI21_X1 U15462 ( .B1(n12968), .B2(n12967), .A(n13011), .ZN(n12970) );
  OAI22_X1 U15463 ( .A1(n12971), .A2(n12970), .B1(n13011), .B2(n12969), .ZN(
        n12973) );
  NAND3_X1 U15464 ( .A1(n13299), .A2(n13006), .A3(n13316), .ZN(n12975) );
  AOI22_X1 U15465 ( .A1(n12973), .A2(n13348), .B1(n12972), .B2(n12975), .ZN(
        n12980) );
  INV_X1 U15466 ( .A(n12976), .ZN(n13315) );
  NOR3_X1 U15467 ( .A1(n12974), .A2(n13006), .A3(n13315), .ZN(n12979) );
  AOI21_X1 U15468 ( .B1(n12977), .B2(n12976), .A(n12975), .ZN(n12978) );
  MUX2_X1 U15469 ( .A(n12981), .B(n13299), .S(n13011), .Z(n12982) );
  INV_X1 U15470 ( .A(n12983), .ZN(n12986) );
  INV_X1 U15471 ( .A(n12984), .ZN(n12985) );
  MUX2_X1 U15472 ( .A(n12986), .B(n12985), .S(n13011), .Z(n12987) );
  NOR2_X1 U15473 ( .A1(n13286), .A2(n12987), .ZN(n12991) );
  MUX2_X1 U15474 ( .A(n12989), .B(n12988), .S(n13011), .Z(n12990) );
  INV_X1 U15475 ( .A(n12992), .ZN(n12993) );
  NAND2_X1 U15476 ( .A1(n12994), .A2(n12993), .ZN(n12996) );
  MUX2_X1 U15477 ( .A(n12996), .B(n12995), .S(n13011), .Z(n12997) );
  XNOR2_X1 U15478 ( .A(n12999), .B(n13011), .ZN(n13000) );
  OAI21_X1 U15479 ( .B1(n13245), .B2(n7925), .A(n13000), .ZN(n13001) );
  NAND3_X1 U15480 ( .A1(n13009), .A2(n13215), .A3(n13004), .ZN(n13007) );
  NAND3_X1 U15481 ( .A1(n13007), .A2(n13006), .A3(n13005), .ZN(n13016) );
  NOR2_X1 U15482 ( .A1(n13027), .A2(n9503), .ZN(n13030) );
  OAI21_X1 U15483 ( .B1(n13031), .B2(n13028), .A(P3_B_REG_SCAN_IN), .ZN(n13029) );
  OAI22_X1 U15484 ( .A1(n6606), .A2(n13031), .B1(n13030), .B2(n13029), .ZN(
        P3_U3296) );
  MUX2_X1 U15485 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n13032), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U15486 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n13033), .S(P3_U3897), .Z(
        P3_U3521) );
  INV_X1 U15487 ( .A(n13201), .ZN(n13195) );
  MUX2_X1 U15488 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n13195), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15489 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n13217), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15490 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n13234), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U15491 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n13218), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U15492 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n13289), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15493 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n6797), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U15494 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13288), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15495 ( .A(n13336), .B(P3_DATAO_REG_19__SCAN_IN), .S(n13043), .Z(
        P3_U3510) );
  MUX2_X1 U15496 ( .A(n13349), .B(P3_DATAO_REG_18__SCAN_IN), .S(n13043), .Z(
        P3_U3509) );
  MUX2_X1 U15497 ( .A(n13358), .B(P3_DATAO_REG_17__SCAN_IN), .S(n13043), .Z(
        P3_U3508) );
  MUX2_X1 U15498 ( .A(n13373), .B(P3_DATAO_REG_16__SCAN_IN), .S(n13043), .Z(
        P3_U3507) );
  MUX2_X1 U15499 ( .A(n13382), .B(P3_DATAO_REG_15__SCAN_IN), .S(n13043), .Z(
        P3_U3506) );
  MUX2_X1 U15500 ( .A(n13392), .B(P3_DATAO_REG_14__SCAN_IN), .S(n13043), .Z(
        P3_U3505) );
  MUX2_X1 U15501 ( .A(n13381), .B(P3_DATAO_REG_13__SCAN_IN), .S(n13043), .Z(
        P3_U3504) );
  MUX2_X1 U15502 ( .A(n13421), .B(P3_DATAO_REG_12__SCAN_IN), .S(n13043), .Z(
        P3_U3503) );
  MUX2_X1 U15503 ( .A(n13034), .B(P3_DATAO_REG_11__SCAN_IN), .S(n13043), .Z(
        P3_U3502) );
  MUX2_X1 U15504 ( .A(n13423), .B(P3_DATAO_REG_10__SCAN_IN), .S(n13043), .Z(
        P3_U3501) );
  MUX2_X1 U15505 ( .A(n13035), .B(P3_DATAO_REG_9__SCAN_IN), .S(n13043), .Z(
        P3_U3500) );
  MUX2_X1 U15506 ( .A(n13036), .B(P3_DATAO_REG_8__SCAN_IN), .S(n13043), .Z(
        P3_U3499) );
  MUX2_X1 U15507 ( .A(n13037), .B(P3_DATAO_REG_7__SCAN_IN), .S(n13043), .Z(
        P3_U3498) );
  MUX2_X1 U15508 ( .A(n13038), .B(P3_DATAO_REG_6__SCAN_IN), .S(n13043), .Z(
        P3_U3497) );
  MUX2_X1 U15509 ( .A(n13039), .B(P3_DATAO_REG_5__SCAN_IN), .S(n13043), .Z(
        P3_U3496) );
  MUX2_X1 U15510 ( .A(n13040), .B(P3_DATAO_REG_4__SCAN_IN), .S(n13043), .Z(
        P3_U3495) );
  MUX2_X1 U15511 ( .A(n13041), .B(P3_DATAO_REG_3__SCAN_IN), .S(n13043), .Z(
        P3_U3494) );
  MUX2_X1 U15512 ( .A(n13042), .B(P3_DATAO_REG_1__SCAN_IN), .S(n13043), .Z(
        P3_U3492) );
  MUX2_X1 U15513 ( .A(n13044), .B(P3_DATAO_REG_0__SCAN_IN), .S(n13043), .Z(
        P3_U3491) );
  NOR3_X1 U15514 ( .A1(n13047), .A2(n13046), .A3(n13045), .ZN(n13048) );
  OAI21_X1 U15515 ( .B1(n6696), .B2(n13048), .A(n13097), .ZN(n13065) );
  OAI21_X1 U15516 ( .B1(n13144), .B2(n13050), .A(n13049), .ZN(n13051) );
  AOI21_X1 U15517 ( .B1(n13052), .B2(n13152), .A(n13051), .ZN(n13064) );
  OAI21_X1 U15518 ( .B1(n13055), .B2(n13054), .A(n13053), .ZN(n13056) );
  NAND2_X1 U15519 ( .A1(n13056), .A2(n13180), .ZN(n13063) );
  INV_X1 U15520 ( .A(n13071), .ZN(n13061) );
  OAI21_X1 U15521 ( .B1(n13059), .B2(n13058), .A(n13057), .ZN(n13060) );
  NAND3_X1 U15522 ( .A1(n13061), .A2(n13173), .A3(n13060), .ZN(n13062) );
  NAND4_X1 U15523 ( .A1(n13065), .A2(n13064), .A3(n13063), .A4(n13062), .ZN(
        P3_U3194) );
  AOI21_X1 U15524 ( .B1(n13394), .B2(n13066), .A(n13086), .ZN(n13079) );
  OAI21_X1 U15525 ( .B1(n13144), .B2(n13068), .A(n13067), .ZN(n13074) );
  OAI21_X1 U15526 ( .B1(n13071), .B2(n13070), .A(n13069), .ZN(n13072) );
  AOI21_X1 U15527 ( .B1(n7406), .B2(n13072), .A(n13146), .ZN(n13073) );
  AOI211_X1 U15528 ( .C1(n13152), .C2(n7518), .A(n13074), .B(n13073), .ZN(
        n13078) );
  XOR2_X1 U15529 ( .A(P3_REG1_REG_13__SCAN_IN), .B(n13075), .Z(n13076) );
  NAND2_X1 U15530 ( .A1(n13076), .A2(n13180), .ZN(n13077) );
  OAI211_X1 U15531 ( .C1(n13079), .C2(n13182), .A(n13078), .B(n13077), .ZN(
        P3_U3195) );
  XNOR2_X1 U15532 ( .A(n13081), .B(n13080), .ZN(n13100) );
  NAND2_X1 U15533 ( .A1(n13083), .A2(n13082), .ZN(n13085) );
  OAI21_X1 U15534 ( .B1(n13086), .B2(n13085), .A(n13084), .ZN(n13098) );
  OAI21_X1 U15535 ( .B1(n13089), .B2(n13088), .A(n13087), .ZN(n13091) );
  NAND3_X1 U15536 ( .A1(n13091), .A2(n13173), .A3(n13090), .ZN(n13094) );
  AOI21_X1 U15537 ( .B1(n15849), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n13092), 
        .ZN(n13093) );
  OAI211_X1 U15538 ( .C1(n13171), .C2(n13095), .A(n13094), .B(n13093), .ZN(
        n13096) );
  AOI21_X1 U15539 ( .B1(n13098), .B2(n13097), .A(n13096), .ZN(n13099) );
  OAI21_X1 U15540 ( .B1(n13101), .B2(n13100), .A(n13099), .ZN(P3_U3196) );
  AOI21_X1 U15541 ( .B1(n13374), .B2(n13102), .A(n13126), .ZN(n13117) );
  OAI21_X1 U15542 ( .B1(n13144), .B2(n13104), .A(n13103), .ZN(n13110) );
  AOI21_X1 U15543 ( .B1(n13107), .B2(n13106), .A(n13105), .ZN(n13108) );
  NOR2_X1 U15544 ( .A1(n13108), .A2(n13146), .ZN(n13109) );
  AOI211_X1 U15545 ( .C1(n13152), .C2(n13111), .A(n13110), .B(n13109), .ZN(
        n13116) );
  OAI21_X1 U15546 ( .B1(n13113), .B2(P3_REG1_REG_15__SCAN_IN), .A(n13112), 
        .ZN(n13114) );
  NAND2_X1 U15547 ( .A1(n13114), .A2(n13180), .ZN(n13115) );
  OAI211_X1 U15548 ( .C1(n13117), .C2(n13182), .A(n13116), .B(n13115), .ZN(
        P3_U3197) );
  NAND2_X1 U15549 ( .A1(n6720), .A2(n13118), .ZN(n13119) );
  XNOR2_X1 U15550 ( .A(n13120), .B(n13119), .ZN(n13131) );
  NAND2_X1 U15551 ( .A1(n15849), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n13121) );
  OAI211_X1 U15552 ( .C1(n13171), .C2(n13123), .A(n13122), .B(n13121), .ZN(
        n13130) );
  OR3_X1 U15553 ( .A1(n13126), .A2(n13125), .A3(n13124), .ZN(n13127) );
  AOI21_X1 U15554 ( .B1(n13128), .B2(n13127), .A(n13182), .ZN(n13129) );
  AOI211_X1 U15555 ( .C1(n13173), .C2(n13131), .A(n13130), .B(n13129), .ZN(
        n13139) );
  INV_X1 U15556 ( .A(n13132), .ZN(n13137) );
  NOR3_X1 U15557 ( .A1(n13135), .A2(n13134), .A3(n13133), .ZN(n13136) );
  OAI21_X1 U15558 ( .B1(n13137), .B2(n13136), .A(n13180), .ZN(n13138) );
  NAND2_X1 U15559 ( .A1(n13139), .A2(n13138), .ZN(P3_U3198) );
  AOI21_X1 U15560 ( .B1(n13351), .B2(n13141), .A(n13140), .ZN(n13157) );
  OAI21_X1 U15561 ( .B1(n13144), .B2(n13143), .A(n13142), .ZN(n13150) );
  AOI211_X1 U15562 ( .C1(n13148), .C2(n13147), .A(n13146), .B(n13145), .ZN(
        n13149) );
  AOI211_X1 U15563 ( .C1(n13152), .C2(n13151), .A(n13150), .B(n13149), .ZN(
        n13156) );
  XOR2_X1 U15564 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n13153), .Z(n13154) );
  NAND2_X1 U15565 ( .A1(n13154), .A2(n13180), .ZN(n13155) );
  OAI211_X1 U15566 ( .C1(n13157), .C2(n13182), .A(n13156), .B(n13155), .ZN(
        P3_U3199) );
  INV_X1 U15567 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13326) );
  XNOR2_X1 U15568 ( .A(n13170), .B(n13326), .ZN(n13165) );
  NAND2_X1 U15569 ( .A1(n13161), .A2(n13160), .ZN(n13162) );
  NAND2_X1 U15570 ( .A1(n13163), .A2(n13162), .ZN(n13167) );
  XNOR2_X1 U15571 ( .A(n13170), .B(n13463), .ZN(n13178) );
  MUX2_X1 U15572 ( .A(n13178), .B(n13165), .S(n13164), .Z(n13166) );
  XNOR2_X1 U15573 ( .A(n13167), .B(n13166), .ZN(n13174) );
  NAND2_X1 U15574 ( .A1(n15849), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n13168) );
  OAI211_X1 U15575 ( .C1(n13171), .C2(n13170), .A(n13169), .B(n13168), .ZN(
        n13172) );
  AOI21_X1 U15576 ( .B1(n13174), .B2(n13173), .A(n13172), .ZN(n13181) );
  NAND2_X1 U15577 ( .A1(n13183), .A2(n13428), .ZN(n13187) );
  INV_X1 U15578 ( .A(P3_B_REG_SCAN_IN), .ZN(n13184) );
  OAI21_X1 U15579 ( .B1(n9503), .B2(n13184), .A(n13420), .ZN(n13202) );
  NOR2_X1 U15580 ( .A1(n13185), .A2(n13202), .ZN(n13502) );
  NOR2_X1 U15581 ( .A1(n13186), .A2(n15855), .ZN(n13205) );
  AOI21_X1 U15582 ( .B1(n13502), .B2(n15870), .A(n13205), .ZN(n13190) );
  OAI211_X1 U15583 ( .C1(n15870), .C2(n13188), .A(n13187), .B(n13190), .ZN(
        P3_U3202) );
  NAND2_X1 U15584 ( .A1(n15873), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n13189) );
  OAI211_X1 U15585 ( .C1(n13507), .C2(n13266), .A(n13190), .B(n13189), .ZN(
        P3_U3203) );
  XNOR2_X1 U15586 ( .A(n13191), .B(n13200), .ZN(n13513) );
  NAND2_X1 U15587 ( .A1(n13194), .A2(n13192), .ZN(n13198) );
  NAND3_X1 U15588 ( .A1(n13194), .A2(n13193), .A3(n13192), .ZN(n13197) );
  OAI22_X1 U15589 ( .A1(n13203), .A2(n13202), .B1(n13201), .B2(n15861), .ZN(
        n13204) );
  AOI21_X1 U15590 ( .B1(n13511), .B2(n13428), .A(n13205), .ZN(n13206) );
  NAND2_X1 U15591 ( .A1(n13207), .A2(n13428), .ZN(n13210) );
  AOI22_X1 U15592 ( .A1(n13208), .A2(n13427), .B1(n15873), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13209) );
  NAND2_X1 U15593 ( .A1(n13210), .A2(n13209), .ZN(n13211) );
  AOI21_X1 U15594 ( .B1(n10679), .B2(n13212), .A(n13211), .ZN(n13213) );
  OAI21_X1 U15595 ( .B1(n13214), .B2(n15873), .A(n13213), .ZN(P3_U3206) );
  XNOR2_X1 U15596 ( .A(n13216), .B(n13215), .ZN(n13222) );
  NAND2_X1 U15597 ( .A1(n13218), .A2(n13422), .ZN(n13219) );
  XNOR2_X1 U15598 ( .A(n13223), .B(n13224), .ZN(n13439) );
  NAND2_X1 U15599 ( .A1(n13438), .A2(n13428), .ZN(n13227) );
  AOI22_X1 U15600 ( .A1(n13225), .A2(n13427), .B1(n15873), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13226) );
  NAND2_X1 U15601 ( .A1(n13227), .A2(n13226), .ZN(n13228) );
  AOI21_X1 U15602 ( .B1(n13439), .B2(n13268), .A(n13228), .ZN(n13229) );
  OAI21_X1 U15603 ( .B1(n13440), .B2(n15873), .A(n13229), .ZN(P3_U3207) );
  XNOR2_X1 U15604 ( .A(n13232), .B(n13230), .ZN(n13445) );
  OAI211_X1 U15605 ( .C1(n13233), .C2(n13232), .A(n13231), .B(n15864), .ZN(
        n13236) );
  NAND2_X1 U15606 ( .A1(n13234), .A2(n13420), .ZN(n13235) );
  OAI211_X1 U15607 ( .C1(n13237), .C2(n15861), .A(n13236), .B(n13235), .ZN(
        n13442) );
  AOI22_X1 U15608 ( .A1(n13238), .A2(n13427), .B1(n15873), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n13239) );
  OAI21_X1 U15609 ( .B1(n13240), .B2(n13266), .A(n13239), .ZN(n13241) );
  AOI21_X1 U15610 ( .B1(n13442), .B2(n15870), .A(n13241), .ZN(n13242) );
  OAI21_X1 U15611 ( .B1(n13243), .B2(n13445), .A(n13242), .ZN(P3_U3208) );
  OAI211_X1 U15612 ( .C1(n13246), .C2(n13245), .A(n13244), .B(n15864), .ZN(
        n13248) );
  NAND2_X1 U15613 ( .A1(n13274), .A2(n13422), .ZN(n13247) );
  OAI211_X1 U15614 ( .C1(n13249), .C2(n15859), .A(n13248), .B(n13247), .ZN(
        n13446) );
  INV_X1 U15615 ( .A(n13446), .ZN(n13256) );
  OAI21_X1 U15616 ( .B1(n6620), .B2(n13251), .A(n13250), .ZN(n13447) );
  AOI22_X1 U15617 ( .A1(n13252), .A2(n13427), .B1(n15873), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n13253) );
  OAI21_X1 U15618 ( .B1(n13519), .B2(n13266), .A(n13253), .ZN(n13254) );
  AOI21_X1 U15619 ( .B1(n13447), .B2(n13411), .A(n13254), .ZN(n13255) );
  OAI21_X1 U15620 ( .B1(n13256), .B2(n15873), .A(n13255), .ZN(P3_U3209) );
  OAI211_X1 U15621 ( .C1(n13258), .C2(n13263), .A(n13257), .B(n15864), .ZN(
        n13261) );
  AOI22_X1 U15622 ( .A1(n13259), .A2(n13420), .B1(n13422), .B2(n13289), .ZN(
        n13260) );
  NAND2_X1 U15623 ( .A1(n13261), .A2(n13260), .ZN(n13450) );
  INV_X1 U15624 ( .A(n13450), .ZN(n13270) );
  XNOR2_X1 U15625 ( .A(n13262), .B(n13263), .ZN(n13451) );
  AOI22_X1 U15626 ( .A1(n13264), .A2(n13427), .B1(n15873), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n13265) );
  OAI21_X1 U15627 ( .B1(n13523), .B2(n13266), .A(n13265), .ZN(n13267) );
  AOI21_X1 U15628 ( .B1(n13451), .B2(n13268), .A(n13267), .ZN(n13269) );
  OAI21_X1 U15629 ( .B1(n13270), .B2(n15873), .A(n13269), .ZN(P3_U3210) );
  XOR2_X1 U15630 ( .A(n13271), .B(n13273), .Z(n13529) );
  INV_X1 U15631 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n13276) );
  XNOR2_X1 U15632 ( .A(n13272), .B(n13273), .ZN(n13275) );
  AOI222_X1 U15633 ( .A1(n15864), .A2(n13275), .B1(n13274), .B2(n13420), .C1(
        n6797), .C2(n13422), .ZN(n13524) );
  MUX2_X1 U15634 ( .A(n13276), .B(n13524), .S(n15870), .Z(n13279) );
  AOI22_X1 U15635 ( .A1(n13526), .A2(n13428), .B1(n13427), .B2(n13277), .ZN(
        n13278) );
  OAI211_X1 U15636 ( .C1(n13529), .C2(n13431), .A(n13279), .B(n13278), .ZN(
        P3_U3211) );
  XOR2_X1 U15637 ( .A(n13280), .B(n13286), .Z(n13535) );
  INV_X1 U15638 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n13291) );
  OAI21_X1 U15639 ( .B1(n13331), .B2(n13282), .A(n13281), .ZN(n13284) );
  AND2_X1 U15640 ( .A1(n13284), .A2(n13283), .ZN(n13287) );
  OAI21_X1 U15641 ( .B1(n13287), .B2(n13286), .A(n13285), .ZN(n13290) );
  AOI222_X1 U15642 ( .A1(n15864), .A2(n13290), .B1(n13289), .B2(n13420), .C1(
        n13288), .C2(n13422), .ZN(n13530) );
  MUX2_X1 U15643 ( .A(n13291), .B(n13530), .S(n15870), .Z(n13294) );
  AOI22_X1 U15644 ( .A1(n13532), .A2(n13428), .B1(n13427), .B2(n13292), .ZN(
        n13293) );
  OAI211_X1 U15645 ( .C1(n13535), .C2(n13431), .A(n13294), .B(n13293), .ZN(
        P3_U3212) );
  INV_X1 U15646 ( .A(n13295), .ZN(n13344) );
  INV_X1 U15647 ( .A(n13296), .ZN(n13298) );
  OAI21_X1 U15648 ( .B1(n13344), .B2(n13298), .A(n13297), .ZN(n13301) );
  NAND3_X1 U15649 ( .A1(n13301), .A2(n13300), .A3(n13299), .ZN(n13303) );
  NAND2_X1 U15650 ( .A1(n13303), .A2(n13302), .ZN(n13541) );
  INV_X1 U15651 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n13310) );
  INV_X1 U15652 ( .A(n13334), .ZN(n13304) );
  NOR2_X1 U15653 ( .A1(n13331), .A2(n13304), .ZN(n13332) );
  OR2_X1 U15654 ( .A1(n13332), .A2(n13305), .ZN(n13320) );
  NAND2_X1 U15655 ( .A1(n13320), .A2(n13306), .ZN(n13308) );
  XNOR2_X1 U15656 ( .A(n13308), .B(n13307), .ZN(n13309) );
  AOI222_X1 U15657 ( .A1(n13336), .A2(n13422), .B1(n6797), .B2(n13420), .C1(
        n15864), .C2(n13309), .ZN(n13536) );
  MUX2_X1 U15658 ( .A(n13310), .B(n13536), .S(n15870), .Z(n13313) );
  AOI22_X1 U15659 ( .A1(n13538), .A2(n13428), .B1(n13427), .B2(n13311), .ZN(
        n13312) );
  OAI211_X1 U15660 ( .C1(n13541), .C2(n13431), .A(n13313), .B(n13312), .ZN(
        P3_U3213) );
  NAND2_X1 U15661 ( .A1(n13295), .A2(n13348), .ZN(n13342) );
  NAND2_X1 U15662 ( .A1(n13342), .A2(n13314), .ZN(n13330) );
  AOI21_X1 U15663 ( .B1(n13330), .B2(n13316), .A(n13315), .ZN(n13317) );
  XNOR2_X1 U15664 ( .A(n13317), .B(n13318), .ZN(n13547) );
  OAI21_X1 U15665 ( .B1(n13332), .B2(n13319), .A(n13318), .ZN(n13321) );
  AND3_X1 U15666 ( .A1(n13321), .A2(n15864), .A3(n13320), .ZN(n13325) );
  OAI22_X1 U15667 ( .A1(n13323), .A2(n15859), .B1(n13322), .B2(n15861), .ZN(
        n13324) );
  NOR2_X1 U15668 ( .A1(n13325), .A2(n13324), .ZN(n13542) );
  MUX2_X1 U15669 ( .A(n13326), .B(n13542), .S(n15870), .Z(n13329) );
  AOI22_X1 U15670 ( .A1(n13544), .A2(n13428), .B1(n13427), .B2(n13327), .ZN(
        n13328) );
  OAI211_X1 U15671 ( .C1(n13547), .C2(n13431), .A(n13329), .B(n13328), .ZN(
        P3_U3214) );
  XNOR2_X1 U15672 ( .A(n13330), .B(n13334), .ZN(n13553) );
  INV_X1 U15673 ( .A(n13331), .ZN(n13335) );
  INV_X1 U15674 ( .A(n13332), .ZN(n13333) );
  OAI21_X1 U15675 ( .B1(n13335), .B2(n13334), .A(n13333), .ZN(n13337) );
  AOI222_X1 U15676 ( .A1(n15864), .A2(n13337), .B1(n13336), .B2(n13420), .C1(
        n13358), .C2(n13422), .ZN(n13548) );
  MUX2_X1 U15677 ( .A(n13338), .B(n13548), .S(n15870), .Z(n13341) );
  AOI22_X1 U15678 ( .A1(n13550), .A2(n13428), .B1(n13427), .B2(n13339), .ZN(
        n13340) );
  OAI211_X1 U15679 ( .C1(n13553), .C2(n13431), .A(n13341), .B(n13340), .ZN(
        P3_U3215) );
  INV_X1 U15680 ( .A(n13348), .ZN(n13345) );
  INV_X1 U15681 ( .A(n13342), .ZN(n13343) );
  AOI21_X1 U15682 ( .B1(n13345), .B2(n13344), .A(n13343), .ZN(n13559) );
  XOR2_X1 U15683 ( .A(n13348), .B(n13347), .Z(n13350) );
  AOI222_X1 U15684 ( .A1(n15864), .A2(n13350), .B1(n13349), .B2(n13420), .C1(
        n13373), .C2(n13422), .ZN(n13554) );
  MUX2_X1 U15685 ( .A(n13351), .B(n13554), .S(n15870), .Z(n13354) );
  AOI22_X1 U15686 ( .A1(n13556), .A2(n13428), .B1(n13352), .B2(n13427), .ZN(
        n13353) );
  OAI211_X1 U15687 ( .C1(n13559), .C2(n13431), .A(n13354), .B(n13353), .ZN(
        P3_U3216) );
  XNOR2_X1 U15688 ( .A(n13355), .B(n13356), .ZN(n13565) );
  XNOR2_X1 U15689 ( .A(n13357), .B(n13356), .ZN(n13359) );
  AOI222_X1 U15690 ( .A1(n15864), .A2(n13359), .B1(n13358), .B2(n13420), .C1(
        n13382), .C2(n13422), .ZN(n13560) );
  MUX2_X1 U15691 ( .A(n13360), .B(n13560), .S(n15870), .Z(n13363) );
  AOI22_X1 U15692 ( .A1(n13562), .A2(n13428), .B1(n13427), .B2(n13361), .ZN(
        n13362) );
  OAI211_X1 U15693 ( .C1(n13565), .C2(n13431), .A(n13363), .B(n13362), .ZN(
        P3_U3217) );
  NOR2_X1 U15694 ( .A1(n13364), .A2(n13379), .ZN(n13378) );
  NOR2_X1 U15695 ( .A1(n13378), .A2(n13365), .ZN(n13366) );
  XNOR2_X1 U15696 ( .A(n13366), .B(n13370), .ZN(n13571) );
  NAND2_X1 U15697 ( .A1(n13390), .A2(n13391), .ZN(n13389) );
  NAND2_X1 U15698 ( .A1(n13389), .A2(n13367), .ZN(n13380) );
  OAI21_X1 U15699 ( .B1(n13380), .B2(n13369), .A(n13368), .ZN(n13371) );
  XNOR2_X1 U15700 ( .A(n13371), .B(n13370), .ZN(n13372) );
  AOI222_X1 U15701 ( .A1(n13392), .A2(n13422), .B1(n13373), .B2(n13420), .C1(
        n15864), .C2(n13372), .ZN(n13566) );
  MUX2_X1 U15702 ( .A(n13374), .B(n13566), .S(n15870), .Z(n13377) );
  AOI22_X1 U15703 ( .A1(n13568), .A2(n13428), .B1(n13427), .B2(n13375), .ZN(
        n13376) );
  OAI211_X1 U15704 ( .C1(n13571), .C2(n13431), .A(n13377), .B(n13376), .ZN(
        P3_U3218) );
  AOI21_X1 U15705 ( .B1(n13364), .B2(n13379), .A(n13378), .ZN(n13577) );
  XNOR2_X1 U15706 ( .A(n13380), .B(n13379), .ZN(n13383) );
  AOI222_X1 U15707 ( .A1(n15864), .A2(n13383), .B1(n13382), .B2(n13420), .C1(
        n13381), .C2(n13422), .ZN(n13572) );
  MUX2_X1 U15708 ( .A(n13384), .B(n13572), .S(n15870), .Z(n13387) );
  AOI22_X1 U15709 ( .A1(n13574), .A2(n13428), .B1(n13427), .B2(n13385), .ZN(
        n13386) );
  OAI211_X1 U15710 ( .C1(n13577), .C2(n13431), .A(n13387), .B(n13386), .ZN(
        P3_U3219) );
  XNOR2_X1 U15711 ( .A(n13388), .B(n13391), .ZN(n13583) );
  OAI21_X1 U15712 ( .B1(n13391), .B2(n13390), .A(n13389), .ZN(n13393) );
  AOI222_X1 U15713 ( .A1(n15864), .A2(n13393), .B1(n13392), .B2(n13420), .C1(
        n13421), .C2(n13422), .ZN(n13578) );
  MUX2_X1 U15714 ( .A(n13394), .B(n13578), .S(n15870), .Z(n13397) );
  AOI22_X1 U15715 ( .A1(n13580), .A2(n13428), .B1(n13427), .B2(n13395), .ZN(
        n13396) );
  OAI211_X1 U15716 ( .C1(n13583), .C2(n13431), .A(n13397), .B(n13396), .ZN(
        P3_U3220) );
  XOR2_X1 U15717 ( .A(n13399), .B(n13405), .Z(n13400) );
  OAI222_X1 U15718 ( .A1(n15859), .A2(n13403), .B1(n15861), .B2(n13402), .C1(
        n13401), .C2(n13400), .ZN(n13483) );
  INV_X1 U15719 ( .A(n13483), .ZN(n13414) );
  INV_X1 U15720 ( .A(n13405), .ZN(n13406) );
  XNOR2_X1 U15721 ( .A(n13404), .B(n13406), .ZN(n13587) );
  INV_X1 U15722 ( .A(n13587), .ZN(n13412) );
  NAND2_X1 U15723 ( .A1(n13484), .A2(n13428), .ZN(n13408) );
  NAND2_X1 U15724 ( .A1(n15873), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n13407) );
  OAI211_X1 U15725 ( .C1(n13409), .C2(n15855), .A(n13408), .B(n13407), .ZN(
        n13410) );
  AOI21_X1 U15726 ( .B1(n13412), .B2(n13411), .A(n13410), .ZN(n13413) );
  OAI21_X1 U15727 ( .B1(n13414), .B2(n15873), .A(n13413), .ZN(P3_U3221) );
  XNOR2_X1 U15728 ( .A(n13415), .B(n13416), .ZN(n13594) );
  XNOR2_X1 U15729 ( .A(n13417), .B(n13418), .ZN(n13419) );
  AOI222_X1 U15730 ( .A1(n13423), .A2(n13422), .B1(n13421), .B2(n13420), .C1(
        n15864), .C2(n13419), .ZN(n13588) );
  MUX2_X1 U15731 ( .A(n13424), .B(n13588), .S(n15870), .Z(n13430) );
  INV_X1 U15732 ( .A(n13425), .ZN(n13426) );
  AOI22_X1 U15733 ( .A1(n13428), .A2(n13590), .B1(n13427), .B2(n13426), .ZN(
        n13429) );
  OAI211_X1 U15734 ( .C1(n13594), .C2(n13431), .A(n13430), .B(n13429), .ZN(
        P3_U3222) );
  NAND2_X1 U15735 ( .A1(n13502), .A2(n15918), .ZN(n13433) );
  NAND2_X1 U15736 ( .A1(n10706), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13432) );
  OAI211_X1 U15737 ( .C1(n13504), .C2(n13496), .A(n13433), .B(n13432), .ZN(
        P3_U3490) );
  NAND2_X1 U15738 ( .A1(n10706), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n13434) );
  OAI211_X1 U15739 ( .C1(n13507), .C2(n13496), .A(n13434), .B(n13433), .ZN(
        P3_U3489) );
  INV_X1 U15740 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n13435) );
  NAND2_X1 U15741 ( .A1(n13511), .A2(n13488), .ZN(n13436) );
  OAI211_X1 U15742 ( .C1(n13513), .C2(n13491), .A(n13437), .B(n13436), .ZN(
        P3_U3488) );
  AOI22_X1 U15743 ( .A1(n13439), .A2(n15899), .B1(n13499), .B2(n13438), .ZN(
        n13441) );
  MUX2_X1 U15744 ( .A(P3_REG1_REG_26__SCAN_IN), .B(n13514), .S(n15918), .Z(
        P3_U3485) );
  AOI21_X1 U15745 ( .B1(n13499), .B2(n13443), .A(n13442), .ZN(n13444) );
  OAI21_X1 U15746 ( .B1(n13508), .B2(n13445), .A(n13444), .ZN(n13515) );
  MUX2_X1 U15747 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n13515), .S(n15918), .Z(
        P3_U3484) );
  INV_X1 U15748 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13448) );
  AOI21_X1 U15749 ( .B1(n15899), .B2(n13447), .A(n13446), .ZN(n13516) );
  MUX2_X1 U15750 ( .A(n13448), .B(n13516), .S(n15918), .Z(n13449) );
  OAI21_X1 U15751 ( .B1(n13519), .B2(n13496), .A(n13449), .ZN(P3_U3483) );
  INV_X1 U15752 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13452) );
  AOI21_X1 U15753 ( .B1(n15899), .B2(n13451), .A(n13450), .ZN(n13520) );
  MUX2_X1 U15754 ( .A(n13452), .B(n13520), .S(n15918), .Z(n13453) );
  OAI21_X1 U15755 ( .B1(n13523), .B2(n13496), .A(n13453), .ZN(P3_U3482) );
  INV_X1 U15756 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13454) );
  MUX2_X1 U15757 ( .A(n13454), .B(n13524), .S(n15918), .Z(n13456) );
  NAND2_X1 U15758 ( .A1(n13526), .A2(n13488), .ZN(n13455) );
  OAI211_X1 U15759 ( .C1(n13529), .C2(n13491), .A(n13456), .B(n13455), .ZN(
        P3_U3481) );
  INV_X1 U15760 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13457) );
  MUX2_X1 U15761 ( .A(n13457), .B(n13530), .S(n15918), .Z(n13459) );
  NAND2_X1 U15762 ( .A1(n13532), .A2(n13488), .ZN(n13458) );
  OAI211_X1 U15763 ( .C1(n13535), .C2(n13491), .A(n13459), .B(n13458), .ZN(
        P3_U3480) );
  MUX2_X1 U15764 ( .A(n13460), .B(n13536), .S(n15918), .Z(n13462) );
  NAND2_X1 U15765 ( .A1(n13538), .A2(n13488), .ZN(n13461) );
  OAI211_X1 U15766 ( .C1(n13491), .C2(n13541), .A(n13462), .B(n13461), .ZN(
        P3_U3479) );
  MUX2_X1 U15767 ( .A(n13463), .B(n13542), .S(n15918), .Z(n13465) );
  NAND2_X1 U15768 ( .A1(n13544), .A2(n13488), .ZN(n13464) );
  OAI211_X1 U15769 ( .C1(n13491), .C2(n13547), .A(n13465), .B(n13464), .ZN(
        P3_U3478) );
  MUX2_X1 U15770 ( .A(n7535), .B(n13548), .S(n15918), .Z(n13467) );
  NAND2_X1 U15771 ( .A1(n13550), .A2(n13488), .ZN(n13466) );
  OAI211_X1 U15772 ( .C1(n13491), .C2(n13553), .A(n13467), .B(n13466), .ZN(
        P3_U3477) );
  MUX2_X1 U15773 ( .A(n13468), .B(n13554), .S(n15918), .Z(n13470) );
  NAND2_X1 U15774 ( .A1(n13556), .A2(n13488), .ZN(n13469) );
  OAI211_X1 U15775 ( .C1(n13559), .C2(n13491), .A(n13470), .B(n13469), .ZN(
        P3_U3476) );
  MUX2_X1 U15776 ( .A(n13471), .B(n13560), .S(n15918), .Z(n13473) );
  NAND2_X1 U15777 ( .A1(n13562), .A2(n13488), .ZN(n13472) );
  OAI211_X1 U15778 ( .C1(n13491), .C2(n13565), .A(n13473), .B(n13472), .ZN(
        P3_U3475) );
  INV_X1 U15779 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13474) );
  MUX2_X1 U15780 ( .A(n13474), .B(n13566), .S(n15918), .Z(n13476) );
  NAND2_X1 U15781 ( .A1(n13568), .A2(n13488), .ZN(n13475) );
  OAI211_X1 U15782 ( .C1(n13491), .C2(n13571), .A(n13476), .B(n13475), .ZN(
        P3_U3474) );
  INV_X1 U15783 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13477) );
  MUX2_X1 U15784 ( .A(n13477), .B(n13572), .S(n15918), .Z(n13479) );
  NAND2_X1 U15785 ( .A1(n13574), .A2(n13488), .ZN(n13478) );
  OAI211_X1 U15786 ( .C1(n13577), .C2(n13491), .A(n13479), .B(n13478), .ZN(
        P3_U3473) );
  MUX2_X1 U15787 ( .A(n13480), .B(n13578), .S(n15918), .Z(n13482) );
  NAND2_X1 U15788 ( .A1(n13580), .A2(n13488), .ZN(n13481) );
  OAI211_X1 U15789 ( .C1(n13583), .C2(n13491), .A(n13482), .B(n13481), .ZN(
        P3_U3472) );
  AOI21_X1 U15790 ( .B1(n13484), .B2(n13499), .A(n13483), .ZN(n13584) );
  MUX2_X1 U15791 ( .A(n13485), .B(n13584), .S(n15918), .Z(n13486) );
  OAI21_X1 U15792 ( .B1(n13491), .B2(n13587), .A(n13486), .ZN(P3_U3471) );
  MUX2_X1 U15793 ( .A(n13487), .B(n13588), .S(n15918), .Z(n13490) );
  NAND2_X1 U15794 ( .A1(n13488), .A2(n13590), .ZN(n13489) );
  OAI211_X1 U15795 ( .C1(n13491), .C2(n13594), .A(n13490), .B(n13489), .ZN(
        P3_U3470) );
  AOI21_X1 U15796 ( .B1(n15879), .B2(n13493), .A(n13492), .ZN(n13595) );
  MUX2_X1 U15797 ( .A(n13494), .B(n13595), .S(n15918), .Z(n13495) );
  OAI21_X1 U15798 ( .B1(n13496), .B2(n13598), .A(n13495), .ZN(P3_U3469) );
  AOI21_X1 U15799 ( .B1(n13499), .B2(n13498), .A(n13497), .ZN(n13500) );
  OAI21_X1 U15800 ( .B1(n13508), .B2(n13501), .A(n13500), .ZN(n13600) );
  MUX2_X1 U15801 ( .A(P3_REG1_REG_8__SCAN_IN), .B(n13600), .S(n15918), .Z(
        P3_U3467) );
  NAND2_X1 U15802 ( .A1(n13502), .A2(n15905), .ZN(n13505) );
  NAND2_X1 U15803 ( .A1(n15906), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n13503) );
  OAI211_X1 U15804 ( .C1(n13504), .C2(n13599), .A(n13505), .B(n13503), .ZN(
        P3_U3458) );
  NAND2_X1 U15805 ( .A1(n15906), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n13506) );
  OAI211_X1 U15806 ( .C1(n13507), .C2(n13599), .A(n13506), .B(n13505), .ZN(
        P3_U3457) );
  NAND2_X1 U15807 ( .A1(n13511), .A2(n10701), .ZN(n13512) );
  MUX2_X1 U15808 ( .A(P3_REG0_REG_26__SCAN_IN), .B(n13514), .S(n15905), .Z(
        P3_U3453) );
  MUX2_X1 U15809 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n13515), .S(n15905), .Z(
        P3_U3452) );
  MUX2_X1 U15810 ( .A(n13517), .B(n13516), .S(n15905), .Z(n13518) );
  OAI21_X1 U15811 ( .B1(n13519), .B2(n13599), .A(n13518), .ZN(P3_U3451) );
  MUX2_X1 U15812 ( .A(n13521), .B(n13520), .S(n15905), .Z(n13522) );
  OAI21_X1 U15813 ( .B1(n13523), .B2(n13599), .A(n13522), .ZN(P3_U3450) );
  MUX2_X1 U15814 ( .A(n13525), .B(n13524), .S(n15905), .Z(n13528) );
  NAND2_X1 U15815 ( .A1(n13526), .A2(n10701), .ZN(n13527) );
  OAI211_X1 U15816 ( .C1(n13529), .C2(n13593), .A(n13528), .B(n13527), .ZN(
        P3_U3449) );
  MUX2_X1 U15817 ( .A(n13531), .B(n13530), .S(n15905), .Z(n13534) );
  NAND2_X1 U15818 ( .A1(n13532), .A2(n10701), .ZN(n13533) );
  OAI211_X1 U15819 ( .C1(n13535), .C2(n13593), .A(n13534), .B(n13533), .ZN(
        P3_U3448) );
  INV_X1 U15820 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13537) );
  MUX2_X1 U15821 ( .A(n13537), .B(n13536), .S(n15905), .Z(n13540) );
  NAND2_X1 U15822 ( .A1(n13538), .A2(n10701), .ZN(n13539) );
  OAI211_X1 U15823 ( .C1(n13541), .C2(n13593), .A(n13540), .B(n13539), .ZN(
        P3_U3447) );
  INV_X1 U15824 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13543) );
  MUX2_X1 U15825 ( .A(n13543), .B(n13542), .S(n15905), .Z(n13546) );
  NAND2_X1 U15826 ( .A1(n13544), .A2(n10701), .ZN(n13545) );
  OAI211_X1 U15827 ( .C1(n13547), .C2(n13593), .A(n13546), .B(n13545), .ZN(
        P3_U3446) );
  MUX2_X1 U15828 ( .A(n13549), .B(n13548), .S(n15905), .Z(n13552) );
  NAND2_X1 U15829 ( .A1(n13550), .A2(n10701), .ZN(n13551) );
  OAI211_X1 U15830 ( .C1(n13553), .C2(n13593), .A(n13552), .B(n13551), .ZN(
        P3_U3444) );
  INV_X1 U15831 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13555) );
  MUX2_X1 U15832 ( .A(n13555), .B(n13554), .S(n15905), .Z(n13558) );
  NAND2_X1 U15833 ( .A1(n13556), .A2(n10701), .ZN(n13557) );
  OAI211_X1 U15834 ( .C1(n13559), .C2(n13593), .A(n13558), .B(n13557), .ZN(
        P3_U3441) );
  MUX2_X1 U15835 ( .A(n13561), .B(n13560), .S(n15905), .Z(n13564) );
  NAND2_X1 U15836 ( .A1(n13562), .A2(n10701), .ZN(n13563) );
  OAI211_X1 U15837 ( .C1(n13565), .C2(n13593), .A(n13564), .B(n13563), .ZN(
        P3_U3438) );
  MUX2_X1 U15838 ( .A(n13567), .B(n13566), .S(n15905), .Z(n13570) );
  NAND2_X1 U15839 ( .A1(n13568), .A2(n10701), .ZN(n13569) );
  OAI211_X1 U15840 ( .C1(n13571), .C2(n13593), .A(n13570), .B(n13569), .ZN(
        P3_U3435) );
  MUX2_X1 U15841 ( .A(n13573), .B(n13572), .S(n15905), .Z(n13576) );
  NAND2_X1 U15842 ( .A1(n13574), .A2(n10701), .ZN(n13575) );
  OAI211_X1 U15843 ( .C1(n13577), .C2(n13593), .A(n13576), .B(n13575), .ZN(
        P3_U3432) );
  MUX2_X1 U15844 ( .A(n13579), .B(n13578), .S(n15905), .Z(n13582) );
  NAND2_X1 U15845 ( .A1(n13580), .A2(n10701), .ZN(n13581) );
  OAI211_X1 U15846 ( .C1(n13583), .C2(n13593), .A(n13582), .B(n13581), .ZN(
        P3_U3429) );
  MUX2_X1 U15847 ( .A(n13585), .B(n13584), .S(n15905), .Z(n13586) );
  OAI21_X1 U15848 ( .B1(n13587), .B2(n13593), .A(n13586), .ZN(P3_U3426) );
  MUX2_X1 U15849 ( .A(n13589), .B(n13588), .S(n15905), .Z(n13592) );
  NAND2_X1 U15850 ( .A1(n10701), .A2(n13590), .ZN(n13591) );
  OAI211_X1 U15851 ( .C1(n13594), .C2(n13593), .A(n13592), .B(n13591), .ZN(
        P3_U3423) );
  MUX2_X1 U15852 ( .A(n13596), .B(n13595), .S(n15905), .Z(n13597) );
  OAI21_X1 U15853 ( .B1(n13599), .B2(n13598), .A(n13597), .ZN(P3_U3420) );
  MUX2_X1 U15854 ( .A(P3_REG0_REG_8__SCAN_IN), .B(n13600), .S(n15905), .Z(
        P3_U3414) );
  MUX2_X1 U15855 ( .A(P3_D_REG_0__SCAN_IN), .B(n9777), .S(n13601), .Z(P3_U3376) );
  INV_X1 U15856 ( .A(n13602), .ZN(n13607) );
  NOR4_X1 U15857 ( .A1(n13603), .A2(P3_IR_REG_30__SCAN_IN), .A3(P3_U3151), 
        .A4(n9015), .ZN(n13604) );
  AOI21_X1 U15858 ( .B1(n13605), .B2(SI_31_), .A(n13604), .ZN(n13606) );
  OAI21_X1 U15859 ( .B1(n13607), .B2(n13611), .A(n13606), .ZN(P3_U3264) );
  INV_X1 U15860 ( .A(n13608), .ZN(n13610) );
  OAI222_X1 U15861 ( .A1(n13612), .A2(P3_U3151), .B1(n13611), .B2(n13610), 
        .C1(n13609), .C2(n13618), .ZN(P3_U3268) );
  INV_X1 U15862 ( .A(SI_26_), .ZN(n13615) );
  INV_X1 U15863 ( .A(n13613), .ZN(n13614) );
  OAI222_X1 U15864 ( .A1(n13616), .A2(P3_U3151), .B1(n13618), .B2(n13615), 
        .C1(n13622), .C2(n13614), .ZN(P3_U3269) );
  INV_X1 U15865 ( .A(n13617), .ZN(n13621) );
  INV_X1 U15866 ( .A(SI_25_), .ZN(n13619) );
  OAI222_X1 U15867 ( .A1(n13622), .A2(n13621), .B1(P3_U3151), .B2(n13620), 
        .C1(n13619), .C2(n13618), .ZN(P3_U3270) );
  INV_X1 U15868 ( .A(n13623), .ZN(n13627) );
  AOI21_X1 U15869 ( .B1(n13625), .B2(n13624), .A(n13796), .ZN(n13626) );
  INV_X1 U15870 ( .A(n14209), .ZN(n13629) );
  OAI22_X1 U15871 ( .A1(n13629), .A2(n13804), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13628), .ZN(n13630) );
  AOI21_X1 U15872 ( .B1(n13631), .B2(n13730), .A(n13630), .ZN(n13632) );
  AND2_X1 U15873 ( .A1(n13634), .A2(n13633), .ZN(n13636) );
  OAI21_X1 U15874 ( .B1(n13637), .B2(n13636), .A(n13635), .ZN(n13638) );
  NAND2_X1 U15875 ( .A1(n13638), .A2(n13798), .ZN(n13643) );
  NAND2_X1 U15876 ( .A1(n6510), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n15714) );
  INV_X1 U15877 ( .A(n15714), .ZN(n13641) );
  INV_X1 U15878 ( .A(n14415), .ZN(n13639) );
  OAI22_X1 U15879 ( .A1(n14412), .A2(n13803), .B1(n13804), .B2(n13639), .ZN(
        n13640) );
  AOI211_X1 U15880 ( .C1(n13770), .C2(n14448), .A(n13641), .B(n13640), .ZN(
        n13642) );
  OAI211_X1 U15881 ( .C1(n14418), .C2(n13733), .A(n13643), .B(n13642), .ZN(
        P2_U3187) );
  OR2_X1 U15882 ( .A1(n13747), .A2(n13644), .ZN(n13749) );
  NAND2_X1 U15883 ( .A1(n13749), .A2(n13645), .ZN(n13647) );
  XNOR2_X1 U15884 ( .A(n13647), .B(n13646), .ZN(n13650) );
  OAI22_X1 U15885 ( .A1(n13650), .A2(n13796), .B1(n13717), .B2(n13758), .ZN(
        n13648) );
  OAI21_X1 U15886 ( .B1(n13650), .B2(n13649), .A(n13648), .ZN(n13654) );
  AOI22_X1 U15887 ( .A1(n14263), .A2(n13770), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(n6510), .ZN(n13651) );
  OAI21_X1 U15888 ( .B1(n14261), .B2(n13804), .A(n13651), .ZN(n13652) );
  AOI21_X1 U15889 ( .B1(n10559), .B2(n13769), .A(n13652), .ZN(n13653) );
  OAI211_X1 U15890 ( .C1(n14273), .C2(n13733), .A(n13654), .B(n13653), .ZN(
        P2_U3188) );
  XNOR2_X1 U15891 ( .A(n13726), .B(n13655), .ZN(n13656) );
  XNOR2_X1 U15892 ( .A(n13725), .B(n13656), .ZN(n13660) );
  OAI22_X1 U15893 ( .A1(n13909), .A2(n14474), .B1(n10517), .B2(n14472), .ZN(
        n14321) );
  NAND2_X1 U15894 ( .A1(n14321), .A2(n13730), .ZN(n13657) );
  NAND2_X1 U15895 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n14177)
         );
  OAI211_X1 U15896 ( .C1(n13804), .C2(n14326), .A(n13657), .B(n14177), .ZN(
        n13658) );
  AOI21_X1 U15897 ( .B1(n14329), .B2(n13808), .A(n13658), .ZN(n13659) );
  OAI21_X1 U15898 ( .B1(n13660), .B2(n13796), .A(n13659), .ZN(P2_U3191) );
  INV_X1 U15899 ( .A(n14539), .ZN(n14299) );
  XNOR2_X1 U15900 ( .A(n13662), .B(n13661), .ZN(n13735) );
  NOR2_X1 U15901 ( .A1(n13725), .A2(n13665), .ZN(n13728) );
  NOR2_X1 U15902 ( .A1(n13728), .A2(n13663), .ZN(n13664) );
  AOI211_X1 U15903 ( .C1(n13665), .C2(n13725), .A(n13735), .B(n13664), .ZN(
        n13724) );
  INV_X1 U15904 ( .A(n13666), .ZN(n13667) );
  NOR2_X1 U15905 ( .A1(n13724), .A2(n13667), .ZN(n13670) );
  OAI211_X1 U15906 ( .C1(n13670), .C2(n13669), .A(n13668), .B(n13798), .ZN(
        n13675) );
  OAI22_X1 U15907 ( .A1(n13671), .A2(n14474), .B1(n13909), .B2(n14472), .ZN(
        n14292) );
  OAI22_X1 U15908 ( .A1(n13804), .A2(n14296), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13672), .ZN(n13673) );
  AOI21_X1 U15909 ( .B1(n14292), .B2(n13730), .A(n13673), .ZN(n13674) );
  OAI211_X1 U15910 ( .C1(n14299), .C2(n13733), .A(n13675), .B(n13674), .ZN(
        P2_U3195) );
  OAI21_X1 U15911 ( .B1(n13678), .B2(n13677), .A(n13676), .ZN(n13679) );
  NAND2_X1 U15912 ( .A1(n13679), .A2(n13798), .ZN(n13684) );
  NAND2_X1 U15913 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n15703)
         );
  INV_X1 U15914 ( .A(n15703), .ZN(n13682) );
  INV_X1 U15915 ( .A(n13680), .ZN(n14455) );
  OAI22_X1 U15916 ( .A1(n14411), .A2(n13803), .B1(n13804), .B2(n14455), .ZN(
        n13681) );
  AOI211_X1 U15917 ( .C1(n13770), .C2(n14450), .A(n13682), .B(n13681), .ZN(
        n13683) );
  OAI211_X1 U15918 ( .C1(n14458), .C2(n13733), .A(n13684), .B(n13683), .ZN(
        P2_U3196) );
  NAND3_X1 U15919 ( .A1(n13685), .A2(n13799), .A3(n10559), .ZN(n13689) );
  OAI21_X1 U15920 ( .B1(n13713), .B2(n13686), .A(n13798), .ZN(n13688) );
  INV_X1 U15921 ( .A(n13783), .ZN(n13687) );
  AOI21_X1 U15922 ( .B1(n13689), .B2(n13688), .A(n13687), .ZN(n13695) );
  AOI22_X1 U15923 ( .A1(n14232), .A2(n13750), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(n6510), .ZN(n13693) );
  NAND2_X1 U15924 ( .A1(n14088), .A2(n14449), .ZN(n13691) );
  OR2_X1 U15925 ( .A1(n14262), .A2(n14472), .ZN(n13690) );
  NAND2_X1 U15926 ( .A1(n13691), .A2(n13690), .ZN(n14237) );
  NAND2_X1 U15927 ( .A1(n14237), .A2(n13730), .ZN(n13692) );
  OAI211_X1 U15928 ( .C1(n14234), .C2(n13733), .A(n13693), .B(n13692), .ZN(
        n13694) );
  OR2_X1 U15929 ( .A1(n13695), .A2(n13694), .ZN(P2_U3197) );
  NAND2_X1 U15930 ( .A1(n13697), .A2(n13696), .ZN(n13701) );
  XNOR2_X1 U15931 ( .A(n13698), .B(n13699), .ZN(n13800) );
  OAI22_X1 U15932 ( .A1(n13800), .A2(n13797), .B1(n13699), .B2(n13698), .ZN(
        n13700) );
  XOR2_X1 U15933 ( .A(n13701), .B(n13700), .Z(n13705) );
  NAND2_X1 U15934 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n15740)
         );
  OAI21_X1 U15935 ( .B1(n13805), .B2(n14412), .A(n15740), .ZN(n13703) );
  OAI22_X1 U15936 ( .A1(n14376), .A2(n13803), .B1(n13804), .B2(n14379), .ZN(
        n13702) );
  AOI211_X1 U15937 ( .C1(n14568), .C2(n13808), .A(n13703), .B(n13702), .ZN(
        n13704) );
  OAI21_X1 U15938 ( .B1(n13705), .B2(n13796), .A(n13704), .ZN(P2_U3198) );
  OAI21_X1 U15939 ( .B1(n13708), .B2(n13707), .A(n13706), .ZN(n13709) );
  NAND2_X1 U15940 ( .A1(n13709), .A2(n13798), .ZN(n13712) );
  AND2_X1 U15941 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n14147) );
  OAI22_X1 U15942 ( .A1(n10517), .A2(n13803), .B1(n13804), .B2(n14365), .ZN(
        n13710) );
  AOI211_X1 U15943 ( .C1(n13770), .C2(n14398), .A(n14147), .B(n13710), .ZN(
        n13711) );
  OAI211_X1 U15944 ( .C1(n7662), .C2(n13733), .A(n13712), .B(n13711), .ZN(
        P2_U3200) );
  AOI211_X1 U15945 ( .C1(n13715), .C2(n13714), .A(n13796), .B(n13713), .ZN(
        n13716) );
  INV_X1 U15946 ( .A(n13716), .ZN(n13723) );
  OAI22_X1 U15947 ( .A1(n13718), .A2(n14474), .B1(n13717), .B2(n14472), .ZN(
        n14246) );
  INV_X1 U15948 ( .A(n14254), .ZN(n13720) );
  OAI22_X1 U15949 ( .A1(n13720), .A2(n13804), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13719), .ZN(n13721) );
  AOI21_X1 U15950 ( .B1(n14246), .B2(n13730), .A(n13721), .ZN(n13722) );
  OAI211_X1 U15951 ( .C1(n14257), .C2(n13733), .A(n13723), .B(n13722), .ZN(
        P2_U3201) );
  INV_X1 U15952 ( .A(n13724), .ZN(n13738) );
  INV_X1 U15953 ( .A(n13725), .ZN(n13727) );
  OAI33_X1 U15954 ( .A1(n13758), .A2(n13907), .A3(n13728), .B1(n13796), .B2(
        n13727), .B3(n13726), .ZN(n13736) );
  OAI22_X1 U15955 ( .A1(n13729), .A2(n14474), .B1(n13907), .B2(n14472), .ZN(
        n14306) );
  AOI22_X1 U15956 ( .A1(n14306), .A2(n13730), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(n6510), .ZN(n13732) );
  NAND2_X1 U15957 ( .A1(n13750), .A2(n14313), .ZN(n13731) );
  OAI211_X1 U15958 ( .C1(n14316), .C2(n13733), .A(n13732), .B(n13731), .ZN(
        n13734) );
  AOI21_X1 U15959 ( .B1(n13736), .B2(n13735), .A(n13734), .ZN(n13737) );
  OAI21_X1 U15960 ( .B1(n13738), .B2(n13796), .A(n13737), .ZN(P2_U3205) );
  XNOR2_X1 U15961 ( .A(n13740), .B(n13739), .ZN(n13746) );
  OAI22_X1 U15962 ( .A1(n13805), .A2(n14475), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13741), .ZN(n13744) );
  INV_X1 U15963 ( .A(n14433), .ZN(n13742) );
  OAI22_X1 U15964 ( .A1(n14427), .A2(n13803), .B1(n13804), .B2(n13742), .ZN(
        n13743) );
  AOI211_X1 U15965 ( .C1(n14432), .C2(n13808), .A(n13744), .B(n13743), .ZN(
        n13745) );
  OAI21_X1 U15966 ( .B1(n13746), .B2(n13796), .A(n13745), .ZN(P2_U3206) );
  INV_X1 U15967 ( .A(n13747), .ZN(n13748) );
  AOI22_X1 U15968 ( .A1(n13748), .A2(n13798), .B1(n13799), .B2(n14263), .ZN(
        n13755) );
  INV_X1 U15969 ( .A(n13749), .ZN(n13754) );
  AOI22_X1 U15970 ( .A1(n14090), .A2(n14449), .B1(n14451), .B2(n14091), .ZN(
        n14279) );
  AOI22_X1 U15971 ( .A1(n14285), .A2(n13750), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13751) );
  OAI21_X1 U15972 ( .B1(n14279), .B2(n13789), .A(n13751), .ZN(n13752) );
  AOI21_X1 U15973 ( .B1(n14284), .B2(n13808), .A(n13752), .ZN(n13753) );
  OAI21_X1 U15974 ( .B1(n13755), .B2(n13754), .A(n13753), .ZN(P2_U3207) );
  INV_X1 U15975 ( .A(n13767), .ZN(n13760) );
  XNOR2_X1 U15976 ( .A(n13757), .B(n13756), .ZN(n13764) );
  OAI22_X1 U15977 ( .A1(n13758), .A2(n13816), .B1(n13761), .B2(n13796), .ZN(
        n13759) );
  NAND3_X1 U15978 ( .A1(n13760), .A2(n13764), .A3(n13759), .ZN(n13774) );
  INV_X1 U15979 ( .A(n13761), .ZN(n13763) );
  NOR2_X1 U15980 ( .A1(n13763), .A2(n13762), .ZN(n13766) );
  INV_X1 U15981 ( .A(n13764), .ZN(n13765) );
  OAI211_X1 U15982 ( .C1(n13767), .C2(n13766), .A(n13798), .B(n13765), .ZN(
        n13773) );
  AOI22_X1 U15983 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(n13768), .B1(n13808), 
        .B2(n13813), .ZN(n13772) );
  AOI22_X1 U15984 ( .A1(n13770), .A2(n14104), .B1(n13769), .B2(n14101), .ZN(
        n13771) );
  NAND4_X1 U15985 ( .A1(n13774), .A2(n13773), .A3(n13772), .A4(n13771), .ZN(
        P2_U3209) );
  XNOR2_X1 U15986 ( .A(n13776), .B(n13775), .ZN(n13780) );
  NAND2_X1 U15987 ( .A1(n6510), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n15753) );
  OAI21_X1 U15988 ( .B1(n13805), .B2(n14376), .A(n15753), .ZN(n13778) );
  OAI22_X1 U15989 ( .A1(n13907), .A2(n13803), .B1(n13804), .B2(n14344), .ZN(
        n13777) );
  AOI211_X1 U15990 ( .C1(n14351), .C2(n13808), .A(n13778), .B(n13777), .ZN(
        n13779) );
  OAI21_X1 U15991 ( .B1(n13780), .B2(n13796), .A(n13779), .ZN(P2_U3210) );
  NAND3_X1 U15992 ( .A1(n13781), .A2(n13799), .A3(n14089), .ZN(n13782) );
  OAI21_X1 U15993 ( .B1(n13783), .B2(n13796), .A(n13782), .ZN(n13786) );
  INV_X1 U15994 ( .A(n13784), .ZN(n13785) );
  NAND2_X1 U15995 ( .A1(n13786), .A2(n13785), .ZN(n13794) );
  OR2_X1 U15996 ( .A1(n13993), .A2(n14474), .ZN(n13788) );
  NAND2_X1 U15997 ( .A1(n14089), .A2(n14451), .ZN(n13787) );
  AND2_X1 U15998 ( .A1(n13788), .A2(n13787), .ZN(n14226) );
  NOR2_X1 U15999 ( .A1(n14226), .A2(n13789), .ZN(n13792) );
  OAI22_X1 U16000 ( .A1(n14219), .A2(n13804), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13790), .ZN(n13791) );
  AOI211_X1 U16001 ( .C1(n14217), .C2(n13808), .A(n13792), .B(n13791), .ZN(
        n13793) );
  OAI211_X1 U16002 ( .C1(n13796), .C2(n13795), .A(n13794), .B(n13793), .ZN(
        P2_U3212) );
  NAND2_X1 U16003 ( .A1(n13798), .A2(n13797), .ZN(n13802) );
  NAND2_X1 U16004 ( .A1(n13799), .A2(n14093), .ZN(n13801) );
  MUX2_X1 U16005 ( .A(n13802), .B(n13801), .S(n13800), .Z(n13810) );
  OAI22_X1 U16006 ( .A1(n13803), .A2(n14361), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6971), .ZN(n13807) );
  OAI22_X1 U16007 ( .A1(n14427), .A2(n13805), .B1(n13804), .B2(n14388), .ZN(
        n13806) );
  AOI211_X1 U16008 ( .C1(n14393), .C2(n13808), .A(n13807), .B(n13806), .ZN(
        n13809) );
  NAND2_X1 U16009 ( .A1(n13810), .A2(n13809), .ZN(P2_U3213) );
  AOI22_X1 U16010 ( .A1(n14102), .A2(n13991), .B1(n14022), .B2(n13813), .ZN(
        n13827) );
  OR2_X1 U16011 ( .A1(n10389), .A2(n6520), .ZN(n13815) );
  NAND2_X1 U16012 ( .A1(n13991), .A2(n13813), .ZN(n13814) );
  NAND2_X1 U16013 ( .A1(n13815), .A2(n13814), .ZN(n13826) );
  NAND2_X1 U16014 ( .A1(n6511), .A2(n10379), .ZN(n13817) );
  AOI22_X1 U16015 ( .A1(n14104), .A2(n13991), .B1(n14022), .B2(n10379), .ZN(
        n13825) );
  OAI22_X1 U16016 ( .A1(n13827), .A2(n13826), .B1(n13824), .B2(n13825), .ZN(
        n13831) );
  OAI211_X1 U16017 ( .C1(n13820), .C2(n14068), .A(n13819), .B(n6511), .ZN(
        n13823) );
  AOI21_X1 U16018 ( .B1(n13819), .B2(n13820), .A(n6520), .ZN(n13821) );
  OAI22_X1 U16019 ( .A1(n13821), .A2(n14068), .B1(n14022), .B2(n13820), .ZN(
        n13822) );
  AOI22_X1 U16020 ( .A1(n13825), .A2(n13824), .B1(n13823), .B2(n13822), .ZN(
        n13830) );
  INV_X1 U16021 ( .A(n13826), .ZN(n13829) );
  INV_X1 U16022 ( .A(n13827), .ZN(n13828) );
  OAI22_X1 U16023 ( .A1(n13831), .A2(n13830), .B1(n13829), .B2(n13828), .ZN(
        n13841) );
  NAND2_X1 U16024 ( .A1(n14101), .A2(n14022), .ZN(n13833) );
  NAND2_X1 U16025 ( .A1(n13991), .A2(n7648), .ZN(n13832) );
  AND2_X1 U16026 ( .A1(n13833), .A2(n13832), .ZN(n13837) );
  NAND2_X1 U16027 ( .A1(n14101), .A2(n6511), .ZN(n13835) );
  NAND2_X1 U16028 ( .A1(n14022), .A2(n7648), .ZN(n13834) );
  NAND2_X1 U16029 ( .A1(n13835), .A2(n13834), .ZN(n13836) );
  NOR2_X1 U16030 ( .A1(n13837), .A2(n13836), .ZN(n13840) );
  INV_X1 U16031 ( .A(n13836), .ZN(n13839) );
  INV_X1 U16032 ( .A(n13837), .ZN(n13838) );
  OAI22_X1 U16033 ( .A1(n13841), .A2(n13840), .B1(n13839), .B2(n13838), .ZN(
        n13846) );
  OAI22_X1 U16034 ( .A1(n13842), .A2(n6560), .B1(n15806), .B2(n6520), .ZN(
        n13847) );
  AOI22_X1 U16035 ( .A1(n13843), .A2(n13991), .B1(n14100), .B2(n14022), .ZN(
        n13844) );
  INV_X1 U16036 ( .A(n13847), .ZN(n13848) );
  OAI22_X1 U16037 ( .A1(n13850), .A2(n6560), .B1(n13849), .B2(n6520), .ZN(
        n13852) );
  OAI22_X1 U16038 ( .A1(n13850), .A2(n6520), .B1(n13849), .B2(n6560), .ZN(
        n13854) );
  INV_X1 U16039 ( .A(n13852), .ZN(n13853) );
  AOI22_X1 U16040 ( .A1(n14022), .A2(n15764), .B1(n14098), .B2(n13991), .ZN(
        n13857) );
  OAI22_X1 U16041 ( .A1(n15824), .A2(n13892), .B1(n13855), .B2(n6520), .ZN(
        n13856) );
  AOI22_X1 U16042 ( .A1(n13858), .A2(n6511), .B1(n14022), .B2(n14097), .ZN(
        n13861) );
  OAI22_X1 U16043 ( .A1(n7911), .A2(n6520), .B1(n13859), .B2(n13892), .ZN(
        n13860) );
  OAI21_X1 U16044 ( .B1(n13862), .B2(n13861), .A(n13860), .ZN(n13864) );
  NAND2_X1 U16045 ( .A1(n13862), .A2(n13861), .ZN(n13863) );
  OAI22_X1 U16046 ( .A1(n10221), .A2(n6520), .B1(n13865), .B2(n13892), .ZN(
        n13867) );
  AOI22_X1 U16047 ( .A1(n7205), .A2(n6511), .B1(n14022), .B2(n14096), .ZN(
        n13866) );
  OAI22_X1 U16048 ( .A1(n13869), .A2(n13892), .B1(n13868), .B2(n6520), .ZN(
        n13872) );
  AOI22_X1 U16049 ( .A1(n13870), .A2(n14022), .B1(n8009), .B2(n13991), .ZN(
        n13871) );
  OAI22_X1 U16050 ( .A1(n7655), .A2(n6520), .B1(n14473), .B2(n13892), .ZN(
        n13874) );
  AOI22_X1 U16051 ( .A1(n14605), .A2(n13991), .B1(n14022), .B2(n14095), .ZN(
        n13873) );
  NOR2_X1 U16052 ( .A1(n13875), .A2(n13874), .ZN(n13876) );
  NOR2_X1 U16053 ( .A1(n13877), .A2(n13876), .ZN(n13881) );
  AOI22_X1 U16054 ( .A1(n14483), .A2(n6511), .B1(n14022), .B2(n14450), .ZN(
        n13880) );
  OAI22_X1 U16055 ( .A1(n14653), .A2(n6520), .B1(n13878), .B2(n13892), .ZN(
        n13879) );
  OAI21_X1 U16056 ( .B1(n13881), .B2(n13880), .A(n13879), .ZN(n13883) );
  NAND2_X1 U16057 ( .A1(n13881), .A2(n13880), .ZN(n13882) );
  OAI22_X1 U16058 ( .A1(n14458), .A2(n6520), .B1(n14475), .B2(n13892), .ZN(
        n13885) );
  OAI22_X1 U16059 ( .A1(n14458), .A2(n13892), .B1(n14475), .B2(n6520), .ZN(
        n13884) );
  INV_X1 U16060 ( .A(n13885), .ZN(n13886) );
  OAI22_X1 U16061 ( .A1(n14645), .A2(n13892), .B1(n14411), .B2(n6520), .ZN(
        n13887) );
  INV_X1 U16062 ( .A(n13887), .ZN(n13891) );
  NAND2_X1 U16063 ( .A1(n13888), .A2(n13887), .ZN(n13890) );
  OAI22_X1 U16064 ( .A1(n14645), .A2(n6520), .B1(n14411), .B2(n13892), .ZN(
        n13889) );
  OAI22_X1 U16065 ( .A1(n14418), .A2(n6520), .B1(n14427), .B2(n13892), .ZN(
        n13893) );
  OAI22_X1 U16066 ( .A1(n14418), .A2(n13892), .B1(n14427), .B2(n6520), .ZN(
        n13894) );
  AOI22_X1 U16067 ( .A1(n14393), .A2(n13991), .B1(n14022), .B2(n14093), .ZN(
        n13896) );
  OAI22_X1 U16068 ( .A1(n14573), .A2(n6520), .B1(n14412), .B2(n13892), .ZN(
        n13895) );
  NAND2_X1 U16069 ( .A1(n13897), .A2(n13896), .ZN(n13898) );
  OAI22_X1 U16070 ( .A1(n7663), .A2(n6520), .B1(n14361), .B2(n13892), .ZN(
        n13900) );
  OAI22_X1 U16071 ( .A1(n7663), .A2(n13892), .B1(n14361), .B2(n6520), .ZN(
        n13901) );
  AOI22_X1 U16072 ( .A1(n14364), .A2(n13991), .B1(n14022), .B2(n14339), .ZN(
        n13902) );
  AOI22_X1 U16073 ( .A1(n14364), .A2(n14022), .B1(n14339), .B2(n6511), .ZN(
        n13903) );
  OAI22_X1 U16074 ( .A1(n10518), .A2(n6520), .B1(n10517), .B2(n13892), .ZN(
        n13906) );
  OAI22_X1 U16075 ( .A1(n10518), .A2(n13892), .B1(n10517), .B2(n6520), .ZN(
        n13904) );
  OAI22_X1 U16076 ( .A1(n14632), .A2(n13892), .B1(n13907), .B2(n6520), .ZN(
        n13928) );
  NOR2_X1 U16077 ( .A1(n13909), .A2(n6520), .ZN(n13908) );
  AOI21_X1 U16078 ( .B1(n14544), .B2(n13991), .A(n13908), .ZN(n13931) );
  NAND2_X1 U16079 ( .A1(n14544), .A2(n14022), .ZN(n13911) );
  OR2_X1 U16080 ( .A1(n13909), .A2(n13892), .ZN(n13910) );
  NAND2_X1 U16081 ( .A1(n13911), .A2(n13910), .ZN(n13930) );
  NOR2_X1 U16082 ( .A1(n14262), .A2(n6520), .ZN(n13912) );
  AOI21_X1 U16083 ( .B1(n14522), .B2(n13991), .A(n13912), .ZN(n13944) );
  NAND2_X1 U16084 ( .A1(n14522), .A2(n14022), .ZN(n13914) );
  OR2_X1 U16085 ( .A1(n14262), .A2(n13892), .ZN(n13913) );
  NAND2_X1 U16086 ( .A1(n13914), .A2(n13913), .ZN(n13943) );
  NAND2_X1 U16087 ( .A1(n13944), .A2(n13943), .ZN(n13948) );
  AND2_X1 U16088 ( .A1(n14090), .A2(n14022), .ZN(n13915) );
  AOI21_X1 U16089 ( .B1(n14528), .B2(n13991), .A(n13915), .ZN(n13940) );
  NAND2_X1 U16090 ( .A1(n14528), .A2(n14022), .ZN(n13917) );
  NAND2_X1 U16091 ( .A1(n14090), .A2(n13991), .ZN(n13916) );
  NAND2_X1 U16092 ( .A1(n13917), .A2(n13916), .ZN(n13939) );
  NAND2_X1 U16093 ( .A1(n13940), .A2(n13939), .ZN(n13918) );
  AND2_X1 U16094 ( .A1(n14263), .A2(n14022), .ZN(n13919) );
  AOI21_X1 U16095 ( .B1(n14284), .B2(n6511), .A(n13919), .ZN(n13950) );
  NAND2_X1 U16096 ( .A1(n14284), .A2(n14022), .ZN(n13921) );
  NAND2_X1 U16097 ( .A1(n14263), .A2(n6511), .ZN(n13920) );
  NAND2_X1 U16098 ( .A1(n13921), .A2(n13920), .ZN(n13949) );
  AND2_X1 U16099 ( .A1(n14091), .A2(n14022), .ZN(n13922) );
  AOI21_X1 U16100 ( .B1(n14539), .B2(n13991), .A(n13922), .ZN(n13936) );
  NAND2_X1 U16101 ( .A1(n14539), .A2(n14022), .ZN(n13924) );
  NAND2_X1 U16102 ( .A1(n14091), .A2(n6511), .ZN(n13923) );
  NAND2_X1 U16103 ( .A1(n13924), .A2(n13923), .ZN(n13935) );
  AND2_X1 U16104 ( .A1(n13936), .A2(n13935), .ZN(n13925) );
  AOI22_X1 U16105 ( .A1(n14329), .A2(n14022), .B1(n14340), .B2(n6511), .ZN(
        n13927) );
  INV_X1 U16106 ( .A(n13929), .ZN(n13934) );
  INV_X1 U16107 ( .A(n13930), .ZN(n13933) );
  INV_X1 U16108 ( .A(n13931), .ZN(n13932) );
  INV_X1 U16109 ( .A(n13935), .ZN(n13938) );
  INV_X1 U16110 ( .A(n13936), .ZN(n13937) );
  NAND2_X1 U16111 ( .A1(n13938), .A2(n13937), .ZN(n13954) );
  INV_X1 U16112 ( .A(n13939), .ZN(n13942) );
  INV_X1 U16113 ( .A(n13940), .ZN(n13941) );
  AND2_X1 U16114 ( .A1(n13942), .A2(n13941), .ZN(n13947) );
  INV_X1 U16115 ( .A(n13943), .ZN(n13946) );
  INV_X1 U16116 ( .A(n13944), .ZN(n13945) );
  OR3_X1 U16117 ( .A1(n13951), .A2(n13950), .A3(n13949), .ZN(n13952) );
  OAI211_X1 U16118 ( .C1(n13955), .C2(n13954), .A(n13953), .B(n13952), .ZN(
        n13956) );
  INV_X1 U16119 ( .A(n13956), .ZN(n13965) );
  AND2_X1 U16120 ( .A1(n14088), .A2(n6511), .ZN(n13957) );
  AOI21_X1 U16121 ( .B1(n14217), .B2(n14022), .A(n13957), .ZN(n14001) );
  NAND2_X1 U16122 ( .A1(n14217), .A2(n6511), .ZN(n13959) );
  NAND2_X1 U16123 ( .A1(n14088), .A2(n14022), .ZN(n13958) );
  NAND2_X1 U16124 ( .A1(n13959), .A2(n13958), .ZN(n14000) );
  NAND2_X1 U16125 ( .A1(n14001), .A2(n14000), .ZN(n13998) );
  OR2_X1 U16126 ( .A1(n14234), .A2(n6520), .ZN(n13961) );
  NAND2_X1 U16127 ( .A1(n14089), .A2(n13991), .ZN(n13960) );
  AND2_X1 U16128 ( .A1(n13961), .A2(n13960), .ZN(n13995) );
  OR2_X1 U16129 ( .A1(n14234), .A2(n13892), .ZN(n13963) );
  NAND2_X1 U16130 ( .A1(n14089), .A2(n14022), .ZN(n13962) );
  NAND2_X1 U16131 ( .A1(n13963), .A2(n13962), .ZN(n13994) );
  NAND2_X1 U16132 ( .A1(n13995), .A2(n13994), .ZN(n13964) );
  NAND2_X1 U16133 ( .A1(n10315), .A2(n11791), .ZN(n14074) );
  NAND3_X1 U16134 ( .A1(n14074), .A2(n14066), .A3(n13966), .ZN(n13967) );
  AOI21_X1 U16135 ( .B1(n14085), .B2(n6511), .A(n13967), .ZN(n13974) );
  NAND2_X1 U16136 ( .A1(n6512), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n13973) );
  NAND2_X1 U16137 ( .A1(n7281), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n13972) );
  NAND2_X1 U16138 ( .A1(n13970), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n13971) );
  AND3_X1 U16139 ( .A1(n13973), .A2(n13972), .A3(n13971), .ZN(n14195) );
  NOR2_X1 U16140 ( .A1(n13974), .A2(n14195), .ZN(n13975) );
  AOI21_X1 U16141 ( .B1(n14060), .B2(n14022), .A(n13975), .ZN(n14015) );
  NAND2_X1 U16142 ( .A1(n14060), .A2(n6511), .ZN(n13977) );
  INV_X1 U16143 ( .A(n14195), .ZN(n14086) );
  NAND2_X1 U16144 ( .A1(n14086), .A2(n14022), .ZN(n13976) );
  NAND2_X1 U16145 ( .A1(n13977), .A2(n13976), .ZN(n14014) );
  NOR2_X1 U16146 ( .A1(n14059), .A2(n13892), .ZN(n13978) );
  AOI21_X1 U16147 ( .B1(n14505), .B2(n14022), .A(n13978), .ZN(n14010) );
  NAND2_X1 U16148 ( .A1(n14505), .A2(n13991), .ZN(n13980) );
  OR2_X1 U16149 ( .A1(n14059), .A2(n6520), .ZN(n13979) );
  NAND2_X1 U16150 ( .A1(n13980), .A2(n13979), .ZN(n14009) );
  INV_X1 U16151 ( .A(n13981), .ZN(n13982) );
  AOI22_X1 U16152 ( .A1(n14085), .A2(n14022), .B1(n13991), .B2(n13982), .ZN(
        n13985) );
  NAND2_X1 U16153 ( .A1(n13983), .A2(n13991), .ZN(n13984) );
  OAI211_X1 U16154 ( .C1(n14025), .C2(n14085), .A(n13985), .B(n13984), .ZN(
        n13986) );
  NOR2_X1 U16155 ( .A1(n14196), .A2(n6520), .ZN(n13987) );
  AOI21_X1 U16156 ( .B1(n14184), .B2(n13991), .A(n13987), .ZN(n14013) );
  NAND2_X1 U16157 ( .A1(n14184), .A2(n14022), .ZN(n13989) );
  NAND2_X1 U16158 ( .A1(n14183), .A2(n6511), .ZN(n13988) );
  NAND2_X1 U16159 ( .A1(n13989), .A2(n13988), .ZN(n14012) );
  NAND2_X1 U16160 ( .A1(n14013), .A2(n14012), .ZN(n13990) );
  INV_X1 U16161 ( .A(n13993), .ZN(n14087) );
  AOI22_X1 U16162 ( .A1(n13992), .A2(n6511), .B1(n14022), .B2(n14087), .ZN(
        n14005) );
  OAI22_X1 U16163 ( .A1(n14511), .A2(n6520), .B1(n13993), .B2(n13892), .ZN(
        n14006) );
  INV_X1 U16164 ( .A(n13994), .ZN(n13997) );
  INV_X1 U16165 ( .A(n13995), .ZN(n13996) );
  NAND3_X1 U16166 ( .A1(n13998), .A2(n13997), .A3(n13996), .ZN(n13999) );
  OAI21_X1 U16167 ( .B1(n14001), .B2(n14000), .A(n13999), .ZN(n14002) );
  AOI21_X1 U16168 ( .B1(n14005), .B2(n14006), .A(n14002), .ZN(n14003) );
  INV_X1 U16169 ( .A(n14004), .ZN(n14020) );
  INV_X1 U16170 ( .A(n14005), .ZN(n14008) );
  INV_X1 U16171 ( .A(n14006), .ZN(n14007) );
  NAND2_X1 U16172 ( .A1(n14008), .A2(n14007), .ZN(n14019) );
  NAND2_X1 U16173 ( .A1(n14010), .A2(n14009), .ZN(n14011) );
  AOI22_X1 U16174 ( .A1(n14017), .A2(n14016), .B1(n14015), .B2(n14014), .ZN(
        n14018) );
  NOR2_X1 U16175 ( .A1(n14085), .A2(n14022), .ZN(n14026) );
  NOR3_X1 U16176 ( .A1(n14025), .A2(n14023), .A3(n13991), .ZN(n14024) );
  AOI21_X1 U16177 ( .B1(n14026), .B2(n14025), .A(n14024), .ZN(n14027) );
  OR2_X1 U16178 ( .A1(n14030), .A2(n14029), .ZN(n14270) );
  INV_X1 U16179 ( .A(n14031), .ZN(n14033) );
  XNOR2_X1 U16180 ( .A(n14588), .B(n14475), .ZN(n14442) );
  AND4_X1 U16181 ( .A1(n14036), .A2(n14065), .A3(n15774), .A4(n14035), .ZN(
        n14040) );
  AND4_X1 U16182 ( .A1(n14040), .A2(n14039), .A3(n14038), .A4(n14037), .ZN(
        n14043) );
  INV_X1 U16183 ( .A(n15765), .ZN(n14041) );
  NAND4_X1 U16184 ( .A1(n14044), .A2(n14043), .A3(n14042), .A4(n14041), .ZN(
        n14045) );
  NOR2_X1 U16185 ( .A1(n14046), .A2(n14045), .ZN(n14048) );
  NAND3_X1 U16186 ( .A1(n14470), .A2(n14048), .A3(n14047), .ZN(n14049) );
  NOR2_X1 U16187 ( .A1(n14442), .A2(n14049), .ZN(n14050) );
  NAND4_X1 U16188 ( .A1(n14409), .A2(n14050), .A3(n14429), .A4(n14374), .ZN(
        n14052) );
  NOR2_X1 U16189 ( .A1(n14052), .A2(n14051), .ZN(n14053) );
  NAND4_X1 U16190 ( .A1(n14300), .A2(n14053), .A3(n14338), .A4(n14394), .ZN(
        n14054) );
  NOR2_X1 U16191 ( .A1(n14054), .A2(n14309), .ZN(n14055) );
  XNOR2_X1 U16192 ( .A(n14329), .B(n14340), .ZN(n14323) );
  NAND4_X1 U16193 ( .A1(n14270), .A2(n14055), .A3(n14282), .A4(n14323), .ZN(
        n14056) );
  NOR2_X1 U16194 ( .A1(n14056), .A2(n14249), .ZN(n14057) );
  XOR2_X1 U16195 ( .A(n14195), .B(n14060), .Z(n14061) );
  XNOR2_X1 U16196 ( .A(n14062), .B(n14076), .ZN(n14063) );
  INV_X1 U16197 ( .A(n14073), .ZN(n14078) );
  AOI21_X1 U16198 ( .B1(n14066), .B2(n14076), .A(n14070), .ZN(n14067) );
  OAI21_X1 U16199 ( .B1(n14068), .B2(n10315), .A(n14067), .ZN(n14069) );
  NAND4_X1 U16200 ( .A1(n14451), .A2(n14071), .A3(n14070), .A4(n15796), .ZN(
        n14072) );
  OAI211_X1 U16201 ( .C1(n10315), .C2(n14073), .A(n14072), .B(P2_B_REG_SCAN_IN), .ZN(n14082) );
  INV_X1 U16202 ( .A(n14074), .ZN(n14081) );
  NOR3_X1 U16203 ( .A1(n14077), .A2(n14076), .A3(n14075), .ZN(n14080) );
  MUX2_X1 U16204 ( .A(n14085), .B(P2_DATAO_REG_31__SCAN_IN), .S(n14103), .Z(
        P2_U3562) );
  MUX2_X1 U16205 ( .A(n14086), .B(P2_DATAO_REG_30__SCAN_IN), .S(n14103), .Z(
        P2_U3561) );
  MUX2_X1 U16206 ( .A(n14183), .B(P2_DATAO_REG_28__SCAN_IN), .S(n14103), .Z(
        P2_U3559) );
  MUX2_X1 U16207 ( .A(n14087), .B(P2_DATAO_REG_27__SCAN_IN), .S(n14103), .Z(
        P2_U3558) );
  MUX2_X1 U16208 ( .A(n14088), .B(P2_DATAO_REG_26__SCAN_IN), .S(n14103), .Z(
        P2_U3557) );
  MUX2_X1 U16209 ( .A(n14089), .B(P2_DATAO_REG_25__SCAN_IN), .S(n14103), .Z(
        P2_U3556) );
  MUX2_X1 U16210 ( .A(n10559), .B(P2_DATAO_REG_24__SCAN_IN), .S(n14103), .Z(
        P2_U3555) );
  MUX2_X1 U16211 ( .A(n14090), .B(P2_DATAO_REG_23__SCAN_IN), .S(n14103), .Z(
        P2_U3554) );
  MUX2_X1 U16212 ( .A(n14263), .B(P2_DATAO_REG_22__SCAN_IN), .S(n14103), .Z(
        P2_U3553) );
  MUX2_X1 U16213 ( .A(n14091), .B(P2_DATAO_REG_21__SCAN_IN), .S(n14103), .Z(
        P2_U3552) );
  MUX2_X1 U16214 ( .A(n14340), .B(P2_DATAO_REG_19__SCAN_IN), .S(n14103), .Z(
        P2_U3550) );
  MUX2_X1 U16215 ( .A(n14092), .B(P2_DATAO_REG_18__SCAN_IN), .S(n14103), .Z(
        P2_U3549) );
  MUX2_X1 U16216 ( .A(n14339), .B(P2_DATAO_REG_17__SCAN_IN), .S(n14103), .Z(
        P2_U3548) );
  MUX2_X1 U16217 ( .A(n14398), .B(P2_DATAO_REG_16__SCAN_IN), .S(n14103), .Z(
        P2_U3547) );
  MUX2_X1 U16218 ( .A(n14093), .B(P2_DATAO_REG_15__SCAN_IN), .S(n14103), .Z(
        P2_U3546) );
  MUX2_X1 U16219 ( .A(n14397), .B(P2_DATAO_REG_14__SCAN_IN), .S(n14103), .Z(
        P2_U3545) );
  MUX2_X1 U16220 ( .A(n14448), .B(P2_DATAO_REG_13__SCAN_IN), .S(n14103), .Z(
        P2_U3544) );
  MUX2_X1 U16221 ( .A(n14094), .B(P2_DATAO_REG_12__SCAN_IN), .S(n14103), .Z(
        P2_U3543) );
  MUX2_X1 U16222 ( .A(n14450), .B(P2_DATAO_REG_11__SCAN_IN), .S(n14103), .Z(
        P2_U3542) );
  MUX2_X1 U16223 ( .A(n14095), .B(P2_DATAO_REG_10__SCAN_IN), .S(n14103), .Z(
        P2_U3541) );
  MUX2_X1 U16224 ( .A(n8009), .B(P2_DATAO_REG_9__SCAN_IN), .S(n14103), .Z(
        P2_U3540) );
  MUX2_X1 U16225 ( .A(n14096), .B(P2_DATAO_REG_8__SCAN_IN), .S(n14103), .Z(
        P2_U3539) );
  MUX2_X1 U16226 ( .A(n14097), .B(P2_DATAO_REG_7__SCAN_IN), .S(n14103), .Z(
        P2_U3538) );
  MUX2_X1 U16227 ( .A(n14098), .B(P2_DATAO_REG_6__SCAN_IN), .S(n14103), .Z(
        P2_U3537) );
  MUX2_X1 U16228 ( .A(n14099), .B(P2_DATAO_REG_5__SCAN_IN), .S(n14103), .Z(
        P2_U3536) );
  MUX2_X1 U16229 ( .A(n14100), .B(P2_DATAO_REG_4__SCAN_IN), .S(n14103), .Z(
        P2_U3535) );
  MUX2_X1 U16230 ( .A(n14101), .B(P2_DATAO_REG_3__SCAN_IN), .S(n14103), .Z(
        P2_U3534) );
  MUX2_X1 U16231 ( .A(n14102), .B(P2_DATAO_REG_2__SCAN_IN), .S(n14103), .Z(
        P2_U3533) );
  MUX2_X1 U16232 ( .A(n14104), .B(P2_DATAO_REG_1__SCAN_IN), .S(n14103), .Z(
        P2_U3532) );
  OAI22_X1 U16233 ( .A1(n15749), .A2(n14105), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7878), .ZN(n14106) );
  AOI21_X1 U16234 ( .B1(n15600), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n14106), .ZN(
        n14115) );
  OAI211_X1 U16235 ( .C1(n14109), .C2(n14108), .A(n15744), .B(n14107), .ZN(
        n14114) );
  OAI211_X1 U16236 ( .C1(n14112), .C2(n14111), .A(n15752), .B(n14110), .ZN(
        n14113) );
  NAND3_X1 U16237 ( .A1(n14115), .A2(n14114), .A3(n14113), .ZN(P2_U3215) );
  NAND2_X1 U16238 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n14116) );
  OAI21_X1 U16239 ( .B1(n15749), .B2(n14117), .A(n14116), .ZN(n14118) );
  AOI21_X1 U16240 ( .B1(n15600), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n14118), .ZN(
        n14127) );
  OAI211_X1 U16241 ( .C1(n14121), .C2(n14120), .A(n15752), .B(n14119), .ZN(
        n14126) );
  OAI211_X1 U16242 ( .C1(n14124), .C2(n14123), .A(n15744), .B(n14122), .ZN(
        n14125) );
  NAND3_X1 U16243 ( .A1(n14127), .A2(n14126), .A3(n14125), .ZN(P2_U3217) );
  NAND2_X1 U16244 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(n6510), .ZN(n14128) );
  OAI21_X1 U16245 ( .B1(n15749), .B2(n14129), .A(n14128), .ZN(n14130) );
  AOI21_X1 U16246 ( .B1(n15600), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n14130), .ZN(
        n14139) );
  OAI211_X1 U16247 ( .C1(n14133), .C2(n14132), .A(n15744), .B(n14131), .ZN(
        n14138) );
  OAI211_X1 U16248 ( .C1(n14136), .C2(n14135), .A(n15752), .B(n14134), .ZN(
        n14137) );
  NAND3_X1 U16249 ( .A1(n14139), .A2(n14138), .A3(n14137), .ZN(P2_U3221) );
  XNOR2_X1 U16250 ( .A(n15713), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n15709) );
  INV_X1 U16251 ( .A(n14141), .ZN(n14142) );
  AOI21_X1 U16252 ( .B1(n14155), .B2(n14142), .A(n15716), .ZN(n15735) );
  XNOR2_X1 U16253 ( .A(n15738), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n15734) );
  NOR2_X1 U16254 ( .A1(n15735), .A2(n15734), .ZN(n15732) );
  INV_X1 U16255 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14564) );
  XNOR2_X1 U16256 ( .A(n14159), .B(n14564), .ZN(n14143) );
  AOI211_X1 U16257 ( .C1(n14144), .C2(n14143), .A(n15733), .B(n14164), .ZN(
        n14148) );
  NOR2_X1 U16258 ( .A1(n15755), .A2(n7564), .ZN(n14146) );
  NOR2_X1 U16259 ( .A1(n15749), .A2(n14159), .ZN(n14145) );
  NOR4_X1 U16260 ( .A1(n14148), .A2(n14147), .A3(n14146), .A4(n14145), .ZN(
        n14163) );
  NAND2_X1 U16261 ( .A1(n14149), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n14150) );
  NAND2_X1 U16262 ( .A1(n14151), .A2(n14150), .ZN(n14153) );
  XNOR2_X1 U16263 ( .A(n14153), .B(n14152), .ZN(n15707) );
  NAND2_X1 U16264 ( .A1(n15707), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n15706) );
  NAND2_X1 U16265 ( .A1(n14153), .A2(n15713), .ZN(n14154) );
  NAND2_X1 U16266 ( .A1(n15706), .A2(n14154), .ZN(n14156) );
  XNOR2_X1 U16267 ( .A(n14156), .B(n15723), .ZN(n15720) );
  NAND2_X1 U16268 ( .A1(n15720), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n15719) );
  NAND2_X1 U16269 ( .A1(n14156), .A2(n14155), .ZN(n14157) );
  NAND2_X1 U16270 ( .A1(n15719), .A2(n14157), .ZN(n15730) );
  INV_X1 U16271 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n14380) );
  XNOR2_X1 U16272 ( .A(n15738), .B(n14380), .ZN(n15729) );
  NAND2_X1 U16273 ( .A1(n15730), .A2(n15729), .ZN(n15728) );
  NAND2_X1 U16274 ( .A1(n15738), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n14158) );
  NAND2_X1 U16275 ( .A1(n15728), .A2(n14158), .ZN(n14161) );
  XNOR2_X1 U16276 ( .A(n14159), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n14160) );
  NAND2_X1 U16277 ( .A1(n14161), .A2(n14160), .ZN(n14169) );
  OAI211_X1 U16278 ( .C1(n14161), .C2(n14160), .A(n14169), .B(n15752), .ZN(
        n14162) );
  NAND2_X1 U16279 ( .A1(n14163), .A2(n14162), .ZN(P2_U3231) );
  NAND2_X1 U16280 ( .A1(n15746), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n15745) );
  INV_X1 U16281 ( .A(n14165), .ZN(n14166) );
  INV_X1 U16282 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14552) );
  NAND2_X1 U16283 ( .A1(n14167), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n14168) );
  NAND2_X1 U16284 ( .A1(n14169), .A2(n14168), .ZN(n14171) );
  XNOR2_X1 U16285 ( .A(n14171), .B(n15748), .ZN(n15743) );
  NAND2_X1 U16286 ( .A1(n15743), .A2(n14345), .ZN(n14173) );
  OR2_X1 U16287 ( .A1(n14171), .A2(n14170), .ZN(n14172) );
  NAND2_X1 U16288 ( .A1(n14173), .A2(n14172), .ZN(n14174) );
  XNOR2_X1 U16289 ( .A(n14174), .B(n14327), .ZN(n14175) );
  OAI211_X1 U16290 ( .C1(n14616), .C2(n14186), .A(n15767), .B(n14178), .ZN(
        n14491) );
  NOR2_X1 U16291 ( .A1(n14616), .A2(n14436), .ZN(n14179) );
  AOI211_X1 U16292 ( .C1(n15783), .C2(P2_REG2_REG_30__SCAN_IN), .A(n14180), 
        .B(n14179), .ZN(n14181) );
  OAI21_X1 U16293 ( .B1(n14461), .B2(n14491), .A(n14181), .ZN(P2_U3235) );
  AOI21_X1 U16294 ( .B1(n14182), .B2(n14496), .A(n14499), .ZN(n14185) );
  XNOR2_X1 U16295 ( .A(n14185), .B(n14498), .ZN(n14200) );
  INV_X1 U16296 ( .A(n14505), .ZN(n14190) );
  AOI22_X1 U16297 ( .A1(n14188), .A2(n15762), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n15783), .ZN(n14189) );
  OAI21_X1 U16298 ( .B1(n14190), .B2(n14436), .A(n14189), .ZN(n14199) );
  XNOR2_X1 U16299 ( .A(n14193), .B(n14494), .ZN(n14198) );
  OAI22_X1 U16300 ( .A1(n14196), .A2(n14472), .B1(n14195), .B2(n14194), .ZN(
        n14197) );
  AOI21_X2 U16301 ( .B1(n14198), .B2(n15759), .A(n14197), .ZN(n14507) );
  AOI22_X1 U16302 ( .A1(n14203), .A2(n15762), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n15783), .ZN(n14204) );
  OAI21_X1 U16303 ( .B1(n14205), .B2(n14436), .A(n14204), .ZN(n14207) );
  INV_X1 U16304 ( .A(n14208), .ZN(n14213) );
  AOI22_X1 U16305 ( .A1(n14209), .A2(n15762), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n15783), .ZN(n14210) );
  OAI21_X1 U16306 ( .B1(n14511), .B2(n14436), .A(n14210), .ZN(n14212) );
  INV_X1 U16307 ( .A(n14514), .ZN(n14229) );
  INV_X1 U16308 ( .A(n14231), .ZN(n14216) );
  AOI211_X1 U16309 ( .C1(n14217), .C2(n14216), .A(n14481), .B(n14215), .ZN(
        n14513) );
  NOR2_X1 U16310 ( .A1(n14619), .A2(n14436), .ZN(n14221) );
  OAI22_X1 U16311 ( .A1(n14219), .A2(n15776), .B1(n14218), .B2(n15781), .ZN(
        n14220) );
  AOI211_X1 U16312 ( .C1(n14513), .C2(n15770), .A(n14221), .B(n14220), .ZN(
        n14228) );
  NOR2_X1 U16313 ( .A1(n14223), .A2(n14222), .ZN(n14225) );
  NAND2_X1 U16314 ( .A1(n14512), .A2(n15781), .ZN(n14227) );
  OAI211_X1 U16315 ( .C1(n14229), .C2(n14421), .A(n14228), .B(n14227), .ZN(
        P2_U3239) );
  XOR2_X1 U16316 ( .A(n14230), .B(n14235), .Z(n14520) );
  AOI211_X1 U16317 ( .C1(n14517), .C2(n14252), .A(n14481), .B(n14231), .ZN(
        n14516) );
  AOI22_X1 U16318 ( .A1(n14232), .A2(n15762), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n15783), .ZN(n14233) );
  OAI21_X1 U16319 ( .B1(n14234), .B2(n14436), .A(n14233), .ZN(n14240) );
  XNOR2_X1 U16320 ( .A(n14236), .B(n14235), .ZN(n14238) );
  AOI21_X1 U16321 ( .B1(n14238), .B2(n15759), .A(n14237), .ZN(n14519) );
  NOR2_X1 U16322 ( .A1(n14519), .A2(n15783), .ZN(n14239) );
  AOI211_X1 U16323 ( .C1(n14516), .C2(n15770), .A(n14240), .B(n14239), .ZN(
        n14241) );
  OAI21_X1 U16324 ( .B1(n14520), .B2(n14421), .A(n14241), .ZN(P2_U3240) );
  NAND2_X1 U16325 ( .A1(n14243), .A2(n14242), .ZN(n14245) );
  XNOR2_X1 U16326 ( .A(n14245), .B(n14244), .ZN(n14247) );
  AOI21_X1 U16327 ( .B1(n14247), .B2(n15759), .A(n14246), .ZN(n14524) );
  OAI21_X1 U16328 ( .B1(n14250), .B2(n14249), .A(n14248), .ZN(n14525) );
  INV_X1 U16329 ( .A(n14525), .ZN(n14259) );
  AOI21_X1 U16330 ( .B1(n14251), .B2(n14522), .A(n14481), .ZN(n14253) );
  AND2_X1 U16331 ( .A1(n14253), .A2(n14252), .ZN(n14521) );
  NAND2_X1 U16332 ( .A1(n14521), .A2(n15770), .ZN(n14256) );
  AOI22_X1 U16333 ( .A1(n14254), .A2(n15762), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n15783), .ZN(n14255) );
  OAI211_X1 U16334 ( .C1(n14257), .C2(n14436), .A(n14256), .B(n14255), .ZN(
        n14258) );
  AOI21_X1 U16335 ( .B1(n14259), .B2(n15771), .A(n14258), .ZN(n14260) );
  OAI21_X1 U16336 ( .B1(n15783), .B2(n14524), .A(n14260), .ZN(P2_U3241) );
  INV_X1 U16337 ( .A(n14261), .ZN(n14269) );
  OR2_X1 U16338 ( .A1(n14262), .A2(n14474), .ZN(n14265) );
  NAND2_X1 U16339 ( .A1(n14263), .A2(n14451), .ZN(n14264) );
  NAND2_X1 U16340 ( .A1(n14265), .A2(n14264), .ZN(n14527) );
  XNOR2_X1 U16341 ( .A(n14266), .B(n14270), .ZN(n14267) );
  NAND2_X1 U16342 ( .A1(n14267), .A2(n15759), .ZN(n14530) );
  INV_X1 U16343 ( .A(n14530), .ZN(n14268) );
  AOI211_X1 U16344 ( .C1(n15762), .C2(n14269), .A(n14527), .B(n14268), .ZN(
        n14277) );
  XNOR2_X1 U16345 ( .A(n14271), .B(n14270), .ZN(n14526) );
  OAI211_X1 U16346 ( .C1(n14283), .C2(n14273), .A(n15767), .B(n14251), .ZN(
        n14529) );
  NOR2_X1 U16347 ( .A1(n14529), .A2(n14461), .ZN(n14275) );
  OAI22_X1 U16348 ( .A1(n14273), .A2(n14436), .B1(n14272), .B2(n15781), .ZN(
        n14274) );
  AOI211_X1 U16349 ( .C1(n14526), .C2(n15771), .A(n14275), .B(n14274), .ZN(
        n14276) );
  OAI21_X1 U16350 ( .B1(n15783), .B2(n14277), .A(n14276), .ZN(P2_U3242) );
  XNOR2_X1 U16351 ( .A(n14278), .B(n14282), .ZN(n14280) );
  OAI21_X1 U16352 ( .B1(n14280), .B2(n14425), .A(n14279), .ZN(n14533) );
  INV_X1 U16353 ( .A(n14533), .ZN(n14290) );
  XOR2_X1 U16354 ( .A(n14282), .B(n14281), .Z(n14535) );
  AOI211_X1 U16355 ( .C1(n14284), .C2(n14294), .A(n14481), .B(n14283), .ZN(
        n14534) );
  NAND2_X1 U16356 ( .A1(n14534), .A2(n15770), .ZN(n14287) );
  AOI22_X1 U16357 ( .A1(n14285), .A2(n15762), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n15783), .ZN(n14286) );
  OAI211_X1 U16358 ( .C1(n14626), .C2(n14436), .A(n14287), .B(n14286), .ZN(
        n14288) );
  AOI21_X1 U16359 ( .B1(n14535), .B2(n15771), .A(n14288), .ZN(n14289) );
  OAI21_X1 U16360 ( .B1(n15783), .B2(n14290), .A(n14289), .ZN(P2_U3243) );
  XNOR2_X1 U16361 ( .A(n14291), .B(n14300), .ZN(n14293) );
  AOI21_X1 U16362 ( .B1(n14293), .B2(n15759), .A(n14292), .ZN(n14541) );
  AOI21_X1 U16363 ( .B1(n6563), .B2(n14539), .A(n14481), .ZN(n14295) );
  AND2_X1 U16364 ( .A1(n14295), .A2(n14294), .ZN(n14538) );
  INV_X1 U16365 ( .A(n14296), .ZN(n14297) );
  AOI22_X1 U16366 ( .A1(n14297), .A2(n15762), .B1(P2_REG2_REG_21__SCAN_IN), 
        .B2(n15783), .ZN(n14298) );
  OAI21_X1 U16367 ( .B1(n14299), .B2(n14436), .A(n14298), .ZN(n14303) );
  XOR2_X1 U16368 ( .A(n14301), .B(n14300), .Z(n14542) );
  NOR2_X1 U16369 ( .A1(n14542), .A2(n14421), .ZN(n14302) );
  AOI211_X1 U16370 ( .C1(n14538), .C2(n15770), .A(n14303), .B(n14302), .ZN(
        n14304) );
  OAI21_X1 U16371 ( .B1(n15783), .B2(n14541), .A(n14304), .ZN(P2_U3244) );
  XNOR2_X1 U16372 ( .A(n14305), .B(n14309), .ZN(n14307) );
  AOI21_X1 U16373 ( .B1(n14307), .B2(n15759), .A(n14306), .ZN(n14546) );
  OAI21_X1 U16374 ( .B1(n14310), .B2(n14309), .A(n14308), .ZN(n14547) );
  INV_X1 U16375 ( .A(n14547), .ZN(n14318) );
  AOI21_X1 U16376 ( .B1(n14325), .B2(n14544), .A(n14481), .ZN(n14312) );
  AND2_X1 U16377 ( .A1(n14312), .A2(n6563), .ZN(n14543) );
  NAND2_X1 U16378 ( .A1(n14543), .A2(n15770), .ZN(n14315) );
  AOI22_X1 U16379 ( .A1(n14313), .A2(n15762), .B1(n15783), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n14314) );
  OAI211_X1 U16380 ( .C1(n14316), .C2(n14436), .A(n14315), .B(n14314), .ZN(
        n14317) );
  AOI21_X1 U16381 ( .B1(n14318), .B2(n15771), .A(n14317), .ZN(n14319) );
  OAI21_X1 U16382 ( .B1(n15783), .B2(n14546), .A(n14319), .ZN(P2_U3245) );
  XOR2_X1 U16383 ( .A(n14320), .B(n14323), .Z(n14322) );
  AOI21_X1 U16384 ( .B1(n14322), .B2(n15759), .A(n14321), .ZN(n14549) );
  XNOR2_X1 U16385 ( .A(n14324), .B(n14323), .ZN(n14550) );
  NOR2_X1 U16386 ( .A1(n14550), .A2(n14421), .ZN(n14332) );
  OAI211_X1 U16387 ( .C1(n14632), .C2(n14348), .A(n15767), .B(n14325), .ZN(
        n14548) );
  OAI22_X1 U16388 ( .A1(n15781), .A2(n14327), .B1(n14326), .B2(n15776), .ZN(
        n14328) );
  AOI21_X1 U16389 ( .B1(n14329), .B2(n15763), .A(n14328), .ZN(n14330) );
  OAI21_X1 U16390 ( .B1(n14548), .B2(n14461), .A(n14330), .ZN(n14331) );
  NOR2_X1 U16391 ( .A1(n14332), .A2(n14331), .ZN(n14333) );
  OAI21_X1 U16392 ( .B1(n15783), .B2(n14549), .A(n14333), .ZN(P2_U3246) );
  NAND2_X1 U16393 ( .A1(n14335), .A2(n14338), .ZN(n14336) );
  NAND2_X1 U16394 ( .A1(n14334), .A2(n14336), .ZN(n14554) );
  INV_X1 U16395 ( .A(n14554), .ZN(n14354) );
  XNOR2_X1 U16396 ( .A(n14337), .B(n14338), .ZN(n14343) );
  NAND2_X1 U16397 ( .A1(n14554), .A2(n14446), .ZN(n14342) );
  AOI22_X1 U16398 ( .A1(n14340), .A2(n14449), .B1(n14339), .B2(n14451), .ZN(
        n14341) );
  OAI211_X1 U16399 ( .C1(n14425), .C2(n14343), .A(n14342), .B(n14341), .ZN(
        n14558) );
  NAND2_X1 U16400 ( .A1(n14558), .A2(n15781), .ZN(n14353) );
  OAI22_X1 U16401 ( .A1(n15781), .A2(n14345), .B1(n14344), .B2(n15776), .ZN(
        n14350) );
  NAND2_X1 U16402 ( .A1(n14362), .A2(n14351), .ZN(n14346) );
  NAND2_X1 U16403 ( .A1(n14346), .A2(n15767), .ZN(n14347) );
  OR2_X1 U16404 ( .A1(n14348), .A2(n14347), .ZN(n14555) );
  NOR2_X1 U16405 ( .A1(n14555), .A2(n14461), .ZN(n14349) );
  AOI211_X1 U16406 ( .C1(n15763), .C2(n14351), .A(n14350), .B(n14349), .ZN(
        n14352) );
  OAI211_X1 U16407 ( .C1(n14354), .C2(n14489), .A(n14353), .B(n14352), .ZN(
        P2_U3247) );
  NAND2_X1 U16408 ( .A1(n14385), .A2(n14355), .ZN(n14372) );
  OAI21_X1 U16409 ( .B1(n14372), .B2(n14374), .A(n7113), .ZN(n14357) );
  XNOR2_X1 U16410 ( .A(n14357), .B(n14359), .ZN(n14563) );
  INV_X1 U16411 ( .A(n14563), .ZN(n14371) );
  XNOR2_X1 U16412 ( .A(n14358), .B(n14359), .ZN(n14360) );
  OAI222_X1 U16413 ( .A1(n14474), .A2(n10517), .B1(n14472), .B2(n14361), .C1(
        n14360), .C2(n14425), .ZN(n14561) );
  INV_X1 U16414 ( .A(n14362), .ZN(n14363) );
  AOI211_X1 U16415 ( .C1(n14364), .C2(n14377), .A(n14481), .B(n14363), .ZN(
        n14562) );
  NAND2_X1 U16416 ( .A1(n14562), .A2(n15770), .ZN(n14368) );
  INV_X1 U16417 ( .A(n14365), .ZN(n14366) );
  AOI22_X1 U16418 ( .A1(n15783), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n14366), 
        .B2(n15762), .ZN(n14367) );
  OAI211_X1 U16419 ( .C1(n7662), .C2(n14436), .A(n14368), .B(n14367), .ZN(
        n14369) );
  AOI21_X1 U16420 ( .B1(n14561), .B2(n15781), .A(n14369), .ZN(n14370) );
  OAI21_X1 U16421 ( .B1(n14371), .B2(n14421), .A(n14370), .ZN(P2_U3248) );
  XNOR2_X1 U16422 ( .A(n14372), .B(n14374), .ZN(n14570) );
  XNOR2_X1 U16423 ( .A(n14373), .B(n14374), .ZN(n14375) );
  OAI222_X1 U16424 ( .A1(n14472), .A2(n14412), .B1(n14474), .B2(n14376), .C1(
        n14375), .C2(n14425), .ZN(n14566) );
  NAND2_X1 U16425 ( .A1(n14566), .A2(n15781), .ZN(n14384) );
  INV_X1 U16426 ( .A(n14377), .ZN(n14378) );
  AOI211_X1 U16427 ( .C1(n14568), .C2(n14390), .A(n14481), .B(n14378), .ZN(
        n14567) );
  NOR2_X1 U16428 ( .A1(n7663), .A2(n14436), .ZN(n14382) );
  OAI22_X1 U16429 ( .A1(n15781), .A2(n14380), .B1(n14379), .B2(n15776), .ZN(
        n14381) );
  AOI211_X1 U16430 ( .C1(n14567), .C2(n15770), .A(n14382), .B(n14381), .ZN(
        n14383) );
  OAI211_X1 U16431 ( .C1(n14570), .C2(n14421), .A(n14384), .B(n14383), .ZN(
        P2_U3249) );
  INV_X1 U16432 ( .A(n14385), .ZN(n14386) );
  AOI21_X1 U16433 ( .B1(n14394), .B2(n14387), .A(n14386), .ZN(n14577) );
  OAI22_X1 U16434 ( .A1(n15781), .A2(n14389), .B1(n14388), .B2(n15776), .ZN(
        n14392) );
  OAI211_X1 U16435 ( .C1(n14573), .C2(n14414), .A(n11714), .B(n14390), .ZN(
        n14572) );
  NOR2_X1 U16436 ( .A1(n14572), .A2(n14461), .ZN(n14391) );
  AOI211_X1 U16437 ( .C1(n15763), .C2(n14393), .A(n14392), .B(n14391), .ZN(
        n14401) );
  XNOR2_X1 U16438 ( .A(n14395), .B(n14394), .ZN(n14396) );
  NAND2_X1 U16439 ( .A1(n14396), .A2(n15759), .ZN(n14575) );
  AOI22_X1 U16440 ( .A1(n14398), .A2(n14449), .B1(n14451), .B2(n14397), .ZN(
        n14571) );
  AOI21_X1 U16441 ( .B1(n14575), .B2(n14571), .A(n15783), .ZN(n14399) );
  INV_X1 U16442 ( .A(n14399), .ZN(n14400) );
  OAI211_X1 U16443 ( .C1(n14577), .C2(n14421), .A(n14401), .B(n14400), .ZN(
        P2_U3250) );
  XNOR2_X1 U16444 ( .A(n14402), .B(n14409), .ZN(n14582) );
  INV_X1 U16445 ( .A(n14403), .ZN(n14471) );
  AOI21_X1 U16446 ( .B1(n14471), .B2(n14405), .A(n14404), .ZN(n14407) );
  NOR2_X1 U16447 ( .A1(n14407), .A2(n14406), .ZN(n14408) );
  XOR2_X1 U16448 ( .A(n14409), .B(n14408), .Z(n14410) );
  OAI222_X1 U16449 ( .A1(n14474), .A2(n14412), .B1(n14472), .B2(n14411), .C1(
        n14410), .C2(n14425), .ZN(n14578) );
  AOI211_X1 U16450 ( .C1(n14580), .C2(n14430), .A(n14481), .B(n14414), .ZN(
        n14579) );
  NAND2_X1 U16451 ( .A1(n14579), .A2(n15770), .ZN(n14417) );
  AOI22_X1 U16452 ( .A1(n15783), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n14415), 
        .B2(n15762), .ZN(n14416) );
  OAI211_X1 U16453 ( .C1(n14418), .C2(n14436), .A(n14417), .B(n14416), .ZN(
        n14419) );
  AOI21_X1 U16454 ( .B1(n14578), .B2(n15781), .A(n14419), .ZN(n14420) );
  OAI21_X1 U16455 ( .B1(n14421), .B2(n14582), .A(n14420), .ZN(P2_U3251) );
  NAND2_X1 U16456 ( .A1(n14469), .A2(n14422), .ZN(n14443) );
  NAND2_X1 U16457 ( .A1(n14445), .A2(n14423), .ZN(n14424) );
  XNOR2_X1 U16458 ( .A(n14424), .B(n14429), .ZN(n14426) );
  OAI222_X1 U16459 ( .A1(n14474), .A2(n14427), .B1(n14472), .B2(n14475), .C1(
        n14426), .C2(n14425), .ZN(n14583) );
  INV_X1 U16460 ( .A(n14583), .ZN(n14439) );
  XNOR2_X1 U16461 ( .A(n14428), .B(n14429), .ZN(n14585) );
  INV_X1 U16462 ( .A(n14460), .ZN(n14431) );
  AOI211_X1 U16463 ( .C1(n14432), .C2(n14431), .A(n14481), .B(n6765), .ZN(
        n14584) );
  NAND2_X1 U16464 ( .A1(n14584), .A2(n15770), .ZN(n14435) );
  AOI22_X1 U16465 ( .A1(n15783), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n14433), 
        .B2(n15762), .ZN(n14434) );
  OAI211_X1 U16466 ( .C1(n14645), .C2(n14436), .A(n14435), .B(n14434), .ZN(
        n14437) );
  AOI21_X1 U16467 ( .B1(n14585), .B2(n15771), .A(n14437), .ZN(n14438) );
  OAI21_X1 U16468 ( .B1(n14439), .B2(n15783), .A(n14438), .ZN(P2_U3252) );
  INV_X1 U16469 ( .A(n14442), .ZN(n14441) );
  XNOR2_X1 U16470 ( .A(n14440), .B(n14441), .ZN(n14447) );
  INV_X1 U16471 ( .A(n14447), .ZN(n14591) );
  NAND2_X1 U16472 ( .A1(n14443), .A2(n14442), .ZN(n14444) );
  NAND3_X1 U16473 ( .A1(n14445), .A2(n15759), .A3(n14444), .ZN(n14454) );
  NAND2_X1 U16474 ( .A1(n14447), .A2(n14446), .ZN(n14453) );
  AOI22_X1 U16475 ( .A1(n14451), .A2(n14450), .B1(n14449), .B2(n14448), .ZN(
        n14452) );
  NAND3_X1 U16476 ( .A1(n14454), .A2(n14453), .A3(n14452), .ZN(n14593) );
  NAND2_X1 U16477 ( .A1(n14593), .A2(n15781), .ZN(n14465) );
  OAI22_X1 U16478 ( .A1(n15781), .A2(n14456), .B1(n14455), .B2(n15776), .ZN(
        n14463) );
  OAI21_X1 U16479 ( .B1(n14457), .B2(n14458), .A(n15767), .ZN(n14459) );
  OR2_X1 U16480 ( .A1(n14460), .A2(n14459), .ZN(n14589) );
  NOR2_X1 U16481 ( .A1(n14589), .A2(n14461), .ZN(n14462) );
  AOI211_X1 U16482 ( .C1(n15763), .C2(n14588), .A(n14463), .B(n14462), .ZN(
        n14464) );
  OAI211_X1 U16483 ( .C1(n14591), .C2(n14489), .A(n14465), .B(n14464), .ZN(
        P2_U3253) );
  NAND2_X1 U16484 ( .A1(n14466), .A2(n14470), .ZN(n14467) );
  NAND2_X1 U16485 ( .A1(n14468), .A2(n14467), .ZN(n14596) );
  OAI21_X1 U16486 ( .B1(n14471), .B2(n14470), .A(n14469), .ZN(n14477) );
  OAI22_X1 U16487 ( .A1(n14475), .A2(n14474), .B1(n14473), .B2(n14472), .ZN(
        n14476) );
  AOI21_X1 U16488 ( .B1(n14477), .B2(n15759), .A(n14476), .ZN(n14478) );
  OAI21_X1 U16489 ( .B1(n14479), .B2(n14596), .A(n14478), .ZN(n14597) );
  NAND2_X1 U16490 ( .A1(n14597), .A2(n15781), .ZN(n14488) );
  INV_X1 U16491 ( .A(n14480), .ZN(n14482) );
  AOI211_X1 U16492 ( .C1(n14483), .C2(n14482), .A(n14481), .B(n14457), .ZN(
        n14598) );
  AOI22_X1 U16493 ( .A1(n15783), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n14484), 
        .B2(n15762), .ZN(n14485) );
  OAI21_X1 U16494 ( .B1(n14653), .B2(n14436), .A(n14485), .ZN(n14486) );
  AOI21_X1 U16495 ( .B1(n14598), .B2(n15770), .A(n14486), .ZN(n14487) );
  OAI211_X1 U16496 ( .C1(n14596), .C2(n14489), .A(n14488), .B(n14487), .ZN(
        P2_U3254) );
  INV_X1 U16497 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n14492) );
  MUX2_X1 U16498 ( .A(n14492), .B(n14613), .S(n15848), .Z(n14493) );
  OAI21_X1 U16499 ( .B1(n14616), .B2(n14602), .A(n14493), .ZN(P2_U3529) );
  NOR2_X1 U16500 ( .A1(n14496), .A2(n14499), .ZN(n14497) );
  AOI21_X1 U16501 ( .B1(n14498), .B2(n14497), .A(n15817), .ZN(n14501) );
  OAI211_X1 U16502 ( .C1(n14509), .C2(n14508), .A(n14507), .B(n14506), .ZN(
        n14617) );
  MUX2_X1 U16503 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n14617), .S(n15848), .Z(
        P2_U3528) );
  INV_X1 U16504 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n14515) );
  AOI21_X1 U16505 ( .B1(n15812), .B2(n14517), .A(n14516), .ZN(n14518) );
  OAI211_X1 U16506 ( .C1(n14520), .C2(n15817), .A(n14519), .B(n14518), .ZN(
        n14620) );
  MUX2_X1 U16507 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14620), .S(n15848), .Z(
        P2_U3524) );
  AOI21_X1 U16508 ( .B1(n15812), .B2(n14522), .A(n14521), .ZN(n14523) );
  OAI211_X1 U16509 ( .C1(n14525), .C2(n15817), .A(n14524), .B(n14523), .ZN(
        n14621) );
  MUX2_X1 U16510 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14621), .S(n15848), .Z(
        P2_U3523) );
  NAND2_X1 U16511 ( .A1(n14526), .A2(n15835), .ZN(n14532) );
  AOI21_X1 U16512 ( .B1(n14528), .B2(n15812), .A(n14527), .ZN(n14531) );
  NAND4_X1 U16513 ( .A1(n14532), .A2(n14531), .A3(n14530), .A4(n14529), .ZN(
        n14622) );
  MUX2_X1 U16514 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14622), .S(n15848), .Z(
        P2_U3522) );
  INV_X1 U16515 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n14536) );
  AOI211_X1 U16516 ( .C1(n14535), .C2(n15835), .A(n14534), .B(n14533), .ZN(
        n14623) );
  MUX2_X1 U16517 ( .A(n14536), .B(n14623), .S(n15848), .Z(n14537) );
  OAI21_X1 U16518 ( .B1(n14626), .B2(n14602), .A(n14537), .ZN(P2_U3521) );
  AOI21_X1 U16519 ( .B1(n15812), .B2(n14539), .A(n14538), .ZN(n14540) );
  OAI211_X1 U16520 ( .C1(n14542), .C2(n15817), .A(n14541), .B(n14540), .ZN(
        n14627) );
  MUX2_X1 U16521 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14627), .S(n15848), .Z(
        P2_U3520) );
  AOI21_X1 U16522 ( .B1(n15812), .B2(n14544), .A(n14543), .ZN(n14545) );
  OAI211_X1 U16523 ( .C1(n14547), .C2(n15817), .A(n14546), .B(n14545), .ZN(
        n14628) );
  MUX2_X1 U16524 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14628), .S(n15848), .Z(
        P2_U3519) );
  OAI211_X1 U16525 ( .C1(n14550), .C2(n15817), .A(n14549), .B(n14548), .ZN(
        n14551) );
  INV_X1 U16526 ( .A(n14551), .ZN(n14629) );
  MUX2_X1 U16527 ( .A(n14552), .B(n14629), .S(n15848), .Z(n14553) );
  OAI21_X1 U16528 ( .B1(n14632), .B2(n14602), .A(n14553), .ZN(P2_U3518) );
  INV_X1 U16529 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14559) );
  NAND2_X1 U16530 ( .A1(n14554), .A2(n15810), .ZN(n14556) );
  OAI211_X1 U16531 ( .C1(n10518), .C2(n15831), .A(n14556), .B(n14555), .ZN(
        n14557) );
  NOR2_X1 U16532 ( .A1(n14558), .A2(n14557), .ZN(n14633) );
  MUX2_X1 U16533 ( .A(n14559), .B(n14633), .S(n15848), .Z(n14560) );
  INV_X1 U16534 ( .A(n14560), .ZN(P2_U3517) );
  AOI211_X1 U16535 ( .C1(n15835), .C2(n14563), .A(n14562), .B(n14561), .ZN(
        n14636) );
  MUX2_X1 U16536 ( .A(n14564), .B(n14636), .S(n15848), .Z(n14565) );
  OAI21_X1 U16537 ( .B1(n7662), .B2(n14602), .A(n14565), .ZN(P2_U3516) );
  AOI211_X1 U16538 ( .C1(n15812), .C2(n14568), .A(n14567), .B(n14566), .ZN(
        n14569) );
  OAI21_X1 U16539 ( .B1(n15817), .B2(n14570), .A(n14569), .ZN(n14639) );
  MUX2_X1 U16540 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14639), .S(n15848), .Z(
        P2_U3515) );
  OAI211_X1 U16541 ( .C1(n14573), .C2(n15831), .A(n14572), .B(n14571), .ZN(
        n14574) );
  INV_X1 U16542 ( .A(n14574), .ZN(n14576) );
  OAI211_X1 U16543 ( .C1(n14577), .C2(n15817), .A(n14576), .B(n14575), .ZN(
        n14640) );
  MUX2_X1 U16544 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n14640), .S(n15848), .Z(
        P2_U3514) );
  AOI211_X1 U16545 ( .C1(n15812), .C2(n14580), .A(n14579), .B(n14578), .ZN(
        n14581) );
  OAI21_X1 U16546 ( .B1(n15817), .B2(n14582), .A(n14581), .ZN(n14641) );
  MUX2_X1 U16547 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n14641), .S(n15848), .Z(
        P2_U3513) );
  INV_X1 U16548 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n14586) );
  AOI211_X1 U16549 ( .C1(n15835), .C2(n14585), .A(n14584), .B(n14583), .ZN(
        n14642) );
  MUX2_X1 U16550 ( .A(n14586), .B(n14642), .S(n15848), .Z(n14587) );
  OAI21_X1 U16551 ( .B1(n14645), .B2(n14602), .A(n14587), .ZN(P2_U3512) );
  INV_X1 U16552 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14594) );
  NAND2_X1 U16553 ( .A1(n14588), .A2(n15812), .ZN(n14590) );
  OAI211_X1 U16554 ( .C1(n14591), .C2(n13811), .A(n14590), .B(n14589), .ZN(
        n14592) );
  NOR2_X1 U16555 ( .A1(n14593), .A2(n14592), .ZN(n14646) );
  MUX2_X1 U16556 ( .A(n14594), .B(n14646), .S(n15848), .Z(n14595) );
  INV_X1 U16557 ( .A(n14595), .ZN(P2_U3511) );
  INV_X1 U16558 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n14600) );
  INV_X1 U16559 ( .A(n14596), .ZN(n14599) );
  AOI211_X1 U16560 ( .C1(n14599), .C2(n15810), .A(n14598), .B(n14597), .ZN(
        n14649) );
  MUX2_X1 U16561 ( .A(n14600), .B(n14649), .S(n15848), .Z(n14601) );
  OAI21_X1 U16562 ( .B1(n14653), .B2(n14602), .A(n14601), .ZN(P2_U3510) );
  INV_X1 U16563 ( .A(n14603), .ZN(n14608) );
  AOI21_X1 U16564 ( .B1(n15812), .B2(n14605), .A(n14604), .ZN(n14606) );
  OAI211_X1 U16565 ( .C1(n14608), .C2(n13811), .A(n14607), .B(n14606), .ZN(
        n14654) );
  MUX2_X1 U16566 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n14654), .S(n15848), .Z(
        P2_U3509) );
  AOI21_X1 U16567 ( .B1(n15812), .B2(n7205), .A(n14609), .ZN(n14610) );
  OAI211_X1 U16568 ( .C1(n13811), .C2(n14612), .A(n14611), .B(n14610), .ZN(
        n14655) );
  MUX2_X1 U16569 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n14655), .S(n15848), .Z(
        P2_U3507) );
  INV_X1 U16570 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n14614) );
  MUX2_X1 U16571 ( .A(n14614), .B(n14613), .S(n15838), .Z(n14615) );
  OAI21_X1 U16572 ( .B1(n14616), .B2(n14652), .A(n14615), .ZN(P2_U3497) );
  MUX2_X1 U16573 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n14617), .S(n15838), .Z(
        P2_U3496) );
  MUX2_X1 U16574 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14620), .S(n15838), .Z(
        P2_U3492) );
  MUX2_X1 U16575 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14621), .S(n15838), .Z(
        P2_U3491) );
  MUX2_X1 U16576 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14622), .S(n15838), .Z(
        P2_U3490) );
  INV_X1 U16577 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n14624) );
  MUX2_X1 U16578 ( .A(n14624), .B(n14623), .S(n15838), .Z(n14625) );
  OAI21_X1 U16579 ( .B1(n14626), .B2(n14652), .A(n14625), .ZN(P2_U3489) );
  MUX2_X1 U16580 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14627), .S(n15838), .Z(
        P2_U3488) );
  MUX2_X1 U16581 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14628), .S(n15838), .Z(
        P2_U3487) );
  INV_X1 U16582 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14630) );
  MUX2_X1 U16583 ( .A(n14630), .B(n14629), .S(n15838), .Z(n14631) );
  OAI21_X1 U16584 ( .B1(n14632), .B2(n14652), .A(n14631), .ZN(P2_U3486) );
  INV_X1 U16585 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n14634) );
  MUX2_X1 U16586 ( .A(n14634), .B(n14633), .S(n15838), .Z(n14635) );
  INV_X1 U16587 ( .A(n14635), .ZN(P2_U3484) );
  MUX2_X1 U16588 ( .A(n14637), .B(n14636), .S(n15838), .Z(n14638) );
  OAI21_X1 U16589 ( .B1(n7662), .B2(n14652), .A(n14638), .ZN(P2_U3481) );
  MUX2_X1 U16590 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14639), .S(n15838), .Z(
        P2_U3478) );
  MUX2_X1 U16591 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n14640), .S(n15838), .Z(
        P2_U3475) );
  MUX2_X1 U16592 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n14641), .S(n15838), .Z(
        P2_U3472) );
  INV_X1 U16593 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14643) );
  MUX2_X1 U16594 ( .A(n14643), .B(n14642), .S(n15838), .Z(n14644) );
  OAI21_X1 U16595 ( .B1(n14645), .B2(n14652), .A(n14644), .ZN(P2_U3469) );
  INV_X1 U16596 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14647) );
  MUX2_X1 U16597 ( .A(n14647), .B(n14646), .S(n15838), .Z(n14648) );
  INV_X1 U16598 ( .A(n14648), .ZN(P2_U3466) );
  INV_X1 U16599 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n14650) );
  MUX2_X1 U16600 ( .A(n14650), .B(n14649), .S(n15838), .Z(n14651) );
  OAI21_X1 U16601 ( .B1(n14653), .B2(n14652), .A(n14651), .ZN(P2_U3463) );
  MUX2_X1 U16602 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n14654), .S(n15838), .Z(
        P2_U3460) );
  MUX2_X1 U16603 ( .A(P2_REG0_REG_8__SCAN_IN), .B(n14655), .S(n15838), .Z(
        P2_U3454) );
  INV_X1 U16604 ( .A(n14656), .ZN(n15426) );
  NAND3_X1 U16605 ( .A1(n14657), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n14659) );
  OAI22_X1 U16606 ( .A1(n14660), .A2(n14659), .B1(n14658), .B2(n14671), .ZN(
        n14661) );
  INV_X1 U16607 ( .A(n14661), .ZN(n14662) );
  OAI21_X1 U16608 ( .B1(n15426), .B2(n14663), .A(n14662), .ZN(P2_U3296) );
  NAND2_X1 U16609 ( .A1(n10297), .A2(n14664), .ZN(n14666) );
  OAI211_X1 U16610 ( .C1(n14667), .C2(n14671), .A(n14666), .B(n14665), .ZN(
        P2_U3299) );
  INV_X1 U16611 ( .A(n14668), .ZN(n15434) );
  OAI222_X1 U16612 ( .A1(n14671), .A2(n14670), .B1(n14673), .B2(n15434), .C1(
        n14669), .C2(n11242), .ZN(P2_U3300) );
  OAI222_X1 U16613 ( .A1(n6510), .A2(n14674), .B1(n14673), .B2(n15437), .C1(
        n14672), .C2(n14671), .ZN(P2_U3301) );
  MUX2_X1 U16614 ( .A(n14675), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XNOR2_X1 U16615 ( .A(n14677), .B(n14676), .ZN(n14726) );
  NAND2_X1 U16616 ( .A1(n14725), .A2(n14726), .ZN(n14783) );
  INV_X1 U16617 ( .A(n14678), .ZN(n14679) );
  XNOR2_X1 U16618 ( .A(n14680), .B(n14679), .ZN(n14781) );
  NAND3_X1 U16619 ( .A1(n14783), .A2(n14781), .A3(n14782), .ZN(n14780) );
  NAND2_X1 U16620 ( .A1(n14780), .A2(n14681), .ZN(n14685) );
  XNOR2_X1 U16621 ( .A(n14683), .B(n14682), .ZN(n14684) );
  XNOR2_X1 U16622 ( .A(n14685), .B(n14684), .ZN(n14690) );
  OAI21_X1 U16623 ( .B1(n15508), .B2(n15229), .A(n14686), .ZN(n14688) );
  OAI22_X1 U16624 ( .A1(n14826), .A2(n15228), .B1(n15226), .B2(n14825), .ZN(
        n14687) );
  AOI211_X1 U16625 ( .C1(n8965), .C2(n14830), .A(n14688), .B(n14687), .ZN(
        n14689) );
  OAI21_X1 U16626 ( .B1(n14690), .B2(n15496), .A(n14689), .ZN(P1_U3215) );
  INV_X1 U16627 ( .A(n14763), .ZN(n14694) );
  NOR3_X1 U16628 ( .A1(n14796), .A2(n14692), .A3(n14691), .ZN(n14693) );
  OAI21_X1 U16629 ( .B1(n14694), .B2(n14693), .A(n14813), .ZN(n14698) );
  INV_X1 U16630 ( .A(n15031), .ZN(n14739) );
  OAI22_X1 U16631 ( .A1(n14739), .A2(n15227), .B1(n15099), .B2(n15225), .ZN(
        n15306) );
  OAI22_X1 U16632 ( .A1(n15068), .A2(n15508), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14695), .ZN(n14696) );
  AOI21_X1 U16633 ( .B1(n15306), .B2(n15500), .A(n14696), .ZN(n14697) );
  OAI211_X1 U16634 ( .C1(n15309), .C2(n15503), .A(n14698), .B(n14697), .ZN(
        P1_U3216) );
  OAI211_X1 U16635 ( .C1(n14701), .C2(n14700), .A(n14699), .B(n14813), .ZN(
        n14706) );
  INV_X1 U16636 ( .A(n14702), .ZN(n15144) );
  OAI22_X1 U16637 ( .A1(n14826), .A2(n15098), .B1(n15177), .B2(n14825), .ZN(
        n14703) );
  AOI211_X1 U16638 ( .C1(n14829), .C2(n15144), .A(n14704), .B(n14703), .ZN(
        n14705) );
  OAI211_X1 U16639 ( .C1(n7851), .C2(n15503), .A(n14706), .B(n14705), .ZN(
        P1_U3219) );
  AOI22_X1 U16640 ( .A1(n14707), .A2(n14856), .B1(n14773), .B2(n14855), .ZN(
        n14716) );
  AOI22_X1 U16641 ( .A1(n14830), .A2(n14709), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n14708), .ZN(n14715) );
  OAI21_X1 U16642 ( .B1(n14712), .B2(n14711), .A(n14710), .ZN(n14713) );
  NAND2_X1 U16643 ( .A1(n14713), .A2(n14813), .ZN(n14714) );
  NAND3_X1 U16644 ( .A1(n14716), .A2(n14715), .A3(n14714), .ZN(P1_U3222) );
  OAI21_X1 U16645 ( .B1(n14718), .B2(n14717), .A(n14794), .ZN(n14719) );
  NAND2_X1 U16646 ( .A1(n14719), .A2(n14813), .ZN(n14723) );
  NOR2_X1 U16647 ( .A1(n15104), .A2(n15508), .ZN(n14721) );
  OAI22_X1 U16648 ( .A1(n15099), .A2(n14826), .B1(n15098), .B2(n14825), .ZN(
        n14720) );
  AOI211_X1 U16649 ( .C1(P1_REG3_REG_21__SCAN_IN), .C2(P1_U3086), .A(n14721), 
        .B(n14720), .ZN(n14722) );
  OAI211_X1 U16650 ( .C1(n15107), .C2(n15503), .A(n14723), .B(n14722), .ZN(
        P1_U3223) );
  OAI21_X1 U16651 ( .B1(n14726), .B2(n14725), .A(n14783), .ZN(n14727) );
  NAND2_X1 U16652 ( .A1(n14727), .A2(n14813), .ZN(n14734) );
  INV_X1 U16653 ( .A(n14728), .ZN(n14732) );
  OAI22_X1 U16654 ( .A1(n14826), .A2(n15226), .B1(n14729), .B2(n14825), .ZN(
        n14730) );
  AOI211_X1 U16655 ( .C1(n14829), .C2(n14732), .A(n14731), .B(n14730), .ZN(
        n14733) );
  OAI211_X1 U16656 ( .C1(n7847), .C2(n15503), .A(n14734), .B(n14733), .ZN(
        P1_U3224) );
  INV_X1 U16657 ( .A(n15030), .ZN(n15296) );
  NOR3_X1 U16658 ( .A1(n14765), .A2(n14736), .A3(n14735), .ZN(n14737) );
  OAI21_X1 U16659 ( .B1(n6619), .B2(n14737), .A(n14813), .ZN(n14743) );
  OAI22_X1 U16660 ( .A1(n15033), .A2(n15508), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14738), .ZN(n14741) );
  NOR2_X1 U16661 ( .A1(n14739), .A2(n14825), .ZN(n14740) );
  AOI211_X1 U16662 ( .C1(n14773), .C2(n15032), .A(n14741), .B(n14740), .ZN(
        n14742) );
  OAI211_X1 U16663 ( .C1(n15296), .C2(n15503), .A(n14743), .B(n14742), .ZN(
        P1_U3225) );
  NAND2_X1 U16664 ( .A1(n6567), .A2(n14744), .ZN(n14745) );
  OAI21_X1 U16665 ( .B1(n6567), .B2(n14744), .A(n14745), .ZN(n14823) );
  NOR2_X1 U16666 ( .A1(n14823), .A2(n14824), .ZN(n14822) );
  INV_X1 U16667 ( .A(n14745), .ZN(n14746) );
  NOR3_X1 U16668 ( .A1(n14822), .A2(n6587), .A3(n14746), .ZN(n14748) );
  INV_X1 U16669 ( .A(n14755), .ZN(n14747) );
  OAI21_X1 U16670 ( .B1(n14748), .B2(n14747), .A(n14813), .ZN(n14753) );
  INV_X1 U16671 ( .A(n14749), .ZN(n15197) );
  OAI22_X1 U16672 ( .A1(n14826), .A2(n15196), .B1(n15228), .B2(n14825), .ZN(
        n14750) );
  AOI211_X1 U16673 ( .C1(n14829), .C2(n15197), .A(n14751), .B(n14750), .ZN(
        n14752) );
  OAI211_X1 U16674 ( .C1(n8968), .C2(n15503), .A(n14753), .B(n14752), .ZN(
        P1_U3226) );
  AND3_X1 U16675 ( .A1(n14755), .A2(n7329), .A3(n14754), .ZN(n14756) );
  OAI21_X1 U16676 ( .B1(n14757), .B2(n14756), .A(n14813), .ZN(n14761) );
  INV_X1 U16677 ( .A(n14758), .ZN(n15181) );
  AND2_X1 U16678 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14946) );
  OAI22_X1 U16679 ( .A1(n14826), .A2(n15177), .B1(n15214), .B2(n14825), .ZN(
        n14759) );
  AOI211_X1 U16680 ( .C1(n14829), .C2(n15181), .A(n14946), .B(n14759), .ZN(
        n14760) );
  OAI211_X1 U16681 ( .C1(n15183), .C2(n15503), .A(n14761), .B(n14760), .ZN(
        P1_U3228) );
  AND3_X1 U16682 ( .A1(n14763), .A2(n14762), .A3(n7743), .ZN(n14764) );
  OAI21_X1 U16683 ( .B1(n14765), .B2(n14764), .A(n14813), .ZN(n14770) );
  OAI22_X1 U16684 ( .A1(n14815), .A2(n15227), .B1(n14766), .B2(n15225), .ZN(
        n15048) );
  OAI22_X1 U16685 ( .A1(n15056), .A2(n15508), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14767), .ZN(n14768) );
  AOI21_X1 U16686 ( .B1(n15048), .B2(n15500), .A(n14768), .ZN(n14769) );
  OAI211_X1 U16687 ( .C1(n7858), .C2(n15503), .A(n14770), .B(n14769), .ZN(
        P1_U3229) );
  XNOR2_X1 U16688 ( .A(n14772), .B(n14771), .ZN(n14779) );
  NAND2_X1 U16689 ( .A1(n15117), .A2(n14773), .ZN(n14775) );
  AOI22_X1 U16690 ( .A1(n14829), .A2(n15125), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14774) );
  OAI211_X1 U16691 ( .C1(n14776), .C2(n14825), .A(n14775), .B(n14774), .ZN(
        n14777) );
  AOI21_X1 U16692 ( .B1(n15324), .B2(n14830), .A(n14777), .ZN(n14778) );
  OAI21_X1 U16693 ( .B1(n14779), .B2(n15496), .A(n14778), .ZN(P1_U3233) );
  NAND2_X1 U16694 ( .A1(n14780), .A2(n14813), .ZN(n14791) );
  AOI21_X1 U16695 ( .B1(n14783), .B2(n14782), .A(n14781), .ZN(n14790) );
  OAI21_X1 U16696 ( .B1(n15508), .B2(n15260), .A(n14784), .ZN(n14787) );
  OAI22_X1 U16697 ( .A1(n14826), .A2(n15213), .B1(n14785), .B2(n14825), .ZN(
        n14786) );
  AOI211_X1 U16698 ( .C1(n14788), .C2(n14830), .A(n14787), .B(n14786), .ZN(
        n14789) );
  OAI21_X1 U16699 ( .B1(n14791), .B2(n14790), .A(n14789), .ZN(P1_U3234) );
  AND3_X1 U16700 ( .A1(n14794), .A2(n14793), .A3(n14792), .ZN(n14795) );
  OAI21_X1 U16701 ( .B1(n14796), .B2(n14795), .A(n14813), .ZN(n14801) );
  AND2_X1 U16702 ( .A1(n15117), .A2(n15257), .ZN(n14797) );
  AOI21_X1 U16703 ( .B1(n14839), .B2(n15256), .A(n14797), .ZN(n15084) );
  INV_X1 U16704 ( .A(n15500), .ZN(n14806) );
  OAI22_X1 U16705 ( .A1(n15084), .A2(n14806), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14798), .ZN(n14799) );
  AOI21_X1 U16706 ( .B1(n15088), .B2(n14829), .A(n14799), .ZN(n14800) );
  OAI211_X1 U16707 ( .C1(n15503), .C2(n15090), .A(n14801), .B(n14800), .ZN(
        P1_U3235) );
  AOI21_X1 U16708 ( .B1(n14804), .B2(n14803), .A(n14802), .ZN(n14809) );
  AOI22_X1 U16709 ( .A1(n15116), .A2(n15256), .B1(n15257), .B2(n14841), .ZN(
        n15156) );
  NAND2_X1 U16710 ( .A1(n14829), .A2(n15162), .ZN(n14805) );
  NAND2_X1 U16711 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14957)
         );
  OAI211_X1 U16712 ( .C1(n15156), .C2(n14806), .A(n14805), .B(n14957), .ZN(
        n14807) );
  AOI21_X1 U16713 ( .B1(n15339), .B2(n14830), .A(n14807), .ZN(n14808) );
  OAI21_X1 U16714 ( .B1(n14809), .B2(n15496), .A(n14808), .ZN(P1_U3238) );
  OAI21_X1 U16715 ( .B1(n14812), .B2(n14811), .A(n14810), .ZN(n14814) );
  NAND2_X1 U16716 ( .A1(n14814), .A2(n14813), .ZN(n14821) );
  OAI22_X1 U16717 ( .A1(n14816), .A2(n15227), .B1(n14815), .B2(n15225), .ZN(
        n15023) );
  INV_X1 U16718 ( .A(n15018), .ZN(n14818) );
  OAI22_X1 U16719 ( .A1(n14818), .A2(n15508), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14817), .ZN(n14819) );
  AOI21_X1 U16720 ( .B1(n15023), .B2(n15500), .A(n14819), .ZN(n14820) );
  OAI211_X1 U16721 ( .C1(n15020), .C2(n15503), .A(n14821), .B(n14820), .ZN(
        P1_U3240) );
  AOI21_X1 U16722 ( .B1(n14824), .B2(n14823), .A(n14822), .ZN(n14833) );
  OAI22_X1 U16723 ( .A1(n14826), .A2(n15214), .B1(n15213), .B2(n14825), .ZN(
        n14827) );
  AOI211_X1 U16724 ( .C1(n14829), .C2(n15215), .A(n14828), .B(n14827), .ZN(
        n14832) );
  NAND2_X1 U16725 ( .A1(n8898), .A2(n14830), .ZN(n14831) );
  OAI211_X1 U16726 ( .C1(n14833), .C2(n15496), .A(n14832), .B(n14831), .ZN(
        P1_U3241) );
  MUX2_X1 U16727 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14834), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16728 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14835), .S(P1_U4016), .Z(
        P1_U3589) );
  INV_X2 U16729 ( .A(n14836), .ZN(P1_U4016) );
  MUX2_X1 U16730 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14982), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16731 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14837), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16732 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n15032), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16733 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14838), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16734 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n15031), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16735 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14839), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16736 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14840), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16737 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n15117), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16738 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n15139), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16739 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n15116), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16740 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n15140), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16741 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14841), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16742 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14842), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16743 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14843), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16744 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n15255), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16745 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14844), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16746 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n15258), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16747 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14845), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16748 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14846), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16749 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14847), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16750 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14848), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16751 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14849), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16752 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14851), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16753 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14852), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16754 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14853), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16755 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14854), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16756 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14855), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16757 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14856), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI22_X1 U16758 ( .A1(n14959), .A2(n6748), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14857), .ZN(n14858) );
  AOI21_X1 U16759 ( .B1(n14962), .B2(n14859), .A(n14858), .ZN(n14867) );
  OAI211_X1 U16760 ( .C1(n14862), .C2(n14861), .A(n14954), .B(n14860), .ZN(
        n14866) );
  OAI211_X1 U16761 ( .C1(n14864), .C2(n14868), .A(n14965), .B(n14863), .ZN(
        n14865) );
  NAND3_X1 U16762 ( .A1(n14867), .A2(n14866), .A3(n14865), .ZN(P1_U3244) );
  INV_X1 U16763 ( .A(n14868), .ZN(n14869) );
  MUX2_X1 U16764 ( .A(n14870), .B(n14869), .S(n14971), .Z(n14875) );
  NAND2_X1 U16765 ( .A1(n14872), .A2(n14871), .ZN(n14873) );
  OAI211_X1 U16766 ( .C1(n14875), .C2(n14874), .A(P1_U4016), .B(n14873), .ZN(
        n14914) );
  INV_X1 U16767 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14877) );
  OAI22_X1 U16768 ( .A1(n14959), .A2(n14877), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14876), .ZN(n14878) );
  AOI21_X1 U16769 ( .B1(n14962), .B2(n14879), .A(n14878), .ZN(n14888) );
  OAI211_X1 U16770 ( .C1(n14882), .C2(n14881), .A(n14965), .B(n14880), .ZN(
        n14887) );
  OAI211_X1 U16771 ( .C1(n14885), .C2(n14884), .A(n14954), .B(n14883), .ZN(
        n14886) );
  NAND4_X1 U16772 ( .A1(n14914), .A2(n14888), .A3(n14887), .A4(n14886), .ZN(
        P1_U3245) );
  INV_X1 U16773 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14890) );
  NAND2_X1 U16774 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n14889) );
  OAI21_X1 U16775 ( .B1(n14959), .B2(n14890), .A(n14889), .ZN(n14891) );
  AOI21_X1 U16776 ( .B1(n14962), .B2(n14892), .A(n14891), .ZN(n14901) );
  OAI211_X1 U16777 ( .C1(n14895), .C2(n14894), .A(n14965), .B(n14893), .ZN(
        n14900) );
  OAI211_X1 U16778 ( .C1(n14898), .C2(n14897), .A(n14954), .B(n14896), .ZN(
        n14899) );
  NAND3_X1 U16779 ( .A1(n14901), .A2(n14900), .A3(n14899), .ZN(P1_U3246) );
  OAI21_X1 U16780 ( .B1(n14959), .B2(n9727), .A(n14902), .ZN(n14903) );
  AOI21_X1 U16781 ( .B1(n14962), .B2(n14904), .A(n14903), .ZN(n14913) );
  OAI211_X1 U16782 ( .C1(n14907), .C2(n14906), .A(n14954), .B(n14905), .ZN(
        n14912) );
  OAI211_X1 U16783 ( .C1(n14910), .C2(n14909), .A(n14965), .B(n14908), .ZN(
        n14911) );
  NAND4_X1 U16784 ( .A1(n14914), .A2(n14913), .A3(n14912), .A4(n14911), .ZN(
        P1_U3247) );
  NAND2_X1 U16785 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n14915) );
  OAI21_X1 U16786 ( .B1(n14959), .B2(n14916), .A(n14915), .ZN(n14917) );
  AOI21_X1 U16787 ( .B1(n14962), .B2(n14918), .A(n14917), .ZN(n14927) );
  OAI211_X1 U16788 ( .C1(n14921), .C2(n14920), .A(n14954), .B(n14919), .ZN(
        n14926) );
  OAI211_X1 U16789 ( .C1(n14924), .C2(n14923), .A(n14965), .B(n14922), .ZN(
        n14925) );
  NAND3_X1 U16790 ( .A1(n14927), .A2(n14926), .A3(n14925), .ZN(P1_U3250) );
  OAI211_X1 U16791 ( .C1(n14930), .C2(n14929), .A(n14928), .B(n14954), .ZN(
        n14940) );
  OAI21_X1 U16792 ( .B1(n14959), .B2(n14932), .A(n14931), .ZN(n14933) );
  AOI21_X1 U16793 ( .B1(n14962), .B2(n14934), .A(n14933), .ZN(n14939) );
  OAI211_X1 U16794 ( .C1(n14937), .C2(n14936), .A(n14935), .B(n14965), .ZN(
        n14938) );
  NAND3_X1 U16795 ( .A1(n14940), .A2(n14939), .A3(n14938), .ZN(P1_U3253) );
  OAI211_X1 U16796 ( .C1(n14943), .C2(n14942), .A(n14941), .B(n14954), .ZN(
        n14953) );
  NOR2_X1 U16797 ( .A1(n14959), .A2(n14944), .ZN(n14945) );
  AOI211_X1 U16798 ( .C1(n14962), .C2(n14947), .A(n14946), .B(n14945), .ZN(
        n14952) );
  OAI211_X1 U16799 ( .C1(n14950), .C2(n14949), .A(n14948), .B(n14965), .ZN(
        n14951) );
  NAND3_X1 U16800 ( .A1(n14953), .A2(n14952), .A3(n14951), .ZN(P1_U3260) );
  OAI211_X1 U16801 ( .C1(n14956), .C2(P1_REG1_REG_18__SCAN_IN), .A(n14955), 
        .B(n14954), .ZN(n14969) );
  OAI21_X1 U16802 ( .B1(n14959), .B2(n14958), .A(n14957), .ZN(n14960) );
  AOI21_X1 U16803 ( .B1(n14962), .B2(n14961), .A(n14960), .ZN(n14968) );
  INV_X1 U16804 ( .A(n14963), .ZN(n14966) );
  OAI211_X1 U16805 ( .C1(n14966), .C2(P1_REG2_REG_18__SCAN_IN), .A(n14965), 
        .B(n14964), .ZN(n14967) );
  NAND3_X1 U16806 ( .A1(n14969), .A2(n14968), .A3(n14967), .ZN(P1_U3261) );
  NAND2_X1 U16807 ( .A1(n15274), .A2(n15001), .ZN(n14970) );
  XNOR2_X1 U16808 ( .A(n14970), .B(n15269), .ZN(n15271) );
  NAND2_X1 U16809 ( .A1(n14971), .A2(P1_B_REG_SCAN_IN), .ZN(n14972) );
  NAND2_X1 U16810 ( .A1(n15256), .A2(n14972), .ZN(n15007) );
  NOR2_X1 U16811 ( .A1(n14973), .A2(n15007), .ZN(n15268) );
  INV_X1 U16812 ( .A(n15268), .ZN(n15272) );
  NOR2_X1 U16813 ( .A1(n15262), .A2(n15272), .ZN(n14980) );
  NOR2_X1 U16814 ( .A1(n14974), .A2(n15517), .ZN(n14975) );
  AOI211_X1 U16815 ( .C1(n15262), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14980), 
        .B(n14975), .ZN(n14976) );
  OAI21_X1 U16816 ( .B1(n15271), .B2(n15236), .A(n14976), .ZN(P1_U3263) );
  XNOR2_X1 U16817 ( .A(n15001), .B(n14977), .ZN(n14978) );
  NAND2_X1 U16818 ( .A1(n14978), .A2(n15555), .ZN(n15273) );
  NOR2_X1 U16819 ( .A1(n15274), .A2(n15517), .ZN(n14979) );
  AOI211_X1 U16820 ( .C1(n15262), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14980), 
        .B(n14979), .ZN(n14981) );
  OAI21_X1 U16821 ( .B1(n15067), .B2(n15273), .A(n14981), .ZN(P1_U3264) );
  NOR2_X1 U16822 ( .A1(n14983), .A2(n14982), .ZN(n14985) );
  OAI22_X1 U16823 ( .A1(n14986), .A2(n14985), .B1(n15009), .B2(n14984), .ZN(
        n14987) );
  XNOR2_X1 U16824 ( .A(n14987), .B(n14993), .ZN(n15280) );
  INV_X1 U16825 ( .A(n14988), .ZN(n14990) );
  NAND2_X1 U16826 ( .A1(n14990), .A2(n14989), .ZN(n14992) );
  INV_X1 U16827 ( .A(n14992), .ZN(n14991) );
  NAND2_X1 U16828 ( .A1(n14993), .A2(n14991), .ZN(n14999) );
  NAND2_X1 U16829 ( .A1(n14992), .A2(n14995), .ZN(n14994) );
  MUX2_X1 U16830 ( .A(n14994), .B(n14995), .S(n14993), .Z(n14998) );
  NAND3_X1 U16831 ( .A1(n15000), .A2(n14996), .A3(n14995), .ZN(n14997) );
  OAI211_X1 U16832 ( .C1(n15000), .C2(n14999), .A(n14998), .B(n14997), .ZN(
        n15281) );
  NAND2_X1 U16833 ( .A1(n15281), .A2(n15242), .ZN(n15014) );
  AOI21_X1 U16834 ( .B1(n15003), .B2(n15002), .A(n15001), .ZN(n15278) );
  INV_X1 U16835 ( .A(n15003), .ZN(n15275) );
  NOR3_X1 U16836 ( .A1(n15005), .A2(n15004), .A3(n15259), .ZN(n15006) );
  AOI21_X1 U16837 ( .B1(n15262), .B2(P1_REG2_REG_29__SCAN_IN), .A(n15006), 
        .ZN(n15011) );
  OAI22_X1 U16838 ( .A1(n15009), .A2(n15225), .B1(n15008), .B2(n15007), .ZN(
        n15276) );
  NAND2_X1 U16839 ( .A1(n15276), .A2(n15232), .ZN(n15010) );
  OAI211_X1 U16840 ( .C1(n15275), .C2(n15517), .A(n15011), .B(n15010), .ZN(
        n15012) );
  AOI21_X1 U16841 ( .B1(n15278), .B2(n15520), .A(n15012), .ZN(n15013) );
  OAI211_X1 U16842 ( .C1(n15245), .C2(n15280), .A(n15014), .B(n15013), .ZN(
        P1_U3356) );
  XNOR2_X1 U16843 ( .A(n6671), .B(n15021), .ZN(n15292) );
  INV_X1 U16844 ( .A(n15029), .ZN(n15017) );
  INV_X1 U16845 ( .A(n15015), .ZN(n15016) );
  AOI211_X1 U16846 ( .C1(n15289), .C2(n15017), .A(n15571), .B(n15016), .ZN(
        n15288) );
  AOI22_X1 U16847 ( .A1(n15018), .A2(n15513), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n15262), .ZN(n15019) );
  OAI21_X1 U16848 ( .B1(n15020), .B2(n15517), .A(n15019), .ZN(n15024) );
  OAI21_X1 U16849 ( .B1(n15292), .B2(n15267), .A(n15025), .ZN(P1_U3267) );
  AOI21_X1 U16850 ( .B1(n15039), .B2(n15027), .A(n15026), .ZN(n15028) );
  INV_X1 U16851 ( .A(n15028), .ZN(n15300) );
  AOI21_X1 U16852 ( .B1(n15030), .B2(n15055), .A(n15029), .ZN(n15293) );
  NOR2_X1 U16853 ( .A1(n15296), .A2(n15517), .ZN(n15037) );
  AOI22_X1 U16854 ( .A1(n15032), .A2(n15256), .B1(n15257), .B2(n15031), .ZN(
        n15294) );
  INV_X1 U16855 ( .A(n15033), .ZN(n15034) );
  AOI22_X1 U16856 ( .A1(n15034), .A2(n15513), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n15262), .ZN(n15035) );
  OAI21_X1 U16857 ( .B1(n15294), .B2(n15262), .A(n15035), .ZN(n15036) );
  AOI211_X1 U16858 ( .C1(n15293), .C2(n15520), .A(n15037), .B(n15036), .ZN(
        n15042) );
  OAI21_X1 U16859 ( .B1(n15040), .B2(n15039), .A(n15038), .ZN(n15298) );
  NAND2_X1 U16860 ( .A1(n15298), .A2(n7490), .ZN(n15041) );
  OAI211_X1 U16861 ( .C1(n15300), .C2(n15267), .A(n15042), .B(n15041), .ZN(
        P1_U3268) );
  XNOR2_X1 U16862 ( .A(n15043), .B(n15044), .ZN(n15301) );
  NAND2_X1 U16863 ( .A1(n15301), .A2(n15552), .ZN(n15052) );
  NOR2_X1 U16864 ( .A1(n15045), .A2(n15044), .ZN(n15047) );
  OR3_X1 U16865 ( .A1(n15047), .A2(n15046), .A3(n15360), .ZN(n15050) );
  INV_X1 U16866 ( .A(n15048), .ZN(n15049) );
  AND2_X1 U16867 ( .A1(n15050), .A2(n15049), .ZN(n15051) );
  NAND2_X1 U16868 ( .A1(n15052), .A2(n15051), .ZN(n15305) );
  INV_X1 U16869 ( .A(n15305), .ZN(n15062) );
  NAND2_X1 U16870 ( .A1(n15066), .A2(n15053), .ZN(n15054) );
  NAND2_X1 U16871 ( .A1(n15055), .A2(n15054), .ZN(n15302) );
  NOR2_X1 U16872 ( .A1(n15302), .A2(n15236), .ZN(n15060) );
  INV_X1 U16873 ( .A(n15056), .ZN(n15057) );
  AOI22_X1 U16874 ( .A1(n15057), .A2(n15513), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n15262), .ZN(n15058) );
  OAI21_X1 U16875 ( .B1(n7858), .B2(n15517), .A(n15058), .ZN(n15059) );
  AOI211_X1 U16876 ( .C1(n15301), .C2(n15521), .A(n15060), .B(n15059), .ZN(
        n15061) );
  OAI21_X1 U16877 ( .B1(n15062), .B2(n15262), .A(n15061), .ZN(P1_U3269) );
  XNOR2_X1 U16878 ( .A(n15063), .B(n15064), .ZN(n15313) );
  XNOR2_X1 U16879 ( .A(n15065), .B(n15064), .ZN(n15311) );
  OAI211_X1 U16880 ( .C1(n15079), .C2(n15309), .A(n15555), .B(n15066), .ZN(
        n15308) );
  NOR2_X1 U16881 ( .A1(n15308), .A2(n15067), .ZN(n15073) );
  INV_X1 U16882 ( .A(n15068), .ZN(n15069) );
  AOI22_X1 U16883 ( .A1(n15069), .A2(n15513), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n15262), .ZN(n15071) );
  NAND2_X1 U16884 ( .A1(n15306), .A2(n15232), .ZN(n15070) );
  OAI211_X1 U16885 ( .C1(n15309), .C2(n15517), .A(n15071), .B(n15070), .ZN(
        n15072) );
  AOI211_X1 U16886 ( .C1(n15311), .C2(n7490), .A(n15073), .B(n15072), .ZN(
        n15074) );
  OAI21_X1 U16887 ( .B1(n15313), .B2(n15267), .A(n15074), .ZN(P1_U3270) );
  OAI21_X1 U16888 ( .B1(n15077), .B2(n15076), .A(n15075), .ZN(n15078) );
  INV_X1 U16889 ( .A(n15078), .ZN(n15318) );
  INV_X1 U16890 ( .A(n15102), .ZN(n15080) );
  AOI21_X1 U16891 ( .B1(n15314), .B2(n15080), .A(n15079), .ZN(n15315) );
  INV_X1 U16892 ( .A(n15315), .ZN(n15087) );
  OAI21_X1 U16893 ( .B1(n15083), .B2(n15081), .A(n15082), .ZN(n15086) );
  INV_X1 U16894 ( .A(n15084), .ZN(n15085) );
  AOI21_X1 U16895 ( .B1(n15086), .B2(n15545), .A(n15085), .ZN(n15317) );
  OAI21_X1 U16896 ( .B1(n15138), .B2(n15087), .A(n15317), .ZN(n15092) );
  AOI22_X1 U16897 ( .A1(n15088), .A2(n15513), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n15262), .ZN(n15089) );
  OAI21_X1 U16898 ( .B1(n15090), .B2(n15517), .A(n15089), .ZN(n15091) );
  AOI21_X1 U16899 ( .B1(n15092), .B2(n15232), .A(n15091), .ZN(n15093) );
  OAI21_X1 U16900 ( .B1(n15318), .B2(n15267), .A(n15093), .ZN(P1_U3271) );
  NAND2_X1 U16901 ( .A1(n15115), .A2(n15122), .ZN(n15114) );
  NAND2_X1 U16902 ( .A1(n15114), .A2(n15096), .ZN(n15097) );
  XOR2_X1 U16903 ( .A(n15108), .B(n15097), .Z(n15101) );
  OAI22_X1 U16904 ( .A1(n15099), .A2(n15227), .B1(n15098), .B2(n15225), .ZN(
        n15100) );
  AOI21_X1 U16905 ( .B1(n15101), .B2(n15545), .A(n15100), .ZN(n15322) );
  INV_X1 U16906 ( .A(n15113), .ZN(n15103) );
  AOI21_X1 U16907 ( .B1(n15319), .B2(n15103), .A(n15102), .ZN(n15320) );
  INV_X1 U16908 ( .A(n15104), .ZN(n15105) );
  AOI22_X1 U16909 ( .A1(n15105), .A2(n15513), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n15262), .ZN(n15106) );
  OAI21_X1 U16910 ( .B1(n15107), .B2(n15517), .A(n15106), .ZN(n15111) );
  XOR2_X1 U16911 ( .A(n15109), .B(n15108), .Z(n15323) );
  NOR2_X1 U16912 ( .A1(n15323), .A2(n15267), .ZN(n15110) );
  AOI211_X1 U16913 ( .C1(n15320), .C2(n15520), .A(n15111), .B(n15110), .ZN(
        n15112) );
  OAI21_X1 U16914 ( .B1(n15262), .B2(n15322), .A(n15112), .ZN(P1_U3272) );
  INV_X1 U16915 ( .A(n15138), .ZN(n15121) );
  AOI21_X1 U16916 ( .B1(n15324), .B2(n15137), .A(n15113), .ZN(n15325) );
  OAI211_X1 U16917 ( .C1(n15115), .C2(n15122), .A(n15114), .B(n15545), .ZN(
        n15119) );
  AOI22_X1 U16918 ( .A1(n15117), .A2(n15256), .B1(n15257), .B2(n15116), .ZN(
        n15118) );
  AND2_X1 U16919 ( .A1(n15119), .A2(n15118), .ZN(n15327) );
  INV_X1 U16920 ( .A(n15327), .ZN(n15120) );
  AOI21_X1 U16921 ( .B1(n15121), .B2(n15325), .A(n15120), .ZN(n15131) );
  OAI21_X1 U16922 ( .B1(n15124), .B2(n8906), .A(n15123), .ZN(n15328) );
  INV_X1 U16923 ( .A(n15328), .ZN(n15129) );
  AOI22_X1 U16924 ( .A1(n15125), .A2(n15513), .B1(P1_REG2_REG_20__SCAN_IN), 
        .B2(n15262), .ZN(n15126) );
  OAI21_X1 U16925 ( .B1(n15127), .B2(n15517), .A(n15126), .ZN(n15128) );
  AOI21_X1 U16926 ( .B1(n15129), .B2(n15242), .A(n15128), .ZN(n15130) );
  OAI21_X1 U16927 ( .B1(n15131), .B2(n15262), .A(n15130), .ZN(P1_U3273) );
  XNOR2_X1 U16928 ( .A(n15133), .B(n15132), .ZN(n15336) );
  OAI21_X1 U16929 ( .B1(n15135), .B2(n15134), .A(n15094), .ZN(n15334) );
  NAND2_X1 U16930 ( .A1(n15330), .A2(n15161), .ZN(n15136) );
  NAND2_X1 U16931 ( .A1(n15137), .A2(n15136), .ZN(n15332) );
  NOR2_X1 U16932 ( .A1(n15332), .A2(n15138), .ZN(n15143) );
  NAND2_X1 U16933 ( .A1(n15139), .A2(n15256), .ZN(n15142) );
  NAND2_X1 U16934 ( .A1(n15140), .A2(n15257), .ZN(n15141) );
  NAND2_X1 U16935 ( .A1(n15142), .A2(n15141), .ZN(n15329) );
  OAI21_X1 U16936 ( .B1(n15143), .B2(n15329), .A(n15232), .ZN(n15146) );
  AOI22_X1 U16937 ( .A1(n15144), .A2(n15513), .B1(n15262), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n15145) );
  OAI211_X1 U16938 ( .C1(n7851), .C2(n15517), .A(n15146), .B(n15145), .ZN(
        n15147) );
  AOI21_X1 U16939 ( .B1(n15334), .B2(n7490), .A(n15147), .ZN(n15148) );
  OAI21_X1 U16940 ( .B1(n15336), .B2(n15267), .A(n15148), .ZN(P1_U3274) );
  XNOR2_X1 U16941 ( .A(n15149), .B(n15153), .ZN(n15341) );
  OAI21_X1 U16942 ( .B1(n15170), .B2(n15151), .A(n15150), .ZN(n15152) );
  INV_X1 U16943 ( .A(n15152), .ZN(n15175) );
  NOR3_X1 U16944 ( .A1(n15175), .A2(n15154), .A3(n15153), .ZN(n15158) );
  NAND2_X1 U16945 ( .A1(n15155), .A2(n15545), .ZN(n15157) );
  OAI21_X1 U16946 ( .B1(n15158), .B2(n15157), .A(n15156), .ZN(n15337) );
  INV_X1 U16947 ( .A(n15337), .ZN(n15165) );
  OR2_X1 U16948 ( .A1(n15180), .A2(n15159), .ZN(n15160) );
  AND3_X1 U16949 ( .A1(n15161), .A2(n15160), .A3(n15555), .ZN(n15338) );
  AOI22_X1 U16950 ( .A1(n15338), .A2(n15163), .B1(n15513), .B2(n15162), .ZN(
        n15164) );
  AOI21_X1 U16951 ( .B1(n15165), .B2(n15164), .A(n15262), .ZN(n15166) );
  INV_X1 U16952 ( .A(n15166), .ZN(n15168) );
  AOI22_X1 U16953 ( .A1(n15339), .A2(n15239), .B1(n15262), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n15167) );
  OAI211_X1 U16954 ( .C1(n15169), .C2(n15341), .A(n15168), .B(n15167), .ZN(
        P1_U3275) );
  NOR2_X1 U16955 ( .A1(n8937), .A2(n15210), .ZN(n15209) );
  NOR2_X1 U16956 ( .A1(n15209), .A2(n15171), .ZN(n15192) );
  NAND2_X1 U16957 ( .A1(n15192), .A2(n15191), .ZN(n15190) );
  AOI21_X1 U16958 ( .B1(n15190), .B2(n15174), .A(n15173), .ZN(n15176) );
  NOR3_X1 U16959 ( .A1(n15176), .A2(n15360), .A3(n15175), .ZN(n15179) );
  OAI22_X1 U16960 ( .A1(n15177), .A2(n15227), .B1(n15214), .B2(n15225), .ZN(
        n15178) );
  NOR2_X1 U16961 ( .A1(n15179), .A2(n15178), .ZN(n15345) );
  AOI21_X1 U16962 ( .B1(n15342), .B2(n15194), .A(n15180), .ZN(n15343) );
  AOI22_X1 U16963 ( .A1(n15262), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n15181), 
        .B2(n15513), .ZN(n15182) );
  OAI21_X1 U16964 ( .B1(n15183), .B2(n15517), .A(n15182), .ZN(n15187) );
  XNOR2_X1 U16965 ( .A(n15185), .B(n15184), .ZN(n15346) );
  NOR2_X1 U16966 ( .A1(n15346), .A2(n15267), .ZN(n15186) );
  AOI211_X1 U16967 ( .C1(n15343), .C2(n15520), .A(n15187), .B(n15186), .ZN(
        n15188) );
  OAI21_X1 U16968 ( .B1(n15345), .B2(n15262), .A(n15188), .ZN(P1_U3276) );
  XNOR2_X1 U16969 ( .A(n15189), .B(n15191), .ZN(n15353) );
  OAI21_X1 U16970 ( .B1(n15192), .B2(n15191), .A(n15190), .ZN(n15347) );
  NAND2_X1 U16971 ( .A1(n15347), .A2(n7490), .ZN(n15205) );
  INV_X1 U16972 ( .A(n15194), .ZN(n15195) );
  AOI211_X1 U16973 ( .C1(n15350), .C2(n15211), .A(n15571), .B(n15195), .ZN(
        n15348) );
  INV_X1 U16974 ( .A(n15348), .ZN(n15200) );
  OAI22_X1 U16975 ( .A1(n15196), .A2(n15227), .B1(n15228), .B2(n15225), .ZN(
        n15349) );
  AOI21_X1 U16976 ( .B1(n15197), .B2(n15513), .A(n15349), .ZN(n15198) );
  OAI21_X1 U16977 ( .B1(n15200), .B2(n15199), .A(n15198), .ZN(n15203) );
  INV_X1 U16978 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n15201) );
  OAI22_X1 U16979 ( .A1(n8968), .A2(n15517), .B1(n15232), .B2(n15201), .ZN(
        n15202) );
  AOI21_X1 U16980 ( .B1(n15203), .B2(n15232), .A(n15202), .ZN(n15204) );
  OAI211_X1 U16981 ( .C1(n15353), .C2(n15267), .A(n15205), .B(n15204), .ZN(
        P1_U3277) );
  NOR2_X1 U16982 ( .A1(n15206), .A2(n15241), .ZN(n15240) );
  NOR2_X1 U16983 ( .A1(n15240), .A2(n15207), .ZN(n15208) );
  XOR2_X1 U16984 ( .A(n15210), .B(n15208), .Z(n15359) );
  AOI21_X1 U16985 ( .B1(n8937), .B2(n15210), .A(n15209), .ZN(n15354) );
  NAND2_X1 U16986 ( .A1(n15354), .A2(n7490), .ZN(n15221) );
  INV_X1 U16987 ( .A(n15211), .ZN(n15212) );
  AOI211_X1 U16988 ( .C1(n8898), .C2(n15235), .A(n15571), .B(n15212), .ZN(
        n15355) );
  OAI22_X1 U16989 ( .A1(n15214), .A2(n15227), .B1(n15213), .B2(n15225), .ZN(
        n15356) );
  AOI22_X1 U16990 ( .A1(n15232), .A2(n15356), .B1(n15215), .B2(n15513), .ZN(
        n15217) );
  NAND2_X1 U16991 ( .A1(n15262), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n15216) );
  OAI211_X1 U16992 ( .C1(n15218), .C2(n15517), .A(n15217), .B(n15216), .ZN(
        n15219) );
  AOI21_X1 U16993 ( .B1(n15355), .B2(n15254), .A(n15219), .ZN(n15220) );
  OAI211_X1 U16994 ( .C1(n15359), .C2(n15267), .A(n15221), .B(n15220), .ZN(
        P1_U3278) );
  OR2_X1 U16995 ( .A1(n15222), .A2(n15241), .ZN(n15223) );
  NAND2_X1 U16996 ( .A1(n15224), .A2(n15223), .ZN(n15361) );
  OAI22_X1 U16997 ( .A1(n15228), .A2(n15227), .B1(n15226), .B2(n15225), .ZN(
        n15363) );
  INV_X1 U16998 ( .A(n15229), .ZN(n15230) );
  AOI22_X1 U16999 ( .A1(n15232), .A2(n15363), .B1(n15230), .B2(n15513), .ZN(
        n15231) );
  OAI21_X1 U17000 ( .B1(n10775), .B2(n15232), .A(n15231), .ZN(n15238) );
  INV_X1 U17001 ( .A(n15252), .ZN(n15233) );
  NAND2_X1 U17002 ( .A1(n15233), .A2(n8965), .ZN(n15234) );
  NAND2_X1 U17003 ( .A1(n15235), .A2(n15234), .ZN(n15365) );
  NOR2_X1 U17004 ( .A1(n15365), .A2(n15236), .ZN(n15237) );
  AOI211_X1 U17005 ( .C1(n15239), .C2(n8965), .A(n15238), .B(n15237), .ZN(
        n15244) );
  INV_X1 U17006 ( .A(n15240), .ZN(n15368) );
  NAND2_X1 U17007 ( .A1(n15206), .A2(n15241), .ZN(n15362) );
  NAND3_X1 U17008 ( .A1(n15368), .A2(n15242), .A3(n15362), .ZN(n15243) );
  OAI211_X1 U17009 ( .C1(n15361), .C2(n15245), .A(n15244), .B(n15243), .ZN(
        P1_U3279) );
  XNOR2_X1 U17010 ( .A(n15246), .B(n15248), .ZN(n15377) );
  OAI21_X1 U17011 ( .B1(n15249), .B2(n15248), .A(n15247), .ZN(n15250) );
  INV_X1 U17012 ( .A(n15250), .ZN(n15375) );
  OAI21_X1 U17013 ( .B1(n15251), .B2(n15372), .A(n15555), .ZN(n15253) );
  NOR2_X1 U17014 ( .A1(n15253), .A2(n15252), .ZN(n15374) );
  NAND2_X1 U17015 ( .A1(n15374), .A2(n15254), .ZN(n15264) );
  AOI22_X1 U17016 ( .A1(n15258), .A2(n15257), .B1(n15256), .B2(n15255), .ZN(
        n15371) );
  OAI22_X1 U17017 ( .A1(n15262), .A2(n15371), .B1(n15260), .B2(n15259), .ZN(
        n15261) );
  AOI21_X1 U17018 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n15262), .A(n15261), 
        .ZN(n15263) );
  OAI211_X1 U17019 ( .C1(n15372), .C2(n15517), .A(n15264), .B(n15263), .ZN(
        n15265) );
  AOI21_X1 U17020 ( .B1(n15375), .B2(n7490), .A(n15265), .ZN(n15266) );
  OAI21_X1 U17021 ( .B1(n15267), .B2(n15377), .A(n15266), .ZN(P1_U3280) );
  AOI21_X1 U17022 ( .B1(n15269), .B2(n15580), .A(n15268), .ZN(n15270) );
  OAI21_X1 U17023 ( .B1(n15271), .B2(n15571), .A(n15270), .ZN(n15400) );
  MUX2_X1 U17024 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15400), .S(n15599), .Z(
        P1_U3559) );
  OAI211_X1 U17025 ( .C1(n15274), .C2(n15569), .A(n15273), .B(n15272), .ZN(
        n15401) );
  MUX2_X1 U17026 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15401), .S(n15599), .Z(
        P1_U3558) );
  NOR2_X1 U17027 ( .A1(n15275), .A2(n15569), .ZN(n15277) );
  NAND2_X1 U17028 ( .A1(n15281), .A2(n15578), .ZN(n15282) );
  MUX2_X1 U17029 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n15402), .S(n15599), .Z(
        P1_U3557) );
  AOI21_X1 U17030 ( .B1(n15580), .B2(n15284), .A(n15283), .ZN(n15285) );
  OAI211_X1 U17031 ( .C1(n15287), .C2(n15560), .A(n15286), .B(n15285), .ZN(
        n15403) );
  MUX2_X1 U17032 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15403), .S(n15599), .Z(
        P1_U3555) );
  AOI21_X1 U17033 ( .B1(n15580), .B2(n15289), .A(n15288), .ZN(n15290) );
  OAI211_X1 U17034 ( .C1(n15292), .C2(n15560), .A(n15291), .B(n15290), .ZN(
        n15404) );
  MUX2_X1 U17035 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15404), .S(n15599), .Z(
        P1_U3554) );
  NAND2_X1 U17036 ( .A1(n15293), .A2(n15555), .ZN(n15295) );
  OAI211_X1 U17037 ( .C1(n15296), .C2(n15569), .A(n15295), .B(n15294), .ZN(
        n15297) );
  AOI21_X1 U17038 ( .B1(n15298), .B2(n15545), .A(n15297), .ZN(n15299) );
  OAI21_X1 U17039 ( .B1(n15300), .B2(n15560), .A(n15299), .ZN(n15405) );
  MUX2_X1 U17040 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15405), .S(n15599), .Z(
        P1_U3553) );
  AND2_X1 U17041 ( .A1(n15301), .A2(n15574), .ZN(n15304) );
  OAI22_X1 U17042 ( .A1(n15302), .A2(n15571), .B1(n7858), .B2(n15569), .ZN(
        n15303) );
  MUX2_X1 U17043 ( .A(n15406), .B(P1_REG1_REG_24__SCAN_IN), .S(n15597), .Z(
        P1_U3552) );
  INV_X1 U17044 ( .A(n15306), .ZN(n15307) );
  OAI211_X1 U17045 ( .C1(n15309), .C2(n15569), .A(n15308), .B(n15307), .ZN(
        n15310) );
  AOI21_X1 U17046 ( .B1(n15311), .B2(n15545), .A(n15310), .ZN(n15312) );
  OAI21_X1 U17047 ( .B1(n15313), .B2(n15560), .A(n15312), .ZN(n15407) );
  MUX2_X1 U17048 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15407), .S(n15599), .Z(
        P1_U3551) );
  AOI22_X1 U17049 ( .A1(n15315), .A2(n15555), .B1(n15314), .B2(n15580), .ZN(
        n15316) );
  OAI211_X1 U17050 ( .C1(n15318), .C2(n15560), .A(n15317), .B(n15316), .ZN(
        n15408) );
  MUX2_X1 U17051 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15408), .S(n15599), .Z(
        P1_U3550) );
  AOI22_X1 U17052 ( .A1(n15320), .A2(n15555), .B1(n15580), .B2(n15319), .ZN(
        n15321) );
  OAI211_X1 U17053 ( .C1(n15560), .C2(n15323), .A(n15322), .B(n15321), .ZN(
        n15409) );
  MUX2_X1 U17054 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15409), .S(n15599), .Z(
        P1_U3549) );
  AOI22_X1 U17055 ( .A1(n15325), .A2(n15555), .B1(n15580), .B2(n15324), .ZN(
        n15326) );
  OAI211_X1 U17056 ( .C1(n15560), .C2(n15328), .A(n15327), .B(n15326), .ZN(
        n15410) );
  MUX2_X1 U17057 ( .A(n15410), .B(P1_REG1_REG_20__SCAN_IN), .S(n15597), .Z(
        P1_U3548) );
  AOI21_X1 U17058 ( .B1(n15330), .B2(n15580), .A(n15329), .ZN(n15331) );
  OAI21_X1 U17059 ( .B1(n15332), .B2(n15571), .A(n15331), .ZN(n15333) );
  AOI21_X1 U17060 ( .B1(n15334), .B2(n15545), .A(n15333), .ZN(n15335) );
  OAI21_X1 U17061 ( .B1(n15560), .B2(n15336), .A(n15335), .ZN(n15411) );
  MUX2_X1 U17062 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15411), .S(n15599), .Z(
        P1_U3547) );
  AOI211_X1 U17063 ( .C1(n15580), .C2(n15339), .A(n15338), .B(n15337), .ZN(
        n15340) );
  OAI21_X1 U17064 ( .B1(n15560), .B2(n15341), .A(n15340), .ZN(n15412) );
  MUX2_X1 U17065 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15412), .S(n15599), .Z(
        P1_U3546) );
  AOI22_X1 U17066 ( .A1(n15343), .A2(n15555), .B1(n15580), .B2(n15342), .ZN(
        n15344) );
  OAI211_X1 U17067 ( .C1(n15560), .C2(n15346), .A(n15345), .B(n15344), .ZN(
        n15413) );
  MUX2_X1 U17068 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15413), .S(n15599), .Z(
        P1_U3545) );
  NAND2_X1 U17069 ( .A1(n15347), .A2(n15545), .ZN(n15352) );
  AOI211_X1 U17070 ( .C1(n15580), .C2(n15350), .A(n15349), .B(n15348), .ZN(
        n15351) );
  OAI211_X1 U17071 ( .C1(n15560), .C2(n15353), .A(n15352), .B(n15351), .ZN(
        n15414) );
  MUX2_X1 U17072 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15414), .S(n15599), .Z(
        P1_U3544) );
  NAND2_X1 U17073 ( .A1(n15354), .A2(n15545), .ZN(n15358) );
  AOI211_X1 U17074 ( .C1(n15580), .C2(n8898), .A(n15356), .B(n15355), .ZN(
        n15357) );
  OAI211_X1 U17075 ( .C1(n15560), .C2(n15359), .A(n15358), .B(n15357), .ZN(
        n15415) );
  MUX2_X1 U17076 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15415), .S(n15599), .Z(
        P1_U3543) );
  OR2_X1 U17077 ( .A1(n15361), .A2(n15360), .ZN(n15370) );
  AND2_X1 U17078 ( .A1(n15362), .A2(n15578), .ZN(n15367) );
  AOI21_X1 U17079 ( .B1(n8965), .B2(n15580), .A(n15363), .ZN(n15364) );
  OAI21_X1 U17080 ( .B1(n15365), .B2(n15571), .A(n15364), .ZN(n15366) );
  AOI21_X1 U17081 ( .B1(n15368), .B2(n15367), .A(n15366), .ZN(n15369) );
  NAND2_X1 U17082 ( .A1(n15370), .A2(n15369), .ZN(n15416) );
  MUX2_X1 U17083 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15416), .S(n15599), .Z(
        P1_U3542) );
  OAI21_X1 U17084 ( .B1(n15372), .B2(n15569), .A(n15371), .ZN(n15373) );
  AOI211_X1 U17085 ( .C1(n15375), .C2(n15545), .A(n15374), .B(n15373), .ZN(
        n15376) );
  OAI21_X1 U17086 ( .B1(n15560), .B2(n15377), .A(n15376), .ZN(n15417) );
  MUX2_X1 U17087 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n15417), .S(n15599), .Z(
        P1_U3541) );
  OAI22_X1 U17088 ( .A1(n15378), .A2(n15571), .B1(n7847), .B2(n15569), .ZN(
        n15379) );
  INV_X1 U17089 ( .A(n15379), .ZN(n15380) );
  OAI21_X1 U17090 ( .B1(n15381), .B2(n15548), .A(n15380), .ZN(n15382) );
  MUX2_X1 U17091 ( .A(n15418), .B(P1_REG1_REG_12__SCAN_IN), .S(n15597), .Z(
        P1_U3540) );
  AOI22_X1 U17092 ( .A1(n15385), .A2(n15555), .B1(n15580), .B2(n15384), .ZN(
        n15386) );
  OAI211_X1 U17093 ( .C1(n15560), .C2(n15388), .A(n15387), .B(n15386), .ZN(
        n15419) );
  MUX2_X1 U17094 ( .A(n15419), .B(P1_REG1_REG_11__SCAN_IN), .S(n15597), .Z(
        P1_U3539) );
  AOI211_X1 U17095 ( .C1(n15580), .C2(n15391), .A(n15390), .B(n15389), .ZN(
        n15392) );
  OAI211_X1 U17096 ( .C1(n15560), .C2(n15394), .A(n15393), .B(n15392), .ZN(
        n15420) );
  MUX2_X1 U17097 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n15420), .S(n15599), .Z(
        P1_U3538) );
  AOI21_X1 U17098 ( .B1(n15580), .B2(n15396), .A(n15395), .ZN(n15397) );
  OAI211_X1 U17099 ( .C1(n15560), .C2(n15399), .A(n15398), .B(n15397), .ZN(
        n15421) );
  MUX2_X1 U17100 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n15421), .S(n15599), .Z(
        P1_U3537) );
  MUX2_X1 U17101 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15400), .S(n15588), .Z(
        P1_U3527) );
  MUX2_X1 U17102 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15401), .S(n15588), .Z(
        P1_U3526) );
  MUX2_X1 U17103 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n15402), .S(n15588), .Z(
        P1_U3525) );
  MUX2_X1 U17104 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15403), .S(n15588), .Z(
        P1_U3523) );
  MUX2_X1 U17105 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15404), .S(n15588), .Z(
        P1_U3522) );
  MUX2_X1 U17106 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15405), .S(n15588), .Z(
        P1_U3521) );
  MUX2_X1 U17107 ( .A(n15406), .B(P1_REG0_REG_24__SCAN_IN), .S(n15587), .Z(
        P1_U3520) );
  MUX2_X1 U17108 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15407), .S(n15588), .Z(
        P1_U3519) );
  MUX2_X1 U17109 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15408), .S(n15588), .Z(
        P1_U3518) );
  MUX2_X1 U17110 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15409), .S(n15588), .Z(
        P1_U3517) );
  MUX2_X1 U17111 ( .A(n15410), .B(P1_REG0_REG_20__SCAN_IN), .S(n15587), .Z(
        P1_U3516) );
  MUX2_X1 U17112 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15411), .S(n15588), .Z(
        P1_U3515) );
  MUX2_X1 U17113 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15412), .S(n15588), .Z(
        P1_U3513) );
  MUX2_X1 U17114 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15413), .S(n15588), .Z(
        P1_U3510) );
  MUX2_X1 U17115 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15414), .S(n15588), .Z(
        P1_U3507) );
  MUX2_X1 U17116 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15415), .S(n15588), .Z(
        P1_U3504) );
  MUX2_X1 U17117 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15416), .S(n15588), .Z(
        P1_U3501) );
  MUX2_X1 U17118 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n15417), .S(n15588), .Z(
        P1_U3498) );
  MUX2_X1 U17119 ( .A(n15418), .B(P1_REG0_REG_12__SCAN_IN), .S(n15587), .Z(
        P1_U3495) );
  MUX2_X1 U17120 ( .A(n15419), .B(P1_REG0_REG_11__SCAN_IN), .S(n15587), .Z(
        P1_U3492) );
  MUX2_X1 U17121 ( .A(P1_REG0_REG_10__SCAN_IN), .B(n15420), .S(n15588), .Z(
        P1_U3489) );
  MUX2_X1 U17122 ( .A(P1_REG0_REG_9__SCAN_IN), .B(n15421), .S(n15588), .Z(
        P1_U3486) );
  NOR4_X1 U17123 ( .A1(n6721), .A2(P1_IR_REG_30__SCAN_IN), .A3(n15422), .A4(
        P1_U3086), .ZN(n15423) );
  AOI21_X1 U17124 ( .B1(n15424), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n15423), 
        .ZN(n15425) );
  OAI21_X1 U17125 ( .B1(n15426), .B2(n15438), .A(n15425), .ZN(P1_U3324) );
  OAI222_X1 U17126 ( .A1(n15435), .A2(n15429), .B1(P1_U3086), .B2(n15427), 
        .C1(n15438), .C2(n15428), .ZN(P1_U3325) );
  OAI222_X1 U17127 ( .A1(n15435), .A2(n15432), .B1(P1_U3086), .B2(n15431), 
        .C1(n15438), .C2(n15430), .ZN(P1_U3326) );
  OAI222_X1 U17128 ( .A1(n15435), .A2(n7803), .B1(n15438), .B2(n15434), .C1(
        P1_U3086), .C2(n15433), .ZN(P1_U3328) );
  OAI222_X1 U17129 ( .A1(n15439), .A2(P1_U3086), .B1(n15438), .B2(n15437), 
        .C1(n15436), .C2(n15435), .ZN(P1_U3329) );
  MUX2_X1 U17130 ( .A(n15441), .B(n15440), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U17131 ( .A(n15442), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U17132 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n15756) );
  AOI21_X1 U17133 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15446) );
  OAI21_X1 U17134 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n15446), 
        .ZN(U28) );
  AOI21_X1 U17135 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n15447) );
  OAI21_X1 U17136 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n15447), 
        .ZN(U29) );
  OAI222_X1 U17137 ( .A1(n15452), .A2(n15451), .B1(n15452), .B2(n15450), .C1(
        n15449), .C2(n15448), .ZN(SUB_1596_U61) );
  AOI21_X1 U17138 ( .B1(n15455), .B2(n15454), .A(n15453), .ZN(SUB_1596_U57) );
  OAI21_X1 U17139 ( .B1(n15457), .B2(n15663), .A(n15456), .ZN(SUB_1596_U55) );
  OAI21_X1 U17140 ( .B1(n15460), .B2(n15459), .A(n15458), .ZN(n15461) );
  XOR2_X1 U17141 ( .A(n15461), .B(n9744), .Z(SUB_1596_U54) );
  AOI21_X1 U17142 ( .B1(n15464), .B2(n15463), .A(n15462), .ZN(n15465) );
  XOR2_X1 U17143 ( .A(n15465), .B(P2_ADDR_REG_10__SCAN_IN), .Z(SUB_1596_U70)
         );
  AOI21_X1 U17144 ( .B1(n15468), .B2(n15467), .A(n15466), .ZN(n15469) );
  XNOR2_X1 U17145 ( .A(n7564), .B(n15469), .ZN(SUB_1596_U63) );
  OAI222_X1 U17146 ( .A1(n15474), .A2(n15473), .B1(n15474), .B2(n15472), .C1(
        n15471), .C2(n15470), .ZN(SUB_1596_U69) );
  OAI21_X1 U17147 ( .B1(n15477), .B2(n15476), .A(n15475), .ZN(n15478) );
  XOR2_X1 U17148 ( .A(n15478), .B(n15705), .Z(SUB_1596_U68) );
  AOI21_X1 U17149 ( .B1(n15481), .B2(n15480), .A(n15479), .ZN(n15482) );
  XNOR2_X1 U17150 ( .A(n7734), .B(n15482), .ZN(SUB_1596_U67) );
  OAI21_X1 U17151 ( .B1(n15485), .B2(n15484), .A(n15483), .ZN(n15486) );
  XOR2_X1 U17152 ( .A(n15486), .B(n9755), .Z(SUB_1596_U66) );
  INV_X1 U17153 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15727) );
  AOI21_X1 U17154 ( .B1(n15489), .B2(n15488), .A(n15487), .ZN(n15490) );
  XNOR2_X1 U17155 ( .A(n15727), .B(n15490), .ZN(SUB_1596_U65) );
  OAI21_X1 U17156 ( .B1(n15493), .B2(n15492), .A(n15491), .ZN(n15494) );
  INV_X1 U17157 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15742) );
  XOR2_X1 U17158 ( .A(n15494), .B(n15742), .Z(SUB_1596_U64) );
  AOI21_X1 U17159 ( .B1(n15495), .B2(n15497), .A(n15496), .ZN(n15506) );
  AOI22_X1 U17160 ( .A1(n15500), .A2(n15499), .B1(P1_U3086), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n15501) );
  OAI21_X1 U17161 ( .B1(n15503), .B2(n15502), .A(n15501), .ZN(n15504) );
  AOI21_X1 U17162 ( .B1(n15506), .B2(n15505), .A(n15504), .ZN(n15507) );
  OAI21_X1 U17163 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(n15508), .A(n15507), .ZN(
        P1_U3218) );
  INV_X1 U17164 ( .A(n15509), .ZN(n15522) );
  INV_X1 U17165 ( .A(n15510), .ZN(n15511) );
  AOI21_X1 U17166 ( .B1(n15552), .B2(n15522), .A(n15511), .ZN(n15525) );
  INV_X1 U17167 ( .A(n15512), .ZN(n15514) );
  AOI22_X1 U17168 ( .A1(n15262), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n15514), 
        .B2(n15513), .ZN(n15515) );
  OAI21_X1 U17169 ( .B1(n15517), .B2(n15516), .A(n15515), .ZN(n15518) );
  INV_X1 U17170 ( .A(n15518), .ZN(n15524) );
  AOI22_X1 U17171 ( .A1(n15522), .A2(n15521), .B1(n15520), .B2(n15519), .ZN(
        n15523) );
  OAI211_X1 U17172 ( .C1(n15262), .C2(n15525), .A(n15524), .B(n15523), .ZN(
        P1_U3286) );
  AND2_X1 U17173 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15531), .ZN(P1_U3294) );
  INV_X1 U17174 ( .A(n15531), .ZN(n15530) );
  NOR2_X1 U17175 ( .A1(n15530), .A2(n15526), .ZN(P1_U3295) );
  AND2_X1 U17176 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15531), .ZN(P1_U3296) );
  AND2_X1 U17177 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15531), .ZN(P1_U3297) );
  AND2_X1 U17178 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15531), .ZN(P1_U3298) );
  AND2_X1 U17179 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15531), .ZN(P1_U3299) );
  AND2_X1 U17180 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15531), .ZN(P1_U3300) );
  AND2_X1 U17181 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15531), .ZN(P1_U3301) );
  AND2_X1 U17182 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15531), .ZN(P1_U3302) );
  AND2_X1 U17183 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15531), .ZN(P1_U3303) );
  AND2_X1 U17184 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15531), .ZN(P1_U3304) );
  AND2_X1 U17185 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15531), .ZN(P1_U3305) );
  AND2_X1 U17186 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15531), .ZN(P1_U3306) );
  AND2_X1 U17187 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15531), .ZN(P1_U3307) );
  AND2_X1 U17188 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15531), .ZN(P1_U3308) );
  AND2_X1 U17189 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15531), .ZN(P1_U3309) );
  NOR2_X1 U17190 ( .A1(n15530), .A2(n15527), .ZN(P1_U3310) );
  AND2_X1 U17191 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15531), .ZN(P1_U3311) );
  AND2_X1 U17192 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15531), .ZN(P1_U3312) );
  AND2_X1 U17193 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15531), .ZN(P1_U3313) );
  NOR2_X1 U17194 ( .A1(n15530), .A2(n15528), .ZN(P1_U3314) );
  AND2_X1 U17195 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15531), .ZN(P1_U3315) );
  AND2_X1 U17196 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15531), .ZN(P1_U3316) );
  AND2_X1 U17197 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15531), .ZN(P1_U3317) );
  AND2_X1 U17198 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15531), .ZN(P1_U3318) );
  AND2_X1 U17199 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15531), .ZN(P1_U3319) );
  AND2_X1 U17200 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15531), .ZN(P1_U3320) );
  NOR2_X1 U17201 ( .A1(n15530), .A2(n15529), .ZN(P1_U3321) );
  AND2_X1 U17202 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15531), .ZN(P1_U3322) );
  AND2_X1 U17203 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15531), .ZN(P1_U3323) );
  INV_X1 U17204 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15532) );
  AOI22_X1 U17205 ( .A1(n15588), .A2(n15533), .B1(n15532), .B2(n15587), .ZN(
        P1_U3459) );
  INV_X1 U17206 ( .A(n15534), .ZN(n15539) );
  OAI22_X1 U17207 ( .A1(n15536), .A2(n15571), .B1(n15535), .B2(n15569), .ZN(
        n15538) );
  AOI211_X1 U17208 ( .C1(n15574), .C2(n15539), .A(n15538), .B(n15537), .ZN(
        n15590) );
  INV_X1 U17209 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15540) );
  AOI22_X1 U17210 ( .A1(n15588), .A2(n15590), .B1(n15540), .B2(n15587), .ZN(
        P1_U3462) );
  INV_X1 U17211 ( .A(n15549), .ZN(n15551) );
  INV_X1 U17212 ( .A(n15541), .ZN(n15542) );
  OAI211_X1 U17213 ( .C1(n8299), .C2(n15569), .A(n15543), .B(n15542), .ZN(
        n15544) );
  AOI21_X1 U17214 ( .B1(n15546), .B2(n15545), .A(n15544), .ZN(n15547) );
  OAI21_X1 U17215 ( .B1(n15549), .B2(n15548), .A(n15547), .ZN(n15550) );
  AOI21_X1 U17216 ( .B1(n15552), .B2(n15551), .A(n15550), .ZN(n15592) );
  AOI22_X1 U17217 ( .A1(n15588), .A2(n15592), .B1(n15553), .B2(n15587), .ZN(
        P1_U3465) );
  AOI22_X1 U17218 ( .A1(n15556), .A2(n15555), .B1(n15580), .B2(n15554), .ZN(
        n15557) );
  OAI211_X1 U17219 ( .C1(n15560), .C2(n15559), .A(n15558), .B(n15557), .ZN(
        n15561) );
  INV_X1 U17220 ( .A(n15561), .ZN(n15594) );
  AOI22_X1 U17221 ( .A1(n15588), .A2(n15594), .B1(n8229), .B2(n15587), .ZN(
        P1_U3471) );
  INV_X1 U17222 ( .A(n15562), .ZN(n15567) );
  OAI22_X1 U17223 ( .A1(n15564), .A2(n15571), .B1(n15563), .B2(n15569), .ZN(
        n15566) );
  AOI211_X1 U17224 ( .C1(n15574), .C2(n15567), .A(n15566), .B(n15565), .ZN(
        n15595) );
  INV_X1 U17225 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15568) );
  AOI22_X1 U17226 ( .A1(n15588), .A2(n15595), .B1(n15568), .B2(n15587), .ZN(
        P1_U3474) );
  OAI22_X1 U17227 ( .A1(n15572), .A2(n15571), .B1(n15570), .B2(n15569), .ZN(
        n15573) );
  AOI21_X1 U17228 ( .B1(n15575), .B2(n15574), .A(n15573), .ZN(n15576) );
  AND2_X1 U17229 ( .A1(n15577), .A2(n15576), .ZN(n15596) );
  AOI22_X1 U17230 ( .A1(n15588), .A2(n15596), .B1(n8314), .B2(n15587), .ZN(
        P1_U3477) );
  AND2_X1 U17231 ( .A1(n15579), .A2(n15578), .ZN(n15585) );
  NAND2_X1 U17232 ( .A1(n15581), .A2(n15580), .ZN(n15582) );
  NAND2_X1 U17233 ( .A1(n15583), .A2(n15582), .ZN(n15584) );
  NOR3_X1 U17234 ( .A1(n15586), .A2(n15585), .A3(n15584), .ZN(n15598) );
  AOI22_X1 U17235 ( .A1(n15588), .A2(n15598), .B1(n8356), .B2(n15587), .ZN(
        P1_U3483) );
  AOI22_X1 U17236 ( .A1(n15599), .A2(n15590), .B1(n15589), .B2(n15597), .ZN(
        P1_U3529) );
  AOI22_X1 U17237 ( .A1(n15599), .A2(n15592), .B1(n15591), .B2(n15597), .ZN(
        P1_U3530) );
  AOI22_X1 U17238 ( .A1(n15599), .A2(n15594), .B1(n15593), .B2(n15597), .ZN(
        P1_U3532) );
  AOI22_X1 U17239 ( .A1(n15599), .A2(n15595), .B1(n8221), .B2(n15597), .ZN(
        P1_U3533) );
  AOI22_X1 U17240 ( .A1(n15599), .A2(n15596), .B1(n10731), .B2(n15597), .ZN(
        P1_U3534) );
  AOI22_X1 U17241 ( .A1(n15599), .A2(n15598), .B1(n8352), .B2(n15597), .ZN(
        P1_U3536) );
  NOR2_X1 U17242 ( .A1(n15600), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U17243 ( .A1(n15600), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n6510), .ZN(n15612) );
  OAI211_X1 U17244 ( .C1(n15603), .C2(n15602), .A(n15744), .B(n15601), .ZN(
        n15608) );
  OAI211_X1 U17245 ( .C1(n15606), .C2(n15605), .A(n15752), .B(n15604), .ZN(
        n15607) );
  OAI211_X1 U17246 ( .C1(n15749), .C2(n15609), .A(n15608), .B(n15607), .ZN(
        n15610) );
  INV_X1 U17247 ( .A(n15610), .ZN(n15611) );
  NAND2_X1 U17248 ( .A1(n15612), .A2(n15611), .ZN(P2_U3216) );
  OAI211_X1 U17249 ( .C1(n15615), .C2(n15614), .A(n15744), .B(n15613), .ZN(
        n15620) );
  OAI211_X1 U17250 ( .C1(n15618), .C2(n15617), .A(n15752), .B(n15616), .ZN(
        n15619) );
  OAI211_X1 U17251 ( .C1(n15749), .C2(n15621), .A(n15620), .B(n15619), .ZN(
        n15622) );
  INV_X1 U17252 ( .A(n15622), .ZN(n15624) );
  OAI211_X1 U17253 ( .C1(n15755), .C2(n15625), .A(n15624), .B(n15623), .ZN(
        P2_U3218) );
  OAI211_X1 U17254 ( .C1(n15628), .C2(n15627), .A(n15744), .B(n15626), .ZN(
        n15633) );
  OAI211_X1 U17255 ( .C1(n15631), .C2(n15630), .A(n15752), .B(n15629), .ZN(
        n15632) );
  OAI211_X1 U17256 ( .C1(n15749), .C2(n15634), .A(n15633), .B(n15632), .ZN(
        n15635) );
  INV_X1 U17257 ( .A(n15635), .ZN(n15637) );
  NAND2_X1 U17258 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(n6510), .ZN(n15636) );
  OAI211_X1 U17259 ( .C1(n15755), .C2(n15922), .A(n15637), .B(n15636), .ZN(
        P2_U3219) );
  OAI211_X1 U17260 ( .C1(n15640), .C2(n15639), .A(n15744), .B(n15638), .ZN(
        n15645) );
  OAI211_X1 U17261 ( .C1(n15643), .C2(n15642), .A(n15752), .B(n15641), .ZN(
        n15644) );
  OAI211_X1 U17262 ( .C1(n15749), .C2(n15646), .A(n15645), .B(n15644), .ZN(
        n15647) );
  INV_X1 U17263 ( .A(n15647), .ZN(n15650) );
  NAND2_X1 U17264 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n15649) );
  OAI211_X1 U17265 ( .C1(n15755), .C2(n7735), .A(n15650), .B(n15649), .ZN(
        P2_U3220) );
  OAI211_X1 U17266 ( .C1(n15653), .C2(n15652), .A(n15744), .B(n15651), .ZN(
        n15658) );
  OAI211_X1 U17267 ( .C1(n15656), .C2(n15655), .A(n15752), .B(n15654), .ZN(
        n15657) );
  OAI211_X1 U17268 ( .C1(n15749), .C2(n15659), .A(n15658), .B(n15657), .ZN(
        n15660) );
  INV_X1 U17269 ( .A(n15660), .ZN(n15662) );
  OAI211_X1 U17270 ( .C1(n15663), .C2(n15755), .A(n15662), .B(n15661), .ZN(
        P2_U3222) );
  NAND2_X1 U17271 ( .A1(n15665), .A2(n15664), .ZN(n15666) );
  NAND2_X1 U17272 ( .A1(n15667), .A2(n15666), .ZN(n15668) );
  NAND2_X1 U17273 ( .A1(n15744), .A2(n15668), .ZN(n15675) );
  NAND2_X1 U17274 ( .A1(n15670), .A2(n15669), .ZN(n15671) );
  NAND2_X1 U17275 ( .A1(n15672), .A2(n15671), .ZN(n15673) );
  NAND2_X1 U17276 ( .A1(n15752), .A2(n15673), .ZN(n15674) );
  OAI211_X1 U17277 ( .C1(n15749), .C2(n15676), .A(n15675), .B(n15674), .ZN(
        n15677) );
  INV_X1 U17278 ( .A(n15677), .ZN(n15679) );
  OAI211_X1 U17279 ( .C1(n9744), .C2(n15755), .A(n15679), .B(n15678), .ZN(
        P2_U3223) );
  INV_X1 U17280 ( .A(n15680), .ZN(n15681) );
  AOI211_X1 U17281 ( .C1(n15684), .C2(n15683), .A(n15682), .B(n15681), .ZN(
        n15689) );
  AOI211_X1 U17282 ( .C1(n15687), .C2(n15686), .A(n15733), .B(n15685), .ZN(
        n15688) );
  AOI211_X1 U17283 ( .C1(n15739), .C2(n15690), .A(n15689), .B(n15688), .ZN(
        n15692) );
  OAI211_X1 U17284 ( .C1(n15693), .C2(n15755), .A(n15692), .B(n15691), .ZN(
        P2_U3224) );
  OAI21_X1 U17285 ( .B1(n15696), .B2(n15695), .A(n15694), .ZN(n15702) );
  OAI21_X1 U17286 ( .B1(n15699), .B2(n15698), .A(n15697), .ZN(n15700) );
  AOI222_X1 U17287 ( .A1(n15702), .A2(n15752), .B1(n15701), .B2(n15739), .C1(
        n15700), .C2(n15744), .ZN(n15704) );
  OAI211_X1 U17288 ( .C1(n15705), .C2(n15755), .A(n15704), .B(n15703), .ZN(
        P2_U3226) );
  OAI211_X1 U17289 ( .C1(n15707), .C2(P2_REG2_REG_14__SCAN_IN), .A(n15706), 
        .B(n15752), .ZN(n15708) );
  INV_X1 U17290 ( .A(n15708), .ZN(n15712) );
  AOI211_X1 U17291 ( .C1(n15710), .C2(n15709), .A(n15733), .B(n6704), .ZN(
        n15711) );
  AOI211_X1 U17292 ( .C1(n15739), .C2(n15713), .A(n15712), .B(n15711), .ZN(
        n15715) );
  OAI211_X1 U17293 ( .C1(n9755), .C2(n15755), .A(n15715), .B(n15714), .ZN(
        P2_U3228) );
  INV_X1 U17294 ( .A(n15716), .ZN(n15717) );
  OAI211_X1 U17295 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n15718), .A(n15717), 
        .B(n15744), .ZN(n15722) );
  OAI211_X1 U17296 ( .C1(n15720), .C2(P2_REG2_REG_15__SCAN_IN), .A(n15719), 
        .B(n15752), .ZN(n15721) );
  OAI211_X1 U17297 ( .C1(n15749), .C2(n15723), .A(n15722), .B(n15721), .ZN(
        n15724) );
  INV_X1 U17298 ( .A(n15724), .ZN(n15726) );
  NAND2_X1 U17299 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(n11242), .ZN(n15725) );
  OAI211_X1 U17300 ( .C1(n15727), .C2(n15755), .A(n15726), .B(n15725), .ZN(
        P2_U3229) );
  OAI211_X1 U17301 ( .C1(n15730), .C2(n15729), .A(n15728), .B(n15752), .ZN(
        n15731) );
  INV_X1 U17302 ( .A(n15731), .ZN(n15737) );
  AOI211_X1 U17303 ( .C1(n15735), .C2(n15734), .A(n15733), .B(n15732), .ZN(
        n15736) );
  AOI211_X1 U17304 ( .C1(n15739), .C2(n15738), .A(n15737), .B(n15736), .ZN(
        n15741) );
  OAI211_X1 U17305 ( .C1(n15742), .C2(n15755), .A(n15741), .B(n15740), .ZN(
        P2_U3230) );
  XNOR2_X1 U17306 ( .A(n15743), .B(n14345), .ZN(n15751) );
  OAI211_X1 U17307 ( .C1(n15746), .C2(P2_REG1_REG_18__SCAN_IN), .A(n15745), 
        .B(n15744), .ZN(n15747) );
  OAI21_X1 U17308 ( .B1(n15749), .B2(n15748), .A(n15747), .ZN(n15750) );
  AOI21_X1 U17309 ( .B1(n15752), .B2(n15751), .A(n15750), .ZN(n15754) );
  OAI211_X1 U17310 ( .C1(n15756), .C2(n15755), .A(n15754), .B(n15753), .ZN(
        P2_U3232) );
  XNOR2_X1 U17311 ( .A(n15757), .B(n15765), .ZN(n15760) );
  AOI21_X1 U17312 ( .B1(n15760), .B2(n15759), .A(n15758), .ZN(n15825) );
  AOI222_X1 U17313 ( .A1(n15764), .A2(n15763), .B1(P2_REG2_REG_6__SCAN_IN), 
        .B2(n15783), .C1(n15762), .C2(n15761), .ZN(n15773) );
  XNOR2_X1 U17314 ( .A(n15766), .B(n15765), .ZN(n15828) );
  INV_X1 U17315 ( .A(n11936), .ZN(n15768) );
  OAI211_X1 U17316 ( .C1(n15824), .C2(n11797), .A(n15768), .B(n15767), .ZN(
        n15823) );
  INV_X1 U17317 ( .A(n15823), .ZN(n15769) );
  AOI22_X1 U17318 ( .A1(n15828), .A2(n15771), .B1(n15770), .B2(n15769), .ZN(
        n15772) );
  OAI211_X1 U17319 ( .C1(n15783), .C2(n15825), .A(n15773), .B(n15772), .ZN(
        P2_U3259) );
  INV_X1 U17320 ( .A(n15774), .ZN(n15779) );
  OAI22_X1 U17321 ( .A1(n15776), .A2(n7270), .B1(n11791), .B2(n15775), .ZN(
        n15778) );
  AOI211_X1 U17322 ( .C1(n15780), .C2(n15779), .A(n15778), .B(n15777), .ZN(
        n15782) );
  AOI22_X1 U17323 ( .A1(n15783), .A2(n11287), .B1(n15782), .B2(n15781), .ZN(
        P2_U3265) );
  AND2_X1 U17324 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15790), .ZN(P2_U3266) );
  AND2_X1 U17325 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15790), .ZN(P2_U3267) );
  AND2_X1 U17326 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15790), .ZN(P2_U3268) );
  AND2_X1 U17327 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15790), .ZN(P2_U3269) );
  AND2_X1 U17328 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15790), .ZN(P2_U3270) );
  NOR2_X1 U17329 ( .A1(n15789), .A2(n15785), .ZN(P2_U3271) );
  AND2_X1 U17330 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15790), .ZN(P2_U3272) );
  NOR2_X1 U17331 ( .A1(n15789), .A2(n15786), .ZN(P2_U3273) );
  AND2_X1 U17332 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15790), .ZN(P2_U3274) );
  AND2_X1 U17333 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15790), .ZN(P2_U3275) );
  AND2_X1 U17334 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15790), .ZN(P2_U3276) );
  AND2_X1 U17335 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15790), .ZN(P2_U3277) );
  AND2_X1 U17336 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15790), .ZN(P2_U3278) );
  AND2_X1 U17337 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15790), .ZN(P2_U3279) );
  AND2_X1 U17338 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15790), .ZN(P2_U3280) );
  AND2_X1 U17339 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15790), .ZN(P2_U3281) );
  NOR2_X1 U17340 ( .A1(n15789), .A2(n15787), .ZN(P2_U3282) );
  AND2_X1 U17341 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15790), .ZN(P2_U3283) );
  AND2_X1 U17342 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15790), .ZN(P2_U3284) );
  AND2_X1 U17343 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15790), .ZN(P2_U3285) );
  AND2_X1 U17344 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15790), .ZN(P2_U3286) );
  AND2_X1 U17345 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15790), .ZN(P2_U3287) );
  AND2_X1 U17346 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15790), .ZN(P2_U3288) );
  AND2_X1 U17347 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15790), .ZN(P2_U3289) );
  AND2_X1 U17348 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15790), .ZN(P2_U3290) );
  AND2_X1 U17349 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15790), .ZN(P2_U3291) );
  NOR2_X1 U17350 ( .A1(n15789), .A2(n15788), .ZN(P2_U3292) );
  AND2_X1 U17351 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15790), .ZN(P2_U3293) );
  AND2_X1 U17352 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15790), .ZN(P2_U3294) );
  AND2_X1 U17353 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15790), .ZN(P2_U3295) );
  AOI22_X1 U17354 ( .A1(n15796), .A2(n15792), .B1(n15791), .B2(n15793), .ZN(
        P2_U3416) );
  AOI22_X1 U17355 ( .A1(n15796), .A2(n15795), .B1(n15794), .B2(n15793), .ZN(
        P2_U3417) );
  INV_X1 U17356 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15797) );
  AOI22_X1 U17357 ( .A1(n15838), .A2(n15798), .B1(n15797), .B2(n7304), .ZN(
        P2_U3430) );
  OAI21_X1 U17358 ( .B1(n15800), .B2(n15831), .A(n15799), .ZN(n15802) );
  AOI211_X1 U17359 ( .C1(n15835), .C2(n15803), .A(n15802), .B(n15801), .ZN(
        n15839) );
  AOI22_X1 U17360 ( .A1(n15838), .A2(n15839), .B1(n15804), .B2(n7304), .ZN(
        P2_U3436) );
  OAI21_X1 U17361 ( .B1(n15806), .B2(n15831), .A(n15805), .ZN(n15808) );
  AOI211_X1 U17362 ( .C1(n15810), .C2(n15809), .A(n15808), .B(n15807), .ZN(
        n15841) );
  AOI22_X1 U17363 ( .A1(n15838), .A2(n15841), .B1(n15811), .B2(n7304), .ZN(
        P2_U3442) );
  NAND2_X1 U17364 ( .A1(n15813), .A2(n15812), .ZN(n15816) );
  INV_X1 U17365 ( .A(n15814), .ZN(n15815) );
  OAI211_X1 U17366 ( .C1(n15818), .C2(n15817), .A(n15816), .B(n15815), .ZN(
        n15819) );
  INV_X1 U17367 ( .A(n15819), .ZN(n15820) );
  AND2_X1 U17368 ( .A1(n15821), .A2(n15820), .ZN(n15843) );
  INV_X1 U17369 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15822) );
  AOI22_X1 U17370 ( .A1(n15838), .A2(n15843), .B1(n15822), .B2(n7304), .ZN(
        P2_U3445) );
  OAI21_X1 U17371 ( .B1(n15824), .B2(n15831), .A(n15823), .ZN(n15827) );
  INV_X1 U17372 ( .A(n15825), .ZN(n15826) );
  AOI211_X1 U17373 ( .C1(n15828), .C2(n15835), .A(n15827), .B(n15826), .ZN(
        n15845) );
  INV_X1 U17374 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15829) );
  AOI22_X1 U17375 ( .A1(n15838), .A2(n15845), .B1(n15829), .B2(n7304), .ZN(
        P2_U3448) );
  OAI21_X1 U17376 ( .B1(n7911), .B2(n15831), .A(n15830), .ZN(n15834) );
  INV_X1 U17377 ( .A(n15832), .ZN(n15833) );
  AOI211_X1 U17378 ( .C1(n15836), .C2(n15835), .A(n15834), .B(n15833), .ZN(
        n15847) );
  INV_X1 U17379 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15837) );
  AOI22_X1 U17380 ( .A1(n15838), .A2(n15847), .B1(n15837), .B2(n7304), .ZN(
        P2_U3451) );
  AOI22_X1 U17381 ( .A1(n15848), .A2(n15839), .B1(n10380), .B2(n7285), .ZN(
        P2_U3501) );
  AOI22_X1 U17382 ( .A1(n15848), .A2(n15841), .B1(n15840), .B2(n7285), .ZN(
        P2_U3503) );
  AOI22_X1 U17383 ( .A1(n15848), .A2(n15843), .B1(n15842), .B2(n7285), .ZN(
        P2_U3504) );
  AOI22_X1 U17384 ( .A1(n15848), .A2(n15845), .B1(n15844), .B2(n7285), .ZN(
        P2_U3505) );
  AOI22_X1 U17385 ( .A1(n15848), .A2(n15847), .B1(n15846), .B2(n7285), .ZN(
        P2_U3506) );
  NOR2_X1 U17386 ( .A1(P3_U3897), .A2(n15849), .ZN(P3_U3150) );
  INV_X1 U17387 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15872) );
  INV_X1 U17388 ( .A(n15850), .ZN(n15869) );
  XNOR2_X1 U17389 ( .A(n15851), .B(n15857), .ZN(n15867) );
  INV_X1 U17390 ( .A(n15867), .ZN(n15880) );
  NOR2_X1 U17391 ( .A1(n15901), .A2(n15852), .ZN(n15878) );
  INV_X1 U17392 ( .A(n15878), .ZN(n15854) );
  OAI22_X1 U17393 ( .A1(n15856), .A2(n15855), .B1(n15854), .B2(n15853), .ZN(
        n15868) );
  XNOR2_X1 U17394 ( .A(n15857), .B(n15858), .ZN(n15863) );
  OAI22_X1 U17395 ( .A1(n15861), .A2(n15860), .B1(n7251), .B2(n15859), .ZN(
        n15862) );
  AOI21_X1 U17396 ( .B1(n15864), .B2(n15863), .A(n15862), .ZN(n15865) );
  OAI21_X1 U17397 ( .B1(n15867), .B2(n15866), .A(n15865), .ZN(n15877) );
  AOI211_X1 U17398 ( .C1(n15869), .C2(n15880), .A(n15868), .B(n15877), .ZN(
        n15871) );
  AOI22_X1 U17399 ( .A1(n15873), .A2(n15872), .B1(n15871), .B2(n15870), .ZN(
        P3_U3231) );
  AOI211_X1 U17400 ( .C1(n15899), .C2(n15876), .A(n15875), .B(n15874), .ZN(
        n15908) );
  AOI22_X1 U17401 ( .A1(n15906), .A2(n12452), .B1(n15908), .B2(n15905), .ZN(
        P3_U3393) );
  AOI211_X1 U17402 ( .C1(n15880), .C2(n15879), .A(n15878), .B(n15877), .ZN(
        n15909) );
  AOI22_X1 U17403 ( .A1(n15906), .A2(n9040), .B1(n15909), .B2(n15905), .ZN(
        P3_U3396) );
  OAI22_X1 U17404 ( .A1(n15882), .A2(n15886), .B1(n15881), .B2(n15901), .ZN(
        n15883) );
  NOR2_X1 U17405 ( .A1(n15884), .A2(n15883), .ZN(n15911) );
  AOI22_X1 U17406 ( .A1(n15906), .A2(n9057), .B1(n15911), .B2(n15905), .ZN(
        P3_U3399) );
  OAI22_X1 U17407 ( .A1(n15887), .A2(n15886), .B1(n15885), .B2(n15901), .ZN(
        n15888) );
  NOR2_X1 U17408 ( .A1(n15889), .A2(n15888), .ZN(n15912) );
  AOI22_X1 U17409 ( .A1(n15906), .A2(n9077), .B1(n15912), .B2(n15905), .ZN(
        P3_U3402) );
  INV_X1 U17410 ( .A(n15890), .ZN(n15894) );
  OAI21_X1 U17411 ( .B1(n15892), .B2(n15901), .A(n15891), .ZN(n15893) );
  AOI21_X1 U17412 ( .B1(n15894), .B2(n15899), .A(n15893), .ZN(n15914) );
  AOI22_X1 U17413 ( .A1(n15906), .A2(n9090), .B1(n15914), .B2(n15905), .ZN(
        P3_U3405) );
  OAI21_X1 U17414 ( .B1(n15896), .B2(n15901), .A(n15895), .ZN(n15897) );
  AOI21_X1 U17415 ( .B1(n15898), .B2(n15899), .A(n15897), .ZN(n15916) );
  AOI22_X1 U17416 ( .A1(n15906), .A2(n9111), .B1(n15916), .B2(n15905), .ZN(
        P3_U3408) );
  AND2_X1 U17417 ( .A1(n15900), .A2(n15899), .ZN(n15903) );
  NOR2_X1 U17418 ( .A1(n15901), .A2(n6956), .ZN(n15902) );
  NOR3_X1 U17419 ( .A1(n15904), .A2(n15903), .A3(n15902), .ZN(n15917) );
  AOI22_X1 U17420 ( .A1(n15906), .A2(n9130), .B1(n15917), .B2(n15905), .ZN(
        P3_U3411) );
  INV_X1 U17421 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15907) );
  AOI22_X1 U17422 ( .A1(n15918), .A2(n15908), .B1(n15907), .B2(n10706), .ZN(
        P3_U3460) );
  AOI22_X1 U17423 ( .A1(n15918), .A2(n15909), .B1(n9619), .B2(n10706), .ZN(
        P3_U3461) );
  AOI22_X1 U17424 ( .A1(n15918), .A2(n15911), .B1(n15910), .B2(n10706), .ZN(
        P3_U3462) );
  AOI22_X1 U17425 ( .A1(n15918), .A2(n15912), .B1(n9073), .B2(n10706), .ZN(
        P3_U3463) );
  AOI22_X1 U17426 ( .A1(n15918), .A2(n15914), .B1(n15913), .B2(n10706), .ZN(
        P3_U3464) );
  AOI22_X1 U17427 ( .A1(n15918), .A2(n15916), .B1(n15915), .B2(n10706), .ZN(
        P3_U3465) );
  AOI22_X1 U17428 ( .A1(n15918), .A2(n15917), .B1(n9648), .B2(n10706), .ZN(
        P3_U3466) );
  AOI21_X1 U17429 ( .B1(n15920), .B2(n15919), .A(n6724), .ZN(SUB_1596_U59) );
  OAI21_X1 U17430 ( .B1(n15923), .B2(n15922), .A(n15921), .ZN(SUB_1596_U58) );
  XOR2_X1 U17431 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15924), .Z(SUB_1596_U53) );
  AOI21_X1 U17432 ( .B1(n15927), .B2(n15926), .A(n15925), .ZN(SUB_1596_U56) );
  AOI21_X1 U17433 ( .B1(n15930), .B2(n15929), .A(n15928), .ZN(n15931) );
  XOR2_X1 U17434 ( .A(n15931), .B(P2_ADDR_REG_3__SCAN_IN), .Z(SUB_1596_U60) );
  AOI21_X1 U17435 ( .B1(n15934), .B2(n15933), .A(n15932), .ZN(SUB_1596_U5) );
  INV_X1 U7308 ( .A(n10381), .ZN(n10373) );
  INV_X1 U7265 ( .A(n10381), .ZN(n13970) );
  CLKBUF_X1 U7274 ( .A(n6560), .Z(n13892) );
  NAND2_X1 U7281 ( .A1(n10724), .A2(n7750), .ZN(n9953) );
  CLKBUF_X1 U7284 ( .A(n8261), .Z(n8780) );
  CLKBUF_X1 U7301 ( .A(n8282), .Z(n8776) );
  CLKBUF_X1 U7316 ( .A(n9069), .Z(n7381) );
  INV_X1 U7320 ( .A(n10643), .ZN(n6512) );
  CLKBUF_X1 U7447 ( .A(n13969), .Z(n7281) );
  CLKBUF_X1 U7590 ( .A(n10586), .Z(n13819) );
  CLKBUF_X1 U9411 ( .A(n10316), .Z(n14077) );
endmodule

