

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput127,
         keyinput126, keyinput125, keyinput124, keyinput123, keyinput122,
         keyinput121, keyinput120, keyinput119, keyinput118, keyinput117,
         keyinput116, keyinput115, keyinput114, keyinput113, keyinput112,
         keyinput111, keyinput110, keyinput109, keyinput108, keyinput107,
         keyinput106, keyinput105, keyinput104, keyinput103, keyinput102,
         keyinput101, keyinput100, keyinput99, keyinput98, keyinput97,
         keyinput96, keyinput95, keyinput94, keyinput93, keyinput92,
         keyinput91, keyinput90, keyinput89, keyinput88, keyinput87,
         keyinput86, keyinput85, keyinput84, keyinput83, keyinput82,
         keyinput81, keyinput80, keyinput79, keyinput78, keyinput77,
         keyinput76, keyinput75, keyinput74, keyinput73, keyinput72,
         keyinput71, keyinput70, keyinput69, keyinput68, keyinput67,
         keyinput66, keyinput65, keyinput64, keyinput63, keyinput62,
         keyinput61, keyinput60, keyinput59, keyinput58, keyinput57,
         keyinput56, keyinput55, keyinput54, keyinput53, keyinput52,
         keyinput51, keyinput50, keyinput49, keyinput48, keyinput47,
         keyinput46, keyinput45, keyinput44, keyinput43, keyinput42,
         keyinput41, keyinput40, keyinput39, keyinput38, keyinput37,
         keyinput36, keyinput35, keyinput34, keyinput33, keyinput32,
         keyinput31, keyinput30, keyinput29, keyinput28, keyinput27,
         keyinput26, keyinput25, keyinput24, keyinput23, keyinput22,
         keyinput21, keyinput20, keyinput19, keyinput18, keyinput17,
         keyinput16, keyinput15, keyinput14, keyinput13, keyinput12,
         keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6,
         keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748;

  NOR2_X1 U7293 ( .A1(n12961), .A2(n12962), .ZN(n12965) );
  NOR2_X1 U7294 ( .A1(n15480), .A2(n12942), .ZN(n12961) );
  NAND2_X1 U7295 ( .A1(n8518), .A2(n8517), .ZN(n13860) );
  INV_X4 U7296 ( .A(n8097), .ZN(n8285) );
  INV_X1 U7297 ( .A(n10731), .ZN(n10405) );
  CLKBUF_X2 U7298 ( .A(n10283), .Z(n10301) );
  INV_X1 U7299 ( .A(n15014), .ZN(n11131) );
  CLKBUF_X1 U7300 ( .A(n9218), .Z(n6547) );
  NAND2_X1 U7301 ( .A1(n7807), .A2(n7806), .ZN(n12043) );
  XNOR2_X1 U7302 ( .A(n8648), .B(n13380), .ZN(n12657) );
  NAND2_X1 U7303 ( .A1(n8148), .A2(n10491), .ZN(n7806) );
  CLKBUF_X1 U7304 ( .A(n12068), .Z(n6553) );
  NAND2_X2 U7305 ( .A1(n8126), .A2(n7997), .ZN(n8133) );
  BUF_X4 U7306 ( .A(n10275), .Z(n6549) );
  XNOR2_X1 U7307 ( .A(n9841), .B(n9840), .ZN(n14235) );
  NAND2_X1 U7308 ( .A1(n7212), .A2(n7210), .ZN(n14629) );
  XNOR2_X1 U7309 ( .A(n9821), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9826) );
  AND2_X1 U7310 ( .A1(n9820), .A2(n9819), .ZN(n6868) );
  INV_X2 U7311 ( .A(n8004), .ZN(n8013) );
  NOR2_X1 U7312 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n9805) );
  INV_X4 U7313 ( .A(n14498), .ZN(n6550) );
  NOR2_X1 U7314 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n9803) );
  AND4_X1 U7315 ( .A1(n9806), .A2(n9805), .A3(n9804), .A4(n9803), .ZN(n9809)
         );
  NOR2_X1 U7316 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n10026) );
  INV_X2 U7318 ( .A(n10283), .ZN(n10216) );
  NAND2_X1 U7319 ( .A1(n14640), .A2(n14235), .ZN(n10709) );
  INV_X2 U7320 ( .A(n11571), .ZN(n12640) );
  NAND2_X1 U7321 ( .A1(n11285), .A2(n11393), .ZN(n9267) );
  NAND2_X2 U7322 ( .A1(n9267), .A2(n9266), .ZN(n11386) );
  OR2_X1 U7323 ( .A1(n8987), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8988) );
  NOR2_X1 U7324 ( .A1(n12068), .A2(n9791), .ZN(n12066) );
  INV_X1 U7325 ( .A(n12777), .ZN(n12746) );
  AND2_X1 U7326 ( .A1(n9826), .A2(n14626), .ZN(n10275) );
  CLKBUF_X2 U7327 ( .A(n9867), .Z(n10237) );
  INV_X1 U7328 ( .A(n10083), .ZN(n9837) );
  BUF_X1 U7329 ( .A(n10083), .Z(n10084) );
  INV_X1 U7330 ( .A(n11383), .ZN(n11571) );
  NAND2_X1 U7331 ( .A1(n7076), .A2(n7077), .ZN(n12624) );
  NOR2_X1 U7332 ( .A1(n12941), .A2(n7477), .ZN(n12960) );
  NOR2_X1 U7333 ( .A1(n12969), .A2(n7187), .ZN(n12972) );
  INV_X1 U7334 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8660) );
  INV_X1 U7335 ( .A(n8133), .ZN(n9624) );
  AND2_X1 U7336 ( .A1(n6997), .A2(n7633), .ZN(n6651) );
  AND3_X1 U7337 ( .A1(n6577), .A2(n7007), .A3(n6676), .ZN(n11781) );
  XNOR2_X1 U7338 ( .A(n12624), .B(n12625), .ZN(n12869) );
  NAND2_X1 U7339 ( .A1(n8354), .A2(n8353), .ZN(n14847) );
  NAND2_X1 U7340 ( .A1(n8257), .A2(n8256), .ZN(n15252) );
  INV_X2 U7341 ( .A(n8013), .ZN(n10486) );
  OAI21_X1 U7342 ( .B1(n12751), .B2(n12750), .A(n12752), .ZN(n14034) );
  NAND2_X1 U7343 ( .A1(n12680), .A2(n6934), .ZN(n14083) );
  INV_X1 U7344 ( .A(n10260), .ZN(n9927) );
  INV_X1 U7345 ( .A(n10179), .ZN(n10278) );
  INV_X1 U7346 ( .A(n8004), .ZN(n7997) );
  AOI22_X1 U7347 ( .A1(n13381), .A2(n9234), .B1(n9216), .B2(SI_31_), .ZN(
        n13257) );
  NAND4_X1 U7349 ( .A1(n8171), .A2(n8170), .A3(n8169), .A4(n8168), .ZN(n13523)
         );
  NAND2_X1 U7350 ( .A1(n6869), .A2(n6863), .ZN(n10373) );
  XNOR2_X1 U7351 ( .A(n9838), .B(P1_IR_REG_22__SCAN_IN), .ZN(n14640) );
  INV_X1 U7352 ( .A(n12902), .ZN(P3_U3897) );
  XNOR2_X1 U7353 ( .A(n8682), .B(n8681), .ZN(n14753) );
  INV_X1 U7355 ( .A(n8013), .ZN(n6546) );
  INV_X2 U7357 ( .A(n8013), .ZN(n10485) );
  NOR2_X2 U7358 ( .A1(n10875), .A2(n11090), .ZN(n11089) );
  OAI211_X2 U7359 ( .C1(n10287), .C2(n10288), .A(n10286), .B(n10285), .ZN(
        n7226) );
  NAND2_X1 U7360 ( .A1(n12657), .A2(n8651), .ZN(n9218) );
  AOI21_X2 U7361 ( .B1(n7372), .B2(n8694), .A(n6606), .ZN(n7376) );
  AND2_X4 U7362 ( .A1(n13388), .A2(n12657), .ZN(n8702) );
  NOR2_X2 U7363 ( .A1(n10956), .A2(n10957), .ZN(n10771) );
  OAI21_X2 U7365 ( .B1(n7641), .B2(n7000), .A(n6651), .ZN(n13466) );
  NAND2_X2 U7366 ( .A1(n8384), .A2(n7645), .ZN(n7641) );
  NOR2_X2 U7367 ( .A1(n14766), .A2(n14703), .ZN(n14706) );
  XNOR2_X1 U7369 ( .A(n12476), .B(n14099), .ZN(n12032) );
  INV_X1 U7370 ( .A(n6781), .ZN(n10758) );
  OAI211_X2 U7371 ( .C1(n8669), .C2(n7689), .A(n7688), .B(n7687), .ZN(n6781)
         );
  OR3_X1 U7372 ( .A1(n9701), .A2(n12403), .A3(n9661), .ZN(n9704) );
  AOI21_X1 U7373 ( .B1(n9658), .B2(n6813), .A(n9657), .ZN(n6812) );
  AOI21_X1 U7374 ( .B1(n9581), .B2(n9577), .A(n9579), .ZN(n6813) );
  OR2_X1 U7375 ( .A1(n9793), .A2(n6909), .ZN(n6907) );
  OAI21_X1 U7376 ( .B1(n13981), .B2(n6950), .A(n6947), .ZN(n14071) );
  NAND2_X1 U7377 ( .A1(n14309), .A2(n6617), .ZN(n14299) );
  NAND2_X1 U7378 ( .A1(n14311), .A2(n14310), .ZN(n14309) );
  AND2_X1 U7379 ( .A1(n7753), .A2(n7752), .ZN(n12609) );
  AOI21_X1 U7380 ( .B1(n15251), .B2(n13843), .A(n13842), .ZN(n13844) );
  AND2_X1 U7381 ( .A1(n13617), .A2(n13616), .ZN(n13842) );
  NOR2_X1 U7382 ( .A1(n13981), .A2(n12742), .ZN(n14035) );
  NAND2_X1 U7383 ( .A1(n7012), .A2(n7014), .ZN(n13483) );
  AOI21_X2 U7384 ( .B1(n14050), .B2(n13979), .A(n13978), .ZN(n13981) );
  NOR2_X1 U7385 ( .A1(n7332), .A2(n14332), .ZN(n7159) );
  AOI21_X1 U7386 ( .B1(n6571), .B2(n12916), .A(n6766), .ZN(n6765) );
  CLKBUF_X1 U7387 ( .A(n12563), .Z(n7109) );
  NAND2_X1 U7388 ( .A1(n9775), .A2(n9774), .ZN(n13727) );
  NAND2_X1 U7389 ( .A1(n14390), .A2(n12561), .ZN(n14372) );
  NAND2_X1 U7390 ( .A1(n10209), .A2(n10208), .ZN(n14334) );
  OR2_X1 U7391 ( .A1(n7825), .A2(n14026), .ZN(n6574) );
  OR2_X1 U7392 ( .A1(n12864), .A2(n7421), .ZN(n7076) );
  NAND2_X1 U7393 ( .A1(n6873), .A2(n7472), .ZN(n14342) );
  NAND2_X1 U7394 ( .A1(n10203), .A2(n10202), .ZN(n14352) );
  OR2_X1 U7395 ( .A1(n12682), .A2(n12681), .ZN(n6934) );
  NAND2_X1 U7396 ( .A1(n8472), .A2(n8471), .ZN(n13875) );
  OR2_X1 U7397 ( .A1(n12845), .A2(n7095), .ZN(n7093) );
  NAND2_X1 U7398 ( .A1(n7129), .A2(n6979), .ZN(n6978) );
  NAND2_X1 U7399 ( .A1(n6954), .A2(n7838), .ZN(n12666) );
  NAND2_X1 U7400 ( .A1(n12441), .A2(n7130), .ZN(n7129) );
  AND2_X1 U7401 ( .A1(n6778), .A2(n6674), .ZN(n12921) );
  NAND2_X1 U7402 ( .A1(n14876), .A2(n7839), .ZN(n6954) );
  NOR2_X1 U7403 ( .A1(n7640), .A2(n8404), .ZN(n7639) );
  XNOR2_X1 U7404 ( .A(n8987), .B(n15645), .ZN(n8986) );
  NAND2_X1 U7405 ( .A1(n6977), .A2(n7794), .ZN(n12229) );
  NAND2_X1 U7406 ( .A1(n7843), .A2(n7849), .ZN(n7838) );
  NOR2_X1 U7407 ( .A1(n7841), .A2(n7840), .ZN(n7839) );
  NAND2_X1 U7408 ( .A1(n7116), .A2(n14097), .ZN(n12552) );
  OR3_X1 U7409 ( .A1(n9478), .A2(n9477), .A3(n7254), .ZN(n7253) );
  NAND2_X1 U7410 ( .A1(n6806), .A2(n6808), .ZN(n8087) );
  AOI22_X1 U7411 ( .A1(n12092), .A2(n9717), .B1(n15264), .B2(n13517), .ZN(
        n12120) );
  AND2_X1 U7412 ( .A1(n7486), .A2(n7485), .ZN(n12910) );
  NAND2_X1 U7413 ( .A1(n8448), .A2(n8447), .ZN(n13893) );
  NAND2_X1 U7414 ( .A1(n6807), .A2(n8452), .ZN(n6806) );
  XNOR2_X1 U7415 ( .A(n8369), .B(n8368), .ZN(n11237) );
  AOI21_X1 U7416 ( .B1(n8049), .B2(n7765), .A(n7764), .ZN(n7763) );
  OAI211_X1 U7417 ( .C1(n11870), .C2(n6960), .A(n6959), .B(n6697), .ZN(n7206)
         );
  NAND2_X1 U7418 ( .A1(n10068), .A2(n10067), .ZN(n12499) );
  NAND2_X1 U7419 ( .A1(n14770), .A2(n10601), .ZN(n14769) );
  NAND2_X1 U7420 ( .A1(n7152), .A2(n8035), .ZN(n8367) );
  NAND2_X1 U7421 ( .A1(n10052), .A2(n10051), .ZN(n12476) );
  NAND2_X1 U7422 ( .A1(n8392), .A2(n8391), .ZN(n13907) );
  NOR2_X1 U7423 ( .A1(n15741), .A2(n14707), .ZN(n14710) );
  NAND2_X1 U7424 ( .A1(n8366), .A2(n8347), .ZN(n8349) );
  NAND2_X1 U7425 ( .A1(n8276), .A2(n8275), .ZN(n12102) );
  AND2_X1 U7426 ( .A1(n6835), .A2(n6834), .ZN(n11864) );
  NAND2_X1 U7427 ( .A1(n7047), .A2(n10016), .ZN(n14870) );
  XNOR2_X1 U7428 ( .A(n8310), .B(n8309), .ZN(n10615) );
  NAND2_X1 U7429 ( .A1(n10031), .A2(n10030), .ZN(n14892) );
  OR2_X1 U7430 ( .A1(n8346), .A2(n10618), .ZN(n8366) );
  AND2_X1 U7431 ( .A1(n8872), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7008) );
  NOR2_X1 U7432 ( .A1(n11058), .A2(n11059), .ZN(n11061) );
  NAND2_X1 U7433 ( .A1(n9923), .A2(n9922), .ZN(n11587) );
  INV_X8 U7434 ( .A(n12779), .ZN(n12743) );
  NAND2_X1 U7435 ( .A1(n8164), .A2(n8163), .ZN(n15227) );
  NAND2_X2 U7436 ( .A1(n9903), .A2(n11133), .ZN(n12779) );
  NOR2_X1 U7437 ( .A1(n13527), .A2(n8105), .ZN(n9426) );
  BUF_X2 U7438 ( .A(P1_U4016), .Z(n6551) );
  INV_X2 U7439 ( .A(n14494), .ZN(n11143) );
  INV_X2 U7440 ( .A(n11440), .ZN(n7324) );
  INV_X2 U7441 ( .A(n15344), .ZN(n11285) );
  NAND2_X1 U7442 ( .A1(n6648), .A2(n9883), .ZN(n14110) );
  INV_X1 U7443 ( .A(n14109), .ZN(n11338) );
  NAND2_X1 U7444 ( .A1(n10370), .A2(n10369), .ZN(n11133) );
  NAND3_X1 U7445 ( .A1(n8101), .A2(n8100), .A3(n8099), .ZN(n13527) );
  OR2_X1 U7446 ( .A1(n10898), .A2(n10897), .ZN(n10924) );
  NAND2_X1 U7447 ( .A1(n9870), .A2(n9869), .ZN(n14933) );
  INV_X1 U7448 ( .A(n14108), .ZN(n11479) );
  CLKBUF_X2 U7450 ( .A(n8134), .Z(n6557) );
  NAND2_X1 U7451 ( .A1(n7740), .A2(n8007), .ZN(n8159) );
  INV_X2 U7452 ( .A(n9610), .ZN(n8148) );
  BUF_X2 U7453 ( .A(n9653), .Z(n9578) );
  NAND4_X1 U7454 ( .A1(n9860), .A2(n9859), .A3(n9858), .A4(n9857), .ZN(n14108)
         );
  INV_X2 U7455 ( .A(n8136), .ZN(n9613) );
  CLKBUF_X2 U7456 ( .A(n8126), .Z(n7128) );
  NAND2_X1 U7457 ( .A1(n9092), .A2(n9097), .ZN(n11687) );
  INV_X2 U7458 ( .A(n9653), .ZN(n6552) );
  XNOR2_X1 U7459 ( .A(n7660), .B(n14692), .ZN(n15745) );
  OAI21_X1 U7460 ( .B1(n10362), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10361) );
  OR2_X2 U7461 ( .A1(n10705), .A2(n10700), .ZN(n15014) );
  NAND2_X1 U7462 ( .A1(n13949), .A2(n7975), .ZN(n8136) );
  INV_X1 U7463 ( .A(n8603), .ZN(n9698) );
  NAND2_X1 U7464 ( .A1(n7973), .A2(n7972), .ZN(n13949) );
  NAND2_X2 U7465 ( .A1(n10709), .A2(n11132), .ZN(n12777) );
  XNOR2_X1 U7466 ( .A(n7987), .B(P2_IR_REG_22__SCAN_IN), .ZN(n9667) );
  INV_X1 U7467 ( .A(n9826), .ZN(n14623) );
  AND2_X2 U7468 ( .A1(n9826), .A2(n9825), .ZN(n10179) );
  OR2_X2 U7469 ( .A1(n12657), .A2(n8651), .ZN(n8699) );
  CLKBUF_X2 U7470 ( .A(n8603), .Z(n6555) );
  INV_X1 U7471 ( .A(n7907), .ZN(n7975) );
  NAND2_X1 U7474 ( .A1(n7971), .A2(n7970), .ZN(n7973) );
  NAND2_X1 U7475 ( .A1(n13385), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8648) );
  XNOR2_X1 U7476 ( .A(n6913), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7907) );
  NAND2_X1 U7477 ( .A1(n9816), .A2(n7146), .ZN(n7212) );
  OAI21_X1 U7478 ( .B1(n8311), .B2(n8083), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8085) );
  AND2_X1 U7479 ( .A1(n10961), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10963) );
  NAND2_X2 U7480 ( .A1(n10485), .A2(P1_U3086), .ZN(n14635) );
  OAI21_X1 U7481 ( .B1(n9839), .B2(n7859), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9838) );
  OAI21_X1 U7482 ( .B1(n8004), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n7995), .ZN(
        n7999) );
  NOR2_X1 U7483 ( .A1(n9147), .A2(n7900), .ZN(n8656) );
  AND3_X2 U7484 ( .A1(n7965), .A2(n7964), .A3(n8082), .ZN(n7986) );
  NAND3_X1 U7485 ( .A1(n9920), .A2(n9809), .A3(n9808), .ZN(n10083) );
  AND3_X1 U7486 ( .A1(n7963), .A2(n7962), .A3(n7961), .ZN(n8082) );
  NAND2_X1 U7487 ( .A1(n7968), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7970) );
  AND4_X2 U7488 ( .A1(n8680), .A2(n8639), .A3(n8640), .A4(n8641), .ZN(n8642)
         );
  NAND2_X1 U7489 ( .A1(n7793), .A2(n8111), .ZN(n8150) );
  AND3_X1 U7490 ( .A1(n9812), .A2(n9811), .A3(n9810), .ZN(n10364) );
  INV_X1 U7491 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8912) );
  INV_X1 U7492 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n14801) );
  INV_X4 U7493 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7494 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n9813) );
  NOR2_X2 U7495 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n8111) );
  NOR2_X1 U7496 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n9814) );
  NOR2_X1 U7497 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n7793) );
  NOR2_X1 U7498 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n7959) );
  NOR2_X1 U7499 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n7958) );
  NOR2_X1 U7500 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n8645) );
  INV_X1 U7501 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n15717) );
  INV_X1 U7502 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9152) );
  INV_X2 U7503 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7739) );
  INV_X1 U7504 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8644) );
  INV_X1 U7505 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n15715) );
  INV_X1 U7506 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8835) );
  INV_X1 U7507 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n14240) );
  OR2_X1 U7508 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), .ZN(
        n7900) );
  NOR2_X2 U7509 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8680) );
  XNOR2_X1 U7510 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8694) );
  NOR2_X1 U7511 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n7964) );
  INV_X1 U7512 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8791) );
  AND4_X1 U7513 ( .A1(n10364), .A2(n9836), .A3(n7736), .A4(n9815), .ZN(n7734)
         );
  NAND2_X1 U7514 ( .A1(n9837), .A2(n9836), .ZN(n9839) );
  NOR2_X1 U7515 ( .A1(n15736), .A2(n15735), .ZN(n15734) );
  NOR2_X2 U7516 ( .A1(n14992), .A2(n14943), .ZN(n7331) );
  AOI21_X2 U7517 ( .B1(n11100), .B2(n11099), .A(n11098), .ZN(n11097) );
  NOR2_X2 U7518 ( .A1(n13820), .A2(n13907), .ZN(n13803) );
  NAND2_X2 U7519 ( .A1(n8080), .A2(n8079), .ZN(n11758) );
  NAND2_X2 U7520 ( .A1(n6555), .A2(n8079), .ZN(n9664) );
  XNOR2_X2 U7521 ( .A(n7992), .B(n7991), .ZN(n8079) );
  NOR2_X2 U7522 ( .A1(n8150), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n8178) );
  NOR2_X2 U7523 ( .A1(n13870), .A2(n13710), .ZN(n13693) );
  OAI211_X1 U7524 ( .C1(n9610), .C2(n10487), .A(n7483), .B(n8113), .ZN(n12068)
         );
  INV_X1 U7525 ( .A(n8126), .ZN(n6554) );
  XNOR2_X1 U7526 ( .A(n8085), .B(n8084), .ZN(n8603) );
  INV_X1 U7527 ( .A(n8133), .ZN(n6556) );
  NAND2_X2 U7528 ( .A1(n7615), .A2(n6555), .ZN(n15256) );
  BUF_X4 U7529 ( .A(n8134), .Z(n6558) );
  INV_X1 U7530 ( .A(n8700), .ZN(n9113) );
  INV_X1 U7531 ( .A(n6547), .ZN(n9224) );
  OR2_X1 U7532 ( .A1(n8649), .A2(n8660), .ZN(n8650) );
  AND2_X1 U7533 ( .A1(n9149), .A2(n6932), .ZN(n8649) );
  NAND2_X1 U7534 ( .A1(n7571), .A2(n7570), .ZN(n7569) );
  OR2_X1 U7535 ( .A1(n13597), .A2(n13596), .ZN(n9605) );
  NAND2_X1 U7536 ( .A1(n6826), .A2(n6828), .ZN(n8063) );
  INV_X1 U7537 ( .A(n6829), .ZN(n6828) );
  NAND2_X1 U7538 ( .A1(n7766), .A2(n8428), .ZN(n7762) );
  AND2_X1 U7539 ( .A1(n8049), .A2(n7767), .ZN(n7766) );
  INV_X1 U7540 ( .A(n8445), .ZN(n7767) );
  AND2_X1 U7541 ( .A1(n10026), .A2(n9807), .ZN(n9808) );
  NAND2_X1 U7542 ( .A1(n10924), .A2(n10923), .ZN(n7244) );
  NAND2_X1 U7543 ( .A1(n6963), .A2(n6962), .ZN(n7482) );
  INV_X1 U7544 ( .A(n11560), .ZN(n6962) );
  OAI21_X1 U7545 ( .B1(n11213), .B2(n11217), .A(n11557), .ZN(n6963) );
  NAND2_X1 U7546 ( .A1(n7922), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7204) );
  NAND2_X1 U7547 ( .A1(n9787), .A2(n9696), .ZN(n9786) );
  NAND2_X1 U7548 ( .A1(n9787), .A2(n6897), .ZN(n6896) );
  INV_X1 U7549 ( .A(n9788), .ZN(n6897) );
  NAND2_X1 U7550 ( .A1(n7316), .A2(n6608), .ZN(n13751) );
  NAND2_X1 U7551 ( .A1(n6978), .A2(n6639), .ZN(n7316) );
  INV_X1 U7552 ( .A(n8702), .ZN(n9080) );
  CLKBUF_X1 U7553 ( .A(n8675), .Z(n10733) );
  INV_X1 U7554 ( .A(n9886), .ZN(n9863) );
  NAND2_X1 U7555 ( .A1(n10372), .A2(n10371), .ZN(n15052) );
  AOI21_X1 U7556 ( .B1(n13075), .B2(n9113), .A(n9112), .ZN(n12798) );
  NAND2_X1 U7557 ( .A1(n7142), .A2(n11440), .ZN(n9872) );
  NAND2_X1 U7558 ( .A1(n9974), .A2(n7577), .ZN(n7576) );
  INV_X1 U7559 ( .A(n9975), .ZN(n7577) );
  INV_X1 U7560 ( .A(n9495), .ZN(n7931) );
  NAND2_X1 U7561 ( .A1(n10033), .A2(n7570), .ZN(n7038) );
  AND2_X1 U7562 ( .A1(n10034), .A2(n7572), .ZN(n7571) );
  NAND2_X1 U7563 ( .A1(n7040), .A2(n7039), .ZN(n10033) );
  OAI21_X1 U7564 ( .B1(n10006), .B2(n7567), .A(n7219), .ZN(n7039) );
  NAND2_X1 U7565 ( .A1(n7041), .A2(n10017), .ZN(n7040) );
  AND2_X1 U7566 ( .A1(n7565), .A2(n7220), .ZN(n7219) );
  NAND2_X1 U7567 ( .A1(n7118), .A2(n10216), .ZN(n7117) );
  NAND2_X1 U7568 ( .A1(n12552), .A2(n12550), .ZN(n7118) );
  NAND2_X1 U7569 ( .A1(n7917), .A2(n7915), .ZN(n9549) );
  INV_X1 U7570 ( .A(n9569), .ZN(n7294) );
  NAND2_X1 U7571 ( .A1(n10204), .A2(n10207), .ZN(n7558) );
  AND2_X1 U7572 ( .A1(n7292), .A2(n9571), .ZN(n7290) );
  NAND2_X1 U7573 ( .A1(n7296), .A2(n7294), .ZN(n7292) );
  NAND2_X1 U7574 ( .A1(n6615), .A2(n7558), .ZN(n7557) );
  AOI21_X1 U7575 ( .B1(n7352), .B2(n7353), .A(n7760), .ZN(n7351) );
  NOR2_X1 U7576 ( .A1(n12617), .A2(n7097), .ZN(n7096) );
  INV_X1 U7577 ( .A(n12616), .ZN(n7097) );
  NOR2_X1 U7578 ( .A1(n10887), .A2(n7949), .ZN(n10889) );
  NOR2_X1 U7579 ( .A1(n6957), .A2(n11219), .ZN(n6956) );
  NOR2_X1 U7580 ( .A1(n7245), .A2(n11211), .ZN(n6957) );
  NAND2_X1 U7581 ( .A1(n7482), .A2(n7481), .ZN(n7207) );
  NAND2_X1 U7582 ( .A1(n11869), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7481) );
  NOR2_X1 U7583 ( .A1(n12910), .A2(n7484), .ZN(n12928) );
  NOR2_X1 U7584 ( .A1(n12396), .A2(n8840), .ZN(n7484) );
  NOR2_X1 U7585 ( .A1(n12990), .A2(n6763), .ZN(n12991) );
  NAND2_X1 U7586 ( .A1(n12646), .A2(n12798), .ZN(n9244) );
  NAND2_X1 U7587 ( .A1(n7390), .A2(n7388), .ZN(n9245) );
  NOR2_X1 U7588 ( .A1(n12798), .A2(n7389), .ZN(n7388) );
  INV_X1 U7589 ( .A(n9193), .ZN(n7389) );
  NAND2_X1 U7590 ( .A1(n7515), .A2(n7516), .ZN(n7510) );
  NAND2_X1 U7591 ( .A1(n7512), .A2(n7515), .ZN(n7509) );
  OAI21_X1 U7592 ( .B1(n7514), .B2(n7513), .A(n10377), .ZN(n7512) );
  NOR2_X1 U7593 ( .A1(n9133), .A2(n7536), .ZN(n7535) );
  INV_X1 U7594 ( .A(n9130), .ZN(n7536) );
  OR2_X1 U7595 ( .A1(n15331), .A2(n12144), .ZN(n9286) );
  AND2_X1 U7596 ( .A1(n6584), .A2(n7885), .ZN(n7884) );
  NOR2_X1 U7597 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n7885) );
  INV_X1 U7598 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8638) );
  OAI21_X1 U7599 ( .B1(n8850), .B2(n8849), .A(n8851), .ZN(n8852) );
  INV_X1 U7600 ( .A(n8848), .ZN(n8849) );
  INV_X1 U7601 ( .A(n8812), .ZN(n7387) );
  NOR2_X1 U7602 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n8639) );
  NOR2_X1 U7603 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n8640) );
  NOR2_X1 U7604 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_5__SCAN_IN), .ZN(
        n8641) );
  NAND2_X1 U7605 ( .A1(n13414), .A2(n7139), .ZN(n8480) );
  NAND2_X1 U7606 ( .A1(n8466), .A2(n7140), .ZN(n7139) );
  INV_X1 U7607 ( .A(n8467), .ZN(n7140) );
  OR2_X1 U7608 ( .A1(n9695), .A2(n9630), .ZN(n9649) );
  INV_X1 U7609 ( .A(n13949), .ZN(n7976) );
  NOR2_X1 U7610 ( .A1(n13732), .A2(n13879), .ZN(n7498) );
  OR2_X1 U7611 ( .A1(n9767), .A2(n7605), .ZN(n7604) );
  INV_X1 U7612 ( .A(n9766), .ZN(n7605) );
  AND2_X1 U7613 ( .A1(n12043), .A2(n8153), .ZN(n6887) );
  NAND2_X1 U7614 ( .A1(n6553), .A2(n7272), .ZN(n9706) );
  NAND2_X1 U7615 ( .A1(n9708), .A2(n9676), .ZN(n9739) );
  NAND2_X1 U7616 ( .A1(n11781), .A2(n13525), .ZN(n9676) );
  NOR2_X1 U7617 ( .A1(n6896), .A2(n6892), .ZN(n6891) );
  INV_X1 U7618 ( .A(n6899), .ZN(n6892) );
  NAND2_X1 U7619 ( .A1(n7498), .A2(n7497), .ZN(n13710) );
  NAND2_X1 U7620 ( .A1(n12291), .A2(n6736), .ZN(n7852) );
  NAND2_X1 U7621 ( .A1(n12713), .A2(n12714), .ZN(n7822) );
  AOI21_X1 U7622 ( .B1(n7833), .B2(n7836), .A(n12761), .ZN(n6951) );
  INV_X1 U7623 ( .A(n11132), .ZN(n9903) );
  NOR2_X1 U7624 ( .A1(n14277), .A2(n7367), .ZN(n7366) );
  NOR2_X1 U7625 ( .A1(n14300), .A2(n7368), .ZN(n7367) );
  NOR2_X1 U7626 ( .A1(n14362), .A2(n7475), .ZN(n7474) );
  INV_X1 U7627 ( .A(n7476), .ZN(n7475) );
  NAND2_X1 U7628 ( .A1(n10700), .A2(n11897), .ZN(n11132) );
  NAND2_X1 U7629 ( .A1(n11727), .A2(n11722), .ZN(n11886) );
  NAND2_X1 U7630 ( .A1(n11082), .A2(n11897), .ZN(n10705) );
  NAND2_X1 U7631 ( .A1(n6818), .A2(n9587), .ZN(n9623) );
  NAND2_X1 U7632 ( .A1(n8062), .A2(n12207), .ZN(n8064) );
  NAND2_X1 U7633 ( .A1(n8063), .A2(SI_24_), .ZN(n8065) );
  NAND3_X1 U7634 ( .A1(n8064), .A2(n7770), .A3(n8065), .ZN(n8503) );
  INV_X1 U7635 ( .A(n8500), .ZN(n7770) );
  OAI21_X1 U7636 ( .B1(n8087), .B2(n7749), .A(n7747), .ZN(n8058) );
  INV_X1 U7637 ( .A(n7748), .ZN(n7747) );
  OAI21_X1 U7638 ( .B1(n8086), .B2(n7749), .A(SI_22_), .ZN(n7748) );
  INV_X1 U7639 ( .A(n8054), .ZN(n7749) );
  XNOR2_X1 U7640 ( .A(n8050), .B(SI_19_), .ZN(n8445) );
  NAND2_X1 U7641 ( .A1(n8049), .A2(n8047), .ZN(n8428) );
  XNOR2_X1 U7642 ( .A(n8045), .B(SI_17_), .ZN(n8405) );
  OAI21_X1 U7643 ( .B1(n8306), .B2(n7353), .A(n7352), .ZN(n8387) );
  INV_X1 U7644 ( .A(SI_11_), .ZN(n8029) );
  NAND2_X1 U7645 ( .A1(n7065), .A2(n7064), .ZN(n8196) );
  AOI21_X1 U7646 ( .B1(n8011), .B2(n7066), .A(n6654), .ZN(n7065) );
  NAND2_X1 U7647 ( .A1(n7300), .A2(n8003), .ZN(n7037) );
  XNOR2_X1 U7648 ( .A(n14647), .B(n7174), .ZN(n14682) );
  XNOR2_X1 U7649 ( .A(n7027), .B(P3_ADDR_REG_5__SCAN_IN), .ZN(n14696) );
  AOI21_X1 U7650 ( .B1(n14705), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n14653), .ZN(
        n14709) );
  AOI21_X1 U7651 ( .B1(n12869), .B2(n13157), .A(n12627), .ZN(n12630) );
  XNOR2_X1 U7652 ( .A(n7244), .B(n10925), .ZN(n10926) );
  OR2_X1 U7653 ( .A1(n10926), .A2(n10910), .ZN(n7166) );
  XNOR2_X1 U7654 ( .A(n7207), .B(n11873), .ZN(n11870) );
  INV_X1 U7655 ( .A(n11902), .ZN(n7685) );
  OR2_X1 U7656 ( .A1(n12354), .A2(n8816), .ZN(n7241) );
  NAND2_X1 U7657 ( .A1(n7196), .A2(n6636), .ZN(n7681) );
  INV_X1 U7658 ( .A(n7185), .ZN(n12394) );
  NAND2_X1 U7659 ( .A1(n7681), .A2(n7680), .ZN(n6751) );
  INV_X1 U7660 ( .A(n12397), .ZN(n7680) );
  XNOR2_X1 U7661 ( .A(n12928), .B(n12929), .ZN(n12911) );
  OR2_X1 U7662 ( .A1(n12987), .A2(n12986), .ZN(n6967) );
  NAND3_X1 U7663 ( .A1(n6966), .A2(P3_REG1_REG_17__SCAN_IN), .A3(n13023), .ZN(
        n13024) );
  NOR2_X1 U7664 ( .A1(n13013), .A2(n12992), .ZN(n12993) );
  AND2_X1 U7665 ( .A1(n13003), .A2(n12991), .ZN(n12992) );
  NOR2_X1 U7666 ( .A1(n13006), .A2(n6735), .ZN(n13031) );
  NAND2_X1 U7667 ( .A1(n9244), .A2(n9245), .ZN(n13070) );
  OR2_X1 U7668 ( .A1(n13355), .A2(n13172), .ZN(n9347) );
  OR2_X1 U7669 ( .A1(n15281), .A2(n15283), .ZN(n8815) );
  NOR2_X1 U7670 ( .A1(n6589), .A2(n7229), .ZN(n11699) );
  NAND3_X1 U7671 ( .A1(n10733), .A2(n10736), .A3(n10731), .ZN(n15298) );
  OR2_X1 U7672 ( .A1(n15421), .A2(n12137), .ZN(n11691) );
  INV_X1 U7673 ( .A(n13107), .ZN(n15363) );
  INV_X1 U7674 ( .A(n8994), .ZN(n9234) );
  INV_X1 U7675 ( .A(n8722), .ZN(n9216) );
  NAND2_X1 U7676 ( .A1(n8675), .A2(n8013), .ZN(n8994) );
  NAND2_X1 U7677 ( .A1(n9114), .A2(n10731), .ZN(n15300) );
  OAI22_X1 U7678 ( .A1(n9191), .A2(n9190), .B1(P2_DATAO_REG_27__SCAN_IN), .B2(
        n13956), .ZN(n9198) );
  NAND2_X1 U7679 ( .A1(n8989), .A2(n7017), .ZN(n9006) );
  INV_X1 U7680 ( .A(n8907), .ZN(n7379) );
  AND2_X1 U7681 ( .A1(n8708), .A2(n15706), .ZN(n8729) );
  XNOR2_X1 U7682 ( .A(n8499), .B(n8488), .ZN(n13397) );
  AND2_X1 U7683 ( .A1(n7647), .A2(n7646), .ZN(n7645) );
  INV_X1 U7684 ( .A(n13439), .ZN(n7646) );
  NAND2_X1 U7685 ( .A1(n14843), .A2(n8365), .ZN(n8384) );
  NAND2_X1 U7686 ( .A1(n9600), .A2(n9599), .ZN(n13597) );
  OAI21_X1 U7687 ( .B1(n6592), .B2(n7594), .A(n13611), .ZN(n7593) );
  XNOR2_X1 U7688 ( .A(n13849), .B(n13637), .ZN(n13628) );
  NAND2_X1 U7689 ( .A1(n13855), .A2(n13424), .ZN(n7298) );
  NAND2_X1 U7690 ( .A1(n6982), .A2(n7781), .ZN(n6980) );
  NAND2_X1 U7691 ( .A1(n13654), .A2(n6982), .ZN(n6981) );
  NAND2_X1 U7692 ( .A1(n7312), .A2(n7311), .ZN(n13702) );
  AND2_X1 U7693 ( .A1(n6565), .A2(n13700), .ZN(n7311) );
  AND2_X1 U7694 ( .A1(n7307), .A2(n7310), .ZN(n7130) );
  AOI21_X1 U7695 ( .B1(n13616), .B2(n12603), .A(n8285), .ZN(n7753) );
  XNOR2_X1 U7696 ( .A(n12603), .B(n9671), .ZN(n9788) );
  NAND2_X1 U7697 ( .A1(n11471), .A2(n11470), .ZN(n11476) );
  AND2_X1 U7698 ( .A1(n13972), .A2(n7811), .ZN(n7810) );
  OR2_X1 U7699 ( .A1(n14073), .A2(n12767), .ZN(n7811) );
  NAND2_X1 U7700 ( .A1(n7822), .A2(n7823), .ZN(n7818) );
  OR2_X1 U7701 ( .A1(n7819), .A2(n7817), .ZN(n7816) );
  INV_X1 U7702 ( .A(n7822), .ZN(n7817) );
  AND2_X1 U7703 ( .A1(n14041), .A2(n7820), .ZN(n7819) );
  OR2_X1 U7704 ( .A1(n7821), .A2(n12708), .ZN(n7820) );
  NAND2_X1 U7705 ( .A1(n6946), .A2(n6951), .ZN(n14072) );
  NAND2_X1 U7706 ( .A1(n13981), .A2(n7833), .ZN(n6946) );
  NAND2_X1 U7707 ( .A1(n7159), .A2(n7158), .ZN(n14260) );
  NOR2_X1 U7708 ( .A1(n14332), .A2(n7332), .ZN(n14281) );
  NOR2_X1 U7709 ( .A1(n12564), .A2(n7701), .ZN(n7700) );
  INV_X1 U7710 ( .A(n12562), .ZN(n7701) );
  AOI21_X1 U7711 ( .B1(n6853), .B2(n6855), .A(n6850), .ZN(n12585) );
  NAND2_X1 U7712 ( .A1(n6671), .A2(n6851), .ZN(n6850) );
  NOR2_X1 U7713 ( .A1(n14445), .A2(n7695), .ZN(n7694) );
  INV_X1 U7714 ( .A(n12556), .ZN(n7695) );
  NAND2_X1 U7715 ( .A1(n7724), .A2(n7720), .ZN(n12029) );
  NOR2_X1 U7716 ( .A1(n12023), .A2(n7937), .ZN(n7720) );
  NAND2_X1 U7717 ( .A1(n11308), .A2(n9911), .ZN(n7690) );
  OAI21_X1 U7718 ( .B1(n14629), .B2(n8013), .A(n6865), .ZN(n9886) );
  NAND2_X1 U7719 ( .A1(n6869), .A2(n6866), .ZN(n6865) );
  NAND2_X1 U7720 ( .A1(n10486), .A2(n6870), .ZN(n6867) );
  INV_X1 U7721 ( .A(n14951), .ZN(n14902) );
  AND2_X1 U7722 ( .A1(n11133), .A2(n12791), .ZN(n11305) );
  OR2_X1 U7723 ( .A1(n10084), .A2(n7738), .ZN(n9816) );
  INV_X1 U7724 ( .A(n7045), .ZN(n7044) );
  OAI21_X1 U7725 ( .B1(n8021), .B2(n7046), .A(n8250), .ZN(n7045) );
  INV_X1 U7726 ( .A(n8023), .ZN(n7046) );
  NAND2_X1 U7727 ( .A1(n14916), .A2(n7653), .ZN(n7032) );
  OR2_X1 U7728 ( .A1(n14916), .A2(n7653), .ZN(n7031) );
  XNOR2_X1 U7729 ( .A(n12630), .B(n12628), .ZN(n12804) );
  NAND2_X1 U7730 ( .A1(n12813), .A2(n12619), .ZN(n12864) );
  AND2_X1 U7731 ( .A1(n9086), .A2(n9085), .ZN(n13090) );
  AND2_X1 U7732 ( .A1(n9229), .A2(n9207), .ZN(n13074) );
  AOI21_X1 U7733 ( .B1(n11226), .B2(n11225), .A(n11224), .ZN(n11547) );
  OR2_X1 U7734 ( .A1(n11549), .A2(n11548), .ZN(n6835) );
  NOR2_X1 U7735 ( .A1(n13009), .A2(n13010), .ZN(n13029) );
  NAND2_X1 U7736 ( .A1(n10386), .A2(n10385), .ZN(n13059) );
  NAND2_X1 U7737 ( .A1(n7791), .A2(n13819), .ZN(n7788) );
  AND2_X1 U7738 ( .A1(n7729), .A2(n7147), .ZN(n14524) );
  AOI21_X1 U7739 ( .B1(n14287), .B2(n15059), .A(n14280), .ZN(n7729) );
  NAND2_X1 U7740 ( .A1(n7143), .A2(n11479), .ZN(n7142) );
  NOR2_X1 U7741 ( .A1(n14109), .A2(n10283), .ZN(n7143) );
  NAND2_X1 U7742 ( .A1(n7107), .A2(n7556), .ZN(n7554) );
  NAND2_X1 U7743 ( .A1(n9925), .A2(n9926), .ZN(n7556) );
  NAND2_X1 U7744 ( .A1(n7555), .A2(n9924), .ZN(n7553) );
  INV_X1 U7745 ( .A(n9926), .ZN(n7555) );
  NAND2_X1 U7746 ( .A1(n6605), .A2(n7576), .ZN(n7575) );
  AND2_X1 U7747 ( .A1(n7576), .A2(n7218), .ZN(n7217) );
  INV_X1 U7748 ( .A(n9988), .ZN(n7218) );
  NAND2_X1 U7749 ( .A1(n7042), .A2(n6631), .ZN(n7041) );
  NAND2_X1 U7750 ( .A1(n10006), .A2(n7565), .ZN(n7042) );
  NAND2_X1 U7751 ( .A1(n7567), .A2(n7565), .ZN(n7564) );
  INV_X1 U7752 ( .A(n9490), .ZN(n7279) );
  NAND2_X1 U7753 ( .A1(n7902), .A2(n7901), .ZN(n9491) );
  NAND2_X1 U7754 ( .A1(n6645), .A2(n7903), .ZN(n7901) );
  NAND2_X1 U7755 ( .A1(n7253), .A2(n7251), .ZN(n7902) );
  NOR2_X1 U7756 ( .A1(n6600), .A2(n7252), .ZN(n7251) );
  NAND2_X1 U7757 ( .A1(n9490), .A2(n7277), .ZN(n7276) );
  NAND2_X1 U7758 ( .A1(n10032), .A2(n10035), .ZN(n7570) );
  AND2_X1 U7759 ( .A1(n10057), .A2(n10056), .ZN(n7061) );
  NOR2_X1 U7760 ( .A1(n7581), .A2(n7062), .ZN(n7580) );
  AND3_X1 U7761 ( .A1(n7117), .A2(n7119), .A3(n12259), .ZN(n7062) );
  NOR2_X1 U7762 ( .A1(n6590), .A2(n7265), .ZN(n7264) );
  NOR2_X1 U7763 ( .A1(n7267), .A2(n9509), .ZN(n7265) );
  INV_X1 U7764 ( .A(n9513), .ZN(n7925) );
  INV_X1 U7765 ( .A(n9529), .ZN(n7909) );
  NAND2_X1 U7766 ( .A1(n10175), .A2(n7070), .ZN(n7069) );
  INV_X1 U7767 ( .A(n10174), .ZN(n7070) );
  NOR2_X1 U7768 ( .A1(n6598), .A2(n7920), .ZN(n7919) );
  OAI21_X1 U7769 ( .B1(n9543), .B2(n7919), .A(n7281), .ZN(n9551) );
  NOR2_X1 U7770 ( .A1(n9546), .A2(n7282), .ZN(n7281) );
  INV_X1 U7771 ( .A(n7918), .ZN(n7282) );
  NOR2_X1 U7772 ( .A1(n7296), .A2(n7294), .ZN(n7293) );
  NAND2_X1 U7773 ( .A1(n7290), .A2(n7293), .ZN(n7289) );
  NAND2_X1 U7774 ( .A1(n6599), .A2(n7935), .ZN(n7933) );
  NAND2_X1 U7775 ( .A1(n7286), .A2(n7285), .ZN(n7284) );
  NAND2_X1 U7776 ( .A1(n7295), .A2(n7292), .ZN(n7285) );
  INV_X1 U7777 ( .A(n7290), .ZN(n7286) );
  NAND2_X1 U7778 ( .A1(n7557), .A2(n10218), .ZN(n7051) );
  INV_X1 U7779 ( .A(n10232), .ZN(n7563) );
  INV_X1 U7780 ( .A(n8068), .ZN(n6825) );
  INV_X1 U7781 ( .A(SI_17_), .ZN(n8044) );
  INV_X1 U7782 ( .A(n8043), .ZN(n7761) );
  INV_X1 U7783 ( .A(n15436), .ZN(n7413) );
  NAND2_X1 U7784 ( .A1(n7021), .A2(n7020), .ZN(n7024) );
  OR2_X1 U7785 ( .A1(n6673), .A2(n7025), .ZN(n7020) );
  INV_X1 U7786 ( .A(n9246), .ZN(n7025) );
  NAND2_X1 U7787 ( .A1(n13330), .A2(n13090), .ZN(n7515) );
  INV_X1 U7788 ( .A(n9144), .ZN(n7547) );
  OR2_X1 U7789 ( .A1(n12409), .A2(n14809), .ZN(n9313) );
  OR2_X1 U7790 ( .A1(n13898), .A2(n9720), .ZN(n7805) );
  INV_X1 U7791 ( .A(n12025), .ZN(n6862) );
  AOI21_X1 U7792 ( .B1(n7773), .B2(n7771), .A(n6659), .ZN(n7352) );
  INV_X1 U7793 ( .A(n7771), .ZN(n7353) );
  INV_X1 U7794 ( .A(n8026), .ZN(n7345) );
  NOR2_X1 U7795 ( .A1(n7348), .A2(n8027), .ZN(n7347) );
  OAI21_X1 U7796 ( .B1(n10486), .B2(P2_DATAO_REG_11__SCAN_IN), .A(n7171), .ZN(
        n8030) );
  NAND2_X1 U7797 ( .A1(n10486), .A2(n10571), .ZN(n7171) );
  AND2_X1 U7798 ( .A1(n7743), .A2(n7742), .ZN(n8002) );
  OAI21_X1 U7799 ( .B1(n14690), .B2(n14689), .A(n6601), .ZN(n7029) );
  INV_X1 U7800 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15566) );
  NAND2_X1 U7801 ( .A1(n15354), .A2(n15344), .ZN(n9266) );
  NAND2_X1 U7802 ( .A1(n7424), .A2(n7425), .ZN(n7423) );
  INV_X1 U7803 ( .A(n12329), .ZN(n7424) );
  NAND3_X1 U7804 ( .A1(n7208), .A2(n12010), .A3(n6623), .ZN(n7104) );
  OR2_X1 U7805 ( .A1(n13070), .A2(n10377), .ZN(n9247) );
  AND2_X1 U7806 ( .A1(n9400), .A2(n13092), .ZN(n7395) );
  NOR2_X1 U7807 ( .A1(n10894), .A2(n7194), .ZN(n10895) );
  AND2_X1 U7808 ( .A1(n6548), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7194) );
  INV_X1 U7809 ( .A(n7207), .ZN(n11912) );
  INV_X1 U7810 ( .A(n7675), .ZN(n6761) );
  AND2_X1 U7811 ( .A1(n7674), .A2(n6580), .ZN(n6764) );
  NOR2_X1 U7812 ( .A1(n12947), .A2(n6838), .ZN(n12968) );
  AND2_X1 U7813 ( .A1(n12954), .A2(n12948), .ZN(n6838) );
  OR2_X1 U7814 ( .A1(n10393), .A2(n13074), .ZN(n9374) );
  NOR2_X1 U7815 ( .A1(n13092), .A2(n7518), .ZN(n7514) );
  OR2_X1 U7816 ( .A1(n13093), .A2(n12830), .ZN(n9243) );
  NAND2_X1 U7817 ( .A1(n9048), .A2(n9047), .ZN(n9064) );
  OR2_X1 U7818 ( .A1(n12832), .A2(n13089), .ZN(n9368) );
  AND2_X1 U7819 ( .A1(n6611), .A2(n7546), .ZN(n7540) );
  AND2_X1 U7820 ( .A1(n7542), .A2(n7544), .ZN(n7541) );
  AOI21_X1 U7821 ( .B1(n6928), .B2(n6588), .A(n7545), .ZN(n7544) );
  NOR2_X1 U7822 ( .A1(n13345), .A2(n12872), .ZN(n7545) );
  OR2_X1 U7823 ( .A1(n13280), .A2(n13157), .ZN(n9357) );
  INV_X1 U7824 ( .A(n9350), .ZN(n7893) );
  NAND2_X1 U7825 ( .A1(n14817), .A2(n6915), .ZN(n6914) );
  NOR2_X1 U7826 ( .A1(n6918), .A2(n6916), .ZN(n6915) );
  INV_X1 U7827 ( .A(n9300), .ZN(n6916) );
  AOI21_X1 U7828 ( .B1(n7878), .B2(n7879), .A(n7877), .ZN(n7876) );
  INV_X1 U7829 ( .A(n7882), .ZN(n7878) );
  INV_X1 U7830 ( .A(n13246), .ZN(n7877) );
  NAND2_X1 U7831 ( .A1(n9314), .A2(n9312), .ZN(n7881) );
  INV_X1 U7832 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n12385) );
  NOR2_X1 U7833 ( .A1(n11992), .A2(n7505), .ZN(n7504) );
  INV_X1 U7834 ( .A(n9118), .ZN(n7505) );
  OR2_X1 U7835 ( .A1(n15343), .A2(n11999), .ZN(n9264) );
  AND2_X1 U7836 ( .A1(n8646), .A2(n9152), .ZN(n7429) );
  INV_X1 U7837 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8646) );
  NAND2_X1 U7838 ( .A1(n8978), .A2(n8977), .ZN(n8987) );
  AND2_X1 U7839 ( .A1(n8637), .A2(n8636), .ZN(n6802) );
  NOR2_X1 U7840 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n8636) );
  AND2_X1 U7841 ( .A1(n8835), .A2(n8877), .ZN(n6803) );
  INV_X1 U7842 ( .A(n7631), .ZN(n7629) );
  NAND2_X1 U7843 ( .A1(n7928), .A2(n7927), .ZN(n9581) );
  NAND2_X1 U7844 ( .A1(n9575), .A2(n7930), .ZN(n7927) );
  OR2_X1 U7845 ( .A1(n9573), .A2(n7929), .ZN(n7928) );
  NOR2_X1 U7846 ( .A1(n9575), .A2(n7930), .ZN(n7929) );
  NOR2_X1 U7847 ( .A1(n7594), .A2(n6900), .ZN(n6899) );
  INV_X1 U7848 ( .A(n9782), .ZN(n6900) );
  INV_X1 U7849 ( .A(n7599), .ZN(n7598) );
  AND2_X1 U7850 ( .A1(n9764), .A2(n7607), .ZN(n7606) );
  INV_X1 U7851 ( .A(n13795), .ZN(n7607) );
  NAND2_X1 U7852 ( .A1(n13831), .A2(n13830), .ZN(n9765) );
  AND2_X1 U7853 ( .A1(n6560), .A2(n12123), .ZN(n7796) );
  NOR2_X1 U7854 ( .A1(n12245), .A2(n7799), .ZN(n7797) );
  AND2_X1 U7855 ( .A1(n9755), .A2(n6904), .ZN(n6903) );
  OR2_X1 U7856 ( .A1(n12073), .A2(n6905), .ZN(n6904) );
  INV_X1 U7857 ( .A(n9754), .ZN(n6905) );
  NAND2_X1 U7858 ( .A1(n13922), .A2(n6984), .ZN(n9708) );
  NOR2_X1 U7859 ( .A1(n8610), .A2(n9789), .ZN(n8097) );
  OR2_X1 U7860 ( .A1(n9667), .A2(n8080), .ZN(n8610) );
  INV_X1 U7861 ( .A(n9783), .ZN(n7170) );
  NOR2_X1 U7862 ( .A1(n8571), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n8585) );
  INV_X1 U7863 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8587) );
  NOR2_X1 U7864 ( .A1(n7829), .A2(n14016), .ZN(n7825) );
  NAND2_X1 U7865 ( .A1(n14944), .A2(n12301), .ZN(n12308) );
  INV_X1 U7866 ( .A(n7833), .ZN(n6949) );
  NAND2_X1 U7867 ( .A1(n14286), .A2(n7333), .ZN(n7332) );
  INV_X1 U7868 ( .A(n7334), .ZN(n7333) );
  OR2_X1 U7869 ( .A1(n14299), .A2(n7368), .ZN(n7365) );
  INV_X1 U7870 ( .A(n7445), .ZN(n7442) );
  NAND2_X1 U7871 ( .A1(n14372), .A2(n14371), .ZN(n12563) );
  AND2_X1 U7872 ( .A1(n14374), .A2(n12587), .ZN(n7476) );
  AND2_X1 U7873 ( .A1(n6854), .A2(n7456), .ZN(n6853) );
  AOI21_X1 U7874 ( .B1(n7718), .B2(n7716), .A(n7715), .ZN(n7714) );
  INV_X1 U7875 ( .A(n12031), .ZN(n7716) );
  INV_X1 U7876 ( .A(n12165), .ZN(n7715) );
  INV_X1 U7877 ( .A(n6586), .ZN(n7467) );
  NOR2_X1 U7878 ( .A1(n6861), .A2(n6860), .ZN(n6859) );
  NOR2_X1 U7879 ( .A1(n12023), .A2(n6862), .ZN(n6860) );
  INV_X1 U7880 ( .A(n7468), .ZN(n6861) );
  NAND2_X1 U7881 ( .A1(n6859), .A2(n6862), .ZN(n6857) );
  NAND2_X1 U7882 ( .A1(n11585), .A2(n11589), .ZN(n7706) );
  AOI21_X1 U7883 ( .B1(n7436), .B2(n7435), .A(n7431), .ZN(n7430) );
  NAND2_X1 U7884 ( .A1(n14299), .A2(n14300), .ZN(n14298) );
  NAND2_X1 U7885 ( .A1(n7329), .A2(n7328), .ZN(n14893) );
  INV_X1 U7886 ( .A(n14870), .ZN(n7328) );
  NOR2_X1 U7887 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n9810) );
  NOR2_X1 U7888 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n9811) );
  AND2_X1 U7889 ( .A1(n8065), .A2(n7769), .ZN(n7768) );
  INV_X1 U7890 ( .A(n8515), .ZN(n7769) );
  NOR2_X1 U7891 ( .A1(n7859), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n7858) );
  INV_X1 U7892 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n10354) );
  NAND2_X1 U7893 ( .A1(n8051), .A2(n11543), .ZN(n6807) );
  NAND2_X1 U7894 ( .A1(n7762), .A2(n7763), .ZN(n8051) );
  NAND2_X1 U7895 ( .A1(n7354), .A2(n7762), .ZN(n6808) );
  AND2_X1 U7896 ( .A1(n7763), .A2(SI_20_), .ZN(n7354) );
  NAND2_X1 U7897 ( .A1(n7149), .A2(SI_18_), .ZN(n8049) );
  OAI21_X1 U7898 ( .B1(n8306), .B2(n6568), .A(n7774), .ZN(n8346) );
  AND2_X1 U7899 ( .A1(n6815), .A2(n6814), .ZN(n7774) );
  INV_X1 U7900 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n15595) );
  NAND2_X1 U7901 ( .A1(n8196), .A2(n8014), .ZN(n8214) );
  NAND2_X1 U7902 ( .A1(n7037), .A2(n8146), .ZN(n7740) );
  XNOR2_X1 U7903 ( .A(n7029), .B(P3_ADDR_REG_3__SCAN_IN), .ZN(n14691) );
  OAI21_X1 U7904 ( .B1(n14682), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6607), .ZN(
        n7027) );
  OAI22_X1 U7905 ( .A1(n14701), .A2(n14651), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n11071), .ZN(n14652) );
  AND2_X1 U7906 ( .A1(n11071), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n14651) );
  OAI21_X1 U7907 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n14656), .A(n14655), .ZN(
        n14657) );
  NAND2_X1 U7908 ( .A1(n14681), .A2(n14680), .ZN(n14655) );
  OAI21_X1 U7909 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n15455), .A(n14663), .ZN(
        n14721) );
  NAND2_X1 U7910 ( .A1(n9288), .A2(n9287), .ZN(n15328) );
  INV_X1 U7911 ( .A(n7090), .ZN(n7088) );
  NOR2_X1 U7912 ( .A1(n12506), .A2(n12425), .ZN(n7090) );
  OR2_X1 U7913 ( .A1(n12183), .A2(n12180), .ZN(n7425) );
  AOI21_X1 U7914 ( .B1(n7426), .B2(n7096), .A(n6579), .ZN(n7094) );
  INV_X1 U7915 ( .A(n7096), .ZN(n7095) );
  NAND2_X1 U7916 ( .A1(n7410), .A2(n7409), .ZN(n7403) );
  AND2_X1 U7917 ( .A1(n7409), .A2(n7405), .ZN(n7404) );
  INV_X1 U7918 ( .A(n7408), .ZN(n7405) );
  INV_X1 U7919 ( .A(n10467), .ZN(n7520) );
  NAND2_X1 U7920 ( .A1(n8675), .A2(n7524), .ZN(n7523) );
  NAND2_X1 U7921 ( .A1(n10485), .A2(SI_1_), .ZN(n7524) );
  NAND2_X1 U7922 ( .A1(n7176), .A2(n7230), .ZN(n7411) );
  NOR2_X1 U7923 ( .A1(n11573), .A2(n11574), .ZN(n7230) );
  AOI21_X1 U7924 ( .B1(n7420), .B2(n7078), .A(n6625), .ZN(n7077) );
  INV_X1 U7925 ( .A(n12863), .ZN(n7078) );
  XNOR2_X1 U7926 ( .A(n13147), .B(n12640), .ZN(n12625) );
  OR2_X1 U7927 ( .A1(n8951), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8972) );
  NOR2_X1 U7928 ( .A1(n13257), .A2(n12895), .ZN(n9402) );
  OR2_X1 U7929 ( .A1(n8700), .A2(n11396), .ZN(n8654) );
  NAND2_X1 U7930 ( .A1(n9162), .A2(n9161), .ZN(n10934) );
  AND2_X1 U7931 ( .A1(n9160), .A2(n9159), .ZN(n9161) );
  OAI21_X1 U7932 ( .B1(n10758), .B2(n10744), .A(n10745), .ZN(n10961) );
  NAND2_X1 U7933 ( .A1(n7186), .A2(n11099), .ZN(n10772) );
  NAND2_X1 U7934 ( .A1(n6772), .A2(n6771), .ZN(n10908) );
  INV_X1 U7935 ( .A(n6770), .ZN(n6772) );
  OAI21_X1 U7936 ( .B1(n10890), .B2(P3_REG2_REG_3__SCAN_IN), .A(n6773), .ZN(
        n6770) );
  NAND2_X1 U7937 ( .A1(n7166), .A2(n6559), .ZN(n7246) );
  OAI21_X1 U7938 ( .B1(n11212), .B2(n11221), .A(n11557), .ZN(n11213) );
  OAI211_X1 U7939 ( .C1(n7166), .C2(n11073), .A(n7479), .B(n6604), .ZN(n11212)
         );
  NAND2_X1 U7940 ( .A1(n6964), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7242) );
  INV_X1 U7941 ( .A(n11213), .ZN(n6964) );
  OAI21_X1 U7942 ( .B1(n7197), .B2(n11554), .A(n6779), .ZN(n7237) );
  INV_X1 U7943 ( .A(n6780), .ZN(n6779) );
  OAI21_X1 U7944 ( .B1(n11550), .B2(n11554), .A(n7683), .ZN(n6780) );
  NAND2_X1 U7945 ( .A1(n11869), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7683) );
  NAND2_X1 U7946 ( .A1(n6958), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7243) );
  INV_X1 U7947 ( .A(n11870), .ZN(n6958) );
  AND2_X1 U7948 ( .A1(n6833), .A2(n6832), .ZN(n12389) );
  NAND2_X1 U7949 ( .A1(n12350), .A2(n12351), .ZN(n6832) );
  NAND2_X1 U7950 ( .A1(n6754), .A2(n6753), .ZN(n7185) );
  AOI21_X1 U7951 ( .B1(n11901), .B2(n7685), .A(n6698), .ZN(n6753) );
  NAND2_X1 U7952 ( .A1(n7241), .A2(n6637), .ZN(n7486) );
  INV_X1 U7953 ( .A(n7206), .ZN(n12381) );
  AOI21_X1 U7954 ( .B1(n12905), .B2(n14765), .A(n12904), .ZN(n12907) );
  NAND2_X1 U7955 ( .A1(n12907), .A2(n12906), .ZN(n12923) );
  AND2_X1 U7956 ( .A1(n6751), .A2(n6731), .ZN(n12919) );
  NAND2_X1 U7957 ( .A1(n6777), .A2(n6776), .ZN(n7232) );
  INV_X1 U7958 ( .A(n12922), .ZN(n6776) );
  INV_X1 U7959 ( .A(n12921), .ZN(n6777) );
  OAI22_X1 U7960 ( .A1(n12911), .A2(n6968), .B1(n6563), .B2(n12931), .ZN(
        n12941) );
  NAND2_X1 U7961 ( .A1(n7478), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n6968) );
  NOR2_X1 U7962 ( .A1(n12926), .A2(n12927), .ZN(n12947) );
  NAND2_X1 U7963 ( .A1(n12953), .A2(n12971), .ZN(n7674) );
  NOR2_X1 U7964 ( .A1(n12950), .A2(n12949), .ZN(n12969) );
  OR2_X1 U7965 ( .A1(n9020), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9035) );
  NAND2_X1 U7966 ( .A1(n13155), .A2(n13150), .ZN(n13140) );
  INV_X1 U7967 ( .A(n13181), .ZN(n7897) );
  INV_X1 U7968 ( .A(n9347), .ZN(n7895) );
  NAND2_X1 U7969 ( .A1(n13198), .A2(n9338), .ZN(n13181) );
  NOR2_X1 U7970 ( .A1(n13202), .A2(n7549), .ZN(n7548) );
  INV_X1 U7971 ( .A(n9139), .ZN(n7549) );
  NAND2_X1 U7972 ( .A1(n13219), .A2(n6930), .ZN(n13198) );
  AND2_X1 U7973 ( .A1(n13202), .A2(n9334), .ZN(n6930) );
  NAND2_X1 U7974 ( .A1(n9138), .A2(n9137), .ZN(n13216) );
  NAND2_X1 U7975 ( .A1(n13221), .A2(n13220), .ZN(n13219) );
  INV_X1 U7976 ( .A(n12897), .ZN(n13232) );
  OAI21_X1 U7977 ( .B1(n9131), .B2(n7533), .A(n7530), .ZN(n13242) );
  AOI21_X1 U7978 ( .B1(n7532), .B2(n7531), .A(n6710), .ZN(n7530) );
  INV_X1 U7979 ( .A(n7535), .ZN(n7531) );
  NOR2_X1 U7980 ( .A1(n12527), .A2(n7883), .ZN(n7882) );
  AND2_X1 U7981 ( .A1(n9324), .A2(n9329), .ZN(n13246) );
  NAND2_X1 U7982 ( .A1(n8865), .A2(n8864), .ZN(n8881) );
  INV_X1 U7983 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8864) );
  INV_X1 U7984 ( .A(n8866), .ZN(n8865) );
  INV_X1 U7985 ( .A(n6917), .ZN(n12463) );
  AOI21_X1 U7986 ( .B1(n12368), .B2(n12367), .A(n6918), .ZN(n6917) );
  OR2_X1 U7987 ( .A1(n8817), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8842) );
  NAND2_X1 U7988 ( .A1(n8815), .A2(n7864), .ZN(n14817) );
  NOR2_X1 U7989 ( .A1(n14814), .A2(n7865), .ZN(n7864) );
  INV_X1 U7990 ( .A(n9302), .ZN(n7865) );
  AOI21_X1 U7991 ( .B1(n7869), .B2(n7871), .A(n7867), .ZN(n7866) );
  INV_X1 U7992 ( .A(n9297), .ZN(n7867) );
  NAND2_X1 U7993 ( .A1(n15320), .A2(n9288), .ZN(n15316) );
  NAND2_X1 U7994 ( .A1(n15316), .A2(n15315), .ZN(n15314) );
  NAND2_X1 U7995 ( .A1(n11422), .A2(n6799), .ZN(n11694) );
  NOR2_X1 U7996 ( .A1(n11697), .A2(n6800), .ZN(n6799) );
  INV_X1 U7997 ( .A(n9121), .ZN(n6800) );
  NAND2_X1 U7998 ( .A1(n11691), .A2(n8714), .ZN(n11423) );
  INV_X1 U7999 ( .A(n11393), .ZN(n15354) );
  NAND2_X1 U8000 ( .A1(n12651), .A2(n9234), .ZN(n7390) );
  NAND2_X1 U8001 ( .A1(n8980), .A2(n8979), .ZN(n13289) );
  NAND2_X1 U8002 ( .A1(n11687), .A2(n11683), .ZN(n15353) );
  OAI21_X1 U8003 ( .B1(n9211), .B2(n9210), .A(n9209), .ZN(n9231) );
  NAND2_X1 U8004 ( .A1(n7019), .A2(n9059), .ZN(n9073) );
  NAND2_X1 U8005 ( .A1(n9058), .A2(n9057), .ZN(n7019) );
  NAND2_X1 U8006 ( .A1(n9006), .A2(n9005), .ZN(n9016) );
  OR2_X1 U8007 ( .A1(n9093), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n9095) );
  AND2_X1 U8008 ( .A1(n8963), .A2(n15717), .ZN(n9090) );
  INV_X1 U8009 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9089) );
  AND2_X1 U8010 ( .A1(n8922), .A2(n8906), .ZN(n8907) );
  AOI21_X1 U8011 ( .B1(n8903), .B2(n7382), .A(n7381), .ZN(n7380) );
  INV_X1 U8012 ( .A(n8905), .ZN(n7381) );
  INV_X1 U8013 ( .A(n8887), .ZN(n7382) );
  AND2_X1 U8014 ( .A1(n8887), .A2(n8874), .ZN(n8875) );
  INV_X1 U8016 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8877) );
  OR2_X1 U8017 ( .A1(n8858), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8890) );
  AND2_X1 U8018 ( .A1(n8851), .A2(n8833), .ZN(n8848) );
  NAND2_X1 U8019 ( .A1(n6991), .A2(n6990), .ZN(n8850) );
  AOI21_X1 U8020 ( .B1(n6992), .B2(n7386), .A(n6713), .ZN(n6990) );
  NAND2_X1 U8021 ( .A1(n8797), .A2(n6992), .ZN(n6991) );
  AND2_X1 U8022 ( .A1(n7383), .A2(n6995), .ZN(n6994) );
  NAND2_X1 U8023 ( .A1(n7385), .A2(n6996), .ZN(n6995) );
  AOI21_X1 U8024 ( .B1(n7385), .B2(n7387), .A(n6656), .ZN(n7383) );
  INV_X1 U8025 ( .A(n15707), .ZN(n6996) );
  XNOR2_X1 U8026 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8794) );
  NAND2_X1 U8027 ( .A1(n6988), .A2(n8745), .ZN(n8760) );
  XNOR2_X1 U8028 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8723) );
  INV_X1 U8029 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7689) );
  XNOR2_X1 U8030 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8667) );
  NAND2_X1 U8031 ( .A1(n8385), .A2(n7643), .ZN(n7642) );
  NOR2_X1 U8032 ( .A1(n13439), .A2(n7644), .ZN(n7643) );
  INV_X1 U8033 ( .A(n11525), .ZN(n7616) );
  NAND2_X1 U8034 ( .A1(n7634), .A2(n6641), .ZN(n6997) );
  INV_X1 U8035 ( .A(n7639), .ZN(n6999) );
  OAI211_X1 U8036 ( .C1(n7005), .C2(n7004), .A(n7002), .B(n8304), .ZN(n7620)
         );
  XNOR2_X1 U8037 ( .A(n8480), .B(n8479), .ZN(n12539) );
  AND2_X1 U8038 ( .A1(n7006), .A2(n8269), .ZN(n7005) );
  INV_X1 U8039 ( .A(n11931), .ZN(n7006) );
  AND2_X1 U8040 ( .A1(n9667), .A2(n8080), .ZN(n10415) );
  AOI21_X1 U8041 ( .B1(n9649), .B2(n9645), .A(n9644), .ZN(n9658) );
  OR2_X1 U8042 ( .A1(n9650), .A2(n6690), .ZN(n6811) );
  OAI22_X1 U8043 ( .A1(n8137), .A2(P2_REG3_REG_3__SCAN_IN), .B1(n8138), .B2(
        n12049), .ZN(n6889) );
  OAI22_X1 U8044 ( .A1(n8137), .A2(n11780), .B1(n10437), .B2(n8138), .ZN(n6986) );
  AOI21_X1 U8045 ( .B1(n7905), .B2(n7904), .A(n7975), .ZN(n7906) );
  NAND2_X1 U8046 ( .A1(n13949), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7905) );
  OR2_X1 U8047 ( .A1(n13949), .A2(n11418), .ZN(n7904) );
  XNOR2_X1 U8048 ( .A(n13531), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n13537) );
  AOI21_X1 U8049 ( .B1(n10454), .B2(n10440), .A(n10439), .ZN(n6744) );
  NOR2_X1 U8050 ( .A1(n10668), .A2(n6748), .ZN(n10679) );
  AND2_X1 U8051 ( .A1(n10669), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6748) );
  INV_X1 U8052 ( .A(n9786), .ZN(n13611) );
  AOI21_X1 U8053 ( .B1(n13651), .B2(n9781), .A(n9780), .ZN(n13640) );
  OR2_X1 U8054 ( .A1(n13677), .A2(n13685), .ZN(n7782) );
  NAND2_X1 U8055 ( .A1(n13654), .A2(n13653), .ZN(n13652) );
  AOI21_X1 U8056 ( .B1(n7599), .B2(n7597), .A(n6610), .ZN(n7596) );
  INV_X1 U8057 ( .A(n9776), .ZN(n7597) );
  OR2_X1 U8058 ( .A1(n13727), .A2(n7598), .ZN(n6884) );
  AOI21_X1 U8059 ( .B1(n7596), .B2(n7598), .A(n6886), .ZN(n6885) );
  INV_X1 U8060 ( .A(n13689), .ZN(n6886) );
  NAND2_X1 U8061 ( .A1(n13702), .A2(n9726), .ZN(n13683) );
  NOR2_X1 U8062 ( .A1(n13700), .A2(n7600), .ZN(n7599) );
  AND2_X1 U8063 ( .A1(n13726), .A2(n9776), .ZN(n7600) );
  NOR2_X1 U8064 ( .A1(n13893), .A2(n13468), .ZN(n7792) );
  NAND2_X1 U8065 ( .A1(n13739), .A2(n13740), .ZN(n13738) );
  INV_X1 U8066 ( .A(n9722), .ZN(n13740) );
  AOI21_X1 U8067 ( .B1(n6562), .B2(n7601), .A(n13760), .ZN(n6910) );
  INV_X1 U8068 ( .A(n7302), .ZN(n7301) );
  OAI21_X1 U8069 ( .B1(n7303), .B2(n9719), .A(n7309), .ZN(n7302) );
  NAND2_X1 U8070 ( .A1(n13907), .A2(n13502), .ZN(n7309) );
  NAND2_X1 U8071 ( .A1(n9765), .A2(n7606), .ZN(n13793) );
  OR2_X1 U8072 ( .A1(n12236), .A2(n15114), .ZN(n7951) );
  NAND2_X1 U8073 ( .A1(n12229), .A2(n6976), .ZN(n6975) );
  OR2_X1 U8074 ( .A1(n12420), .A2(n12443), .ZN(n6976) );
  NOR2_X1 U8075 ( .A1(n8279), .A2(n8278), .ZN(n8317) );
  OAI22_X1 U8076 ( .A1(n12125), .A2(n9756), .B1(n12214), .B2(n15112), .ZN(
        n12243) );
  NAND2_X1 U8077 ( .A1(n12074), .A2(n12073), .ZN(n12076) );
  AND2_X1 U8078 ( .A1(n7803), .A2(n9715), .ZN(n7802) );
  NAND2_X1 U8079 ( .A1(n11844), .A2(n9714), .ZN(n7804) );
  NAND2_X1 U8080 ( .A1(n6877), .A2(n9749), .ZN(n11842) );
  NAND2_X1 U8081 ( .A1(n6878), .A2(n9744), .ZN(n11823) );
  NAND2_X1 U8082 ( .A1(n8148), .A2(n10479), .ZN(n7007) );
  CLKBUF_X1 U8083 ( .A(n8097), .Z(n13690) );
  OR2_X1 U8084 ( .A1(n11758), .A2(n6555), .ZN(n11824) );
  NAND2_X1 U8085 ( .A1(n9617), .A2(n9732), .ZN(n13819) );
  NAND2_X1 U8086 ( .A1(n9784), .A2(n6592), .ZN(n13848) );
  XNOR2_X1 U8087 ( .A(n9667), .B(n11758), .ZN(n7615) );
  NAND2_X1 U8088 ( .A1(n8057), .A2(n8056), .ZN(n8470) );
  INV_X1 U8089 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8312) );
  NAND2_X1 U8090 ( .A1(n9973), .A2(n9972), .ZN(n11734) );
  NAND2_X1 U8091 ( .A1(n7854), .A2(n12291), .ZN(n7851) );
  NAND2_X1 U8092 ( .A1(n6943), .A2(n6630), .ZN(n6942) );
  INV_X1 U8093 ( .A(n7852), .ZN(n6943) );
  NOR2_X1 U8094 ( .A1(n7852), .A2(n6945), .ZN(n6944) );
  INV_X1 U8095 ( .A(n11645), .ZN(n6945) );
  AND2_X1 U8096 ( .A1(n7814), .A2(n13998), .ZN(n7813) );
  NAND2_X1 U8097 ( .A1(n7816), .A2(n7818), .ZN(n7814) );
  AND2_X1 U8098 ( .A1(n7834), .A2(n14008), .ZN(n7833) );
  NAND2_X1 U8099 ( .A1(n7835), .A2(n14034), .ZN(n7834) );
  INV_X1 U8100 ( .A(n6953), .ZN(n11177) );
  AOI22_X1 U8101 ( .A1(n12743), .A2(n11134), .B1(n11137), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n6952) );
  NAND2_X1 U8102 ( .A1(n11177), .A2(n11176), .ZN(n11175) );
  INV_X1 U8103 ( .A(n12709), .ZN(n7824) );
  NOR2_X1 U8104 ( .A1(n12477), .A2(n12478), .ZN(n7844) );
  OAI22_X1 U8105 ( .A1(n11143), .A2(n11135), .B1(n11144), .B2(n12779), .ZN(
        n11142) );
  AND4_X1 U8106 ( .A1(n10247), .A2(n10246), .A3(n10245), .A4(n10244), .ZN(
        n14076) );
  AND4_X1 U8107 ( .A1(n9934), .A2(n9933), .A3(n9932), .A4(n9931), .ZN(n11595)
         );
  OR2_X1 U8108 ( .A1(n14299), .A2(n7364), .ZN(n7363) );
  OR2_X1 U8109 ( .A1(n7366), .A2(n12566), .ZN(n7362) );
  NAND2_X1 U8110 ( .A1(n7369), .A2(n12565), .ZN(n7364) );
  AND2_X1 U8111 ( .A1(n14308), .A2(n12593), .ZN(n14291) );
  INV_X1 U8112 ( .A(n6872), .ZN(n14324) );
  OAI21_X1 U8113 ( .B1(n14342), .B2(n12589), .A(n12590), .ZN(n6872) );
  AND2_X1 U8114 ( .A1(n7699), .A2(n14344), .ZN(n7698) );
  OR2_X1 U8115 ( .A1(n7700), .A2(n7705), .ZN(n7699) );
  XNOR2_X1 U8116 ( .A(n14060), .B(n10309), .ZN(n14362) );
  NAND2_X1 U8117 ( .A1(n7109), .A2(n12562), .ZN(n14356) );
  NAND2_X1 U8118 ( .A1(n14388), .A2(n7476), .ZN(n14373) );
  NAND2_X1 U8119 ( .A1(n12559), .A2(n7732), .ZN(n7731) );
  NOR2_X1 U8120 ( .A1(n14406), .A2(n7733), .ZN(n7732) );
  INV_X1 U8121 ( .A(n12558), .ZN(n7733) );
  NAND2_X1 U8122 ( .A1(n7731), .A2(n7730), .ZN(n14390) );
  AND2_X1 U8123 ( .A1(n12586), .A2(n12560), .ZN(n7730) );
  OR2_X1 U8124 ( .A1(n14387), .A2(n12586), .ZN(n14388) );
  AND2_X1 U8125 ( .A1(n7460), .A2(n12582), .ZN(n7459) );
  OR2_X1 U8126 ( .A1(n12583), .A2(n7461), .ZN(n7460) );
  NAND2_X1 U8127 ( .A1(n12578), .A2(n12579), .ZN(n7461) );
  NAND2_X1 U8128 ( .A1(n12580), .A2(n12579), .ZN(n7457) );
  NAND2_X1 U8129 ( .A1(n14423), .A2(n14420), .ZN(n12559) );
  NAND2_X1 U8130 ( .A1(n6849), .A2(n12577), .ZN(n14438) );
  NAND2_X1 U8131 ( .A1(n6855), .A2(n6854), .ZN(n6849) );
  AND2_X1 U8132 ( .A1(n10121), .A2(n10120), .ZN(n14463) );
  NAND2_X1 U8133 ( .A1(n12555), .A2(n12554), .ZN(n14456) );
  INV_X1 U8134 ( .A(n14475), .ZN(n14489) );
  NOR2_X1 U8135 ( .A1(n14489), .A2(n7465), .ZN(n7464) );
  INV_X1 U8136 ( .A(n12575), .ZN(n7465) );
  NAND2_X1 U8137 ( .A1(n10074), .A2(n10073), .ZN(n12672) );
  NAND2_X1 U8138 ( .A1(n12265), .A2(n12259), .ZN(n12576) );
  NOR2_X1 U8139 ( .A1(n12032), .A2(n7469), .ZN(n7468) );
  INV_X1 U8140 ( .A(n12026), .ZN(n7469) );
  NAND2_X1 U8141 ( .A1(n14883), .A2(n12031), .ZN(n7719) );
  NAND2_X1 U8142 ( .A1(n6858), .A2(n12025), .ZN(n14890) );
  NAND2_X1 U8143 ( .A1(n12024), .A2(n12023), .ZN(n6858) );
  NOR2_X1 U8144 ( .A1(n11941), .A2(n7722), .ZN(n7721) );
  INV_X1 U8145 ( .A(n11885), .ZN(n7722) );
  AND2_X1 U8146 ( .A1(n11885), .A2(n10311), .ZN(n11722) );
  AND2_X1 U8147 ( .A1(n7430), .A2(n7434), .ZN(n6845) );
  NAND2_X1 U8148 ( .A1(n11584), .A2(n7430), .ZN(n6847) );
  AND2_X1 U8149 ( .A1(n9938), .A2(n9937), .ZN(n15008) );
  NAND2_X1 U8150 ( .A1(n11334), .A2(n11317), .ZN(n11586) );
  NOR2_X1 U8151 ( .A1(n11588), .A2(n11583), .ZN(n7436) );
  INV_X1 U8152 ( .A(n7435), .ZN(n7434) );
  AND2_X1 U8153 ( .A1(n12777), .A2(n10710), .ZN(n11306) );
  XNOR2_X1 U8154 ( .A(n14933), .B(n14108), .ZN(n11335) );
  INV_X1 U8155 ( .A(n14933), .ZN(n11478) );
  OR2_X1 U8156 ( .A1(n14110), .A2(n11143), .ZN(n11112) );
  INV_X1 U8157 ( .A(n14462), .ZN(n14479) );
  NAND2_X1 U8158 ( .A1(n10138), .A2(n10137), .ZN(n14574) );
  NAND2_X1 U8159 ( .A1(n10130), .A2(n10129), .ZN(n14580) );
  INV_X1 U8160 ( .A(n15052), .ZN(n15002) );
  XNOR2_X1 U8161 ( .A(n9598), .B(n9597), .ZN(n13942) );
  AOI21_X1 U8162 ( .B1(n9623), .B2(n9622), .A(n9592), .ZN(n9606) );
  OR2_X1 U8163 ( .A1(n14616), .A2(n14617), .ZN(n9821) );
  XNOR2_X1 U8164 ( .A(n9823), .B(P1_IR_REG_29__SCAN_IN), .ZN(n9825) );
  NAND2_X1 U8165 ( .A1(n14617), .A2(n9819), .ZN(n6870) );
  NAND2_X1 U8166 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n6871) );
  NOR2_X1 U8167 ( .A1(n7737), .A2(n14617), .ZN(n7146) );
  AND2_X1 U8168 ( .A1(n8503), .A2(n8502), .ZN(n13965) );
  NAND2_X1 U8169 ( .A1(n8065), .A2(n8064), .ZN(n8501) );
  AND2_X1 U8170 ( .A1(n8054), .A2(n8055), .ZN(n7750) );
  OAI21_X1 U8171 ( .B1(n9839), .B2(n6655), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9842) );
  NAND2_X1 U8172 ( .A1(n9837), .A2(n6638), .ZN(n10366) );
  AND2_X1 U8173 ( .A1(n7776), .A2(n8307), .ZN(n8329) );
  NAND2_X1 U8174 ( .A1(n8306), .A2(n8034), .ZN(n7776) );
  XNOR2_X1 U8175 ( .A(n7048), .B(SI_10_), .ZN(n10565) );
  NAND2_X1 U8176 ( .A1(n7946), .A2(n8270), .ZN(n7048) );
  NAND2_X1 U8177 ( .A1(n7349), .A2(n8028), .ZN(n8270) );
  OR2_X1 U8178 ( .A1(n7349), .A2(n8028), .ZN(n7946) );
  INV_X1 U8179 ( .A(SI_9_), .ZN(n8024) );
  OR2_X1 U8180 ( .A1(n7661), .A2(n14737), .ZN(n7660) );
  AOI21_X1 U8181 ( .B1(n14739), .B2(n14738), .A(n7662), .ZN(n7661) );
  XNOR2_X1 U8182 ( .A(n14682), .B(n7225), .ZN(n14683) );
  INV_X1 U8183 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7225) );
  NAND2_X1 U8184 ( .A1(n15737), .A2(n14699), .ZN(n14700) );
  NAND2_X1 U8185 ( .A1(n14769), .A2(n14712), .ZN(n14714) );
  XNOR2_X1 U8186 ( .A(n14658), .B(n14657), .ZN(n14715) );
  NAND2_X1 U8187 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7656) );
  XNOR2_X1 U8188 ( .A(n14714), .B(n7036), .ZN(n7125) );
  INV_X1 U8189 ( .A(n14713), .ZN(n7036) );
  AOI21_X1 U8190 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n14662), .A(n14661), .ZN(
        n14679) );
  NOR2_X1 U8191 ( .A1(n14717), .A2(n14716), .ZN(n14661) );
  AND2_X1 U8192 ( .A1(n7026), .A2(n14921), .ZN(n14726) );
  OAI21_X1 U8193 ( .B1(n14922), .B2(n14923), .A(n7649), .ZN(n7026) );
  INV_X1 U8194 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7649) );
  OR2_X1 U8195 ( .A1(n7030), .A2(n14789), .ZN(n7650) );
  INV_X1 U8196 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7651) );
  OR2_X1 U8197 ( .A1(n14732), .A2(n14731), .ZN(n14797) );
  AND2_X1 U8198 ( .A1(n7082), .A2(n6692), .ZN(n7080) );
  AND2_X1 U8199 ( .A1(n7083), .A2(n12861), .ZN(n7082) );
  OAI22_X1 U8200 ( .A1(n12796), .A2(n6564), .B1(n12797), .B2(n7084), .ZN(n7083) );
  NOR2_X1 U8201 ( .A1(n12888), .A2(n6564), .ZN(n7084) );
  AND2_X1 U8202 ( .A1(n9042), .A2(n9041), .ZN(n13131) );
  NAND2_X1 U8203 ( .A1(n9019), .A2(n9018), .ZN(n12808) );
  NAND2_X1 U8204 ( .A1(n7402), .A2(n7406), .ZN(n7400) );
  NAND2_X1 U8205 ( .A1(n7407), .A2(n7409), .ZN(n7406) );
  INV_X1 U8206 ( .A(n7410), .ZN(n7407) );
  NAND2_X1 U8207 ( .A1(n7416), .A2(n12635), .ZN(n12826) );
  NAND2_X1 U8208 ( .A1(n12853), .A2(n12854), .ZN(n7416) );
  AND3_X1 U8209 ( .A1(n8733), .A2(n8732), .A3(n8731), .ZN(n11746) );
  INV_X1 U8210 ( .A(n13363), .ZN(n12850) );
  INV_X1 U8211 ( .A(n13171), .ZN(n12871) );
  INV_X1 U8212 ( .A(n13147), .ZN(n13280) );
  AND2_X1 U8213 ( .A1(n11278), .A2(n11285), .ZN(n11279) );
  AOI21_X1 U8214 ( .B1(n7417), .B2(n7419), .A(n6650), .ZN(n7414) );
  AND2_X1 U8215 ( .A1(n10952), .A2(n10951), .ZN(n15425) );
  NAND2_X1 U8216 ( .A1(n12518), .A2(n12517), .ZN(n12611) );
  NAND2_X1 U8217 ( .A1(n8893), .A2(n8892), .ZN(n13248) );
  OAI211_X1 U8218 ( .C1(n8699), .C2(n13032), .A(n8975), .B(n8974), .ZN(n13172)
         );
  NAND4_X1 U8219 ( .A1(n8742), .A2(n8741), .A3(n8740), .A4(n8739), .ZN(n15331)
         );
  INV_X1 U8220 ( .A(n11699), .ZN(n15421) );
  XNOR2_X1 U8221 ( .A(n8747), .B(P3_IR_REG_6__SCAN_IN), .ZN(n11210) );
  INV_X1 U8222 ( .A(n7684), .ZN(n11555) );
  NOR2_X1 U8223 ( .A1(n11547), .A2(n11546), .ZN(n11549) );
  NAND2_X1 U8224 ( .A1(n6756), .A2(n6755), .ZN(n7686) );
  INV_X1 U8225 ( .A(n7489), .ZN(n11917) );
  OR2_X1 U8226 ( .A1(n12347), .A2(n8819), .ZN(n7196) );
  INV_X1 U8227 ( .A(n7241), .ZN(n12382) );
  XNOR2_X1 U8228 ( .A(n7185), .B(n14760), .ZN(n12347) );
  OR2_X1 U8229 ( .A1(n12903), .A2(n8862), .ZN(n6778) );
  INV_X1 U8230 ( .A(n7240), .ZN(n12930) );
  XNOR2_X1 U8231 ( .A(n12919), .B(n12929), .ZN(n12903) );
  NAND2_X1 U8232 ( .A1(n6965), .A2(n13003), .ZN(n6966) );
  NAND2_X1 U8233 ( .A1(n6967), .A2(n13007), .ZN(n13023) );
  NOR2_X1 U8234 ( .A1(n13002), .A2(n7114), .ZN(n7113) );
  NAND2_X1 U8235 ( .A1(n7233), .A2(n7115), .ZN(n7114) );
  NAND2_X1 U8236 ( .A1(n13041), .A2(n13003), .ZN(n7115) );
  NAND2_X1 U8237 ( .A1(n13019), .A2(n13018), .ZN(n7135) );
  AND2_X1 U8238 ( .A1(n7669), .A2(n7671), .ZN(n13019) );
  OR2_X1 U8239 ( .A1(n13020), .A2(n6720), .ZN(n7134) );
  NAND2_X1 U8240 ( .A1(n12993), .A2(n7672), .ZN(n7671) );
  NOR2_X1 U8241 ( .A1(n13015), .A2(n13223), .ZN(n7672) );
  NAND2_X1 U8242 ( .A1(n7175), .A2(n6721), .ZN(n6766) );
  NOR2_X1 U8243 ( .A1(n6732), .A2(n7132), .ZN(n7131) );
  NOR2_X1 U8244 ( .A1(n13029), .A2(n6614), .ZN(n13035) );
  INV_X1 U8245 ( .A(n6769), .ZN(n6768) );
  OAI211_X1 U8246 ( .C1(n7671), .C2(n13038), .A(n7666), .B(n12995), .ZN(n6769)
         );
  OAI21_X1 U8247 ( .B1(n13013), .B2(n13037), .A(n7664), .ZN(n7666) );
  INV_X1 U8248 ( .A(n7665), .ZN(n7664) );
  NAND2_X1 U8249 ( .A1(n13073), .A2(n6785), .ZN(n13262) );
  NOR2_X1 U8250 ( .A1(n6700), .A2(n6786), .ZN(n6785) );
  NAND2_X1 U8251 ( .A1(n9146), .A2(n7160), .ZN(n13080) );
  NAND2_X1 U8252 ( .A1(n6570), .A2(n10380), .ZN(n7160) );
  OR2_X1 U8253 ( .A1(n8722), .A2(n12503), .ZN(n9076) );
  NOR2_X1 U8254 ( .A1(n10390), .A2(n10389), .ZN(n10391) );
  INV_X1 U8255 ( .A(n15405), .ZN(n10389) );
  INV_X1 U8256 ( .A(n13064), .ZN(n10390) );
  NOR2_X1 U8257 ( .A1(n13262), .A2(n6784), .ZN(n13326) );
  AND2_X1 U8258 ( .A1(n13263), .A2(n15405), .ZN(n6784) );
  NAND2_X1 U8259 ( .A1(n8996), .A2(n8995), .ZN(n13349) );
  OR2_X1 U8260 ( .A1(n8722), .A2(n11601), .ZN(n8995) );
  AND2_X1 U8261 ( .A1(n8915), .A2(n8914), .ZN(n13367) );
  AND2_X1 U8262 ( .A1(n9158), .A2(n9157), .ZN(n13379) );
  OR2_X1 U8263 ( .A1(n10520), .A2(P3_D_REG_0__SCAN_IN), .ZN(n9158) );
  XNOR2_X1 U8264 ( .A(n8662), .B(n8661), .ZN(n12652) );
  OR2_X1 U8265 ( .A1(n8656), .A2(n8660), .ZN(n8662) );
  MUX2_X1 U8266 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8657), .S(
        P3_IR_REG_27__SCAN_IN), .Z(n8658) );
  NAND2_X1 U8267 ( .A1(n6842), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8657) );
  NAND2_X1 U8268 ( .A1(n13390), .A2(n13391), .ZN(n7203) );
  NAND2_X1 U8269 ( .A1(n13483), .A2(n7631), .ZN(n13390) );
  INV_X1 U8270 ( .A(n14840), .ZN(n7164) );
  NAND2_X1 U8271 ( .A1(n10512), .A2(n8148), .ZN(n7320) );
  OR2_X1 U8272 ( .A1(n8415), .A2(n9791), .ZN(n8106) );
  NAND2_X1 U8273 ( .A1(n8091), .A2(n8090), .ZN(n13879) );
  NAND2_X1 U8274 ( .A1(n8414), .A2(n8413), .ZN(n13903) );
  NAND2_X1 U8275 ( .A1(n7151), .A2(n8488), .ZN(n7150) );
  INV_X1 U8276 ( .A(n8499), .ZN(n7151) );
  NAND2_X1 U8277 ( .A1(n8455), .A2(n8454), .ZN(n13887) );
  OR2_X1 U8278 ( .A1(n8139), .A2(n8117), .ZN(n8119) );
  OR2_X1 U8279 ( .A1(n8137), .A2(n13528), .ZN(n8118) );
  NAND2_X1 U8280 ( .A1(n11348), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15124) );
  CLKBUF_X1 U8281 ( .A(n13506), .Z(n14848) );
  INV_X1 U8282 ( .A(n8079), .ZN(n9789) );
  OAI21_X1 U8283 ( .B1(n13720), .B2(n8137), .A(n8096), .ZN(n13742) );
  NAND2_X1 U8284 ( .A1(n15161), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n15160) );
  XNOR2_X1 U8285 ( .A(n13555), .B(n13568), .ZN(n15171) );
  NAND2_X1 U8286 ( .A1(n15171), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n15170) );
  OR2_X1 U8287 ( .A1(n13559), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6746) );
  XNOR2_X1 U8288 ( .A(n13578), .B(n13581), .ZN(n13559) );
  NAND2_X1 U8289 ( .A1(n8538), .A2(n8537), .ZN(n13849) );
  AND2_X1 U8290 ( .A1(n13770), .A2(n6555), .ZN(n13835) );
  AND2_X1 U8291 ( .A1(n12603), .A2(n15251), .ZN(n7751) );
  XNOR2_X1 U8292 ( .A(n9731), .B(n9788), .ZN(n7791) );
  OAI21_X1 U8293 ( .B1(n7790), .B2(n15277), .A(n7789), .ZN(n7787) );
  NAND2_X1 U8294 ( .A1(n15277), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7789) );
  NAND2_X1 U8295 ( .A1(n9795), .A2(n9794), .ZN(n6908) );
  AND2_X1 U8296 ( .A1(n10550), .A2(n10554), .ZN(n10369) );
  OAI21_X1 U8297 ( .B1(n14072), .B2(n12767), .A(n7810), .ZN(n13970) );
  NAND2_X1 U8298 ( .A1(n11476), .A2(n7831), .ZN(n14939) );
  AND2_X1 U8299 ( .A1(n11485), .A2(n11475), .ZN(n7831) );
  NAND2_X1 U8300 ( .A1(n10104), .A2(n10103), .ZN(n14591) );
  NAND2_X1 U8301 ( .A1(n14641), .A2(n10563), .ZN(n14060) );
  INV_X1 U8302 ( .A(n14935), .ZN(n14961) );
  OAI21_X1 U8303 ( .B1(n7226), .B2(n7058), .A(n7056), .ZN(n7053) );
  NAND2_X1 U8304 ( .A1(n10306), .A2(n10357), .ZN(n7058) );
  INV_X1 U8305 ( .A(n7057), .ZN(n7056) );
  OAI21_X1 U8306 ( .B1(n6572), .B2(n12372), .A(n10376), .ZN(n7057) );
  NAND2_X1 U8307 ( .A1(n10338), .A2(n10337), .ZN(n10353) );
  INV_X1 U8308 ( .A(n13992), .ZN(n14409) );
  NAND2_X1 U8309 ( .A1(n10173), .A2(n10172), .ZN(n14381) );
  NAND2_X1 U8310 ( .A1(n10004), .A2(n10003), .ZN(n14952) );
  NAND2_X1 U8311 ( .A1(n9886), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7437) );
  NAND2_X1 U8312 ( .A1(n10136), .A2(n14129), .ZN(n7438) );
  NAND2_X1 U8313 ( .A1(n7447), .A2(n7168), .ZN(n14515) );
  NAND2_X1 U8314 ( .A1(n7169), .A2(n14257), .ZN(n7168) );
  NAND2_X1 U8315 ( .A1(n7944), .A2(n14514), .ZN(n7371) );
  OAI21_X1 U8316 ( .B1(n14525), .B2(n15055), .A(n14523), .ZN(n7728) );
  NOR2_X1 U8317 ( .A1(n15742), .A2(n15743), .ZN(n15741) );
  INV_X1 U8318 ( .A(n7125), .ZN(n14772) );
  OR2_X1 U8319 ( .A1(n14772), .A2(n7658), .ZN(n7655) );
  OR2_X1 U8320 ( .A1(n14772), .A2(n14773), .ZN(n7659) );
  NOR2_X1 U8321 ( .A1(n6581), .A2(n14912), .ZN(n14911) );
  INV_X1 U8322 ( .A(n14911), .ZN(n7034) );
  NAND2_X1 U8323 ( .A1(n14718), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7035) );
  XNOR2_X1 U8324 ( .A(n7652), .B(n14723), .ZN(n14920) );
  NAND2_X1 U8325 ( .A1(n14920), .A2(n14919), .ZN(n14918) );
  NAND2_X1 U8326 ( .A1(n7123), .A2(n7122), .ZN(n14927) );
  INV_X1 U8327 ( .A(n14725), .ZN(n7122) );
  INV_X1 U8328 ( .A(n14726), .ZN(n7123) );
  NOR2_X1 U8329 ( .A1(n14790), .A2(n14791), .ZN(n14789) );
  NAND2_X1 U8330 ( .A1(n7609), .A2(n9653), .ZN(n9418) );
  INV_X1 U8331 ( .A(n11106), .ZN(n10316) );
  OAI21_X1 U8332 ( .B1(n10283), .B2(n11588), .A(n7108), .ZN(n9926) );
  NAND2_X1 U8333 ( .A1(n10283), .A2(n11587), .ZN(n7108) );
  NOR2_X1 U8334 ( .A1(n9444), .A2(n9445), .ZN(n7256) );
  NOR2_X1 U8335 ( .A1(n9447), .A2(n9446), .ZN(n7260) );
  INV_X1 U8336 ( .A(n9444), .ZN(n7258) );
  INV_X1 U8337 ( .A(n9445), .ZN(n7262) );
  NAND2_X1 U8338 ( .A1(n7554), .A2(n7553), .ZN(n9943) );
  INV_X1 U8339 ( .A(n7550), .ZN(n7552) );
  INV_X1 U8340 ( .A(n9482), .ZN(n7255) );
  NOR2_X1 U8341 ( .A1(n7255), .A2(n9483), .ZN(n7252) );
  NAND2_X1 U8342 ( .A1(n10005), .A2(n7566), .ZN(n7565) );
  INV_X1 U8343 ( .A(n10007), .ZN(n7566) );
  INV_X1 U8344 ( .A(n10018), .ZN(n7220) );
  INV_X1 U8345 ( .A(n9987), .ZN(n7215) );
  AND2_X1 U8346 ( .A1(n10007), .A2(n7568), .ZN(n7567) );
  NAND2_X1 U8347 ( .A1(n7275), .A2(n7274), .ZN(n9501) );
  AND2_X1 U8348 ( .A1(n9492), .A2(n7279), .ZN(n7278) );
  NAND2_X1 U8349 ( .A1(n7038), .A2(n6634), .ZN(n10054) );
  OAI21_X1 U8350 ( .B1(n10033), .B2(n7571), .A(n6653), .ZN(n10056) );
  INV_X1 U8351 ( .A(n10055), .ZN(n7216) );
  NAND2_X1 U8352 ( .A1(n10069), .A2(n10070), .ZN(n7063) );
  NAND2_X1 U8353 ( .A1(n10092), .A2(n10301), .ZN(n7119) );
  INV_X1 U8354 ( .A(n9509), .ZN(n7266) );
  INV_X1 U8355 ( .A(n10106), .ZN(n7228) );
  NAND2_X1 U8356 ( .A1(n7926), .A2(n7923), .ZN(n9520) );
  NAND2_X1 U8357 ( .A1(n7925), .A2(n7924), .ZN(n7923) );
  INV_X1 U8358 ( .A(n9512), .ZN(n7924) );
  NOR2_X1 U8359 ( .A1(n10165), .A2(n7589), .ZN(n7588) );
  INV_X1 U8360 ( .A(n10154), .ZN(n7589) );
  OAI22_X1 U8361 ( .A1(n9530), .A2(n7908), .B1(n9529), .B2(n9528), .ZN(n9538)
         );
  NOR2_X1 U8362 ( .A1(n7909), .A2(n7910), .ZN(n7908) );
  NAND2_X1 U8363 ( .A1(n9538), .A2(n9537), .ZN(n9536) );
  AND2_X1 U8364 ( .A1(n9546), .A2(n7916), .ZN(n7915) );
  NAND2_X1 U8365 ( .A1(n7919), .A2(n7918), .ZN(n7916) );
  NAND2_X1 U8366 ( .A1(n6598), .A2(n7920), .ZN(n7918) );
  NAND2_X1 U8367 ( .A1(n7072), .A2(n10174), .ZN(n7071) );
  INV_X1 U8368 ( .A(n9568), .ZN(n7296) );
  NOR2_X1 U8369 ( .A1(n6599), .A2(n7935), .ZN(n7934) );
  AND2_X1 U8370 ( .A1(n9555), .A2(n9554), .ZN(n7280) );
  AND2_X1 U8371 ( .A1(n10219), .A2(n7558), .ZN(n7227) );
  AOI21_X1 U8372 ( .B1(n7557), .B2(n6627), .A(n7050), .ZN(n7049) );
  INV_X1 U8373 ( .A(n10217), .ZN(n7050) );
  AND2_X1 U8374 ( .A1(n7690), .A2(n11335), .ZN(n10318) );
  NOR2_X1 U8375 ( .A1(n8060), .A2(n8468), .ZN(n6827) );
  AOI21_X1 U8376 ( .B1(n7772), .B2(n6568), .A(n6666), .ZN(n7771) );
  AOI21_X1 U8377 ( .B1(n7779), .B2(SI_13_), .A(n8327), .ZN(n7777) );
  NOR2_X1 U8378 ( .A1(n7779), .A2(SI_13_), .ZN(n7775) );
  OR2_X1 U8379 ( .A1(n9056), .A2(n7890), .ZN(n7889) );
  INV_X1 U8380 ( .A(n9252), .ZN(n7890) );
  AND2_X1 U8381 ( .A1(n13175), .A2(n6791), .ZN(n6790) );
  NAND2_X1 U8382 ( .A1(n9383), .A2(n9142), .ZN(n6791) );
  INV_X1 U8383 ( .A(n9576), .ZN(n7930) );
  INV_X1 U8384 ( .A(n7288), .ZN(n7287) );
  OAI21_X1 U8385 ( .B1(n7291), .B2(n9572), .A(n7289), .ZN(n7288) );
  NAND2_X1 U8386 ( .A1(n8073), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8070) );
  INV_X1 U8387 ( .A(n13843), .ZN(n7754) );
  NOR2_X1 U8388 ( .A1(n7562), .A2(n7561), .ZN(n10235) );
  AOI21_X1 U8389 ( .B1(n10231), .B2(n10230), .A(n7563), .ZN(n7562) );
  NAND2_X1 U8390 ( .A1(n7704), .A2(n7361), .ZN(n7360) );
  INV_X1 U8391 ( .A(n12563), .ZN(n7361) );
  NOR2_X1 U8392 ( .A1(n14415), .A2(n7457), .ZN(n7456) );
  NOR2_X1 U8393 ( .A1(n7745), .A2(n9588), .ZN(n6819) );
  INV_X1 U8394 ( .A(n8503), .ZN(n6817) );
  NAND2_X1 U8395 ( .A1(n6821), .A2(n6824), .ZN(n6820) );
  INV_X1 U8396 ( .A(n7768), .ZN(n6821) );
  NOR2_X1 U8397 ( .A1(n8050), .A2(SI_19_), .ZN(n7764) );
  NOR2_X1 U8398 ( .A1(n8445), .A2(n8427), .ZN(n7765) );
  AOI21_X1 U8399 ( .B1(n7759), .B2(n7761), .A(n6649), .ZN(n7757) );
  NAND2_X1 U8400 ( .A1(n7777), .A2(n7778), .ZN(n6814) );
  NAND2_X1 U8401 ( .A1(n8034), .A2(SI_13_), .ZN(n7778) );
  INV_X1 U8402 ( .A(n8010), .ZN(n7066) );
  INV_X1 U8403 ( .A(n7221), .ZN(n14647) );
  OAI21_X1 U8404 ( .B1(n14691), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n7028), .ZN(
        n7221) );
  AND2_X1 U8405 ( .A1(n12641), .A2(n13090), .ZN(n12642) );
  INV_X1 U8406 ( .A(n15431), .ZN(n7412) );
  INV_X1 U8407 ( .A(n12622), .ZN(n7422) );
  AOI21_X1 U8408 ( .B1(n7148), .B2(n6616), .A(n9401), .ZN(n9376) );
  OR2_X1 U8409 ( .A1(n9371), .A2(n10405), .ZN(n7022) );
  NAND2_X1 U8410 ( .A1(n7188), .A2(n6841), .ZN(n10767) );
  NAND2_X1 U8411 ( .A1(n10764), .A2(n10766), .ZN(n6841) );
  OR2_X1 U8412 ( .A1(n10764), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7188) );
  OR2_X1 U8413 ( .A1(n11907), .A2(n11906), .ZN(n6833) );
  OR2_X1 U8414 ( .A1(n11916), .A2(n11861), .ZN(n6960) );
  OR2_X1 U8415 ( .A1(n9064), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9078) );
  NOR2_X1 U8416 ( .A1(n7889), .A2(n6928), .ZN(n6927) );
  INV_X1 U8417 ( .A(n9357), .ZN(n6925) );
  INV_X1 U8418 ( .A(n7888), .ZN(n7887) );
  OAI21_X1 U8419 ( .B1(n7889), .B2(n6587), .A(n9368), .ZN(n7888) );
  OR2_X1 U8420 ( .A1(n9035), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9049) );
  NAND2_X1 U8421 ( .A1(n13140), .A2(n7546), .ZN(n7543) );
  OAI21_X1 U8422 ( .B1(n13182), .B2(n6789), .A(n6787), .ZN(n13152) );
  AOI21_X1 U8423 ( .B1(n6790), .B2(n6788), .A(n6711), .ZN(n6787) );
  INV_X1 U8424 ( .A(n6790), .ZN(n6789) );
  INV_X1 U8425 ( .A(n9142), .ZN(n6788) );
  AND2_X1 U8426 ( .A1(n9347), .A2(n9346), .ZN(n9383) );
  INV_X1 U8427 ( .A(n9313), .ZN(n6918) );
  NAND2_X1 U8428 ( .A1(n12361), .A2(n9392), .ZN(n9131) );
  AND2_X1 U8429 ( .A1(n7527), .A2(n6797), .ZN(n6796) );
  OR2_X1 U8430 ( .A1(n15295), .A2(n6585), .ZN(n6797) );
  INV_X1 U8431 ( .A(n7528), .ZN(n7527) );
  OAI21_X1 U8432 ( .B1(n15283), .B2(n7529), .A(n14814), .ZN(n7528) );
  INV_X1 U8433 ( .A(n9128), .ZN(n7529) );
  NAND2_X1 U8434 ( .A1(n6796), .A2(n6585), .ZN(n6794) );
  AND2_X1 U8435 ( .A1(n9288), .A2(n9286), .ZN(n6921) );
  AND2_X1 U8436 ( .A1(n7869), .A2(n6680), .ZN(n6919) );
  INV_X1 U8437 ( .A(n7870), .ZN(n7869) );
  OAI21_X1 U8438 ( .B1(n15315), .B2(n7871), .A(n9296), .ZN(n7870) );
  INV_X1 U8439 ( .A(n9293), .ZN(n7871) );
  INV_X1 U8440 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8715) );
  NAND2_X1 U8441 ( .A1(n15339), .A2(n9387), .ZN(n9119) );
  NAND2_X1 U8442 ( .A1(n15423), .A2(n15348), .ZN(n9254) );
  NAND2_X1 U8443 ( .A1(n6805), .A2(n6804), .ZN(n9253) );
  NAND2_X1 U8444 ( .A1(n9254), .A2(n9253), .ZN(n9387) );
  NAND2_X1 U8445 ( .A1(n15359), .A2(n11365), .ZN(n9116) );
  NAND2_X1 U8446 ( .A1(n6929), .A2(n9357), .ZN(n13128) );
  NOR2_X1 U8447 ( .A1(n8929), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n8963) );
  NAND2_X1 U8448 ( .A1(n8643), .A2(n8642), .ZN(n8929) );
  AND2_X1 U8449 ( .A1(n6994), .A2(n6688), .ZN(n6992) );
  INV_X1 U8450 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n8778) );
  INV_X1 U8451 ( .A(n8709), .ZN(n7374) );
  CLKBUF_X3 U8452 ( .A(n6552), .Z(n9632) );
  INV_X1 U8453 ( .A(n9785), .ZN(n7594) );
  INV_X1 U8454 ( .A(n6983), .ZN(n6982) );
  OAI21_X1 U8455 ( .B1(n13653), .B2(n7781), .A(n7299), .ZN(n6983) );
  NAND2_X1 U8456 ( .A1(n13644), .A2(n13513), .ZN(n7299) );
  AND2_X1 U8457 ( .A1(n13893), .A2(n13468), .ZN(n7315) );
  AOI21_X1 U8458 ( .B1(n6602), .B2(n7305), .A(n7304), .ZN(n7303) );
  INV_X1 U8459 ( .A(n9718), .ZN(n7305) );
  NOR2_X1 U8460 ( .A1(n13829), .A2(n13796), .ZN(n7304) );
  NOR2_X1 U8461 ( .A1(n7308), .A2(n9718), .ZN(n7307) );
  INV_X1 U8462 ( .A(n12449), .ZN(n7308) );
  OR3_X1 U8463 ( .A1(n8377), .A2(n8375), .A3(n8376), .ZN(n8394) );
  NAND2_X1 U8464 ( .A1(n11849), .A2(n7493), .ZN(n12098) );
  INV_X1 U8465 ( .A(n7921), .ZN(n7610) );
  XNOR2_X1 U8466 ( .A(n8588), .B(n8587), .ZN(n10416) );
  INV_X1 U8467 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7622) );
  OR2_X1 U8468 ( .A1(n8407), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n8408) );
  OR2_X1 U8469 ( .A1(n8254), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8271) );
  NOR2_X1 U8470 ( .A1(n12319), .A2(n7848), .ZN(n7847) );
  NAND2_X1 U8471 ( .A1(n14297), .A2(n7335), .ZN(n7334) );
  NAND2_X1 U8472 ( .A1(n6876), .A2(n7444), .ZN(n7443) );
  INV_X1 U8473 ( .A(n14291), .ZN(n6876) );
  NAND2_X1 U8474 ( .A1(n10307), .A2(n7446), .ZN(n7445) );
  NOR2_X1 U8475 ( .A1(n14329), .A2(n7696), .ZN(n7358) );
  NAND2_X1 U8476 ( .A1(n7360), .A2(n7698), .ZN(n7359) );
  NAND2_X1 U8477 ( .A1(n7456), .A2(n6852), .ZN(n6851) );
  INV_X1 U8478 ( .A(n12577), .ZN(n6852) );
  NOR2_X1 U8479 ( .A1(n7339), .A2(n14574), .ZN(n7338) );
  INV_X1 U8480 ( .A(n7340), .ZN(n7339) );
  NOR2_X1 U8481 ( .A1(n14580), .A2(n14585), .ZN(n7340) );
  NAND2_X1 U8482 ( .A1(n11309), .A2(n11308), .ZN(n11326) );
  NAND2_X1 U8483 ( .A1(n11143), .A2(n11144), .ZN(n11106) );
  NAND2_X1 U8484 ( .A1(n14517), .A2(n14266), .ZN(n7453) );
  INV_X1 U8485 ( .A(n14952), .ZN(n7330) );
  XNOR2_X1 U8486 ( .A(n9589), .B(n9583), .ZN(n8551) );
  NAND2_X1 U8487 ( .A1(n8052), .A2(SI_21_), .ZN(n8054) );
  OR2_X1 U8488 ( .A1(n10028), .A2(n10027), .ZN(n10045) );
  NAND2_X1 U8489 ( .A1(n7348), .A2(n8027), .ZN(n7346) );
  NOR2_X1 U8490 ( .A1(n7347), .A2(n7345), .ZN(n7344) );
  AND2_X1 U8491 ( .A1(n8305), .A2(n8032), .ZN(n8290) );
  NAND2_X1 U8492 ( .A1(n8253), .A2(n8026), .ZN(n7349) );
  XNOR2_X1 U8493 ( .A(n8005), .B(SI_3_), .ZN(n8146) );
  AOI21_X1 U8494 ( .B1(n8109), .B2(n8108), .A(n8000), .ZN(n8132) );
  INV_X1 U8495 ( .A(SI_2_), .ZN(n7741) );
  NOR2_X1 U8496 ( .A1(n14654), .A2(n7126), .ZN(n14681) );
  AND2_X1 U8497 ( .A1(n15566), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n7126) );
  NOR2_X1 U8498 ( .A1(n12642), .A2(n6564), .ZN(n7408) );
  OR2_X1 U8499 ( .A1(n12796), .A2(n12642), .ZN(n7409) );
  NAND2_X1 U8500 ( .A1(n7199), .A2(n7198), .ZN(n7209) );
  INV_X1 U8501 ( .A(n7176), .ZN(n15433) );
  AND2_X1 U8502 ( .A1(n7423), .A2(n7103), .ZN(n7102) );
  INV_X1 U8503 ( .A(n12331), .ZN(n7103) );
  AND2_X1 U8504 ( .A1(n12827), .A2(n7418), .ZN(n7417) );
  OR2_X1 U8505 ( .A1(n12854), .A2(n7419), .ZN(n7418) );
  INV_X1 U8506 ( .A(n12635), .ZN(n7419) );
  INV_X1 U8507 ( .A(n12870), .ZN(n15422) );
  NOR2_X1 U8508 ( .A1(n9402), .A2(n9401), .ZN(n7392) );
  NOR2_X1 U8509 ( .A1(n7394), .A2(n9247), .ZN(n7393) );
  NAND2_X1 U8510 ( .A1(n6616), .A2(n7395), .ZN(n7394) );
  AND2_X1 U8511 ( .A1(n8672), .A2(n8673), .ZN(n7075) );
  AND2_X1 U8512 ( .A1(n8671), .A2(n8670), .ZN(n7074) );
  AOI21_X1 U8513 ( .B1(n7682), .B2(P3_REG2_REG_1__SCAN_IN), .A(n6658), .ZN(
        n10741) );
  NAND2_X1 U8514 ( .A1(n10767), .A2(n10777), .ZN(n11099) );
  NOR2_X1 U8515 ( .A1(n11089), .A2(n10896), .ZN(n10898) );
  OR2_X1 U8516 ( .A1(n11092), .A2(n10876), .ZN(n6775) );
  OAI21_X1 U8517 ( .B1(n11097), .B2(n10884), .A(n7950), .ZN(n10917) );
  AND2_X1 U8518 ( .A1(n10908), .A2(n10907), .ZN(n11057) );
  OR2_X1 U8519 ( .A1(n11204), .A2(n11203), .ZN(n11205) );
  OAI21_X1 U8520 ( .B1(n11067), .B2(n11066), .A(n7942), .ZN(n11226) );
  NAND2_X1 U8521 ( .A1(n7197), .A2(n11550), .ZN(n7684) );
  INV_X1 U8522 ( .A(n7482), .ZN(n11868) );
  NAND2_X1 U8523 ( .A1(n11859), .A2(n11860), .ZN(n6834) );
  INV_X1 U8524 ( .A(n7237), .ZN(n11899) );
  NOR2_X1 U8525 ( .A1(n11905), .A2(n11904), .ZN(n11907) );
  INV_X1 U8526 ( .A(n6833), .ZN(n12349) );
  XNOR2_X1 U8527 ( .A(n7206), .B(n14760), .ZN(n12354) );
  INV_X1 U8528 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15455) );
  OR2_X1 U8529 ( .A1(n12911), .A2(n8863), .ZN(n7240) );
  NAND2_X1 U8530 ( .A1(n12923), .A2(n6839), .ZN(n12926) );
  NAND2_X1 U8531 ( .A1(n6840), .A2(n12929), .ZN(n6839) );
  INV_X1 U8532 ( .A(n12925), .ZN(n6840) );
  NAND2_X1 U8533 ( .A1(n7677), .A2(n12971), .ZN(n7676) );
  NAND2_X1 U8534 ( .A1(n6758), .A2(n6757), .ZN(n12990) );
  NAND2_X1 U8535 ( .A1(n12979), .A2(n6762), .ZN(n6757) );
  NAND2_X1 U8536 ( .A1(n6760), .A2(n6764), .ZN(n6758) );
  AND2_X1 U8537 ( .A1(n12970), .A2(n12971), .ZN(n7187) );
  AND2_X1 U8538 ( .A1(n12954), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7477) );
  INV_X1 U8539 ( .A(n13001), .ZN(n6836) );
  INV_X1 U8540 ( .A(n6837), .ZN(n13000) );
  NOR2_X1 U8541 ( .A1(n7235), .A2(n7234), .ZN(n7233) );
  INV_X1 U8542 ( .A(n12996), .ZN(n7234) );
  NOR2_X1 U8543 ( .A1(n13012), .A2(n14730), .ZN(n7235) );
  NAND2_X1 U8544 ( .A1(n12993), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n13017) );
  INV_X1 U8545 ( .A(n13015), .ZN(n7670) );
  INV_X1 U8546 ( .A(n13039), .ZN(n7132) );
  NAND2_X1 U8547 ( .A1(n13041), .A2(n13042), .ZN(n7105) );
  OAI21_X1 U8548 ( .B1(n7670), .B2(n13037), .A(n7673), .ZN(n7665) );
  OAI21_X1 U8549 ( .B1(n9196), .B2(n9195), .A(n9371), .ZN(n10387) );
  AOI21_X1 U8550 ( .B1(n7509), .B2(n7510), .A(n7507), .ZN(n7506) );
  INV_X1 U8551 ( .A(n13070), .ZN(n7507) );
  OAI21_X1 U8552 ( .B1(n13100), .B2(n7510), .A(n7509), .ZN(n13071) );
  NOR2_X1 U8553 ( .A1(n13074), .A2(n15300), .ZN(n6786) );
  NAND2_X1 U8554 ( .A1(n13100), .A2(n7514), .ZN(n7511) );
  XNOR2_X1 U8555 ( .A(n13088), .B(n13092), .ZN(n7193) );
  NOR2_X1 U8556 ( .A1(n13090), .A2(n15300), .ZN(n7191) );
  AND2_X1 U8557 ( .A1(n9242), .A2(n9243), .ZN(n13092) );
  OAI21_X1 U8558 ( .B1(n6929), .B2(n6926), .A(n6923), .ZN(n13091) );
  INV_X1 U8559 ( .A(n6927), .ZN(n6926) );
  AND2_X1 U8560 ( .A1(n7887), .A2(n6924), .ZN(n6923) );
  NAND2_X1 U8561 ( .A1(n6927), .A2(n6925), .ZN(n6924) );
  NAND2_X1 U8562 ( .A1(n7539), .A2(n7537), .ZN(n13102) );
  NAND2_X1 U8563 ( .A1(n7538), .A2(n6611), .ZN(n7537) );
  INV_X1 U8564 ( .A(n7541), .ZN(n7538) );
  NAND2_X1 U8565 ( .A1(n13102), .A2(n13101), .ZN(n13100) );
  NAND2_X1 U8566 ( .A1(n13116), .A2(n9252), .ZN(n13099) );
  NAND2_X1 U8567 ( .A1(n7543), .A2(n7544), .ZN(n13114) );
  NAND2_X1 U8568 ( .A1(n13130), .A2(n6587), .ZN(n13116) );
  NAND2_X1 U8569 ( .A1(n9010), .A2(n9009), .ZN(n9020) );
  AND2_X1 U8570 ( .A1(n9357), .A2(n9358), .ZN(n13144) );
  AOI21_X1 U8571 ( .B1(n7894), .B2(n8976), .A(n7893), .ZN(n7892) );
  OR2_X1 U8572 ( .A1(n13182), .A2(n9383), .ZN(n13183) );
  INV_X1 U8573 ( .A(n9383), .ZN(n13184) );
  NAND2_X1 U8574 ( .A1(n8934), .A2(n8933), .ZN(n8951) );
  INV_X1 U8575 ( .A(n8935), .ZN(n8934) );
  INV_X1 U8576 ( .A(n13186), .ZN(n13218) );
  OR2_X1 U8577 ( .A1(n8916), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8935) );
  AOI21_X1 U8578 ( .B1(n7876), .B2(n7880), .A(n7874), .ZN(n7873) );
  NAND2_X1 U8579 ( .A1(n6914), .A2(n6566), .ZN(n7872) );
  INV_X1 U8580 ( .A(n9329), .ZN(n7874) );
  NAND2_X1 U8581 ( .A1(n8895), .A2(n8894), .ZN(n8916) );
  INV_X1 U8582 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n8894) );
  INV_X1 U8583 ( .A(n8896), .ZN(n8895) );
  INV_X1 U8584 ( .A(n12898), .ZN(n13245) );
  NAND2_X1 U8585 ( .A1(n9131), .A2(n7535), .ZN(n7534) );
  INV_X1 U8586 ( .A(n8842), .ZN(n8841) );
  NAND2_X1 U8587 ( .A1(n14817), .A2(n9300), .ZN(n12368) );
  INV_X1 U8588 ( .A(n6792), .ZN(n12361) );
  AOI21_X1 U8589 ( .B1(n15294), .B2(n6796), .A(n6793), .ZN(n6792) );
  NAND2_X1 U8590 ( .A1(n6794), .A2(n7525), .ZN(n6793) );
  AOI21_X1 U8591 ( .B1(n7527), .B2(n7529), .A(n6701), .ZN(n7525) );
  NAND2_X1 U8592 ( .A1(n15284), .A2(n15283), .ZN(n7526) );
  INV_X1 U8593 ( .A(n6795), .ZN(n15284) );
  AOI21_X1 U8594 ( .B1(n15294), .B2(n15295), .A(n6585), .ZN(n6795) );
  NAND2_X1 U8595 ( .A1(n8783), .A2(n8782), .ZN(n8801) );
  INV_X1 U8596 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n11556) );
  NAND2_X1 U8597 ( .A1(n15327), .A2(n9124), .ZN(n15309) );
  NOR2_X1 U8598 ( .A1(n8751), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8764) );
  NAND2_X1 U8599 ( .A1(n11705), .A2(n9286), .ZN(n15322) );
  NAND2_X1 U8600 ( .A1(n15322), .A2(n15321), .ZN(n15320) );
  NAND2_X1 U8601 ( .A1(n11694), .A2(n6798), .ZN(n11708) );
  AND2_X1 U8602 ( .A1(n11709), .A2(n9122), .ZN(n6798) );
  OR2_X1 U8603 ( .A1(n8736), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8751) );
  AOI21_X1 U8604 ( .B1(n11697), .B2(n8735), .A(n8734), .ZN(n9278) );
  NAND2_X1 U8605 ( .A1(n7863), .A2(n11697), .ZN(n11692) );
  NOR2_X1 U8606 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8716) );
  NAND2_X1 U8607 ( .A1(n9119), .A2(n9118), .ZN(n11993) );
  AND2_X1 U8608 ( .A1(n9264), .A2(n9263), .ZN(n11992) );
  INV_X1 U8609 ( .A(n9387), .ZN(n15341) );
  INV_X1 U8610 ( .A(n15300), .ZN(n15358) );
  OAI211_X1 U8611 ( .C1(n13377), .C2(n11360), .A(n11359), .B(n11358), .ZN(
        n11363) );
  NOR2_X1 U8612 ( .A1(n13053), .A2(n13052), .ZN(n13319) );
  NAND2_X1 U8613 ( .A1(n15314), .A2(n9293), .ZN(n15303) );
  AND2_X1 U8614 ( .A1(n10934), .A2(n9166), .ZN(n10950) );
  AND2_X1 U8615 ( .A1(n7898), .A2(n8646), .ZN(n6932) );
  NOR2_X1 U8616 ( .A1(n7900), .A2(n7899), .ZN(n7898) );
  NAND2_X1 U8617 ( .A1(n8661), .A2(n9152), .ZN(n7899) );
  OAI21_X1 U8618 ( .B1(n9198), .B2(n9197), .A(n9199), .ZN(n9211) );
  AND2_X1 U8619 ( .A1(n7429), .A2(n7428), .ZN(n7427) );
  INV_X1 U8620 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7428) );
  OAI21_X1 U8621 ( .B1(n9073), .B2(n9072), .A(n9074), .ZN(n9191) );
  XNOR2_X1 U8622 ( .A(n9148), .B(P3_IR_REG_26__SCAN_IN), .ZN(n9162) );
  OR2_X1 U8623 ( .A1(n9031), .A2(n13966), .ZN(n7396) );
  OAI21_X1 U8624 ( .B1(n9016), .B2(n9015), .A(n9017), .ZN(n9028) );
  NAND2_X1 U8625 ( .A1(n9165), .A2(n9164), .ZN(n10933) );
  AND2_X1 U8626 ( .A1(n8977), .A2(n8959), .ZN(n8960) );
  AND2_X1 U8627 ( .A1(n8957), .A2(n8943), .ZN(n8944) );
  NAND2_X1 U8628 ( .A1(n8852), .A2(n10065), .ZN(n8872) );
  NAND2_X1 U8629 ( .A1(n7167), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n7009) );
  OAI21_X1 U8630 ( .B1(n8760), .B2(n8759), .A(n8761), .ZN(n8777) );
  AND2_X1 U8631 ( .A1(n10499), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8759) );
  NAND2_X1 U8632 ( .A1(n6989), .A2(n8725), .ZN(n8744) );
  XNOR2_X1 U8633 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8743) );
  AND2_X1 U8634 ( .A1(n8680), .A2(n8707), .ZN(n8708) );
  XNOR2_X1 U8635 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8709) );
  INV_X1 U8636 ( .A(n8694), .ZN(n7375) );
  NAND2_X1 U8637 ( .A1(n8531), .A2(n7632), .ZN(n7631) );
  INV_X1 U8638 ( .A(n8533), .ZN(n7632) );
  AND2_X1 U8639 ( .A1(n6670), .A2(n7015), .ZN(n7014) );
  NAND2_X1 U8640 ( .A1(n13430), .A2(n8530), .ZN(n7015) );
  NAND2_X1 U8641 ( .A1(n7624), .A2(n7625), .ZN(n7145) );
  NAND2_X1 U8642 ( .A1(n7628), .A2(n6677), .ZN(n7624) );
  NAND2_X1 U8643 ( .A1(n8550), .A2(n7630), .ZN(n7625) );
  AND2_X1 U8644 ( .A1(n13430), .A2(n13456), .ZN(n7010) );
  INV_X1 U8645 ( .A(n8507), .ZN(n8521) );
  NAND2_X1 U8646 ( .A1(n7648), .A2(n7644), .ZN(n7647) );
  INV_X1 U8647 ( .A(n7642), .ZN(n7640) );
  XNOR2_X1 U8648 ( .A(n15227), .B(n6558), .ZN(n11616) );
  NAND2_X1 U8649 ( .A1(n7141), .A2(n11398), .ZN(n11399) );
  AND2_X1 U8650 ( .A1(n11406), .A2(n8172), .ZN(n7141) );
  NAND2_X1 U8651 ( .A1(n8234), .A2(n11516), .ZN(n11444) );
  NAND2_X1 U8652 ( .A1(n8335), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8377) );
  AND2_X1 U8653 ( .A1(n11794), .A2(n8300), .ZN(n7621) );
  XNOR2_X1 U8654 ( .A(n8415), .B(n11781), .ZN(n8141) );
  NAND2_X1 U8655 ( .A1(n7013), .A2(n13430), .ZN(n13484) );
  OR2_X1 U8656 ( .A1(n13453), .A2(n8530), .ZN(n7013) );
  XNOR2_X1 U8657 ( .A(n13829), .B(n6558), .ZN(n8385) );
  AND2_X1 U8658 ( .A1(n7112), .A2(n13628), .ZN(n7111) );
  AND4_X1 U8659 ( .A1(n8513), .A2(n8512), .A3(n8511), .A4(n8510), .ZN(n13426)
         );
  INV_X1 U8660 ( .A(n8139), .ZN(n9601) );
  NOR2_X1 U8661 ( .A1(n6744), .A2(n6743), .ZN(n10854) );
  NOR2_X1 U8662 ( .A1(n10578), .A2(n11766), .ZN(n6743) );
  NAND2_X1 U8663 ( .A1(n10679), .A2(n10678), .ZN(n10813) );
  NAND2_X1 U8664 ( .A1(n15147), .A2(n15146), .ZN(n15145) );
  NAND2_X1 U8665 ( .A1(n15145), .A2(n6749), .ZN(n13553) );
  OR2_X1 U8666 ( .A1(n15148), .A2(n13551), .ZN(n6749) );
  AND2_X1 U8667 ( .A1(n13849), .A2(n9730), .ZN(n7297) );
  INV_X1 U8668 ( .A(n7755), .ZN(n13625) );
  NAND2_X1 U8669 ( .A1(n13678), .A2(n9779), .ZN(n13651) );
  NAND2_X1 U8670 ( .A1(n6881), .A2(n9777), .ZN(n6880) );
  INV_X1 U8671 ( .A(n6885), .ZN(n6881) );
  NAND2_X1 U8672 ( .A1(n7784), .A2(n13669), .ZN(n7783) );
  NAND2_X1 U8673 ( .A1(n9725), .A2(n7314), .ZN(n7313) );
  INV_X1 U8674 ( .A(n9723), .ZN(n7314) );
  NAND2_X1 U8675 ( .A1(n13739), .A2(n6629), .ZN(n7312) );
  INV_X1 U8676 ( .A(n7498), .ZN(n13718) );
  NOR2_X1 U8677 ( .A1(n8441), .A2(n8440), .ZN(n8456) );
  AND2_X1 U8678 ( .A1(n8456), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8458) );
  INV_X1 U8679 ( .A(n13887), .ZN(n7499) );
  OR2_X1 U8680 ( .A1(n8433), .A2(n15652), .ZN(n8441) );
  AND2_X1 U8681 ( .A1(n7301), .A2(n6686), .ZN(n6979) );
  INV_X1 U8682 ( .A(n7604), .ZN(n6912) );
  INV_X1 U8683 ( .A(n7602), .ZN(n7601) );
  OAI21_X1 U8684 ( .B1(n7606), .B2(n7604), .A(n7603), .ZN(n7602) );
  OR2_X1 U8685 ( .A1(n13903), .A2(n13797), .ZN(n7603) );
  NOR2_X1 U8686 ( .A1(n8394), .A2(n8393), .ZN(n8416) );
  NAND2_X1 U8687 ( .A1(n7306), .A2(n7303), .ZN(n13794) );
  NAND2_X1 U8688 ( .A1(n12441), .A2(n7307), .ZN(n7306) );
  NAND2_X1 U8689 ( .A1(n9765), .A2(n9764), .ZN(n13791) );
  INV_X1 U8690 ( .A(n7614), .ZN(n13831) );
  NAND2_X1 U8691 ( .A1(n7496), .A2(n13829), .ZN(n13820) );
  OR2_X1 U8692 ( .A1(n12243), .A2(n9757), .ZN(n9759) );
  NAND2_X1 U8693 ( .A1(n7795), .A2(n6560), .ZN(n7794) );
  NAND2_X1 U8694 ( .A1(n12120), .A2(n7796), .ZN(n6977) );
  INV_X1 U8695 ( .A(n7797), .ZN(n7795) );
  NAND2_X1 U8696 ( .A1(n12119), .A2(n7798), .ZN(n12244) );
  NOR2_X1 U8697 ( .A1(n12102), .A2(n7492), .ZN(n7491) );
  INV_X1 U8698 ( .A(n7493), .ZN(n7492) );
  AOI21_X1 U8699 ( .B1(n6903), .B2(n6905), .A(n6620), .ZN(n6902) );
  NAND2_X1 U8700 ( .A1(n12120), .A2(n12123), .ZN(n12119) );
  OR2_X1 U8701 ( .A1(n8260), .A2(n7977), .ZN(n8279) );
  OAI21_X1 U8702 ( .B1(n11844), .B2(n6987), .A(n7800), .ZN(n12079) );
  INV_X1 U8703 ( .A(n7802), .ZN(n6987) );
  AOI21_X1 U8704 ( .B1(n7802), .B2(n7801), .A(n6647), .ZN(n7800) );
  INV_X1 U8705 ( .A(n9714), .ZN(n7801) );
  NAND2_X1 U8706 ( .A1(n11849), .A2(n11807), .ZN(n12084) );
  AND2_X1 U8707 ( .A1(n11848), .A2(n11852), .ZN(n11849) );
  NOR2_X1 U8708 ( .A1(n11834), .A2(n11815), .ZN(n11848) );
  INV_X1 U8709 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8201) );
  NAND2_X1 U8710 ( .A1(n11826), .A2(n9712), .ZN(n11293) );
  NAND2_X1 U8711 ( .A1(n9747), .A2(n9746), .ZN(n11291) );
  AND2_X1 U8712 ( .A1(n9713), .A2(n9673), .ZN(n11294) );
  OAI21_X1 U8713 ( .B1(n11762), .B2(n6974), .A(n6972), .ZN(n11826) );
  INV_X1 U8714 ( .A(n6973), .ZN(n6972) );
  OAI21_X1 U8715 ( .B1(n11763), .B2(n6974), .A(n11827), .ZN(n6973) );
  INV_X1 U8716 ( .A(n9710), .ZN(n6974) );
  NAND2_X1 U8717 ( .A1(n11761), .A2(n9710), .ZN(n11828) );
  OR2_X1 U8718 ( .A1(n11836), .A2(n11837), .ZN(n11834) );
  AND2_X1 U8719 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8185) );
  NAND2_X1 U8720 ( .A1(n6879), .A2(n9742), .ZN(n11760) );
  NAND2_X1 U8721 ( .A1(n11767), .A2(n11771), .ZN(n11836) );
  NAND2_X1 U8722 ( .A1(n11762), .A2(n11763), .ZN(n11761) );
  AND2_X1 U8723 ( .A1(n9709), .A2(n9677), .ZN(n11191) );
  NAND2_X1 U8724 ( .A1(n7272), .A2(n15222), .ZN(n9737) );
  XNOR2_X1 U8725 ( .A(n7609), .B(n6553), .ZN(n9705) );
  OAI211_X1 U8726 ( .C1(n7592), .C2(n6896), .A(n6895), .B(n6603), .ZN(n12607)
         );
  NAND2_X1 U8727 ( .A1(n6894), .A2(n9788), .ZN(n6893) );
  NAND2_X1 U8728 ( .A1(n9784), .A2(n9783), .ZN(n13627) );
  INV_X1 U8729 ( .A(n12043), .ZN(n11194) );
  INV_X1 U8730 ( .A(n15251), .ZN(n15263) );
  OR2_X1 U8731 ( .A1(n9790), .A2(n9789), .ZN(n15255) );
  AOI21_X1 U8732 ( .B1(n11951), .B2(n15217), .A(n7269), .ZN(n15214) );
  NAND2_X1 U8733 ( .A1(n7967), .A2(n7922), .ZN(n7921) );
  NAND2_X1 U8734 ( .A1(n7972), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6913) );
  NAND2_X1 U8735 ( .A1(n8071), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7969) );
  NAND2_X1 U8736 ( .A1(n8574), .A2(n8572), .ZN(n8579) );
  INV_X1 U8737 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8572) );
  OR2_X1 U8738 ( .A1(n8311), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n8351) );
  OR2_X1 U8739 ( .A1(n8238), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8254) );
  INV_X1 U8740 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8217) );
  INV_X1 U8741 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U8742 ( .A1(n7856), .A2(n6736), .ZN(n7855) );
  INV_X1 U8743 ( .A(n10177), .ZN(n10197) );
  NAND2_X1 U8744 ( .A1(n10197), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n10196) );
  AND2_X1 U8745 ( .A1(n13990), .A2(n13988), .ZN(n12708) );
  NOR2_X1 U8746 ( .A1(n10038), .A2(n10037), .ZN(n10058) );
  NOR2_X1 U8747 ( .A1(n14083), .A2(n7828), .ZN(n6933) );
  OR2_X1 U8748 ( .A1(n14016), .A2(n14084), .ZN(n7828) );
  INV_X1 U8749 ( .A(n10196), .ZN(n10211) );
  NAND2_X1 U8750 ( .A1(n10211), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n10210) );
  INV_X4 U8751 ( .A(n11135), .ZN(n12753) );
  OR2_X1 U8752 ( .A1(n12779), .A2(n11136), .ZN(n11139) );
  OR2_X1 U8753 ( .A1(n10155), .A2(n14043), .ZN(n10166) );
  NAND2_X1 U8754 ( .A1(n12488), .A2(n12489), .ZN(n7849) );
  INV_X1 U8755 ( .A(n7847), .ZN(n7841) );
  INV_X1 U8756 ( .A(n7849), .ZN(n7840) );
  OR2_X1 U8757 ( .A1(n12319), .A2(n7850), .ZN(n7846) );
  NAND2_X1 U8758 ( .A1(n14876), .A2(n7847), .ZN(n7845) );
  NAND2_X1 U8759 ( .A1(n6939), .A2(n11645), .ZN(n11667) );
  OR2_X1 U8760 ( .A1(n11647), .A2(n11646), .ZN(n6939) );
  AOI21_X1 U8761 ( .B1(n6951), .B2(n6949), .A(n6948), .ZN(n6947) );
  INV_X1 U8762 ( .A(n6951), .ZN(n6950) );
  INV_X1 U8763 ( .A(n14073), .ZN(n6948) );
  OR2_X1 U8764 ( .A1(n14083), .A2(n14084), .ZN(n7830) );
  AND3_X1 U8765 ( .A1(n10082), .A2(n10081), .A3(n10080), .ZN(n12670) );
  INV_X1 U8766 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n15651) );
  NAND2_X1 U8767 ( .A1(n10300), .A2(n10299), .ZN(n10344) );
  NAND2_X1 U8768 ( .A1(n10267), .A2(n10266), .ZN(n14249) );
  NAND2_X1 U8769 ( .A1(n10274), .A2(n10273), .ZN(n14261) );
  NAND2_X1 U8770 ( .A1(n7439), .A2(n7440), .ZN(n12598) );
  AOI21_X1 U8771 ( .B1(n7441), .B2(n14300), .A(n6635), .ZN(n7440) );
  NAND2_X1 U8772 ( .A1(n14291), .A2(n7441), .ZN(n7439) );
  NOR2_X1 U8773 ( .A1(n14332), .A2(n7334), .ZN(n14293) );
  AND2_X1 U8774 ( .A1(n14298), .A2(n12565), .ZN(n14278) );
  NAND2_X1 U8775 ( .A1(n14273), .A2(n6874), .ZN(n14287) );
  NAND2_X1 U8776 ( .A1(n7443), .A2(n7441), .ZN(n14273) );
  NAND2_X1 U8777 ( .A1(n6875), .A2(n12594), .ZN(n6874) );
  NAND2_X1 U8778 ( .A1(n7443), .A2(n7445), .ZN(n6875) );
  NOR2_X1 U8779 ( .A1(n14332), .A2(n14535), .ZN(n14314) );
  AND2_X1 U8780 ( .A1(n14323), .A2(n12591), .ZN(n7945) );
  NAND2_X1 U8781 ( .A1(n14324), .A2(n14329), .ZN(n14323) );
  AND2_X1 U8782 ( .A1(n7359), .A2(n7358), .ZN(n14327) );
  NAND2_X1 U8783 ( .A1(n7359), .A2(n7702), .ZN(n14328) );
  INV_X1 U8784 ( .A(n7473), .ZN(n7472) );
  NAND2_X1 U8785 ( .A1(n14388), .A2(n7474), .ZN(n6873) );
  OAI22_X1 U8786 ( .A1(n14362), .A2(n12588), .B1(n14095), .B2(n14551), .ZN(
        n7473) );
  NAND2_X1 U8787 ( .A1(n14467), .A2(n7336), .ZN(n14395) );
  NOR2_X1 U8788 ( .A1(n14566), .A2(n7337), .ZN(n7336) );
  INV_X1 U8789 ( .A(n7338), .ZN(n7337) );
  NAND2_X1 U8790 ( .A1(n14467), .A2(n7340), .ZN(n14429) );
  NAND2_X1 U8791 ( .A1(n7458), .A2(n12579), .ZN(n14421) );
  OR2_X1 U8792 ( .A1(n14438), .A2(n12578), .ZN(n7458) );
  NAND2_X1 U8793 ( .A1(n14467), .A2(n14444), .ZN(n14439) );
  NOR2_X1 U8794 ( .A1(n10088), .A2(n10087), .ZN(n10094) );
  AND2_X1 U8795 ( .A1(n10094), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10115) );
  INV_X1 U8796 ( .A(n7464), .ZN(n7463) );
  OR2_X1 U8797 ( .A1(n10076), .A2(n10075), .ZN(n10088) );
  NAND2_X1 U8798 ( .A1(n7711), .A2(n7713), .ZN(n12258) );
  INV_X1 U8799 ( .A(n7718), .ZN(n7717) );
  AOI21_X1 U8800 ( .B1(n7468), .B2(n7467), .A(n6644), .ZN(n7466) );
  OR2_X1 U8801 ( .A1(n10019), .A2(n15586), .ZN(n10038) );
  NOR2_X1 U8802 ( .A1(n9990), .A2(n10794), .ZN(n10008) );
  OR2_X1 U8803 ( .A1(n9965), .A2(n11678), .ZN(n9978) );
  OR2_X1 U8804 ( .A1(n9978), .A2(n9977), .ZN(n9990) );
  OAI21_X1 U8805 ( .B1(n6847), .B2(n11591), .A(n6846), .ZN(n14983) );
  AOI21_X1 U8806 ( .B1(n6845), .B2(n11717), .A(n6843), .ZN(n6846) );
  OAI21_X1 U8807 ( .B1(n11591), .B2(n6844), .A(n6661), .ZN(n6843) );
  INV_X1 U8808 ( .A(n6591), .ZN(n6844) );
  NAND2_X1 U8809 ( .A1(n7709), .A2(n7707), .ZN(n11592) );
  NAND2_X1 U8810 ( .A1(n7708), .A2(n6595), .ZN(n7707) );
  NAND2_X1 U8811 ( .A1(n7706), .A2(n11590), .ZN(n7708) );
  AOI22_X1 U8812 ( .A1(n9886), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n10136), .B2(
        n14148), .ZN(n9869) );
  NOR2_X1 U8813 ( .A1(n11331), .A2(n14933), .ZN(n11330) );
  NAND2_X1 U8814 ( .A1(n11143), .A2(n11463), .ZN(n11117) );
  NAND2_X1 U8815 ( .A1(n7324), .A2(n7321), .ZN(n11331) );
  INV_X1 U8816 ( .A(n11117), .ZN(n7321) );
  NAND2_X1 U8817 ( .A1(n10317), .A2(n11106), .ZN(n10707) );
  INV_X1 U8818 ( .A(n7453), .ZN(n7448) );
  INV_X1 U8819 ( .A(n14254), .ZN(n7169) );
  INV_X1 U8820 ( .A(n14060), .ZN(n14551) );
  NAND2_X1 U8821 ( .A1(n11886), .A2(n11885), .ZN(n11940) );
  NAND2_X1 U8822 ( .A1(n11303), .A2(n11313), .ZN(n14951) );
  AND2_X1 U8823 ( .A1(n9819), .A2(n7737), .ZN(n7736) );
  NAND2_X1 U8824 ( .A1(n9606), .A2(n9594), .ZN(n9609) );
  XNOR2_X1 U8825 ( .A(n9623), .B(n9622), .ZN(n13948) );
  XNOR2_X1 U8826 ( .A(n8551), .B(SI_27_), .ZN(n13954) );
  AND2_X1 U8827 ( .A1(n10368), .A2(n9816), .ZN(n10554) );
  OAI21_X1 U8828 ( .B1(n10366), .B2(n10365), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n10367) );
  NAND2_X1 U8829 ( .A1(n6823), .A2(n8068), .ZN(n8536) );
  NAND2_X1 U8830 ( .A1(n8503), .A2(n8065), .ZN(n8516) );
  NAND2_X1 U8831 ( .A1(n10362), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10363) );
  INV_X1 U8832 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7860) );
  NAND2_X1 U8833 ( .A1(n8087), .A2(n8086), .ZN(n8089) );
  NAND2_X1 U8834 ( .A1(n6807), .A2(n6808), .ZN(n8453) );
  OAI21_X1 U8835 ( .B1(n8428), .B2(n8048), .A(n8049), .ZN(n8446) );
  NAND2_X1 U8836 ( .A1(n7758), .A2(n8043), .ZN(n8406) );
  NAND2_X1 U8837 ( .A1(n8387), .A2(n8386), .ZN(n7758) );
  AND2_X1 U8838 ( .A1(n10014), .A2(n10002), .ZN(n10976) );
  XNOR2_X1 U8839 ( .A(n8216), .B(n8215), .ZN(n10508) );
  NOR2_X1 U8840 ( .A1(n9952), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n9955) );
  OR2_X1 U8841 ( .A1(n9935), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9952) );
  NAND2_X1 U8842 ( .A1(n7067), .A2(n8010), .ZN(n8177) );
  NAND2_X1 U8843 ( .A1(n8008), .A2(n8159), .ZN(n7067) );
  AND2_X1 U8844 ( .A1(n7200), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14684) );
  INV_X1 U8845 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7200) );
  XNOR2_X1 U8846 ( .A(n14684), .B(n7127), .ZN(n14687) );
  XNOR2_X1 U8847 ( .A(n7663), .B(P1_ADDR_REG_1__SCAN_IN), .ZN(n7127) );
  AOI22_X1 U8848 ( .A1(n14684), .A2(n14645), .B1(P3_ADDR_REG_1__SCAN_IN), .B2(
        n15651), .ZN(n14690) );
  NAND2_X1 U8849 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7663), .ZN(n14645) );
  XNOR2_X1 U8850 ( .A(n14696), .B(n7173), .ZN(n14698) );
  NOR2_X1 U8851 ( .A1(n15734), .A2(n14695), .ZN(n14697) );
  NOR2_X1 U8852 ( .A1(n14650), .A2(n14649), .ZN(n14701) );
  INV_X1 U8853 ( .A(n7027), .ZN(n14648) );
  NOR2_X1 U8854 ( .A1(n14660), .A2(n14659), .ZN(n14717) );
  NOR2_X1 U8855 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n14715), .ZN(n14659) );
  AOI22_X1 U8856 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14665), .B1(n14721), 
        .B2(n14664), .ZN(n14676) );
  XNOR2_X1 U8857 ( .A(n15328), .B(n12640), .ZN(n12108) );
  INV_X1 U8858 ( .A(n12505), .ZN(n7089) );
  AND2_X1 U8859 ( .A1(n12508), .A2(n7087), .ZN(n7086) );
  NAND2_X1 U8860 ( .A1(n7088), .A2(n12505), .ZN(n7087) );
  NAND2_X1 U8861 ( .A1(n7085), .A2(n12505), .ZN(n12509) );
  NAND2_X1 U8862 ( .A1(n12427), .A2(n7090), .ZN(n7085) );
  NOR2_X1 U8863 ( .A1(n12181), .A2(n7425), .ZN(n12330) );
  AND2_X1 U8864 ( .A1(n7094), .A2(n7092), .ZN(n7091) );
  INV_X1 U8865 ( .A(n12811), .ZN(n7092) );
  NAND2_X1 U8866 ( .A1(n7093), .A2(n7094), .ZN(n12812) );
  AND2_X1 U8867 ( .A1(n8013), .A2(n7520), .ZN(n7519) );
  NAND2_X1 U8868 ( .A1(n12862), .A2(n12622), .ZN(n12819) );
  AND4_X1 U8869 ( .A1(n8871), .A2(n8870), .A3(n8869), .A4(n8868), .ZN(n12428)
         );
  AND2_X1 U8870 ( .A1(n8839), .A2(n8838), .ZN(n12409) );
  NAND2_X1 U8871 ( .A1(n9046), .A2(n9045), .ZN(n12832) );
  OR2_X1 U8872 ( .A1(n8722), .A2(n12344), .ZN(n9045) );
  INV_X1 U8873 ( .A(n13367), .ZN(n12841) );
  INV_X1 U8874 ( .A(n7199), .ZN(n11742) );
  AND2_X1 U8875 ( .A1(n9055), .A2(n9054), .ZN(n13089) );
  NAND2_X1 U8876 ( .A1(n12632), .A2(n12631), .ZN(n12853) );
  NAND2_X1 U8877 ( .A1(n9034), .A2(n9033), .ZN(n12858) );
  OR2_X1 U8878 ( .A1(n8722), .A2(n12207), .ZN(n9033) );
  INV_X1 U8879 ( .A(n7411), .ZN(n11740) );
  NOR2_X1 U8880 ( .A1(n12012), .A2(n12013), .ZN(n12181) );
  NAND2_X1 U8881 ( .A1(n7208), .A2(n12010), .ZN(n12012) );
  NAND2_X1 U8882 ( .A1(n12864), .A2(n12863), .ZN(n12862) );
  NAND2_X1 U8883 ( .A1(n12427), .A2(n12426), .ZN(n12507) );
  NAND2_X1 U8884 ( .A1(n7098), .A2(n12616), .ZN(n12880) );
  NAND2_X1 U8885 ( .A1(n12845), .A2(n12844), .ZN(n7098) );
  NAND2_X1 U8886 ( .A1(n10943), .A2(n10942), .ZN(n15439) );
  NAND2_X1 U8887 ( .A1(n9063), .A2(n9062), .ZN(n13093) );
  OR2_X1 U8888 ( .A1(n8722), .A2(n12455), .ZN(n9062) );
  INV_X1 U8889 ( .A(n12830), .ZN(n13104) );
  NAND2_X1 U8890 ( .A1(n9001), .A2(n9000), .ZN(n13171) );
  INV_X1 U8891 ( .A(n13156), .ZN(n13187) );
  NAND4_X1 U8892 ( .A1(n8690), .A2(n8689), .A3(n8688), .A4(n8687), .ZN(n15343)
         );
  NAND2_X1 U8893 ( .A1(n8702), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8690) );
  OR2_X1 U8894 ( .A1(n8699), .A2(n10757), .ZN(n8655) );
  NAND2_X1 U8895 ( .A1(n8702), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8653) );
  NAND2_X1 U8896 ( .A1(n7074), .A2(n7075), .ZN(n15359) );
  INV_X1 U8897 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14685) );
  INV_X1 U8898 ( .A(n7166), .ZN(n11072) );
  XNOR2_X1 U8899 ( .A(n11057), .B(n7480), .ZN(n10909) );
  NOR2_X1 U8900 ( .A1(n10909), .A2(n10911), .ZN(n11058) );
  INV_X1 U8901 ( .A(n7246), .ZN(n11074) );
  INV_X1 U8902 ( .A(n7242), .ZN(n11558) );
  INV_X1 U8903 ( .A(n7197), .ZN(n11551) );
  XNOR2_X1 U8904 ( .A(n7237), .B(n11873), .ZN(n11856) );
  INV_X1 U8905 ( .A(n7243), .ZN(n11914) );
  NAND2_X1 U8906 ( .A1(n12398), .A2(n12397), .ZN(n6752) );
  INV_X1 U8907 ( .A(n7681), .ZN(n12398) );
  INV_X1 U8908 ( .A(n12383), .ZN(n7485) );
  INV_X1 U8909 ( .A(n7486), .ZN(n12384) );
  INV_X1 U8910 ( .A(n7232), .ZN(n12953) );
  NOR2_X1 U8911 ( .A1(n7673), .A2(n13037), .ZN(n7668) );
  XNOR2_X1 U8912 ( .A(n10387), .B(n6616), .ZN(n13064) );
  NAND2_X1 U8913 ( .A1(n7192), .A2(n7189), .ZN(n13266) );
  NOR2_X1 U8914 ( .A1(n7191), .A2(n7190), .ZN(n7189) );
  NAND2_X1 U8915 ( .A1(n7193), .A2(n10380), .ZN(n7192) );
  NOR2_X1 U8916 ( .A1(n13089), .A2(n15298), .ZN(n7190) );
  AOI21_X1 U8917 ( .B1(n13140), .B2(n9144), .A(n6588), .ZN(n13126) );
  AOI21_X1 U8918 ( .B1(n11685), .B2(n9234), .A(n9007), .ZN(n13147) );
  NAND2_X1 U8919 ( .A1(n7896), .A2(n9347), .ZN(n13174) );
  NAND2_X1 U8920 ( .A1(n7897), .A2(n9346), .ZN(n7896) );
  NAND2_X1 U8921 ( .A1(n9140), .A2(n9139), .ZN(n13201) );
  NAND2_X1 U8922 ( .A1(n13219), .A2(n9334), .ZN(n13196) );
  NAND2_X1 U8923 ( .A1(n7875), .A2(n7879), .ZN(n13247) );
  NAND2_X1 U8924 ( .A1(n12463), .A2(n7882), .ZN(n7875) );
  OAI21_X1 U8925 ( .B1(n12463), .B2(n9314), .A(n9312), .ZN(n12525) );
  NAND2_X1 U8926 ( .A1(n8861), .A2(n8860), .ZN(n14821) );
  NAND2_X1 U8927 ( .A1(n8815), .A2(n9302), .ZN(n14815) );
  NAND2_X1 U8928 ( .A1(n11422), .A2(n9121), .ZN(n11696) );
  NAND2_X1 U8929 ( .A1(n15336), .A2(n13290), .ZN(n13249) );
  NAND2_X1 U8930 ( .A1(n13081), .A2(n11688), .ZN(n15323) );
  OR2_X1 U8931 ( .A1(n11361), .A2(n15368), .ZN(n15326) );
  NAND2_X1 U8932 ( .A1(n9236), .A2(n9235), .ZN(n13322) );
  NAND2_X1 U8933 ( .A1(n12655), .A2(n9234), .ZN(n9236) );
  NOR2_X1 U8934 ( .A1(n13080), .A2(n7938), .ZN(n13329) );
  INV_X1 U8935 ( .A(n12832), .ZN(n13337) );
  INV_X1 U8936 ( .A(n12858), .ZN(n13341) );
  NAND2_X1 U8937 ( .A1(n8967), .A2(n8966), .ZN(n13355) );
  AND2_X1 U8938 ( .A1(n8950), .A2(n8949), .ZN(n13359) );
  AND2_X1 U8939 ( .A1(n8932), .A2(n8931), .ZN(n13363) );
  NAND2_X1 U8940 ( .A1(n8880), .A2(n8879), .ZN(n13375) );
  AND3_X1 U8941 ( .A1(n8750), .A2(n8749), .A3(n8748), .ZN(n12144) );
  OAI211_X1 U8942 ( .C1(n10922), .C2(n10733), .A(n8713), .B(n8712), .ZN(n12137) );
  INV_X1 U8943 ( .A(n11365), .ZN(n11432) );
  NAND2_X1 U8944 ( .A1(n10933), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13378) );
  NAND2_X1 U8945 ( .A1(n9149), .A2(n6931), .ZN(n13385) );
  AND2_X1 U8946 ( .A1(n6932), .A2(n8647), .ZN(n6931) );
  INV_X1 U8947 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8647) );
  INV_X1 U8948 ( .A(n8651), .ZN(n13388) );
  XNOR2_X1 U8949 ( .A(n9153), .B(n9152), .ZN(n12346) );
  NAND2_X1 U8950 ( .A1(n6582), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9153) );
  NAND2_X1 U8951 ( .A1(n9151), .A2(n6582), .ZN(n12209) );
  XNOR2_X1 U8952 ( .A(n9098), .B(n7886), .ZN(n11683) );
  NAND2_X1 U8953 ( .A1(n8989), .A2(n8988), .ZN(n8992) );
  NAND2_X1 U8954 ( .A1(n9096), .A2(n9095), .ZN(n11542) );
  OAI21_X1 U8955 ( .B1(n7223), .B2(n8902), .A(n7380), .ZN(n8908) );
  NAND2_X1 U8956 ( .A1(n7223), .A2(n8887), .ZN(n8904) );
  NAND2_X1 U8957 ( .A1(n6993), .A2(n6994), .ZN(n8832) );
  OR2_X1 U8958 ( .A1(n8797), .A2(n7386), .ZN(n6993) );
  NAND2_X1 U8959 ( .A1(n7384), .A2(n8812), .ZN(n8826) );
  NAND2_X1 U8960 ( .A1(n8811), .A2(n8810), .ZN(n7384) );
  INV_X1 U8961 ( .A(n11210), .ZN(n14747) );
  NOR2_X1 U8962 ( .A1(n8729), .A2(n6969), .ZN(n10922) );
  OAI21_X1 U8963 ( .B1(n8708), .B2(n6971), .A(n6970), .ZN(n6969) );
  NAND2_X1 U8964 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n6971) );
  NAND2_X1 U8965 ( .A1(n8660), .A2(n15706), .ZN(n6970) );
  OR2_X1 U8966 ( .A1(n8680), .A2(n8660), .ZN(n8682) );
  NAND2_X1 U8967 ( .A1(n8683), .A2(n8684), .ZN(n8695) );
  NAND2_X1 U8968 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8669) );
  NAND2_X1 U8969 ( .A1(n8660), .A2(n7689), .ZN(n7687) );
  INV_X1 U8970 ( .A(n8667), .ZN(n8664) );
  NAND2_X1 U8971 ( .A1(n8345), .A2(n8344), .ZN(n14841) );
  NAND2_X1 U8972 ( .A1(n13397), .A2(n7231), .ZN(n13403) );
  AND2_X1 U8973 ( .A1(n13669), .A2(n8285), .ZN(n7231) );
  NAND2_X1 U8974 ( .A1(n11639), .A2(n8269), .ZN(n11930) );
  NAND2_X1 U8975 ( .A1(n8145), .A2(n8144), .ZN(n11526) );
  NAND2_X1 U8976 ( .A1(n7635), .A2(n7634), .ZN(n13406) );
  AND2_X1 U8977 ( .A1(n7635), .A2(n7638), .ZN(n13408) );
  NAND2_X1 U8978 ( .A1(n7001), .A2(n7636), .ZN(n7635) );
  NAND2_X1 U8979 ( .A1(n7626), .A2(n7144), .ZN(n8633) );
  NAND2_X1 U8980 ( .A1(n7012), .A2(n7011), .ZN(n7626) );
  AOI21_X1 U8981 ( .B1(n13483), .B2(n6628), .A(n7145), .ZN(n7144) );
  AND2_X1 U8982 ( .A1(n6677), .A2(n7014), .ZN(n7011) );
  INV_X1 U8983 ( .A(n7620), .ZN(n15111) );
  NAND2_X1 U8984 ( .A1(n7641), .A2(n7642), .ZN(n13437) );
  AOI22_X1 U8985 ( .A1(n8384), .A2(n7647), .B1(n8385), .B2(n13495), .ZN(n13438) );
  AND2_X1 U8986 ( .A1(n7641), .A2(n7639), .ZN(n13448) );
  AOI21_X1 U8987 ( .B1(n7634), .B2(n7637), .A(n8451), .ZN(n7633) );
  INV_X1 U8988 ( .A(n15109), .ZN(n7619) );
  NAND2_X1 U8989 ( .A1(n8334), .A2(n8333), .ZN(n12420) );
  NOR2_X1 U8990 ( .A1(n12539), .A2(n6699), .ZN(n12547) );
  NAND2_X1 U8991 ( .A1(n8125), .A2(n8124), .ZN(n11378) );
  NOR2_X1 U8992 ( .A1(n13446), .A2(n8426), .ZN(n13475) );
  NAND2_X1 U8993 ( .A1(n8432), .A2(n8431), .ZN(n13898) );
  OAI21_X1 U8994 ( .B1(n8618), .B2(n8612), .A(n13784), .ZN(n13506) );
  XNOR2_X1 U8995 ( .A(n8384), .B(n8385), .ZN(n13497) );
  NAND2_X1 U8996 ( .A1(n6811), .A2(n9658), .ZN(n6810) );
  INV_X1 U8997 ( .A(n13426), .ZN(n13685) );
  NOR2_X1 U8998 ( .A1(n6624), .A2(n6986), .ZN(n6985) );
  INV_X1 U8999 ( .A(n7906), .ZN(n8101) );
  OR2_X1 U9000 ( .A1(n8136), .A2(n8098), .ZN(n8100) );
  AND2_X1 U9001 ( .A1(n6750), .A2(n8112), .ZN(n13531) );
  INV_X1 U9002 ( .A(n8111), .ZN(n6750) );
  NOR3_X1 U9003 ( .A1(n15129), .A2(n6744), .A3(n10441), .ZN(n10447) );
  NOR2_X1 U9004 ( .A1(n10816), .A2(n10815), .ZN(n11037) );
  NAND2_X1 U9005 ( .A1(n10813), .A2(n6747), .ZN(n10816) );
  OR2_X1 U9006 ( .A1(n10814), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6747) );
  XNOR2_X1 U9007 ( .A(n13553), .B(n15164), .ZN(n15161) );
  NAND2_X1 U9008 ( .A1(n15170), .A2(n13556), .ZN(n15185) );
  NAND2_X1 U9009 ( .A1(n15185), .A2(n15184), .ZN(n15183) );
  XNOR2_X1 U9010 ( .A(n6745), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n13588) );
  NAND2_X1 U9011 ( .A1(n6746), .A2(n6609), .ZN(n6745) );
  INV_X1 U9012 ( .A(n7613), .ZN(n7317) );
  AOI21_X1 U9013 ( .B1(n12609), .B2(n13835), .A(n12608), .ZN(n7613) );
  NOR2_X1 U9014 ( .A1(n12607), .A2(n13832), .ZN(n7183) );
  NAND2_X1 U9015 ( .A1(n13848), .A2(n9785), .ZN(n13612) );
  NAND2_X1 U9016 ( .A1(n13652), .A2(n7780), .ZN(n13636) );
  AND2_X1 U9017 ( .A1(n8505), .A2(n8504), .ZN(n13677) );
  NAND2_X1 U9018 ( .A1(n6883), .A2(n6885), .ZN(n13687) );
  NAND2_X1 U9019 ( .A1(n6884), .A2(n7596), .ZN(n13688) );
  NAND2_X1 U9020 ( .A1(n13727), .A2(n7596), .ZN(n6883) );
  NAND2_X1 U9021 ( .A1(n7595), .A2(n7599), .ZN(n13704) );
  NAND2_X1 U9022 ( .A1(n13727), .A2(n9776), .ZN(n7595) );
  OR2_X1 U9023 ( .A1(n12210), .A2(n9610), .ZN(n8472) );
  OR2_X1 U9024 ( .A1(n13727), .A2(n13726), .ZN(n13881) );
  NAND2_X1 U9025 ( .A1(n13738), .A2(n9723), .ZN(n13715) );
  NAND2_X1 U9026 ( .A1(n7129), .A2(n7301), .ZN(n13776) );
  NAND2_X1 U9027 ( .A1(n13793), .A2(n9766), .ZN(n13775) );
  AOI21_X1 U9028 ( .B1(n12441), .B2(n12449), .A(n6602), .ZN(n13813) );
  NAND2_X1 U9029 ( .A1(n12076), .A2(n9754), .ZN(n12090) );
  INV_X1 U9030 ( .A(n13828), .ZN(n13734) );
  NAND2_X1 U9031 ( .A1(n7804), .A2(n7802), .ZN(n11607) );
  NAND2_X1 U9032 ( .A1(n7804), .A2(n9715), .ZN(n11605) );
  NAND2_X1 U9033 ( .A1(n15210), .A2(n8611), .ZN(n13784) );
  AOI21_X1 U9034 ( .B1(n13524), .B2(n13816), .A(n7268), .ZN(n11788) );
  AND2_X1 U9035 ( .A1(n8615), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15210) );
  NAND2_X1 U9036 ( .A1(n8076), .A2(n8073), .ZN(n13955) );
  XNOR2_X1 U9037 ( .A(n8580), .B(P2_IR_REG_26__SCAN_IN), .ZN(n13957) );
  OAI21_X1 U9038 ( .B1(n8579), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8580) );
  NAND2_X1 U9039 ( .A1(n7988), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7989) );
  INV_X1 U9040 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n15645) );
  NAND2_X1 U9041 ( .A1(n7986), .A2(n8178), .ZN(n7990) );
  INV_X1 U9042 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8084) );
  INV_X1 U9043 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11236) );
  INV_X1 U9044 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11183) );
  INV_X1 U9045 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n15544) );
  INV_X1 U9046 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10571) );
  INV_X1 U9047 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10499) );
  INV_X1 U9048 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10490) );
  INV_X1 U9049 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10497) );
  INV_X1 U9050 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10493) );
  INV_X1 U9051 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10488) );
  INV_X1 U9052 ( .A(n13531), .ZN(n13532) );
  NAND2_X1 U9053 ( .A1(n11476), .A2(n11475), .ZN(n14937) );
  NAND2_X1 U9054 ( .A1(n14061), .A2(n12708), .ZN(n13989) );
  AOI21_X1 U9055 ( .B1(n7810), .B2(n12767), .A(n12775), .ZN(n7809) );
  AOI21_X1 U9056 ( .B1(n6940), .B2(n6937), .A(n6936), .ZN(n6935) );
  INV_X1 U9057 ( .A(n6944), .ZN(n6937) );
  INV_X1 U9058 ( .A(n14946), .ZN(n6936) );
  NAND2_X1 U9059 ( .A1(n6938), .A2(n6940), .ZN(n14945) );
  NAND2_X1 U9060 ( .A1(n11647), .A2(n6944), .ZN(n6938) );
  NAND2_X1 U9061 ( .A1(n7812), .A2(n7816), .ZN(n13999) );
  OR2_X1 U9062 ( .A1(n14061), .A2(n7818), .ZN(n7812) );
  OAI21_X1 U9063 ( .B1(n13981), .B2(n7836), .A(n7833), .ZN(n14006) );
  NAND2_X1 U9064 ( .A1(n7832), .A2(n7835), .ZN(n14007) );
  NAND2_X1 U9065 ( .A1(n13981), .A2(n7837), .ZN(n7832) );
  AOI21_X1 U9066 ( .B1(n7829), .B2(n14084), .A(n14016), .ZN(n7826) );
  NAND2_X1 U9067 ( .A1(n14083), .A2(n7829), .ZN(n7827) );
  AND2_X1 U9068 ( .A1(n7830), .A2(n12680), .ZN(n14017) );
  NAND2_X1 U9069 ( .A1(n13989), .A2(n7823), .ZN(n14042) );
  NAND2_X1 U9070 ( .A1(n7845), .A2(n7846), .ZN(n12479) );
  AOI21_X1 U9071 ( .B1(n14876), .B2(n14873), .A(n14874), .ZN(n12320) );
  NAND2_X1 U9072 ( .A1(n11149), .A2(n11148), .ZN(n11471) );
  OR2_X1 U9073 ( .A1(n14297), .A2(n14902), .ZN(n14528) );
  NAND2_X1 U9074 ( .A1(n11153), .A2(n11158), .ZN(n14935) );
  NAND2_X1 U9075 ( .A1(n10179), .A2(n9856), .ZN(n9857) );
  NAND2_X1 U9076 ( .A1(n10179), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n7692) );
  NAND2_X1 U9077 ( .A1(n10260), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7691) );
  NAND2_X1 U9078 ( .A1(n6549), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7693) );
  NAND2_X1 U9079 ( .A1(n9893), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9883) );
  NAND2_X1 U9080 ( .A1(n10179), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n9882) );
  NAND2_X1 U9081 ( .A1(n9893), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9894) );
  INV_X1 U9082 ( .A(n10344), .ZN(n14504) );
  INV_X1 U9083 ( .A(n14249), .ZN(n14507) );
  INV_X1 U9084 ( .A(n14260), .ZN(n14241) );
  AOI21_X1 U9085 ( .B1(n12571), .B2(n15052), .A(n12570), .ZN(n14519) );
  NAND2_X1 U9086 ( .A1(n12567), .A2(n14256), .ZN(n12571) );
  NAND2_X1 U9087 ( .A1(n7697), .A2(n7704), .ZN(n14345) );
  OAI21_X1 U9088 ( .B1(n7109), .B2(n7705), .A(n7698), .ZN(n14343) );
  NAND2_X1 U9089 ( .A1(n7109), .A2(n7700), .ZN(n7697) );
  AND2_X1 U9090 ( .A1(n14373), .A2(n12588), .ZN(n14363) );
  AND2_X1 U9091 ( .A1(n14361), .A2(n14360), .ZN(n14556) );
  OR2_X1 U9092 ( .A1(n14357), .A2(n15002), .ZN(n14361) );
  AND2_X1 U9093 ( .A1(n14388), .A2(n12587), .ZN(n14375) );
  NAND2_X1 U9094 ( .A1(n7731), .A2(n12560), .ZN(n14392) );
  NAND2_X1 U9095 ( .A1(n7454), .A2(n7459), .ZN(n14416) );
  NAND2_X1 U9096 ( .A1(n14438), .A2(n7455), .ZN(n7454) );
  INV_X1 U9097 ( .A(n7457), .ZN(n7455) );
  NAND2_X1 U9098 ( .A1(n12559), .A2(n12558), .ZN(n14407) );
  NAND2_X1 U9099 ( .A1(n14456), .A2(n12556), .ZN(n14446) );
  NAND2_X1 U9100 ( .A1(n12576), .A2(n12575), .ZN(n14488) );
  NAND2_X1 U9101 ( .A1(n7470), .A2(n12026), .ZN(n12027) );
  NAND2_X1 U9102 ( .A1(n7471), .A2(n6586), .ZN(n7470) );
  AND2_X1 U9103 ( .A1(n7719), .A2(n6621), .ZN(n12033) );
  NAND2_X1 U9104 ( .A1(n7718), .A2(n7719), .ZN(n14785) );
  AND2_X1 U9105 ( .A1(n7724), .A2(n7723), .ZN(n11888) );
  NAND2_X1 U9106 ( .A1(n10565), .A2(n10237), .ZN(n7047) );
  OR2_X1 U9107 ( .A1(n6550), .A2(n11313), .ZN(n15009) );
  NAND2_X1 U9108 ( .A1(n6847), .A2(n6848), .ZN(n11718) );
  NOR2_X1 U9109 ( .A1(n6845), .A2(n6591), .ZN(n6848) );
  NAND2_X1 U9110 ( .A1(n7710), .A2(n11589), .ZN(n15000) );
  OR2_X1 U9111 ( .A1(n11586), .A2(n11585), .ZN(n7710) );
  INV_X1 U9112 ( .A(n7432), .ZN(n14999) );
  AOI21_X1 U9113 ( .B1(n11584), .B2(n7433), .A(n7434), .ZN(n7432) );
  INV_X1 U9114 ( .A(n7436), .ZN(n7433) );
  OR2_X1 U9115 ( .A1(n6550), .A2(n11307), .ZN(n14490) );
  OR2_X1 U9116 ( .A1(n14265), .A2(n11311), .ZN(n14383) );
  NAND2_X1 U9117 ( .A1(n11305), .A2(n11304), .ZN(n15005) );
  NAND2_X1 U9118 ( .A1(n14265), .A2(n15005), .ZN(n14498) );
  INV_X1 U9119 ( .A(n15009), .ZN(n14889) );
  INV_X1 U9120 ( .A(n14383), .ZN(n15017) );
  OR2_X1 U9121 ( .A1(n10550), .A2(n10554), .ZN(n10832) );
  INV_X1 U9122 ( .A(n9825), .ZN(n14626) );
  NOR2_X1 U9123 ( .A1(n6868), .A2(n6864), .ZN(n6863) );
  INV_X1 U9124 ( .A(n6870), .ZN(n6864) );
  NOR2_X1 U9125 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n7211) );
  INV_X1 U9126 ( .A(n10554), .ZN(n14634) );
  INV_X1 U9127 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n10360) );
  NAND2_X1 U9128 ( .A1(n8483), .A2(n8482), .ZN(n8485) );
  XNOR2_X1 U9129 ( .A(n10187), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14641) );
  XNOR2_X1 U9130 ( .A(n9844), .B(n9843), .ZN(n11897) );
  INV_X1 U9131 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11234) );
  INV_X1 U9132 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n15512) );
  INV_X1 U9133 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11240) );
  INV_X1 U9134 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n15628) );
  INV_X1 U9135 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10566) );
  INV_X1 U9136 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10519) );
  NAND2_X1 U9137 ( .A1(n7043), .A2(n8023), .ZN(n8251) );
  INV_X1 U9138 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10504) );
  XNOR2_X1 U9139 ( .A(n14687), .B(n13529), .ZN(n15747) );
  INV_X1 U9140 ( .A(n7660), .ZN(n14693) );
  XNOR2_X1 U9141 ( .A(n14683), .B(n10442), .ZN(n15736) );
  XNOR2_X1 U9142 ( .A(n14697), .B(n7172), .ZN(n15739) );
  INV_X1 U9143 ( .A(n14698), .ZN(n7172) );
  XNOR2_X1 U9144 ( .A(n14700), .B(n7247), .ZN(n14768) );
  XNOR2_X1 U9145 ( .A(n14706), .B(n14704), .ZN(n15742) );
  INV_X1 U9146 ( .A(n14711), .ZN(n7248) );
  NAND2_X1 U9147 ( .A1(n7125), .A2(n7124), .ZN(n7654) );
  NAND2_X1 U9148 ( .A1(n7222), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7224) );
  NAND2_X1 U9149 ( .A1(n7658), .A2(n7656), .ZN(n7124) );
  INV_X1 U9150 ( .A(n7652), .ZN(n14722) );
  INV_X1 U9151 ( .A(n7650), .ZN(n14794) );
  NAND2_X1 U9152 ( .A1(n7082), .A2(n6626), .ZN(n7081) );
  NAND2_X1 U9153 ( .A1(n7400), .A2(n12861), .ZN(n7398) );
  NAND2_X1 U9154 ( .A1(n12639), .A2(n6569), .ZN(n7397) );
  INV_X1 U9155 ( .A(n6835), .ZN(n11858) );
  INV_X1 U9156 ( .A(n7686), .ZN(n11903) );
  INV_X1 U9157 ( .A(n7196), .ZN(n12395) );
  INV_X1 U9158 ( .A(n6778), .ZN(n12920) );
  NAND2_X1 U9159 ( .A1(n6966), .A2(n13023), .ZN(n12989) );
  AOI21_X1 U9160 ( .B1(n7135), .B2(n12995), .A(n7134), .ZN(n13027) );
  NAND2_X1 U9161 ( .A1(n6767), .A2(n6765), .ZN(P3_U3201) );
  NAND2_X1 U9162 ( .A1(n6768), .A2(n7667), .ZN(n6767) );
  NOR2_X1 U9163 ( .A1(n6704), .A2(n7179), .ZN(n7178) );
  NOR2_X1 U9164 ( .A1(n15419), .A2(n10392), .ZN(n7179) );
  MUX2_X1 U9165 ( .A(n13264), .B(n13326), .S(n15419), .Z(n13265) );
  NOR2_X1 U9166 ( .A1(n6705), .A2(n7181), .ZN(n7180) );
  NOR2_X1 U9167 ( .A1(n15407), .A2(n10410), .ZN(n7181) );
  OAI21_X1 U9168 ( .B1(n13326), .B2(n15409), .A(n6782), .ZN(P3_U3455) );
  AOI21_X1 U9169 ( .B1(n12646), .B2(n10411), .A(n6783), .ZN(n6782) );
  NOR2_X1 U9170 ( .A1(n15407), .A2(n13327), .ZN(n6783) );
  OAI21_X1 U9171 ( .B1(n13329), .B2(n15409), .A(n7161), .ZN(P3_U3454) );
  INV_X1 U9172 ( .A(n7162), .ZN(n7161) );
  OAI21_X1 U9173 ( .B1(n13330), .B2(n13376), .A(n7163), .ZN(n7162) );
  OR2_X1 U9174 ( .A1(n15407), .A2(n15657), .ZN(n7163) );
  NAND2_X1 U9175 ( .A1(n7202), .A2(n7201), .ZN(P2_U3186) );
  INV_X1 U9176 ( .A(n13396), .ZN(n7201) );
  INV_X1 U9177 ( .A(n7270), .ZN(P2_U3532) );
  AOI21_X1 U9178 ( .B1(n13526), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n7271), .ZN(
        n7270) );
  NOR2_X1 U9179 ( .A1(n13526), .A2(n7272), .ZN(n7271) );
  INV_X1 U9180 ( .A(n6746), .ZN(n13579) );
  NAND2_X1 U9181 ( .A1(n7184), .A2(n7182), .ZN(P2_U3236) );
  NAND2_X1 U9182 ( .A1(n7318), .A2(n13770), .ZN(n7184) );
  NOR2_X1 U9183 ( .A1(n7183), .A2(n7317), .ZN(n7182) );
  NAND2_X1 U9184 ( .A1(n7788), .A2(n7790), .ZN(n7318) );
  INV_X1 U9185 ( .A(n7787), .ZN(n7786) );
  AND2_X1 U9186 ( .A1(n6908), .A2(n9792), .ZN(n9796) );
  NAND2_X1 U9187 ( .A1(n6907), .A2(n15270), .ZN(n6906) );
  OAI21_X1 U9188 ( .B1(n14624), .B2(n13967), .A(n7249), .ZN(P2_U3297) );
  INV_X1 U9189 ( .A(n7250), .ZN(n7249) );
  OAI22_X1 U9190 ( .A1(n7975), .A2(P2_U3088), .B1(n13947), .B2(n13964), .ZN(
        n7250) );
  INV_X1 U9191 ( .A(n7156), .ZN(n7155) );
  OAI21_X1 U9192 ( .B1(n14286), .B2(n14864), .A(n13977), .ZN(n7156) );
  OAI211_X1 U9193 ( .C1(n7059), .C2(n12372), .A(n7055), .B(n7054), .ZN(
        P1_U3242) );
  NAND2_X1 U9194 ( .A1(n6672), .A2(n10357), .ZN(n7054) );
  NAND2_X1 U9195 ( .A1(n15105), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n7325) );
  OAI21_X1 U9196 ( .B1(n7371), .B2(n7327), .A(n15107), .ZN(n7326) );
  NOR2_X1 U9197 ( .A1(n14515), .A2(n14599), .ZN(n7327) );
  NAND2_X1 U9198 ( .A1(n15105), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n7725) );
  NAND2_X1 U9199 ( .A1(n14603), .A2(n15107), .ZN(n7726) );
  NAND2_X1 U9200 ( .A1(n15096), .A2(n15093), .ZN(n7452) );
  AOI21_X1 U9201 ( .B1(n7371), .B2(n15096), .A(n6738), .ZN(n7450) );
  NAND2_X1 U9202 ( .A1(n7657), .A2(n7655), .ZN(n14774) );
  AND2_X1 U9203 ( .A1(n7659), .A2(n6583), .ZN(n14776) );
  NOR2_X1 U9204 ( .A1(n14915), .A2(n14916), .ZN(n14914) );
  AND2_X1 U9205 ( .A1(n7034), .A2(n7035), .ZN(n14915) );
  INV_X1 U9206 ( .A(n14927), .ZN(n14926) );
  BUF_X2 U9207 ( .A(n9578), .Z(n9566) );
  INV_X1 U9208 ( .A(n14517), .ZN(n7158) );
  NAND2_X1 U9209 ( .A1(n7244), .A2(n10925), .ZN(n6559) );
  OR2_X1 U9210 ( .A1(n12253), .A2(n12121), .ZN(n6560) );
  INV_X1 U9211 ( .A(n11781), .ZN(n13922) );
  AND2_X1 U9212 ( .A1(n9321), .A2(n9320), .ZN(n9396) );
  INV_X1 U9213 ( .A(n9396), .ZN(n12527) );
  AND2_X1 U9214 ( .A1(n13407), .A2(n7638), .ZN(n7634) );
  INV_X1 U9215 ( .A(n11697), .ZN(n6801) );
  OR2_X1 U9216 ( .A1(n8033), .A2(n6830), .ZN(n8307) );
  NAND3_X2 U9217 ( .A1(n7110), .A2(n9894), .A3(n9896), .ZN(n11168) );
  INV_X1 U9218 ( .A(n7836), .ZN(n7835) );
  OAI21_X1 U9219 ( .B1(n14034), .B2(n12741), .A(n12752), .ZN(n7836) );
  OAI211_X1 U9220 ( .C1(n10777), .C2(n10733), .A(n8685), .B(n8686), .ZN(n15348) );
  INV_X1 U9221 ( .A(n15348), .ZN(n6805) );
  NOR2_X1 U9222 ( .A1(n13907), .A2(n13502), .ZN(n9719) );
  INV_X1 U9223 ( .A(n9486), .ZN(n7903) );
  INV_X1 U9224 ( .A(n9791), .ZN(n8105) );
  INV_X1 U9225 ( .A(n7386), .ZN(n7385) );
  OAI21_X1 U9226 ( .B1(n8810), .B2(n7387), .A(n8825), .ZN(n7386) );
  AND2_X1 U9227 ( .A1(n6669), .A2(n7276), .ZN(n6561) );
  NAND2_X1 U9228 ( .A1(n13830), .A2(n6912), .ZN(n6562) );
  OR2_X1 U9229 ( .A1(n12929), .A2(n12928), .ZN(n6563) );
  INV_X1 U9230 ( .A(n11073), .ZN(n7245) );
  NAND2_X1 U9231 ( .A1(n6955), .A2(n6956), .ZN(n11557) );
  AND2_X1 U9232 ( .A1(n12638), .A2(n12830), .ZN(n6564) );
  INV_X1 U9233 ( .A(n10925), .ZN(n7480) );
  AND2_X1 U9234 ( .A1(n6665), .A2(n7313), .ZN(n6565) );
  NAND2_X1 U9235 ( .A1(n8316), .A2(n8315), .ZN(n12253) );
  AND2_X1 U9236 ( .A1(n7876), .A2(n6703), .ZN(n6566) );
  AND3_X1 U9237 ( .A1(n9639), .A2(n9786), .A3(n7111), .ZN(n6567) );
  NOR2_X1 U9238 ( .A1(n7777), .A2(n7775), .ZN(n6568) );
  NOR2_X1 U9239 ( .A1(n7399), .A2(n15434), .ZN(n6569) );
  XOR2_X1 U9240 ( .A(n10378), .B(n9145), .Z(n6570) );
  INV_X1 U9241 ( .A(n7637), .ZN(n7636) );
  NAND2_X1 U9242 ( .A1(n13474), .A2(n8425), .ZN(n7637) );
  XOR2_X1 U9243 ( .A(n13035), .B(n13034), .Z(n6571) );
  OR2_X1 U9244 ( .A1(n10297), .A2(n7060), .ZN(n6572) );
  AND2_X1 U9245 ( .A1(n7119), .A2(n7063), .ZN(n6573) );
  NAND2_X1 U9246 ( .A1(n9818), .A2(n9817), .ZN(n14517) );
  AND2_X1 U9247 ( .A1(n9855), .A2(n9854), .ZN(n14297) );
  INV_X1 U9248 ( .A(n10032), .ZN(n7572) );
  AND2_X1 U9249 ( .A1(n7754), .A2(n7495), .ZN(n6575) );
  AND2_X1 U9250 ( .A1(n7448), .A2(n14257), .ZN(n6576) );
  OR2_X1 U9251 ( .A1(n8133), .A2(n10495), .ZN(n6577) );
  NAND2_X1 U9252 ( .A1(n8295), .A2(n8294), .ZN(n12214) );
  NAND2_X1 U9253 ( .A1(n13483), .A2(n7627), .ZN(n6578) );
  NAND2_X1 U9254 ( .A1(n8487), .A2(n8486), .ZN(n13870) );
  INV_X1 U9255 ( .A(n13870), .ZN(n7784) );
  AND2_X1 U9256 ( .A1(n12878), .A2(n13218), .ZN(n6579) );
  NAND2_X1 U9257 ( .A1(n7534), .A2(n7532), .ZN(n12526) );
  INV_X1 U9258 ( .A(n12646), .ZN(n13328) );
  NAND2_X1 U9259 ( .A1(n7390), .A2(n9193), .ZN(n12646) );
  AND2_X1 U9260 ( .A1(n7676), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n6580) );
  INV_X1 U9261 ( .A(n10891), .ZN(n6773) );
  INV_X2 U9262 ( .A(n8675), .ZN(n7522) );
  AND3_X1 U9263 ( .A1(n7654), .A2(n7657), .A3(n7224), .ZN(n6581) );
  NAND2_X1 U9264 ( .A1(n9149), .A2(n8646), .ZN(n6582) );
  OR2_X1 U9265 ( .A1(n14713), .A2(n14714), .ZN(n6583) );
  INV_X1 U9266 ( .A(n6549), .ZN(n9861) );
  AND4_X1 U9267 ( .A1(n8645), .A2(n15717), .A3(n8644), .A4(n15715), .ZN(n6584)
         );
  INV_X1 U9268 ( .A(n8137), .ZN(n8492) );
  NAND2_X1 U9269 ( .A1(n8675), .A2(n10485), .ZN(n8722) );
  INV_X1 U9270 ( .A(n13519), .ZN(n7319) );
  AND2_X1 U9271 ( .A1(n15311), .A2(n12018), .ZN(n6585) );
  AND2_X1 U9272 ( .A1(n8178), .A2(n8081), .ZN(n8180) );
  INV_X1 U9273 ( .A(n13447), .ZN(n6998) );
  NAND2_X1 U9274 ( .A1(n8111), .A2(n7952), .ZN(n8129) );
  OR2_X1 U9275 ( .A1(n14892), .A2(n14100), .ZN(n6586) );
  AND2_X1 U9276 ( .A1(n13117), .A2(n9248), .ZN(n6587) );
  INV_X1 U9277 ( .A(n7781), .ZN(n7780) );
  NOR2_X1 U9278 ( .A1(n9729), .A2(n13668), .ZN(n7781) );
  AND2_X1 U9279 ( .A1(n9357), .A2(n12896), .ZN(n6588) );
  NOR2_X1 U9280 ( .A1(n9080), .A2(n8703), .ZN(n6589) );
  AND2_X1 U9281 ( .A1(n9513), .A2(n9512), .ZN(n6590) );
  AND2_X1 U9282 ( .A1(n15008), .A2(n11595), .ZN(n6591) );
  NOR2_X1 U9283 ( .A1(n13628), .A2(n7170), .ZN(n6592) );
  OR2_X1 U9284 ( .A1(n9218), .A2(n10756), .ZN(n6593) );
  AND2_X1 U9285 ( .A1(n9613), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6594) );
  NAND2_X1 U9286 ( .A1(n15008), .A2(n14106), .ZN(n6595) );
  NAND2_X1 U9287 ( .A1(n13783), .A2(n13797), .ZN(n6596) );
  AND2_X1 U9288 ( .A1(n9814), .A2(n9813), .ZN(n9836) );
  AND2_X1 U9289 ( .A1(n9494), .A2(n9493), .ZN(n6597) );
  AND2_X1 U9290 ( .A1(n9541), .A2(n9540), .ZN(n6598) );
  AND2_X1 U9291 ( .A1(n9565), .A2(n9564), .ZN(n6599) );
  NOR2_X1 U9292 ( .A1(n7903), .A2(n6645), .ZN(n6600) );
  INV_X1 U9293 ( .A(n12164), .ZN(n7712) );
  NAND2_X1 U9294 ( .A1(n14646), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n6601) );
  AND2_X1 U9295 ( .A1(n14847), .A2(n13500), .ZN(n6602) );
  AND2_X1 U9296 ( .A1(n6890), .A2(n6893), .ZN(n6603) );
  OR2_X1 U9297 ( .A1(n6559), .A2(n11073), .ZN(n6604) );
  AND2_X1 U9298 ( .A1(n7578), .A2(n9975), .ZN(n6605) );
  INV_X1 U9299 ( .A(n8642), .ZN(n8772) );
  AND2_X1 U9300 ( .A1(n10495), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6606) );
  OR2_X1 U9301 ( .A1(n14647), .A2(n7174), .ZN(n6607) );
  NAND2_X1 U9302 ( .A1(n8797), .A2(n15707), .ZN(n8811) );
  OR2_X1 U9303 ( .A1(n13767), .A2(n13515), .ZN(n6608) );
  OAI21_X1 U9304 ( .B1(n14624), .B2(n9610), .A(n9611), .ZN(n13593) );
  XNOR2_X1 U9305 ( .A(n9842), .B(P1_IR_REG_21__SCAN_IN), .ZN(n10700) );
  OR2_X1 U9306 ( .A1(n13581), .A2(n13578), .ZN(n6609) );
  AND2_X1 U9307 ( .A1(n13875), .A2(n13684), .ZN(n6610) );
  NAND2_X1 U9308 ( .A1(n13341), .A2(n13131), .ZN(n6611) );
  AND2_X1 U9309 ( .A1(n14339), .A2(n14094), .ZN(n6612) );
  AND2_X1 U9310 ( .A1(n8249), .A2(n8248), .ZN(n6613) );
  AND2_X1 U9311 ( .A1(n13031), .A2(n13030), .ZN(n6614) );
  NAND2_X1 U9312 ( .A1(n13183), .A2(n9142), .ZN(n13169) );
  INV_X1 U9313 ( .A(n13593), .ZN(n13841) );
  INV_X1 U9314 ( .A(n9312), .ZN(n7883) );
  NAND2_X1 U9315 ( .A1(n10229), .A2(n10228), .ZN(n14535) );
  INV_X1 U9316 ( .A(n14535), .ZN(n7335) );
  AND2_X1 U9317 ( .A1(n10206), .A2(n7559), .ZN(n6615) );
  NAND2_X1 U9318 ( .A1(n8373), .A2(n8372), .ZN(n13912) );
  AND2_X1 U9319 ( .A1(n9374), .A2(n9375), .ZN(n6616) );
  INV_X1 U9320 ( .A(n14257), .ZN(n7449) );
  INV_X1 U9321 ( .A(n13875), .ZN(n7497) );
  INV_X1 U9322 ( .A(n14034), .ZN(n7837) );
  NAND4_X1 U9323 ( .A1(n8655), .A2(n8654), .A3(n6593), .A4(n8653), .ZN(n15344)
         );
  OR2_X1 U9324 ( .A1(n7335), .A2(n14325), .ZN(n6617) );
  AND2_X1 U9325 ( .A1(n13455), .A2(n13456), .ZN(n13453) );
  AND2_X1 U9326 ( .A1(n7410), .A2(n7408), .ZN(n6618) );
  AND4_X1 U9327 ( .A1(n12193), .A2(n7138), .A3(n12005), .A4(n12004), .ZN(n6619) );
  AND2_X1 U9328 ( .A1(n12102), .A2(n13517), .ZN(n6620) );
  NAND2_X1 U9329 ( .A1(n14892), .A2(n12030), .ZN(n6621) );
  XNOR2_X1 U9330 ( .A(n11611), .B(n7319), .ZN(n11604) );
  INV_X1 U9331 ( .A(n11604), .ZN(n7803) );
  OR2_X1 U9332 ( .A1(n11168), .A2(n11463), .ZN(n11111) );
  NAND2_X1 U9333 ( .A1(n7320), .A2(n8240), .ZN(n11611) );
  NAND2_X1 U9334 ( .A1(n10114), .A2(n10113), .ZN(n14585) );
  AND2_X1 U9335 ( .A1(n12565), .A2(n10308), .ZN(n14300) );
  INV_X1 U9336 ( .A(n14300), .ZN(n7444) );
  OR2_X1 U9337 ( .A1(n9538), .A2(n9537), .ZN(n6622) );
  NOR2_X1 U9338 ( .A1(n12329), .A2(n12013), .ZN(n6623) );
  NOR2_X1 U9339 ( .A1(n8139), .A2(n10424), .ZN(n6624) );
  INV_X1 U9340 ( .A(n7880), .ZN(n7879) );
  OAI21_X1 U9341 ( .B1(n12527), .B2(n7881), .A(n9321), .ZN(n7880) );
  AND2_X1 U9342 ( .A1(n12623), .A2(n12871), .ZN(n6625) );
  AND2_X1 U9343 ( .A1(n10163), .A2(n10162), .ZN(n14401) );
  INV_X1 U9344 ( .A(n14401), .ZN(n14566) );
  OR2_X1 U9345 ( .A1(n12797), .A2(n6564), .ZN(n6626) );
  AND2_X1 U9346 ( .A1(n7052), .A2(n10218), .ZN(n6627) );
  NOR2_X1 U9347 ( .A1(n12594), .A2(n7442), .ZN(n7441) );
  AND2_X1 U9348 ( .A1(n7627), .A2(n7630), .ZN(n6628) );
  INV_X1 U9349 ( .A(n12565), .ZN(n7368) );
  AND2_X1 U9350 ( .A1(n9725), .A2(n13740), .ZN(n6629) );
  AND2_X1 U9351 ( .A1(n11646), .A2(n11645), .ZN(n6630) );
  AND2_X1 U9352 ( .A1(n7564), .A2(n10018), .ZN(n6631) );
  NOR2_X1 U9353 ( .A1(n14035), .A2(n14034), .ZN(n6632) );
  INV_X1 U9354 ( .A(n7799), .ZN(n7798) );
  AND2_X1 U9355 ( .A1(n7413), .A2(n7412), .ZN(n6633) );
  AND2_X1 U9356 ( .A1(n7569), .A2(n10055), .ZN(n6634) );
  AND2_X1 U9357 ( .A1(n14286), .A2(n14076), .ZN(n6635) );
  OR2_X1 U9358 ( .A1(n7487), .A2(n12394), .ZN(n6636) );
  OR2_X1 U9359 ( .A1(n7487), .A2(n12381), .ZN(n6637) );
  AND2_X1 U9360 ( .A1(n9836), .A2(n9840), .ZN(n6638) );
  AND2_X1 U9361 ( .A1(n6596), .A2(n7805), .ZN(n6639) );
  INV_X1 U9362 ( .A(n7518), .ZN(n7517) );
  INV_X1 U9363 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9840) );
  INV_X1 U9364 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n15706) );
  INV_X1 U9365 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n7663) );
  NAND2_X1 U9366 ( .A1(n8675), .A2(n7519), .ZN(n6640) );
  AND2_X1 U9367 ( .A1(n6999), .A2(n6998), .ZN(n6641) );
  AND2_X1 U9368 ( .A1(n7543), .A2(n7541), .ZN(n6642) );
  INV_X1 U9369 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7737) );
  NAND2_X1 U9370 ( .A1(n7312), .A2(n6565), .ZN(n6643) );
  NAND3_X2 U9371 ( .A1(n9865), .A2(n7438), .A3(n7437), .ZN(n11440) );
  NOR2_X1 U9372 ( .A1(n12476), .A2(n14099), .ZN(n6644) );
  INV_X1 U9373 ( .A(n7702), .ZN(n7696) );
  NAND2_X1 U9374 ( .A1(n14352), .A2(n7703), .ZN(n7702) );
  AND2_X1 U9375 ( .A1(n9485), .A2(n9484), .ZN(n6645) );
  NOR2_X1 U9376 ( .A1(n14595), .A2(n14097), .ZN(n6646) );
  NOR2_X1 U9377 ( .A1(n11611), .A2(n7319), .ZN(n6647) );
  INV_X1 U9378 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9819) );
  INV_X1 U9379 ( .A(n7516), .ZN(n7513) );
  OR2_X1 U9380 ( .A1(n13093), .A2(n13104), .ZN(n7516) );
  INV_X1 U9381 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10495) );
  AND3_X1 U9382 ( .A1(n9884), .A2(n9882), .A3(n9885), .ZN(n6648) );
  AND2_X1 U9383 ( .A1(n8045), .A2(n8044), .ZN(n6649) );
  AND2_X1 U9384 ( .A1(n12637), .A2(n13089), .ZN(n6650) );
  INV_X1 U9385 ( .A(n13644), .ZN(n13855) );
  AND2_X1 U9386 ( .A1(n8078), .A2(n8077), .ZN(n13644) );
  AND2_X1 U9387 ( .A1(n6882), .A2(n6880), .ZN(n6652) );
  INV_X1 U9388 ( .A(n7937), .ZN(n7723) );
  AND2_X1 U9389 ( .A1(n7216), .A2(n7570), .ZN(n6653) );
  AND2_X1 U9390 ( .A1(n8012), .A2(SI_5_), .ZN(n6654) );
  NAND2_X1 U9391 ( .A1(n9843), .A2(n9840), .ZN(n6655) );
  INV_X1 U9392 ( .A(n7533), .ZN(n7532) );
  NAND2_X1 U9393 ( .A1(n12527), .A2(n9132), .ZN(n7533) );
  INV_X1 U9394 ( .A(n6941), .ZN(n6940) );
  NAND2_X1 U9395 ( .A1(n7851), .A2(n6942), .ZN(n6941) );
  AND2_X1 U9396 ( .A1(n10566), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n6656) );
  NAND2_X1 U9397 ( .A1(n9776), .A2(n13881), .ZN(n6657) );
  AND2_X1 U9398 ( .A1(n8680), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n6658) );
  INV_X1 U9399 ( .A(n7760), .ZN(n7759) );
  OAI21_X1 U9400 ( .B1(n8386), .B2(n7761), .A(n8405), .ZN(n7760) );
  AND2_X1 U9401 ( .A1(n8040), .A2(n8039), .ZN(n6659) );
  AND2_X1 U9402 ( .A1(n9465), .A2(n9464), .ZN(n6660) );
  INV_X1 U9403 ( .A(n12844), .ZN(n7426) );
  OR2_X1 U9404 ( .A1(n11719), .A2(n14105), .ZN(n6661) );
  AND2_X1 U9405 ( .A1(n9375), .A2(n10731), .ZN(n6662) );
  INV_X1 U9406 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10573) );
  AND2_X1 U9407 ( .A1(n6597), .A2(n7931), .ZN(n6663) );
  INV_X1 U9408 ( .A(n14522), .ZN(n14286) );
  NAND2_X1 U9409 ( .A1(n10239), .A2(n10238), .ZN(n14522) );
  INV_X1 U9410 ( .A(n7402), .ZN(n7401) );
  OAI21_X1 U9411 ( .B1(n7410), .B2(n7404), .A(n7403), .ZN(n7402) );
  NOR2_X1 U9412 ( .A1(n10069), .A2(n10070), .ZN(n6664) );
  NAND2_X1 U9413 ( .A1(n13879), .A2(n13469), .ZN(n6665) );
  NAND2_X2 U9414 ( .A1(n8625), .A2(n13955), .ZN(n8126) );
  INV_X1 U9415 ( .A(n7705), .ZN(n7704) );
  NAND2_X1 U9416 ( .A1(n8037), .A2(n8036), .ZN(n6666) );
  INV_X1 U9417 ( .A(n10204), .ZN(n7559) );
  AND2_X1 U9418 ( .A1(n7596), .A2(n9777), .ZN(n6667) );
  XOR2_X1 U9419 ( .A(n13593), .B(n9734), .Z(n6668) );
  INV_X1 U9420 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7922) );
  INV_X1 U9421 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7968) );
  OR2_X1 U9422 ( .A1(n6597), .A2(n7931), .ZN(n6669) );
  INV_X1 U9423 ( .A(n10005), .ZN(n7568) );
  AND2_X1 U9424 ( .A1(n13490), .A2(n8532), .ZN(n6670) );
  OR2_X1 U9425 ( .A1(n7459), .A2(n14415), .ZN(n6671) );
  INV_X1 U9426 ( .A(n7628), .ZN(n7627) );
  OR2_X1 U9427 ( .A1(n13391), .A2(n7629), .ZN(n7628) );
  INV_X1 U9428 ( .A(n7843), .ZN(n7842) );
  NAND2_X1 U9429 ( .A1(n7846), .A2(n7844), .ZN(n7843) );
  INV_X1 U9430 ( .A(n7854), .ZN(n7853) );
  NAND2_X1 U9431 ( .A1(n11674), .A2(n11666), .ZN(n7854) );
  NAND2_X1 U9432 ( .A1(n10353), .A2(n10352), .ZN(n6672) );
  INV_X1 U9433 ( .A(n10175), .ZN(n7072) );
  INV_X1 U9434 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8661) );
  INV_X1 U9435 ( .A(n9778), .ZN(n13679) );
  AND3_X1 U9436 ( .A1(n9370), .A2(n9369), .A3(n13092), .ZN(n6673) );
  OR2_X1 U9437 ( .A1(n12929), .A2(n12919), .ZN(n6674) );
  OR2_X1 U9438 ( .A1(n8035), .A2(SI_14_), .ZN(n6675) );
  OR2_X1 U9439 ( .A1(n7128), .A2(n10730), .ZN(n6676) );
  AND2_X1 U9440 ( .A1(n8549), .A2(n8561), .ZN(n6677) );
  AND3_X1 U9441 ( .A1(n8791), .A2(n8638), .A3(n8912), .ZN(n6678) );
  INV_X1 U9442 ( .A(n12566), .ZN(n7369) );
  AND2_X1 U9443 ( .A1(n9249), .A2(n9252), .ZN(n13117) );
  INV_X1 U9444 ( .A(n13117), .ZN(n7542) );
  AND2_X1 U9445 ( .A1(n13130), .A2(n9248), .ZN(n6679) );
  NOR2_X1 U9446 ( .A1(n13175), .A2(n7895), .ZN(n7894) );
  OR2_X1 U9447 ( .A1(n15321), .A2(n6922), .ZN(n6680) );
  AND2_X1 U9448 ( .A1(n6595), .A2(n11589), .ZN(n6681) );
  NAND4_X1 U9449 ( .A1(n8756), .A2(n8755), .A3(n8754), .A4(n8753), .ZN(n15310)
         );
  OR2_X1 U9450 ( .A1(n7358), .A2(n6612), .ZN(n6682) );
  INV_X1 U9451 ( .A(n9492), .ZN(n7277) );
  NAND3_X1 U9452 ( .A1(n7966), .A2(n7986), .A3(n7610), .ZN(n8071) );
  AND2_X1 U9453 ( .A1(n7236), .A2(n7113), .ZN(n6683) );
  INV_X1 U9454 ( .A(n9792), .ZN(n9793) );
  NOR2_X1 U9455 ( .A1(n12609), .A2(n7751), .ZN(n9792) );
  AND2_X1 U9456 ( .A1(n7453), .A2(n7449), .ZN(n6684) );
  AND2_X1 U9457 ( .A1(n7164), .A2(n8344), .ZN(n6685) );
  NAND2_X1 U9458 ( .A1(n13903), .A2(n13442), .ZN(n6686) );
  AND2_X1 U9459 ( .A1(n6759), .A2(n7678), .ZN(n6687) );
  NAND2_X1 U9460 ( .A1(n10573), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6688) );
  AND2_X1 U9461 ( .A1(n6857), .A2(n7466), .ZN(n6689) );
  AND2_X1 U9462 ( .A1(n9652), .A2(n9651), .ZN(n6690) );
  AND2_X1 U9463 ( .A1(n6575), .A2(n13841), .ZN(n6691) );
  INV_X1 U9464 ( .A(n7421), .ZN(n7420) );
  OR2_X1 U9465 ( .A1(n12820), .A2(n7422), .ZN(n7421) );
  INV_X1 U9466 ( .A(n9719), .ZN(n7310) );
  NAND2_X1 U9467 ( .A1(n12797), .A2(n12888), .ZN(n6692) );
  INV_X1 U9468 ( .A(n11211), .ZN(n7479) );
  INV_X1 U9469 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n15461) );
  INV_X1 U9470 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7967) );
  INV_X1 U9471 ( .A(n14874), .ZN(n7850) );
  INV_X1 U9472 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7991) );
  NOR2_X1 U9473 ( .A1(n7921), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n6693) );
  OR2_X1 U9474 ( .A1(n7266), .A2(n9508), .ZN(n6694) );
  INV_X1 U9475 ( .A(n8699), .ZN(n9203) );
  NAND2_X1 U9476 ( .A1(n7177), .A2(n10086), .ZN(n14595) );
  INV_X1 U9477 ( .A(n14595), .ZN(n7116) );
  NAND2_X1 U9478 ( .A1(n11886), .A2(n7721), .ZN(n7724) );
  XNOR2_X1 U9479 ( .A(n8558), .B(n8557), .ZN(n12536) );
  AND2_X1 U9480 ( .A1(n7827), .A2(n7826), .ZN(n6695) );
  INV_X1 U9481 ( .A(n12802), .ZN(n13330) );
  NAND2_X1 U9482 ( .A1(n9077), .A2(n9076), .ZN(n12802) );
  AND2_X1 U9483 ( .A1(n14467), .A2(n7338), .ZN(n6696) );
  XOR2_X1 U9484 ( .A(n12640), .B(n13248), .Z(n12610) );
  INV_X1 U9485 ( .A(n14760), .ZN(n7487) );
  INV_X1 U9486 ( .A(n13495), .ZN(n7644) );
  NAND2_X1 U9487 ( .A1(n14756), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n6697) );
  AND2_X1 U9488 ( .A1(n14756), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6698) );
  OR2_X1 U9489 ( .A1(n13448), .A2(n13447), .ZN(n7001) );
  NAND2_X1 U9490 ( .A1(n7526), .A2(n9128), .ZN(n14807) );
  NAND2_X1 U9491 ( .A1(n9131), .A2(n9130), .ZN(n12458) );
  OR2_X1 U9492 ( .A1(n13418), .A2(n13690), .ZN(n6699) );
  AND2_X1 U9493 ( .A1(n13072), .A2(n15360), .ZN(n6700) );
  AND2_X1 U9494 ( .A1(n15282), .A2(n12334), .ZN(n6701) );
  INV_X1 U9495 ( .A(n11873), .ZN(n11913) );
  INV_X1 U9496 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7886) );
  NAND2_X1 U9497 ( .A1(n9626), .A2(n9625), .ZN(n12603) );
  INV_X1 U9498 ( .A(n12603), .ZN(n7495) );
  INV_X1 U9499 ( .A(n8348), .ZN(n8035) );
  AND2_X1 U9500 ( .A1(n14591), .A2(n14478), .ZN(n6702) );
  INV_X1 U9501 ( .A(n12931), .ZN(n7478) );
  AND4_X1 U9502 ( .A1(n9853), .A2(n9852), .A3(n9851), .A4(n9850), .ZN(n14275)
         );
  INV_X1 U9503 ( .A(n14275), .ZN(n7446) );
  OR2_X1 U9504 ( .A1(n12367), .A2(n6918), .ZN(n6703) );
  AND2_X1 U9505 ( .A1(n10393), .A2(n9187), .ZN(n6704) );
  AND2_X1 U9506 ( .A1(n10393), .A2(n10411), .ZN(n6705) );
  INV_X1 U9507 ( .A(n7500), .ZN(n13748) );
  INV_X1 U9508 ( .A(SI_12_), .ZN(n6830) );
  AND2_X1 U9509 ( .A1(n7470), .A2(n7468), .ZN(n6706) );
  AND2_X1 U9510 ( .A1(n12576), .A2(n7464), .ZN(n6707) );
  AND2_X1 U9511 ( .A1(n7896), .A2(n7894), .ZN(n6708) );
  INV_X1 U9512 ( .A(n7496), .ZN(n13823) );
  NOR2_X2 U9513 ( .A1(n12445), .A2(n14847), .ZN(n7496) );
  INV_X1 U9514 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7174) );
  AND2_X1 U9515 ( .A1(n12862), .A2(n7420), .ZN(n6709) );
  INV_X1 U9516 ( .A(n13202), .ZN(n13195) );
  AND2_X1 U9517 ( .A1(n9338), .A2(n9341), .ZN(n13202) );
  INV_X1 U9518 ( .A(n7823), .ZN(n7821) );
  NAND2_X1 U9519 ( .A1(n12704), .A2(n7824), .ZN(n7823) );
  NOR2_X1 U9520 ( .A1(n13375), .A2(n13244), .ZN(n6710) );
  AND2_X1 U9521 ( .A1(n13289), .A2(n13187), .ZN(n6711) );
  AND2_X1 U9522 ( .A1(n7534), .A2(n9132), .ZN(n6712) );
  AND2_X1 U9523 ( .A1(n10571), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n6713) );
  AND2_X1 U9524 ( .A1(n6978), .A2(n6596), .ZN(n6714) );
  INV_X1 U9525 ( .A(n9288), .ZN(n6922) );
  INV_X1 U9526 ( .A(n11916), .ZN(n7488) );
  AND2_X1 U9527 ( .A1(n12119), .A2(n7797), .ZN(n6715) );
  OR2_X1 U9528 ( .A1(n12614), .A2(n13245), .ZN(n6716) );
  INV_X1 U9529 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n15654) );
  AND2_X1 U9530 ( .A1(n7240), .A2(n6563), .ZN(n6717) );
  INV_X1 U9531 ( .A(n8307), .ZN(n7779) );
  AND2_X1 U9532 ( .A1(n6752), .A2(n6751), .ZN(n6718) );
  AND2_X1 U9533 ( .A1(n10408), .A2(n10407), .ZN(n15409) );
  INV_X1 U9534 ( .A(n6557), .ZN(n8415) );
  NOR2_X2 U9535 ( .A1(n8618), .A2(n8606), .ZN(n15120) );
  AND2_X1 U9536 ( .A1(n11444), .A2(n8247), .ZN(n6719) );
  NAND2_X1 U9537 ( .A1(n11292), .A2(n9713), .ZN(n11844) );
  INV_X1 U9538 ( .A(n12396), .ZN(n14765) );
  OAI21_X1 U9539 ( .B1(n7620), .B2(n7619), .A(n15108), .ZN(n12055) );
  XNOR2_X1 U9540 ( .A(n10363), .B(P1_IR_REG_24__SCAN_IN), .ZN(n10550) );
  INV_X1 U9541 ( .A(n14873), .ZN(n7848) );
  AND2_X1 U9542 ( .A1(n13041), .A2(n13030), .ZN(n6720) );
  NAND2_X1 U9543 ( .A1(n7855), .A2(n7853), .ZN(n12292) );
  NAND2_X1 U9544 ( .A1(n7331), .A2(n7330), .ZN(n11937) );
  INV_X1 U9545 ( .A(n11937), .ZN(n7329) );
  INV_X1 U9546 ( .A(n7331), .ZN(n11938) );
  NAND2_X1 U9547 ( .A1(n6802), .A2(n6803), .ZN(n8910) );
  AND2_X1 U9548 ( .A1(n7131), .A2(n7105), .ZN(n6721) );
  INV_X1 U9549 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7247) );
  INV_X1 U9550 ( .A(n7745), .ZN(n7744) );
  NOR2_X1 U9551 ( .A1(n8534), .A2(n12455), .ZN(n7745) );
  NOR2_X1 U9552 ( .A1(n8535), .A2(SI_26_), .ZN(n6722) );
  INV_X1 U9553 ( .A(n8468), .ZN(n8056) );
  NAND4_X1 U9554 ( .A1(n8643), .A2(n8642), .A3(n6584), .A4(n7886), .ZN(n6723)
         );
  NOR2_X1 U9555 ( .A1(n6722), .A2(n6825), .ZN(n6824) );
  NAND2_X1 U9556 ( .A1(n7845), .A2(n7842), .ZN(n6724) );
  NOR2_X1 U9557 ( .A1(n7677), .A2(n12971), .ZN(n6725) );
  AND2_X1 U9558 ( .A1(n7489), .A2(n7488), .ZN(n6726) );
  AND2_X1 U9559 ( .A1(n7242), .A2(n11557), .ZN(n6727) );
  AND2_X1 U9560 ( .A1(n11694), .A2(n9122), .ZN(n6728) );
  AND2_X1 U9561 ( .A1(n7686), .A2(n7685), .ZN(n6729) );
  AND2_X1 U9562 ( .A1(n7684), .A2(n11553), .ZN(n6730) );
  INV_X1 U9563 ( .A(n7679), .ZN(n7677) );
  NAND2_X1 U9564 ( .A1(n12954), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7679) );
  OR2_X1 U9565 ( .A1(n12396), .A2(n12365), .ZN(n6731) );
  INV_X1 U9566 ( .A(n15096), .ZN(n7451) );
  INV_X1 U9567 ( .A(n15282), .ZN(n7100) );
  NAND2_X1 U9568 ( .A1(n9698), .A2(n9667), .ZN(n9617) );
  AND2_X2 U9569 ( .A1(n11197), .A2(n11196), .ZN(n15279) );
  NAND4_X1 U9570 ( .A1(n8679), .A2(n8678), .A3(n8676), .A4(n8677), .ZN(n15423)
         );
  INV_X1 U9571 ( .A(n15423), .ZN(n6804) );
  AND2_X1 U9572 ( .A1(n15280), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n6732) );
  AND2_X1 U9573 ( .A1(n12999), .A2(n12998), .ZN(n6733) );
  AND2_X1 U9574 ( .A1(n13506), .A2(n13922), .ZN(n6734) );
  AND2_X1 U9575 ( .A1(n13008), .A2(n13007), .ZN(n6735) );
  NAND2_X1 U9576 ( .A1(n11653), .A2(n11654), .ZN(n6736) );
  AND2_X1 U9577 ( .A1(n15279), .A2(n13819), .ZN(n6737) );
  AND2_X1 U9578 ( .A1(n7451), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6738) );
  AND2_X1 U9579 ( .A1(n11414), .A2(n15120), .ZN(n6739) );
  AND2_X1 U9580 ( .A1(n7246), .A2(n7245), .ZN(n6740) );
  XNOR2_X1 U9581 ( .A(n8965), .B(n9089), .ZN(n13033) );
  NAND2_X1 U9582 ( .A1(n8140), .A2(n6985), .ZN(n13525) );
  INV_X1 U9583 ( .A(n13525), .ZN(n6984) );
  NOR2_X1 U9584 ( .A1(n9822), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n14616) );
  NAND2_X1 U9585 ( .A1(n6775), .A2(n6774), .ZN(n6741) );
  AND2_X1 U9586 ( .A1(n8104), .A2(n8103), .ZN(n6742) );
  INV_X1 U9587 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7653) );
  INV_X1 U9588 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7173) );
  INV_X1 U9589 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7662) );
  INV_X1 U9590 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7608) );
  INV_X1 U9591 ( .A(n13127), .ZN(n6928) );
  NOR2_X1 U9592 ( .A1(n13127), .A2(n7547), .ZN(n7546) );
  NAND2_X1 U9593 ( .A1(n13128), .A2(n13127), .ZN(n13130) );
  XNOR2_X1 U9594 ( .A(n13031), .B(n13030), .ZN(n13009) );
  XNOR2_X1 U9595 ( .A(n12968), .B(n12977), .ZN(n12950) );
  NAND2_X1 U9596 ( .A1(n11900), .A2(n7685), .ZN(n6754) );
  INV_X1 U9597 ( .A(n11901), .ZN(n6755) );
  INV_X1 U9598 ( .A(n11900), .ZN(n6756) );
  NAND2_X1 U9599 ( .A1(n6764), .A2(n7675), .ZN(n7678) );
  INV_X1 U9600 ( .A(n12979), .ZN(n6759) );
  NOR2_X1 U9601 ( .A1(n6761), .A2(n12981), .ZN(n6760) );
  INV_X1 U9602 ( .A(n12981), .ZN(n6762) );
  AND2_X1 U9603 ( .A1(n12998), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n6763) );
  NAND2_X1 U9604 ( .A1(n6774), .A2(n11092), .ZN(n6771) );
  INV_X1 U9605 ( .A(n10890), .ZN(n6774) );
  INV_X1 U9606 ( .A(n6775), .ZN(n11091) );
  OAI21_X1 U9607 ( .B1(n6781), .B2(n10988), .A(n10739), .ZN(n10960) );
  AND3_X2 U9608 ( .A1(n7884), .A2(n8643), .A3(n8642), .ZN(n9149) );
  NAND4_X1 U9609 ( .A1(n7884), .A2(n8643), .A3(n8642), .A4(n7429), .ZN(n9147)
         );
  NAND2_X1 U9611 ( .A1(n6809), .A2(n9609), .ZN(n14624) );
  NAND2_X1 U9612 ( .A1(n9608), .A2(n9607), .ZN(n6809) );
  NAND3_X1 U9613 ( .A1(n7273), .A2(n6812), .A3(n6810), .ZN(n9701) );
  INV_X1 U9614 ( .A(n7773), .ZN(n7772) );
  NAND3_X1 U9615 ( .A1(n6815), .A2(n6675), .A3(n6814), .ZN(n7773) );
  NAND2_X1 U9616 ( .A1(n7775), .A2(n6816), .ZN(n6815) );
  INV_X1 U9617 ( .A(n8034), .ZN(n6816) );
  NAND2_X1 U9618 ( .A1(n6817), .A2(n6824), .ZN(n6822) );
  NAND3_X1 U9619 ( .A1(n6822), .A2(n7744), .A3(n6820), .ZN(n9589) );
  NAND2_X1 U9620 ( .A1(n7768), .A2(n8503), .ZN(n6823) );
  NAND3_X1 U9621 ( .A1(n6822), .A2(n6819), .A3(n6820), .ZN(n6818) );
  NAND2_X1 U9622 ( .A1(n8057), .A2(n6827), .ZN(n6826) );
  OAI21_X1 U9623 ( .B1(n8058), .B2(n8060), .A(n8061), .ZN(n6829) );
  NAND2_X1 U9624 ( .A1(n8470), .A2(n8058), .ZN(n8483) );
  OAI21_X1 U9625 ( .B1(n8013), .B2(P1_DATAO_REG_12__SCAN_IN), .A(n6831), .ZN(
        n8033) );
  NAND2_X1 U9626 ( .A1(n8013), .A2(n15628), .ZN(n6831) );
  OAI22_X2 U9627 ( .A1(n12389), .A2(n12388), .B1(n12387), .B2(n14760), .ZN(
        n12390) );
  OR2_X2 U9629 ( .A1(n12997), .A2(n6733), .ZN(n6837) );
  NAND4_X1 U9630 ( .A1(n7884), .A2(n8642), .A3(n7427), .A4(n8643), .ZN(n6842)
         );
  OAI21_X1 U9631 ( .B1(n12265), .B2(n7463), .A(n7462), .ZN(n14455) );
  AOI21_X1 U9632 ( .B1(n7462), .B2(n7463), .A(n6702), .ZN(n6854) );
  NAND2_X1 U9633 ( .A1(n12265), .A2(n7462), .ZN(n6855) );
  NAND2_X1 U9634 ( .A1(n12024), .A2(n6859), .ZN(n6856) );
  NAND2_X1 U9635 ( .A1(n6689), .A2(n6856), .ZN(n12169) );
  NOR2_X1 U9636 ( .A1(n6867), .A2(n6868), .ZN(n6866) );
  NAND2_X2 U9637 ( .A1(n10373), .A2(n14629), .ZN(n10563) );
  OR2_X1 U9638 ( .A1(n9820), .A2(n6871), .ZN(n6869) );
  NAND2_X2 U9639 ( .A1(n7322), .A2(n9891), .ZN(n14494) );
  NAND2_X1 U9640 ( .A1(n11842), .A2(n9750), .ZN(n9752) );
  NAND2_X1 U9641 ( .A1(n11291), .A2(n9748), .ZN(n6877) );
  NAND2_X1 U9642 ( .A1(n11760), .A2(n9743), .ZN(n6878) );
  NAND2_X1 U9643 ( .A1(n11187), .A2(n11188), .ZN(n6879) );
  NAND2_X1 U9644 ( .A1(n13727), .A2(n6667), .ZN(n6882) );
  NAND3_X1 U9645 ( .A1(n6882), .A2(n6880), .A3(n13679), .ZN(n13678) );
  NAND2_X1 U9646 ( .A1(n6888), .A2(n6887), .ZN(n9709) );
  NAND2_X2 U9647 ( .A1(n6888), .A2(n8153), .ZN(n13524) );
  NOR2_X2 U9648 ( .A1(n6889), .A2(n6594), .ZN(n6888) );
  NAND2_X1 U9649 ( .A1(n13640), .A2(n6899), .ZN(n6898) );
  NAND2_X1 U9650 ( .A1(n6891), .A2(n13640), .ZN(n6890) );
  NAND2_X1 U9651 ( .A1(n13640), .A2(n9782), .ZN(n9784) );
  NAND2_X1 U9652 ( .A1(n7592), .A2(n6898), .ZN(n13610) );
  INV_X1 U9653 ( .A(n9787), .ZN(n6894) );
  NAND3_X1 U9654 ( .A1(n7592), .A2(n6898), .A3(n9788), .ZN(n6895) );
  NAND2_X1 U9655 ( .A1(n12074), .A2(n6903), .ZN(n6901) );
  NAND2_X1 U9656 ( .A1(n6901), .A2(n6902), .ZN(n12125) );
  NAND2_X1 U9657 ( .A1(n7788), .A2(n7790), .ZN(n6909) );
  OAI211_X1 U9658 ( .C1(n6908), .C2(n9800), .A(n6906), .B(n9801), .ZN(P2_U3496) );
  OAI21_X1 U9659 ( .B1(n7614), .B2(n6562), .A(n7601), .ZN(n13761) );
  NAND2_X1 U9660 ( .A1(n6911), .A2(n6910), .ZN(n9769) );
  NAND2_X1 U9661 ( .A1(n7614), .A2(n7601), .ZN(n6911) );
  NAND2_X2 U9662 ( .A1(n13949), .A2(n7907), .ZN(n8138) );
  NAND2_X1 U9663 ( .A1(n6920), .A2(n6919), .ZN(n7868) );
  NAND2_X1 U9664 ( .A1(n11705), .A2(n6921), .ZN(n6920) );
  NAND2_X1 U9665 ( .A1(n13143), .A2(n9358), .ZN(n6929) );
  NAND3_X1 U9666 ( .A1(n9253), .A2(n9254), .A3(n15342), .ZN(n15340) );
  NAND2_X1 U9667 ( .A1(n14939), .A2(n11486), .ZN(n11490) );
  OAI21_X2 U9668 ( .B1(n6574), .B2(n6933), .A(n14025), .ZN(n14024) );
  OAI21_X2 U9669 ( .B1(n11647), .B2(n6941), .A(n6935), .ZN(n14944) );
  OAI21_X1 U9670 ( .B1(n11136), .B2(n12776), .A(n6952), .ZN(n6953) );
  NAND2_X4 U9671 ( .A1(n12753), .A2(n14399), .ZN(n12776) );
  OAI22_X2 U9672 ( .A1(n12666), .A2(n12665), .B1(n12664), .B2(n12663), .ZN(
        n14859) );
  OAI21_X2 U9673 ( .B1(n14954), .B2(n14957), .A(n14955), .ZN(n14876) );
  NAND3_X1 U9674 ( .A1(n7166), .A2(n6559), .A3(n7479), .ZN(n6955) );
  NAND2_X1 U9675 ( .A1(n11915), .A2(n7488), .ZN(n6959) );
  INV_X1 U9676 ( .A(n11915), .ZN(n6961) );
  NAND2_X1 U9677 ( .A1(n7243), .A2(n6961), .ZN(n7489) );
  INV_X1 U9678 ( .A(n6967), .ZN(n6965) );
  NAND3_X1 U9680 ( .A1(n6981), .A2(n6980), .A3(n7298), .ZN(n13622) );
  NAND2_X2 U9681 ( .A1(n7976), .A2(n7907), .ZN(n8137) );
  NOR2_X2 U9682 ( .A1(n9721), .A2(n7792), .ZN(n13739) );
  NAND2_X1 U9683 ( .A1(n8744), .A2(n8743), .ZN(n6988) );
  NAND2_X1 U9684 ( .A1(n8724), .A2(n8723), .ZN(n6989) );
  NAND2_X1 U9685 ( .A1(n6998), .A2(n7634), .ZN(n7000) );
  INV_X1 U9686 ( .A(n7001), .ZN(n13446) );
  NAND2_X1 U9687 ( .A1(n7986), .A2(n7966), .ZN(n8074) );
  NAND3_X1 U9688 ( .A1(n7986), .A2(n7966), .A3(n7967), .ZN(n8073) );
  INV_X1 U9689 ( .A(n11639), .ZN(n7003) );
  NAND2_X1 U9690 ( .A1(n7003), .A2(n7621), .ZN(n7002) );
  INV_X1 U9691 ( .A(n7621), .ZN(n7004) );
  NAND2_X1 U9692 ( .A1(n11928), .A2(n7621), .ZN(n11792) );
  NAND2_X1 U9693 ( .A1(n11639), .A2(n7005), .ZN(n11928) );
  NAND2_X1 U9694 ( .A1(n7009), .A2(n8872), .ZN(n8853) );
  NAND2_X1 U9695 ( .A1(n7009), .A2(n7008), .ZN(n8873) );
  NAND2_X1 U9696 ( .A1(n13455), .A2(n7010), .ZN(n7012) );
  INV_X1 U9697 ( .A(n8988), .ZN(n7016) );
  NOR2_X1 U9698 ( .A1(n7016), .A2(n8991), .ZN(n7017) );
  NAND2_X1 U9699 ( .A1(n8345), .A2(n6685), .ZN(n14843) );
  NAND3_X1 U9700 ( .A1(n8145), .A2(n7616), .A3(n8144), .ZN(n11398) );
  NAND2_X1 U9701 ( .A1(n9032), .A2(n14636), .ZN(n7018) );
  NAND2_X1 U9702 ( .A1(n7396), .A2(n7018), .ZN(n9058) );
  NAND2_X1 U9703 ( .A1(n7396), .A2(n9032), .ZN(n9043) );
  INV_X1 U9704 ( .A(n9247), .ZN(n7021) );
  NAND3_X1 U9705 ( .A1(n7024), .A2(n7023), .A3(n7022), .ZN(n7148) );
  NAND3_X1 U9706 ( .A1(n9247), .A2(n9371), .A3(n10405), .ZN(n7023) );
  NAND2_X1 U9707 ( .A1(n9194), .A2(n9245), .ZN(n9371) );
  NAND2_X1 U9708 ( .A1(n14922), .A2(n14923), .ZN(n14921) );
  NAND2_X2 U9709 ( .A1(n14918), .A2(n14724), .ZN(n14922) );
  NAND2_X1 U9710 ( .A1(n7029), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n7028) );
  OAI21_X2 U9711 ( .B1(n14727), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n14929), .ZN(
        n14790) );
  AOI21_X1 U9712 ( .B1(n14790), .B2(n14791), .A(n7651), .ZN(n7030) );
  NAND3_X1 U9713 ( .A1(n7034), .A2(n7035), .A3(n7031), .ZN(n7033) );
  AND2_X2 U9714 ( .A1(n7033), .A2(n7032), .ZN(n7652) );
  XNOR2_X1 U9715 ( .A(n7037), .B(n8147), .ZN(n10491) );
  NAND2_X1 U9716 ( .A1(n8236), .A2(n8021), .ZN(n7043) );
  OAI21_X2 U9717 ( .B1(n8236), .B2(n7046), .A(n7044), .ZN(n8253) );
  OAI21_X1 U9718 ( .B1(n10205), .B2(n7051), .A(n7049), .ZN(n10221) );
  NAND2_X1 U9719 ( .A1(n10195), .A2(n10194), .ZN(n10205) );
  INV_X1 U9720 ( .A(n7558), .ZN(n7052) );
  INV_X1 U9721 ( .A(n7053), .ZN(n7055) );
  NAND3_X1 U9722 ( .A1(n7226), .A2(n10297), .A3(n10305), .ZN(n7059) );
  INV_X1 U9723 ( .A(n10306), .ZN(n7060) );
  NAND2_X1 U9724 ( .A1(n7580), .A2(n7579), .ZN(n10107) );
  OAI211_X1 U9725 ( .C1(n7061), .C2(n6664), .A(n7117), .B(n6573), .ZN(n7579)
         );
  NAND3_X1 U9726 ( .A1(n8159), .A2(n8008), .A3(n8011), .ZN(n7064) );
  NAND3_X1 U9727 ( .A1(n7590), .A2(n7591), .A3(n7069), .ZN(n7068) );
  NAND2_X1 U9728 ( .A1(n7068), .A2(n7071), .ZN(n10190) );
  NAND2_X1 U9729 ( .A1(n7411), .A2(n11739), .ZN(n7199) );
  NAND2_X1 U9730 ( .A1(n7121), .A2(n6633), .ZN(n7176) );
  NAND3_X1 U9731 ( .A1(n7074), .A2(n7075), .A3(n11365), .ZN(n7073) );
  OR2_X1 U9732 ( .A1(n11386), .A2(n7073), .ZN(n15362) );
  INV_X1 U9733 ( .A(n12624), .ZN(n12626) );
  NAND2_X1 U9734 ( .A1(n12887), .A2(n7080), .ZN(n7079) );
  OAI211_X1 U9735 ( .C1(n12887), .C2(n7081), .A(n7079), .B(n12803), .ZN(
        P3_U3154) );
  NAND2_X1 U9736 ( .A1(n12887), .A2(n12888), .ZN(n12639) );
  OAI21_X1 U9737 ( .B1(n12427), .B2(n7089), .A(n7086), .ZN(n12518) );
  NAND2_X1 U9738 ( .A1(n7093), .A2(n7091), .ZN(n12813) );
  NAND2_X1 U9739 ( .A1(n7104), .A2(n7102), .ZN(n7101) );
  NAND2_X1 U9740 ( .A1(n12406), .A2(n7099), .ZN(n12407) );
  NAND2_X1 U9741 ( .A1(n7101), .A2(n7100), .ZN(n7099) );
  NAND2_X1 U9742 ( .A1(n7104), .A2(n7423), .ZN(n12332) );
  NOR2_X1 U9743 ( .A1(n11388), .A2(n11279), .ZN(n11385) );
  NAND2_X1 U9744 ( .A1(n7195), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7197) );
  NOR2_X1 U9745 ( .A1(n11856), .A2(n11862), .ZN(n11900) );
  OAI21_X1 U9746 ( .B1(n12611), .B2(n12610), .A(n12899), .ZN(n12612) );
  NAND2_X1 U9747 ( .A1(n9945), .A2(n9944), .ZN(n7550) );
  AOI21_X2 U9748 ( .B1(n10253), .B2(n10252), .A(n10251), .ZN(n10256) );
  OAI21_X1 U9749 ( .B1(n7213), .B2(n7214), .A(n10125), .ZN(n10149) );
  OAI21_X1 U9750 ( .B1(n7573), .B2(n7215), .A(n9989), .ZN(n10006) );
  NAND4_X2 U9751 ( .A1(n9862), .A2(n7693), .A3(n7691), .A4(n7692), .ZN(n14109)
         );
  INV_X1 U9752 ( .A(n12657), .ZN(n8652) );
  NAND2_X1 U9753 ( .A1(n11386), .A2(n9116), .ZN(n11271) );
  NAND2_X1 U9754 ( .A1(n7106), .A2(n6640), .ZN(n11393) );
  NAND2_X1 U9755 ( .A1(n11572), .A2(n11699), .ZN(n11739) );
  INV_X1 U9756 ( .A(n11741), .ZN(n7198) );
  NAND2_X1 U9757 ( .A1(n7238), .A2(n9162), .ZN(n10520) );
  OAI22_X1 U9758 ( .A1(n15362), .A2(n11571), .B1(n11271), .B2(n11383), .ZN(
        n11388) );
  NOR2_X1 U9759 ( .A1(n11385), .A2(n11280), .ZN(n15432) );
  NAND2_X1 U9760 ( .A1(n7521), .A2(n7523), .ZN(n7106) );
  NAND2_X1 U9761 ( .A1(n7522), .A2(n6781), .ZN(n7521) );
  NAND2_X1 U9762 ( .A1(n12804), .A2(n12872), .ZN(n12632) );
  NAND2_X1 U9763 ( .A1(n13013), .A2(n7670), .ZN(n7669) );
  NAND2_X1 U9764 ( .A1(n9772), .A2(n9771), .ZN(n13731) );
  NAND2_X1 U9765 ( .A1(n9769), .A2(n9768), .ZN(n13747) );
  NAND2_X1 U9766 ( .A1(n9741), .A2(n9740), .ZN(n11188) );
  OAI21_X1 U9767 ( .B1(n12239), .B2(n9760), .A(n9761), .ZN(n12450) );
  NOR2_X1 U9768 ( .A1(n7401), .A2(n6618), .ZN(n7399) );
  OAI211_X1 U9769 ( .C1(n12639), .C2(n7398), .A(n7397), .B(n12647), .ZN(
        P3_U3160) );
  XNOR2_X1 U9770 ( .A(n13070), .B(n12640), .ZN(n7410) );
  OAI21_X1 U9771 ( .B1(n9880), .B2(n9879), .A(n9878), .ZN(n9881) );
  NAND2_X1 U9772 ( .A1(n8873), .A2(n8872), .ZN(n8876) );
  NAND2_X1 U9773 ( .A1(n9376), .A2(n6662), .ZN(n7133) );
  OR2_X1 U9774 ( .A1(n10278), .A2(n11537), .ZN(n9915) );
  NAND2_X1 U9775 ( .A1(n7575), .A2(n9988), .ZN(n7574) );
  INV_X1 U9776 ( .A(n9974), .ZN(n7578) );
  NAND2_X1 U9777 ( .A1(n9913), .A2(n9914), .ZN(n7107) );
  AND2_X1 U9778 ( .A1(n9897), .A2(n9895), .ZN(n7110) );
  NAND2_X1 U9779 ( .A1(n7727), .A2(n14524), .ZN(n14603) );
  OR2_X1 U9780 ( .A1(n14279), .A2(n15002), .ZN(n7147) );
  NAND2_X1 U9781 ( .A1(n7355), .A2(n6682), .ZN(n14311) );
  NOR2_X1 U9782 ( .A1(n7357), .A2(n6612), .ZN(n7356) );
  NAND2_X1 U9783 ( .A1(n11592), .A2(n11591), .ZN(n11724) );
  NAND2_X1 U9784 ( .A1(n11205), .A2(n11221), .ZN(n11550) );
  INV_X1 U9785 ( .A(n7360), .ZN(n7357) );
  NAND2_X1 U9786 ( .A1(n11113), .A2(n7690), .ZN(n11316) );
  NAND2_X1 U9787 ( .A1(n7756), .A2(n7757), .ZN(n8046) );
  NAND2_X1 U9788 ( .A1(n6668), .A2(n6567), .ZN(n9697) );
  NOR2_X1 U9789 ( .A1(n9788), .A2(n9694), .ZN(n7112) );
  INV_X1 U9790 ( .A(n8349), .ZN(n7152) );
  NAND2_X1 U9791 ( .A1(n11237), .A2(n10237), .ZN(n7177) );
  NAND2_X1 U9792 ( .A1(n12611), .A2(n12610), .ZN(n7120) );
  NAND2_X1 U9793 ( .A1(n12612), .A2(n7120), .ZN(n12836) );
  INV_X1 U9794 ( .A(n15432), .ZN(n7121) );
  XNOR2_X2 U9795 ( .A(n7650), .B(n14793), .ZN(n14734) );
  NAND2_X1 U9796 ( .A1(n7239), .A2(n6716), .ZN(n12845) );
  NOR2_X1 U9797 ( .A1(n14931), .A2(n14930), .ZN(n14727) );
  OAI21_X1 U9798 ( .B1(n10771), .B2(n10770), .A(n10769), .ZN(n11100) );
  NOR2_X2 U9799 ( .A1(n10084), .A2(n7735), .ZN(n9820) );
  NAND3_X1 U9800 ( .A1(n7579), .A2(n7228), .A3(n7580), .ZN(n7582) );
  NOR2_X1 U9801 ( .A1(n14768), .A2(n14767), .ZN(n14766) );
  NAND2_X1 U9802 ( .A1(n15739), .A2(n15738), .ZN(n15737) );
  NOR2_X1 U9803 ( .A1(n14739), .A2(n14738), .ZN(n14737) );
  NAND2_X1 U9804 ( .A1(n6583), .A2(n14775), .ZN(n7222) );
  OAI21_X1 U9805 ( .B1(n10256), .B2(n10255), .A(n10254), .ZN(n10286) );
  OAI21_X1 U9806 ( .B1(n9716), .B2(n15252), .A(n12077), .ZN(n12092) );
  NAND2_X1 U9807 ( .A1(n11786), .A2(n11785), .ZN(n11784) );
  NAND2_X1 U9808 ( .A1(n12079), .A2(n12078), .ZN(n12077) );
  NAND2_X1 U9809 ( .A1(n11189), .A2(n9709), .ZN(n11762) );
  INV_X1 U9810 ( .A(n9739), .ZN(n11786) );
  NAND2_X1 U9811 ( .A1(n7891), .A2(n7892), .ZN(n13165) );
  NAND2_X1 U9812 ( .A1(n13235), .A2(n13234), .ZN(n13233) );
  NAND2_X1 U9813 ( .A1(n11190), .A2(n11191), .ZN(n11189) );
  OAI21_X1 U9814 ( .B1(n13091), .B2(n9071), .A(n9242), .ZN(n9087) );
  NOR3_X1 U9815 ( .A1(n9240), .A2(n9402), .A3(n9239), .ZN(n9241) );
  NAND2_X1 U9816 ( .A1(n7136), .A2(n8711), .ZN(n8724) );
  NAND2_X1 U9817 ( .A1(n8876), .A2(n8875), .ZN(n8888) );
  NAND2_X1 U9818 ( .A1(n8945), .A2(n8944), .ZN(n8958) );
  XNOR2_X1 U9819 ( .A(n7391), .B(n13033), .ZN(n9403) );
  NAND2_X1 U9820 ( .A1(n7133), .A2(n9377), .ZN(n9378) );
  NOR2_X1 U9821 ( .A1(n12991), .A2(n13003), .ZN(n13013) );
  OAI21_X1 U9822 ( .B1(n9379), .B2(n9378), .A(n9382), .ZN(n9404) );
  NAND2_X1 U9823 ( .A1(n7373), .A2(n7154), .ZN(n7136) );
  NAND2_X1 U9824 ( .A1(n14051), .A2(n14052), .ZN(n14050) );
  NAND2_X1 U9825 ( .A1(n14062), .A2(n14063), .ZN(n14061) );
  NAND2_X1 U9826 ( .A1(n7815), .A2(n7813), .ZN(n13997) );
  NOR2_X1 U9827 ( .A1(n12678), .A2(n12679), .ZN(n12683) );
  INV_X1 U9828 ( .A(n12108), .ZN(n12193) );
  NAND2_X1 U9829 ( .A1(n12108), .A2(n7137), .ZN(n12008) );
  NAND2_X1 U9830 ( .A1(n7138), .A2(n15310), .ZN(n7137) );
  INV_X1 U9831 ( .A(n12195), .ZN(n7138) );
  INV_X1 U9832 ( .A(n8633), .ZN(n8608) );
  NAND2_X1 U9833 ( .A1(n11627), .A2(n8194), .ZN(n11372) );
  INV_X1 U9834 ( .A(n7165), .ZN(n11371) );
  OAI21_X2 U9835 ( .B1(n13466), .B2(n13462), .A(n13463), .ZN(n13416) );
  NAND2_X1 U9836 ( .A1(n8072), .A2(n8071), .ZN(n8625) );
  NAND2_X1 U9837 ( .A1(n8190), .A2(n11617), .ZN(n11627) );
  OR2_X2 U9838 ( .A1(n12129), .A2(n12253), .ZN(n12249) );
  NAND2_X1 U9839 ( .A1(n7490), .A2(n12132), .ZN(n12129) );
  NAND2_X1 U9840 ( .A1(n7500), .A2(n7499), .ZN(n13732) );
  NAND2_X1 U9841 ( .A1(n13803), .A2(n13783), .ZN(n13780) );
  NOR2_X2 U9842 ( .A1(n13860), .A2(n13671), .ZN(n13662) );
  INV_X1 U9843 ( .A(n9426), .ZN(n9675) );
  NOR2_X2 U9844 ( .A1(n13646), .A2(n13849), .ZN(n7755) );
  AOI21_X1 U9845 ( .B1(n9976), .B2(n7576), .A(n7574), .ZN(n7573) );
  OAI21_X1 U9846 ( .B1(n9904), .B2(n9903), .A(n9902), .ZN(n9906) );
  INV_X1 U9847 ( .A(n8046), .ZN(n7149) );
  NAND2_X1 U9848 ( .A1(n9087), .A2(n9145), .ZN(n9196) );
  MUX2_X1 U9849 ( .A(P2_IR_REG_0__SCAN_IN), .B(n6742), .S(n8126), .Z(n9791) );
  NAND2_X1 U9850 ( .A1(n13403), .A2(n7150), .ZN(n13455) );
  INV_X1 U9851 ( .A(n12267), .ZN(n12265) );
  INV_X1 U9852 ( .A(n7323), .ZN(n7322) );
  NAND2_X1 U9853 ( .A1(n7153), .A2(n8779), .ZN(n8795) );
  NAND2_X1 U9854 ( .A1(n9030), .A2(n9029), .ZN(n9031) );
  NAND2_X1 U9855 ( .A1(n8777), .A2(n8776), .ZN(n7153) );
  NAND2_X1 U9856 ( .A1(n7376), .A2(n8684), .ZN(n7154) );
  NAND2_X1 U9857 ( .A1(n7157), .A2(n7155), .ZN(P1_U3214) );
  NAND2_X1 U9858 ( .A1(n13973), .A2(n14961), .ZN(n7157) );
  NAND2_X1 U9859 ( .A1(n14071), .A2(n12768), .ZN(n13971) );
  INV_X1 U9860 ( .A(n7728), .ZN(n7727) );
  NAND2_X1 U9861 ( .A1(n7726), .A2(n7725), .ZN(P1_U3555) );
  NAND2_X1 U9862 ( .A1(n7511), .A2(n7516), .ZN(n10378) );
  NAND2_X1 U9863 ( .A1(n13199), .A2(n9141), .ZN(n13182) );
  NAND2_X1 U9864 ( .A1(n7623), .A2(n7622), .ZN(n8571) );
  NOR2_X1 U9865 ( .A1(n11372), .A2(n11373), .ZN(n7165) );
  NAND2_X1 U9866 ( .A1(n8157), .A2(n8172), .ZN(n11525) );
  INV_X1 U9867 ( .A(n8152), .ZN(n7807) );
  NOR2_X1 U9868 ( .A1(n12965), .A2(n12964), .ZN(n12987) );
  NAND2_X1 U9869 ( .A1(n8986), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8989) );
  NAND2_X1 U9870 ( .A1(n8961), .A2(n8960), .ZN(n8978) );
  INV_X1 U9871 ( .A(n8683), .ZN(n7372) );
  INV_X1 U9872 ( .A(n8852), .ZN(n7167) );
  AOI21_X1 U9873 ( .B1(n7380), .B2(n8902), .A(n7379), .ZN(n7378) );
  NAND2_X1 U9874 ( .A1(n8958), .A2(n8957), .ZN(n8961) );
  NAND2_X1 U9875 ( .A1(n7936), .A2(n9405), .ZN(n9408) );
  AOI21_X1 U9876 ( .B1(n7376), .B2(n7375), .A(n7374), .ZN(n7373) );
  NAND2_X1 U9877 ( .A1(n7326), .A2(n7325), .ZN(P1_U3557) );
  NAND2_X1 U9878 ( .A1(n7868), .A2(n7866), .ZN(n15281) );
  OR2_X2 U9879 ( .A1(n6583), .A2(n14775), .ZN(n7657) );
  OAI21_X1 U9880 ( .B1(n11603), .B2(n7803), .A(n9753), .ZN(n12074) );
  NAND2_X1 U9881 ( .A1(n9752), .A2(n9751), .ZN(n11603) );
  NAND2_X1 U9882 ( .A1(n13050), .A2(n13049), .ZN(n7175) );
  XNOR2_X1 U9883 ( .A(n10895), .B(n10888), .ZN(n11090) );
  AOI21_X1 U9884 ( .B1(n10149), .B2(n12581), .A(n10148), .ZN(n10150) );
  NOR2_X1 U9885 ( .A1(n10231), .A2(n10230), .ZN(n7561) );
  AND2_X1 U9886 ( .A1(n7582), .A2(n10105), .ZN(n7214) );
  NAND2_X1 U9887 ( .A1(n13152), .A2(n9143), .ZN(n13155) );
  OAI211_X1 U9888 ( .C1(n7504), .C2(n7503), .A(n11423), .B(n7501), .ZN(n11422)
         );
  NAND2_X1 U9889 ( .A1(n7508), .A2(n7506), .ZN(n13069) );
  OAI21_X1 U9890 ( .B1(n10409), .B2(n15417), .A(n7178), .ZN(P3_U3488) );
  OAI21_X1 U9891 ( .B1(n10409), .B2(n15409), .A(n7180), .ZN(P3_U3456) );
  OAI21_X2 U9892 ( .B1(n13667), .B2(n13679), .A(n7782), .ZN(n13654) );
  NAND2_X1 U9893 ( .A1(n11293), .A2(n11294), .ZN(n11292) );
  NOR2_X1 U9894 ( .A1(n13751), .A2(n7315), .ZN(n9721) );
  AOI21_X1 U9895 ( .B1(n13622), .B2(n13628), .A(n7297), .ZN(n13605) );
  NAND2_X1 U9896 ( .A1(n13605), .A2(n9786), .ZN(n13608) );
  NAND2_X1 U9897 ( .A1(n12994), .A2(n12995), .ZN(n7236) );
  INV_X1 U9898 ( .A(n7593), .ZN(n7592) );
  INV_X1 U9899 ( .A(n11206), .ZN(n7195) );
  NAND2_X1 U9900 ( .A1(n10768), .A2(n6548), .ZN(n7186) );
  NAND2_X1 U9901 ( .A1(n7232), .A2(n6725), .ZN(n7675) );
  AOI21_X1 U9902 ( .B1(n7232), .B2(n7679), .A(n12977), .ZN(n12979) );
  NAND2_X1 U9903 ( .A1(n14927), .A2(n14925), .ZN(n14930) );
  OAI21_X1 U9904 ( .B1(n12450), .B2(n9762), .A(n9763), .ZN(n7614) );
  NAND2_X1 U9905 ( .A1(n9759), .A2(n9758), .ZN(n12239) );
  INV_X1 U9906 ( .A(n11111), .ZN(n9904) );
  AOI21_X1 U9907 ( .B1(n10250), .B2(n10249), .A(n10248), .ZN(n10251) );
  NAND2_X1 U9908 ( .A1(n10151), .A2(n7588), .ZN(n7585) );
  NAND3_X1 U9909 ( .A1(n6578), .A2(n7203), .A3(n15120), .ZN(n7202) );
  NOR2_X2 U9910 ( .A1(n12547), .A2(n8481), .ZN(n8499) );
  NAND2_X1 U9911 ( .A1(n7205), .A2(n7204), .ZN(n8072) );
  NAND2_X1 U9912 ( .A1(n8070), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n7205) );
  NAND2_X1 U9913 ( .A1(n11371), .A2(n8212), .ZN(n8234) );
  NAND2_X1 U9914 ( .A1(n10150), .A2(n7588), .ZN(n7584) );
  NOR2_X1 U9915 ( .A1(n10314), .A2(n10283), .ZN(n9902) );
  OAI21_X1 U9916 ( .B1(n14235), .B2(n14640), .A(n10709), .ZN(n9845) );
  NAND2_X1 U9917 ( .A1(n9964), .A2(n9963), .ZN(n9976) );
  INV_X1 U9918 ( .A(n7209), .ZN(n12011) );
  NAND2_X1 U9919 ( .A1(n7209), .A2(n6619), .ZN(n7208) );
  OAI21_X1 U9920 ( .B1(n10265), .B2(n10487), .A(n9892), .ZN(n7323) );
  NOR2_X1 U9921 ( .A1(n9820), .A2(n7211), .ZN(n7210) );
  NAND2_X1 U9922 ( .A1(n10123), .A2(n10122), .ZN(n7213) );
  OAI21_X1 U9923 ( .B1(n9976), .B2(n6605), .A(n7217), .ZN(n9989) );
  OAI21_X1 U9924 ( .B1(n10235), .B2(n10234), .A(n10233), .ZN(n10236) );
  NAND2_X1 U9925 ( .A1(n14928), .A2(n15165), .ZN(n14925) );
  XNOR2_X1 U9926 ( .A(n14710), .B(n7248), .ZN(n14770) );
  NAND2_X1 U9927 ( .A1(n9404), .A2(n9410), .ZN(n9405) );
  AOI21_X2 U9928 ( .B1(n8214), .B2(n8020), .A(n7941), .ZN(n8236) );
  NAND2_X1 U9929 ( .A1(n13416), .A2(n13415), .ZN(n13414) );
  NAND2_X1 U9930 ( .A1(n8571), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7987) );
  NAND2_X1 U9931 ( .A1(n9728), .A2(n7783), .ZN(n13667) );
  OAI21_X1 U9932 ( .B1(n10205), .B2(n6615), .A(n7227), .ZN(n10220) );
  INV_X1 U9933 ( .A(n10093), .ZN(n7581) );
  NAND2_X1 U9934 ( .A1(n10235), .A2(n10234), .ZN(n7560) );
  NAND2_X1 U9935 ( .A1(n10236), .A2(n7560), .ZN(n10250) );
  OR2_X1 U9936 ( .A1(n9149), .A2(n8660), .ZN(n9150) );
  NAND3_X1 U9937 ( .A1(n8706), .A2(n8704), .A3(n8705), .ZN(n7229) );
  INV_X1 U9938 ( .A(n11271), .ZN(n15355) );
  AOI21_X2 U9939 ( .B1(n10917), .B2(n10916), .A(n10915), .ZN(n11067) );
  OAI21_X1 U9940 ( .B1(n11205), .B2(n11221), .A(n11550), .ZN(n11206) );
  NOR2_X1 U9941 ( .A1(n10741), .A2(n10740), .ZN(n10887) );
  NAND2_X1 U9942 ( .A1(n9154), .A2(n12346), .ZN(n7238) );
  NAND2_X1 U9943 ( .A1(n12836), .A2(n12835), .ZN(n7239) );
  INV_X1 U9944 ( .A(n8385), .ZN(n7648) );
  NAND2_X2 U9945 ( .A1(n8291), .A2(n8290), .ZN(n8306) );
  NOR2_X1 U9946 ( .A1(n12626), .A2(n12625), .ZN(n12627) );
  XNOR2_X1 U9947 ( .A(n12960), .B(n12977), .ZN(n12942) );
  NAND2_X2 U9948 ( .A1(n7976), .A2(n7975), .ZN(n8139) );
  AND2_X1 U9949 ( .A1(n9483), .A2(n7255), .ZN(n7254) );
  NAND3_X1 U9950 ( .A1(n7986), .A2(n6693), .A3(n7966), .ZN(n7972) );
  NOR2_X1 U9951 ( .A1(n7256), .A2(n7260), .ZN(n7259) );
  NAND3_X1 U9952 ( .A1(n7261), .A2(n7259), .A3(n7257), .ZN(n9449) );
  NAND3_X1 U9953 ( .A1(n7948), .A2(n9439), .A3(n7258), .ZN(n7257) );
  NAND3_X1 U9954 ( .A1(n7948), .A2(n7262), .A3(n9439), .ZN(n7261) );
  NAND3_X1 U9955 ( .A1(n9504), .A2(n6694), .A3(n9503), .ZN(n7263) );
  NAND2_X1 U9956 ( .A1(n7263), .A2(n7264), .ZN(n7926) );
  INV_X1 U9957 ( .A(n9508), .ZN(n7267) );
  NAND2_X1 U9958 ( .A1(n7609), .A2(n8285), .ZN(n8122) );
  AND2_X1 U9959 ( .A1(n7609), .A2(n13814), .ZN(n7268) );
  AND2_X1 U9960 ( .A1(n7609), .A2(n13816), .ZN(n7269) );
  INV_X1 U9961 ( .A(n7609), .ZN(n7272) );
  AOI21_X1 U9962 ( .B1(n15113), .B2(n7609), .A(n6734), .ZN(n11380) );
  AOI21_X1 U9963 ( .B1(n15115), .B2(n7609), .A(n6739), .ZN(n11417) );
  NAND2_X1 U9964 ( .A1(n9646), .A2(n9658), .ZN(n7273) );
  NAND2_X1 U9965 ( .A1(n9491), .A2(n6561), .ZN(n7275) );
  AOI21_X1 U9966 ( .B1(n6561), .B2(n7278), .A(n6663), .ZN(n7274) );
  OAI22_X1 U9967 ( .A1(n9556), .A2(n7280), .B1(n9554), .B2(n9555), .ZN(n9561)
         );
  NOR2_X1 U9968 ( .A1(n9561), .A2(n9560), .ZN(n9562) );
  NAND2_X1 U9969 ( .A1(n9570), .A2(n7284), .ZN(n7283) );
  NAND2_X1 U9970 ( .A1(n7283), .A2(n7287), .ZN(n9573) );
  AOI21_X1 U9971 ( .B1(n7293), .B2(n7292), .A(n9571), .ZN(n7291) );
  INV_X1 U9972 ( .A(n9572), .ZN(n7295) );
  MUX2_X1 U9973 ( .A(n10493), .B(n10507), .S(n8013), .Z(n8005) );
  NAND2_X1 U9974 ( .A1(n8001), .A2(n8131), .ZN(n7300) );
  XNOR2_X1 U9975 ( .A(n8002), .B(n7741), .ZN(n8131) );
  NOR2_X2 U9976 ( .A1(n14893), .A2(n14892), .ZN(n14894) );
  NAND4_X1 U9977 ( .A1(n14801), .A2(n7739), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7341) );
  NAND4_X1 U9978 ( .A1(n7994), .A2(n14240), .A3(n7993), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7342) );
  NAND2_X1 U9979 ( .A1(n8253), .A2(n7344), .ZN(n7343) );
  NAND2_X1 U9980 ( .A1(n7343), .A2(n7346), .ZN(n8291) );
  INV_X1 U9981 ( .A(n8028), .ZN(n7348) );
  NAND2_X1 U9982 ( .A1(n8306), .A2(n7352), .ZN(n7350) );
  NAND2_X1 U9983 ( .A1(n7350), .A2(n7351), .ZN(n7756) );
  NAND2_X1 U9984 ( .A1(n7698), .A2(n7356), .ZN(n7355) );
  NAND3_X1 U9985 ( .A1(n7363), .A2(n12597), .A3(n7362), .ZN(n14256) );
  NAND2_X1 U9986 ( .A1(n7365), .A2(n7366), .ZN(n7370) );
  INV_X1 U9987 ( .A(n7370), .ZN(n14276) );
  OAI21_X1 U9988 ( .B1(n8684), .B2(n7375), .A(n7376), .ZN(n8710) );
  NAND2_X1 U9989 ( .A1(n8888), .A2(n7380), .ZN(n7377) );
  NAND2_X1 U9990 ( .A1(n7377), .A2(n7378), .ZN(n8923) );
  NAND3_X1 U9991 ( .A1(n9382), .A2(n7393), .A3(n7392), .ZN(n7391) );
  NAND2_X1 U9992 ( .A1(n12853), .A2(n7417), .ZN(n7415) );
  NAND2_X2 U9993 ( .A1(n7415), .A2(n7414), .ZN(n12887) );
  INV_X1 U9994 ( .A(n15001), .ZN(n7431) );
  NAND2_X1 U9995 ( .A1(n11583), .A2(n11588), .ZN(n7435) );
  INV_X1 U9996 ( .A(n12598), .ZN(n12596) );
  AOI21_X1 U9997 ( .B1(n14254), .B2(n6684), .A(n6576), .ZN(n7447) );
  OAI21_X1 U9998 ( .B1(n14515), .B2(n7452), .A(n7450), .ZN(P1_U3525) );
  INV_X1 U9999 ( .A(n14890), .ZN(n7471) );
  AND2_X1 U10000 ( .A1(n11778), .A2(n11194), .ZN(n11767) );
  MUX2_X1 U10001 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8773), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n8774) );
  MUX2_X1 U10002 ( .A(n8789), .B(P3_IR_REG_31__SCAN_IN), .S(n8791), .Z(n8793)
         );
  MUX2_X1 U10003 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8928), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n8930) );
  NAND2_X1 U10004 ( .A1(n6556), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7483) );
  INV_X1 U10005 ( .A(n7494), .ZN(n7490) );
  NAND2_X1 U10006 ( .A1(n7491), .A2(n11849), .ZN(n7494) );
  NOR2_X1 U10007 ( .A1(n15252), .A2(n11611), .ZN(n7493) );
  NAND2_X1 U10008 ( .A1(n8074), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8075) );
  NOR2_X2 U10009 ( .A1(n8150), .A2(n7957), .ZN(n7966) );
  NAND2_X1 U10010 ( .A1(n7755), .A2(n6575), .ZN(n7752) );
  NAND2_X1 U10011 ( .A1(n7755), .A2(n6691), .ZN(n13600) );
  NAND2_X1 U10012 ( .A1(n7755), .A2(n7754), .ZN(n13616) );
  INV_X1 U10013 ( .A(n7752), .ZN(n13601) );
  NOR2_X2 U10014 ( .A1(n13765), .A2(n13893), .ZN(n7500) );
  INV_X1 U10015 ( .A(n9119), .ZN(n7502) );
  NAND2_X1 U10016 ( .A1(n7502), .A2(n9120), .ZN(n7501) );
  INV_X1 U10017 ( .A(n9120), .ZN(n7503) );
  NAND2_X1 U10018 ( .A1(n11995), .A2(n9120), .ZN(n11424) );
  NAND2_X1 U10019 ( .A1(n7504), .A2(n9119), .ZN(n11995) );
  NAND2_X1 U10020 ( .A1(n13100), .A2(n7509), .ZN(n7508) );
  NAND2_X1 U10021 ( .A1(n13100), .A2(n7517), .ZN(n13088) );
  NOR2_X1 U10022 ( .A1(n13337), .A2(n13089), .ZN(n7518) );
  NAND2_X1 U10023 ( .A1(n13140), .A2(n7540), .ZN(n7539) );
  NAND2_X1 U10024 ( .A1(n9140), .A2(n7548), .ZN(n13199) );
  NAND2_X1 U10025 ( .A1(n7550), .A2(n9960), .ZN(n9962) );
  NAND2_X1 U10026 ( .A1(n7552), .A2(n7551), .ZN(n9964) );
  INV_X1 U10027 ( .A(n9960), .ZN(n7551) );
  NAND3_X1 U10028 ( .A1(n7554), .A2(n9939), .A3(n7553), .ZN(n9941) );
  INV_X1 U10029 ( .A(n12259), .ZN(n7583) );
  NAND2_X1 U10030 ( .A1(n9839), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9841) );
  AND2_X1 U10031 ( .A1(n10128), .A2(n9839), .ZN(n14222) );
  NAND2_X1 U10032 ( .A1(n10151), .A2(n10154), .ZN(n7587) );
  NAND2_X1 U10033 ( .A1(n10150), .A2(n10154), .ZN(n7586) );
  NAND3_X1 U10034 ( .A1(n7585), .A2(n7584), .A3(n10164), .ZN(n7591) );
  NAND3_X1 U10035 ( .A1(n7587), .A2(n7586), .A3(n10165), .ZN(n7590) );
  NAND3_X1 U10036 ( .A1(n13949), .A2(n7975), .A3(P2_REG0_REG_1__SCAN_IN), .ZN(
        n8115) );
  NAND2_X1 U10037 ( .A1(n6552), .A2(n7609), .ZN(n9417) );
  NAND2_X1 U10038 ( .A1(n7612), .A2(n7611), .ZN(n9738) );
  INV_X1 U10039 ( .A(n12065), .ZN(n7611) );
  INV_X1 U10040 ( .A(n9705), .ZN(n7612) );
  XNOR2_X1 U10041 ( .A(n9705), .B(n9426), .ZN(n12064) );
  XNOR2_X1 U10042 ( .A(n9705), .B(n12065), .ZN(n15218) );
  NAND4_X1 U10043 ( .A1(n9678), .A2(n11191), .A3(n9705), .A4(n11786), .ZN(
        n9681) );
  NAND2_X4 U10044 ( .A1(n8659), .A2(n8658), .ZN(n12946) );
  INV_X1 U10045 ( .A(n8680), .ZN(n7688) );
  NOR2_X1 U10046 ( .A1(n10746), .A2(n10963), .ZN(n10748) );
  OR2_X2 U10047 ( .A1(n14381), .A2(n14395), .ZN(n14376) );
  NOR2_X4 U10048 ( .A1(n14482), .A2(n14591), .ZN(n14467) );
  NOR2_X2 U10049 ( .A1(n15012), .A2(n11719), .ZN(n14994) );
  NAND2_X1 U10050 ( .A1(n7945), .A2(n12592), .ZN(n14308) );
  NAND2_X1 U10051 ( .A1(n12264), .A2(n12263), .ZN(n12267) );
  NAND2_X2 U10052 ( .A1(n15256), .A2(n11758), .ZN(n8134) );
  OAI21_X2 U10053 ( .B1(n11444), .B2(n6613), .A(n7617), .ZN(n11639) );
  AND2_X1 U10054 ( .A1(n7618), .A2(n11634), .ZN(n7617) );
  OR2_X1 U10055 ( .A1(n8247), .A2(n6613), .ZN(n7618) );
  INV_X1 U10056 ( .A(n7988), .ZN(n7623) );
  NAND3_X1 U10057 ( .A1(n7986), .A2(n7991), .A3(n8178), .ZN(n7988) );
  INV_X1 U10058 ( .A(n8561), .ZN(n7630) );
  NAND2_X1 U10059 ( .A1(n8438), .A2(n8439), .ZN(n7638) );
  OR2_X1 U10060 ( .A1(n14775), .A2(n14773), .ZN(n7658) );
  INV_X1 U10061 ( .A(n7659), .ZN(n14771) );
  NOR2_X2 U10062 ( .A1(n15746), .A2(n14688), .ZN(n14739) );
  NAND3_X1 U10063 ( .A1(n7671), .A2(n7669), .A3(n7668), .ZN(n7667) );
  INV_X1 U10064 ( .A(n13038), .ZN(n7673) );
  NAND3_X1 U10065 ( .A1(n7675), .A2(n7676), .A3(n7674), .ZN(n12955) );
  INV_X1 U10066 ( .A(n7678), .ZN(n12978) );
  INV_X1 U10067 ( .A(n10960), .ZN(n7682) );
  INV_X1 U10068 ( .A(n7690), .ZN(n11108) );
  OAI21_X1 U10069 ( .B1(n11113), .B2(n7690), .A(n11316), .ZN(n11116) );
  NAND2_X1 U10070 ( .A1(n14456), .A2(n7694), .ZN(n14450) );
  INV_X1 U10071 ( .A(n14358), .ZN(n7703) );
  NOR2_X1 U10072 ( .A1(n14060), .A2(n14095), .ZN(n7705) );
  NAND2_X1 U10073 ( .A1(n11586), .A2(n6681), .ZN(n7709) );
  NAND2_X1 U10074 ( .A1(n14883), .A2(n7714), .ZN(n7713) );
  AOI21_X1 U10075 ( .B1(n7714), .B2(n7717), .A(n7712), .ZN(n7711) );
  INV_X1 U10076 ( .A(n7724), .ZN(n11939) );
  NAND2_X1 U10077 ( .A1(n9837), .A2(n7734), .ZN(n9822) );
  NAND4_X1 U10078 ( .A1(n10364), .A2(n9836), .A3(n7737), .A4(n9815), .ZN(n7735) );
  NAND3_X1 U10079 ( .A1(n10364), .A2(n9836), .A3(n9815), .ZN(n7738) );
  NAND2_X1 U10080 ( .A1(n8004), .A2(n10495), .ZN(n7742) );
  NAND2_X1 U10081 ( .A1(n7997), .A2(n10481), .ZN(n7743) );
  NAND2_X1 U10082 ( .A1(n8089), .A2(n7750), .ZN(n7746) );
  NAND2_X1 U10083 ( .A1(n8058), .A2(n7746), .ZN(n10186) );
  NAND2_X1 U10084 ( .A1(n7791), .A2(n6737), .ZN(n7785) );
  OAI211_X1 U10085 ( .C1(n9796), .C2(n15277), .A(n7786), .B(n7785), .ZN(
        P2_U3528) );
  INV_X1 U10086 ( .A(n9736), .ZN(n7790) );
  NOR2_X1 U10087 ( .A1(n12132), .A2(n15112), .ZN(n7799) );
  NAND2_X1 U10088 ( .A1(n7808), .A2(n7809), .ZN(n12783) );
  NAND2_X1 U10089 ( .A1(n14072), .A2(n7810), .ZN(n7808) );
  NAND2_X1 U10090 ( .A1(n14061), .A2(n7816), .ZN(n7815) );
  INV_X1 U10091 ( .A(n7830), .ZN(n14082) );
  INV_X1 U10092 ( .A(n12683), .ZN(n7829) );
  NAND2_X1 U10093 ( .A1(n7855), .A2(n11666), .ZN(n11672) );
  INV_X1 U10094 ( .A(n11667), .ZN(n7856) );
  INV_X1 U10095 ( .A(n9839), .ZN(n7857) );
  NAND2_X1 U10096 ( .A1(n7857), .A2(n7858), .ZN(n10358) );
  NAND3_X1 U10097 ( .A1(n9843), .A2(n9840), .A3(n7860), .ZN(n7859) );
  INV_X1 U10098 ( .A(n11689), .ZN(n7863) );
  NAND3_X1 U10099 ( .A1(n7862), .A2(n7861), .A3(n11706), .ZN(n11705) );
  NAND2_X1 U10100 ( .A1(n6801), .A2(n9278), .ZN(n7861) );
  NAND2_X1 U10101 ( .A1(n11689), .A2(n9278), .ZN(n7862) );
  NAND2_X1 U10102 ( .A1(n11692), .A2(n9278), .ZN(n11707) );
  NAND2_X1 U10103 ( .A1(n7872), .A2(n7873), .ZN(n13235) );
  NAND3_X1 U10104 ( .A1(n8643), .A2(n8642), .A3(n6584), .ZN(n9097) );
  NAND2_X1 U10105 ( .A1(n13181), .A2(n7894), .ZN(n7891) );
  INV_X1 U10106 ( .A(n9528), .ZN(n7910) );
  INV_X1 U10107 ( .A(n7911), .ZN(n9476) );
  AOI21_X1 U10108 ( .B1(n9466), .B2(n7913), .A(n7912), .ZN(n7911) );
  NOR2_X1 U10109 ( .A1(n9471), .A2(n7914), .ZN(n7912) );
  AOI21_X1 U10110 ( .B1(n9471), .B2(n7914), .A(n6660), .ZN(n7913) );
  INV_X1 U10111 ( .A(n9470), .ZN(n7914) );
  NAND2_X1 U10112 ( .A1(n9543), .A2(n7918), .ZN(n7917) );
  INV_X1 U10113 ( .A(n9542), .ZN(n7920) );
  OAI21_X1 U10114 ( .B1(n7932), .B2(n9563), .A(n7933), .ZN(n9570) );
  OR2_X1 U10115 ( .A1(n9562), .A2(n7934), .ZN(n7932) );
  INV_X1 U10116 ( .A(n9567), .ZN(n7935) );
  NAND2_X1 U10117 ( .A1(n14984), .A2(n11726), .ZN(n11729) );
  NAND2_X1 U10118 ( .A1(n12596), .A2(n12595), .ZN(n14254) );
  OAI21_X1 U10119 ( .B1(n9409), .B2(n9408), .A(n9407), .ZN(n9415) );
  INV_X1 U10120 ( .A(n9893), .ZN(n10257) );
  INV_X1 U10121 ( .A(n12607), .ZN(n9795) );
  AND2_X1 U10122 ( .A1(n13198), .A2(n13197), .ZN(n13299) );
  INV_X1 U10123 ( .A(n11490), .ZN(n11493) );
  OR2_X1 U10124 ( .A1(n9403), .A2(n10396), .ZN(n7936) );
  OR2_X1 U10125 ( .A1(n15409), .A2(n15353), .ZN(n13376) );
  INV_X1 U10126 ( .A(n13376), .ZN(n10411) );
  INV_X2 U10127 ( .A(n15372), .ZN(n13255) );
  NAND2_X2 U10128 ( .A1(n11363), .A2(n15326), .ZN(n15372) );
  AND2_X1 U10129 ( .A1(n14952), .A2(n12302), .ZN(n7937) );
  INV_X1 U10130 ( .A(n8080), .ZN(n12053) );
  NAND2_X2 U10131 ( .A1(n11757), .A2(n13784), .ZN(n13770) );
  INV_X1 U10132 ( .A(n15270), .ZN(n9800) );
  AND2_X1 U10133 ( .A1(n13085), .A2(n15381), .ZN(n7938) );
  AND2_X1 U10134 ( .A1(n14110), .A2(n11143), .ZN(n7939) );
  INV_X1 U10135 ( .A(n13967), .ZN(n13951) );
  INV_X1 U10136 ( .A(n13951), .ZN(n12649) );
  NAND2_X1 U10137 ( .A1(n9638), .A2(n9637), .ZN(n7940) );
  NOR2_X1 U10138 ( .A1(n8019), .A2(n8018), .ZN(n7941) );
  AND2_X1 U10139 ( .A1(n11225), .A2(n11065), .ZN(n7942) );
  INV_X1 U10140 ( .A(n14814), .ZN(n8831) );
  INV_X1 U10141 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8375) );
  INV_X1 U10142 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7994) );
  INV_X1 U10143 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10037) );
  INV_X1 U10144 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9977) );
  INV_X1 U10145 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13943) );
  INV_X1 U10146 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10065) );
  INV_X1 U10147 ( .A(n15366), .ZN(n10380) );
  NAND2_X1 U10148 ( .A1(n9648), .A2(n9647), .ZN(n7943) );
  NOR2_X1 U10149 ( .A1(n14513), .A2(n14512), .ZN(n7944) );
  INV_X1 U10150 ( .A(n14310), .ZN(n12592) );
  AND2_X1 U10151 ( .A1(n10166), .A2(n14001), .ZN(n7947) );
  OR2_X1 U10152 ( .A1(n9438), .A2(n9437), .ZN(n7948) );
  AND2_X1 U10153 ( .A1(n6548), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7949) );
  AND2_X1 U10154 ( .A1(n10916), .A2(n10883), .ZN(n7950) );
  INV_X1 U10155 ( .A(SI_26_), .ZN(n12455) );
  INV_X1 U10156 ( .A(n11975), .ZN(n9407) );
  AND2_X1 U10157 ( .A1(n15256), .A2(n15255), .ZN(n15249) );
  INV_X1 U10158 ( .A(n15249), .ZN(n9794) );
  AND2_X1 U10159 ( .A1(n9653), .A2(n8105), .ZN(n9420) );
  NAND2_X1 U10160 ( .A1(n9426), .A2(n6552), .ZN(n9427) );
  NAND2_X1 U10161 ( .A1(n9430), .A2(n9429), .ZN(n9431) );
  NAND2_X1 U10162 ( .A1(n11111), .A2(n10283), .ZN(n9905) );
  OAI21_X1 U10163 ( .B1(n9711), .B2(n9653), .A(n9452), .ZN(n9453) );
  OAI21_X1 U10164 ( .B1(n11451), .B2(n9653), .A(n9469), .ZN(n9470) );
  AOI21_X1 U10165 ( .B1(n9476), .B2(n9475), .A(n9474), .ZN(n9478) );
  OAI21_X1 U10166 ( .B1(n9716), .B2(n9653), .A(n9481), .ZN(n9482) );
  NAND2_X1 U10167 ( .A1(n9515), .A2(n9514), .ZN(n9521) );
  NAND2_X1 U10168 ( .A1(n10193), .A2(n10192), .ZN(n10194) );
  INV_X1 U10169 ( .A(n14750), .ZN(n10888) );
  INV_X1 U10170 ( .A(n9049), .ZN(n9048) );
  NAND2_X1 U10171 ( .A1(n9028), .A2(n9027), .ZN(n9030) );
  INV_X1 U10172 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8933) );
  INV_X1 U10173 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8782) );
  INV_X1 U10174 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n8796) );
  INV_X1 U10175 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8393) );
  NAND2_X1 U10176 ( .A1(n13870), .A2(n13398), .ZN(n9727) );
  INV_X1 U10177 ( .A(n11673), .ZN(n11674) );
  INV_X1 U10178 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9928) );
  INV_X1 U10179 ( .A(n11491), .ZN(n11492) );
  INV_X1 U10180 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14043) );
  INV_X1 U10181 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n15586) );
  INV_X1 U10182 ( .A(SI_15_), .ZN(n8039) );
  INV_X1 U10183 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9802) );
  INV_X1 U10184 ( .A(n8972), .ZN(n8971) );
  INV_X1 U10185 ( .A(n9008), .ZN(n9010) );
  INV_X1 U10186 ( .A(n11542), .ZN(n11274) );
  OR2_X1 U10187 ( .A1(n9078), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9107) );
  INV_X1 U10188 ( .A(n10377), .ZN(n9145) );
  OR2_X1 U10189 ( .A1(n8881), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8896) );
  NAND2_X1 U10190 ( .A1(n8841), .A2(n12385), .ZN(n8866) );
  OR2_X1 U10191 ( .A1(n8801), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8817) );
  OR2_X1 U10192 ( .A1(n10520), .A2(n9177), .ZN(n10399) );
  AND2_X1 U10193 ( .A1(n8941), .A2(n8924), .ZN(n8925) );
  INV_X1 U10194 ( .A(n8126), .ZN(n8237) );
  INV_X1 U10195 ( .A(n8490), .ZN(n8508) );
  INV_X1 U10196 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8440) );
  OR2_X1 U10197 ( .A1(n8138), .A2(n8114), .ZN(n8116) );
  NAND2_X1 U10198 ( .A1(n7497), .A2(n13684), .ZN(n9726) );
  INV_X1 U10199 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8081) );
  NAND2_X1 U10200 ( .A1(n11493), .A2(n11492), .ZN(n11531) );
  NOR2_X1 U10201 ( .A1(n10293), .A2(n10296), .ZN(n10297) );
  INV_X1 U10202 ( .A(n10210), .ZN(n10223) );
  OR2_X1 U10203 ( .A1(n10141), .A2(n9827), .ZN(n10155) );
  OR2_X1 U10204 ( .A1(n11008), .A2(n11007), .ZN(n11025) );
  INV_X1 U10205 ( .A(n14640), .ZN(n11082) );
  AND2_X1 U10206 ( .A1(n8305), .A2(n8308), .ZN(n8034) );
  NAND2_X1 U10207 ( .A1(n8004), .A2(n10488), .ZN(n7995) );
  NOR2_X1 U10208 ( .A1(n14709), .A2(n14708), .ZN(n14654) );
  NAND2_X1 U10209 ( .A1(n8971), .A2(n8970), .ZN(n8981) );
  OR2_X1 U10210 ( .A1(n8981), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9008) );
  INV_X1 U10211 ( .A(n13141), .ZN(n12872) );
  NAND2_X1 U10212 ( .A1(n10948), .A2(n11283), .ZN(n12891) );
  INV_X1 U10213 ( .A(n11683), .ZN(n9411) );
  AND2_X1 U10214 ( .A1(n9070), .A2(n9069), .ZN(n12830) );
  AND3_X1 U10215 ( .A1(n8985), .A2(n8984), .A3(n8983), .ZN(n13156) );
  INV_X1 U10216 ( .A(n11219), .ZN(n11221) );
  OR2_X1 U10217 ( .A1(n10752), .A2(n10734), .ZN(n10742) );
  NOR2_X1 U10218 ( .A1(n10384), .A2(n10383), .ZN(n10385) );
  INV_X1 U10219 ( .A(n12899), .ZN(n13231) );
  AND2_X1 U10220 ( .A1(n8764), .A2(n11556), .ZN(n8783) );
  INV_X1 U10221 ( .A(n13379), .ZN(n10401) );
  OR2_X1 U10222 ( .A1(n8722), .A2(n12653), .ZN(n9193) );
  AND2_X1 U10223 ( .A1(n9104), .A2(n9179), .ZN(n13107) );
  AND2_X1 U10224 ( .A1(n9380), .A2(n10397), .ZN(n15366) );
  OAI21_X1 U10225 ( .B1(n9735), .B2(n13690), .A(n15120), .ZN(n8609) );
  AND2_X1 U10226 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n7978) );
  NAND2_X1 U10227 ( .A1(n9662), .A2(n9698), .ZN(n9663) );
  AND2_X1 U10228 ( .A1(n8473), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8489) );
  AND2_X1 U10229 ( .A1(n8458), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8473) );
  NAND2_X1 U10230 ( .A1(n13770), .A2(n11769), .ZN(n13828) );
  INV_X1 U10231 ( .A(n13677), .ZN(n13865) );
  INV_X1 U10232 ( .A(n13819), .ZN(n13799) );
  AND2_X1 U10233 ( .A1(n8585), .A2(n8587), .ZN(n8574) );
  INV_X1 U10234 ( .A(n14936), .ZN(n11485) );
  INV_X1 U10235 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14001) );
  INV_X1 U10236 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10794) );
  INV_X1 U10237 ( .A(n14359), .ZN(n14396) );
  NAND2_X1 U10238 ( .A1(n10115), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10141) );
  OR2_X1 U10239 ( .A1(n11156), .A2(n11155), .ZN(n11501) );
  INV_X1 U10240 ( .A(n10351), .ZN(n10352) );
  OR2_X1 U10241 ( .A1(n10278), .A2(n14283), .ZN(n10245) );
  NOR2_X1 U10242 ( .A1(n10166), .A2(n14001), .ZN(n10176) );
  INV_X1 U10243 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14646) );
  INV_X1 U10244 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n11678) );
  OR2_X1 U10245 ( .A1(n11151), .A2(n10373), .ZN(n14462) );
  NAND2_X1 U10246 ( .A1(n11131), .A2(n11311), .ZN(n11303) );
  NOR2_X1 U10247 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n14696), .ZN(n14649) );
  OAI21_X1 U10248 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n14667), .A(n14666), 
        .ZN(n14674) );
  INV_X1 U10249 ( .A(n15434), .ZN(n12861) );
  OR2_X1 U10250 ( .A1(n13054), .A2(n8700), .ZN(n9229) );
  AND3_X1 U10251 ( .A1(n9014), .A2(n9013), .A3(n9012), .ZN(n13157) );
  INV_X1 U10252 ( .A(n13051), .ZN(n12916) );
  INV_X1 U10253 ( .A(n10742), .ZN(n10738) );
  INV_X1 U10254 ( .A(n13033), .ZN(n13042) );
  INV_X1 U10255 ( .A(n15298), .ZN(n15360) );
  NOR2_X1 U10256 ( .A1(n11363), .A2(n11362), .ZN(n15336) );
  INV_X1 U10257 ( .A(n15326), .ZN(n15369) );
  INV_X1 U10258 ( .A(n13317), .ZN(n9187) );
  INV_X1 U10259 ( .A(n15353), .ZN(n13290) );
  AND2_X1 U10260 ( .A1(n10394), .A2(n9178), .ZN(n11359) );
  NAND2_X1 U10261 ( .A1(n13107), .A2(n10388), .ZN(n15405) );
  OR2_X1 U10262 ( .A1(n10520), .A2(P3_D_REG_1__SCAN_IN), .ZN(n9156) );
  INV_X1 U10263 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13380) );
  INV_X1 U10264 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8834) );
  INV_X1 U10265 ( .A(n14741), .ZN(n14761) );
  AND2_X1 U10266 ( .A1(n13512), .A2(n13496), .ZN(n8607) );
  AND2_X1 U10267 ( .A1(n8317), .A2(n7978), .ZN(n8335) );
  AND2_X1 U10268 ( .A1(n14845), .A2(n13814), .ZN(n15113) );
  AND4_X1 U10269 ( .A1(n7985), .A2(n7984), .A3(n7983), .A4(n7982), .ZN(n13424)
         );
  OR2_X1 U10270 ( .A1(n8136), .A2(n8135), .ZN(n8140) );
  OR2_X1 U10271 ( .A1(n10434), .A2(n10435), .ZN(n15136) );
  INV_X1 U10272 ( .A(n15136), .ZN(n15190) );
  AND2_X1 U10273 ( .A1(n10436), .A2(n10435), .ZN(n15198) );
  AND2_X1 U10274 ( .A1(n13793), .A2(n13792), .ZN(n13807) );
  INV_X1 U10275 ( .A(n15209), .ZN(n11196) );
  INV_X1 U10276 ( .A(n13807), .ZN(n13910) );
  AND2_X1 U10277 ( .A1(n15211), .A2(n9799), .ZN(n11197) );
  AND2_X1 U10278 ( .A1(n8581), .A2(n13957), .ZN(n15205) );
  AND2_X1 U10279 ( .A1(n8412), .A2(n8429), .ZN(n13545) );
  INV_X1 U10280 ( .A(n14965), .ZN(n14068) );
  AND2_X1 U10281 ( .A1(n14960), .A2(n14479), .ZN(n14087) );
  INV_X1 U10282 ( .A(n12372), .ZN(n10357) );
  AND4_X1 U10283 ( .A1(n9835), .A2(n9834), .A3(n9833), .A4(n9832), .ZN(n14274)
         );
  AND2_X1 U10284 ( .A1(n10161), .A2(n10160), .ZN(n13992) );
  AND2_X1 U10285 ( .A1(n11015), .A2(n11014), .ZN(n11020) );
  AND2_X1 U10286 ( .A1(n10647), .A2(n14629), .ZN(n14233) );
  INV_X1 U10287 ( .A(n14976), .ZN(n14206) );
  INV_X1 U10288 ( .A(n14235), .ZN(n11311) );
  NAND2_X1 U10289 ( .A1(n12569), .A2(n12568), .ZN(n12570) );
  INV_X1 U10290 ( .A(n14464), .ZN(n14477) );
  INV_X1 U10291 ( .A(n14490), .ZN(n14898) );
  NAND2_X1 U10292 ( .A1(n14508), .A2(n15052), .ZN(n14514) );
  AND2_X1 U10293 ( .A1(n15081), .A2(n15055), .ZN(n14599) );
  INV_X1 U10294 ( .A(n14599), .ZN(n15093) );
  AND2_X1 U10295 ( .A1(n11300), .A2(n11303), .ZN(n11156) );
  XNOR2_X1 U10296 ( .A(n10355), .B(n10354), .ZN(n10561) );
  INV_X1 U10297 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9843) );
  AND2_X1 U10298 ( .A1(n10049), .A2(n10071), .ZN(n11246) );
  AND2_X1 U10299 ( .A1(n10752), .A2(n10751), .ZN(n15280) );
  INV_X1 U10300 ( .A(n15425), .ZN(n12882) );
  INV_X1 U10301 ( .A(n15439), .ZN(n12848) );
  AND2_X1 U10302 ( .A1(n9229), .A2(n9228), .ZN(n11665) );
  NAND2_X1 U10303 ( .A1(n9026), .A2(n9025), .ZN(n13141) );
  INV_X1 U10304 ( .A(n12428), .ZN(n12901) );
  OR2_X2 U10305 ( .A1(n10934), .A2(n13378), .ZN(n12902) );
  NAND2_X1 U10306 ( .A1(n10738), .A2(n10737), .ZN(n13040) );
  INV_X1 U10307 ( .A(n13049), .ZN(n13004) );
  AND2_X1 U10308 ( .A1(n13160), .A2(n13159), .ZN(n13286) );
  AND2_X1 U10309 ( .A1(n12461), .A2(n12460), .ZN(n14825) );
  INV_X1 U10310 ( .A(n15323), .ZN(n13214) );
  NAND2_X1 U10311 ( .A1(n12802), .A2(n9187), .ZN(n9188) );
  NAND2_X1 U10312 ( .A1(n15419), .A2(n13290), .ZN(n13317) );
  AND2_X2 U10313 ( .A1(n11359), .A2(n9185), .ZN(n15419) );
  INV_X2 U10314 ( .A(n15409), .ZN(n15407) );
  INV_X1 U10315 ( .A(SI_13_), .ZN(n10560) );
  INV_X1 U10316 ( .A(n15166), .ZN(n15196) );
  NAND2_X1 U10317 ( .A1(n8608), .A2(n8607), .ZN(n8635) );
  INV_X1 U10318 ( .A(n15120), .ZN(n13481) );
  INV_X1 U10319 ( .A(n13424), .ZN(n13513) );
  OAI21_X1 U10320 ( .B1(n13706), .B2(n8137), .A(n8478), .ZN(n13684) );
  NAND2_X1 U10321 ( .A1(n10444), .A2(n10443), .ZN(n15204) );
  NAND2_X1 U10322 ( .A1(n13770), .A2(n11759), .ZN(n13832) );
  INV_X1 U10323 ( .A(n15279), .ZN(n15277) );
  NAND2_X1 U10324 ( .A1(n9800), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9801) );
  AND4_X1 U10325 ( .A1(n15234), .A2(n15233), .A3(n15232), .A4(n15231), .ZN(
        n15273) );
  AND2_X2 U10326 ( .A1(n11197), .A2(n15209), .ZN(n15270) );
  INV_X1 U10327 ( .A(n15207), .ZN(n15206) );
  NOR2_X1 U10328 ( .A1(n15212), .A2(n15205), .ZN(n15207) );
  INV_X1 U10329 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12212) );
  INV_X1 U10330 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11238) );
  INV_X1 U10331 ( .A(n12476), .ZN(n14781) );
  AND2_X1 U10332 ( .A1(n11502), .A2(n12372), .ZN(n14965) );
  INV_X1 U10333 ( .A(n14090), .ZN(n14864) );
  INV_X1 U10334 ( .A(n14076), .ZN(n14301) );
  OAI21_X1 U10335 ( .B1(n14378), .B2(n10278), .A(n10171), .ZN(n14359) );
  INV_X1 U10336 ( .A(n12670), .ZN(n14480) );
  INV_X1 U10337 ( .A(n14233), .ZN(n14974) );
  OR2_X1 U10338 ( .A1(n10844), .A2(n10649), .ZN(n14972) );
  AND2_X2 U10339 ( .A1(n11156), .A2(n10834), .ZN(n15107) );
  AND2_X2 U10340 ( .A1(n11302), .A2(n11156), .ZN(n15096) );
  AND2_X1 U10341 ( .A1(n10561), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12791) );
  INV_X1 U10342 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n15594) );
  INV_X1 U10343 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n11088) );
  NAND2_X1 U10344 ( .A1(n9415), .A2(n9414), .ZN(P3_U3296) );
  AND2_X1 U10345 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10418), .ZN(P2_U3947) );
  NOR2_X1 U10346 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n7956) );
  NOR2_X1 U10347 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .ZN(n7955) );
  NOR2_X1 U10348 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n7954) );
  NOR2_X1 U10349 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), 
        .ZN(n7953) );
  NAND4_X1 U10350 ( .A1(n7956), .A2(n7955), .A3(n7954), .A4(n7953), .ZN(n7957)
         );
  NOR2_X1 U10351 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), 
        .ZN(n7960) );
  NAND4_X1 U10352 ( .A1(n7960), .A2(n7959), .A3(n7958), .A4(n8312), .ZN(n8083)
         );
  INV_X1 U10353 ( .A(n8083), .ZN(n7965) );
  NOR2_X1 U10354 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7963) );
  NOR2_X1 U10355 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n7962) );
  NOR2_X1 U10356 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7961) );
  NAND2_X1 U10357 ( .A1(n7969), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n7971) );
  NAND2_X1 U10358 ( .A1(n9613), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n7985) );
  INV_X1 U10359 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n7974) );
  OR2_X1 U10360 ( .A1(n8139), .A2(n7974), .ZN(n7984) );
  NAND2_X1 U10361 ( .A1(n8185), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8202) );
  NOR2_X1 U10362 ( .A1(n8202), .A2(n8201), .ZN(n8224) );
  NAND2_X1 U10363 ( .A1(n8224), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8260) );
  NAND2_X1 U10364 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_8__SCAN_IN), 
        .ZN(n7977) );
  INV_X1 U10365 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8278) );
  INV_X1 U10366 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8376) );
  NAND2_X1 U10367 ( .A1(n8416), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8433) );
  INV_X1 U10368 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n15652) );
  NAND2_X1 U10369 ( .A1(n8489), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8490) );
  NAND2_X1 U10370 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n8508), .ZN(n8507) );
  NAND2_X1 U10371 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(n8521), .ZN(n8520) );
  INV_X1 U10372 ( .A(n8520), .ZN(n7979) );
  NAND2_X1 U10373 ( .A1(n7979), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8541) );
  INV_X1 U10374 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n7980) );
  NAND2_X1 U10375 ( .A1(n8520), .A2(n7980), .ZN(n7981) );
  NAND2_X1 U10376 ( .A1(n8541), .A2(n7981), .ZN(n13641) );
  OR2_X1 U10377 ( .A1(n8137), .A2(n13641), .ZN(n7983) );
  INV_X1 U10378 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n13642) );
  OR2_X1 U10379 ( .A1(n8138), .A2(n13642), .ZN(n7982) );
  XNOR2_X2 U10380 ( .A(n7989), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8080) );
  NAND2_X1 U10381 ( .A1(n7990), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7992) );
  NOR2_X1 U10382 ( .A1(n13424), .A2(n13690), .ZN(n8533) );
  INV_X1 U10383 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7993) );
  INV_X1 U10384 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10470) );
  XNOR2_X1 U10385 ( .A(n7999), .B(SI_1_), .ZN(n8109) );
  AND2_X1 U10386 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n7996) );
  NAND2_X1 U10387 ( .A1(n8013), .A2(n7996), .ZN(n9901) );
  AND2_X1 U10388 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7998) );
  NAND2_X1 U10389 ( .A1(n8004), .A2(n7998), .ZN(n8103) );
  NAND2_X1 U10390 ( .A1(n9901), .A2(n8103), .ZN(n8108) );
  INV_X1 U10391 ( .A(SI_1_), .ZN(n10466) );
  NOR2_X1 U10392 ( .A1(n7999), .A2(n10466), .ZN(n8000) );
  INV_X1 U10393 ( .A(n8132), .ZN(n8001) );
  INV_X1 U10394 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10481) );
  NAND2_X1 U10395 ( .A1(n8002), .A2(SI_2_), .ZN(n8003) );
  INV_X1 U10396 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10507) );
  INV_X1 U10397 ( .A(n8005), .ZN(n8006) );
  NAND2_X1 U10398 ( .A1(n8006), .A2(SI_3_), .ZN(n8007) );
  MUX2_X1 U10399 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n10485), .Z(n8009) );
  XNOR2_X1 U10400 ( .A(n8009), .B(SI_4_), .ZN(n8158) );
  INV_X1 U10401 ( .A(n8158), .ZN(n8008) );
  NAND2_X1 U10402 ( .A1(n8009), .A2(SI_4_), .ZN(n8010) );
  MUX2_X1 U10403 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n6546), .Z(n8012) );
  XNOR2_X1 U10404 ( .A(n8012), .B(SI_5_), .ZN(n8176) );
  INV_X1 U10405 ( .A(n8176), .ZN(n8011) );
  MUX2_X1 U10406 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n10486), .Z(n8015) );
  XNOR2_X1 U10407 ( .A(n8015), .B(SI_6_), .ZN(n8195) );
  INV_X1 U10408 ( .A(n8195), .ZN(n8014) );
  NAND2_X1 U10409 ( .A1(n8015), .A2(SI_6_), .ZN(n8213) );
  MUX2_X1 U10410 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n10486), .Z(n8017) );
  NAND2_X1 U10411 ( .A1(n8017), .A2(SI_7_), .ZN(n8016) );
  AND2_X1 U10412 ( .A1(n8213), .A2(n8016), .ZN(n8020) );
  INV_X1 U10413 ( .A(n8016), .ZN(n8019) );
  XNOR2_X1 U10414 ( .A(n8017), .B(SI_7_), .ZN(n8215) );
  INV_X1 U10415 ( .A(n8215), .ZN(n8018) );
  MUX2_X1 U10416 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10486), .Z(n8022) );
  XNOR2_X1 U10417 ( .A(n8022), .B(SI_8_), .ZN(n8235) );
  INV_X1 U10418 ( .A(n8235), .ZN(n8021) );
  NAND2_X1 U10419 ( .A1(n8022), .A2(SI_8_), .ZN(n8023) );
  MUX2_X1 U10420 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10486), .Z(n8025) );
  XNOR2_X1 U10421 ( .A(n8025), .B(n8024), .ZN(n8250) );
  NAND2_X1 U10422 ( .A1(n8025), .A2(SI_9_), .ZN(n8026) );
  MUX2_X1 U10423 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10486), .Z(n8028) );
  INV_X1 U10424 ( .A(SI_10_), .ZN(n8027) );
  NAND2_X1 U10425 ( .A1(n8030), .A2(n8029), .ZN(n8305) );
  INV_X1 U10426 ( .A(n8030), .ZN(n8031) );
  NAND2_X1 U10427 ( .A1(n8031), .A2(SI_11_), .ZN(n8032) );
  NAND2_X1 U10428 ( .A1(n8033), .A2(n6830), .ZN(n8308) );
  MUX2_X1 U10429 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n10486), .Z(n8327) );
  MUX2_X1 U10430 ( .A(n11088), .B(n15544), .S(n10485), .Z(n8348) );
  MUX2_X1 U10431 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n10486), .Z(n8038) );
  XNOR2_X1 U10432 ( .A(n8038), .B(SI_15_), .ZN(n8368) );
  INV_X1 U10433 ( .A(n8368), .ZN(n8037) );
  NAND2_X1 U10434 ( .A1(n8035), .A2(SI_14_), .ZN(n8036) );
  INV_X1 U10435 ( .A(n8038), .ZN(n8040) );
  MUX2_X1 U10436 ( .A(n15512), .B(n11183), .S(n10486), .Z(n8042) );
  XNOR2_X1 U10437 ( .A(n8042), .B(SI_16_), .ZN(n8386) );
  INV_X1 U10438 ( .A(SI_16_), .ZN(n8041) );
  NAND2_X1 U10439 ( .A1(n8042), .A2(n8041), .ZN(n8043) );
  MUX2_X1 U10440 ( .A(n11234), .B(n11236), .S(n10485), .Z(n8045) );
  INV_X1 U10441 ( .A(SI_18_), .ZN(n11185) );
  NAND2_X1 U10442 ( .A1(n8046), .A2(n11185), .ZN(n8047) );
  MUX2_X1 U10443 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n10486), .Z(n8427) );
  INV_X1 U10444 ( .A(n8427), .ZN(n8048) );
  MUX2_X1 U10445 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10485), .Z(n8050) );
  INV_X1 U10446 ( .A(SI_20_), .ZN(n11543) );
  MUX2_X1 U10447 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n10485), .Z(n8452) );
  MUX2_X1 U10448 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n6546), .Z(n8052) );
  OAI21_X1 U10449 ( .B1(SI_21_), .B2(n8052), .A(n8054), .ZN(n8053) );
  INV_X1 U10450 ( .A(n8053), .ZN(n8086) );
  INV_X1 U10451 ( .A(SI_22_), .ZN(n8055) );
  INV_X1 U10452 ( .A(n10186), .ZN(n8057) );
  INV_X1 U10453 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n15584) );
  MUX2_X1 U10454 ( .A(n15584), .B(n12212), .S(n10485), .Z(n8468) );
  MUX2_X1 U10455 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10486), .Z(n8059) );
  NAND2_X1 U10456 ( .A1(n8059), .A2(SI_23_), .ZN(n8061) );
  OAI21_X1 U10457 ( .B1(SI_23_), .B2(n8059), .A(n8061), .ZN(n8060) );
  INV_X1 U10458 ( .A(n8060), .ZN(n8482) );
  INV_X1 U10459 ( .A(n8063), .ZN(n8062) );
  INV_X1 U10460 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n14636) );
  INV_X1 U10461 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13966) );
  MUX2_X1 U10462 ( .A(n14636), .B(n13966), .S(n10486), .Z(n8500) );
  MUX2_X1 U10463 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n10485), .Z(n8066) );
  XNOR2_X1 U10464 ( .A(n8066), .B(SI_25_), .ZN(n8515) );
  INV_X1 U10465 ( .A(n8066), .ZN(n8067) );
  INV_X1 U10466 ( .A(SI_25_), .ZN(n12344) );
  NAND2_X1 U10467 ( .A1(n8067), .A2(n12344), .ZN(n8068) );
  INV_X1 U10468 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14632) );
  INV_X1 U10469 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13959) );
  MUX2_X1 U10470 ( .A(n14632), .B(n13959), .S(n10485), .Z(n8534) );
  XNOR2_X1 U10471 ( .A(n8534), .B(SI_26_), .ZN(n8069) );
  XNOR2_X1 U10472 ( .A(n8536), .B(n8069), .ZN(n13958) );
  MUX2_X1 U10473 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8075), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n8076) );
  NAND2_X2 U10474 ( .A1(n8126), .A2(n10485), .ZN(n9610) );
  NAND2_X1 U10475 ( .A1(n13958), .A2(n8148), .ZN(n8078) );
  NAND2_X1 U10476 ( .A1(n9624), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8077) );
  NAND2_X1 U10477 ( .A1(n8180), .A2(n8082), .ZN(n8311) );
  XNOR2_X1 U10478 ( .A(n13644), .B(n6558), .ZN(n8531) );
  OR2_X1 U10479 ( .A1(n8087), .A2(n8086), .ZN(n8088) );
  NAND2_X1 U10480 ( .A1(n8089), .A2(n8088), .ZN(n12052) );
  OR2_X1 U10481 ( .A1(n12052), .A2(n9610), .ZN(n8091) );
  NAND2_X1 U10482 ( .A1(n9624), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8090) );
  XNOR2_X1 U10483 ( .A(n13879), .B(n6558), .ZN(n8466) );
  NOR2_X1 U10484 ( .A1(n8458), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8092) );
  OR2_X1 U10485 ( .A1(n8473), .A2(n8092), .ZN(n13720) );
  INV_X1 U10486 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n13721) );
  NAND2_X1 U10487 ( .A1(n9613), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8094) );
  NAND2_X1 U10488 ( .A1(n9601), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8093) );
  OAI211_X1 U10489 ( .C1(n13721), .C2(n8138), .A(n8094), .B(n8093), .ZN(n8095)
         );
  INV_X1 U10490 ( .A(n8095), .ZN(n8096) );
  NAND2_X1 U10491 ( .A1(n13742), .A2(n8285), .ZN(n8467) );
  INV_X1 U10492 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11418) );
  INV_X1 U10493 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10621) );
  INV_X1 U10494 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n8098) );
  INV_X1 U10495 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10620) );
  OR2_X1 U10496 ( .A1(n8139), .A2(n10620), .ZN(n8099) );
  INV_X1 U10497 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n13534) );
  NAND2_X1 U10498 ( .A1(n10486), .A2(SI_0_), .ZN(n8102) );
  INV_X1 U10499 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8663) );
  NAND2_X1 U10500 ( .A1(n8102), .A2(n8663), .ZN(n8104) );
  INV_X1 U10501 ( .A(n8610), .ZN(n8604) );
  NAND2_X1 U10502 ( .A1(n9791), .A2(n8604), .ZN(n15213) );
  NAND2_X1 U10503 ( .A1(n9675), .A2(n15213), .ZN(n11414) );
  INV_X1 U10504 ( .A(n11414), .ZN(n8107) );
  NAND2_X1 U10505 ( .A1(n8107), .A2(n8106), .ZN(n11351) );
  XNOR2_X1 U10506 ( .A(n8109), .B(n8108), .ZN(n10487) );
  NAND2_X1 U10507 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8110) );
  MUX2_X1 U10508 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8110), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8112) );
  NAND2_X1 U10509 ( .A1(n6554), .A2(n13531), .ZN(n8113) );
  XNOR2_X1 U10510 ( .A(n6557), .B(n6553), .ZN(n8121) );
  INV_X1 U10511 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n8114) );
  AND2_X1 U10512 ( .A1(n8116), .A2(n8115), .ZN(n8120) );
  INV_X1 U10513 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n8117) );
  INV_X1 U10514 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n13528) );
  XNOR2_X1 U10515 ( .A(n8121), .B(n8122), .ZN(n11352) );
  NAND2_X1 U10516 ( .A1(n11351), .A2(n11352), .ZN(n8125) );
  INV_X1 U10517 ( .A(n8121), .ZN(n8123) );
  NAND2_X1 U10518 ( .A1(n8123), .A2(n8122), .ZN(n8124) );
  NOR2_X1 U10519 ( .A1(n8111), .A2(n13943), .ZN(n8127) );
  MUX2_X1 U10520 ( .A(n13943), .B(n8127), .S(P2_IR_REG_2__SCAN_IN), .Z(n8128)
         );
  INV_X1 U10521 ( .A(n8128), .ZN(n8130) );
  NAND2_X1 U10522 ( .A1(n8130), .A2(n8129), .ZN(n10730) );
  XNOR2_X1 U10523 ( .A(n8132), .B(n8131), .ZN(n10479) );
  INV_X1 U10524 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n8135) );
  INV_X1 U10525 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11780) );
  INV_X1 U10526 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10437) );
  INV_X1 U10527 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10424) );
  NAND2_X1 U10528 ( .A1(n13525), .A2(n8285), .ZN(n8142) );
  XNOR2_X1 U10529 ( .A(n8141), .B(n8142), .ZN(n11377) );
  NAND2_X1 U10530 ( .A1(n11378), .A2(n11377), .ZN(n8145) );
  INV_X1 U10531 ( .A(n8141), .ZN(n8143) );
  NAND2_X1 U10532 ( .A1(n8143), .A2(n8142), .ZN(n8144) );
  INV_X1 U10533 ( .A(n8146), .ZN(n8147) );
  NAND2_X1 U10534 ( .A1(n8129), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8149) );
  MUX2_X1 U10535 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8149), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n8151) );
  NAND2_X1 U10536 ( .A1(n8151), .A2(n8150), .ZN(n10492) );
  OAI22_X1 U10537 ( .A1(n8133), .A2(n10493), .B1(n7128), .B2(n10492), .ZN(
        n8152) );
  XNOR2_X1 U10538 ( .A(n12043), .B(n6558), .ZN(n8154) );
  INV_X1 U10539 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n12049) );
  INV_X1 U10540 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10428) );
  OR2_X1 U10541 ( .A1(n8139), .A2(n10428), .ZN(n8153) );
  AND2_X1 U10542 ( .A1(n13524), .A2(n8285), .ZN(n8155) );
  NAND2_X1 U10543 ( .A1(n8154), .A2(n8155), .ZN(n8172) );
  INV_X1 U10544 ( .A(n8154), .ZN(n11407) );
  INV_X1 U10545 ( .A(n8155), .ZN(n8156) );
  NAND2_X1 U10546 ( .A1(n11407), .A2(n8156), .ZN(n8157) );
  XNOR2_X1 U10547 ( .A(n8159), .B(n8158), .ZN(n10496) );
  NAND2_X1 U10548 ( .A1(n10496), .A2(n8148), .ZN(n8164) );
  NAND2_X1 U10549 ( .A1(n8150), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8161) );
  INV_X1 U10550 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8160) );
  XNOR2_X1 U10551 ( .A(n8161), .B(n8160), .ZN(n10578) );
  OAI22_X1 U10552 ( .A1(n8133), .A2(n10497), .B1(n7128), .B2(n10578), .ZN(
        n8162) );
  INV_X1 U10553 ( .A(n8162), .ZN(n8163) );
  NAND2_X1 U10554 ( .A1(n9613), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8171) );
  INV_X1 U10555 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10577) );
  OR2_X1 U10556 ( .A1(n8139), .A2(n10577), .ZN(n8170) );
  INV_X1 U10557 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11766) );
  OR2_X1 U10558 ( .A1(n8138), .A2(n11766), .ZN(n8169) );
  INV_X1 U10559 ( .A(n8185), .ZN(n8167) );
  INV_X1 U10560 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n12042) );
  INV_X1 U10561 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n8165) );
  NAND2_X1 U10562 ( .A1(n12042), .A2(n8165), .ZN(n8166) );
  NAND2_X1 U10563 ( .A1(n8167), .A2(n8166), .ZN(n11770) );
  OR2_X1 U10564 ( .A1(n8137), .A2(n11770), .ZN(n8168) );
  NAND2_X1 U10565 ( .A1(n13523), .A2(n8285), .ZN(n8173) );
  XNOR2_X1 U10566 ( .A(n11616), .B(n8173), .ZN(n11406) );
  INV_X1 U10567 ( .A(n11616), .ZN(n8174) );
  NAND2_X1 U10568 ( .A1(n8174), .A2(n8173), .ZN(n8175) );
  NAND2_X1 U10569 ( .A1(n11399), .A2(n8175), .ZN(n8190) );
  XNOR2_X1 U10570 ( .A(n8177), .B(n8176), .ZN(n10482) );
  NAND2_X1 U10571 ( .A1(n10482), .A2(n8148), .ZN(n8184) );
  NOR2_X1 U10572 ( .A1(n8178), .A2(n13943), .ZN(n8179) );
  MUX2_X1 U10573 ( .A(n13943), .B(n8179), .S(P2_IR_REG_5__SCAN_IN), .Z(n8181)
         );
  OR2_X1 U10574 ( .A1(n8181), .A2(n8180), .ZN(n10860) );
  OAI22_X1 U10575 ( .A1(n8133), .A2(n10490), .B1(n7128), .B2(n10860), .ZN(
        n8182) );
  INV_X1 U10576 ( .A(n8182), .ZN(n8183) );
  NAND2_X1 U10577 ( .A1(n8184), .A2(n8183), .ZN(n11837) );
  XNOR2_X1 U10578 ( .A(n11837), .B(n6558), .ZN(n8191) );
  NAND2_X1 U10579 ( .A1(n9613), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8189) );
  INV_X1 U10580 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10579) );
  OR2_X1 U10581 ( .A1(n8139), .A2(n10579), .ZN(n8188) );
  INV_X1 U10582 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11833) );
  OR2_X1 U10583 ( .A1(n8138), .A2(n11833), .ZN(n8187) );
  OAI21_X1 U10584 ( .B1(n8185), .B2(P2_REG3_REG_5__SCAN_IN), .A(n8202), .ZN(
        n11838) );
  OR2_X1 U10585 ( .A1(n8137), .A2(n11838), .ZN(n8186) );
  NAND4_X1 U10586 ( .A1(n8189), .A2(n8188), .A3(n8187), .A4(n8186), .ZN(n13522) );
  NAND2_X1 U10587 ( .A1(n13522), .A2(n8285), .ZN(n8192) );
  XNOR2_X1 U10588 ( .A(n8191), .B(n8192), .ZN(n11617) );
  INV_X1 U10589 ( .A(n8191), .ZN(n8193) );
  NAND2_X1 U10590 ( .A1(n8193), .A2(n8192), .ZN(n8194) );
  XNOR2_X1 U10591 ( .A(n8196), .B(n8195), .ZN(n10498) );
  NAND2_X1 U10592 ( .A1(n10498), .A2(n8148), .ZN(n8200) );
  OR2_X1 U10593 ( .A1(n8180), .A2(n13943), .ZN(n8197) );
  XNOR2_X1 U10594 ( .A(n8197), .B(n8217), .ZN(n10874) );
  OAI22_X1 U10595 ( .A1(n8133), .A2(n10499), .B1(n7128), .B2(n10874), .ZN(
        n8198) );
  INV_X1 U10596 ( .A(n8198), .ZN(n8199) );
  NAND2_X1 U10597 ( .A1(n8200), .A2(n8199), .ZN(n11815) );
  XNOR2_X1 U10598 ( .A(n11815), .B(n6558), .ZN(n11515) );
  NAND2_X1 U10599 ( .A1(n9613), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8207) );
  INV_X1 U10600 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10583) );
  OR2_X1 U10601 ( .A1(n8139), .A2(n10583), .ZN(n8206) );
  INV_X1 U10602 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11814) );
  OR2_X1 U10603 ( .A1(n8138), .A2(n11814), .ZN(n8205) );
  AND2_X1 U10604 ( .A1(n8202), .A2(n8201), .ZN(n8203) );
  OR2_X1 U10605 ( .A1(n8203), .A2(n8224), .ZN(n11816) );
  OR2_X1 U10606 ( .A1(n8137), .A2(n11816), .ZN(n8204) );
  NAND4_X1 U10607 ( .A1(n8207), .A2(n8206), .A3(n8205), .A4(n8204), .ZN(n13521) );
  AND2_X1 U10608 ( .A1(n13521), .A2(n8285), .ZN(n8208) );
  NAND2_X1 U10609 ( .A1(n11515), .A2(n8208), .ZN(n8212) );
  INV_X1 U10610 ( .A(n11515), .ZN(n8210) );
  INV_X1 U10611 ( .A(n8208), .ZN(n8209) );
  NAND2_X1 U10612 ( .A1(n8210), .A2(n8209), .ZN(n8211) );
  NAND2_X1 U10613 ( .A1(n8212), .A2(n8211), .ZN(n11373) );
  NAND2_X1 U10614 ( .A1(n8214), .A2(n8213), .ZN(n8216) );
  NAND2_X1 U10615 ( .A1(n10508), .A2(n8148), .ZN(n8222) );
  INV_X1 U10616 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10511) );
  NAND2_X1 U10617 ( .A1(n8180), .A2(n8217), .ZN(n8238) );
  NAND2_X1 U10618 ( .A1(n8238), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8219) );
  INV_X1 U10619 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n8218) );
  XNOR2_X1 U10620 ( .A(n8219), .B(n8218), .ZN(n10602) );
  OAI22_X1 U10621 ( .A1(n8133), .A2(n10511), .B1(n7128), .B2(n10602), .ZN(
        n8220) );
  INV_X1 U10622 ( .A(n8220), .ZN(n8221) );
  NAND2_X1 U10623 ( .A1(n8222), .A2(n8221), .ZN(n15245) );
  XNOR2_X1 U10624 ( .A(n15245), .B(n6558), .ZN(n8230) );
  NAND2_X1 U10625 ( .A1(n9601), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8229) );
  INV_X1 U10626 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n8223) );
  OR2_X1 U10627 ( .A1(n8136), .A2(n8223), .ZN(n8228) );
  OR2_X1 U10628 ( .A1(n8224), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8225) );
  NAND2_X1 U10629 ( .A1(n8260), .A2(n8225), .ZN(n11851) );
  OR2_X1 U10630 ( .A1(n8137), .A2(n11851), .ZN(n8227) );
  INV_X1 U10631 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11847) );
  OR2_X1 U10632 ( .A1(n8138), .A2(n11847), .ZN(n8226) );
  NAND4_X1 U10633 ( .A1(n8229), .A2(n8228), .A3(n8227), .A4(n8226), .ZN(n13520) );
  AND2_X1 U10634 ( .A1(n13520), .A2(n8285), .ZN(n8231) );
  NAND2_X1 U10635 ( .A1(n8230), .A2(n8231), .ZN(n8246) );
  INV_X1 U10636 ( .A(n8230), .ZN(n11450) );
  INV_X1 U10637 ( .A(n8231), .ZN(n8232) );
  NAND2_X1 U10638 ( .A1(n11450), .A2(n8232), .ZN(n8233) );
  AND2_X1 U10639 ( .A1(n8246), .A2(n8233), .ZN(n11516) );
  XNOR2_X1 U10640 ( .A(n8236), .B(n8235), .ZN(n10512) );
  NAND2_X1 U10641 ( .A1(n8254), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8239) );
  XNOR2_X1 U10642 ( .A(n8239), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10669) );
  AOI22_X1 U10643 ( .A1(n9624), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8237), .B2(
        n10669), .ZN(n8240) );
  XNOR2_X1 U10644 ( .A(n11611), .B(n6558), .ZN(n11633) );
  NAND2_X1 U10645 ( .A1(n9601), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8245) );
  INV_X1 U10646 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11805) );
  OR2_X1 U10647 ( .A1(n8138), .A2(n11805), .ZN(n8244) );
  INV_X1 U10648 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8259) );
  XNOR2_X1 U10649 ( .A(n8260), .B(n8259), .ZN(n11806) );
  OR2_X1 U10650 ( .A1(n8137), .A2(n11806), .ZN(n8243) );
  INV_X1 U10651 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n8241) );
  OR2_X1 U10652 ( .A1(n8136), .A2(n8241), .ZN(n8242) );
  NAND4_X1 U10653 ( .A1(n8245), .A2(n8244), .A3(n8243), .A4(n8242), .ZN(n13519) );
  NAND2_X1 U10654 ( .A1(n13519), .A2(n8285), .ZN(n8248) );
  XNOR2_X1 U10655 ( .A(n11633), .B(n8248), .ZN(n11452) );
  AND2_X1 U10656 ( .A1(n11452), .A2(n8246), .ZN(n8247) );
  INV_X1 U10657 ( .A(n11633), .ZN(n8249) );
  OR2_X1 U10658 ( .A1(n8251), .A2(n8250), .ZN(n8252) );
  NAND2_X1 U10659 ( .A1(n8253), .A2(n8252), .ZN(n10518) );
  OR2_X1 U10660 ( .A1(n10518), .A2(n9610), .ZN(n8257) );
  NAND2_X1 U10661 ( .A1(n8271), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8255) );
  XNOR2_X1 U10662 ( .A(n8255), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10814) );
  AOI22_X1 U10663 ( .A1(n9624), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n10814), 
        .B2(n8237), .ZN(n8256) );
  XNOR2_X1 U10664 ( .A(n15252), .B(n6558), .ZN(n8266) );
  NAND2_X1 U10665 ( .A1(n9613), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8265) );
  INV_X1 U10666 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10673) );
  OR2_X1 U10667 ( .A1(n8139), .A2(n10673), .ZN(n8264) );
  INV_X1 U10668 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n12083) );
  OR2_X1 U10669 ( .A1(n8138), .A2(n12083), .ZN(n8263) );
  INV_X1 U10670 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8258) );
  OAI21_X1 U10671 ( .B1(n8260), .B2(n8259), .A(n8258), .ZN(n8261) );
  NAND2_X1 U10672 ( .A1(n8261), .A2(n8279), .ZN(n12082) );
  OR2_X1 U10673 ( .A1(n8137), .A2(n12082), .ZN(n8262) );
  NAND4_X1 U10674 ( .A1(n8265), .A2(n8264), .A3(n8263), .A4(n8262), .ZN(n13518) );
  NAND2_X1 U10675 ( .A1(n13518), .A2(n8285), .ZN(n8267) );
  XNOR2_X1 U10676 ( .A(n8266), .B(n8267), .ZN(n11634) );
  INV_X1 U10677 ( .A(n8266), .ZN(n8268) );
  NAND2_X1 U10678 ( .A1(n8268), .A2(n8267), .ZN(n8269) );
  NAND2_X1 U10679 ( .A1(n10565), .A2(n8148), .ZN(n8276) );
  INV_X1 U10680 ( .A(n8271), .ZN(n8273) );
  INV_X1 U10681 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8272) );
  NAND2_X1 U10682 ( .A1(n8273), .A2(n8272), .ZN(n8292) );
  NAND2_X1 U10683 ( .A1(n8292), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8274) );
  XNOR2_X1 U10684 ( .A(n8274), .B(P2_IR_REG_10__SCAN_IN), .ZN(n11040) );
  AOI22_X1 U10685 ( .A1(n11040), .A2(n8237), .B1(P1_DATAO_REG_10__SCAN_IN), 
        .B2(n9624), .ZN(n8275) );
  XNOR2_X1 U10686 ( .A(n12102), .B(n6558), .ZN(n8286) );
  NAND2_X1 U10687 ( .A1(n9613), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8284) );
  INV_X1 U10688 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8277) );
  OR2_X1 U10689 ( .A1(n8139), .A2(n8277), .ZN(n8283) );
  INV_X1 U10690 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n12097) );
  OR2_X1 U10691 ( .A1(n8138), .A2(n12097), .ZN(n8282) );
  AND2_X1 U10692 ( .A1(n8279), .A2(n8278), .ZN(n8280) );
  OR2_X1 U10693 ( .A1(n8280), .A2(n8317), .ZN(n12096) );
  OR2_X1 U10694 ( .A1(n8137), .A2(n12096), .ZN(n8281) );
  NAND4_X1 U10695 ( .A1(n8284), .A2(n8283), .A3(n8282), .A4(n8281), .ZN(n13517) );
  AND2_X1 U10696 ( .A1(n13517), .A2(n8285), .ZN(n8287) );
  NAND2_X1 U10697 ( .A1(n8286), .A2(n8287), .ZN(n8300) );
  INV_X1 U10698 ( .A(n8286), .ZN(n11793) );
  INV_X1 U10699 ( .A(n8287), .ZN(n8288) );
  NAND2_X1 U10700 ( .A1(n11793), .A2(n8288), .ZN(n8289) );
  NAND2_X1 U10701 ( .A1(n8300), .A2(n8289), .ZN(n11931) );
  XNOR2_X1 U10702 ( .A(n8291), .B(n8290), .ZN(n10570) );
  NAND2_X1 U10703 ( .A1(n10570), .A2(n8148), .ZN(n8295) );
  OAI21_X1 U10704 ( .B1(n8292), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8293) );
  XNOR2_X1 U10705 ( .A(n8293), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11044) );
  AOI22_X1 U10706 ( .A1(n11044), .A2(n8237), .B1(n9624), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n8294) );
  XNOR2_X1 U10707 ( .A(n12214), .B(n6558), .ZN(n8301) );
  NAND2_X1 U10708 ( .A1(n9613), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8299) );
  INV_X1 U10709 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11041) );
  OR2_X1 U10710 ( .A1(n8139), .A2(n11041), .ZN(n8298) );
  INV_X1 U10711 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n13549) );
  OR2_X1 U10712 ( .A1(n8138), .A2(n13549), .ZN(n8297) );
  XNOR2_X1 U10713 ( .A(n8317), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n11796) );
  OR2_X1 U10714 ( .A1(n8137), .A2(n11796), .ZN(n8296) );
  NAND4_X1 U10715 ( .A1(n8299), .A2(n8298), .A3(n8297), .A4(n8296), .ZN(n15112) );
  NAND2_X1 U10716 ( .A1(n15112), .A2(n8285), .ZN(n8302) );
  XNOR2_X1 U10717 ( .A(n8301), .B(n8302), .ZN(n11794) );
  INV_X1 U10718 ( .A(n8301), .ZN(n8303) );
  NAND2_X1 U10719 ( .A1(n8303), .A2(n8302), .ZN(n8304) );
  NAND2_X1 U10720 ( .A1(n8306), .A2(n8305), .ZN(n8310) );
  AND2_X1 U10721 ( .A1(n8308), .A2(n8307), .ZN(n8309) );
  NAND2_X1 U10722 ( .A1(n10615), .A2(n8148), .ZN(n8316) );
  NAND2_X1 U10723 ( .A1(n8311), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8313) );
  XNOR2_X1 U10724 ( .A(n8313), .B(n8312), .ZN(n15135) );
  OAI22_X1 U10725 ( .A1(n8133), .A2(n15461), .B1(n7128), .B2(n15135), .ZN(
        n8314) );
  INV_X1 U10726 ( .A(n8314), .ZN(n8315) );
  XNOR2_X1 U10727 ( .A(n12253), .B(n8415), .ZN(n8323) );
  NAND2_X1 U10728 ( .A1(n9613), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8322) );
  INV_X1 U10729 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n13564) );
  OR2_X1 U10730 ( .A1(n8139), .A2(n13564), .ZN(n8321) );
  INV_X1 U10731 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n13550) );
  OR2_X1 U10732 ( .A1(n8138), .A2(n13550), .ZN(n8320) );
  AOI21_X1 U10733 ( .B1(n8317), .B2(P2_REG3_REG_11__SCAN_IN), .A(
        P2_REG3_REG_12__SCAN_IN), .ZN(n8318) );
  OR2_X1 U10734 ( .A1(n8335), .A2(n8318), .ZN(n15123) );
  OR2_X1 U10735 ( .A1(n8137), .A2(n15123), .ZN(n8319) );
  NAND4_X1 U10736 ( .A1(n8322), .A2(n8321), .A3(n8320), .A4(n8319), .ZN(n13516) );
  NAND2_X1 U10737 ( .A1(n13516), .A2(n8285), .ZN(n8324) );
  NAND2_X1 U10738 ( .A1(n8323), .A2(n8324), .ZN(n15109) );
  INV_X1 U10739 ( .A(n8323), .ZN(n8326) );
  INV_X1 U10740 ( .A(n8324), .ZN(n8325) );
  NAND2_X1 U10741 ( .A1(n8326), .A2(n8325), .ZN(n15108) );
  XNOR2_X1 U10742 ( .A(n8327), .B(n10560), .ZN(n8328) );
  XNOR2_X1 U10743 ( .A(n8329), .B(n8328), .ZN(n10627) );
  NAND2_X1 U10744 ( .A1(n10627), .A2(n8148), .ZN(n8334) );
  NAND2_X1 U10745 ( .A1(n8351), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8331) );
  INV_X1 U10746 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8330) );
  XNOR2_X1 U10747 ( .A(n8331), .B(n8330), .ZN(n15148) );
  OAI22_X1 U10748 ( .A1(n8133), .A2(n15654), .B1(n15148), .B2(n7128), .ZN(
        n8332) );
  INV_X1 U10749 ( .A(n8332), .ZN(n8333) );
  XNOR2_X1 U10750 ( .A(n12420), .B(n6558), .ZN(n8343) );
  NAND2_X1 U10751 ( .A1(n9613), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8340) );
  INV_X1 U10752 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n13565) );
  OR2_X1 U10753 ( .A1(n8139), .A2(n13565), .ZN(n8339) );
  INV_X1 U10754 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n13551) );
  OR2_X1 U10755 ( .A1(n8138), .A2(n13551), .ZN(n8338) );
  OR2_X1 U10756 ( .A1(n8335), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8336) );
  NAND2_X1 U10757 ( .A1(n8377), .A2(n8336), .ZN(n12233) );
  OR2_X1 U10758 ( .A1(n8137), .A2(n12233), .ZN(n8337) );
  NAND4_X1 U10759 ( .A1(n8340), .A2(n8339), .A3(n8338), .A4(n8337), .ZN(n15114) );
  NAND2_X1 U10760 ( .A1(n15114), .A2(n8285), .ZN(n8341) );
  XNOR2_X1 U10761 ( .A(n8343), .B(n8341), .ZN(n12056) );
  NAND2_X1 U10762 ( .A1(n12055), .A2(n12056), .ZN(n8345) );
  INV_X1 U10763 ( .A(n8341), .ZN(n8342) );
  NAND2_X1 U10764 ( .A1(n8343), .A2(n8342), .ZN(n8344) );
  INV_X1 U10765 ( .A(SI_14_), .ZN(n10618) );
  NAND2_X1 U10766 ( .A1(n8346), .A2(n10618), .ZN(n8347) );
  NAND2_X1 U10767 ( .A1(n8349), .A2(n8348), .ZN(n8350) );
  NAND2_X1 U10768 ( .A1(n8367), .A2(n8350), .ZN(n11087) );
  OR2_X1 U10769 ( .A1(n11087), .A2(n9610), .ZN(n8354) );
  OR2_X1 U10770 ( .A1(n8351), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n8370) );
  NAND2_X1 U10771 ( .A1(n8370), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8352) );
  XNOR2_X1 U10772 ( .A(n8352), .B(P2_IR_REG_14__SCAN_IN), .ZN(n13552) );
  AOI22_X1 U10773 ( .A1(n8237), .A2(n13552), .B1(n9624), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n8353) );
  XNOR2_X1 U10774 ( .A(n14847), .B(n8415), .ZN(n8360) );
  NAND2_X1 U10775 ( .A1(n9613), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8359) );
  INV_X1 U10776 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n13566) );
  OR2_X1 U10777 ( .A1(n8139), .A2(n13566), .ZN(n8358) );
  XNOR2_X1 U10778 ( .A(n8377), .B(n8376), .ZN(n14850) );
  OR2_X1 U10779 ( .A1(n8137), .A2(n14850), .ZN(n8357) );
  INV_X1 U10780 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8355) );
  OR2_X1 U10781 ( .A1(n8138), .A2(n8355), .ZN(n8356) );
  NAND4_X1 U10782 ( .A1(n8359), .A2(n8358), .A3(n8357), .A4(n8356), .ZN(n13815) );
  NAND2_X1 U10783 ( .A1(n13815), .A2(n8285), .ZN(n8361) );
  NAND2_X1 U10784 ( .A1(n8360), .A2(n8361), .ZN(n8365) );
  INV_X1 U10785 ( .A(n8360), .ZN(n8363) );
  INV_X1 U10786 ( .A(n8361), .ZN(n8362) );
  NAND2_X1 U10787 ( .A1(n8363), .A2(n8362), .ZN(n8364) );
  NAND2_X1 U10788 ( .A1(n8365), .A2(n8364), .ZN(n14840) );
  NAND2_X1 U10789 ( .A1(n8367), .A2(n8366), .ZN(n8369) );
  NAND2_X1 U10790 ( .A1(n11237), .A2(n8148), .ZN(n8373) );
  NOR2_X1 U10791 ( .A1(n8370), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n8389) );
  OR2_X1 U10792 ( .A1(n8389), .A2(n13943), .ZN(n8371) );
  XNOR2_X1 U10793 ( .A(n8371), .B(P2_IR_REG_15__SCAN_IN), .ZN(n15169) );
  AOI22_X1 U10794 ( .A1(n15169), .A2(n8237), .B1(n9624), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n8372) );
  INV_X1 U10795 ( .A(n13912), .ZN(n13829) );
  NAND2_X1 U10796 ( .A1(n9613), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8383) );
  INV_X1 U10797 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8374) );
  OR2_X1 U10798 ( .A1(n8139), .A2(n8374), .ZN(n8382) );
  OAI21_X1 U10799 ( .B1(n8377), .B2(n8376), .A(n8375), .ZN(n8378) );
  NAND2_X1 U10800 ( .A1(n8378), .A2(n8394), .ZN(n13824) );
  OR2_X1 U10801 ( .A1(n8137), .A2(n13824), .ZN(n8381) );
  INV_X1 U10802 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8379) );
  OR2_X1 U10803 ( .A1(n8138), .A2(n8379), .ZN(n8380) );
  NAND4_X1 U10804 ( .A1(n8383), .A2(n8382), .A3(n8381), .A4(n8380), .ZN(n13796) );
  NAND2_X1 U10805 ( .A1(n13796), .A2(n8285), .ZN(n13495) );
  XNOR2_X1 U10806 ( .A(n8387), .B(n8386), .ZN(n11181) );
  NAND2_X1 U10807 ( .A1(n11181), .A2(n8148), .ZN(n8392) );
  INV_X1 U10808 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8388) );
  NAND2_X1 U10809 ( .A1(n8389), .A2(n8388), .ZN(n8407) );
  NAND2_X1 U10810 ( .A1(n8407), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8390) );
  XNOR2_X1 U10811 ( .A(n8390), .B(P2_IR_REG_16__SCAN_IN), .ZN(n13547) );
  AOI22_X1 U10812 ( .A1(n13547), .A2(n8237), .B1(n9624), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n8391) );
  XNOR2_X1 U10813 ( .A(n13907), .B(n8415), .ZN(n8402) );
  AND2_X1 U10814 ( .A1(n8394), .A2(n8393), .ZN(n8395) );
  NOR2_X1 U10815 ( .A1(n8416), .A2(n8395), .ZN(n13804) );
  NAND2_X1 U10816 ( .A1(n13804), .A2(n8492), .ZN(n8400) );
  NAND2_X1 U10817 ( .A1(n9601), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8399) );
  NAND2_X1 U10818 ( .A1(n9613), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8398) );
  INV_X1 U10819 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8396) );
  OR2_X1 U10820 ( .A1(n8138), .A2(n8396), .ZN(n8397) );
  NAND4_X1 U10821 ( .A1(n8400), .A2(n8399), .A3(n8398), .A4(n8397), .ZN(n13817) );
  NAND2_X1 U10822 ( .A1(n13817), .A2(n8285), .ZN(n8401) );
  NAND2_X1 U10823 ( .A1(n8402), .A2(n8401), .ZN(n8403) );
  OAI21_X1 U10824 ( .B1(n8402), .B2(n8401), .A(n8403), .ZN(n13439) );
  INV_X1 U10825 ( .A(n8403), .ZN(n8404) );
  XNOR2_X1 U10826 ( .A(n8406), .B(n8405), .ZN(n11233) );
  NAND2_X1 U10827 ( .A1(n11233), .A2(n8148), .ZN(n8414) );
  NAND2_X1 U10828 ( .A1(n8408), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8411) );
  INV_X1 U10829 ( .A(n8411), .ZN(n8409) );
  NAND2_X1 U10830 ( .A1(n8409), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n8412) );
  INV_X1 U10831 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8410) );
  NAND2_X1 U10832 ( .A1(n8411), .A2(n8410), .ZN(n8429) );
  AOI22_X1 U10833 ( .A1(n13545), .A2(n8237), .B1(n9624), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n8413) );
  XNOR2_X1 U10834 ( .A(n13903), .B(n8415), .ZN(n8424) );
  OR2_X1 U10835 ( .A1(n8416), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8417) );
  NAND2_X1 U10836 ( .A1(n8433), .A2(n8417), .ZN(n13785) );
  INV_X1 U10837 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13571) );
  OR2_X1 U10838 ( .A1(n8139), .A2(n13571), .ZN(n8420) );
  INV_X1 U10839 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8418) );
  OR2_X1 U10840 ( .A1(n8136), .A2(n8418), .ZN(n8419) );
  AND2_X1 U10841 ( .A1(n8420), .A2(n8419), .ZN(n8422) );
  INV_X1 U10842 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13786) );
  OR2_X1 U10843 ( .A1(n8138), .A2(n13786), .ZN(n8421) );
  OAI211_X1 U10844 ( .C1(n13785), .C2(n8137), .A(n8422), .B(n8421), .ZN(n13797) );
  NAND2_X1 U10845 ( .A1(n13797), .A2(n8285), .ZN(n8423) );
  NAND2_X1 U10846 ( .A1(n8424), .A2(n8423), .ZN(n8425) );
  OAI21_X1 U10847 ( .B1(n8424), .B2(n8423), .A(n8425), .ZN(n13447) );
  INV_X1 U10848 ( .A(n8425), .ZN(n8426) );
  XNOR2_X1 U10849 ( .A(n8428), .B(n8427), .ZN(n11465) );
  NAND2_X1 U10850 ( .A1(n11465), .A2(n8148), .ZN(n8432) );
  NAND2_X1 U10851 ( .A1(n8429), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8430) );
  XNOR2_X1 U10852 ( .A(n8430), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13581) );
  AOI22_X1 U10853 ( .A1(n13581), .A2(n8237), .B1(n9624), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n8431) );
  XNOR2_X1 U10854 ( .A(n13898), .B(n6558), .ZN(n8438) );
  NAND2_X1 U10855 ( .A1(n8433), .A2(n15652), .ZN(n8434) );
  NAND2_X1 U10856 ( .A1(n8441), .A2(n8434), .ZN(n13768) );
  INV_X1 U10857 ( .A(n8138), .ZN(n9612) );
  AOI22_X1 U10858 ( .A1(n9601), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n9612), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n8436) );
  NAND2_X1 U10859 ( .A1(n9613), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8435) );
  OAI211_X1 U10860 ( .C1(n13768), .C2(n8137), .A(n8436), .B(n8435), .ZN(n13515) );
  NAND2_X1 U10861 ( .A1(n13515), .A2(n8285), .ZN(n8437) );
  XNOR2_X1 U10862 ( .A(n8438), .B(n8437), .ZN(n13474) );
  INV_X1 U10863 ( .A(n8437), .ZN(n8439) );
  AND2_X1 U10864 ( .A1(n8441), .A2(n8440), .ZN(n8442) );
  OR2_X1 U10865 ( .A1(n8442), .A2(n8456), .ZN(n13410) );
  AOI22_X1 U10866 ( .A1(n9613), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n9601), .B2(
        P2_REG1_REG_19__SCAN_IN), .ZN(n8444) );
  NAND2_X1 U10867 ( .A1(n9612), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8443) );
  OAI211_X1 U10868 ( .C1(n13410), .C2(n8137), .A(n8444), .B(n8443), .ZN(n13741) );
  AND2_X1 U10869 ( .A1(n13741), .A2(n8285), .ZN(n8450) );
  XNOR2_X1 U10870 ( .A(n8446), .B(n8445), .ZN(n11628) );
  NAND2_X1 U10871 ( .A1(n11628), .A2(n8148), .ZN(n8448) );
  AOI22_X1 U10872 ( .A1(n9624), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9698), 
        .B2(n8237), .ZN(n8447) );
  XNOR2_X1 U10873 ( .A(n13893), .B(n6558), .ZN(n8449) );
  NOR2_X1 U10874 ( .A1(n8449), .A2(n8450), .ZN(n8451) );
  AOI21_X1 U10875 ( .B1(n8450), .B2(n8449), .A(n8451), .ZN(n13407) );
  XNOR2_X1 U10876 ( .A(n8453), .B(n8452), .ZN(n11896) );
  NAND2_X1 U10877 ( .A1(n11896), .A2(n8148), .ZN(n8455) );
  NAND2_X1 U10878 ( .A1(n9624), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8454) );
  XNOR2_X1 U10879 ( .A(n13887), .B(n6558), .ZN(n8465) );
  NOR2_X1 U10880 ( .A1(n8456), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8457) );
  OR2_X1 U10881 ( .A1(n8458), .A2(n8457), .ZN(n13737) );
  INV_X1 U10882 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8461) );
  NAND2_X1 U10883 ( .A1(n9612), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8460) );
  NAND2_X1 U10884 ( .A1(n9601), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8459) );
  OAI211_X1 U10885 ( .C1(n8136), .C2(n8461), .A(n8460), .B(n8459), .ZN(n8462)
         );
  INV_X1 U10886 ( .A(n8462), .ZN(n8463) );
  OAI21_X1 U10887 ( .B1(n13737), .B2(n8137), .A(n8463), .ZN(n13514) );
  AND2_X1 U10888 ( .A1(n13514), .A2(n8285), .ZN(n8464) );
  NOR2_X1 U10889 ( .A1(n8465), .A2(n8464), .ZN(n13462) );
  NAND2_X1 U10890 ( .A1(n8465), .A2(n8464), .ZN(n13463) );
  XNOR2_X1 U10891 ( .A(n8466), .B(n8467), .ZN(n13415) );
  NAND2_X1 U10892 ( .A1(n10186), .A2(n8468), .ZN(n8469) );
  NAND2_X1 U10893 ( .A1(n8470), .A2(n8469), .ZN(n12210) );
  NAND2_X1 U10894 ( .A1(n9624), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8471) );
  XNOR2_X1 U10895 ( .A(n13875), .B(n6558), .ZN(n8479) );
  NOR2_X1 U10896 ( .A1(n8473), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8474) );
  OR2_X1 U10897 ( .A1(n8489), .A2(n8474), .ZN(n13706) );
  INV_X1 U10898 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13707) );
  NAND2_X1 U10899 ( .A1(n9613), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8476) );
  NAND2_X1 U10900 ( .A1(n9601), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8475) );
  OAI211_X1 U10901 ( .C1(n13707), .C2(n8138), .A(n8476), .B(n8475), .ZN(n8477)
         );
  INV_X1 U10902 ( .A(n8477), .ZN(n8478) );
  INV_X1 U10903 ( .A(n13684), .ZN(n13418) );
  AND2_X1 U10904 ( .A1(n8480), .A2(n8479), .ZN(n8481) );
  OR2_X1 U10905 ( .A1(n8483), .A2(n8482), .ZN(n8484) );
  AND2_X1 U10906 ( .A1(n8485), .A2(n8484), .ZN(n12402) );
  NAND2_X1 U10907 ( .A1(n12402), .A2(n8148), .ZN(n8487) );
  NAND2_X1 U10908 ( .A1(n9624), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8486) );
  XNOR2_X1 U10909 ( .A(n13870), .B(n6558), .ZN(n8488) );
  OR2_X1 U10910 ( .A1(n8489), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8491) );
  AND2_X1 U10911 ( .A1(n8491), .A2(n8490), .ZN(n13694) );
  NAND2_X1 U10912 ( .A1(n13694), .A2(n8492), .ZN(n8498) );
  INV_X1 U10913 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8495) );
  NAND2_X1 U10914 ( .A1(n9613), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8494) );
  NAND2_X1 U10915 ( .A1(n9601), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8493) );
  OAI211_X1 U10916 ( .C1(n8495), .C2(n8138), .A(n8494), .B(n8493), .ZN(n8496)
         );
  INV_X1 U10917 ( .A(n8496), .ZN(n8497) );
  NAND2_X1 U10918 ( .A1(n8498), .A2(n8497), .ZN(n13669) );
  NAND2_X1 U10919 ( .A1(n8501), .A2(n8500), .ZN(n8502) );
  NAND2_X1 U10920 ( .A1(n13965), .A2(n8148), .ZN(n8505) );
  NAND2_X1 U10921 ( .A1(n9624), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8504) );
  XNOR2_X1 U10922 ( .A(n13677), .B(n6558), .ZN(n13428) );
  NAND2_X1 U10923 ( .A1(n9613), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8513) );
  INV_X1 U10924 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8506) );
  OR2_X1 U10925 ( .A1(n8139), .A2(n8506), .ZN(n8512) );
  OAI21_X1 U10926 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n8508), .A(n8507), .ZN(
        n13674) );
  OR2_X1 U10927 ( .A1(n8137), .A2(n13674), .ZN(n8511) );
  INV_X1 U10928 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8509) );
  OR2_X1 U10929 ( .A1(n8138), .A2(n8509), .ZN(n8510) );
  OR2_X1 U10930 ( .A1(n13426), .A2(n13690), .ZN(n8514) );
  NOR2_X1 U10931 ( .A1(n13428), .A2(n8514), .ZN(n8530) );
  AOI21_X1 U10932 ( .B1(n13428), .B2(n8514), .A(n8530), .ZN(n13456) );
  XNOR2_X1 U10933 ( .A(n8516), .B(n8515), .ZN(n12794) );
  NAND2_X1 U10934 ( .A1(n12794), .A2(n8148), .ZN(n8518) );
  NAND2_X1 U10935 ( .A1(n9624), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8517) );
  XNOR2_X1 U10936 ( .A(n13860), .B(n6558), .ZN(n8526) );
  NAND2_X1 U10937 ( .A1(n9613), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8525) );
  INV_X1 U10938 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8519) );
  OR2_X1 U10939 ( .A1(n8139), .A2(n8519), .ZN(n8524) );
  INV_X1 U10940 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13658) );
  OR2_X1 U10941 ( .A1(n8138), .A2(n13658), .ZN(n8523) );
  OAI21_X1 U10942 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n8521), .A(n8520), .ZN(
        n13657) );
  OR2_X1 U10943 ( .A1(n8137), .A2(n13657), .ZN(n8522) );
  NAND4_X1 U10944 ( .A1(n8525), .A2(n8524), .A3(n8523), .A4(n8522), .ZN(n13668) );
  AND2_X1 U10945 ( .A1(n13668), .A2(n8285), .ZN(n8527) );
  NAND2_X1 U10946 ( .A1(n8526), .A2(n8527), .ZN(n8532) );
  INV_X1 U10947 ( .A(n8526), .ZN(n13489) );
  INV_X1 U10948 ( .A(n8527), .ZN(n8528) );
  NAND2_X1 U10949 ( .A1(n13489), .A2(n8528), .ZN(n8529) );
  AND2_X1 U10950 ( .A1(n8532), .A2(n8529), .ZN(n13430) );
  XNOR2_X1 U10951 ( .A(n8531), .B(n8533), .ZN(n13490) );
  INV_X1 U10952 ( .A(n8534), .ZN(n8535) );
  MUX2_X1 U10953 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n10485), .Z(n9583) );
  NAND2_X1 U10954 ( .A1(n13954), .A2(n8148), .ZN(n8538) );
  NAND2_X1 U10955 ( .A1(n9624), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8537) );
  XNOR2_X1 U10956 ( .A(n13849), .B(n6558), .ZN(n8548) );
  NAND2_X1 U10957 ( .A1(n9613), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8546) );
  INV_X1 U10958 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n15559) );
  OR2_X1 U10959 ( .A1(n8139), .A2(n15559), .ZN(n8545) );
  INV_X1 U10960 ( .A(n8541), .ZN(n8539) );
  NAND2_X1 U10961 ( .A1(n8539), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8565) );
  INV_X1 U10962 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8540) );
  NAND2_X1 U10963 ( .A1(n8541), .A2(n8540), .ZN(n8542) );
  NAND2_X1 U10964 ( .A1(n8565), .A2(n8542), .ZN(n13629) );
  OR2_X1 U10965 ( .A1(n8137), .A2(n13629), .ZN(n8544) );
  INV_X1 U10966 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13630) );
  OR2_X1 U10967 ( .A1(n8138), .A2(n13630), .ZN(n8543) );
  NAND4_X1 U10968 ( .A1(n8546), .A2(n8545), .A3(n8544), .A4(n8543), .ZN(n13637) );
  AND2_X1 U10969 ( .A1(n13637), .A2(n8285), .ZN(n8547) );
  NAND2_X1 U10970 ( .A1(n8548), .A2(n8547), .ZN(n8549) );
  OAI21_X1 U10971 ( .B1(n8548), .B2(n8547), .A(n8549), .ZN(n13391) );
  INV_X1 U10972 ( .A(n8549), .ZN(n8550) );
  INV_X1 U10973 ( .A(n8551), .ZN(n8552) );
  NAND2_X1 U10974 ( .A1(n8552), .A2(SI_27_), .ZN(n8554) );
  NAND2_X1 U10975 ( .A1(n9589), .A2(n9583), .ZN(n8553) );
  NAND2_X1 U10976 ( .A1(n8554), .A2(n8553), .ZN(n8558) );
  MUX2_X1 U10977 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n6546), .Z(n8555) );
  NAND2_X1 U10978 ( .A1(n8555), .A2(SI_28_), .ZN(n9585) );
  NOR2_X1 U10979 ( .A1(n8555), .A2(SI_28_), .ZN(n9584) );
  INV_X1 U10980 ( .A(n9584), .ZN(n8556) );
  NAND2_X1 U10981 ( .A1(n9585), .A2(n8556), .ZN(n8557) );
  NAND2_X1 U10982 ( .A1(n12536), .A2(n8148), .ZN(n8560) );
  NAND2_X1 U10983 ( .A1(n9624), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8559) );
  NAND2_X2 U10984 ( .A1(n8560), .A2(n8559), .ZN(n13843) );
  XNOR2_X1 U10985 ( .A(n13843), .B(n6558), .ZN(n8561) );
  NAND2_X1 U10986 ( .A1(n9613), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8570) );
  INV_X1 U10987 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8562) );
  OR2_X1 U10988 ( .A1(n8139), .A2(n8562), .ZN(n8569) );
  INV_X1 U10989 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13614) );
  OR2_X1 U10990 ( .A1(n8138), .A2(n13614), .ZN(n8568) );
  INV_X1 U10991 ( .A(n8565), .ZN(n8563) );
  NAND2_X1 U10992 ( .A1(n8563), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n12604) );
  INV_X1 U10993 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8564) );
  NAND2_X1 U10994 ( .A1(n8565), .A2(n8564), .ZN(n8566) );
  NAND2_X1 U10995 ( .A1(n12604), .A2(n8566), .ZN(n13613) );
  OR2_X1 U10996 ( .A1(n8137), .A2(n13613), .ZN(n8567) );
  NAND4_X1 U10997 ( .A1(n8570), .A2(n8569), .A3(n8568), .A4(n8567), .ZN(n13512) );
  NAND2_X1 U10998 ( .A1(n8579), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8573) );
  XNOR2_X1 U10999 ( .A(n8573), .B(P2_IR_REG_25__SCAN_IN), .ZN(n8584) );
  INV_X1 U11000 ( .A(n8584), .ZN(n13961) );
  INV_X1 U11001 ( .A(n8574), .ZN(n8575) );
  NAND2_X1 U11002 ( .A1(n8575), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8576) );
  MUX2_X1 U11003 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8576), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8577) );
  NAND2_X1 U11004 ( .A1(n8577), .A2(n8579), .ZN(n13968) );
  XNOR2_X1 U11005 ( .A(n13968), .B(P2_B_REG_SCAN_IN), .ZN(n8578) );
  NAND2_X1 U11006 ( .A1(n13961), .A2(n8578), .ZN(n8581) );
  INV_X1 U11007 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15489) );
  NAND2_X1 U11008 ( .A1(n15205), .A2(n15489), .ZN(n8583) );
  OR2_X1 U11009 ( .A1(n13957), .A2(n8584), .ZN(n8582) );
  NAND2_X1 U11010 ( .A1(n8583), .A2(n8582), .ZN(n9797) );
  INV_X1 U11011 ( .A(n9797), .ZN(n8613) );
  INV_X1 U11012 ( .A(n13968), .ZN(n8589) );
  NAND3_X1 U11013 ( .A1(n13957), .A2(n8589), .A3(n8584), .ZN(n10413) );
  INV_X1 U11014 ( .A(n8585), .ZN(n8586) );
  NAND2_X1 U11015 ( .A1(n8586), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8588) );
  AND2_X1 U11016 ( .A1(n10413), .A2(n10416), .ZN(n8615) );
  NAND2_X1 U11017 ( .A1(n8613), .A2(n15210), .ZN(n11756) );
  INV_X1 U11018 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15208) );
  NAND2_X1 U11019 ( .A1(n15205), .A2(n15208), .ZN(n8591) );
  OR2_X1 U11020 ( .A1(n8589), .A2(n13957), .ZN(n8590) );
  NAND2_X1 U11021 ( .A1(n8591), .A2(n8590), .ZN(n15209) );
  NOR2_X1 U11022 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .ZN(
        n15723) );
  NOR4_X1 U11023 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8594) );
  NOR4_X1 U11024 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8593) );
  NOR4_X1 U11025 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n8592) );
  AND4_X1 U11026 ( .A1(n15723), .A2(n8594), .A3(n8593), .A4(n8592), .ZN(n8600)
         );
  NOR4_X1 U11027 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n8598) );
  NOR4_X1 U11028 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n8597) );
  NOR4_X1 U11029 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n8596) );
  NOR4_X1 U11030 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n8595) );
  AND4_X1 U11031 ( .A1(n8598), .A2(n8597), .A3(n8596), .A4(n8595), .ZN(n8599)
         );
  NAND2_X1 U11032 ( .A1(n8600), .A2(n8599), .ZN(n8601) );
  NAND2_X1 U11033 ( .A1(n15205), .A2(n8601), .ZN(n11754) );
  NAND2_X1 U11034 ( .A1(n11196), .A2(n11754), .ZN(n8602) );
  OR2_X1 U11035 ( .A1(n11756), .A2(n8602), .ZN(n8618) );
  AND2_X2 U11036 ( .A1(n8604), .A2(n9664), .ZN(n15251) );
  INV_X1 U11037 ( .A(n10415), .ZN(n8605) );
  NAND2_X1 U11038 ( .A1(n15263), .A2(n8605), .ZN(n8606) );
  NOR2_X1 U11039 ( .A1(n13481), .A2(n13690), .ZN(n13496) );
  INV_X1 U11040 ( .A(n13512), .ZN(n9735) );
  INV_X1 U11041 ( .A(n8609), .ZN(n8632) );
  NOR2_X1 U11042 ( .A1(n8610), .A2(n8079), .ZN(n11769) );
  INV_X1 U11043 ( .A(n11769), .ZN(n8612) );
  NAND2_X1 U11044 ( .A1(n13690), .A2(n9698), .ZN(n9798) );
  INV_X1 U11045 ( .A(n9798), .ZN(n8611) );
  NAND3_X1 U11046 ( .A1(n11196), .A2(n8613), .A3(n11754), .ZN(n8614) );
  NAND2_X1 U11047 ( .A1(n8614), .A2(n9798), .ZN(n8617) );
  NAND2_X1 U11048 ( .A1(n10415), .A2(n9664), .ZN(n11753) );
  AND2_X1 U11049 ( .A1(n8615), .A2(n11753), .ZN(n8616) );
  NAND2_X1 U11050 ( .A1(n8617), .A2(n8616), .ZN(n11348) );
  NOR2_X2 U11051 ( .A1(n8618), .A2(n9664), .ZN(n14845) );
  NAND2_X1 U11052 ( .A1(n9613), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8624) );
  INV_X1 U11053 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8619) );
  OR2_X1 U11054 ( .A1(n8139), .A2(n8619), .ZN(n8623) );
  INV_X1 U11055 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8620) );
  OR2_X1 U11056 ( .A1(n8138), .A2(n8620), .ZN(n8622) );
  OR2_X1 U11057 ( .A1(n8137), .A2(n12604), .ZN(n8621) );
  NAND4_X1 U11058 ( .A1(n8624), .A2(n8623), .A3(n8622), .A4(n8621), .ZN(n13511) );
  AND2_X2 U11059 ( .A1(n10415), .A2(n8625), .ZN(n13816) );
  NAND2_X1 U11060 ( .A1(n13511), .A2(n13816), .ZN(n8627) );
  INV_X1 U11061 ( .A(n8625), .ZN(n10419) );
  AND2_X2 U11062 ( .A1(n10415), .A2(n10419), .ZN(n13814) );
  NAND2_X1 U11063 ( .A1(n13637), .A2(n13814), .ZN(n8626) );
  NAND2_X1 U11064 ( .A1(n8627), .A2(n8626), .ZN(n13607) );
  AOI22_X1 U11065 ( .A1(n14845), .A2(n13607), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n8628) );
  OAI21_X1 U11066 ( .B1(n13613), .B2(n15124), .A(n8628), .ZN(n8629) );
  AOI21_X1 U11067 ( .B1(n13843), .B2(n13506), .A(n8629), .ZN(n8630) );
  INV_X1 U11068 ( .A(n8630), .ZN(n8631) );
  AOI21_X1 U11069 ( .B1(n8633), .B2(n8632), .A(n8631), .ZN(n8634) );
  NAND2_X1 U11070 ( .A1(n8635), .A2(n8634), .ZN(P2_U3192) );
  INV_X1 U11071 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n9186) );
  NOR2_X1 U11072 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), 
        .ZN(n8637) );
  XNOR2_X2 U11073 ( .A(n8650), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8651) );
  INV_X1 U11074 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10756) );
  INV_X1 U11075 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10757) );
  NAND2_X2 U11076 ( .A1(n8652), .A2(n8651), .ZN(n8700) );
  INV_X1 U11077 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11396) );
  INV_X1 U11078 ( .A(n8656), .ZN(n8659) );
  NAND2_X1 U11079 ( .A1(n8663), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8665) );
  NAND2_X1 U11080 ( .A1(n8664), .A2(n8665), .ZN(n8668) );
  INV_X1 U11081 ( .A(n8665), .ZN(n8666) );
  NAND2_X1 U11082 ( .A1(n8667), .A2(n8666), .ZN(n8684) );
  AND2_X1 U11083 ( .A1(n8668), .A2(n8684), .ZN(n10467) );
  NAND2_X1 U11084 ( .A1(n8702), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8673) );
  INV_X1 U11085 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n15714) );
  OR2_X1 U11086 ( .A1(n8700), .A2(n15714), .ZN(n8672) );
  INV_X1 U11087 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10762) );
  OR2_X1 U11088 ( .A1(n6547), .A2(n10762), .ZN(n8671) );
  INV_X1 U11089 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10763) );
  OR2_X1 U11090 ( .A1(n8699), .A2(n10763), .ZN(n8670) );
  INV_X1 U11091 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9898) );
  XNOR2_X1 U11092 ( .A(n9898), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8674) );
  MUX2_X1 U11093 ( .A(n8674), .B(SI_0_), .S(n10486), .Z(n10464) );
  MUX2_X1 U11094 ( .A(P3_IR_REG_0__SCAN_IN), .B(n10464), .S(n8675), .Z(n11365)
         );
  INV_X1 U11095 ( .A(n9116), .ZN(n15357) );
  NAND2_X1 U11096 ( .A1(n15362), .A2(n9267), .ZN(n15342) );
  NAND2_X1 U11097 ( .A1(n8702), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8679) );
  INV_X1 U11098 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10765) );
  OR2_X1 U11099 ( .A1(n6547), .A2(n10765), .ZN(n8678) );
  INV_X1 U11100 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n11286) );
  OR2_X1 U11101 ( .A1(n8700), .A2(n11286), .ZN(n8677) );
  INV_X1 U11102 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10766) );
  OR2_X1 U11103 ( .A1(n8699), .A2(n10766), .ZN(n8676) );
  INV_X1 U11104 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8681) );
  INV_X1 U11105 ( .A(n14753), .ZN(n10777) );
  NAND2_X1 U11106 ( .A1(n10488), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8683) );
  XNOR2_X1 U11107 ( .A(n8695), .B(n8694), .ZN(n14751) );
  OR2_X1 U11108 ( .A1(n8994), .A2(n14751), .ZN(n8686) );
  OR2_X1 U11109 ( .A1(n8722), .A2(SI_2_), .ZN(n8685) );
  NAND2_X1 U11110 ( .A1(n15340), .A2(n9253), .ZN(n11991) );
  INV_X1 U11111 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10875) );
  OR2_X1 U11112 ( .A1(n6547), .A2(n10875), .ZN(n8689) );
  OR2_X1 U11113 ( .A1(n8700), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8688) );
  INV_X1 U11114 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10876) );
  OR2_X1 U11115 ( .A1(n8699), .A2(n10876), .ZN(n8687) );
  INV_X1 U11116 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8693) );
  OR3_X1 U11117 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n8691) );
  NAND2_X1 U11118 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n8691), .ZN(n8692) );
  XNOR2_X1 U11119 ( .A(n8693), .B(n8692), .ZN(n14750) );
  XNOR2_X1 U11120 ( .A(n8710), .B(n8709), .ZN(n14748) );
  OR2_X1 U11121 ( .A1(n8994), .A2(n14748), .ZN(n8697) );
  OR2_X1 U11122 ( .A1(n8722), .A2(SI_3_), .ZN(n8696) );
  OAI211_X1 U11123 ( .C1(n10888), .C2(n10733), .A(n8697), .B(n8696), .ZN(
        n11999) );
  NAND2_X1 U11124 ( .A1(n15343), .A2(n11999), .ZN(n9263) );
  NAND2_X1 U11125 ( .A1(n11991), .A2(n11992), .ZN(n8698) );
  NAND2_X1 U11126 ( .A1(n8698), .A2(n9264), .ZN(n11421) );
  NAND2_X1 U11127 ( .A1(n9203), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8706) );
  INV_X1 U11128 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10921) );
  OR2_X1 U11129 ( .A1(n6547), .A2(n10921), .ZN(n8705) );
  AND2_X1 U11130 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8701) );
  NOR2_X1 U11131 ( .A1(n8716), .A2(n8701), .ZN(n12136) );
  OR2_X1 U11132 ( .A1(n8700), .A2(n12136), .ZN(n8704) );
  INV_X1 U11133 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8703) );
  NOR2_X1 U11134 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n8707) );
  OR2_X1 U11135 ( .A1(n8722), .A2(SI_4_), .ZN(n8713) );
  NAND2_X1 U11136 ( .A1(n10493), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8711) );
  XNOR2_X1 U11137 ( .A(n8724), .B(n8723), .ZN(n10477) );
  OR2_X1 U11138 ( .A1(n8994), .A2(n10477), .ZN(n8712) );
  NAND2_X1 U11139 ( .A1(n15421), .A2(n12137), .ZN(n8714) );
  INV_X1 U11140 ( .A(n11423), .ZN(n11420) );
  NAND2_X1 U11141 ( .A1(n11421), .A2(n11420), .ZN(n11689) );
  NAND2_X1 U11142 ( .A1(n8702), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8721) );
  INV_X1 U11143 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10911) );
  OR2_X1 U11144 ( .A1(n8699), .A2(n10911), .ZN(n8720) );
  INV_X1 U11145 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10910) );
  OR2_X1 U11146 ( .A1(n6547), .A2(n10910), .ZN(n8719) );
  NAND2_X1 U11147 ( .A1(n8716), .A2(n8715), .ZN(n8736) );
  OR2_X1 U11148 ( .A1(n8716), .A2(n8715), .ZN(n8717) );
  AND2_X1 U11149 ( .A1(n8736), .A2(n8717), .ZN(n11744) );
  OR2_X1 U11150 ( .A1(n8700), .A2(n11744), .ZN(n8718) );
  NAND4_X1 U11151 ( .A1(n8721), .A2(n8720), .A3(n8719), .A4(n8718), .ZN(n11983) );
  OR2_X1 U11152 ( .A1(n8722), .A2(SI_5_), .ZN(n8733) );
  NAND2_X1 U11153 ( .A1(n10497), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8725) );
  XNOR2_X1 U11154 ( .A(n8744), .B(n8743), .ZN(n10475) );
  OR2_X1 U11155 ( .A1(n8994), .A2(n10475), .ZN(n8732) );
  NOR2_X1 U11156 ( .A1(n8729), .A2(n8660), .ZN(n8726) );
  MUX2_X1 U11157 ( .A(n8660), .B(n8726), .S(P3_IR_REG_5__SCAN_IN), .Z(n8727)
         );
  INV_X1 U11158 ( .A(n8727), .ZN(n8730) );
  INV_X1 U11159 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8728) );
  NAND2_X1 U11160 ( .A1(n8729), .A2(n8728), .ZN(n8757) );
  NAND2_X1 U11161 ( .A1(n8730), .A2(n8757), .ZN(n10925) );
  NAND2_X1 U11162 ( .A1(n7522), .A2(n10925), .ZN(n8731) );
  XNOR2_X1 U11163 ( .A(n11983), .B(n11746), .ZN(n11697) );
  INV_X1 U11164 ( .A(n11691), .ZN(n8735) );
  INV_X1 U11165 ( .A(n11746), .ZN(n9281) );
  NOR2_X1 U11166 ( .A1(n11983), .A2(n9281), .ZN(n8734) );
  NAND2_X1 U11167 ( .A1(n9203), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8742) );
  INV_X1 U11168 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11209) );
  OR2_X1 U11169 ( .A1(n6547), .A2(n11209), .ZN(n8741) );
  NAND2_X1 U11170 ( .A1(n8736), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8737) );
  AND2_X1 U11171 ( .A1(n8751), .A2(n8737), .ZN(n12143) );
  OR2_X1 U11172 ( .A1(n8700), .A2(n12143), .ZN(n8740) );
  INV_X1 U11173 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n8738) );
  OR2_X1 U11174 ( .A1(n9080), .A2(n8738), .ZN(n8739) );
  INV_X1 U11175 ( .A(SI_6_), .ZN(n14742) );
  OR2_X1 U11176 ( .A1(n8722), .A2(n14742), .ZN(n8750) );
  NAND2_X1 U11177 ( .A1(n10490), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8745) );
  XNOR2_X1 U11178 ( .A(n10499), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8746) );
  XNOR2_X1 U11179 ( .A(n8760), .B(n8746), .ZN(n14744) );
  OR2_X1 U11180 ( .A1(n8994), .A2(n14744), .ZN(n8749) );
  NAND2_X1 U11181 ( .A1(n8757), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8747) );
  NAND2_X1 U11182 ( .A1(n7522), .A2(n11210), .ZN(n8748) );
  NAND2_X1 U11183 ( .A1(n15331), .A2(n12144), .ZN(n9284) );
  NAND2_X1 U11184 ( .A1(n9286), .A2(n9284), .ZN(n11709) );
  INV_X1 U11185 ( .A(n11709), .ZN(n11706) );
  NAND2_X1 U11186 ( .A1(n8702), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8756) );
  INV_X1 U11187 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11217) );
  OR2_X1 U11188 ( .A1(n6547), .A2(n11217), .ZN(n8755) );
  AND2_X1 U11189 ( .A1(n8751), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8752) );
  NOR2_X1 U11190 ( .A1(n8764), .A2(n8752), .ZN(n15325) );
  OR2_X1 U11191 ( .A1(n8700), .A2(n15325), .ZN(n8754) );
  INV_X1 U11192 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11218) );
  OR2_X1 U11193 ( .A1(n8699), .A2(n11218), .ZN(n8753) );
  OAI21_X1 U11194 ( .B1(n8757), .B2(P3_IR_REG_6__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8758) );
  XNOR2_X1 U11195 ( .A(n8758), .B(P3_IR_REG_7__SCAN_IN), .ZN(n11219) );
  OR2_X1 U11196 ( .A1(n8722), .A2(SI_7_), .ZN(n8763) );
  NAND2_X1 U11197 ( .A1(n10504), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8761) );
  XNOR2_X1 U11198 ( .A(n8778), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n8775) );
  XNOR2_X1 U11199 ( .A(n8777), .B(n8775), .ZN(n10473) );
  OR2_X1 U11200 ( .A1(n8994), .A2(n10473), .ZN(n8762) );
  OAI211_X1 U11201 ( .C1(n11219), .C2(n10733), .A(n8763), .B(n8762), .ZN(
        n15324) );
  OR2_X1 U11202 ( .A1(n15310), .A2(n15324), .ZN(n9288) );
  NAND2_X1 U11203 ( .A1(n15310), .A2(n15324), .ZN(n9287) );
  INV_X1 U11204 ( .A(n15328), .ZN(n15321) );
  NAND2_X1 U11205 ( .A1(n9203), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8771) );
  NOR2_X1 U11206 ( .A1(n8764), .A2(n11556), .ZN(n8765) );
  OR2_X1 U11207 ( .A1(n8783), .A2(n8765), .ZN(n15313) );
  INV_X1 U11208 ( .A(n15313), .ZN(n8766) );
  OR2_X1 U11209 ( .A1(n8700), .A2(n8766), .ZN(n8770) );
  INV_X1 U11210 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n8767) );
  OR2_X1 U11211 ( .A1(n9080), .A2(n8767), .ZN(n8769) );
  INV_X1 U11212 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11559) );
  OR2_X1 U11213 ( .A1(n6547), .A2(n11559), .ZN(n8768) );
  NAND4_X1 U11214 ( .A1(n8771), .A2(n8770), .A3(n8769), .A4(n8768), .ZN(n15330) );
  NAND2_X1 U11215 ( .A1(n8772), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8773) );
  OR2_X1 U11216 ( .A1(n8772), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8790) );
  NAND2_X1 U11217 ( .A1(n8774), .A2(n8790), .ZN(n11869) );
  INV_X1 U11218 ( .A(SI_8_), .ZN(n10469) );
  OR2_X1 U11219 ( .A1(n8722), .A2(n10469), .ZN(n8781) );
  INV_X1 U11220 ( .A(n8775), .ZN(n8776) );
  NAND2_X1 U11221 ( .A1(n8778), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8779) );
  XNOR2_X1 U11222 ( .A(n8795), .B(n8794), .ZN(n10468) );
  OR2_X1 U11223 ( .A1(n8994), .A2(n10468), .ZN(n8780) );
  OAI211_X1 U11224 ( .C1(n10733), .C2(n11869), .A(n8781), .B(n8780), .ZN(
        n12198) );
  XNOR2_X1 U11225 ( .A(n15330), .B(n12198), .ZN(n15315) );
  INV_X1 U11226 ( .A(n12198), .ZN(n15317) );
  OR2_X1 U11227 ( .A1(n15330), .A2(n15317), .ZN(n9293) );
  NAND2_X1 U11228 ( .A1(n8702), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8788) );
  OR2_X1 U11229 ( .A1(n8783), .A2(n8782), .ZN(n8784) );
  AND2_X1 U11230 ( .A1(n8801), .A2(n8784), .ZN(n15301) );
  OR2_X1 U11231 ( .A1(n8700), .A2(n15301), .ZN(n8787) );
  INV_X1 U11232 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11862) );
  OR2_X1 U11233 ( .A1(n8699), .A2(n11862), .ZN(n8786) );
  INV_X1 U11234 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11861) );
  OR2_X1 U11235 ( .A1(n6547), .A2(n11861), .ZN(n8785) );
  NAND4_X1 U11236 ( .A1(n8788), .A2(n8787), .A3(n8786), .A4(n8785), .ZN(n15311) );
  NAND2_X1 U11237 ( .A1(n8790), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8789) );
  INV_X1 U11238 ( .A(n8790), .ZN(n8792) );
  NAND2_X1 U11239 ( .A1(n8792), .A2(n8791), .ZN(n8911) );
  NAND2_X1 U11240 ( .A1(n8793), .A2(n8911), .ZN(n11873) );
  OR2_X1 U11241 ( .A1(n8722), .A2(SI_9_), .ZN(n8799) );
  NAND2_X1 U11242 ( .A1(n8795), .A2(n8794), .ZN(n8797) );
  NAND2_X1 U11243 ( .A1(n8796), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n15707) );
  XNOR2_X1 U11244 ( .A(n10519), .B(P1_DATAO_REG_9__SCAN_IN), .ZN(n8809) );
  XNOR2_X1 U11245 ( .A(n8811), .B(n8809), .ZN(n10471) );
  OR2_X1 U11246 ( .A1(n8994), .A2(n10471), .ZN(n8798) );
  OAI211_X1 U11247 ( .C1(n11913), .C2(n10733), .A(n8799), .B(n8798), .ZN(
        n15304) );
  NAND2_X1 U11248 ( .A1(n15311), .A2(n15304), .ZN(n9296) );
  OR2_X1 U11249 ( .A1(n15311), .A2(n15304), .ZN(n9297) );
  NAND2_X1 U11250 ( .A1(n8702), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8807) );
  INV_X1 U11251 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n8800) );
  OR2_X1 U11252 ( .A1(n6547), .A2(n8800), .ZN(n8806) );
  NAND2_X1 U11253 ( .A1(n8801), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8802) );
  AND2_X1 U11254 ( .A1(n8817), .A2(n8802), .ZN(n15288) );
  OR2_X1 U11255 ( .A1(n8700), .A2(n15288), .ZN(n8805) );
  INV_X1 U11256 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n8803) );
  OR2_X1 U11257 ( .A1(n8699), .A2(n8803), .ZN(n8804) );
  NAND4_X1 U11258 ( .A1(n8807), .A2(n8806), .A3(n8805), .A4(n8804), .ZN(n14810) );
  NAND2_X1 U11259 ( .A1(n8911), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8808) );
  XNOR2_X1 U11260 ( .A(n8808), .B(n8835), .ZN(n14756) );
  INV_X1 U11261 ( .A(n14756), .ZN(n12351) );
  INV_X1 U11262 ( .A(n8809), .ZN(n8810) );
  NAND2_X1 U11263 ( .A1(n10519), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8812) );
  XNOR2_X1 U11264 ( .A(n10566), .B(P1_DATAO_REG_10__SCAN_IN), .ZN(n8824) );
  XNOR2_X1 U11265 ( .A(n8826), .B(n8824), .ZN(n14754) );
  OR2_X1 U11266 ( .A1(n8994), .A2(n14754), .ZN(n8814) );
  OR2_X1 U11267 ( .A1(n8722), .A2(SI_10_), .ZN(n8813) );
  OAI211_X1 U11268 ( .C1(n12351), .C2(n10733), .A(n8814), .B(n8813), .ZN(
        n15287) );
  OR2_X1 U11269 ( .A1(n14810), .A2(n15287), .ZN(n9301) );
  NAND2_X1 U11270 ( .A1(n14810), .A2(n15287), .ZN(n9302) );
  NAND2_X1 U11271 ( .A1(n9301), .A2(n9302), .ZN(n15283) );
  NAND2_X1 U11272 ( .A1(n8702), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8823) );
  INV_X1 U11273 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n8816) );
  OR2_X1 U11274 ( .A1(n6547), .A2(n8816), .ZN(n8822) );
  NAND2_X1 U11275 ( .A1(n8817), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8818) );
  AND2_X1 U11276 ( .A1(n8842), .A2(n8818), .ZN(n12335) );
  OR2_X1 U11277 ( .A1(n8700), .A2(n12335), .ZN(n8821) );
  INV_X1 U11278 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n8819) );
  OR2_X1 U11279 ( .A1(n8699), .A2(n8819), .ZN(n8820) );
  NAND4_X1 U11280 ( .A1(n8823), .A2(n8822), .A3(n8821), .A4(n8820), .ZN(n15282) );
  INV_X1 U11281 ( .A(n8824), .ZN(n8825) );
  XNOR2_X1 U11282 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8827) );
  XNOR2_X1 U11283 ( .A(n8832), .B(n8827), .ZN(n14757) );
  NAND2_X1 U11284 ( .A1(n14757), .A2(n9234), .ZN(n8830) );
  OAI21_X1 U11285 ( .B1(n8911), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8828) );
  XNOR2_X1 U11286 ( .A(n8828), .B(n8834), .ZN(n14760) );
  NAND2_X1 U11287 ( .A1(n7522), .A2(n14760), .ZN(n8829) );
  OAI211_X1 U11288 ( .C1(SI_11_), .C2(n8722), .A(n8830), .B(n8829), .ZN(n14818) );
  OR2_X1 U11289 ( .A1(n15282), .A2(n14818), .ZN(n9300) );
  NAND2_X1 U11290 ( .A1(n15282), .A2(n14818), .ZN(n9308) );
  NAND2_X1 U11291 ( .A1(n9300), .A2(n9308), .ZN(n14814) );
  NAND2_X1 U11292 ( .A1(n15628), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8851) );
  NAND2_X1 U11293 ( .A1(n15461), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8833) );
  XNOR2_X1 U11294 ( .A(n8850), .B(n8848), .ZN(n14763) );
  NAND2_X1 U11295 ( .A1(n14763), .A2(n9234), .ZN(n8839) );
  NAND2_X1 U11296 ( .A1(n8835), .A2(n8834), .ZN(n8836) );
  NOR2_X1 U11297 ( .A1(n8911), .A2(n8836), .ZN(n8856) );
  OR2_X1 U11298 ( .A1(n8856), .A2(n8660), .ZN(n8837) );
  XNOR2_X1 U11299 ( .A(n8837), .B(P3_IR_REG_12__SCAN_IN), .ZN(n12396) );
  AOI22_X1 U11300 ( .A1(n9216), .A2(SI_12_), .B1(n7522), .B2(n12396), .ZN(
        n8838) );
  NAND2_X1 U11301 ( .A1(n8702), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8847) );
  INV_X1 U11302 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12365) );
  OR2_X1 U11303 ( .A1(n8699), .A2(n12365), .ZN(n8846) );
  INV_X1 U11304 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n8840) );
  OR2_X1 U11305 ( .A1(n6547), .A2(n8840), .ZN(n8845) );
  NAND2_X1 U11306 ( .A1(n8842), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8843) );
  AND2_X1 U11307 ( .A1(n8866), .A2(n8843), .ZN(n12411) );
  OR2_X1 U11308 ( .A1(n8700), .A2(n12411), .ZN(n8844) );
  NAND4_X1 U11309 ( .A1(n8847), .A2(n8846), .A3(n8845), .A4(n8844), .ZN(n14809) );
  NAND2_X1 U11310 ( .A1(n12409), .A2(n14809), .ZN(n9310) );
  NAND2_X1 U11311 ( .A1(n9313), .A2(n9310), .ZN(n9392) );
  INV_X1 U11312 ( .A(n9392), .ZN(n12367) );
  NAND2_X1 U11313 ( .A1(n8853), .A2(n15654), .ZN(n8854) );
  NAND2_X1 U11314 ( .A1(n8873), .A2(n8854), .ZN(n10559) );
  NAND2_X1 U11315 ( .A1(n10559), .A2(n9234), .ZN(n8861) );
  INV_X1 U11316 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8855) );
  NAND2_X1 U11317 ( .A1(n8856), .A2(n8855), .ZN(n8858) );
  NAND2_X1 U11318 ( .A1(n8858), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8857) );
  MUX2_X1 U11319 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8857), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n8859) );
  NAND2_X1 U11320 ( .A1(n8859), .A2(n8890), .ZN(n12924) );
  AOI22_X1 U11321 ( .A1(n9216), .A2(n10560), .B1(n7522), .B2(n12924), .ZN(
        n8860) );
  NAND2_X1 U11322 ( .A1(n8702), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8871) );
  INV_X1 U11323 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n8862) );
  OR2_X1 U11324 ( .A1(n8699), .A2(n8862), .ZN(n8870) );
  INV_X1 U11325 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n8863) );
  OR2_X1 U11326 ( .A1(n6547), .A2(n8863), .ZN(n8869) );
  NAND2_X1 U11327 ( .A1(n8866), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8867) );
  AND2_X1 U11328 ( .A1(n8881), .A2(n8867), .ZN(n12464) );
  OR2_X1 U11329 ( .A1(n8700), .A2(n12464), .ZN(n8868) );
  NOR2_X1 U11330 ( .A1(n14821), .A2(n12901), .ZN(n9314) );
  NAND2_X1 U11331 ( .A1(n14821), .A2(n12901), .ZN(n9312) );
  NAND2_X1 U11332 ( .A1(n11088), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8887) );
  NAND2_X1 U11333 ( .A1(n15544), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8874) );
  OAI21_X1 U11334 ( .B1(n8876), .B2(n8875), .A(n7223), .ZN(n10617) );
  NAND2_X1 U11335 ( .A1(n10617), .A2(n9234), .ZN(n8880) );
  NAND2_X1 U11336 ( .A1(n8890), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8878) );
  XNOR2_X1 U11337 ( .A(n8878), .B(n8877), .ZN(n12954) );
  AOI22_X1 U11338 ( .A1(n9216), .A2(n10618), .B1(n7522), .B2(n12954), .ZN(
        n8879) );
  NAND2_X1 U11339 ( .A1(n9203), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8886) );
  INV_X1 U11340 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13315) );
  OR2_X1 U11341 ( .A1(n6547), .A2(n13315), .ZN(n8885) );
  NAND2_X1 U11342 ( .A1(n8881), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8882) );
  AND2_X1 U11343 ( .A1(n8896), .A2(n8882), .ZN(n12530) );
  OR2_X1 U11344 ( .A1(n8700), .A2(n12530), .ZN(n8884) );
  INV_X1 U11345 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13373) );
  OR2_X1 U11346 ( .A1(n9080), .A2(n13373), .ZN(n8883) );
  NAND4_X1 U11347 ( .A1(n8886), .A2(n8885), .A3(n8884), .A4(n8883), .ZN(n12900) );
  OR2_X1 U11348 ( .A1(n13375), .A2(n12900), .ZN(n9321) );
  NAND2_X1 U11349 ( .A1(n13375), .A2(n12900), .ZN(n9320) );
  NAND2_X1 U11350 ( .A1(n11240), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8905) );
  NAND2_X1 U11351 ( .A1(n11238), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8889) );
  NAND2_X1 U11352 ( .A1(n8905), .A2(n8889), .ZN(n8902) );
  XNOR2_X1 U11353 ( .A(n8904), .B(n8902), .ZN(n10779) );
  NAND2_X1 U11354 ( .A1(n10779), .A2(n9234), .ZN(n8893) );
  OAI21_X1 U11355 ( .B1(n8890), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8891) );
  XNOR2_X1 U11356 ( .A(n8891), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12977) );
  AOI22_X1 U11357 ( .A1(n9216), .A2(SI_15_), .B1(n7522), .B2(n12977), .ZN(
        n8892) );
  NAND2_X1 U11358 ( .A1(n8702), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8901) );
  INV_X1 U11359 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n15480) );
  OR2_X1 U11360 ( .A1(n6547), .A2(n15480), .ZN(n8900) );
  INV_X1 U11361 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13251) );
  OR2_X1 U11362 ( .A1(n8699), .A2(n13251), .ZN(n8899) );
  NAND2_X1 U11363 ( .A1(n8896), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8897) );
  AND2_X1 U11364 ( .A1(n8916), .A2(n8897), .ZN(n13250) );
  OR2_X1 U11365 ( .A1(n8700), .A2(n13250), .ZN(n8898) );
  NAND4_X1 U11366 ( .A1(n8901), .A2(n8900), .A3(n8899), .A4(n8898), .ZN(n12899) );
  OR2_X1 U11367 ( .A1(n13248), .A2(n13231), .ZN(n9324) );
  NAND2_X1 U11368 ( .A1(n13248), .A2(n13231), .ZN(n9329) );
  INV_X1 U11369 ( .A(n8902), .ZN(n8903) );
  NAND2_X1 U11370 ( .A1(n15512), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8922) );
  NAND2_X1 U11371 ( .A1(n11183), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8906) );
  OR2_X1 U11372 ( .A1(n8908), .A2(n8907), .ZN(n8909) );
  AND2_X1 U11373 ( .A1(n8923), .A2(n8909), .ZN(n11055) );
  NAND2_X1 U11374 ( .A1(n11055), .A2(n9234), .ZN(n8915) );
  OAI21_X1 U11375 ( .B1(n8911), .B2(n8910), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8913) );
  XNOR2_X1 U11376 ( .A(n8913), .B(n8912), .ZN(n12998) );
  INV_X1 U11377 ( .A(n12998), .ZN(n12976) );
  AOI22_X1 U11378 ( .A1(n9216), .A2(SI_16_), .B1(n7522), .B2(n12976), .ZN(
        n8914) );
  NAND2_X1 U11379 ( .A1(n9224), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8921) );
  INV_X1 U11380 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13237) );
  OR2_X1 U11381 ( .A1(n8699), .A2(n13237), .ZN(n8920) );
  NAND2_X1 U11382 ( .A1(n8916), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8917) );
  AND2_X1 U11383 ( .A1(n8935), .A2(n8917), .ZN(n13236) );
  OR2_X1 U11384 ( .A1(n8700), .A2(n13236), .ZN(n8919) );
  INV_X1 U11385 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13365) );
  OR2_X1 U11386 ( .A1(n9080), .A2(n13365), .ZN(n8918) );
  NAND4_X1 U11387 ( .A1(n8921), .A2(n8920), .A3(n8919), .A4(n8918), .ZN(n12898) );
  NAND2_X1 U11388 ( .A1(n13367), .A2(n12898), .ZN(n9331) );
  NAND2_X1 U11389 ( .A1(n12841), .A2(n13245), .ZN(n9330) );
  NAND2_X1 U11390 ( .A1(n9331), .A2(n9330), .ZN(n13229) );
  INV_X1 U11391 ( .A(n13229), .ZN(n13234) );
  NAND2_X1 U11392 ( .A1(n13233), .A2(n9330), .ZN(n13221) );
  NAND2_X1 U11393 ( .A1(n8923), .A2(n8922), .ZN(n8926) );
  NAND2_X1 U11394 ( .A1(n11234), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8941) );
  NAND2_X1 U11395 ( .A1(n11236), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8924) );
  NAND2_X1 U11396 ( .A1(n8926), .A2(n8925), .ZN(n8942) );
  OR2_X1 U11397 ( .A1(n8926), .A2(n8925), .ZN(n8927) );
  AND2_X1 U11398 ( .A1(n8942), .A2(n8927), .ZN(n11173) );
  NAND2_X1 U11399 ( .A1(n11173), .A2(n9234), .ZN(n8932) );
  NAND2_X1 U11400 ( .A1(n8929), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8928) );
  INV_X1 U11401 ( .A(n8963), .ZN(n8947) );
  NAND2_X1 U11402 ( .A1(n8930), .A2(n8947), .ZN(n13007) );
  INV_X1 U11403 ( .A(n13007), .ZN(n13003) );
  AOI22_X1 U11404 ( .A1(n9216), .A2(SI_17_), .B1(n7522), .B2(n13003), .ZN(
        n8931) );
  NAND2_X1 U11405 ( .A1(n9203), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8940) );
  NAND2_X1 U11406 ( .A1(n8935), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8936) );
  AND2_X1 U11407 ( .A1(n8951), .A2(n8936), .ZN(n13222) );
  OR2_X1 U11408 ( .A1(n8700), .A2(n13222), .ZN(n8939) );
  INV_X1 U11409 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13304) );
  OR2_X1 U11410 ( .A1(n6547), .A2(n13304), .ZN(n8938) );
  INV_X1 U11411 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13361) );
  OR2_X1 U11412 ( .A1(n9080), .A2(n13361), .ZN(n8937) );
  NAND4_X1 U11413 ( .A1(n8940), .A2(n8939), .A3(n8938), .A4(n8937), .ZN(n12897) );
  NAND2_X1 U11414 ( .A1(n13363), .A2(n12897), .ZN(n9335) );
  NAND2_X1 U11415 ( .A1(n12850), .A2(n13232), .ZN(n9334) );
  NAND2_X1 U11416 ( .A1(n9335), .A2(n9334), .ZN(n13215) );
  INV_X1 U11417 ( .A(n13215), .ZN(n13220) );
  NAND2_X1 U11418 ( .A1(n8942), .A2(n8941), .ZN(n8945) );
  INV_X1 U11419 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11469) );
  NAND2_X1 U11420 ( .A1(n11469), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8957) );
  INV_X1 U11421 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11466) );
  NAND2_X1 U11422 ( .A1(n11466), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8943) );
  OR2_X1 U11423 ( .A1(n8945), .A2(n8944), .ZN(n8946) );
  NAND2_X1 U11424 ( .A1(n8958), .A2(n8946), .ZN(n11184) );
  OR2_X1 U11425 ( .A1(n11184), .A2(n8994), .ZN(n8950) );
  NAND2_X1 U11426 ( .A1(n8947), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8948) );
  XNOR2_X1 U11427 ( .A(n8948), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13030) );
  AOI22_X1 U11428 ( .A1(n9216), .A2(SI_18_), .B1(n7522), .B2(n13030), .ZN(
        n8949) );
  NAND2_X1 U11429 ( .A1(n8951), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8952) );
  NAND2_X1 U11430 ( .A1(n8972), .A2(n8952), .ZN(n13205) );
  NAND2_X1 U11431 ( .A1(n9113), .A2(n13205), .ZN(n8956) );
  INV_X1 U11432 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13207) );
  OR2_X1 U11433 ( .A1(n8699), .A2(n13207), .ZN(n8955) );
  INV_X1 U11434 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13300) );
  OR2_X1 U11435 ( .A1(n6547), .A2(n13300), .ZN(n8954) );
  INV_X1 U11436 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13357) );
  OR2_X1 U11437 ( .A1(n9080), .A2(n13357), .ZN(n8953) );
  NAND4_X1 U11438 ( .A1(n8956), .A2(n8955), .A3(n8954), .A4(n8953), .ZN(n13186) );
  NAND2_X1 U11439 ( .A1(n13359), .A2(n13186), .ZN(n9338) );
  INV_X1 U11440 ( .A(n13359), .ZN(n13210) );
  NAND2_X1 U11441 ( .A1(n13210), .A2(n13218), .ZN(n9341) );
  NAND2_X1 U11442 ( .A1(n15594), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8977) );
  INV_X1 U11443 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12650) );
  NAND2_X1 U11444 ( .A1(n12650), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8959) );
  OR2_X1 U11445 ( .A1(n8961), .A2(n8960), .ZN(n8962) );
  NAND2_X1 U11446 ( .A1(n8978), .A2(n8962), .ZN(n11232) );
  NAND2_X1 U11447 ( .A1(n11232), .A2(n9234), .ZN(n8967) );
  INV_X1 U11448 ( .A(SI_19_), .ZN(n11231) );
  INV_X1 U11449 ( .A(n9090), .ZN(n8964) );
  NAND2_X1 U11450 ( .A1(n8964), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8965) );
  AOI22_X1 U11451 ( .A1(n9216), .A2(n11231), .B1(n7522), .B2(n13033), .ZN(
        n8966) );
  INV_X1 U11452 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13032) );
  INV_X1 U11453 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13296) );
  OR2_X1 U11454 ( .A1(n6547), .A2(n13296), .ZN(n8969) );
  INV_X1 U11455 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13353) );
  OR2_X1 U11456 ( .A1(n9080), .A2(n13353), .ZN(n8968) );
  AND2_X1 U11457 ( .A1(n8969), .A2(n8968), .ZN(n8975) );
  INV_X1 U11458 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8970) );
  NAND2_X1 U11459 ( .A1(n8972), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8973) );
  NAND2_X1 U11460 ( .A1(n8981), .A2(n8973), .ZN(n13190) );
  NAND2_X1 U11461 ( .A1(n13190), .A2(n9113), .ZN(n8974) );
  NAND2_X1 U11462 ( .A1(n13355), .A2(n13172), .ZN(n9346) );
  INV_X1 U11463 ( .A(n9346), .ZN(n8976) );
  XNOR2_X1 U11464 ( .A(n8986), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n11541) );
  NAND2_X1 U11465 ( .A1(n11541), .A2(n9234), .ZN(n8980) );
  OR2_X1 U11466 ( .A1(n8722), .A2(n11543), .ZN(n8979) );
  NAND2_X1 U11467 ( .A1(n8981), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8982) );
  NAND2_X1 U11468 ( .A1(n9008), .A2(n8982), .ZN(n13176) );
  NAND2_X1 U11469 ( .A1(n13176), .A2(n9113), .ZN(n8985) );
  AOI22_X1 U11470 ( .A1(n9203), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n9224), .B2(
        P3_REG1_REG_20__SCAN_IN), .ZN(n8984) );
  NAND2_X1 U11471 ( .A1(n8702), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8983) );
  XNOR2_X1 U11472 ( .A(n13289), .B(n13156), .ZN(n13175) );
  OR2_X1 U11473 ( .A1(n13289), .A2(n13156), .ZN(n9350) );
  INV_X1 U11474 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12022) );
  NAND2_X1 U11475 ( .A1(n12022), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9005) );
  INV_X1 U11476 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12054) );
  NAND2_X1 U11477 ( .A1(n12054), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8990) );
  NAND2_X1 U11478 ( .A1(n9005), .A2(n8990), .ZN(n8991) );
  NAND2_X1 U11479 ( .A1(n8992), .A2(n8991), .ZN(n8993) );
  NAND2_X1 U11480 ( .A1(n9006), .A2(n8993), .ZN(n11602) );
  OR2_X1 U11481 ( .A1(n11602), .A2(n8994), .ZN(n8996) );
  INV_X1 U11482 ( .A(SI_21_), .ZN(n11601) );
  XNOR2_X1 U11483 ( .A(n9008), .B(P3_REG3_REG_21__SCAN_IN), .ZN(n13161) );
  NAND2_X1 U11484 ( .A1(n13161), .A2(n9113), .ZN(n9001) );
  INV_X1 U11485 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n13162) );
  NAND2_X1 U11486 ( .A1(n8702), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8998) );
  NAND2_X1 U11487 ( .A1(n9224), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8997) );
  OAI211_X1 U11488 ( .C1(n8699), .C2(n13162), .A(n8998), .B(n8997), .ZN(n8999)
         );
  INV_X1 U11489 ( .A(n8999), .ZN(n9000) );
  NAND2_X1 U11490 ( .A1(n13349), .A2(n12871), .ZN(n9002) );
  NAND2_X1 U11491 ( .A1(n13165), .A2(n9002), .ZN(n9004) );
  OR2_X1 U11492 ( .A1(n13349), .A2(n12871), .ZN(n9003) );
  NAND2_X1 U11493 ( .A1(n9004), .A2(n9003), .ZN(n13143) );
  XNOR2_X1 U11494 ( .A(n12212), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n9015) );
  XNOR2_X1 U11495 ( .A(n9016), .B(n9015), .ZN(n11685) );
  NOR2_X1 U11496 ( .A1(n8722), .A2(n8055), .ZN(n9007) );
  OAI21_X1 U11497 ( .B1(n9008), .B2(P3_REG3_REG_21__SCAN_IN), .A(
        P3_REG3_REG_22__SCAN_IN), .ZN(n9011) );
  NOR2_X1 U11498 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(P3_REG3_REG_22__SCAN_IN), 
        .ZN(n9009) );
  NAND2_X1 U11499 ( .A1(n9011), .A2(n9020), .ZN(n13145) );
  NAND2_X1 U11500 ( .A1(n13145), .A2(n9113), .ZN(n9014) );
  AOI22_X1 U11501 ( .A1(n9203), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n9224), .B2(
        P3_REG1_REG_22__SCAN_IN), .ZN(n9013) );
  INV_X1 U11502 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n15447) );
  OR2_X1 U11503 ( .A1(n9080), .A2(n15447), .ZN(n9012) );
  NAND2_X1 U11504 ( .A1(n13280), .A2(n13157), .ZN(n9358) );
  NAND2_X1 U11505 ( .A1(n12212), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n9017) );
  XNOR2_X1 U11506 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n9027) );
  XNOR2_X1 U11507 ( .A(n9028), .B(n9027), .ZN(n11974) );
  NAND2_X1 U11508 ( .A1(n11974), .A2(n9234), .ZN(n9019) );
  INV_X1 U11509 ( .A(SI_23_), .ZN(n11977) );
  OR2_X1 U11510 ( .A1(n8722), .A2(n11977), .ZN(n9018) );
  NAND2_X1 U11511 ( .A1(n9020), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9021) );
  NAND2_X1 U11512 ( .A1(n9035), .A2(n9021), .ZN(n13135) );
  NAND2_X1 U11513 ( .A1(n13135), .A2(n9113), .ZN(n9026) );
  INV_X1 U11514 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n15481) );
  NAND2_X1 U11515 ( .A1(n9203), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n9023) );
  NAND2_X1 U11516 ( .A1(n8702), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n9022) );
  OAI211_X1 U11517 ( .C1(n6547), .C2(n15481), .A(n9023), .B(n9022), .ZN(n9024)
         );
  INV_X1 U11518 ( .A(n9024), .ZN(n9025) );
  XNOR2_X1 U11519 ( .A(n12808), .B(n13141), .ZN(n13127) );
  OR2_X1 U11520 ( .A1(n12808), .A2(n12872), .ZN(n9248) );
  INV_X1 U11521 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n15676) );
  NAND2_X1 U11522 ( .A1(n15676), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9029) );
  NAND2_X1 U11523 ( .A1(n9031), .A2(n13966), .ZN(n9032) );
  XNOR2_X1 U11524 ( .A(n9043), .B(n14636), .ZN(n12206) );
  NAND2_X1 U11525 ( .A1(n12206), .A2(n9234), .ZN(n9034) );
  INV_X1 U11526 ( .A(SI_24_), .ZN(n12207) );
  NAND2_X1 U11527 ( .A1(n9035), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9036) );
  NAND2_X1 U11528 ( .A1(n9049), .A2(n9036), .ZN(n13121) );
  NAND2_X1 U11529 ( .A1(n13121), .A2(n9113), .ZN(n9042) );
  INV_X1 U11530 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n9039) );
  NAND2_X1 U11531 ( .A1(n8702), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n9038) );
  NAND2_X1 U11532 ( .A1(n9224), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9037) );
  OAI211_X1 U11533 ( .C1(n8699), .C2(n9039), .A(n9038), .B(n9037), .ZN(n9040)
         );
  INV_X1 U11534 ( .A(n9040), .ZN(n9041) );
  OR2_X1 U11535 ( .A1(n12858), .A2(n13131), .ZN(n9249) );
  NAND2_X1 U11536 ( .A1(n12858), .A2(n13131), .ZN(n9252) );
  INV_X1 U11537 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13963) );
  INV_X1 U11538 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12795) );
  AOI22_X1 U11539 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .B1(n13963), .B2(n12795), .ZN(n9044) );
  XNOR2_X1 U11540 ( .A(n9058), .B(n9044), .ZN(n12343) );
  NAND2_X1 U11541 ( .A1(n12343), .A2(n9234), .ZN(n9046) );
  INV_X1 U11542 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9047) );
  NAND2_X1 U11543 ( .A1(n9049), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9050) );
  NAND2_X1 U11544 ( .A1(n9064), .A2(n9050), .ZN(n13109) );
  NAND2_X1 U11545 ( .A1(n13109), .A2(n9113), .ZN(n9055) );
  INV_X1 U11546 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n15621) );
  NAND2_X1 U11547 ( .A1(n9203), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9052) );
  INV_X1 U11548 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n15613) );
  OR2_X1 U11549 ( .A1(n9080), .A2(n15613), .ZN(n9051) );
  OAI211_X1 U11550 ( .C1(n6547), .C2(n15621), .A(n9052), .B(n9051), .ZN(n9053)
         );
  INV_X1 U11551 ( .A(n9053), .ZN(n9054) );
  NAND2_X1 U11552 ( .A1(n12832), .A2(n13089), .ZN(n9367) );
  INV_X1 U11553 ( .A(n9367), .ZN(n9056) );
  NAND2_X1 U11554 ( .A1(n13963), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9057) );
  NAND2_X1 U11555 ( .A1(n12795), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9059) );
  AOI22_X1 U11556 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n13959), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n14632), .ZN(n9060) );
  INV_X1 U11557 ( .A(n9060), .ZN(n9061) );
  XNOR2_X1 U11558 ( .A(n9073), .B(n9061), .ZN(n12454) );
  NAND2_X1 U11559 ( .A1(n12454), .A2(n9234), .ZN(n9063) );
  NAND2_X1 U11560 ( .A1(n9064), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9065) );
  NAND2_X1 U11561 ( .A1(n9078), .A2(n9065), .ZN(n13094) );
  NAND2_X1 U11562 ( .A1(n13094), .A2(n9113), .ZN(n9070) );
  INV_X1 U11563 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n15543) );
  NAND2_X1 U11564 ( .A1(n9224), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9067) );
  NAND2_X1 U11565 ( .A1(n8702), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n9066) );
  OAI211_X1 U11566 ( .C1(n15543), .C2(n8699), .A(n9067), .B(n9066), .ZN(n9068)
         );
  INV_X1 U11567 ( .A(n9068), .ZN(n9069) );
  INV_X1 U11568 ( .A(n9243), .ZN(n9071) );
  NAND2_X1 U11569 ( .A1(n13093), .A2(n12830), .ZN(n9242) );
  AND2_X1 U11570 ( .A1(n14632), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9072) );
  NAND2_X1 U11571 ( .A1(n13959), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9074) );
  XNOR2_X1 U11572 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n9075) );
  XNOR2_X1 U11573 ( .A(n9191), .B(n9075), .ZN(n12502) );
  NAND2_X1 U11574 ( .A1(n12502), .A2(n9234), .ZN(n9077) );
  INV_X1 U11575 ( .A(SI_27_), .ZN(n12503) );
  NAND2_X1 U11576 ( .A1(n9078), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9079) );
  NAND2_X1 U11577 ( .A1(n9107), .A2(n9079), .ZN(n13082) );
  NAND2_X1 U11578 ( .A1(n13082), .A2(n9113), .ZN(n9086) );
  INV_X1 U11579 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n9083) );
  NAND2_X1 U11580 ( .A1(n9224), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9082) );
  INV_X1 U11581 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n15657) );
  OR2_X1 U11582 ( .A1(n9080), .A2(n15657), .ZN(n9081) );
  OAI211_X1 U11583 ( .C1(n8699), .C2(n9083), .A(n9082), .B(n9081), .ZN(n9084)
         );
  INV_X1 U11584 ( .A(n9084), .ZN(n9085) );
  XNOR2_X1 U11585 ( .A(n12802), .B(n13090), .ZN(n10377) );
  OR2_X1 U11586 ( .A1(n9087), .A2(n9145), .ZN(n9088) );
  NAND2_X1 U11587 ( .A1(n9196), .A2(n9088), .ZN(n13085) );
  NAND2_X1 U11588 ( .A1(n9090), .A2(n9089), .ZN(n9093) );
  NAND2_X1 U11589 ( .A1(n9095), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9091) );
  MUX2_X1 U11590 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9091), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n9092) );
  NAND2_X1 U11591 ( .A1(n9093), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9094) );
  MUX2_X1 U11592 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9094), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n9096) );
  NAND2_X1 U11593 ( .A1(n11687), .A2(n11542), .ZN(n9099) );
  NAND2_X1 U11594 ( .A1(n9097), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9098) );
  NAND2_X1 U11595 ( .A1(n9099), .A2(n11683), .ZN(n9180) );
  NAND2_X1 U11596 ( .A1(n11542), .A2(n9411), .ZN(n9100) );
  NAND2_X1 U11597 ( .A1(n9100), .A2(n13042), .ZN(n9101) );
  NAND2_X1 U11598 ( .A1(n11687), .A2(n9101), .ZN(n9102) );
  NAND2_X1 U11599 ( .A1(n9180), .A2(n9102), .ZN(n10937) );
  AND2_X1 U11600 ( .A1(n10937), .A2(n15353), .ZN(n11125) );
  NAND2_X1 U11601 ( .A1(n11542), .A2(n13033), .ZN(n11273) );
  INV_X1 U11602 ( .A(n11273), .ZN(n9410) );
  NAND2_X1 U11603 ( .A1(n11125), .A2(n9410), .ZN(n9104) );
  AND2_X1 U11604 ( .A1(n13033), .A2(n9411), .ZN(n9103) );
  NAND2_X1 U11605 ( .A1(n11274), .A2(n9103), .ZN(n9179) );
  INV_X1 U11606 ( .A(n9107), .ZN(n9106) );
  INV_X1 U11607 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n9105) );
  NAND2_X1 U11608 ( .A1(n9106), .A2(n9105), .ZN(n13054) );
  NAND2_X1 U11609 ( .A1(n9107), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9108) );
  NAND2_X1 U11610 ( .A1(n13054), .A2(n9108), .ZN(n13075) );
  INV_X1 U11611 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n9111) );
  NAND2_X1 U11612 ( .A1(n8702), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9110) );
  NAND2_X1 U11613 ( .A1(n9224), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9109) );
  OAI211_X1 U11614 ( .C1(n8699), .C2(n9111), .A(n9110), .B(n9109), .ZN(n9112)
         );
  INV_X1 U11615 ( .A(n12652), .ZN(n10735) );
  NAND2_X1 U11616 ( .A1(n10735), .A2(n10764), .ZN(n10736) );
  NAND2_X1 U11617 ( .A1(n10733), .A2(n10736), .ZN(n9114) );
  NOR2_X4 U11618 ( .A1(n11687), .A2(n11683), .ZN(n10731) );
  OAI22_X1 U11619 ( .A1(n12798), .A2(n15300), .B1(n12830), .B2(n15298), .ZN(
        n9115) );
  AOI21_X1 U11620 ( .B1(n13085), .B2(n15363), .A(n9115), .ZN(n9146) );
  OR2_X1 U11621 ( .A1(n15344), .A2(n11393), .ZN(n9117) );
  NAND2_X1 U11622 ( .A1(n11271), .A2(n9117), .ZN(n15339) );
  OR2_X1 U11623 ( .A1(n15423), .A2(n6805), .ZN(n9118) );
  INV_X1 U11624 ( .A(n11999), .ZN(n15424) );
  NAND2_X1 U11625 ( .A1(n15343), .A2(n15424), .ZN(n9120) );
  INV_X1 U11626 ( .A(n12137), .ZN(n11580) );
  NAND2_X1 U11627 ( .A1(n15421), .A2(n11580), .ZN(n9121) );
  OR2_X1 U11628 ( .A1(n11983), .A2(n11746), .ZN(n9122) );
  INV_X1 U11629 ( .A(n12144), .ZN(n11984) );
  NAND2_X1 U11630 ( .A1(n15331), .A2(n11984), .ZN(n9123) );
  NAND2_X1 U11631 ( .A1(n11708), .A2(n9123), .ZN(n15329) );
  NAND2_X1 U11632 ( .A1(n15329), .A2(n15328), .ZN(n15327) );
  INV_X1 U11633 ( .A(n15324), .ZN(n12111) );
  NAND2_X1 U11634 ( .A1(n15310), .A2(n12111), .ZN(n9124) );
  OR2_X1 U11635 ( .A1(n15330), .A2(n12198), .ZN(n9125) );
  NAND2_X1 U11636 ( .A1(n15309), .A2(n9125), .ZN(n9127) );
  NAND2_X1 U11637 ( .A1(n15330), .A2(n12198), .ZN(n9126) );
  NAND2_X1 U11638 ( .A1(n9127), .A2(n9126), .ZN(n15294) );
  XNOR2_X1 U11639 ( .A(n15311), .B(n15304), .ZN(n15295) );
  INV_X1 U11640 ( .A(n15304), .ZN(n12018) );
  INV_X1 U11641 ( .A(n15287), .ZN(n12185) );
  NAND2_X1 U11642 ( .A1(n14810), .A2(n12185), .ZN(n9128) );
  INV_X1 U11643 ( .A(n14818), .ZN(n12334) );
  INV_X1 U11644 ( .A(n12409), .ZN(n9129) );
  NAND2_X1 U11645 ( .A1(n9129), .A2(n14809), .ZN(n9130) );
  NOR2_X1 U11646 ( .A1(n14821), .A2(n12428), .ZN(n9133) );
  NAND2_X1 U11647 ( .A1(n14821), .A2(n12428), .ZN(n9132) );
  INV_X1 U11648 ( .A(n12900), .ZN(n13244) );
  OR2_X1 U11649 ( .A1(n13248), .A2(n12899), .ZN(n9134) );
  NAND2_X1 U11650 ( .A1(n13242), .A2(n9134), .ZN(n9136) );
  NAND2_X1 U11651 ( .A1(n13248), .A2(n12899), .ZN(n9135) );
  NAND2_X1 U11652 ( .A1(n9136), .A2(n9135), .ZN(n13228) );
  NAND2_X1 U11653 ( .A1(n13228), .A2(n13229), .ZN(n9138) );
  NAND2_X1 U11654 ( .A1(n12841), .A2(n12898), .ZN(n9137) );
  NAND2_X1 U11655 ( .A1(n13216), .A2(n13215), .ZN(n9140) );
  NAND2_X1 U11656 ( .A1(n12850), .A2(n12897), .ZN(n9139) );
  NAND2_X1 U11657 ( .A1(n13359), .A2(n13218), .ZN(n9141) );
  INV_X1 U11658 ( .A(n13172), .ZN(n13204) );
  OR2_X1 U11659 ( .A1(n13355), .A2(n13204), .ZN(n9142) );
  OR2_X1 U11660 ( .A1(n13349), .A2(n13171), .ZN(n9143) );
  NAND2_X1 U11661 ( .A1(n13349), .A2(n13171), .ZN(n13150) );
  NAND2_X1 U11662 ( .A1(n13147), .A2(n13157), .ZN(n9144) );
  INV_X1 U11663 ( .A(n13157), .ZN(n12896) );
  INV_X1 U11664 ( .A(n12808), .ZN(n13345) );
  NAND2_X1 U11665 ( .A1(n9368), .A2(n9367), .ZN(n13101) );
  INV_X1 U11666 ( .A(n11687), .ZN(n9261) );
  NAND2_X1 U11667 ( .A1(n9261), .A2(n11274), .ZN(n9380) );
  NAND2_X1 U11668 ( .A1(n13042), .A2(n9411), .ZN(n10397) );
  NAND2_X1 U11669 ( .A1(n11542), .A2(n13042), .ZN(n15368) );
  OR2_X1 U11670 ( .A1(n15368), .A2(n9411), .ZN(n10388) );
  INV_X1 U11671 ( .A(n10388), .ZN(n15381) );
  NAND2_X1 U11672 ( .A1(n9147), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9148) );
  INV_X1 U11673 ( .A(n9149), .ZN(n9164) );
  MUX2_X1 U11674 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9150), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n9151) );
  XNOR2_X1 U11675 ( .A(n12209), .B(P3_B_REG_SCAN_IN), .ZN(n9154) );
  INV_X1 U11676 ( .A(n9162), .ZN(n12457) );
  NAND2_X1 U11677 ( .A1(n12457), .A2(n12346), .ZN(n9155) );
  AND2_X1 U11678 ( .A1(n9156), .A2(n9155), .ZN(n13377) );
  NAND2_X1 U11679 ( .A1(n12457), .A2(n12209), .ZN(n9157) );
  NAND2_X1 U11680 ( .A1(n13377), .A2(n13379), .ZN(n10394) );
  INV_X1 U11681 ( .A(n12346), .ZN(n9160) );
  INV_X1 U11682 ( .A(n12209), .ZN(n9159) );
  NAND2_X1 U11683 ( .A1(n6723), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9163) );
  MUX2_X1 U11684 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9163), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n9165) );
  INV_X1 U11685 ( .A(n13378), .ZN(n9166) );
  NOR2_X1 U11686 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .ZN(
        n9170) );
  NOR4_X1 U11687 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_25__SCAN_IN), .ZN(n9169) );
  NOR4_X1 U11688 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .A3(
        P3_D_REG_24__SCAN_IN), .A4(P3_D_REG_29__SCAN_IN), .ZN(n9168) );
  NOR4_X1 U11689 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_20__SCAN_IN), .A4(P3_D_REG_19__SCAN_IN), .ZN(n9167) );
  NAND4_X1 U11690 ( .A1(n9170), .A2(n9169), .A3(n9168), .A4(n9167), .ZN(n9176)
         );
  NOR4_X1 U11691 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n9174) );
  NOR4_X1 U11692 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_14__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n9173) );
  NOR4_X1 U11693 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9172) );
  NOR4_X1 U11694 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n9171) );
  NAND4_X1 U11695 ( .A1(n9174), .A2(n9173), .A3(n9172), .A4(n9171), .ZN(n9175)
         );
  NOR2_X1 U11696 ( .A1(n9176), .A2(n9175), .ZN(n9177) );
  AND2_X1 U11697 ( .A1(n10950), .A2(n10399), .ZN(n9178) );
  INV_X1 U11698 ( .A(n13377), .ZN(n9184) );
  NAND2_X1 U11699 ( .A1(n10731), .A2(n11273), .ZN(n11356) );
  NAND2_X1 U11700 ( .A1(n10405), .A2(n9179), .ZN(n11360) );
  NAND2_X1 U11701 ( .A1(n11356), .A2(n11360), .ZN(n9183) );
  NAND3_X1 U11702 ( .A1(n9180), .A2(n11273), .A3(n10397), .ZN(n9181) );
  NAND2_X1 U11703 ( .A1(n9181), .A2(n10405), .ZN(n9182) );
  OAI22_X1 U11704 ( .A1(n9184), .A2(n9183), .B1(n10401), .B2(n9182), .ZN(n9185) );
  MUX2_X1 U11705 ( .A(n9186), .B(n13329), .S(n15419), .Z(n9189) );
  NAND2_X1 U11706 ( .A1(n9189), .A2(n9188), .ZN(P3_U3486) );
  INV_X1 U11707 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13956) );
  AND2_X1 U11708 ( .A1(n13956), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9190) );
  INV_X1 U11709 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12538) );
  XNOR2_X1 U11710 ( .A(n12538), .B(P1_DATAO_REG_28__SCAN_IN), .ZN(n9192) );
  XNOR2_X1 U11711 ( .A(n9198), .B(n9192), .ZN(n12651) );
  INV_X1 U11712 ( .A(SI_28_), .ZN(n12653) );
  INV_X1 U11713 ( .A(n9245), .ZN(n9195) );
  NAND2_X1 U11714 ( .A1(n12802), .A2(n13090), .ZN(n13067) );
  NAND2_X1 U11715 ( .A1(n9244), .A2(n13067), .ZN(n9194) );
  AND2_X1 U11716 ( .A1(n12538), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9197) );
  INV_X1 U11717 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n15457) );
  NAND2_X1 U11718 ( .A1(n15457), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9199) );
  INV_X1 U11719 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14628) );
  NAND2_X1 U11720 ( .A1(n14628), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n9209) );
  INV_X1 U11721 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13950) );
  NAND2_X1 U11722 ( .A1(n13950), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9200) );
  AND2_X1 U11723 ( .A1(n9209), .A2(n9200), .ZN(n9208) );
  XNOR2_X1 U11724 ( .A(n9211), .B(n9208), .ZN(n13386) );
  NAND2_X1 U11725 ( .A1(n13386), .A2(n9234), .ZN(n9202) );
  INV_X1 U11726 ( .A(SI_29_), .ZN(n13389) );
  OR2_X1 U11727 ( .A1(n8722), .A2(n13389), .ZN(n9201) );
  NAND2_X1 U11728 ( .A1(n9202), .A2(n9201), .ZN(n10393) );
  INV_X1 U11729 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n10392) );
  NAND2_X1 U11730 ( .A1(n9203), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9205) );
  NAND2_X1 U11731 ( .A1(n8702), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9204) );
  OAI211_X1 U11732 ( .C1(n10392), .C2(n6547), .A(n9205), .B(n9204), .ZN(n9206)
         );
  INV_X1 U11733 ( .A(n9206), .ZN(n9207) );
  INV_X1 U11734 ( .A(n9208), .ZN(n9210) );
  INV_X1 U11735 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n15515) );
  NAND2_X1 U11736 ( .A1(n15515), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n9213) );
  INV_X1 U11737 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13947) );
  NAND2_X1 U11738 ( .A1(n13947), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9212) );
  AND2_X1 U11739 ( .A1(n9213), .A2(n9212), .ZN(n9230) );
  NAND2_X1 U11740 ( .A1(n9231), .A2(n9230), .ZN(n9233) );
  NAND2_X1 U11741 ( .A1(n9233), .A2(n9213), .ZN(n9215) );
  XOR2_X1 U11742 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .Z(n9214) );
  XNOR2_X1 U11743 ( .A(n9215), .B(n9214), .ZN(n13381) );
  INV_X1 U11744 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n9221) );
  NAND2_X1 U11745 ( .A1(n8702), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n9220) );
  INV_X1 U11746 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n9217) );
  OR2_X1 U11747 ( .A1(n6547), .A2(n9217), .ZN(n9219) );
  OAI211_X1 U11748 ( .C1(n8699), .C2(n9221), .A(n9220), .B(n9219), .ZN(n9222)
         );
  INV_X1 U11749 ( .A(n9222), .ZN(n9223) );
  NAND2_X1 U11750 ( .A1(n9229), .A2(n9223), .ZN(n12895) );
  NAND2_X1 U11751 ( .A1(n13257), .A2(n12895), .ZN(n9382) );
  NAND2_X1 U11752 ( .A1(n10393), .A2(n13074), .ZN(n9375) );
  INV_X1 U11753 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n13058) );
  NAND2_X1 U11754 ( .A1(n8702), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9226) );
  NAND2_X1 U11755 ( .A1(n9224), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9225) );
  OAI211_X1 U11756 ( .C1(n8699), .C2(n13058), .A(n9226), .B(n9225), .ZN(n9227)
         );
  INV_X1 U11757 ( .A(n9227), .ZN(n9228) );
  INV_X1 U11758 ( .A(n12895), .ZN(n13053) );
  OR2_X1 U11759 ( .A1(n9231), .A2(n9230), .ZN(n9232) );
  AND2_X1 U11760 ( .A1(n9233), .A2(n9232), .ZN(n12655) );
  INV_X1 U11761 ( .A(SI_30_), .ZN(n15514) );
  OR2_X1 U11762 ( .A1(n8722), .A2(n15514), .ZN(n9235) );
  OAI21_X1 U11763 ( .B1(n11665), .B2(n13053), .A(n13322), .ZN(n9237) );
  NAND3_X1 U11764 ( .A1(n9382), .A2(n9375), .A3(n9237), .ZN(n9238) );
  AOI21_X1 U11765 ( .B1(n10387), .B2(n9374), .A(n9238), .ZN(n9240) );
  NOR3_X1 U11766 ( .A1(n13257), .A2(n11665), .A3(n13322), .ZN(n9239) );
  XNOR2_X1 U11767 ( .A(n9241), .B(n13042), .ZN(n9381) );
  MUX2_X1 U11768 ( .A(n9243), .B(n9242), .S(n10731), .Z(n9246) );
  INV_X1 U11769 ( .A(n13101), .ZN(n9366) );
  NAND2_X1 U11770 ( .A1(n9249), .A2(n9248), .ZN(n9250) );
  NAND2_X1 U11771 ( .A1(n9250), .A2(n9252), .ZN(n9251) );
  MUX2_X1 U11772 ( .A(n9252), .B(n9251), .S(n10405), .Z(n9365) );
  NAND2_X1 U11773 ( .A1(n9264), .A2(n9253), .ZN(n9256) );
  NAND2_X1 U11774 ( .A1(n9263), .A2(n9254), .ZN(n9255) );
  MUX2_X1 U11775 ( .A(n9256), .B(n9255), .S(n10731), .Z(n9265) );
  NAND2_X1 U11776 ( .A1(n15359), .A2(n11432), .ZN(n9384) );
  NAND2_X1 U11777 ( .A1(n9384), .A2(n9261), .ZN(n9257) );
  NAND2_X1 U11778 ( .A1(n9257), .A2(n9267), .ZN(n9259) );
  NAND2_X1 U11779 ( .A1(n9266), .A2(n9384), .ZN(n9258) );
  MUX2_X1 U11780 ( .A(n9259), .B(n9258), .S(n10731), .Z(n9260) );
  NOR2_X1 U11781 ( .A1(n9265), .A2(n9260), .ZN(n9262) );
  NAND2_X1 U11782 ( .A1(n9262), .A2(n9261), .ZN(n9274) );
  OR2_X1 U11783 ( .A1(n15359), .A2(n11432), .ZN(n11384) );
  NAND2_X1 U11784 ( .A1(n9262), .A2(n11384), .ZN(n9273) );
  MUX2_X1 U11785 ( .A(n9264), .B(n9263), .S(n10405), .Z(n9272) );
  INV_X1 U11786 ( .A(n9265), .ZN(n9270) );
  MUX2_X1 U11787 ( .A(n9267), .B(n9266), .S(n10405), .Z(n9268) );
  NAND2_X1 U11788 ( .A1(n9268), .A2(n15341), .ZN(n9269) );
  NAND2_X1 U11789 ( .A1(n9270), .A2(n9269), .ZN(n9271) );
  NAND4_X1 U11790 ( .A1(n9274), .A2(n9273), .A3(n9272), .A4(n9271), .ZN(n9275)
         );
  NAND2_X1 U11791 ( .A1(n9275), .A2(n11420), .ZN(n9277) );
  NAND3_X1 U11792 ( .A1(n15421), .A2(n12137), .A3(n10405), .ZN(n9276) );
  AOI21_X1 U11793 ( .B1(n9277), .B2(n9276), .A(n6801), .ZN(n9280) );
  AOI21_X1 U11794 ( .B1(n9278), .B2(n9286), .A(n10405), .ZN(n9279) );
  OR2_X1 U11795 ( .A1(n9280), .A2(n9279), .ZN(n9285) );
  NAND2_X1 U11796 ( .A1(n11983), .A2(n9281), .ZN(n9282) );
  AOI21_X1 U11797 ( .B1(n9284), .B2(n9282), .A(n10731), .ZN(n9283) );
  AOI21_X1 U11798 ( .B1(n9285), .B2(n9284), .A(n9283), .ZN(n9291) );
  OAI21_X1 U11799 ( .B1(n10731), .B2(n9286), .A(n15321), .ZN(n9290) );
  MUX2_X1 U11800 ( .A(n9288), .B(n9287), .S(n10405), .Z(n9289) );
  OAI211_X1 U11801 ( .C1(n9291), .C2(n9290), .A(n15315), .B(n9289), .ZN(n9295)
         );
  INV_X1 U11802 ( .A(n15295), .ZN(n15302) );
  NAND2_X1 U11803 ( .A1(n15330), .A2(n15317), .ZN(n9292) );
  MUX2_X1 U11804 ( .A(n9293), .B(n9292), .S(n10731), .Z(n9294) );
  NAND3_X1 U11805 ( .A1(n9295), .A2(n15302), .A3(n9294), .ZN(n9299) );
  NOR2_X1 U11806 ( .A1(n15283), .A2(n14814), .ZN(n9390) );
  MUX2_X1 U11807 ( .A(n9297), .B(n9296), .S(n10405), .Z(n9298) );
  NAND3_X1 U11808 ( .A1(n9299), .A2(n9390), .A3(n9298), .ZN(n9307) );
  OAI211_X1 U11809 ( .C1(n14814), .C2(n9301), .A(n9313), .B(n9300), .ZN(n9304)
         );
  NOR2_X1 U11810 ( .A1(n14814), .A2(n9302), .ZN(n9303) );
  MUX2_X1 U11811 ( .A(n9304), .B(n9303), .S(n10731), .Z(n9305) );
  INV_X1 U11812 ( .A(n9305), .ZN(n9306) );
  NAND2_X1 U11813 ( .A1(n9307), .A2(n9306), .ZN(n9311) );
  AOI21_X1 U11814 ( .B1(n9310), .B2(n9308), .A(n10405), .ZN(n9309) );
  AOI21_X1 U11815 ( .B1(n9311), .B2(n9310), .A(n9309), .ZN(n9318) );
  OR2_X1 U11816 ( .A1(n9314), .A2(n7883), .ZN(n9393) );
  INV_X1 U11817 ( .A(n9393), .ZN(n12462) );
  OAI21_X1 U11818 ( .B1(n9313), .B2(n10405), .A(n12462), .ZN(n9317) );
  MUX2_X1 U11819 ( .A(n7883), .B(n9314), .S(n10405), .Z(n9315) );
  INV_X1 U11820 ( .A(n9315), .ZN(n9316) );
  OAI21_X1 U11821 ( .B1(n9318), .B2(n9317), .A(n9316), .ZN(n9319) );
  NAND2_X1 U11822 ( .A1(n9319), .A2(n9396), .ZN(n9323) );
  MUX2_X1 U11823 ( .A(n9321), .B(n9320), .S(n10731), .Z(n9322) );
  NAND3_X1 U11824 ( .A1(n9323), .A2(n13246), .A3(n9322), .ZN(n9328) );
  NAND2_X1 U11825 ( .A1(n9331), .A2(n9324), .ZN(n9325) );
  NAND2_X1 U11826 ( .A1(n9325), .A2(n10405), .ZN(n9327) );
  INV_X1 U11827 ( .A(n9330), .ZN(n9326) );
  AOI21_X1 U11828 ( .B1(n9328), .B2(n9327), .A(n9326), .ZN(n9333) );
  AOI21_X1 U11829 ( .B1(n9330), .B2(n9329), .A(n10405), .ZN(n9332) );
  OAI22_X1 U11830 ( .A1(n9333), .A2(n9332), .B1(n9331), .B2(n10405), .ZN(n9340) );
  INV_X1 U11831 ( .A(n9334), .ZN(n9339) );
  INV_X1 U11832 ( .A(n9335), .ZN(n9336) );
  NAND2_X1 U11833 ( .A1(n9341), .A2(n9336), .ZN(n9337) );
  NAND4_X1 U11834 ( .A1(n9346), .A2(n10731), .A3(n9338), .A4(n9337), .ZN(n9343) );
  AOI22_X1 U11835 ( .A1(n9340), .A2(n13220), .B1(n9339), .B2(n9343), .ZN(n9345) );
  NAND3_X1 U11836 ( .A1(n9347), .A2(n9341), .A3(n10405), .ZN(n9342) );
  NAND2_X1 U11837 ( .A1(n9343), .A2(n9342), .ZN(n9344) );
  OAI21_X1 U11838 ( .B1(n9345), .B2(n13195), .A(n9344), .ZN(n9349) );
  INV_X1 U11839 ( .A(n13175), .ZN(n13170) );
  MUX2_X1 U11840 ( .A(n9347), .B(n9346), .S(n10405), .Z(n9348) );
  NAND3_X1 U11841 ( .A1(n9349), .A2(n13170), .A3(n9348), .ZN(n9353) );
  NAND2_X1 U11842 ( .A1(n13289), .A2(n13156), .ZN(n9351) );
  MUX2_X1 U11843 ( .A(n9351), .B(n9350), .S(n10731), .Z(n9352) );
  XNOR2_X1 U11844 ( .A(n13349), .B(n13171), .ZN(n13151) );
  NAND3_X1 U11845 ( .A1(n9353), .A2(n9352), .A3(n13151), .ZN(n9356) );
  OR3_X1 U11846 ( .A1(n13349), .A2(n12871), .A3(n10731), .ZN(n9355) );
  NAND3_X1 U11847 ( .A1(n13349), .A2(n12871), .A3(n10731), .ZN(n9354) );
  NAND4_X1 U11848 ( .A1(n9356), .A2(n13144), .A3(n9355), .A4(n9354), .ZN(n9360) );
  MUX2_X1 U11849 ( .A(n9358), .B(n9357), .S(n10731), .Z(n9359) );
  NAND3_X1 U11850 ( .A1(n9360), .A2(n13127), .A3(n9359), .ZN(n9362) );
  NAND3_X1 U11851 ( .A1(n12808), .A2(n12872), .A3(n10731), .ZN(n9361) );
  NAND2_X1 U11852 ( .A1(n9362), .A2(n9361), .ZN(n9363) );
  NAND2_X1 U11853 ( .A1(n9363), .A2(n13117), .ZN(n9364) );
  NAND3_X1 U11854 ( .A1(n9366), .A2(n9365), .A3(n9364), .ZN(n9370) );
  MUX2_X1 U11855 ( .A(n9368), .B(n9367), .S(n10405), .Z(n9369) );
  XNOR2_X1 U11856 ( .A(n13322), .B(n11665), .ZN(n9401) );
  INV_X1 U11857 ( .A(n13322), .ZN(n13261) );
  AOI21_X1 U11858 ( .B1(n13322), .B2(n10731), .A(n11665), .ZN(n9372) );
  AOI21_X1 U11859 ( .B1(n13261), .B2(n10405), .A(n9372), .ZN(n9373) );
  AOI21_X1 U11860 ( .B1(n9376), .B2(n9374), .A(n9373), .ZN(n9379) );
  INV_X1 U11861 ( .A(n9402), .ZN(n9377) );
  OAI22_X1 U11862 ( .A1(n9381), .A2(n9380), .B1(n15368), .B2(n9404), .ZN(n9409) );
  INV_X1 U11863 ( .A(n11384), .ZN(n9386) );
  INV_X1 U11864 ( .A(n9384), .ZN(n9385) );
  NOR2_X1 U11865 ( .A1(n9386), .A2(n9385), .ZN(n11127) );
  INV_X1 U11866 ( .A(n11386), .ZN(n15356) );
  NAND4_X1 U11867 ( .A1(n11127), .A2(n11420), .A3(n15356), .A4(n11992), .ZN(
        n9388) );
  NOR4_X1 U11868 ( .A1(n9388), .A2(n15328), .A3(n9387), .A4(n11709), .ZN(n9389) );
  NAND4_X1 U11869 ( .A1(n9389), .A2(n11697), .A3(n15302), .A4(n15315), .ZN(
        n9394) );
  INV_X1 U11870 ( .A(n9390), .ZN(n9391) );
  NOR4_X1 U11871 ( .A1(n9394), .A2(n9393), .A3(n9392), .A4(n9391), .ZN(n9395)
         );
  NAND4_X1 U11872 ( .A1(n13234), .A2(n13246), .A3(n9396), .A4(n9395), .ZN(
        n9397) );
  NOR4_X1 U11873 ( .A1(n13184), .A2(n13195), .A3(n13215), .A4(n9397), .ZN(
        n9398) );
  NAND4_X1 U11874 ( .A1(n13144), .A2(n9398), .A3(n13170), .A4(n13151), .ZN(
        n9399) );
  NOR4_X1 U11875 ( .A1(n13101), .A2(n7542), .A3(n6928), .A4(n9399), .ZN(n9400)
         );
  NAND2_X1 U11876 ( .A1(n11687), .A2(n11274), .ZN(n10396) );
  INV_X1 U11877 ( .A(n10933), .ZN(n9406) );
  NAND2_X1 U11878 ( .A1(n9406), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11975) );
  NAND2_X1 U11879 ( .A1(n10950), .A2(n9410), .ZN(n11281) );
  NOR3_X1 U11880 ( .A1(n15298), .A2(n12652), .A3(n11281), .ZN(n9413) );
  OAI21_X1 U11881 ( .B1(n11975), .B2(n9411), .A(P3_B_REG_SCAN_IN), .ZN(n9412)
         );
  OR2_X1 U11882 ( .A1(n9413), .A2(n9412), .ZN(n9414) );
  INV_X1 U11883 ( .A(n11758), .ZN(n9421) );
  AND3_X2 U11884 ( .A1(n9617), .A2(n9664), .A3(n9421), .ZN(n9653) );
  NAND2_X1 U11885 ( .A1(n6553), .A2(n9578), .ZN(n9416) );
  NAND2_X1 U11886 ( .A1(n9417), .A2(n9416), .ZN(n9429) );
  NAND2_X1 U11887 ( .A1(n6553), .A2(n6552), .ZN(n9419) );
  AND2_X1 U11888 ( .A1(n9419), .A2(n9418), .ZN(n9430) );
  NAND2_X1 U11889 ( .A1(n6552), .A2(n9421), .ZN(n9424) );
  NAND2_X1 U11890 ( .A1(n13527), .A2(n9420), .ZN(n9423) );
  INV_X1 U11891 ( .A(n9667), .ZN(n12211) );
  NAND2_X1 U11892 ( .A1(n9698), .A2(n12211), .ZN(n9790) );
  NAND3_X1 U11893 ( .A1(n9791), .A2(n9421), .A3(n9790), .ZN(n9422) );
  OAI211_X1 U11894 ( .C1(n13527), .C2(n9424), .A(n9423), .B(n9422), .ZN(n9425)
         );
  INV_X1 U11895 ( .A(n9425), .ZN(n9428) );
  OAI211_X1 U11896 ( .C1(n9429), .C2(n9430), .A(n9428), .B(n9427), .ZN(n9432)
         );
  NAND2_X1 U11897 ( .A1(n9432), .A2(n9431), .ZN(n9438) );
  NAND2_X1 U11898 ( .A1(n13525), .A2(n6552), .ZN(n9434) );
  NAND2_X1 U11899 ( .A1(n13922), .A2(n9578), .ZN(n9433) );
  NAND2_X1 U11900 ( .A1(n9434), .A2(n9433), .ZN(n9437) );
  AOI22_X1 U11901 ( .A1(n13525), .A2(n9578), .B1(n13922), .B2(n6552), .ZN(
        n9435) );
  AOI21_X1 U11902 ( .B1(n9438), .B2(n9437), .A(n9435), .ZN(n9436) );
  INV_X1 U11903 ( .A(n9436), .ZN(n9439) );
  NAND2_X1 U11904 ( .A1(n13524), .A2(n9578), .ZN(n9441) );
  NAND2_X1 U11905 ( .A1(n12043), .A2(n6552), .ZN(n9440) );
  NAND2_X1 U11906 ( .A1(n9441), .A2(n9440), .ZN(n9445) );
  AOI22_X1 U11907 ( .A1(n15227), .A2(n9578), .B1(n13523), .B2(n6552), .ZN(
        n9447) );
  NAND2_X1 U11908 ( .A1(n15227), .A2(n6552), .ZN(n9443) );
  NAND2_X1 U11909 ( .A1(n13523), .A2(n9578), .ZN(n9442) );
  NAND2_X1 U11910 ( .A1(n9443), .A2(n9442), .ZN(n9446) );
  AOI22_X1 U11911 ( .A1(n13524), .A2(n6552), .B1(n12043), .B2(n9578), .ZN(
        n9444) );
  NAND2_X1 U11912 ( .A1(n9447), .A2(n9446), .ZN(n9448) );
  NAND2_X1 U11913 ( .A1(n9449), .A2(n9448), .ZN(n9461) );
  NAND2_X1 U11914 ( .A1(n11837), .A2(n6552), .ZN(n9451) );
  NAND2_X1 U11915 ( .A1(n13522), .A2(n9566), .ZN(n9450) );
  NAND2_X1 U11916 ( .A1(n9451), .A2(n9450), .ZN(n9460) );
  NAND2_X1 U11917 ( .A1(n9461), .A2(n9460), .ZN(n9454) );
  INV_X1 U11918 ( .A(n13522), .ZN(n9711) );
  NAND2_X1 U11919 ( .A1(n11837), .A2(n9566), .ZN(n9452) );
  NAND2_X1 U11920 ( .A1(n9454), .A2(n9453), .ZN(n9459) );
  AND2_X1 U11921 ( .A1(n13521), .A2(n9566), .ZN(n9455) );
  AOI21_X1 U11922 ( .B1(n11815), .B2(n9632), .A(n9455), .ZN(n9463) );
  NAND2_X1 U11923 ( .A1(n11815), .A2(n9566), .ZN(n9457) );
  NAND2_X1 U11924 ( .A1(n13521), .A2(n6552), .ZN(n9456) );
  NAND2_X1 U11925 ( .A1(n9457), .A2(n9456), .ZN(n9462) );
  NAND2_X1 U11926 ( .A1(n9463), .A2(n9462), .ZN(n9458) );
  OAI211_X1 U11927 ( .C1(n9461), .C2(n9460), .A(n9459), .B(n9458), .ZN(n9466)
         );
  INV_X1 U11928 ( .A(n9462), .ZN(n9465) );
  INV_X1 U11929 ( .A(n9463), .ZN(n9464) );
  NAND2_X1 U11930 ( .A1(n15245), .A2(n9632), .ZN(n9468) );
  NAND2_X1 U11931 ( .A1(n13520), .A2(n9566), .ZN(n9467) );
  NAND2_X1 U11932 ( .A1(n9468), .A2(n9467), .ZN(n9471) );
  INV_X1 U11933 ( .A(n13520), .ZN(n11451) );
  NAND2_X1 U11934 ( .A1(n15245), .A2(n9566), .ZN(n9469) );
  NAND2_X1 U11935 ( .A1(n11611), .A2(n9566), .ZN(n9473) );
  NAND2_X1 U11936 ( .A1(n13519), .A2(n9632), .ZN(n9472) );
  NAND2_X1 U11937 ( .A1(n9473), .A2(n9472), .ZN(n9475) );
  AOI22_X1 U11938 ( .A1(n11611), .A2(n9632), .B1(n9566), .B2(n13519), .ZN(
        n9474) );
  NOR2_X1 U11939 ( .A1(n9476), .A2(n9475), .ZN(n9477) );
  NAND2_X1 U11940 ( .A1(n15252), .A2(n9632), .ZN(n9480) );
  NAND2_X1 U11941 ( .A1(n13518), .A2(n9566), .ZN(n9479) );
  NAND2_X1 U11942 ( .A1(n9480), .A2(n9479), .ZN(n9483) );
  INV_X1 U11943 ( .A(n13518), .ZN(n9716) );
  NAND2_X1 U11944 ( .A1(n15252), .A2(n9566), .ZN(n9481) );
  NAND2_X1 U11945 ( .A1(n12102), .A2(n9566), .ZN(n9485) );
  NAND2_X1 U11946 ( .A1(n13517), .A2(n9632), .ZN(n9484) );
  AOI22_X1 U11947 ( .A1(n12102), .A2(n9632), .B1(n9566), .B2(n13517), .ZN(
        n9486) );
  NAND2_X1 U11948 ( .A1(n12214), .A2(n9632), .ZN(n9488) );
  NAND2_X1 U11949 ( .A1(n15112), .A2(n9566), .ZN(n9487) );
  NAND2_X1 U11950 ( .A1(n9488), .A2(n9487), .ZN(n9492) );
  INV_X1 U11951 ( .A(n15112), .ZN(n11927) );
  NAND2_X1 U11952 ( .A1(n12214), .A2(n9655), .ZN(n9489) );
  OAI21_X1 U11953 ( .B1(n11927), .B2(n9653), .A(n9489), .ZN(n9490) );
  NAND2_X1 U11954 ( .A1(n12253), .A2(n9655), .ZN(n9494) );
  NAND2_X1 U11955 ( .A1(n13516), .A2(n9632), .ZN(n9493) );
  AOI22_X1 U11956 ( .A1(n12253), .A2(n9632), .B1(n9566), .B2(n13516), .ZN(
        n9495) );
  NAND2_X1 U11957 ( .A1(n12420), .A2(n9632), .ZN(n9497) );
  NAND2_X1 U11958 ( .A1(n15114), .A2(n9655), .ZN(n9496) );
  NAND2_X1 U11959 ( .A1(n9497), .A2(n9496), .ZN(n9500) );
  AOI22_X1 U11960 ( .A1(n12420), .A2(n9655), .B1(n15114), .B2(n9632), .ZN(
        n9498) );
  AOI21_X1 U11961 ( .B1(n9501), .B2(n9500), .A(n9498), .ZN(n9499) );
  INV_X1 U11962 ( .A(n9499), .ZN(n9504) );
  NOR2_X1 U11963 ( .A1(n9501), .A2(n9500), .ZN(n9502) );
  INV_X1 U11964 ( .A(n9502), .ZN(n9503) );
  NAND2_X1 U11965 ( .A1(n14847), .A2(n9655), .ZN(n9506) );
  NAND2_X1 U11966 ( .A1(n13815), .A2(n9632), .ZN(n9505) );
  NAND2_X1 U11967 ( .A1(n9506), .A2(n9505), .ZN(n9509) );
  INV_X1 U11968 ( .A(n13815), .ZN(n13500) );
  NAND2_X1 U11969 ( .A1(n14847), .A2(n9632), .ZN(n9507) );
  OAI21_X1 U11970 ( .B1(n13500), .B2(n9632), .A(n9507), .ZN(n9508) );
  NAND2_X1 U11971 ( .A1(n13912), .A2(n9632), .ZN(n9511) );
  NAND2_X1 U11972 ( .A1(n13796), .A2(n9655), .ZN(n9510) );
  NAND2_X1 U11973 ( .A1(n9511), .A2(n9510), .ZN(n9513) );
  AOI22_X1 U11974 ( .A1(n13912), .A2(n9566), .B1(n13796), .B2(n9632), .ZN(
        n9512) );
  NAND2_X1 U11975 ( .A1(n13907), .A2(n9655), .ZN(n9515) );
  NAND2_X1 U11976 ( .A1(n13817), .A2(n9632), .ZN(n9514) );
  NAND2_X1 U11977 ( .A1(n9520), .A2(n9521), .ZN(n9519) );
  NAND2_X1 U11978 ( .A1(n13907), .A2(n9632), .ZN(n9517) );
  NAND2_X1 U11979 ( .A1(n13817), .A2(n9655), .ZN(n9516) );
  NAND2_X1 U11980 ( .A1(n9517), .A2(n9516), .ZN(n9518) );
  NAND2_X1 U11981 ( .A1(n9519), .A2(n9518), .ZN(n9525) );
  INV_X1 U11982 ( .A(n9520), .ZN(n9523) );
  INV_X1 U11983 ( .A(n9521), .ZN(n9522) );
  NAND2_X1 U11984 ( .A1(n9523), .A2(n9522), .ZN(n9524) );
  NAND2_X1 U11985 ( .A1(n9525), .A2(n9524), .ZN(n9530) );
  NAND2_X1 U11986 ( .A1(n13903), .A2(n9632), .ZN(n9527) );
  NAND2_X1 U11987 ( .A1(n13797), .A2(n9655), .ZN(n9526) );
  NAND2_X1 U11988 ( .A1(n9527), .A2(n9526), .ZN(n9529) );
  AOI22_X1 U11989 ( .A1(n13903), .A2(n9578), .B1(n13797), .B2(n9632), .ZN(
        n9528) );
  NAND2_X1 U11990 ( .A1(n13898), .A2(n9578), .ZN(n9532) );
  NAND2_X1 U11991 ( .A1(n13515), .A2(n9632), .ZN(n9531) );
  NAND2_X1 U11992 ( .A1(n9532), .A2(n9531), .ZN(n9537) );
  NAND2_X1 U11993 ( .A1(n13898), .A2(n9632), .ZN(n9534) );
  NAND2_X1 U11994 ( .A1(n13515), .A2(n9655), .ZN(n9533) );
  NAND2_X1 U11995 ( .A1(n9534), .A2(n9533), .ZN(n9535) );
  NAND2_X1 U11996 ( .A1(n9536), .A2(n9535), .ZN(n9539) );
  NAND2_X1 U11997 ( .A1(n9539), .A2(n6622), .ZN(n9543) );
  NAND2_X1 U11998 ( .A1(n13893), .A2(n9632), .ZN(n9541) );
  NAND2_X1 U11999 ( .A1(n13741), .A2(n9655), .ZN(n9540) );
  AOI22_X1 U12000 ( .A1(n13893), .A2(n9578), .B1(n13741), .B2(n9632), .ZN(
        n9542) );
  NAND2_X1 U12001 ( .A1(n13887), .A2(n9655), .ZN(n9545) );
  NAND2_X1 U12002 ( .A1(n13514), .A2(n9632), .ZN(n9544) );
  NAND2_X1 U12003 ( .A1(n9545), .A2(n9544), .ZN(n9546) );
  INV_X1 U12004 ( .A(n13514), .ZN(n13417) );
  NAND2_X1 U12005 ( .A1(n13887), .A2(n9632), .ZN(n9547) );
  OAI21_X1 U12006 ( .B1(n13417), .B2(n9632), .A(n9547), .ZN(n9548) );
  NAND2_X1 U12007 ( .A1(n9549), .A2(n9548), .ZN(n9550) );
  NAND2_X1 U12008 ( .A1(n9551), .A2(n9550), .ZN(n9556) );
  NAND2_X1 U12009 ( .A1(n13879), .A2(n9632), .ZN(n9553) );
  NAND2_X1 U12010 ( .A1(n13742), .A2(n9655), .ZN(n9552) );
  NAND2_X1 U12011 ( .A1(n9553), .A2(n9552), .ZN(n9555) );
  AOI22_X1 U12012 ( .A1(n13879), .A2(n9655), .B1(n13742), .B2(n9632), .ZN(
        n9554) );
  NAND2_X1 U12013 ( .A1(n13875), .A2(n9655), .ZN(n9558) );
  NAND2_X1 U12014 ( .A1(n13684), .A2(n9632), .ZN(n9557) );
  NAND2_X1 U12015 ( .A1(n9558), .A2(n9557), .ZN(n9560) );
  AOI22_X1 U12016 ( .A1(n13875), .A2(n9632), .B1(n9578), .B2(n13684), .ZN(
        n9559) );
  AOI21_X1 U12017 ( .B1(n9561), .B2(n9560), .A(n9559), .ZN(n9563) );
  NAND2_X1 U12018 ( .A1(n13870), .A2(n9632), .ZN(n9565) );
  NAND2_X1 U12019 ( .A1(n13669), .A2(n9655), .ZN(n9564) );
  AOI22_X1 U12020 ( .A1(n13870), .A2(n9566), .B1(n13669), .B2(n9632), .ZN(
        n9567) );
  OAI22_X1 U12021 ( .A1(n13677), .A2(n9632), .B1(n13426), .B2(n9653), .ZN(
        n9569) );
  AOI22_X1 U12022 ( .A1(n13865), .A2(n9632), .B1(n9578), .B2(n13685), .ZN(
        n9568) );
  AOI22_X1 U12023 ( .A1(n13860), .A2(n9632), .B1(n9655), .B2(n13668), .ZN(
        n9571) );
  AOI22_X1 U12024 ( .A1(n13860), .A2(n9655), .B1(n13668), .B2(n9632), .ZN(
        n9572) );
  OAI22_X1 U12025 ( .A1(n13644), .A2(n9632), .B1(n13424), .B2(n9653), .ZN(
        n9576) );
  AOI22_X1 U12026 ( .A1(n13855), .A2(n9632), .B1(n9578), .B2(n13513), .ZN(
        n9574) );
  INV_X1 U12027 ( .A(n9574), .ZN(n9575) );
  AOI22_X1 U12028 ( .A1(n13849), .A2(n9632), .B1(n9578), .B2(n13637), .ZN(
        n9580) );
  INV_X1 U12029 ( .A(n9580), .ZN(n9577) );
  AOI22_X1 U12030 ( .A1(n13849), .A2(n9578), .B1(n13637), .B2(n9632), .ZN(
        n9579) );
  NOR2_X1 U12031 ( .A1(n9581), .A2(n9577), .ZN(n9646) );
  INV_X1 U12032 ( .A(n9583), .ZN(n9582) );
  OAI21_X1 U12033 ( .B1(n12503), .B2(n9582), .A(n9585), .ZN(n9588) );
  NOR2_X1 U12034 ( .A1(n9583), .A2(SI_27_), .ZN(n9586) );
  AOI21_X1 U12035 ( .B1(n9586), .B2(n9585), .A(n9584), .ZN(n9587) );
  MUX2_X1 U12036 ( .A(n14628), .B(n13950), .S(n10486), .Z(n9590) );
  XNOR2_X1 U12037 ( .A(n9590), .B(SI_29_), .ZN(n9622) );
  INV_X1 U12038 ( .A(n9590), .ZN(n9591) );
  NOR2_X1 U12039 ( .A1(n9591), .A2(SI_29_), .ZN(n9592) );
  MUX2_X1 U12040 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6546), .Z(n9593) );
  NAND2_X1 U12041 ( .A1(n9593), .A2(SI_30_), .ZN(n9595) );
  OAI21_X1 U12042 ( .B1(SI_30_), .B2(n9593), .A(n9595), .ZN(n9607) );
  INV_X1 U12043 ( .A(n9607), .ZN(n9594) );
  NAND2_X1 U12044 ( .A1(n9609), .A2(n9595), .ZN(n9598) );
  MUX2_X1 U12045 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10485), .Z(n9596) );
  XNOR2_X1 U12046 ( .A(n9596), .B(SI_31_), .ZN(n9597) );
  NAND2_X1 U12047 ( .A1(n13942), .A2(n8148), .ZN(n9600) );
  NAND2_X1 U12048 ( .A1(n9624), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n9599) );
  INV_X1 U12049 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9604) );
  NAND2_X1 U12050 ( .A1(n9612), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9603) );
  NAND2_X1 U12051 ( .A1(n9601), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9602) );
  OAI211_X1 U12052 ( .C1(n8136), .C2(n9604), .A(n9603), .B(n9602), .ZN(n13509)
         );
  INV_X1 U12053 ( .A(n13509), .ZN(n13596) );
  NAND2_X1 U12054 ( .A1(n13597), .A2(n13596), .ZN(n9656) );
  NAND2_X1 U12055 ( .A1(n9656), .A2(n9605), .ZN(n9695) );
  INV_X1 U12056 ( .A(n9606), .ZN(n9608) );
  NAND2_X1 U12057 ( .A1(n9624), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n9611) );
  INV_X1 U12058 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n15503) );
  NAND2_X1 U12059 ( .A1(n9612), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9615) );
  NAND2_X1 U12060 ( .A1(n9613), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9614) );
  OAI211_X1 U12061 ( .C1(n8139), .C2(n15503), .A(n9615), .B(n9614), .ZN(n13510) );
  AND2_X1 U12062 ( .A1(n13510), .A2(n9578), .ZN(n9616) );
  AOI21_X1 U12063 ( .B1(n13593), .B2(n9632), .A(n9616), .ZN(n9641) );
  NAND2_X1 U12064 ( .A1(n13593), .A2(n9655), .ZN(n9621) );
  OAI211_X1 U12065 ( .C1(n9617), .C2(n9789), .A(n8080), .B(n9664), .ZN(n9618)
         );
  AOI21_X1 U12066 ( .B1(n13509), .B2(n9632), .A(n9618), .ZN(n9619) );
  INV_X1 U12067 ( .A(n13510), .ZN(n9734) );
  OR2_X1 U12068 ( .A1(n9619), .A2(n9734), .ZN(n9620) );
  NAND2_X1 U12069 ( .A1(n9621), .A2(n9620), .ZN(n9640) );
  NAND2_X1 U12070 ( .A1(n13948), .A2(n8148), .ZN(n9626) );
  NAND2_X1 U12071 ( .A1(n9624), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n9625) );
  AND2_X1 U12072 ( .A1(n13511), .A2(n9655), .ZN(n9627) );
  AOI21_X1 U12073 ( .B1(n12603), .B2(n9632), .A(n9627), .ZN(n9636) );
  NAND2_X1 U12074 ( .A1(n12603), .A2(n9655), .ZN(n9629) );
  NAND2_X1 U12075 ( .A1(n13511), .A2(n9632), .ZN(n9628) );
  NAND2_X1 U12076 ( .A1(n9629), .A2(n9628), .ZN(n9635) );
  AOI22_X1 U12077 ( .A1(n9641), .A2(n9640), .B1(n9636), .B2(n9635), .ZN(n9630)
         );
  INV_X1 U12078 ( .A(n9695), .ZN(n9639) );
  AND2_X1 U12079 ( .A1(n13512), .A2(n9632), .ZN(n9631) );
  AOI21_X1 U12080 ( .B1(n13843), .B2(n9578), .A(n9631), .ZN(n9648) );
  NAND2_X1 U12081 ( .A1(n13843), .A2(n9632), .ZN(n9634) );
  NAND2_X1 U12082 ( .A1(n13512), .A2(n9655), .ZN(n9633) );
  NAND2_X1 U12083 ( .A1(n9634), .A2(n9633), .ZN(n9647) );
  INV_X1 U12084 ( .A(n9635), .ZN(n9638) );
  INV_X1 U12085 ( .A(n9636), .ZN(n9637) );
  NAND3_X1 U12086 ( .A1(n9639), .A2(n7943), .A3(n7940), .ZN(n9645) );
  INV_X1 U12087 ( .A(n9640), .ZN(n9643) );
  INV_X1 U12088 ( .A(n9641), .ZN(n9642) );
  AND2_X1 U12089 ( .A1(n9643), .A2(n9642), .ZN(n9644) );
  INV_X1 U12090 ( .A(n9647), .ZN(n9652) );
  INV_X1 U12091 ( .A(n9648), .ZN(n9651) );
  INV_X1 U12092 ( .A(n9649), .ZN(n9650) );
  NAND2_X1 U12093 ( .A1(n13509), .A2(n9653), .ZN(n9654) );
  OAI22_X1 U12094 ( .A1(n9656), .A2(n9655), .B1(n13597), .B2(n9654), .ZN(n9657) );
  INV_X1 U12095 ( .A(n10416), .ZN(n10412) );
  NAND2_X1 U12096 ( .A1(n10412), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12403) );
  NAND2_X1 U12097 ( .A1(n6555), .A2(n8080), .ZN(n9659) );
  OAI211_X1 U12098 ( .C1(n9667), .C2(n11758), .A(n9664), .B(n9659), .ZN(n9660)
         );
  INV_X1 U12099 ( .A(n9660), .ZN(n9661) );
  MUX2_X1 U12100 ( .A(n9667), .B(n8080), .S(n9789), .Z(n9662) );
  NOR2_X1 U12101 ( .A1(n12403), .A2(n9663), .ZN(n9670) );
  INV_X1 U12102 ( .A(n13955), .ZN(n10435) );
  INV_X1 U12103 ( .A(n9664), .ZN(n9665) );
  NAND4_X1 U12104 ( .A1(n15210), .A2(n10435), .A3(n13814), .A4(n9665), .ZN(
        n9666) );
  OAI211_X1 U12105 ( .C1(n9667), .C2(n12403), .A(n9666), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9668) );
  INV_X1 U12106 ( .A(n9668), .ZN(n9669) );
  AOI21_X1 U12107 ( .B1(n9701), .B2(n9670), .A(n9669), .ZN(n9703) );
  INV_X1 U12108 ( .A(n13511), .ZN(n9671) );
  XNOR2_X1 U12109 ( .A(n13855), .B(n13513), .ZN(n13639) );
  INV_X1 U12110 ( .A(n13669), .ZN(n13398) );
  XNOR2_X1 U12111 ( .A(n13870), .B(n13398), .ZN(n13689) );
  XNOR2_X1 U12112 ( .A(n13875), .B(n13684), .ZN(n13700) );
  NAND2_X1 U12113 ( .A1(n13887), .A2(n13417), .ZN(n9723) );
  OR2_X1 U12114 ( .A1(n13887), .A2(n13417), .ZN(n9672) );
  NAND2_X1 U12115 ( .A1(n9723), .A2(n9672), .ZN(n9722) );
  OR2_X1 U12116 ( .A1(n13893), .A2(n13741), .ZN(n9771) );
  NAND2_X1 U12117 ( .A1(n13893), .A2(n13741), .ZN(n9770) );
  NAND2_X1 U12118 ( .A1(n9771), .A2(n9770), .ZN(n13752) );
  INV_X1 U12119 ( .A(n13796), .ZN(n12442) );
  XNOR2_X1 U12120 ( .A(n13912), .B(n12442), .ZN(n13830) );
  XNOR2_X1 U12121 ( .A(n13907), .B(n13817), .ZN(n13795) );
  INV_X1 U12122 ( .A(n13516), .ZN(n12121) );
  XNOR2_X1 U12123 ( .A(n12253), .B(n12121), .ZN(n12245) );
  XNOR2_X1 U12124 ( .A(n12214), .B(n15112), .ZN(n12123) );
  XNOR2_X1 U12125 ( .A(n15252), .B(n9716), .ZN(n12073) );
  XNOR2_X1 U12126 ( .A(n15245), .B(n13520), .ZN(n11843) );
  INV_X1 U12127 ( .A(n13521), .ZN(n11620) );
  NAND2_X1 U12128 ( .A1(n11815), .A2(n11620), .ZN(n9713) );
  OR2_X1 U12129 ( .A1(n11815), .A2(n11620), .ZN(n9673) );
  NAND2_X1 U12130 ( .A1(n13527), .A2(n8105), .ZN(n9674) );
  NAND2_X1 U12131 ( .A1(n9675), .A2(n9674), .ZN(n15217) );
  NOR2_X1 U12132 ( .A1(n15217), .A2(n8079), .ZN(n9678) );
  NAND2_X1 U12133 ( .A1(n11194), .A2(n13524), .ZN(n9677) );
  INV_X1 U12134 ( .A(n13523), .ZN(n9679) );
  NAND2_X1 U12135 ( .A1(n15227), .A2(n9679), .ZN(n9710) );
  OR2_X1 U12136 ( .A1(n15227), .A2(n9679), .ZN(n9680) );
  NAND2_X1 U12137 ( .A1(n9710), .A2(n9680), .ZN(n9743) );
  NOR2_X1 U12138 ( .A1(n9681), .A2(n9743), .ZN(n9682) );
  XNOR2_X1 U12139 ( .A(n11837), .B(n13522), .ZN(n11827) );
  NAND4_X1 U12140 ( .A1(n11843), .A2(n11294), .A3(n9682), .A4(n11827), .ZN(
        n9683) );
  NOR2_X1 U12141 ( .A1(n12073), .A2(n9683), .ZN(n9684) );
  XNOR2_X1 U12142 ( .A(n12102), .B(n13517), .ZN(n12091) );
  NAND4_X1 U12143 ( .A1(n12123), .A2(n9684), .A3(n7803), .A4(n12091), .ZN(
        n9685) );
  NOR2_X1 U12144 ( .A1(n12245), .A2(n9685), .ZN(n9686) );
  XNOR2_X1 U12145 ( .A(n14847), .B(n13815), .ZN(n12449) );
  XNOR2_X1 U12146 ( .A(n12420), .B(n15114), .ZN(n12237) );
  NAND4_X1 U12147 ( .A1(n13795), .A2(n9686), .A3(n12449), .A4(n12237), .ZN(
        n9687) );
  NOR2_X1 U12148 ( .A1(n13830), .A2(n9687), .ZN(n9688) );
  XNOR2_X1 U12149 ( .A(n13898), .B(n13515), .ZN(n13760) );
  XNOR2_X1 U12150 ( .A(n13903), .B(n13797), .ZN(n13777) );
  NAND4_X1 U12151 ( .A1(n13752), .A2(n9688), .A3(n13760), .A4(n13777), .ZN(
        n9689) );
  NOR2_X1 U12152 ( .A1(n9722), .A2(n9689), .ZN(n9690) );
  XNOR2_X1 U12153 ( .A(n13879), .B(n13742), .ZN(n13726) );
  NAND3_X1 U12154 ( .A1(n13700), .A2(n9690), .A3(n13726), .ZN(n9691) );
  NOR2_X1 U12155 ( .A1(n13689), .A2(n9691), .ZN(n9693) );
  NAND2_X1 U12156 ( .A1(n13677), .A2(n13426), .ZN(n9692) );
  NAND2_X1 U12157 ( .A1(n13865), .A2(n13685), .ZN(n9779) );
  NAND2_X1 U12158 ( .A1(n9692), .A2(n9779), .ZN(n9778) );
  XNOR2_X1 U12159 ( .A(n13860), .B(n13668), .ZN(n13653) );
  NAND4_X1 U12160 ( .A1(n13639), .A2(n9693), .A3(n9778), .A4(n13653), .ZN(
        n9694) );
  NAND2_X1 U12161 ( .A1(n13843), .A2(n13512), .ZN(n9787) );
  OR2_X1 U12162 ( .A1(n13843), .A2(n13512), .ZN(n9696) );
  XOR2_X1 U12163 ( .A(n9698), .B(n9697), .Z(n9699) );
  NOR3_X1 U12164 ( .A1(n9699), .A2(n8080), .A3(n12403), .ZN(n9700) );
  OAI21_X1 U12165 ( .B1(n9701), .B2(n9789), .A(n9700), .ZN(n9702) );
  NAND3_X1 U12166 ( .A1(n9704), .A2(n9703), .A3(n9702), .ZN(P2_U3328) );
  INV_X1 U12167 ( .A(n13860), .ZN(n9729) );
  INV_X1 U12168 ( .A(n13893), .ZN(n13750) );
  INV_X1 U12169 ( .A(n13741), .ZN(n13468) );
  INV_X1 U12170 ( .A(n13898), .ZN(n13767) );
  INV_X1 U12171 ( .A(n13515), .ZN(n9720) );
  INV_X1 U12172 ( .A(n13903), .ZN(n13783) );
  INV_X1 U12173 ( .A(n13797), .ZN(n13442) );
  INV_X1 U12174 ( .A(n15114), .ZN(n12443) );
  INV_X1 U12175 ( .A(n12253), .ZN(n15118) );
  INV_X1 U12176 ( .A(n12214), .ZN(n12132) );
  NAND2_X1 U12177 ( .A1(n9705), .A2(n9426), .ZN(n9707) );
  INV_X1 U12178 ( .A(n6553), .ZN(n15222) );
  NAND2_X1 U12179 ( .A1(n9707), .A2(n9706), .ZN(n11785) );
  NAND2_X1 U12180 ( .A1(n11784), .A2(n9708), .ZN(n11190) );
  INV_X1 U12181 ( .A(n9743), .ZN(n11763) );
  NAND2_X1 U12182 ( .A1(n11837), .A2(n9711), .ZN(n9712) );
  OR2_X1 U12183 ( .A1(n15245), .A2(n11451), .ZN(n9714) );
  NAND2_X1 U12184 ( .A1(n15245), .A2(n11451), .ZN(n9715) );
  INV_X1 U12185 ( .A(n12073), .ZN(n12078) );
  INV_X1 U12186 ( .A(n13517), .ZN(n12122) );
  NAND2_X1 U12187 ( .A1(n12102), .A2(n12122), .ZN(n9717) );
  INV_X1 U12188 ( .A(n12102), .ZN(n15264) );
  INV_X1 U12189 ( .A(n12420), .ZN(n12236) );
  NOR2_X1 U12190 ( .A1(n13912), .A2(n12442), .ZN(n9718) );
  INV_X1 U12191 ( .A(n13817), .ZN(n13502) );
  INV_X1 U12192 ( .A(n13907), .ZN(n13806) );
  INV_X1 U12193 ( .A(n13879), .ZN(n9724) );
  NAND2_X1 U12194 ( .A1(n9724), .A2(n13742), .ZN(n9725) );
  INV_X1 U12195 ( .A(n13742), .ZN(n13469) );
  NAND2_X1 U12196 ( .A1(n13683), .A2(n9727), .ZN(n9728) );
  INV_X1 U12197 ( .A(n13637), .ZN(n9730) );
  OAI21_X1 U12198 ( .B1(n9735), .B2(n13843), .A(n13608), .ZN(n9731) );
  NAND2_X1 U12199 ( .A1(n8080), .A2(n9789), .ZN(n9732) );
  INV_X1 U12200 ( .A(n13814), .ZN(n13425) );
  INV_X1 U12201 ( .A(P2_B_REG_SCAN_IN), .ZN(n9733) );
  OAI21_X1 U12202 ( .B1(n13955), .B2(n9733), .A(n13816), .ZN(n13595) );
  OAI22_X1 U12203 ( .A1(n9735), .A2(n13425), .B1(n9734), .B2(n13595), .ZN(
        n9736) );
  AND2_X1 U12204 ( .A1(n13527), .A2(n9791), .ZN(n12065) );
  NAND2_X1 U12205 ( .A1(n9738), .A2(n9737), .ZN(n11777) );
  NAND2_X1 U12206 ( .A1(n11777), .A2(n9739), .ZN(n9741) );
  OR2_X1 U12207 ( .A1(n13525), .A2(n13922), .ZN(n9740) );
  INV_X1 U12208 ( .A(n11191), .ZN(n11187) );
  OR2_X1 U12209 ( .A1(n13524), .A2(n12043), .ZN(n9742) );
  OR2_X1 U12210 ( .A1(n15227), .A2(n13523), .ZN(n9744) );
  INV_X1 U12211 ( .A(n11827), .ZN(n9745) );
  NAND2_X1 U12212 ( .A1(n11823), .A2(n9745), .ZN(n9747) );
  OR2_X1 U12213 ( .A1(n11837), .A2(n13522), .ZN(n9746) );
  INV_X1 U12214 ( .A(n11294), .ZN(n9748) );
  OR2_X1 U12215 ( .A1(n11815), .A2(n13521), .ZN(n9749) );
  INV_X1 U12216 ( .A(n11843), .ZN(n9750) );
  OR2_X1 U12217 ( .A1(n15245), .A2(n13520), .ZN(n9751) );
  NAND2_X1 U12218 ( .A1(n11611), .A2(n13519), .ZN(n9753) );
  NAND2_X1 U12219 ( .A1(n15252), .A2(n13518), .ZN(n9754) );
  OR2_X1 U12220 ( .A1(n12102), .A2(n13517), .ZN(n9755) );
  AND2_X1 U12221 ( .A1(n12214), .A2(n15112), .ZN(n9756) );
  NOR2_X1 U12222 ( .A1(n12253), .A2(n13516), .ZN(n9757) );
  NAND2_X1 U12223 ( .A1(n12253), .A2(n13516), .ZN(n9758) );
  AND2_X1 U12224 ( .A1(n12420), .A2(n15114), .ZN(n9760) );
  OR2_X1 U12225 ( .A1(n12420), .A2(n15114), .ZN(n9761) );
  NOR2_X1 U12226 ( .A1(n14847), .A2(n13815), .ZN(n9762) );
  NAND2_X1 U12227 ( .A1(n14847), .A2(n13815), .ZN(n9763) );
  OR2_X1 U12228 ( .A1(n13912), .A2(n13796), .ZN(n9764) );
  NAND2_X1 U12229 ( .A1(n13907), .A2(n13817), .ZN(n9766) );
  AND2_X1 U12230 ( .A1(n13903), .A2(n13797), .ZN(n9767) );
  INV_X1 U12231 ( .A(n13760), .ZN(n13762) );
  OR2_X1 U12232 ( .A1(n13898), .A2(n13515), .ZN(n9768) );
  NAND2_X1 U12233 ( .A1(n13747), .A2(n9770), .ZN(n9772) );
  NAND2_X1 U12234 ( .A1(n13887), .A2(n13514), .ZN(n9773) );
  NAND2_X1 U12235 ( .A1(n13731), .A2(n9773), .ZN(n9775) );
  OR2_X1 U12236 ( .A1(n13887), .A2(n13514), .ZN(n9774) );
  NAND2_X1 U12237 ( .A1(n13879), .A2(n13742), .ZN(n9776) );
  NAND2_X1 U12238 ( .A1(n13870), .A2(n13669), .ZN(n9777) );
  OR2_X1 U12239 ( .A1(n13860), .A2(n13668), .ZN(n9781) );
  AND2_X1 U12240 ( .A1(n13860), .A2(n13668), .ZN(n9780) );
  OR2_X1 U12241 ( .A1(n13644), .A2(n13424), .ZN(n9782) );
  NAND2_X1 U12242 ( .A1(n13644), .A2(n13424), .ZN(n9783) );
  NAND2_X1 U12243 ( .A1(n13849), .A2(n13637), .ZN(n9785) );
  AND2_X1 U12244 ( .A1(n12066), .A2(n11781), .ZN(n11778) );
  INV_X1 U12245 ( .A(n15227), .ZN(n11771) );
  INV_X1 U12246 ( .A(n15245), .ZN(n11852) );
  INV_X1 U12247 ( .A(n11611), .ZN(n11807) );
  OR2_X2 U12248 ( .A1(n12249), .A2(n12420), .ZN(n12445) );
  OR2_X2 U12249 ( .A1(n13898), .A2(n13780), .ZN(n13765) );
  NAND2_X1 U12250 ( .A1(n13677), .A2(n13693), .ZN(n13671) );
  NAND2_X1 U12251 ( .A1(n13644), .A2(n13662), .ZN(n13646) );
  AND2_X1 U12252 ( .A1(n15210), .A2(n9797), .ZN(n15211) );
  AND3_X1 U12253 ( .A1(n11754), .A2(n9798), .A3(n11753), .ZN(n9799) );
  NOR2_X2 U12254 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9888) );
  AND2_X2 U12255 ( .A1(n9888), .A2(n9802), .ZN(n9920) );
  NOR2_X1 U12256 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n9806) );
  NOR2_X1 U12258 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), 
        .ZN(n9807) );
  NOR2_X1 U12259 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n9812) );
  NOR2_X1 U12260 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n9815) );
  NAND2_X2 U12261 ( .A1(n10563), .A2(n8013), .ZN(n10265) );
  INV_X2 U12262 ( .A(n10265), .ZN(n9867) );
  NAND2_X1 U12263 ( .A1(n12536), .A2(n10237), .ZN(n9818) );
  INV_X2 U12264 ( .A(n9863), .ZN(n10298) );
  NAND2_X1 U12265 ( .A1(n10298), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9817) );
  NAND2_X1 U12266 ( .A1(n9822), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9823) );
  NAND2_X1 U12267 ( .A1(n6549), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9835) );
  AND2_X4 U12268 ( .A1(n14623), .A2(n9825), .ZN(n10260) );
  INV_X1 U12269 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9824) );
  OR2_X1 U12270 ( .A1(n9927), .A2(n9824), .ZN(n9834) );
  NAND2_X1 U12271 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9929) );
  NOR2_X1 U12272 ( .A1(n9929), .A2(n9928), .ZN(n9946) );
  NAND2_X1 U12273 ( .A1(n9946), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9965) );
  NAND2_X1 U12274 ( .A1(n10008), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10019) );
  NAND2_X1 U12275 ( .A1(n10058), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10076) );
  INV_X1 U12276 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n10075) );
  INV_X1 U12277 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n10087) );
  NAND2_X1 U12278 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n9827) );
  NAND2_X1 U12279 ( .A1(n10176), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n10177) );
  NAND2_X1 U12280 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n10223), .ZN(n10222) );
  INV_X1 U12281 ( .A(n10222), .ZN(n9828) );
  NAND2_X1 U12282 ( .A1(n9828), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n10241) );
  INV_X1 U12283 ( .A(n10241), .ZN(n9829) );
  NAND2_X1 U12284 ( .A1(n9829), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n10276) );
  INV_X1 U12285 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9830) );
  XNOR2_X1 U12286 ( .A(n10276), .B(n9830), .ZN(n12784) );
  OR2_X1 U12287 ( .A1(n10278), .A2(n12784), .ZN(n9833) );
  AND2_X4 U12288 ( .A1(n14623), .A2(n14626), .ZN(n9893) );
  INV_X1 U12289 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9831) );
  OR2_X1 U12290 ( .A1(n10257), .A2(n9831), .ZN(n9832) );
  INV_X1 U12291 ( .A(n10700), .ZN(n12021) );
  NAND2_X1 U12292 ( .A1(n9845), .A2(n12021), .ZN(n10270) );
  NAND2_X1 U12293 ( .A1(n10366), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9844) );
  OR2_X1 U12294 ( .A1(n9845), .A2(n11897), .ZN(n9846) );
  NAND2_X2 U12295 ( .A1(n9846), .A2(n10270), .ZN(n10283) );
  MUX2_X1 U12296 ( .A(n7158), .B(n14274), .S(n10283), .Z(n10255) );
  INV_X1 U12297 ( .A(n10255), .ZN(n10288) );
  NAND2_X1 U12298 ( .A1(n9893), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9853) );
  INV_X1 U12299 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9847) );
  OR2_X1 U12300 ( .A1(n9861), .A2(n9847), .ZN(n9852) );
  INV_X1 U12301 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14075) );
  NAND2_X1 U12302 ( .A1(n10222), .A2(n14075), .ZN(n9848) );
  NAND2_X1 U12303 ( .A1(n10241), .A2(n9848), .ZN(n14294) );
  OR2_X1 U12304 ( .A1(n10278), .A2(n14294), .ZN(n9851) );
  INV_X1 U12305 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9849) );
  OR2_X1 U12306 ( .A1(n9927), .A2(n9849), .ZN(n9850) );
  NAND2_X1 U12307 ( .A1(n13958), .A2(n9867), .ZN(n9855) );
  NAND2_X1 U12308 ( .A1(n10298), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9854) );
  MUX2_X1 U12309 ( .A(n14275), .B(n14297), .S(n10216), .Z(n10234) );
  NAND2_X1 U12310 ( .A1(n6549), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9860) );
  NAND2_X1 U12311 ( .A1(n10260), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9859) );
  NAND2_X1 U12312 ( .A1(n9893), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9858) );
  INV_X1 U12313 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9856) );
  NAND2_X1 U12314 ( .A1(n9893), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9862) );
  INV_X1 U12315 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n11437) );
  INV_X1 U12316 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10631) );
  INV_X1 U12317 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14127) );
  INV_X4 U12318 ( .A(n10563), .ZN(n10136) );
  OR2_X1 U12319 ( .A1(n9888), .A2(n14617), .ZN(n9864) );
  XNOR2_X1 U12320 ( .A(n9864), .B(P1_IR_REG_2__SCAN_IN), .ZN(n14129) );
  NAND2_X1 U12321 ( .A1(n10479), .A2(n9867), .ZN(n9865) );
  NAND2_X1 U12322 ( .A1(n10283), .A2(n14109), .ZN(n9866) );
  NAND2_X1 U12323 ( .A1(n9866), .A2(n7324), .ZN(n9871) );
  NAND2_X1 U12324 ( .A1(n10491), .A2(n9867), .ZN(n9870) );
  INV_X1 U12325 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n14617) );
  OR2_X1 U12326 ( .A1(n9920), .A2(n14617), .ZN(n9868) );
  XNOR2_X1 U12327 ( .A(n9868), .B(P1_IR_REG_3__SCAN_IN), .ZN(n14148) );
  AOI21_X1 U12328 ( .B1(n9872), .B2(n9871), .A(n14933), .ZN(n9880) );
  OAI21_X1 U12329 ( .B1(n10283), .B2(n14109), .A(n11440), .ZN(n9875) );
  NAND3_X1 U12330 ( .A1(n10283), .A2(n14108), .A3(n14109), .ZN(n9873) );
  NAND2_X1 U12331 ( .A1(n9873), .A2(n7324), .ZN(n9874) );
  AOI21_X1 U12332 ( .B1(n9875), .B2(n9874), .A(n11478), .ZN(n9879) );
  NAND3_X1 U12333 ( .A1(n11478), .A2(n14108), .A3(n10283), .ZN(n9877) );
  NAND3_X1 U12334 ( .A1(n11479), .A2(n10216), .A3(n14933), .ZN(n9876) );
  AND2_X1 U12335 ( .A1(n9877), .A2(n9876), .ZN(n9878) );
  INV_X1 U12336 ( .A(n9881), .ZN(n9914) );
  NAND2_X1 U12337 ( .A1(n6549), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9885) );
  NAND2_X1 U12338 ( .A1(n10260), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9884) );
  NAND2_X1 U12339 ( .A1(n9886), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9892) );
  NAND2_X1 U12340 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9887) );
  MUX2_X1 U12341 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9887), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n9890) );
  INV_X1 U12342 ( .A(n9888), .ZN(n9889) );
  NAND2_X1 U12343 ( .A1(n9890), .A2(n9889), .ZN(n10650) );
  INV_X1 U12344 ( .A(n10650), .ZN(n14113) );
  NAND2_X1 U12345 ( .A1(n10136), .A2(n14113), .ZN(n9891) );
  MUX2_X1 U12346 ( .A(n14494), .B(n14110), .S(n10283), .Z(n9908) );
  NAND2_X1 U12347 ( .A1(n10179), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9897) );
  NAND2_X1 U12348 ( .A1(n6549), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9896) );
  NAND2_X1 U12349 ( .A1(n10260), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9895) );
  INV_X1 U12350 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14123) );
  INV_X1 U12351 ( .A(SI_0_), .ZN(n9899) );
  OAI21_X1 U12352 ( .B1(n10486), .B2(n9899), .A(n9898), .ZN(n9900) );
  NAND2_X1 U12353 ( .A1(n9901), .A2(n9900), .ZN(n14642) );
  MUX2_X1 U12354 ( .A(n14123), .B(n14642), .S(n10563), .Z(n11463) );
  AND2_X1 U12355 ( .A1(n11168), .A2(n11463), .ZN(n10314) );
  NAND2_X1 U12356 ( .A1(n9906), .A2(n9905), .ZN(n9907) );
  OAI21_X1 U12357 ( .B1(n10316), .B2(n9908), .A(n9907), .ZN(n9910) );
  NAND2_X1 U12358 ( .A1(n14110), .A2(n14494), .ZN(n10317) );
  NAND2_X1 U12359 ( .A1(n9908), .A2(n10317), .ZN(n9909) );
  NAND2_X1 U12360 ( .A1(n9910), .A2(n9909), .ZN(n9912) );
  NAND2_X1 U12361 ( .A1(n11338), .A2(n7324), .ZN(n11308) );
  NAND2_X1 U12362 ( .A1(n14109), .A2(n11440), .ZN(n9911) );
  NAND2_X1 U12363 ( .A1(n9912), .A2(n10318), .ZN(n9913) );
  NAND2_X1 U12364 ( .A1(n9893), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9918) );
  NAND2_X1 U12365 ( .A1(n6549), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9917) );
  NAND2_X1 U12366 ( .A1(n10260), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9916) );
  OAI21_X1 U12367 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n9929), .ZN(n11537) );
  NAND4_X1 U12368 ( .A1(n9918), .A2(n9917), .A3(n9916), .A4(n9915), .ZN(n14107) );
  NAND2_X1 U12369 ( .A1(n10496), .A2(n10237), .ZN(n9923) );
  INV_X1 U12370 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9919) );
  NAND2_X1 U12371 ( .A1(n9920), .A2(n9919), .ZN(n9935) );
  NAND2_X1 U12372 ( .A1(n9935), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9921) );
  XNOR2_X1 U12373 ( .A(n9921), .B(P1_IR_REG_4__SCAN_IN), .ZN(n14161) );
  AOI22_X1 U12374 ( .A1(n10298), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n10136), 
        .B2(n14161), .ZN(n9922) );
  MUX2_X1 U12375 ( .A(n14107), .B(n11587), .S(n10216), .Z(n9924) );
  INV_X1 U12376 ( .A(n9924), .ZN(n9925) );
  NAND2_X1 U12377 ( .A1(n9893), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9934) );
  INV_X1 U12378 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10657) );
  OR2_X1 U12379 ( .A1(n9861), .A2(n10657), .ZN(n9933) );
  INV_X1 U12380 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10629) );
  OR2_X1 U12381 ( .A1(n9927), .A2(n10629), .ZN(n9932) );
  AND2_X1 U12382 ( .A1(n9929), .A2(n9928), .ZN(n9930) );
  OR2_X1 U12383 ( .A1(n9930), .A2(n9946), .ZN(n15004) );
  OR2_X1 U12384 ( .A1(n10278), .A2(n15004), .ZN(n9931) );
  NAND2_X1 U12385 ( .A1(n10482), .A2(n10237), .ZN(n9938) );
  NAND2_X1 U12386 ( .A1(n9952), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9936) );
  XNOR2_X1 U12387 ( .A(n9936), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10798) );
  AOI22_X1 U12388 ( .A1(n10298), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n10136), 
        .B2(n10798), .ZN(n9937) );
  MUX2_X1 U12389 ( .A(n11595), .B(n15008), .S(n10283), .Z(n9942) );
  INV_X1 U12390 ( .A(n9942), .ZN(n9939) );
  INV_X1 U12391 ( .A(n11595), .ZN(n14106) );
  INV_X1 U12392 ( .A(n15008), .ZN(n15016) );
  MUX2_X1 U12393 ( .A(n14106), .B(n15016), .S(n10216), .Z(n9940) );
  NAND2_X1 U12394 ( .A1(n9941), .A2(n9940), .ZN(n9945) );
  NAND2_X1 U12395 ( .A1(n9943), .A2(n9942), .ZN(n9944) );
  NAND2_X1 U12396 ( .A1(n6549), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9951) );
  NAND2_X1 U12397 ( .A1(n10260), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9950) );
  NAND2_X1 U12398 ( .A1(n9893), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9949) );
  OR2_X1 U12399 ( .A1(n9946), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9947) );
  NAND2_X1 U12400 ( .A1(n9965), .A2(n9947), .ZN(n11660) );
  OR2_X1 U12401 ( .A1(n10278), .A2(n11660), .ZN(n9948) );
  NAND4_X1 U12402 ( .A1(n9951), .A2(n9950), .A3(n9949), .A4(n9948), .ZN(n14105) );
  NAND2_X1 U12403 ( .A1(n10498), .A2(n10237), .ZN(n9959) );
  NOR2_X1 U12404 ( .A1(n9955), .A2(n14617), .ZN(n9953) );
  MUX2_X1 U12405 ( .A(n14617), .B(n9953), .S(P1_IR_REG_6__SCAN_IN), .Z(n9957)
         );
  INV_X1 U12406 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9954) );
  NAND2_X1 U12407 ( .A1(n9955), .A2(n9954), .ZN(n10028) );
  INV_X1 U12408 ( .A(n10028), .ZN(n9956) );
  NOR2_X1 U12409 ( .A1(n9957), .A2(n9956), .ZN(n14179) );
  AOI22_X1 U12410 ( .A1(n10298), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n10136), 
        .B2(n14179), .ZN(n9958) );
  NAND2_X1 U12411 ( .A1(n9959), .A2(n9958), .ZN(n11719) );
  MUX2_X1 U12412 ( .A(n14105), .B(n11719), .S(n10216), .Z(n9960) );
  MUX2_X1 U12413 ( .A(n14105), .B(n11719), .S(n10301), .Z(n9961) );
  NAND2_X1 U12414 ( .A1(n9962), .A2(n9961), .ZN(n9963) );
  NAND2_X1 U12415 ( .A1(n9893), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9970) );
  NAND2_X1 U12416 ( .A1(n6549), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9969) );
  NAND2_X1 U12417 ( .A1(n10260), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9968) );
  NAND2_X1 U12418 ( .A1(n9965), .A2(n11678), .ZN(n9966) );
  NAND2_X1 U12419 ( .A1(n9978), .A2(n9966), .ZN(n14988) );
  OR2_X1 U12420 ( .A1(n10278), .A2(n14988), .ZN(n9967) );
  NAND4_X1 U12421 ( .A1(n9970), .A2(n9969), .A3(n9968), .A4(n9967), .ZN(n14104) );
  NAND2_X1 U12422 ( .A1(n10508), .A2(n10237), .ZN(n9973) );
  NAND2_X1 U12423 ( .A1(n10028), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9971) );
  XNOR2_X1 U12424 ( .A(n9971), .B(P1_IR_REG_7__SCAN_IN), .ZN(n14194) );
  AOI22_X1 U12425 ( .A1(n10298), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n10136), 
        .B2(n14194), .ZN(n9972) );
  MUX2_X1 U12426 ( .A(n14104), .B(n11734), .S(n10301), .Z(n9975) );
  MUX2_X1 U12427 ( .A(n14104), .B(n11734), .S(n10216), .Z(n9974) );
  NAND2_X1 U12428 ( .A1(n6549), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9983) );
  NAND2_X1 U12429 ( .A1(n9893), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9982) );
  NAND2_X1 U12430 ( .A1(n10260), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9981) );
  NAND2_X1 U12431 ( .A1(n9978), .A2(n9977), .ZN(n9979) );
  NAND2_X1 U12432 ( .A1(n9990), .A2(n9979), .ZN(n14950) );
  OR2_X1 U12433 ( .A1(n10278), .A2(n14950), .ZN(n9980) );
  NAND4_X1 U12434 ( .A1(n9983), .A2(n9982), .A3(n9981), .A4(n9980), .ZN(n14103) );
  NAND2_X1 U12435 ( .A1(n10512), .A2(n10237), .ZN(n9986) );
  OR2_X1 U12436 ( .A1(n10028), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9984) );
  NAND2_X1 U12437 ( .A1(n9984), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9999) );
  XNOR2_X1 U12438 ( .A(n9999), .B(P1_IR_REG_8__SCAN_IN), .ZN(n14205) );
  AOI22_X1 U12439 ( .A1(n10298), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n14205), 
        .B2(n10136), .ZN(n9985) );
  NAND2_X1 U12440 ( .A1(n9986), .A2(n9985), .ZN(n14943) );
  MUX2_X1 U12441 ( .A(n14103), .B(n14943), .S(n10216), .Z(n9988) );
  MUX2_X1 U12442 ( .A(n14103), .B(n14943), .S(n10301), .Z(n9987) );
  NAND2_X1 U12443 ( .A1(n9893), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9997) );
  NAND2_X1 U12444 ( .A1(n6549), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9996) );
  INV_X1 U12445 ( .A(n10008), .ZN(n9992) );
  NAND2_X1 U12446 ( .A1(n9990), .A2(n10794), .ZN(n9991) );
  NAND2_X1 U12447 ( .A1(n9992), .A2(n9991), .ZN(n14966) );
  OR2_X1 U12448 ( .A1(n10278), .A2(n14966), .ZN(n9995) );
  INV_X1 U12449 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9993) );
  OR2_X1 U12450 ( .A1(n9927), .A2(n9993), .ZN(n9994) );
  NAND4_X1 U12451 ( .A1(n9997), .A2(n9996), .A3(n9995), .A4(n9994), .ZN(n14102) );
  OR2_X1 U12452 ( .A1(n10518), .A2(n10265), .ZN(n10004) );
  INV_X1 U12453 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9998) );
  NAND2_X1 U12454 ( .A1(n9999), .A2(n9998), .ZN(n10000) );
  NAND2_X1 U12455 ( .A1(n10000), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10001) );
  NAND2_X1 U12456 ( .A1(n10001), .A2(n15595), .ZN(n10014) );
  OR2_X1 U12457 ( .A1(n10001), .A2(n15595), .ZN(n10002) );
  AOI22_X1 U12458 ( .A1(n10976), .A2(n10136), .B1(n10298), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n10003) );
  MUX2_X1 U12459 ( .A(n14102), .B(n14952), .S(n10301), .Z(n10007) );
  MUX2_X1 U12460 ( .A(n14102), .B(n14952), .S(n10216), .Z(n10005) );
  NAND2_X1 U12461 ( .A1(n6549), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10013) );
  NAND2_X1 U12462 ( .A1(n10260), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10012) );
  NAND2_X1 U12463 ( .A1(n9893), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n10011) );
  OR2_X1 U12464 ( .A1(n10008), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10009) );
  NAND2_X1 U12465 ( .A1(n10019), .A2(n10009), .ZN(n14882) );
  OR2_X1 U12466 ( .A1(n10278), .A2(n14882), .ZN(n10010) );
  NAND4_X1 U12467 ( .A1(n10013), .A2(n10012), .A3(n10011), .A4(n10010), .ZN(
        n14101) );
  NAND2_X1 U12468 ( .A1(n10014), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10015) );
  XNOR2_X1 U12469 ( .A(n10015), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11002) );
  AOI22_X1 U12470 ( .A1(n11002), .A2(n10136), .B1(P2_DATAO_REG_10__SCAN_IN), 
        .B2(n10298), .ZN(n10016) );
  MUX2_X1 U12471 ( .A(n14101), .B(n14870), .S(n10216), .Z(n10018) );
  MUX2_X1 U12472 ( .A(n14101), .B(n14870), .S(n10301), .Z(n10017) );
  NAND2_X1 U12473 ( .A1(n6549), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10024) );
  NAND2_X1 U12474 ( .A1(n10260), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10023) );
  NAND2_X1 U12475 ( .A1(n9893), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n10022) );
  NAND2_X1 U12476 ( .A1(n10019), .A2(n15586), .ZN(n10020) );
  NAND2_X1 U12477 ( .A1(n10038), .A2(n10020), .ZN(n14886) );
  OR2_X1 U12478 ( .A1(n10278), .A2(n14886), .ZN(n10021) );
  NAND4_X1 U12479 ( .A1(n10024), .A2(n10023), .A3(n10022), .A4(n10021), .ZN(
        n14100) );
  NAND2_X1 U12480 ( .A1(n10570), .A2(n10237), .ZN(n10031) );
  INV_X1 U12481 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n10025) );
  NAND3_X1 U12482 ( .A1(n10026), .A2(n15595), .A3(n10025), .ZN(n10027) );
  NAND2_X1 U12483 ( .A1(n10045), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10029) );
  XNOR2_X1 U12484 ( .A(n10029), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11024) );
  AOI22_X1 U12485 ( .A1(n10298), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n11024), 
        .B2(n10136), .ZN(n10030) );
  MUX2_X1 U12486 ( .A(n14100), .B(n14892), .S(n10301), .Z(n10034) );
  MUX2_X1 U12487 ( .A(n14100), .B(n14892), .S(n10216), .Z(n10032) );
  INV_X1 U12488 ( .A(n10034), .ZN(n10035) );
  INV_X1 U12489 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10036) );
  OR2_X1 U12490 ( .A1(n9861), .A2(n10036), .ZN(n10044) );
  NAND2_X1 U12491 ( .A1(n10260), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10043) );
  NAND2_X1 U12492 ( .A1(n9893), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10042) );
  INV_X1 U12493 ( .A(n10058), .ZN(n10040) );
  NAND2_X1 U12494 ( .A1(n10038), .A2(n10037), .ZN(n10039) );
  NAND2_X1 U12495 ( .A1(n10040), .A2(n10039), .ZN(n12481) );
  OR2_X1 U12496 ( .A1(n10278), .A2(n12481), .ZN(n10041) );
  NAND4_X1 U12497 ( .A1(n10044), .A2(n10043), .A3(n10042), .A4(n10041), .ZN(
        n14099) );
  NAND2_X1 U12498 ( .A1(n10615), .A2(n10237), .ZN(n10052) );
  NOR2_X1 U12499 ( .A1(n10045), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n10048) );
  OR2_X1 U12500 ( .A1(n10048), .A2(n14617), .ZN(n10046) );
  INV_X1 U12501 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10047) );
  MUX2_X1 U12502 ( .A(n10046), .B(P1_IR_REG_31__SCAN_IN), .S(n10047), .Z(
        n10049) );
  NAND2_X1 U12503 ( .A1(n10048), .A2(n10047), .ZN(n10071) );
  NOR2_X1 U12504 ( .A1(n9863), .A2(n15628), .ZN(n10050) );
  AOI21_X1 U12505 ( .B1(n11246), .B2(n10136), .A(n10050), .ZN(n10051) );
  MUX2_X1 U12506 ( .A(n14099), .B(n12476), .S(n10216), .Z(n10055) );
  MUX2_X1 U12507 ( .A(n14099), .B(n12476), .S(n10301), .Z(n10053) );
  NAND2_X1 U12508 ( .A1(n10054), .A2(n10053), .ZN(n10057) );
  OR2_X1 U12509 ( .A1(n10058), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10059) );
  AND2_X1 U12510 ( .A1(n10076), .A2(n10059), .ZN(n12172) );
  NAND2_X1 U12511 ( .A1(n12172), .A2(n10179), .ZN(n10063) );
  NAND2_X1 U12512 ( .A1(n9893), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n10062) );
  INV_X1 U12513 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n12173) );
  OR2_X1 U12514 ( .A1(n9861), .A2(n12173), .ZN(n10061) );
  INV_X1 U12515 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11257) );
  OR2_X1 U12516 ( .A1(n9927), .A2(n11257), .ZN(n10060) );
  NAND4_X1 U12517 ( .A1(n10063), .A2(n10062), .A3(n10061), .A4(n10060), .ZN(
        n14098) );
  NAND2_X1 U12518 ( .A1(n10627), .A2(n10237), .ZN(n10068) );
  NAND2_X1 U12519 ( .A1(n10071), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10064) );
  XNOR2_X1 U12520 ( .A(n10064), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11261) );
  NOR2_X1 U12521 ( .A1(n9863), .A2(n10065), .ZN(n10066) );
  AOI21_X1 U12522 ( .B1(n11261), .B2(n10136), .A(n10066), .ZN(n10067) );
  MUX2_X1 U12523 ( .A(n14098), .B(n12499), .S(n10301), .Z(n10070) );
  INV_X1 U12524 ( .A(n14098), .ZN(n12491) );
  INV_X1 U12525 ( .A(n12499), .ZN(n12492) );
  MUX2_X1 U12526 ( .A(n12491), .B(n12492), .S(n10216), .Z(n10069) );
  OR2_X1 U12527 ( .A1(n11087), .A2(n10265), .ZN(n10074) );
  OAI21_X1 U12528 ( .B1(n10071), .B2(P1_IR_REG_13__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10072) );
  XNOR2_X1 U12529 ( .A(n10072), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11264) );
  AOI22_X1 U12530 ( .A1(n11264), .A2(n10136), .B1(n10298), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n10073) );
  NAND2_X1 U12531 ( .A1(n10076), .A2(n10075), .ZN(n10077) );
  NAND2_X1 U12532 ( .A1(n10088), .A2(n10077), .ZN(n14869) );
  OR2_X1 U12533 ( .A1(n14869), .A2(n10278), .ZN(n10082) );
  NAND2_X1 U12534 ( .A1(n9893), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n10079) );
  INV_X1 U12535 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n15528) );
  OR2_X1 U12536 ( .A1(n9927), .A2(n15528), .ZN(n10078) );
  AND2_X1 U12537 ( .A1(n10079), .A2(n10078), .ZN(n10081) );
  INV_X1 U12538 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11265) );
  OR2_X1 U12539 ( .A1(n9861), .A2(n11265), .ZN(n10080) );
  XNOR2_X1 U12540 ( .A(n12672), .B(n12670), .ZN(n12259) );
  NAND2_X1 U12541 ( .A1(n10084), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10085) );
  XNOR2_X1 U12542 ( .A(n10085), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11965) );
  AOI22_X1 U12543 ( .A1(n10298), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n10136), 
        .B2(n11965), .ZN(n10086) );
  AND2_X1 U12544 ( .A1(n10088), .A2(n10087), .ZN(n10089) );
  OR2_X1 U12545 ( .A1(n10089), .A2(n10094), .ZN(n14485) );
  AOI22_X1 U12546 ( .A1(n6549), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9893), .B2(
        P1_REG0_REG_15__SCAN_IN), .ZN(n10091) );
  INV_X1 U12547 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n15527) );
  OR2_X1 U12548 ( .A1(n9927), .A2(n15527), .ZN(n10090) );
  OAI211_X1 U12549 ( .C1(n14485), .C2(n10278), .A(n10091), .B(n10090), .ZN(
        n14097) );
  INV_X1 U12550 ( .A(n14097), .ZN(n14461) );
  NAND2_X1 U12551 ( .A1(n14595), .A2(n14461), .ZN(n10310) );
  NAND2_X1 U12552 ( .A1(n12672), .A2(n12670), .ZN(n12548) );
  NAND2_X1 U12553 ( .A1(n10310), .A2(n12548), .ZN(n10092) );
  OR2_X1 U12554 ( .A1(n12672), .A2(n12670), .ZN(n12550) );
  MUX2_X1 U12555 ( .A(n10310), .B(n12552), .S(n10301), .Z(n10093) );
  NOR2_X1 U12556 ( .A1(n10094), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10095) );
  OR2_X1 U12557 ( .A1(n10115), .A2(n10095), .ZN(n14469) );
  AOI22_X1 U12558 ( .A1(n6549), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n10260), 
        .B2(P1_REG1_REG_16__SCAN_IN), .ZN(n10097) );
  INV_X1 U12559 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n15445) );
  OR2_X1 U12560 ( .A1(n10257), .A2(n15445), .ZN(n10096) );
  OAI211_X1 U12561 ( .C1(n14469), .C2(n10278), .A(n10097), .B(n10096), .ZN(
        n14478) );
  NAND2_X1 U12562 ( .A1(n11181), .A2(n10237), .ZN(n10104) );
  OR2_X1 U12563 ( .A1(n10084), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n10099) );
  NAND2_X1 U12564 ( .A1(n10099), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10098) );
  INV_X1 U12565 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n10100) );
  MUX2_X1 U12566 ( .A(n10098), .B(P1_IR_REG_31__SCAN_IN), .S(n10100), .Z(
        n10102) );
  INV_X1 U12567 ( .A(n10099), .ZN(n10101) );
  NAND2_X1 U12568 ( .A1(n10101), .A2(n10100), .ZN(n10109) );
  NAND2_X1 U12569 ( .A1(n10102), .A2(n10109), .ZN(n12151) );
  INV_X1 U12570 ( .A(n12151), .ZN(n12155) );
  AOI22_X1 U12571 ( .A1(n10298), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n10136), 
        .B2(n12155), .ZN(n10103) );
  MUX2_X1 U12572 ( .A(n14478), .B(n14591), .S(n10216), .Z(n10106) );
  INV_X1 U12573 ( .A(n14478), .ZN(n14447) );
  INV_X1 U12574 ( .A(n14591), .ZN(n14468) );
  MUX2_X1 U12575 ( .A(n14447), .B(n14468), .S(n10301), .Z(n10105) );
  NAND2_X1 U12576 ( .A1(n10107), .A2(n10106), .ZN(n10123) );
  NAND2_X1 U12577 ( .A1(n11233), .A2(n10237), .ZN(n10114) );
  NAND2_X1 U12578 ( .A1(n10109), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10108) );
  MUX2_X1 U12579 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10108), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n10112) );
  INV_X1 U12580 ( .A(n10109), .ZN(n10111) );
  INV_X1 U12581 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n10110) );
  NAND2_X1 U12582 ( .A1(n10111), .A2(n10110), .ZN(n10126) );
  NAND2_X1 U12583 ( .A1(n10112), .A2(n10126), .ZN(n12163) );
  INV_X1 U12584 ( .A(n12163), .ZN(n12278) );
  AOI22_X1 U12585 ( .A1(n10298), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n10136), 
        .B2(n12278), .ZN(n10113) );
  OR2_X1 U12586 ( .A1(n10115), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10116) );
  AND2_X1 U12587 ( .A1(n10141), .A2(n10116), .ZN(n14442) );
  NAND2_X1 U12588 ( .A1(n14442), .A2(n10179), .ZN(n10121) );
  INV_X1 U12589 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n12152) );
  NAND2_X1 U12590 ( .A1(n10260), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n10118) );
  INV_X1 U12591 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n15598) );
  OR2_X1 U12592 ( .A1(n10257), .A2(n15598), .ZN(n10117) );
  OAI211_X1 U12593 ( .C1(n9861), .C2(n12152), .A(n10118), .B(n10117), .ZN(
        n10119) );
  INV_X1 U12594 ( .A(n10119), .ZN(n10120) );
  NAND2_X1 U12595 ( .A1(n14585), .A2(n14463), .ZN(n10124) );
  OR2_X1 U12596 ( .A1(n14585), .A2(n14463), .ZN(n12557) );
  MUX2_X1 U12597 ( .A(n10124), .B(n12557), .S(n10301), .Z(n10122) );
  MUX2_X1 U12598 ( .A(n10124), .B(n12557), .S(n10216), .Z(n10125) );
  NAND2_X1 U12599 ( .A1(n11465), .A2(n10237), .ZN(n10130) );
  NAND2_X1 U12600 ( .A1(n10126), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10127) );
  MUX2_X1 U12601 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10127), .S(
        P1_IR_REG_18__SCAN_IN), .Z(n10128) );
  AOI22_X1 U12602 ( .A1(n10298), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n14222), 
        .B2(n10136), .ZN(n10129) );
  XNOR2_X1 U12603 ( .A(n10141), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n14431) );
  NAND2_X1 U12604 ( .A1(n14431), .A2(n10179), .ZN(n10135) );
  INV_X1 U12605 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14224) );
  NAND2_X1 U12606 ( .A1(n9893), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n10132) );
  NAND2_X1 U12607 ( .A1(n10260), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n10131) );
  OAI211_X1 U12608 ( .C1(n9861), .C2(n14224), .A(n10132), .B(n10131), .ZN(
        n10133) );
  INV_X1 U12609 ( .A(n10133), .ZN(n10134) );
  NAND2_X1 U12610 ( .A1(n10135), .A2(n10134), .ZN(n14408) );
  NAND2_X1 U12611 ( .A1(n14580), .A2(n14408), .ZN(n12580) );
  NAND2_X1 U12612 ( .A1(n11628), .A2(n10237), .ZN(n10138) );
  AOI22_X1 U12613 ( .A1(n10298), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n11311), 
        .B2(n10136), .ZN(n10137) );
  INV_X1 U12614 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n10140) );
  INV_X1 U12615 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n10139) );
  OAI21_X1 U12616 ( .B1(n10141), .B2(n10140), .A(n10139), .ZN(n10142) );
  NAND2_X1 U12617 ( .A1(n10142), .A2(n10155), .ZN(n14411) );
  OR2_X1 U12618 ( .A1(n14411), .A2(n10278), .ZN(n10147) );
  INV_X1 U12619 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n15675) );
  NAND2_X1 U12620 ( .A1(n6549), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n10144) );
  NAND2_X1 U12621 ( .A1(n9893), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n10143) );
  OAI211_X1 U12622 ( .C1(n9927), .C2(n15675), .A(n10144), .B(n10143), .ZN(
        n10145) );
  INV_X1 U12623 ( .A(n10145), .ZN(n10146) );
  NAND2_X1 U12624 ( .A1(n10147), .A2(n10146), .ZN(n14096) );
  XNOR2_X1 U12625 ( .A(n14574), .B(n14096), .ZN(n14415) );
  OAI21_X1 U12626 ( .B1(n10149), .B2(n12580), .A(n14415), .ZN(n10151) );
  NOR2_X1 U12627 ( .A1(n14580), .A2(n14408), .ZN(n12581) );
  MUX2_X1 U12628 ( .A(n14408), .B(n14580), .S(n10301), .Z(n10148) );
  NAND2_X1 U12629 ( .A1(n14096), .A2(n10216), .ZN(n10153) );
  INV_X1 U12630 ( .A(n14096), .ZN(n14427) );
  NAND2_X1 U12631 ( .A1(n14427), .A2(n10301), .ZN(n10152) );
  MUX2_X1 U12632 ( .A(n10153), .B(n10152), .S(n14574), .Z(n10154) );
  NAND2_X1 U12633 ( .A1(n10155), .A2(n14043), .ZN(n10156) );
  NAND2_X1 U12634 ( .A1(n10166), .A2(n10156), .ZN(n14046) );
  INV_X1 U12635 ( .A(n14046), .ZN(n14397) );
  NAND2_X1 U12636 ( .A1(n14397), .A2(n10179), .ZN(n10161) );
  INV_X1 U12637 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n15555) );
  NAND2_X1 U12638 ( .A1(n10260), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n10158) );
  NAND2_X1 U12639 ( .A1(n6549), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n10157) );
  OAI211_X1 U12640 ( .C1(n10257), .C2(n15555), .A(n10158), .B(n10157), .ZN(
        n10159) );
  INV_X1 U12641 ( .A(n10159), .ZN(n10160) );
  NAND2_X1 U12642 ( .A1(n11896), .A2(n10237), .ZN(n10163) );
  NAND2_X1 U12643 ( .A1(n10298), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n10162) );
  MUX2_X1 U12644 ( .A(n13992), .B(n14401), .S(n10216), .Z(n10165) );
  MUX2_X1 U12645 ( .A(n14409), .B(n14566), .S(n10301), .Z(n10164) );
  OR2_X1 U12646 ( .A1(n7947), .A2(n10176), .ZN(n14378) );
  INV_X1 U12647 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n10169) );
  NAND2_X1 U12648 ( .A1(n10260), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n10168) );
  INV_X1 U12649 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n15617) );
  OR2_X1 U12650 ( .A1(n10257), .A2(n15617), .ZN(n10167) );
  OAI211_X1 U12651 ( .C1(n9861), .C2(n10169), .A(n10168), .B(n10167), .ZN(
        n10170) );
  INV_X1 U12652 ( .A(n10170), .ZN(n10171) );
  OR2_X1 U12653 ( .A1(n12052), .A2(n10265), .ZN(n10173) );
  NAND2_X1 U12654 ( .A1(n10298), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n10172) );
  MUX2_X1 U12655 ( .A(n14359), .B(n14381), .S(n10301), .Z(n10175) );
  MUX2_X1 U12656 ( .A(n14381), .B(n14359), .S(n10301), .Z(n10174) );
  OR2_X1 U12657 ( .A1(n10176), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n10178) );
  AND2_X1 U12658 ( .A1(n10178), .A2(n10177), .ZN(n14366) );
  NAND2_X1 U12659 ( .A1(n14366), .A2(n10179), .ZN(n10185) );
  INV_X1 U12660 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n10182) );
  NAND2_X1 U12661 ( .A1(n9893), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n10181) );
  NAND2_X1 U12662 ( .A1(n10260), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n10180) );
  OAI211_X1 U12663 ( .C1(n9861), .C2(n10182), .A(n10181), .B(n10180), .ZN(
        n10183) );
  INV_X1 U12664 ( .A(n10183), .ZN(n10184) );
  NAND2_X1 U12665 ( .A1(n10185), .A2(n10184), .ZN(n14095) );
  OR2_X1 U12666 ( .A1(n10186), .A2(n6546), .ZN(n10187) );
  MUX2_X1 U12667 ( .A(n14095), .B(n14551), .S(n10216), .Z(n10191) );
  NAND2_X1 U12668 ( .A1(n10190), .A2(n10191), .ZN(n10189) );
  MUX2_X1 U12669 ( .A(n14095), .B(n14551), .S(n10301), .Z(n10188) );
  NAND2_X1 U12670 ( .A1(n10189), .A2(n10188), .ZN(n10195) );
  INV_X1 U12671 ( .A(n10190), .ZN(n10193) );
  INV_X1 U12672 ( .A(n10191), .ZN(n10192) );
  NAND2_X1 U12673 ( .A1(n9893), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n10201) );
  NAND2_X1 U12674 ( .A1(n6549), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n10200) );
  NAND2_X1 U12675 ( .A1(n10260), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n10199) );
  OAI21_X1 U12676 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n10197), .A(n10196), 
        .ZN(n14348) );
  OR2_X1 U12677 ( .A1(n10278), .A2(n14348), .ZN(n10198) );
  NAND4_X1 U12678 ( .A1(n10201), .A2(n10200), .A3(n10199), .A4(n10198), .ZN(
        n14358) );
  NAND2_X1 U12679 ( .A1(n12402), .A2(n9867), .ZN(n10203) );
  NAND2_X1 U12680 ( .A1(n10298), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n10202) );
  MUX2_X1 U12681 ( .A(n14358), .B(n14352), .S(n10301), .Z(n10206) );
  MUX2_X1 U12682 ( .A(n14352), .B(n14358), .S(n10301), .Z(n10204) );
  INV_X1 U12683 ( .A(n10206), .ZN(n10207) );
  NAND2_X1 U12684 ( .A1(n13965), .A2(n9867), .ZN(n10209) );
  NAND2_X1 U12685 ( .A1(n10298), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n10208) );
  NAND2_X1 U12686 ( .A1(n6549), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n10215) );
  NAND2_X1 U12687 ( .A1(n9893), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n10214) );
  NAND2_X1 U12688 ( .A1(n10260), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n10213) );
  OAI21_X1 U12689 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n10211), .A(n10210), 
        .ZN(n14335) );
  OR2_X1 U12690 ( .A1(n10278), .A2(n14335), .ZN(n10212) );
  NAND4_X1 U12691 ( .A1(n10215), .A2(n10214), .A3(n10213), .A4(n10212), .ZN(
        n14094) );
  MUX2_X1 U12692 ( .A(n14334), .B(n14094), .S(n10301), .Z(n10218) );
  MUX2_X1 U12693 ( .A(n14334), .B(n14094), .S(n10216), .Z(n10217) );
  INV_X1 U12694 ( .A(n10218), .ZN(n10219) );
  NAND2_X1 U12695 ( .A1(n10221), .A2(n10220), .ZN(n10231) );
  NAND2_X1 U12696 ( .A1(n9893), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n10227) );
  NAND2_X1 U12697 ( .A1(n6549), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n10226) );
  NAND2_X1 U12698 ( .A1(n10260), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n10225) );
  OAI21_X1 U12699 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n10223), .A(n10222), 
        .ZN(n14315) );
  OR2_X1 U12700 ( .A1(n10278), .A2(n14315), .ZN(n10224) );
  NAND4_X1 U12701 ( .A1(n10227), .A2(n10226), .A3(n10225), .A4(n10224), .ZN(
        n14325) );
  NAND2_X1 U12702 ( .A1(n12794), .A2(n9867), .ZN(n10229) );
  NAND2_X1 U12703 ( .A1(n10298), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n10228) );
  MUX2_X1 U12704 ( .A(n14325), .B(n14535), .S(n10301), .Z(n10230) );
  MUX2_X1 U12705 ( .A(n14535), .B(n14325), .S(n10301), .Z(n10232) );
  INV_X1 U12706 ( .A(n14297), .ZN(n10307) );
  MUX2_X1 U12707 ( .A(n7446), .B(n10307), .S(n10301), .Z(n10233) );
  INV_X1 U12708 ( .A(n10250), .ZN(n10253) );
  NAND2_X1 U12709 ( .A1(n13954), .A2(n10237), .ZN(n10239) );
  NAND2_X1 U12710 ( .A1(n10298), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n10238) );
  NAND2_X1 U12711 ( .A1(n6549), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n10247) );
  INV_X1 U12712 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10240) );
  OR2_X1 U12713 ( .A1(n10257), .A2(n10240), .ZN(n10246) );
  INV_X1 U12714 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n13974) );
  NAND2_X1 U12715 ( .A1(n10241), .A2(n13974), .ZN(n10242) );
  NAND2_X1 U12716 ( .A1(n10276), .A2(n10242), .ZN(n14283) );
  INV_X1 U12717 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10243) );
  OR2_X1 U12718 ( .A1(n9927), .A2(n10243), .ZN(n10244) );
  MUX2_X1 U12719 ( .A(n14286), .B(n14076), .S(n10301), .Z(n10249) );
  INV_X1 U12720 ( .A(n10249), .ZN(n10252) );
  MUX2_X1 U12721 ( .A(n14301), .B(n14522), .S(n10301), .Z(n10248) );
  INV_X1 U12722 ( .A(n10256), .ZN(n10287) );
  INV_X1 U12723 ( .A(n14274), .ZN(n14266) );
  MUX2_X1 U12724 ( .A(n14266), .B(n14517), .S(n10301), .Z(n10254) );
  INV_X1 U12725 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n15540) );
  NAND2_X1 U12726 ( .A1(n6549), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n10259) );
  INV_X1 U12727 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n15630) );
  OR2_X1 U12728 ( .A1(n10257), .A2(n15630), .ZN(n10258) );
  OAI211_X1 U12729 ( .C1(n9927), .C2(n15540), .A(n10259), .B(n10258), .ZN(
        n14246) );
  INV_X1 U12730 ( .A(n11897), .ZN(n10303) );
  NAND2_X1 U12731 ( .A1(n10700), .A2(n10303), .ZN(n10371) );
  INV_X1 U12732 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n10263) );
  NAND2_X1 U12733 ( .A1(n10260), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n10262) );
  NAND2_X1 U12734 ( .A1(n9893), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n10261) );
  OAI211_X1 U12735 ( .C1(n9861), .C2(n10263), .A(n10262), .B(n10261), .ZN(
        n14262) );
  OAI21_X1 U12736 ( .B1(n14246), .B2(n10371), .A(n14262), .ZN(n10264) );
  INV_X1 U12737 ( .A(n10264), .ZN(n10268) );
  OR2_X1 U12738 ( .A1(n14624), .A2(n10265), .ZN(n10267) );
  NAND2_X1 U12739 ( .A1(n10298), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n10266) );
  MUX2_X1 U12740 ( .A(n10268), .B(n14249), .S(n10301), .Z(n10292) );
  NAND2_X1 U12741 ( .A1(n10301), .A2(n14246), .ZN(n10271) );
  INV_X1 U12742 ( .A(n14262), .ZN(n10269) );
  AOI21_X1 U12743 ( .B1(n10271), .B2(n10270), .A(n10269), .ZN(n10272) );
  AOI21_X1 U12744 ( .B1(n14249), .B2(n10216), .A(n10272), .ZN(n10294) );
  NAND2_X1 U12745 ( .A1(n13948), .A2(n9867), .ZN(n10274) );
  NAND2_X1 U12746 ( .A1(n10298), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n10273) );
  NAND2_X1 U12747 ( .A1(n6549), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n10282) );
  INV_X1 U12748 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n15641) );
  OR2_X1 U12749 ( .A1(n9927), .A2(n15641), .ZN(n10281) );
  NAND2_X1 U12750 ( .A1(n9893), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n10280) );
  INV_X1 U12751 ( .A(n10276), .ZN(n10277) );
  NAND2_X1 U12752 ( .A1(n10277), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n14264) );
  OR2_X1 U12753 ( .A1(n10278), .A2(n14264), .ZN(n10279) );
  NAND4_X1 U12754 ( .A1(n10282), .A2(n10281), .A3(n10280), .A4(n10279), .ZN(
        n14093) );
  MUX2_X1 U12755 ( .A(n14261), .B(n14093), .S(n10301), .Z(n10290) );
  INV_X1 U12756 ( .A(n10290), .ZN(n10284) );
  MUX2_X1 U12757 ( .A(n14093), .B(n14261), .S(n10301), .Z(n10289) );
  AOI22_X1 U12758 ( .A1(n10292), .A2(n10294), .B1(n10284), .B2(n10289), .ZN(
        n10285) );
  INV_X1 U12759 ( .A(n10289), .ZN(n10291) );
  NAND2_X1 U12760 ( .A1(n10291), .A2(n10290), .ZN(n10295) );
  AOI21_X1 U12761 ( .B1(n10294), .B2(n10295), .A(n10292), .ZN(n10293) );
  NOR2_X1 U12762 ( .A1(n10295), .A2(n10294), .ZN(n10296) );
  NAND2_X1 U12763 ( .A1(n13942), .A2(n9867), .ZN(n10300) );
  NAND2_X1 U12764 ( .A1(n10298), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n10299) );
  NOR2_X1 U12765 ( .A1(n10344), .A2(n10301), .ZN(n10340) );
  NAND2_X1 U12766 ( .A1(n14640), .A2(n10700), .ZN(n11151) );
  NAND2_X1 U12767 ( .A1(n11151), .A2(n10705), .ZN(n10302) );
  OR2_X1 U12768 ( .A1(n11132), .A2(n14235), .ZN(n11329) );
  NAND2_X1 U12769 ( .A1(n10302), .A2(n11329), .ZN(n10341) );
  NAND2_X1 U12770 ( .A1(n12021), .A2(n10303), .ZN(n10714) );
  NAND2_X1 U12771 ( .A1(n10341), .A2(n10714), .ZN(n10343) );
  NAND2_X1 U12772 ( .A1(n10344), .A2(n10301), .ZN(n10350) );
  NOR2_X1 U12773 ( .A1(n10350), .A2(n14246), .ZN(n10304) );
  AOI211_X1 U12774 ( .C1(n10340), .C2(n14246), .A(n10343), .B(n10304), .ZN(
        n10305) );
  XOR2_X1 U12775 ( .A(n14246), .B(n10344), .Z(n10333) );
  NOR2_X1 U12776 ( .A1(n10333), .A2(n10341), .ZN(n10306) );
  XNOR2_X1 U12777 ( .A(n14249), .B(n14262), .ZN(n10330) );
  NAND2_X1 U12778 ( .A1(n10307), .A2(n14275), .ZN(n12565) );
  OR2_X1 U12779 ( .A1(n10307), .A2(n14275), .ZN(n10308) );
  INV_X1 U12780 ( .A(n14094), .ZN(n12748) );
  XNOR2_X1 U12781 ( .A(n14334), .B(n12748), .ZN(n14329) );
  XNOR2_X1 U12782 ( .A(n14352), .B(n14358), .ZN(n14344) );
  INV_X1 U12783 ( .A(n14095), .ZN(n10309) );
  XNOR2_X1 U12784 ( .A(n14381), .B(n14396), .ZN(n14374) );
  INV_X1 U12785 ( .A(n14415), .ZN(n14406) );
  NAND2_X1 U12786 ( .A1(n12552), .A2(n10310), .ZN(n14475) );
  XNOR2_X1 U12787 ( .A(n14591), .B(n14447), .ZN(n14459) );
  XNOR2_X1 U12788 ( .A(n12499), .B(n14098), .ZN(n12164) );
  INV_X1 U12789 ( .A(n14101), .ZN(n12321) );
  XNOR2_X1 U12790 ( .A(n14870), .B(n12321), .ZN(n12023) );
  XNOR2_X1 U12791 ( .A(n14952), .B(n14102), .ZN(n11935) );
  INV_X1 U12792 ( .A(n14103), .ZN(n12296) );
  OR2_X1 U12793 ( .A1(n14943), .A2(n12296), .ZN(n11885) );
  NAND2_X1 U12794 ( .A1(n14943), .A2(n12296), .ZN(n10311) );
  INV_X1 U12795 ( .A(n14105), .ZN(n10312) );
  NAND2_X1 U12796 ( .A1(n11719), .A2(n10312), .ZN(n11723) );
  OR2_X1 U12797 ( .A1(n11719), .A2(n10312), .ZN(n10313) );
  NAND2_X1 U12798 ( .A1(n11723), .A2(n10313), .ZN(n11717) );
  XNOR2_X1 U12799 ( .A(n15016), .B(n11595), .ZN(n15001) );
  XNOR2_X1 U12800 ( .A(n11587), .B(n14107), .ZN(n11318) );
  INV_X1 U12801 ( .A(n10314), .ZN(n10315) );
  AND2_X1 U12802 ( .A1(n11111), .A2(n10315), .ZN(n11081) );
  NAND4_X1 U12803 ( .A1(n10318), .A2(n11318), .A3(n11081), .A4(n10707), .ZN(
        n10319) );
  NOR3_X1 U12804 ( .A1(n11717), .A2(n15001), .A3(n10319), .ZN(n10320) );
  XNOR2_X1 U12805 ( .A(n11734), .B(n14104), .ZN(n14985) );
  NAND4_X1 U12806 ( .A1(n11935), .A2(n11722), .A3(n10320), .A4(n14985), .ZN(
        n10321) );
  NOR2_X1 U12807 ( .A1(n12023), .A2(n10321), .ZN(n10322) );
  XNOR2_X1 U12808 ( .A(n14892), .B(n14100), .ZN(n14891) );
  NAND4_X1 U12809 ( .A1(n12164), .A2(n10322), .A3(n12032), .A4(n14891), .ZN(
        n10323) );
  OR4_X1 U12810 ( .A1(n14475), .A2(n14459), .A3(n12259), .A4(n10323), .ZN(
        n10324) );
  INV_X1 U12811 ( .A(n14408), .ZN(n14448) );
  XNOR2_X1 U12812 ( .A(n14580), .B(n14448), .ZN(n14422) );
  XNOR2_X1 U12813 ( .A(n14585), .B(n14463), .ZN(n14445) );
  OR4_X1 U12814 ( .A1(n14406), .A2(n10324), .A3(n14422), .A4(n14445), .ZN(
        n10325) );
  NOR2_X1 U12815 ( .A1(n14374), .A2(n10325), .ZN(n10326) );
  XNOR2_X1 U12816 ( .A(n14566), .B(n14409), .ZN(n12586) );
  NAND4_X1 U12817 ( .A1(n14344), .A2(n14362), .A3(n10326), .A4(n12586), .ZN(
        n10327) );
  NOR2_X1 U12818 ( .A1(n14329), .A2(n10327), .ZN(n10329) );
  NAND2_X1 U12819 ( .A1(n14535), .A2(n14325), .ZN(n12593) );
  OR2_X1 U12820 ( .A1(n14535), .A2(n14325), .ZN(n10328) );
  NAND2_X1 U12821 ( .A1(n12593), .A2(n10328), .ZN(n14310) );
  NAND4_X1 U12822 ( .A1(n10330), .A2(n14300), .A3(n10329), .A4(n14310), .ZN(
        n10332) );
  NAND2_X1 U12823 ( .A1(n14517), .A2(n14274), .ZN(n14255) );
  OR2_X1 U12824 ( .A1(n14517), .A2(n14274), .ZN(n10331) );
  NAND2_X1 U12825 ( .A1(n14255), .A2(n10331), .ZN(n12595) );
  INV_X1 U12826 ( .A(n14093), .ZN(n12786) );
  XNOR2_X1 U12827 ( .A(n14261), .B(n12786), .ZN(n14257) );
  NOR3_X1 U12828 ( .A1(n10332), .A2(n12595), .A3(n14257), .ZN(n10335) );
  XNOR2_X1 U12829 ( .A(n14522), .B(n14301), .ZN(n12594) );
  INV_X1 U12830 ( .A(n10333), .ZN(n10334) );
  NAND3_X1 U12831 ( .A1(n10335), .A2(n12594), .A3(n10334), .ZN(n10336) );
  XNOR2_X1 U12832 ( .A(n10336), .B(n11311), .ZN(n10338) );
  INV_X1 U12833 ( .A(n10714), .ZN(n10337) );
  INV_X1 U12834 ( .A(n14246), .ZN(n10346) );
  INV_X1 U12835 ( .A(n10341), .ZN(n10339) );
  NAND2_X1 U12836 ( .A1(n10346), .A2(n10339), .ZN(n10349) );
  XOR2_X1 U12837 ( .A(n10341), .B(n10340), .Z(n10342) );
  NAND4_X1 U12838 ( .A1(n10342), .A2(n14504), .A3(n10714), .A4(n14246), .ZN(
        n10348) );
  INV_X1 U12839 ( .A(n10343), .ZN(n10345) );
  NAND4_X1 U12840 ( .A1(n10350), .A2(n10346), .A3(n10345), .A4(n10344), .ZN(
        n10347) );
  OAI211_X1 U12841 ( .C1(n10350), .C2(n10349), .A(n10348), .B(n10347), .ZN(
        n10351) );
  NAND2_X1 U12842 ( .A1(n10358), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10355) );
  INV_X1 U12843 ( .A(n10561), .ZN(n10356) );
  NAND2_X1 U12844 ( .A1(n10356), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12372) );
  INV_X1 U12845 ( .A(n10358), .ZN(n10359) );
  NAND2_X1 U12846 ( .A1(n10359), .A2(n10354), .ZN(n10362) );
  XNOR2_X1 U12847 ( .A(n10361), .B(n10360), .ZN(n10551) );
  INV_X1 U12848 ( .A(n10551), .ZN(n10370) );
  INV_X1 U12849 ( .A(n10364), .ZN(n10365) );
  MUX2_X1 U12850 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10367), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n10368) );
  NAND2_X1 U12851 ( .A1(n14640), .A2(n11311), .ZN(n10372) );
  INV_X1 U12852 ( .A(n11151), .ZN(n10562) );
  NAND2_X1 U12853 ( .A1(n15052), .A2(n10562), .ZN(n11499) );
  NAND2_X1 U12854 ( .A1(n11305), .A2(n11499), .ZN(n11157) );
  NOR3_X1 U12855 ( .A1(n11157), .A2(n14629), .A3(n14462), .ZN(n10375) );
  OAI21_X1 U12856 ( .B1(n12372), .B2(n14640), .A(P1_B_REG_SCAN_IN), .ZN(n10374) );
  OR2_X1 U12857 ( .A1(n10375), .A2(n10374), .ZN(n10376) );
  OAI21_X1 U12858 ( .B1(n12798), .B2(n13328), .A(n13069), .ZN(n10379) );
  XNOR2_X1 U12859 ( .A(n10379), .B(n6616), .ZN(n10381) );
  NAND2_X1 U12860 ( .A1(n10381), .A2(n10380), .ZN(n10386) );
  AND2_X1 U12861 ( .A1(n10735), .A2(P3_B_REG_SCAN_IN), .ZN(n10382) );
  OR2_X1 U12862 ( .A1(n15300), .A2(n10382), .ZN(n13052) );
  NOR2_X1 U12863 ( .A1(n11665), .A2(n13052), .ZN(n10384) );
  NOR2_X1 U12864 ( .A1(n12798), .A2(n15298), .ZN(n10383) );
  NOR2_X1 U12865 ( .A1(n13059), .A2(n10391), .ZN(n10409) );
  INV_X1 U12866 ( .A(n10393), .ZN(n13062) );
  INV_X1 U12867 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n10410) );
  INV_X1 U12868 ( .A(n10394), .ZN(n10395) );
  NAND2_X1 U12869 ( .A1(n10395), .A2(n10399), .ZN(n10949) );
  INV_X1 U12870 ( .A(n10396), .ZN(n11272) );
  INV_X1 U12871 ( .A(n10397), .ZN(n10398) );
  NAND2_X1 U12872 ( .A1(n11272), .A2(n10398), .ZN(n10944) );
  INV_X1 U12873 ( .A(n10399), .ZN(n10400) );
  NOR2_X1 U12874 ( .A1(n13377), .A2(n10400), .ZN(n10402) );
  NAND2_X1 U12875 ( .A1(n10402), .A2(n10401), .ZN(n10947) );
  INV_X1 U12876 ( .A(n10937), .ZN(n10403) );
  OAI22_X1 U12877 ( .A1(n10949), .A2(n10944), .B1(n10947), .B2(n10403), .ZN(
        n10404) );
  NAND2_X1 U12878 ( .A1(n10404), .A2(n10950), .ZN(n10408) );
  INV_X1 U12879 ( .A(n10949), .ZN(n10406) );
  NOR2_X1 U12880 ( .A1(n11281), .A2(n10405), .ZN(n10941) );
  NAND2_X1 U12881 ( .A1(n10406), .A2(n10941), .ZN(n10407) );
  NOR2_X1 U12882 ( .A1(n10413), .A2(n10412), .ZN(n10418) );
  INV_X1 U12883 ( .A(n12791), .ZN(n10414) );
  NOR2_X1 U12884 ( .A1(n11133), .A2(n10414), .ZN(P1_U4016) );
  INV_X2 U12885 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X2 U12886 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  AOI21_X1 U12887 ( .B1(n10416), .B2(n10415), .A(n8237), .ZN(n10417) );
  OR2_X1 U12888 ( .A1(n10418), .A2(n10417), .ZN(n10444) );
  NAND2_X1 U12889 ( .A1(n10419), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13952) );
  INV_X1 U12890 ( .A(n13952), .ZN(n10420) );
  NAND2_X1 U12891 ( .A1(n10444), .A2(n10420), .ZN(n10434) );
  XNOR2_X1 U12892 ( .A(n10730), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n10721) );
  NAND2_X1 U12893 ( .A1(n13531), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10423) );
  NAND2_X1 U12894 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n10421) );
  AOI21_X1 U12895 ( .B1(n13532), .B2(n8117), .A(n10421), .ZN(n10422) );
  NAND2_X1 U12896 ( .A1(n10423), .A2(n10422), .ZN(n13536) );
  NAND2_X1 U12897 ( .A1(n13536), .A2(n10423), .ZN(n10720) );
  NAND2_X1 U12898 ( .A1(n10721), .A2(n10720), .ZN(n10426) );
  OR2_X1 U12899 ( .A1(n10730), .A2(n10424), .ZN(n10425) );
  NAND2_X1 U12900 ( .A1(n10426), .A2(n10425), .ZN(n10449) );
  MUX2_X1 U12901 ( .A(n10428), .B(P2_REG1_REG_3__SCAN_IN), .S(n10492), .Z(
        n10427) );
  NAND2_X1 U12902 ( .A1(n10449), .A2(n10427), .ZN(n10450) );
  OR2_X1 U12903 ( .A1(n10492), .A2(n10428), .ZN(n10432) );
  NAND2_X1 U12904 ( .A1(n10450), .A2(n10432), .ZN(n10430) );
  MUX2_X1 U12905 ( .A(n10577), .B(P2_REG1_REG_4__SCAN_IN), .S(n10578), .Z(
        n10429) );
  NAND2_X1 U12906 ( .A1(n10430), .A2(n10429), .ZN(n10849) );
  MUX2_X1 U12907 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10577), .S(n10578), .Z(
        n10431) );
  NAND3_X1 U12908 ( .A1(n10450), .A2(n10432), .A3(n10431), .ZN(n10433) );
  AND3_X1 U12909 ( .A1(n15190), .A2(n10849), .A3(n10433), .ZN(n10448) );
  INV_X1 U12910 ( .A(n10434), .ZN(n10436) );
  INV_X1 U12911 ( .A(n15198), .ZN(n15129) );
  NOR3_X1 U12912 ( .A1(n13537), .A2(n13534), .A3(n10621), .ZN(n13538) );
  AOI21_X1 U12913 ( .B1(n13531), .B2(P2_REG2_REG_1__SCAN_IN), .A(n13538), .ZN(
        n10724) );
  MUX2_X1 U12914 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10437), .S(n10730), .Z(
        n10723) );
  NOR2_X1 U12915 ( .A1(n10724), .A2(n10723), .ZN(n10722) );
  NOR2_X1 U12916 ( .A1(n10730), .A2(n10437), .ZN(n10456) );
  MUX2_X1 U12917 ( .A(n12049), .B(P2_REG2_REG_3__SCAN_IN), .S(n10492), .Z(
        n10455) );
  OAI21_X1 U12918 ( .B1(n10722), .B2(n10456), .A(n10455), .ZN(n10454) );
  INV_X1 U12919 ( .A(n10492), .ZN(n10438) );
  NAND2_X1 U12920 ( .A1(n10438), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10440) );
  MUX2_X1 U12921 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11766), .S(n10578), .Z(
        n10439) );
  AND3_X1 U12922 ( .A1(n10454), .A2(n10440), .A3(n10439), .ZN(n10441) );
  OR2_X1 U12923 ( .A1(n10444), .A2(P2_U3088), .ZN(n15166) );
  INV_X1 U12924 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10442) );
  NAND2_X1 U12925 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n11404) );
  OAI21_X1 U12926 ( .B1(n15166), .B2(n10442), .A(n11404), .ZN(n10446) );
  AND2_X1 U12927 ( .A1(n8625), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10443) );
  NOR2_X1 U12928 ( .A1(n15204), .A2(n10578), .ZN(n10445) );
  OR4_X1 U12929 ( .A1(n10448), .A2(n10447), .A3(n10446), .A4(n10445), .ZN(
        P2_U3218) );
  INV_X1 U12930 ( .A(n10449), .ZN(n10453) );
  MUX2_X1 U12931 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10428), .S(n10492), .Z(
        n10452) );
  INV_X1 U12932 ( .A(n10450), .ZN(n10451) );
  AOI211_X1 U12933 ( .C1(n10453), .C2(n10452), .A(n10451), .B(n15136), .ZN(
        n10463) );
  INV_X1 U12934 ( .A(n10454), .ZN(n10458) );
  NOR3_X1 U12935 ( .A1(n10722), .A2(n10456), .A3(n10455), .ZN(n10457) );
  NOR3_X1 U12936 ( .A1(n15129), .A2(n10458), .A3(n10457), .ZN(n10462) );
  INV_X1 U12937 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10459) );
  OAI22_X1 U12938 ( .A1(n15166), .A2(n10459), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12042), .ZN(n10461) );
  NOR2_X1 U12939 ( .A1(n15204), .A2(n10492), .ZN(n10460) );
  OR4_X1 U12940 ( .A1(n10463), .A2(n10462), .A3(n10461), .A4(n10460), .ZN(
        P2_U3217) );
  INV_X1 U12941 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10998) );
  NAND2_X1 U12942 ( .A1(n10464), .A2(P3_U3151), .ZN(n10465) );
  OAI21_X1 U12943 ( .B1(n10998), .B2(P3_U3151), .A(n10465), .ZN(P3_U3295) );
  NOR2_X2 U12944 ( .A1(n6546), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14762) );
  INV_X1 U12945 ( .A(n14762), .ZN(n14743) );
  NAND2_X1 U12946 ( .A1(n10486), .A2(P3_U3151), .ZN(n14741) );
  OAI222_X1 U12947 ( .A1(n6781), .A2(P3_U3151), .B1(n14743), .B2(n10467), .C1(
        n10466), .C2(n14741), .ZN(P3_U3294) );
  OAI222_X1 U12948 ( .A1(P3_U3151), .A2(n11869), .B1(n14741), .B2(n10469), 
        .C1(n14743), .C2(n10468), .ZN(P3_U3287) );
  NAND2_X2 U12949 ( .A1(n7997), .A2(P1_U3086), .ZN(n14638) );
  OAI222_X1 U12950 ( .A1(n14635), .A2(n10470), .B1(n14638), .B2(n10487), .C1(
        P1_U3086), .C2(n10650), .ZN(P1_U3354) );
  AOI222_X1 U12951 ( .A1(n10471), .A2(n14762), .B1(SI_9_), .B2(n14761), .C1(
        n11913), .C2(P3_STATE_REG_SCAN_IN), .ZN(n10472) );
  INV_X1 U12952 ( .A(n10472), .ZN(P3_U3286) );
  AOI222_X1 U12953 ( .A1(n10473), .A2(n14762), .B1(SI_7_), .B2(n14761), .C1(
        n11219), .C2(P3_STATE_REG_SCAN_IN), .ZN(n10474) );
  INV_X1 U12954 ( .A(n10474), .ZN(P3_U3288) );
  AOI222_X1 U12955 ( .A1(n10475), .A2(n14762), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n7480), .C1(SI_5_), .C2(n14761), .ZN(n10476) );
  INV_X1 U12956 ( .A(n10476), .ZN(P3_U3290) );
  AOI222_X1 U12957 ( .A1(n10477), .A2(n14762), .B1(n10922), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_4_), .C2(n14761), .ZN(n10478) );
  INV_X1 U12958 ( .A(n10478), .ZN(P3_U3291) );
  INV_X1 U12959 ( .A(n10479), .ZN(n10494) );
  INV_X1 U12960 ( .A(n14129), .ZN(n10480) );
  OAI222_X1 U12961 ( .A1(n14635), .A2(n10481), .B1(n14638), .B2(n10494), .C1(
        P1_U3086), .C2(n10480), .ZN(P1_U3353) );
  INV_X1 U12962 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10484) );
  INV_X1 U12963 ( .A(n10482), .ZN(n10489) );
  INV_X1 U12964 ( .A(n10798), .ZN(n10483) );
  OAI222_X1 U12965 ( .A1(n14635), .A2(n10484), .B1(n14638), .B2(n10489), .C1(
        P1_U3086), .C2(n10483), .ZN(P1_U3350) );
  NOR2_X1 U12966 ( .A1(n10486), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13945) );
  INV_X2 U12967 ( .A(n13945), .ZN(n13964) );
  NAND2_X1 U12968 ( .A1(n10486), .A2(P2_U3088), .ZN(n13967) );
  OAI222_X1 U12969 ( .A1(n13964), .A2(n10488), .B1(n12649), .B2(n10487), .C1(
        P2_U3088), .C2(n13532), .ZN(P2_U3326) );
  OAI222_X1 U12970 ( .A1(n13964), .A2(n10490), .B1(n13967), .B2(n10489), .C1(
        P2_U3088), .C2(n10860), .ZN(P2_U3322) );
  INV_X1 U12971 ( .A(n10491), .ZN(n10506) );
  OAI222_X1 U12972 ( .A1(n13964), .A2(n10493), .B1(n13967), .B2(n10506), .C1(
        P2_U3088), .C2(n10492), .ZN(P2_U3324) );
  OAI222_X1 U12973 ( .A1(n13964), .A2(n10495), .B1(n13967), .B2(n10494), .C1(
        P2_U3088), .C2(n10730), .ZN(P2_U3325) );
  INV_X1 U12974 ( .A(n10496), .ZN(n10500) );
  OAI222_X1 U12975 ( .A1(n13964), .A2(n10497), .B1(n13967), .B2(n10500), .C1(
        P2_U3088), .C2(n10578), .ZN(P2_U3323) );
  INV_X1 U12976 ( .A(n10498), .ZN(n10503) );
  OAI222_X1 U12977 ( .A1(n13964), .A2(n10499), .B1(n13967), .B2(n10503), .C1(
        P2_U3088), .C2(n10874), .ZN(P2_U3321) );
  INV_X1 U12978 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10501) );
  INV_X1 U12979 ( .A(n14161), .ZN(n14153) );
  OAI222_X1 U12980 ( .A1(n14635), .A2(n10501), .B1(n14638), .B2(n10500), .C1(
        P1_U3086), .C2(n14153), .ZN(P1_U3351) );
  INV_X1 U12981 ( .A(n14179), .ZN(n10502) );
  OAI222_X1 U12982 ( .A1(n14635), .A2(n10504), .B1(n14638), .B2(n10503), .C1(
        P1_U3086), .C2(n10502), .ZN(P1_U3349) );
  INV_X1 U12983 ( .A(n14148), .ZN(n10505) );
  OAI222_X1 U12984 ( .A1(n14635), .A2(n10507), .B1(n14638), .B2(n10506), .C1(
        P1_U3086), .C2(n10505), .ZN(P1_U3352) );
  INV_X1 U12985 ( .A(n10508), .ZN(n10510) );
  INV_X1 U12986 ( .A(n14635), .ZN(n14620) );
  AOI22_X1 U12987 ( .A1(n14194), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n14620), .ZN(n10509) );
  OAI21_X1 U12988 ( .B1(n10510), .B2(n14638), .A(n10509), .ZN(P1_U3348) );
  OAI222_X1 U12989 ( .A1(n13964), .A2(n10511), .B1(n13967), .B2(n10510), .C1(
        P2_U3088), .C2(n10602), .ZN(P2_U3320) );
  INV_X1 U12990 ( .A(n10512), .ZN(n10515) );
  AOI22_X1 U12991 ( .A1(n14205), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n14620), .ZN(n10513) );
  OAI21_X1 U12992 ( .B1(n10515), .B2(n14638), .A(n10513), .ZN(P1_U3347) );
  INV_X1 U12993 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10516) );
  INV_X1 U12994 ( .A(n10669), .ZN(n10514) );
  OAI222_X1 U12995 ( .A1(n13964), .A2(n10516), .B1(n13967), .B2(n10515), .C1(
        P2_U3088), .C2(n10514), .ZN(P2_U3319) );
  INV_X1 U12996 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10517) );
  INV_X1 U12997 ( .A(n10814), .ZN(n10817) );
  OAI222_X1 U12998 ( .A1(n13964), .A2(n10517), .B1(n13967), .B2(n10518), .C1(
        n10817), .C2(P2_U3088), .ZN(P2_U3318) );
  INV_X1 U12999 ( .A(n10976), .ZN(n10970) );
  OAI222_X1 U13000 ( .A1(n14635), .A2(n10519), .B1(n14638), .B2(n10518), .C1(
        n10970), .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U13001 ( .A(n10520), .ZN(n10521) );
  NOR2_X1 U13002 ( .A1(n10521), .A2(n13378), .ZN(n10523) );
  CLKBUF_X1 U13003 ( .A(n10523), .Z(n10548) );
  INV_X1 U13004 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10522) );
  NOR2_X1 U13005 ( .A1(n10548), .A2(n10522), .ZN(P3_U3252) );
  INV_X1 U13006 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10524) );
  NOR2_X1 U13007 ( .A1(n10548), .A2(n10524), .ZN(P3_U3258) );
  INV_X1 U13008 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10525) );
  NOR2_X1 U13009 ( .A1(n10548), .A2(n10525), .ZN(P3_U3256) );
  INV_X1 U13010 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10526) );
  NOR2_X1 U13011 ( .A1(n10548), .A2(n10526), .ZN(P3_U3249) );
  INV_X1 U13012 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10527) );
  NOR2_X1 U13013 ( .A1(n10548), .A2(n10527), .ZN(P3_U3255) );
  INV_X1 U13014 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10528) );
  NOR2_X1 U13015 ( .A1(n10548), .A2(n10528), .ZN(P3_U3254) );
  INV_X1 U13016 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10529) );
  NOR2_X1 U13017 ( .A1(n10548), .A2(n10529), .ZN(P3_U3253) );
  INV_X1 U13018 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10530) );
  NOR2_X1 U13019 ( .A1(n10523), .A2(n10530), .ZN(P3_U3262) );
  INV_X1 U13020 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10531) );
  NOR2_X1 U13021 ( .A1(n10548), .A2(n10531), .ZN(P3_U3251) );
  INV_X1 U13022 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10532) );
  NOR2_X1 U13023 ( .A1(n10548), .A2(n10532), .ZN(P3_U3257) );
  INV_X1 U13024 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10533) );
  NOR2_X1 U13025 ( .A1(n10548), .A2(n10533), .ZN(P3_U3259) );
  INV_X1 U13026 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10534) );
  NOR2_X1 U13027 ( .A1(n10523), .A2(n10534), .ZN(P3_U3241) );
  INV_X1 U13028 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n15472) );
  NOR2_X1 U13029 ( .A1(n10523), .A2(n15472), .ZN(P3_U3240) );
  INV_X1 U13030 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10535) );
  NOR2_X1 U13031 ( .A1(n10523), .A2(n10535), .ZN(P3_U3239) );
  INV_X1 U13032 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10536) );
  NOR2_X1 U13033 ( .A1(n10523), .A2(n10536), .ZN(P3_U3238) );
  INV_X1 U13034 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10537) );
  NOR2_X1 U13035 ( .A1(n10523), .A2(n10537), .ZN(P3_U3237) );
  INV_X1 U13036 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10538) );
  NOR2_X1 U13037 ( .A1(n10523), .A2(n10538), .ZN(P3_U3236) );
  INV_X1 U13038 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n15603) );
  NOR2_X1 U13039 ( .A1(n10523), .A2(n15603), .ZN(P3_U3235) );
  INV_X1 U13040 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n15710) );
  NOR2_X1 U13041 ( .A1(n10523), .A2(n15710), .ZN(P3_U3234) );
  INV_X1 U13042 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10539) );
  NOR2_X1 U13043 ( .A1(n10548), .A2(n10539), .ZN(P3_U3250) );
  INV_X1 U13044 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10540) );
  NOR2_X1 U13045 ( .A1(n10523), .A2(n10540), .ZN(P3_U3242) );
  INV_X1 U13046 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10541) );
  NOR2_X1 U13047 ( .A1(n10548), .A2(n10541), .ZN(P3_U3248) );
  INV_X1 U13048 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10542) );
  NOR2_X1 U13049 ( .A1(n10548), .A2(n10542), .ZN(P3_U3247) );
  INV_X1 U13050 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10543) );
  NOR2_X1 U13051 ( .A1(n10548), .A2(n10543), .ZN(P3_U3246) );
  INV_X1 U13052 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10544) );
  NOR2_X1 U13053 ( .A1(n10523), .A2(n10544), .ZN(P3_U3245) );
  INV_X1 U13054 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10545) );
  NOR2_X1 U13055 ( .A1(n10548), .A2(n10545), .ZN(P3_U3244) );
  INV_X1 U13056 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10546) );
  NOR2_X1 U13057 ( .A1(n10548), .A2(n10546), .ZN(P3_U3243) );
  INV_X1 U13058 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n15602) );
  NOR2_X1 U13059 ( .A1(n10548), .A2(n15602), .ZN(P3_U3261) );
  INV_X1 U13060 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10547) );
  NOR2_X1 U13061 ( .A1(n10548), .A2(n10547), .ZN(P3_U3263) );
  INV_X1 U13062 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10549) );
  NOR2_X1 U13063 ( .A1(n10548), .A2(n10549), .ZN(P3_U3260) );
  INV_X1 U13064 ( .A(n10550), .ZN(n14639) );
  NAND3_X1 U13065 ( .A1(n14639), .A2(n10551), .A3(P1_B_REG_SCAN_IN), .ZN(
        n10553) );
  INV_X1 U13066 ( .A(P1_B_REG_SCAN_IN), .ZN(n14244) );
  AOI21_X1 U13067 ( .B1(n10550), .B2(n14244), .A(n14634), .ZN(n10552) );
  NAND2_X1 U13068 ( .A1(n10553), .A2(n10552), .ZN(n10831) );
  NAND2_X1 U13069 ( .A1(n11305), .A2(n10831), .ZN(n15022) );
  INV_X1 U13070 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10828) );
  INV_X1 U13071 ( .A(n10832), .ZN(n10555) );
  AOI22_X1 U13072 ( .A1(n15022), .A2(n10828), .B1(n12791), .B2(n10555), .ZN(
        P1_U3445) );
  NAND2_X1 U13073 ( .A1(n15114), .A2(P2_U3947), .ZN(n10556) );
  OAI21_X1 U13074 ( .B1(n10065), .B2(P2_U3947), .A(n10556), .ZN(P2_U3544) );
  INV_X1 U13075 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n15458) );
  NAND2_X1 U13076 ( .A1(n15344), .A2(P3_U3897), .ZN(n10557) );
  OAI21_X1 U13077 ( .B1(P3_U3897), .B2(n15458), .A(n10557), .ZN(P3_U3492) );
  INV_X1 U13078 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n15597) );
  NAND2_X1 U13079 ( .A1(n15423), .A2(P3_U3897), .ZN(n10558) );
  OAI21_X1 U13080 ( .B1(P3_U3897), .B2(n15597), .A(n10558), .ZN(P3_U3493) );
  OAI222_X1 U13081 ( .A1(P3_U3151), .A2(n12924), .B1(n14741), .B2(n10560), 
        .C1(n14743), .C2(n10559), .ZN(P3_U3282) );
  INV_X1 U13082 ( .A(n11305), .ZN(n11160) );
  NAND2_X1 U13083 ( .A1(n11160), .A2(n12372), .ZN(n10646) );
  NAND2_X1 U13084 ( .A1(n10562), .A2(n10561), .ZN(n10564) );
  NAND2_X1 U13085 ( .A1(n10564), .A2(n10563), .ZN(n10644) );
  NAND2_X1 U13086 ( .A1(n10646), .A2(n10644), .ZN(n14980) );
  INV_X1 U13087 ( .A(n14980), .ZN(n14212) );
  NOR2_X1 U13088 ( .A1(n14212), .A2(n6551), .ZN(P1_U3085) );
  INV_X1 U13089 ( .A(n11002), .ZN(n10985) );
  INV_X1 U13090 ( .A(n10565), .ZN(n10567) );
  OAI222_X1 U13091 ( .A1(P1_U3086), .A2(n10985), .B1(n14635), .B2(n10566), 
        .C1(n14638), .C2(n10567), .ZN(P1_U3345) );
  INV_X1 U13092 ( .A(n11040), .ZN(n10824) );
  INV_X1 U13093 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10568) );
  OAI222_X1 U13094 ( .A1(P2_U3088), .A2(n10824), .B1(n13964), .B2(n10568), 
        .C1(n13967), .C2(n10567), .ZN(P2_U3317) );
  NAND2_X1 U13095 ( .A1(n6551), .A2(n11168), .ZN(n10569) );
  OAI21_X1 U13096 ( .B1(n6551), .B2(n8663), .A(n10569), .ZN(P1_U3560) );
  INV_X1 U13097 ( .A(n10570), .ZN(n10572) );
  INV_X1 U13098 ( .A(n11044), .ZN(n13563) );
  OAI222_X1 U13099 ( .A1(n13964), .A2(n10571), .B1(n12649), .B2(n10572), .C1(
        n13563), .C2(P2_U3088), .ZN(P2_U3316) );
  INV_X1 U13100 ( .A(n11024), .ZN(n11021) );
  OAI222_X1 U13101 ( .A1(n14635), .A2(n10573), .B1(n14638), .B2(n10572), .C1(
        n11021), .C2(P1_U3086), .ZN(P1_U3344) );
  INV_X1 U13102 ( .A(n10860), .ZN(n10582) );
  MUX2_X1 U13103 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11833), .S(n10860), .Z(
        n10853) );
  NOR2_X1 U13104 ( .A1(n10854), .A2(n10853), .ZN(n10852) );
  AOI21_X1 U13105 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n10582), .A(n10852), .ZN(
        n10868) );
  MUX2_X1 U13106 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11814), .S(n10874), .Z(
        n10867) );
  NOR2_X1 U13107 ( .A1(n10868), .A2(n10867), .ZN(n10866) );
  NOR2_X1 U13108 ( .A1(n10874), .A2(n11814), .ZN(n10575) );
  MUX2_X1 U13109 ( .A(n11847), .B(P2_REG2_REG_7__SCAN_IN), .S(n10602), .Z(
        n10574) );
  OAI21_X1 U13110 ( .B1(n10866), .B2(n10575), .A(n10574), .ZN(n10599) );
  OR3_X1 U13111 ( .A1(n10866), .A2(n10575), .A3(n10574), .ZN(n10576) );
  NAND3_X1 U13112 ( .A1(n10599), .A2(n15198), .A3(n10576), .ZN(n10595) );
  INV_X1 U13113 ( .A(n15204), .ZN(n15168) );
  INV_X1 U13114 ( .A(n10602), .ZN(n10596) );
  INV_X1 U13115 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14704) );
  NAND2_X1 U13116 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n11513) );
  OAI21_X1 U13117 ( .B1(n15166), .B2(n14704), .A(n11513), .ZN(n10593) );
  OR2_X1 U13118 ( .A1(n10578), .A2(n10577), .ZN(n10848) );
  NAND2_X1 U13119 ( .A1(n10849), .A2(n10848), .ZN(n10581) );
  MUX2_X1 U13120 ( .A(n10579), .B(P2_REG1_REG_5__SCAN_IN), .S(n10860), .Z(
        n10580) );
  NAND2_X1 U13121 ( .A1(n10581), .A2(n10580), .ZN(n10863) );
  NAND2_X1 U13122 ( .A1(n10582), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10862) );
  NAND2_X1 U13123 ( .A1(n10863), .A2(n10862), .ZN(n10585) );
  MUX2_X1 U13124 ( .A(n10583), .B(P2_REG1_REG_6__SCAN_IN), .S(n10874), .Z(
        n10584) );
  NAND2_X1 U13125 ( .A1(n10585), .A2(n10584), .ZN(n10865) );
  OR2_X1 U13126 ( .A1(n10874), .A2(n10583), .ZN(n10590) );
  NAND2_X1 U13127 ( .A1(n10865), .A2(n10590), .ZN(n10588) );
  INV_X1 U13128 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10586) );
  MUX2_X1 U13129 ( .A(n10586), .B(P2_REG1_REG_7__SCAN_IN), .S(n10602), .Z(
        n10587) );
  NAND2_X1 U13130 ( .A1(n10588), .A2(n10587), .ZN(n10608) );
  MUX2_X1 U13131 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10586), .S(n10602), .Z(
        n10589) );
  NAND3_X1 U13132 ( .A1(n10865), .A2(n10590), .A3(n10589), .ZN(n10591) );
  AND3_X1 U13133 ( .A1(n15190), .A2(n10608), .A3(n10591), .ZN(n10592) );
  AOI211_X1 U13134 ( .C1(n15168), .C2(n10596), .A(n10593), .B(n10592), .ZN(
        n10594) );
  NAND2_X1 U13135 ( .A1(n10595), .A2(n10594), .ZN(P2_U3221) );
  NAND2_X1 U13136 ( .A1(n10596), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10598) );
  MUX2_X1 U13137 ( .A(n11805), .B(P2_REG2_REG_8__SCAN_IN), .S(n10669), .Z(
        n10597) );
  AOI21_X1 U13138 ( .B1(n10599), .B2(n10598), .A(n10597), .ZN(n10668) );
  NAND3_X1 U13139 ( .A1(n10599), .A2(n10598), .A3(n10597), .ZN(n10600) );
  NAND2_X1 U13140 ( .A1(n10600), .A2(n15198), .ZN(n10613) );
  INV_X1 U13141 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10601) );
  NAND2_X1 U13142 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n11448) );
  OAI21_X1 U13143 ( .B1(n15166), .B2(n10601), .A(n11448), .ZN(n10611) );
  OR2_X1 U13144 ( .A1(n10602), .A2(n10586), .ZN(n10607) );
  NAND2_X1 U13145 ( .A1(n10608), .A2(n10607), .ZN(n10605) );
  INV_X1 U13146 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10603) );
  MUX2_X1 U13147 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10603), .S(n10669), .Z(
        n10604) );
  NAND2_X1 U13148 ( .A1(n10605), .A2(n10604), .ZN(n10667) );
  MUX2_X1 U13149 ( .A(n10603), .B(P2_REG1_REG_8__SCAN_IN), .S(n10669), .Z(
        n10606) );
  NAND3_X1 U13150 ( .A1(n10608), .A2(n10607), .A3(n10606), .ZN(n10609) );
  AND3_X1 U13151 ( .A1(n15190), .A2(n10667), .A3(n10609), .ZN(n10610) );
  AOI211_X1 U13152 ( .C1(n15168), .C2(n10669), .A(n10611), .B(n10610), .ZN(
        n10612) );
  OAI21_X1 U13153 ( .B1(n10668), .B2(n10613), .A(n10612), .ZN(P2_U3222) );
  INV_X1 U13154 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n15541) );
  NAND2_X1 U13155 ( .A1(n11983), .A2(P3_U3897), .ZN(n10614) );
  OAI21_X1 U13156 ( .B1(P3_U3897), .B2(n15541), .A(n10614), .ZN(P3_U3496) );
  INV_X1 U13157 ( .A(n10615), .ZN(n10616) );
  OAI222_X1 U13158 ( .A1(n13964), .A2(n15461), .B1(n12649), .B2(n10616), .C1(
        n15135), .C2(P2_U3088), .ZN(P2_U3315) );
  INV_X1 U13159 ( .A(n11246), .ZN(n11033) );
  OAI222_X1 U13160 ( .A1(n14635), .A2(n15628), .B1(n14638), .B2(n10616), .C1(
        n11033), .C2(P1_U3086), .ZN(P1_U3343) );
  OAI222_X1 U13161 ( .A1(P3_U3151), .A2(n12954), .B1(n14741), .B2(n10618), 
        .C1(n14743), .C2(n10617), .ZN(P3_U3281) );
  NAND2_X1 U13162 ( .A1(n15198), .A2(n10621), .ZN(n10619) );
  OAI211_X1 U13163 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n15136), .A(n10619), .B(
        n15204), .ZN(n10623) );
  OAI22_X1 U13164 ( .A1(n15129), .A2(n10621), .B1(n10620), .B2(n15136), .ZN(
        n10622) );
  MUX2_X1 U13165 ( .A(n10623), .B(n10622), .S(n13534), .Z(n10626) );
  INV_X1 U13166 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10624) );
  OAI22_X1 U13167 ( .A1(n15166), .A2(n10624), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11418), .ZN(n10625) );
  OR2_X1 U13168 ( .A1(n10626), .A2(n10625), .ZN(P2_U3214) );
  INV_X1 U13169 ( .A(n10627), .ZN(n10628) );
  OAI222_X1 U13170 ( .A1(P2_U3088), .A2(n15148), .B1(n12649), .B2(n10628), 
        .C1(n15654), .C2(n13964), .ZN(P2_U3314) );
  INV_X1 U13171 ( .A(n11261), .ZN(n11256) );
  OAI222_X1 U13172 ( .A1(P1_U3086), .A2(n11256), .B1(n14635), .B2(n10065), 
        .C1(n10628), .C2(n14638), .ZN(P1_U3342) );
  MUX2_X1 U13173 ( .A(n10629), .B(P1_REG1_REG_5__SCAN_IN), .S(n10798), .Z(
        n10643) );
  INV_X1 U13174 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10630) );
  MUX2_X1 U13175 ( .A(n10630), .B(P1_REG1_REG_1__SCAN_IN), .S(n10650), .Z(
        n14114) );
  AND2_X1 U13176 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14115) );
  NAND2_X1 U13177 ( .A1(n14114), .A2(n14115), .ZN(n14132) );
  NAND2_X1 U13178 ( .A1(n14113), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n14131) );
  NAND2_X1 U13179 ( .A1(n14132), .A2(n14131), .ZN(n10633) );
  MUX2_X1 U13180 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10631), .S(n14129), .Z(
        n10632) );
  NAND2_X1 U13181 ( .A1(n10633), .A2(n10632), .ZN(n14140) );
  NAND2_X1 U13182 ( .A1(n14129), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n14139) );
  NAND2_X1 U13183 ( .A1(n14140), .A2(n14139), .ZN(n10636) );
  INV_X1 U13184 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10634) );
  MUX2_X1 U13185 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10634), .S(n14148), .Z(
        n10635) );
  NAND2_X1 U13186 ( .A1(n10636), .A2(n10635), .ZN(n14158) );
  NAND2_X1 U13187 ( .A1(n14148), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n14157) );
  NAND2_X1 U13188 ( .A1(n14158), .A2(n14157), .ZN(n10639) );
  INV_X1 U13189 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10637) );
  MUX2_X1 U13190 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10637), .S(n14161), .Z(
        n10638) );
  NAND2_X1 U13191 ( .A1(n10639), .A2(n10638), .ZN(n14160) );
  NAND2_X1 U13192 ( .A1(n14161), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10640) );
  NAND2_X1 U13193 ( .A1(n14160), .A2(n10640), .ZN(n10642) );
  OR2_X1 U13194 ( .A1(n10642), .A2(n10643), .ZN(n10800) );
  INV_X1 U13195 ( .A(n10800), .ZN(n10641) );
  AOI21_X1 U13196 ( .B1(n10643), .B2(n10642), .A(n10641), .ZN(n10665) );
  INV_X1 U13197 ( .A(n10644), .ZN(n10645) );
  NAND2_X1 U13198 ( .A1(n10646), .A2(n10645), .ZN(n10844) );
  INV_X1 U13199 ( .A(n10844), .ZN(n10647) );
  INV_X1 U13200 ( .A(n10373), .ZN(n10839) );
  OR2_X1 U13201 ( .A1(n10844), .A2(n10839), .ZN(n14976) );
  AND2_X1 U13202 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n11505) );
  NOR2_X1 U13203 ( .A1(n14980), .A2(n7173), .ZN(n10648) );
  AOI211_X1 U13204 ( .C1(n14206), .C2(n10798), .A(n11505), .B(n10648), .ZN(
        n10664) );
  INV_X1 U13205 ( .A(n14629), .ZN(n10840) );
  NAND2_X1 U13206 ( .A1(n10839), .A2(n10840), .ZN(n10649) );
  INV_X1 U13207 ( .A(n14972), .ZN(n14232) );
  XNOR2_X1 U13208 ( .A(n10650), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n14117) );
  AND2_X1 U13209 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10651) );
  NAND2_X1 U13210 ( .A1(n14117), .A2(n10651), .ZN(n14116) );
  NAND2_X1 U13211 ( .A1(n14113), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10652) );
  NAND2_X1 U13212 ( .A1(n14116), .A2(n10652), .ZN(n14134) );
  MUX2_X1 U13213 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n11437), .S(n14129), .Z(
        n14135) );
  NAND2_X1 U13214 ( .A1(n14134), .A2(n14135), .ZN(n14145) );
  NAND2_X1 U13215 ( .A1(n14129), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14144) );
  NAND2_X1 U13216 ( .A1(n14145), .A2(n14144), .ZN(n10654) );
  INV_X1 U13217 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n14143) );
  MUX2_X1 U13218 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n14143), .S(n14148), .Z(
        n10653) );
  NAND2_X1 U13219 ( .A1(n10654), .A2(n10653), .ZN(n14165) );
  NAND2_X1 U13220 ( .A1(n14148), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n14164) );
  NAND2_X1 U13221 ( .A1(n14165), .A2(n14164), .ZN(n10656) );
  INV_X1 U13222 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n14162) );
  MUX2_X1 U13223 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n14162), .S(n14161), .Z(
        n10655) );
  NAND2_X1 U13224 ( .A1(n10656), .A2(n10655), .ZN(n14167) );
  NAND2_X1 U13225 ( .A1(n14161), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10661) );
  NAND2_X1 U13226 ( .A1(n14167), .A2(n10661), .ZN(n10659) );
  MUX2_X1 U13227 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10657), .S(n10798), .Z(
        n10658) );
  NAND2_X1 U13228 ( .A1(n10659), .A2(n10658), .ZN(n14176) );
  MUX2_X1 U13229 ( .A(n10657), .B(P1_REG2_REG_5__SCAN_IN), .S(n10798), .Z(
        n10660) );
  NAND3_X1 U13230 ( .A1(n14167), .A2(n10661), .A3(n10660), .ZN(n10662) );
  NAND3_X1 U13231 ( .A1(n14232), .A2(n14176), .A3(n10662), .ZN(n10663) );
  OAI211_X1 U13232 ( .C1(n10665), .C2(n14974), .A(n10664), .B(n10663), .ZN(
        P1_U3248) );
  NOR2_X1 U13233 ( .A1(n15136), .A2(n10673), .ZN(n10671) );
  NAND2_X1 U13234 ( .A1(n10669), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10666) );
  NAND2_X1 U13235 ( .A1(n10667), .A2(n10666), .ZN(n10674) );
  NOR3_X1 U13236 ( .A1(n10679), .A2(n12083), .A3(n15129), .ZN(n10670) );
  AOI211_X1 U13237 ( .C1(n10671), .C2(n10674), .A(n15168), .B(n10670), .ZN(
        n10684) );
  AND2_X1 U13238 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n10677) );
  MUX2_X1 U13239 ( .A(n10673), .B(P2_REG1_REG_9__SCAN_IN), .S(n10814), .Z(
        n10672) );
  OR2_X1 U13240 ( .A1(n10674), .A2(n10672), .ZN(n10819) );
  NAND3_X1 U13241 ( .A1(n10674), .A2(n10817), .A3(n10673), .ZN(n10675) );
  AOI21_X1 U13242 ( .B1(n10819), .B2(n10675), .A(n15136), .ZN(n10676) );
  AOI211_X1 U13243 ( .C1(n15196), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n10677), .B(
        n10676), .ZN(n10683) );
  NOR3_X1 U13244 ( .A1(n10679), .A2(n10814), .A3(P2_REG2_REG_9__SCAN_IN), .ZN(
        n10681) );
  MUX2_X1 U13245 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n12083), .S(n10814), .Z(
        n10678) );
  INV_X1 U13246 ( .A(n10813), .ZN(n10680) );
  OAI21_X1 U13247 ( .B1(n10681), .B2(n10680), .A(n15198), .ZN(n10682) );
  OAI211_X1 U13248 ( .C1(n10684), .C2(n10817), .A(n10683), .B(n10682), .ZN(
        P2_U3223) );
  NOR4_X1 U13249 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n10688) );
  NOR4_X1 U13250 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n10687) );
  NOR4_X1 U13251 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n10686) );
  NOR4_X1 U13252 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n10685) );
  AND4_X1 U13253 ( .A1(n10688), .A2(n10687), .A3(n10686), .A4(n10685), .ZN(
        n10693) );
  NOR2_X1 U13254 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .ZN(
        n15721) );
  NOR4_X1 U13255 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n10691) );
  NOR4_X1 U13256 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n10690) );
  NOR4_X1 U13257 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n10689) );
  AND4_X1 U13258 ( .A1(n15721), .A2(n10691), .A3(n10690), .A4(n10689), .ZN(
        n10692) );
  NAND2_X1 U13259 ( .A1(n10693), .A2(n10692), .ZN(n10829) );
  INV_X1 U13260 ( .A(n10829), .ZN(n10694) );
  NOR2_X1 U13261 ( .A1(n10831), .A2(n10694), .ZN(n10695) );
  NOR2_X1 U13262 ( .A1(n11157), .A2(n10695), .ZN(n10697) );
  OAI21_X1 U13263 ( .B1(n10831), .B2(P1_D_REG_0__SCAN_IN), .A(n10832), .ZN(
        n10696) );
  AND2_X1 U13264 ( .A1(n10697), .A2(n10696), .ZN(n11302) );
  OR2_X1 U13265 ( .A1(n10831), .A2(P1_D_REG_1__SCAN_IN), .ZN(n10699) );
  NAND2_X1 U13266 ( .A1(n10551), .A2(n14634), .ZN(n10698) );
  NAND2_X1 U13267 ( .A1(n10699), .A2(n10698), .ZN(n11300) );
  INV_X1 U13268 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15696) );
  INV_X1 U13269 ( .A(n10707), .ZN(n10701) );
  INV_X1 U13270 ( .A(n11463), .ZN(n11134) );
  NAND2_X1 U13271 ( .A1(n11168), .A2(n11134), .ZN(n10702) );
  NAND2_X1 U13272 ( .A1(n10701), .A2(n10702), .ZN(n11107) );
  INV_X1 U13273 ( .A(n10702), .ZN(n10703) );
  NAND2_X1 U13274 ( .A1(n10707), .A2(n10703), .ZN(n10704) );
  NAND2_X1 U13275 ( .A1(n11107), .A2(n10704), .ZN(n14495) );
  INV_X1 U13276 ( .A(n14495), .ZN(n10718) );
  OR2_X1 U13277 ( .A1(n10705), .A2(n14235), .ZN(n15055) );
  NAND2_X1 U13278 ( .A1(n11134), .A2(n14494), .ZN(n10706) );
  NAND2_X1 U13279 ( .A1(n11117), .A2(n10706), .ZN(n10715) );
  INV_X1 U13280 ( .A(n14110), .ZN(n11144) );
  XNOR2_X1 U13281 ( .A(n10715), .B(n11144), .ZN(n10708) );
  MUX2_X1 U13282 ( .A(n10708), .B(n10707), .S(n11168), .Z(n10713) );
  OR2_X1 U13283 ( .A1(n10709), .A2(n11132), .ZN(n10710) );
  NAND2_X1 U13284 ( .A1(n11306), .A2(n14235), .ZN(n15081) );
  INV_X1 U13285 ( .A(n15081), .ZN(n15059) );
  NAND2_X1 U13286 ( .A1(n14495), .A2(n15059), .ZN(n10712) );
  OR2_X1 U13287 ( .A1(n11151), .A2(n10839), .ZN(n14464) );
  AOI22_X1 U13288 ( .A1(n14109), .A2(n14477), .B1(n14479), .B2(n11168), .ZN(
        n10711) );
  OAI211_X1 U13289 ( .C1(n10713), .C2(n15002), .A(n10712), .B(n10711), .ZN(
        n14497) );
  INV_X1 U13290 ( .A(n14497), .ZN(n10717) );
  OR2_X1 U13291 ( .A1(n14640), .A2(n10714), .ZN(n11313) );
  NOR2_X1 U13292 ( .A1(n10715), .A2(n15014), .ZN(n14496) );
  AOI21_X1 U13293 ( .B1(n14494), .B2(n14951), .A(n14496), .ZN(n10716) );
  OAI211_X1 U13294 ( .C1(n10718), .C2(n15055), .A(n10717), .B(n10716), .ZN(
        n10835) );
  NAND2_X1 U13295 ( .A1(n10835), .A2(n15096), .ZN(n10719) );
  OAI21_X1 U13296 ( .B1(n15096), .B2(n15696), .A(n10719), .ZN(P1_U3462) );
  XOR2_X1 U13297 ( .A(n10721), .B(n10720), .Z(n10726) );
  AOI211_X1 U13298 ( .C1(n10724), .C2(n10723), .A(n10722), .B(n15129), .ZN(
        n10725) );
  AOI21_X1 U13299 ( .B1(n15190), .B2(n10726), .A(n10725), .ZN(n10729) );
  OAI22_X1 U13300 ( .A1(n15166), .A2(n7662), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11780), .ZN(n10727) );
  INV_X1 U13301 ( .A(n10727), .ZN(n10728) );
  OAI211_X1 U13302 ( .C1(n10730), .C2(n15204), .A(n10729), .B(n10728), .ZN(
        P2_U3216) );
  NAND2_X1 U13303 ( .A1(n10731), .A2(n10933), .ZN(n10732) );
  NAND2_X1 U13304 ( .A1(n10733), .A2(n10732), .ZN(n10752) );
  OR2_X1 U13305 ( .A1(n10950), .A2(n9407), .ZN(n10751) );
  INV_X1 U13306 ( .A(n10751), .ZN(n10734) );
  MUX2_X1 U13307 ( .A(n10738), .B(P3_U3897), .S(n10735), .Z(n13041) );
  INV_X1 U13308 ( .A(n10736), .ZN(n10737) );
  NOR2_X1 U13309 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n10763), .ZN(n10988) );
  NAND2_X1 U13310 ( .A1(n8680), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10739) );
  AOI22_X1 U13311 ( .A1(P3_REG2_REG_2__SCAN_IN), .A2(n10777), .B1(n6548), .B2(
        n10766), .ZN(n10740) );
  AOI21_X1 U13312 ( .B1(n10741), .B2(n10740), .A(n10887), .ZN(n10755) );
  NOR2_X1 U13313 ( .A1(n10742), .A2(n10764), .ZN(n13049) );
  NOR2_X1 U13314 ( .A1(n10762), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10744) );
  INV_X1 U13315 ( .A(n10744), .ZN(n10743) );
  NOR2_X1 U13316 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10743), .ZN(n10746) );
  NAND2_X1 U13317 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10744), .ZN(n10745) );
  AOI22_X1 U13318 ( .A1(P3_REG1_REG_2__SCAN_IN), .A2(n10777), .B1(n6548), .B2(
        n10765), .ZN(n10747) );
  NOR2_X1 U13319 ( .A1(n10748), .A2(n10747), .ZN(n10894) );
  AOI21_X1 U13320 ( .B1(n10748), .B2(n10747), .A(n10894), .ZN(n10749) );
  INV_X1 U13321 ( .A(n10749), .ZN(n10750) );
  NAND2_X1 U13322 ( .A1(n13049), .A2(n10750), .ZN(n10754) );
  AOI22_X1 U13323 ( .A1(n15280), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10753) );
  OAI211_X1 U13324 ( .C1(n13040), .C2(n10755), .A(n10754), .B(n10753), .ZN(
        n10776) );
  MUX2_X1 U13325 ( .A(n10757), .B(n10756), .S(n12946), .Z(n10759) );
  NAND2_X1 U13326 ( .A1(n10759), .A2(n10758), .ZN(n10773) );
  INV_X1 U13327 ( .A(n10759), .ZN(n10760) );
  NAND2_X1 U13328 ( .A1(n10760), .A2(n6781), .ZN(n10761) );
  NAND2_X1 U13329 ( .A1(n10773), .A2(n10761), .ZN(n10956) );
  MUX2_X1 U13330 ( .A(n10763), .B(n10762), .S(n12946), .Z(n10989) );
  NAND2_X1 U13331 ( .A1(n10989), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10957) );
  INV_X1 U13332 ( .A(n10773), .ZN(n10770) );
  INV_X1 U13333 ( .A(n10767), .ZN(n10768) );
  INV_X1 U13334 ( .A(n10772), .ZN(n10769) );
  INV_X1 U13335 ( .A(n10771), .ZN(n10958) );
  NAND3_X1 U13336 ( .A1(n10958), .A2(n10773), .A3(n10772), .ZN(n10774) );
  NAND2_X1 U13337 ( .A1(P3_U3897), .A2(n12652), .ZN(n13051) );
  AOI21_X1 U13338 ( .B1(n11100), .B2(n10774), .A(n13051), .ZN(n10775) );
  AOI211_X1 U13339 ( .C1(n13041), .C2(n10777), .A(n10776), .B(n10775), .ZN(
        n10778) );
  INV_X1 U13340 ( .A(n10778), .ZN(P3_U3184) );
  AOI222_X1 U13341 ( .A1(n10779), .A2(n14762), .B1(SI_15_), .B2(n14761), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n12977), .ZN(n10780) );
  INV_X1 U13342 ( .A(n10780), .ZN(P3_U3280) );
  INV_X1 U13343 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n14174) );
  MUX2_X1 U13344 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n14174), .S(n14179), .Z(
        n10782) );
  NAND2_X1 U13345 ( .A1(n10798), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n14175) );
  NAND2_X1 U13346 ( .A1(n14176), .A2(n14175), .ZN(n10781) );
  NAND2_X1 U13347 ( .A1(n10782), .A2(n10781), .ZN(n14192) );
  NAND2_X1 U13348 ( .A1(n14179), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n14191) );
  NAND2_X1 U13349 ( .A1(n14192), .A2(n14191), .ZN(n10785) );
  INV_X1 U13350 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10783) );
  MUX2_X1 U13351 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10783), .S(n14194), .Z(
        n10784) );
  NAND2_X1 U13352 ( .A1(n10785), .A2(n10784), .ZN(n14202) );
  NAND2_X1 U13353 ( .A1(n14194), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n14201) );
  NAND2_X1 U13354 ( .A1(n14202), .A2(n14201), .ZN(n10787) );
  INV_X1 U13355 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11733) );
  MUX2_X1 U13356 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n11733), .S(n14205), .Z(
        n10786) );
  NAND2_X1 U13357 ( .A1(n10787), .A2(n10786), .ZN(n14204) );
  NAND2_X1 U13358 ( .A1(n14205), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10792) );
  NAND2_X1 U13359 ( .A1(n14204), .A2(n10792), .ZN(n10789) );
  MUX2_X1 U13360 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10790), .S(n10976), .Z(
        n10788) );
  NAND2_X1 U13361 ( .A1(n10789), .A2(n10788), .ZN(n10981) );
  INV_X1 U13362 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10790) );
  MUX2_X1 U13363 ( .A(n10790), .B(P1_REG2_REG_9__SCAN_IN), .S(n10976), .Z(
        n10791) );
  NAND3_X1 U13364 ( .A1(n14204), .A2(n10792), .A3(n10791), .ZN(n10793) );
  NAND3_X1 U13365 ( .A1(n14232), .A2(n10981), .A3(n10793), .ZN(n10797) );
  NOR2_X1 U13366 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10794), .ZN(n10795) );
  AOI21_X1 U13367 ( .B1(n14212), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n10795), .ZN(
        n10796) );
  OAI211_X1 U13368 ( .C1(n14976), .C2(n10970), .A(n10797), .B(n10796), .ZN(
        n10812) );
  OR2_X1 U13369 ( .A1(n10798), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n10799) );
  AND2_X1 U13370 ( .A1(n10800), .A2(n10799), .ZN(n14173) );
  INV_X1 U13371 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10801) );
  MUX2_X1 U13372 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10801), .S(n14179), .Z(
        n14172) );
  NAND2_X1 U13373 ( .A1(n14173), .A2(n14172), .ZN(n14187) );
  NAND2_X1 U13374 ( .A1(n14179), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n14186) );
  NAND2_X1 U13375 ( .A1(n14187), .A2(n14186), .ZN(n10804) );
  INV_X1 U13376 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10802) );
  MUX2_X1 U13377 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10802), .S(n14194), .Z(
        n10803) );
  NAND2_X1 U13378 ( .A1(n10804), .A2(n10803), .ZN(n14189) );
  NAND2_X1 U13379 ( .A1(n14194), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10805) );
  AND2_X1 U13380 ( .A1(n14189), .A2(n10805), .ZN(n14208) );
  INV_X1 U13381 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n15102) );
  MUX2_X1 U13382 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n15102), .S(n14205), .Z(
        n14209) );
  NAND2_X1 U13383 ( .A1(n14208), .A2(n14209), .ZN(n14207) );
  OR2_X1 U13384 ( .A1(n14205), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10808) );
  NAND2_X1 U13385 ( .A1(n14207), .A2(n10808), .ZN(n10806) );
  MUX2_X1 U13386 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9993), .S(n10976), .Z(
        n10807) );
  NAND2_X1 U13387 ( .A1(n10806), .A2(n10807), .ZN(n10972) );
  INV_X1 U13388 ( .A(n10807), .ZN(n10809) );
  NAND3_X1 U13389 ( .A1(n14207), .A2(n10809), .A3(n10808), .ZN(n10810) );
  AOI21_X1 U13390 ( .B1(n10972), .B2(n10810), .A(n14974), .ZN(n10811) );
  OR2_X1 U13391 ( .A1(n10812), .A2(n10811), .ZN(P1_U3252) );
  MUX2_X1 U13392 ( .A(n12097), .B(P2_REG2_REG_10__SCAN_IN), .S(n11040), .Z(
        n10815) );
  AOI211_X1 U13393 ( .C1(n10816), .C2(n10815), .A(n15129), .B(n11037), .ZN(
        n10827) );
  NAND2_X1 U13394 ( .A1(n10817), .A2(n10673), .ZN(n10818) );
  NAND2_X1 U13395 ( .A1(n10819), .A2(n10818), .ZN(n10822) );
  MUX2_X1 U13396 ( .A(n8277), .B(P2_REG1_REG_10__SCAN_IN), .S(n11040), .Z(
        n10821) );
  OR2_X1 U13397 ( .A1(n10822), .A2(n10821), .ZN(n11047) );
  INV_X1 U13398 ( .A(n11047), .ZN(n10820) );
  AOI211_X1 U13399 ( .C1(n10822), .C2(n10821), .A(n15136), .B(n10820), .ZN(
        n10826) );
  NAND2_X1 U13400 ( .A1(n15196), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n10823) );
  NAND2_X1 U13401 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n11925)
         );
  OAI211_X1 U13402 ( .C1(n15204), .C2(n10824), .A(n10823), .B(n11925), .ZN(
        n10825) );
  OR3_X1 U13403 ( .A1(n10827), .A2(n10826), .A3(n10825), .ZN(P2_U3224) );
  NOR2_X1 U13404 ( .A1(n10829), .A2(n10828), .ZN(n10830) );
  OR2_X1 U13405 ( .A1(n10831), .A2(n10830), .ZN(n10833) );
  NAND2_X1 U13406 ( .A1(n10833), .A2(n10832), .ZN(n11154) );
  NOR2_X1 U13407 ( .A1(n11154), .A2(n11157), .ZN(n10834) );
  NAND2_X1 U13408 ( .A1(n10835), .A2(n15107), .ZN(n10836) );
  OAI21_X1 U13409 ( .B1(n15107), .B2(n10630), .A(n10836), .ZN(P1_U3529) );
  INV_X1 U13410 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10837) );
  NAND2_X1 U13411 ( .A1(n10840), .A2(n10837), .ZN(n10838) );
  NAND2_X1 U13412 ( .A1(n10839), .A2(n10838), .ZN(n14124) );
  INV_X1 U13413 ( .A(n14124), .ZN(n10841) );
  OAI21_X1 U13414 ( .B1(n10840), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10841), .ZN(
        n10842) );
  MUX2_X1 U13415 ( .A(n10842), .B(n10841), .S(P1_IR_REG_0__SCAN_IN), .Z(n10843) );
  INV_X1 U13416 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11457) );
  OAI22_X1 U13417 ( .A1(n10844), .A2(n10843), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11457), .ZN(n10846) );
  NOR3_X1 U13418 ( .A1(n14974), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n14123), .ZN(
        n10845) );
  AOI211_X1 U13419 ( .C1(n14212), .C2(P1_ADDR_REG_0__SCAN_IN), .A(n10846), .B(
        n10845), .ZN(n10847) );
  INV_X1 U13420 ( .A(n10847), .ZN(P1_U3243) );
  MUX2_X1 U13421 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n10579), .S(n10860), .Z(
        n10850) );
  NAND3_X1 U13422 ( .A1(n10850), .A2(n10849), .A3(n10848), .ZN(n10851) );
  NAND3_X1 U13423 ( .A1(n15190), .A2(n10863), .A3(n10851), .ZN(n10859) );
  NAND2_X1 U13424 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n11621) );
  AOI211_X1 U13425 ( .C1(n10854), .C2(n10853), .A(n10852), .B(n15129), .ZN(
        n10855) );
  INV_X1 U13426 ( .A(n10855), .ZN(n10856) );
  NAND2_X1 U13427 ( .A1(n11621), .A2(n10856), .ZN(n10857) );
  AOI21_X1 U13428 ( .B1(n15196), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n10857), .ZN(
        n10858) );
  OAI211_X1 U13429 ( .C1(n15204), .C2(n10860), .A(n10859), .B(n10858), .ZN(
        P2_U3219) );
  MUX2_X1 U13430 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10583), .S(n10874), .Z(
        n10861) );
  NAND3_X1 U13431 ( .A1(n10863), .A2(n10862), .A3(n10861), .ZN(n10864) );
  NAND3_X1 U13432 ( .A1(n15190), .A2(n10865), .A3(n10864), .ZN(n10873) );
  NAND2_X1 U13433 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n11369) );
  AOI211_X1 U13434 ( .C1(n10868), .C2(n10867), .A(n10866), .B(n15129), .ZN(
        n10869) );
  INV_X1 U13435 ( .A(n10869), .ZN(n10870) );
  NAND2_X1 U13436 ( .A1(n11369), .A2(n10870), .ZN(n10871) );
  AOI21_X1 U13437 ( .B1(n15196), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n10871), .ZN(
        n10872) );
  OAI211_X1 U13438 ( .C1(n15204), .C2(n10874), .A(n10873), .B(n10872), .ZN(
        P2_U3220) );
  INV_X1 U13439 ( .A(n13041), .ZN(n12935) );
  INV_X1 U13440 ( .A(n10922), .ZN(n10905) );
  MUX2_X1 U13441 ( .A(n10876), .B(n10875), .S(n12946), .Z(n10877) );
  NAND2_X1 U13442 ( .A1(n10877), .A2(n10888), .ZN(n10880) );
  INV_X1 U13443 ( .A(n10877), .ZN(n10878) );
  NAND2_X1 U13444 ( .A1(n10878), .A2(n14750), .ZN(n10879) );
  NAND2_X1 U13445 ( .A1(n10880), .A2(n10879), .ZN(n11098) );
  INV_X1 U13446 ( .A(n10880), .ZN(n10884) );
  INV_X1 U13447 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10906) );
  MUX2_X1 U13448 ( .A(n10906), .B(n10921), .S(n12946), .Z(n10881) );
  NAND2_X1 U13449 ( .A1(n10881), .A2(n10922), .ZN(n10916) );
  INV_X1 U13450 ( .A(n10881), .ZN(n10882) );
  NAND2_X1 U13451 ( .A1(n10882), .A2(n10905), .ZN(n10883) );
  INV_X1 U13452 ( .A(n10917), .ZN(n10886) );
  NOR3_X1 U13453 ( .A1(n11097), .A2(n10884), .A3(n7950), .ZN(n10885) );
  OAI21_X1 U13454 ( .B1(n10886), .B2(n10885), .A(n12916), .ZN(n10904) );
  INV_X1 U13455 ( .A(n13040), .ZN(n12995) );
  MUX2_X1 U13456 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n10906), .S(n10922), .Z(
        n10891) );
  NOR2_X1 U13457 ( .A1(n10888), .A2(n10889), .ZN(n10890) );
  XNOR2_X1 U13458 ( .A(n10889), .B(n10888), .ZN(n11092) );
  OAI21_X1 U13459 ( .B1(n6773), .B2(n6741), .A(n10908), .ZN(n10902) );
  INV_X1 U13460 ( .A(n15280), .ZN(n13012) );
  INV_X1 U13461 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10892) );
  NOR2_X1 U13462 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10892), .ZN(n11577) );
  INV_X1 U13463 ( .A(n11577), .ZN(n10893) );
  OAI21_X1 U13464 ( .B1(n13012), .B2(n7174), .A(n10893), .ZN(n10901) );
  NOR2_X1 U13465 ( .A1(n10888), .A2(n10895), .ZN(n10896) );
  MUX2_X1 U13466 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n10921), .S(n10922), .Z(
        n10897) );
  NAND2_X1 U13467 ( .A1(n10898), .A2(n10897), .ZN(n10899) );
  AOI21_X1 U13468 ( .B1(n10924), .B2(n10899), .A(n13004), .ZN(n10900) );
  AOI211_X1 U13469 ( .C1(n12995), .C2(n10902), .A(n10901), .B(n10900), .ZN(
        n10903) );
  OAI211_X1 U13470 ( .C1(n12935), .C2(n10905), .A(n10904), .B(n10903), .ZN(
        P3_U3186) );
  OR2_X1 U13471 ( .A1(n10922), .A2(n10906), .ZN(n10907) );
  AOI21_X1 U13472 ( .B1(n10911), .B2(n10909), .A(n11058), .ZN(n10932) );
  MUX2_X1 U13473 ( .A(n10911), .B(n10910), .S(n12946), .Z(n10912) );
  NAND2_X1 U13474 ( .A1(n10912), .A2(n7480), .ZN(n11062) );
  INV_X1 U13475 ( .A(n10912), .ZN(n10913) );
  NAND2_X1 U13476 ( .A1(n10913), .A2(n10925), .ZN(n10914) );
  NAND2_X1 U13477 ( .A1(n11062), .A2(n10914), .ZN(n10915) );
  AND3_X1 U13478 ( .A1(n10917), .A2(n10916), .A3(n10915), .ZN(n10918) );
  OAI21_X1 U13479 ( .B1(n11067), .B2(n10918), .A(n12916), .ZN(n10931) );
  INV_X1 U13480 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n10920) );
  AND2_X1 U13481 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n11743) );
  INV_X1 U13482 ( .A(n11743), .ZN(n10919) );
  OAI21_X1 U13483 ( .B1(n13012), .B2(n10920), .A(n10919), .ZN(n10929) );
  OR2_X1 U13484 ( .A1(n10922), .A2(n10921), .ZN(n10923) );
  AOI21_X1 U13485 ( .B1(n10910), .B2(n10926), .A(n11072), .ZN(n10927) );
  NOR2_X1 U13486 ( .A1(n10927), .A2(n13004), .ZN(n10928) );
  AOI211_X1 U13487 ( .C1(n13041), .C2(n7480), .A(n10929), .B(n10928), .ZN(
        n10930) );
  OAI211_X1 U13488 ( .C1(n10932), .C2(n13040), .A(n10931), .B(n10930), .ZN(
        P3_U3187) );
  INV_X1 U13489 ( .A(n10944), .ZN(n10936) );
  NAND3_X1 U13490 ( .A1(n11356), .A2(n10934), .A3(n10933), .ZN(n10935) );
  AOI21_X1 U13491 ( .B1(n10947), .B2(n10936), .A(n10935), .ZN(n10939) );
  NAND2_X1 U13492 ( .A1(n10949), .A2(n10937), .ZN(n10938) );
  NAND2_X1 U13493 ( .A1(n10939), .A2(n10938), .ZN(n10940) );
  NAND2_X1 U13494 ( .A1(n10940), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10943) );
  NAND2_X1 U13495 ( .A1(n10947), .A2(n10941), .ZN(n10942) );
  NOR2_X1 U13496 ( .A1(n15439), .A2(P3_U3151), .ZN(n11397) );
  INV_X1 U13497 ( .A(n11127), .ZN(n10954) );
  INV_X1 U13498 ( .A(n11125), .ZN(n10945) );
  OAI22_X1 U13499 ( .A1(n10949), .A2(n10945), .B1(n10947), .B2(n10944), .ZN(
        n10946) );
  NAND2_X1 U13500 ( .A1(n10946), .A2(n10950), .ZN(n15434) );
  NOR2_X1 U13501 ( .A1(n15300), .A2(n11281), .ZN(n10948) );
  INV_X1 U13502 ( .A(n10947), .ZN(n11283) );
  NAND2_X1 U13503 ( .A1(n10949), .A2(n15368), .ZN(n10952) );
  NAND2_X1 U13504 ( .A1(n10950), .A2(n13290), .ZN(n11361) );
  INV_X1 U13505 ( .A(n11361), .ZN(n10951) );
  OAI22_X1 U13506 ( .A1(n11285), .A2(n12891), .B1(n12882), .B2(n11432), .ZN(
        n10953) );
  AOI21_X1 U13507 ( .B1(n10954), .B2(n12861), .A(n10953), .ZN(n10955) );
  OAI21_X1 U13508 ( .B1(n11397), .B2(n15714), .A(n10955), .ZN(P3_U3172) );
  INV_X1 U13509 ( .A(n10956), .ZN(n10959) );
  INV_X1 U13510 ( .A(n10957), .ZN(n10996) );
  OAI21_X1 U13511 ( .B1(n10959), .B2(n10996), .A(n10958), .ZN(n10968) );
  XNOR2_X1 U13512 ( .A(n10960), .B(P3_REG2_REG_1__SCAN_IN), .ZN(n10966) );
  NOR2_X1 U13513 ( .A1(n10961), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10962) );
  OAI21_X1 U13514 ( .B1(n10963), .B2(n10962), .A(n13049), .ZN(n10965) );
  AOI22_X1 U13515 ( .A1(n15280), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10964) );
  OAI211_X1 U13516 ( .C1(n13040), .C2(n10966), .A(n10965), .B(n10964), .ZN(
        n10967) );
  AOI21_X1 U13517 ( .B1(n12916), .B2(n10968), .A(n10967), .ZN(n10969) );
  OAI21_X1 U13518 ( .B1(n6781), .B2(n12935), .A(n10969), .ZN(P3_U3183) );
  NAND2_X1 U13519 ( .A1(n10970), .A2(n9993), .ZN(n10971) );
  NAND2_X1 U13520 ( .A1(n10972), .A2(n10971), .ZN(n10975) );
  INV_X1 U13521 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n15536) );
  MUX2_X1 U13522 ( .A(n15536), .B(P1_REG1_REG_10__SCAN_IN), .S(n11002), .Z(
        n10974) );
  OR2_X1 U13523 ( .A1(n10975), .A2(n10974), .ZN(n11004) );
  INV_X1 U13524 ( .A(n11004), .ZN(n10973) );
  AOI211_X1 U13525 ( .C1(n10975), .C2(n10974), .A(n14974), .B(n10973), .ZN(
        n10987) );
  NAND2_X1 U13526 ( .A1(n10976), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10980) );
  NAND2_X1 U13527 ( .A1(n10981), .A2(n10980), .ZN(n10978) );
  INV_X1 U13528 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11890) );
  MUX2_X1 U13529 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n11890), .S(n11002), .Z(
        n10977) );
  NAND2_X1 U13530 ( .A1(n10978), .A2(n10977), .ZN(n11001) );
  MUX2_X1 U13531 ( .A(n11890), .B(P1_REG2_REG_10__SCAN_IN), .S(n11002), .Z(
        n10979) );
  NAND3_X1 U13532 ( .A1(n10981), .A2(n10980), .A3(n10979), .ZN(n10982) );
  NAND3_X1 U13533 ( .A1(n14232), .A2(n11001), .A3(n10982), .ZN(n10984) );
  AND2_X1 U13534 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n14871) );
  AOI21_X1 U13535 ( .B1(n14212), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n14871), 
        .ZN(n10983) );
  OAI211_X1 U13536 ( .C1(n14976), .C2(n10985), .A(n10984), .B(n10983), .ZN(
        n10986) );
  OR2_X1 U13537 ( .A1(n10987), .A2(n10986), .ZN(P1_U3253) );
  NAND3_X1 U13538 ( .A1(n13004), .A2(n13051), .A3(n13040), .ZN(n10995) );
  AOI22_X1 U13539 ( .A1(n12995), .A2(n10988), .B1(n13049), .B2(n10744), .ZN(
        n10993) );
  NOR2_X1 U13540 ( .A1(n13051), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10991) );
  INV_X1 U13541 ( .A(n10989), .ZN(n10990) );
  AOI22_X1 U13542 ( .A1(n10991), .A2(n10990), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10992) );
  OAI211_X1 U13543 ( .C1(n14685), .C2(n13012), .A(n10993), .B(n10992), .ZN(
        n10994) );
  AOI21_X1 U13544 ( .B1(n10996), .B2(n10995), .A(n10994), .ZN(n10997) );
  OAI21_X1 U13545 ( .B1(n10998), .B2(n12935), .A(n10997), .ZN(P3_U3182) );
  INV_X1 U13546 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n15643) );
  NAND2_X1 U13547 ( .A1(n13187), .A2(P3_U3897), .ZN(n10999) );
  OAI21_X1 U13548 ( .B1(P3_U3897), .B2(n15643), .A(n10999), .ZN(P3_U3511) );
  NAND2_X1 U13549 ( .A1(n11002), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n11000) );
  AND2_X1 U13550 ( .A1(n11001), .A2(n11000), .ZN(n11008) );
  NOR2_X1 U13551 ( .A1(n14972), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11006) );
  NAND2_X1 U13552 ( .A1(n11002), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n11003) );
  AND2_X1 U13553 ( .A1(n11004), .A2(n11003), .ZN(n11015) );
  INV_X1 U13554 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n14908) );
  NOR3_X1 U13555 ( .A1(n11015), .A2(n14974), .A3(n14908), .ZN(n11005) );
  AOI211_X1 U13556 ( .C1(n11008), .C2(n11006), .A(n14206), .B(n11005), .ZN(
        n11019) );
  INV_X1 U13557 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n11012) );
  INV_X1 U13558 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11009) );
  MUX2_X1 U13559 ( .A(n11009), .B(P1_REG2_REG_11__SCAN_IN), .S(n11024), .Z(
        n11007) );
  OAI21_X1 U13560 ( .B1(n11024), .B2(n11009), .A(n11008), .ZN(n11010) );
  NAND3_X1 U13561 ( .A1(n11025), .A2(n14232), .A3(n11010), .ZN(n11011) );
  NAND2_X1 U13562 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n12323)
         );
  OAI211_X1 U13563 ( .C1(n11012), .C2(n14980), .A(n11011), .B(n12323), .ZN(
        n11013) );
  INV_X1 U13564 ( .A(n11013), .ZN(n11018) );
  NOR3_X1 U13565 ( .A1(n11015), .A2(n11024), .A3(P1_REG1_REG_11__SCAN_IN), 
        .ZN(n11016) );
  MUX2_X1 U13566 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n14908), .S(n11024), .Z(
        n11014) );
  OAI21_X1 U13567 ( .B1(n11016), .B2(n11020), .A(n14233), .ZN(n11017) );
  OAI211_X1 U13568 ( .C1(n11019), .C2(n11021), .A(n11018), .B(n11017), .ZN(
        P1_U3254) );
  AOI21_X1 U13569 ( .B1(n14908), .B2(n11021), .A(n11020), .ZN(n11023) );
  INV_X1 U13570 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n14787) );
  AOI22_X1 U13571 ( .A1(n11246), .A2(n14787), .B1(P1_REG1_REG_12__SCAN_IN), 
        .B2(n11033), .ZN(n11022) );
  NOR2_X1 U13572 ( .A1(n11023), .A2(n11022), .ZN(n11248) );
  AOI21_X1 U13573 ( .B1(n11023), .B2(n11022), .A(n11248), .ZN(n11036) );
  AOI22_X1 U13574 ( .A1(n11246), .A2(n10036), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n11033), .ZN(n11028) );
  NAND2_X1 U13575 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n11024), .ZN(n11026) );
  NAND2_X1 U13576 ( .A1(n11026), .A2(n11025), .ZN(n11027) );
  NOR2_X1 U13577 ( .A1(n11028), .A2(n11027), .ZN(n11241) );
  AOI21_X1 U13578 ( .B1(n11028), .B2(n11027), .A(n11241), .ZN(n11029) );
  OR2_X1 U13579 ( .A1(n11029), .A2(n14972), .ZN(n11032) );
  NOR2_X1 U13580 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10037), .ZN(n11030) );
  AOI21_X1 U13581 ( .B1(n14212), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n11030), 
        .ZN(n11031) );
  OAI211_X1 U13582 ( .C1(n14976), .C2(n11033), .A(n11032), .B(n11031), .ZN(
        n11034) );
  INV_X1 U13583 ( .A(n11034), .ZN(n11035) );
  OAI21_X1 U13584 ( .B1(n11036), .B2(n14974), .A(n11035), .ZN(P1_U3255) );
  AOI21_X1 U13585 ( .B1(n11040), .B2(P2_REG2_REG_10__SCAN_IN), .A(n11037), 
        .ZN(n11039) );
  MUX2_X1 U13586 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n13549), .S(n11044), .Z(
        n11038) );
  NAND2_X1 U13587 ( .A1(n11039), .A2(n11038), .ZN(n15128) );
  OAI21_X1 U13588 ( .B1(n11039), .B2(n11038), .A(n15128), .ZN(n11053) );
  NAND2_X1 U13589 ( .A1(n11040), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n11046) );
  NAND2_X1 U13590 ( .A1(n11047), .A2(n11046), .ZN(n11043) );
  MUX2_X1 U13591 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n11041), .S(n11044), .Z(
        n11042) );
  NAND2_X1 U13592 ( .A1(n11043), .A2(n11042), .ZN(n13562) );
  MUX2_X1 U13593 ( .A(n11041), .B(P2_REG1_REG_11__SCAN_IN), .S(n11044), .Z(
        n11045) );
  NAND3_X1 U13594 ( .A1(n11047), .A2(n11046), .A3(n11045), .ZN(n11048) );
  NAND3_X1 U13595 ( .A1(n15190), .A2(n13562), .A3(n11048), .ZN(n11051) );
  NAND2_X1 U13596 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n11797)
         );
  INV_X1 U13597 ( .A(n11797), .ZN(n11049) );
  AOI21_X1 U13598 ( .B1(n15196), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n11049), 
        .ZN(n11050) );
  OAI211_X1 U13599 ( .C1(n15204), .C2(n13563), .A(n11051), .B(n11050), .ZN(
        n11052) );
  AOI21_X1 U13600 ( .B1(n11053), .B2(n15198), .A(n11052), .ZN(n11054) );
  INV_X1 U13601 ( .A(n11054), .ZN(P2_U3225) );
  AOI222_X1 U13602 ( .A1(n11055), .A2(n14762), .B1(n12976), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_16_), .C2(n14761), .ZN(n11056) );
  INV_X1 U13603 ( .A(n11056), .ZN(P3_U3279) );
  NOR2_X1 U13604 ( .A1(n7480), .A2(n11057), .ZN(n11059) );
  AOI22_X1 U13605 ( .A1(n11210), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n11202), 
        .B2(n14747), .ZN(n11060) );
  NOR2_X1 U13606 ( .A1(n11061), .A2(n11060), .ZN(n11204) );
  AOI21_X1 U13607 ( .B1(n11061), .B2(n11060), .A(n11204), .ZN(n11080) );
  INV_X1 U13608 ( .A(n11062), .ZN(n11066) );
  INV_X1 U13609 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11202) );
  MUX2_X1 U13610 ( .A(n11202), .B(n11209), .S(n12946), .Z(n11063) );
  NAND2_X1 U13611 ( .A1(n11063), .A2(n11210), .ZN(n11225) );
  INV_X1 U13612 ( .A(n11063), .ZN(n11064) );
  NAND2_X1 U13613 ( .A1(n11064), .A2(n14747), .ZN(n11065) );
  INV_X1 U13614 ( .A(n11226), .ZN(n11069) );
  NOR3_X1 U13615 ( .A1(n11067), .A2(n11066), .A3(n7942), .ZN(n11068) );
  OAI21_X1 U13616 ( .B1(n11069), .B2(n11068), .A(n12916), .ZN(n11079) );
  INV_X1 U13617 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n11071) );
  INV_X1 U13618 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n11070) );
  OR2_X1 U13619 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11070), .ZN(n11985) );
  OAI21_X1 U13620 ( .B1(n13012), .B2(n11071), .A(n11985), .ZN(n11077) );
  AOI22_X1 U13621 ( .A1(n11210), .A2(P3_REG1_REG_6__SCAN_IN), .B1(n11209), 
        .B2(n14747), .ZN(n11073) );
  AOI21_X1 U13622 ( .B1(n11074), .B2(n11073), .A(n6740), .ZN(n11075) );
  NOR2_X1 U13623 ( .A1(n11075), .A2(n13004), .ZN(n11076) );
  AOI211_X1 U13624 ( .C1(n13041), .C2(n11210), .A(n11077), .B(n11076), .ZN(
        n11078) );
  OAI211_X1 U13625 ( .C1(n11080), .C2(n13040), .A(n11079), .B(n11078), .ZN(
        P3_U3188) );
  INV_X1 U13626 ( .A(n15107), .ZN(n15105) );
  INV_X1 U13627 ( .A(n11081), .ZN(n11460) );
  NAND2_X1 U13628 ( .A1(n14599), .A2(n15002), .ZN(n11085) );
  NAND2_X1 U13629 ( .A1(n14110), .A2(n14477), .ZN(n11458) );
  NAND3_X1 U13630 ( .A1(n11134), .A2(n12021), .A3(n11082), .ZN(n11083) );
  NAND2_X1 U13631 ( .A1(n11458), .A2(n11083), .ZN(n11084) );
  AOI21_X1 U13632 ( .B1(n11460), .B2(n11085), .A(n11084), .ZN(n15025) );
  NAND2_X1 U13633 ( .A1(n15105), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n11086) );
  OAI21_X1 U13634 ( .B1(n15105), .B2(n15025), .A(n11086), .ZN(P1_U3528) );
  INV_X1 U13635 ( .A(n13552), .ZN(n15164) );
  OAI222_X1 U13636 ( .A1(n13964), .A2(n15544), .B1(n12649), .B2(n11087), .C1(
        n15164), .C2(P2_U3088), .ZN(P2_U3313) );
  INV_X1 U13637 ( .A(n11264), .ZN(n11964) );
  OAI222_X1 U13638 ( .A1(n14635), .A2(n11088), .B1(n14638), .B2(n11087), .C1(
        n11964), .C2(P1_U3086), .ZN(P1_U3341) );
  AOI21_X1 U13639 ( .B1(n10875), .B2(n11090), .A(n11089), .ZN(n11096) );
  INV_X1 U13640 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n15440) );
  NOR2_X1 U13641 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15440), .ZN(n15426) );
  AOI21_X1 U13642 ( .B1(n10876), .B2(n11092), .A(n11091), .ZN(n11093) );
  NOR2_X1 U13643 ( .A1(n13040), .A2(n11093), .ZN(n11094) );
  AOI211_X1 U13644 ( .C1(n15280), .C2(P3_ADDR_REG_3__SCAN_IN), .A(n15426), .B(
        n11094), .ZN(n11095) );
  OAI21_X1 U13645 ( .B1(n11096), .B2(n13004), .A(n11095), .ZN(n11104) );
  INV_X1 U13646 ( .A(n11097), .ZN(n11102) );
  NAND3_X1 U13647 ( .A1(n11100), .A2(n11099), .A3(n11098), .ZN(n11101) );
  AOI21_X1 U13648 ( .B1(n11102), .B2(n11101), .A(n13051), .ZN(n11103) );
  AOI211_X1 U13649 ( .C1(n13041), .C2(n10888), .A(n11104), .B(n11103), .ZN(
        n11105) );
  INV_X1 U13650 ( .A(n11105), .ZN(P3_U3185) );
  INV_X1 U13651 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n11122) );
  NAND2_X1 U13652 ( .A1(n11107), .A2(n11106), .ZN(n11109) );
  NAND2_X1 U13653 ( .A1(n11109), .A2(n11108), .ZN(n11309) );
  OAI21_X1 U13654 ( .B1(n11109), .B2(n11108), .A(n11309), .ZN(n11110) );
  INV_X1 U13655 ( .A(n11110), .ZN(n11443) );
  AOI21_X2 U13656 ( .B1(n11112), .B2(n11111), .A(n7939), .ZN(n11113) );
  OAI22_X1 U13657 ( .A1(n11144), .A2(n14462), .B1(n11479), .B2(n14464), .ZN(
        n11115) );
  NOR2_X1 U13658 ( .A1(n11443), .A2(n15081), .ZN(n11114) );
  AOI211_X1 U13659 ( .C1(n15052), .C2(n11116), .A(n11115), .B(n11114), .ZN(
        n11436) );
  NAND2_X1 U13660 ( .A1(n11440), .A2(n11117), .ZN(n11118) );
  NAND3_X1 U13661 ( .A1(n11331), .A2(n11131), .A3(n11118), .ZN(n11438) );
  INV_X1 U13662 ( .A(n11438), .ZN(n11119) );
  AOI21_X1 U13663 ( .B1(n11440), .B2(n14951), .A(n11119), .ZN(n11120) );
  OAI211_X1 U13664 ( .C1(n11443), .C2(n15055), .A(n11436), .B(n11120), .ZN(
        n11123) );
  NAND2_X1 U13665 ( .A1(n11123), .A2(n15096), .ZN(n11121) );
  OAI21_X1 U13666 ( .B1(n15096), .B2(n11122), .A(n11121), .ZN(P1_U3465) );
  NAND2_X1 U13667 ( .A1(n11123), .A2(n15107), .ZN(n11124) );
  OAI21_X1 U13668 ( .B1(n15107), .B2(n10631), .A(n11124), .ZN(P1_U3530) );
  NOR2_X1 U13669 ( .A1(n10380), .A2(n11125), .ZN(n11126) );
  OAI22_X1 U13670 ( .A1(n11127), .A2(n11126), .B1(n11285), .B2(n15300), .ZN(
        n11434) );
  INV_X1 U13671 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11128) );
  OAI22_X1 U13672 ( .A1(n11432), .A2(n13376), .B1(n15407), .B2(n11128), .ZN(
        n11129) );
  AOI21_X1 U13673 ( .B1(n11434), .B2(n15407), .A(n11129), .ZN(n11130) );
  INV_X1 U13674 ( .A(n11130), .ZN(P3_U3390) );
  NAND2_X1 U13675 ( .A1(n11131), .A2(n14235), .ZN(n14399) );
  NAND2_X2 U13676 ( .A1(n11133), .A2(n11132), .ZN(n11135) );
  INV_X1 U13677 ( .A(n11133), .ZN(n11137) );
  INV_X1 U13678 ( .A(n11168), .ZN(n11136) );
  NAND2_X1 U13679 ( .A1(n11137), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n11138) );
  OAI211_X1 U13680 ( .C1(n11135), .C2(n11463), .A(n11139), .B(n11138), .ZN(
        n11176) );
  INV_X1 U13681 ( .A(n11176), .ZN(n11140) );
  NAND2_X1 U13682 ( .A1(n11140), .A2(n12777), .ZN(n11141) );
  NAND2_X1 U13683 ( .A1(n11175), .A2(n11141), .ZN(n11166) );
  XNOR2_X1 U13684 ( .A(n11142), .B(n12746), .ZN(n11147) );
  OAI22_X1 U13685 ( .A1(n12776), .A2(n11144), .B1(n11143), .B2(n12779), .ZN(
        n11145) );
  XNOR2_X1 U13686 ( .A(n11145), .B(n11147), .ZN(n11167) );
  NAND2_X1 U13687 ( .A1(n11166), .A2(n11167), .ZN(n11149) );
  INV_X1 U13688 ( .A(n11145), .ZN(n11146) );
  NAND2_X1 U13689 ( .A1(n11147), .A2(n11146), .ZN(n11148) );
  OAI22_X1 U13690 ( .A1(n7324), .A2(n11135), .B1(n12779), .B2(n11338), .ZN(
        n11150) );
  XNOR2_X1 U13691 ( .A(n11150), .B(n12746), .ZN(n11474) );
  OAI22_X1 U13692 ( .A1(n12776), .A2(n11338), .B1(n7324), .B2(n12779), .ZN(
        n11472) );
  XNOR2_X1 U13693 ( .A(n11474), .B(n11472), .ZN(n11470) );
  XNOR2_X1 U13694 ( .A(n11471), .B(n11470), .ZN(n11164) );
  NAND3_X1 U13695 ( .A1(n11305), .A2(n14902), .A3(n11151), .ZN(n11152) );
  NOR2_X1 U13696 ( .A1(n11300), .A2(n11152), .ZN(n11153) );
  INV_X1 U13697 ( .A(n11154), .ZN(n11158) );
  AND2_X1 U13698 ( .A1(n11154), .A2(n11303), .ZN(n11155) );
  NOR2_X1 U13699 ( .A1(n11501), .A2(n11157), .ZN(n11178) );
  NOR2_X1 U13700 ( .A1(n11300), .A2(n11157), .ZN(n11159) );
  AND2_X1 U13701 ( .A1(n11159), .A2(n11158), .ZN(n14960) );
  INV_X1 U13702 ( .A(n14960), .ZN(n14862) );
  OR2_X1 U13703 ( .A1(n14862), .A2(n14464), .ZN(n14085) );
  INV_X1 U13704 ( .A(n14085), .ZN(n14054) );
  AOI22_X1 U13705 ( .A1(n14054), .A2(n14108), .B1(n14087), .B2(n14110), .ZN(
        n11162) );
  NOR2_X1 U13706 ( .A1(n11501), .A2(n11160), .ZN(n14953) );
  AND2_X1 U13707 ( .A1(n14953), .A2(n14951), .ZN(n14090) );
  NAND2_X1 U13708 ( .A1(n14090), .A2(n11440), .ZN(n11161) );
  OAI211_X1 U13709 ( .C1(n11178), .C2(n14127), .A(n11162), .B(n11161), .ZN(
        n11163) );
  AOI21_X1 U13710 ( .B1(n11164), .B2(n14961), .A(n11163), .ZN(n11165) );
  INV_X1 U13711 ( .A(n11165), .ZN(P1_U3237) );
  XOR2_X1 U13712 ( .A(n11167), .B(n11166), .Z(n11172) );
  INV_X1 U13713 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n14111) );
  AOI22_X1 U13714 ( .A1(n14054), .A2(n14109), .B1(n14087), .B2(n11168), .ZN(
        n11169) );
  OAI21_X1 U13715 ( .B1(n11178), .B2(n14111), .A(n11169), .ZN(n11170) );
  AOI21_X1 U13716 ( .B1(n14090), .B2(n14494), .A(n11170), .ZN(n11171) );
  OAI21_X1 U13717 ( .B1(n14935), .B2(n11172), .A(n11171), .ZN(P1_U3222) );
  AOI222_X1 U13718 ( .A1(n11173), .A2(n14762), .B1(SI_17_), .B2(n14761), .C1(
        n13003), .C2(P3_STATE_REG_SCAN_IN), .ZN(n11174) );
  INV_X1 U13719 ( .A(n11174), .ZN(P3_U3278) );
  OAI21_X1 U13720 ( .B1(n11177), .B2(n11176), .A(n11175), .ZN(n14121) );
  OAI22_X1 U13721 ( .A1(n11178), .A2(n11457), .B1(n14862), .B2(n11458), .ZN(
        n11179) );
  AOI21_X1 U13722 ( .B1(n14961), .B2(n14121), .A(n11179), .ZN(n11180) );
  OAI21_X1 U13723 ( .B1(n11463), .B2(n14864), .A(n11180), .ZN(P1_U3232) );
  INV_X1 U13724 ( .A(n11181), .ZN(n11182) );
  OAI222_X1 U13725 ( .A1(n14635), .A2(n15512), .B1(n14638), .B2(n11182), .C1(
        n12151), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U13726 ( .A(n13547), .ZN(n15188) );
  OAI222_X1 U13727 ( .A1(n13964), .A2(n11183), .B1(n12649), .B2(n11182), .C1(
        n15188), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U13728 ( .A(n13030), .ZN(n11186) );
  OAI222_X1 U13729 ( .A1(P3_U3151), .A2(n11186), .B1(n14741), .B2(n11185), 
        .C1(n14743), .C2(n11184), .ZN(P3_U3277) );
  XNOR2_X1 U13730 ( .A(n11188), .B(n11187), .ZN(n12047) );
  OAI21_X1 U13731 ( .B1(n11191), .B2(n11190), .A(n11189), .ZN(n11192) );
  AOI222_X1 U13732 ( .A1(n13819), .A2(n11192), .B1(n13523), .B2(n13816), .C1(
        n13525), .C2(n13814), .ZN(n12048) );
  OAI21_X1 U13733 ( .B1(n11778), .B2(n11194), .A(n13690), .ZN(n11193) );
  OR2_X1 U13734 ( .A1(n11767), .A2(n11193), .ZN(n12045) );
  OAI211_X1 U13735 ( .C1(n11194), .C2(n15263), .A(n12048), .B(n12045), .ZN(
        n11195) );
  AOI21_X1 U13736 ( .B1(n9794), .B2(n12047), .A(n11195), .ZN(n11201) );
  OR2_X1 U13737 ( .A1(n15279), .A2(n10428), .ZN(n11198) );
  OAI21_X1 U13738 ( .B1(n11201), .B2(n15277), .A(n11198), .ZN(P2_U3502) );
  INV_X1 U13739 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n11199) );
  OR2_X1 U13740 ( .A1(n15270), .A2(n11199), .ZN(n11200) );
  OAI21_X1 U13741 ( .B1(n11201), .B2(n9800), .A(n11200), .ZN(P2_U3439) );
  NOR2_X1 U13742 ( .A1(n11210), .A2(n11202), .ZN(n11203) );
  AOI21_X1 U13743 ( .B1(n11206), .B2(n11218), .A(n11551), .ZN(n11230) );
  INV_X1 U13744 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n11208) );
  AND2_X1 U13745 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n12109) );
  INV_X1 U13746 ( .A(n12109), .ZN(n11207) );
  OAI21_X1 U13747 ( .B1(n13012), .B2(n11208), .A(n11207), .ZN(n11216) );
  NOR2_X1 U13748 ( .A1(n11210), .A2(n11209), .ZN(n11211) );
  AOI21_X1 U13749 ( .B1(n11213), .B2(n11217), .A(n11558), .ZN(n11214) );
  NOR2_X1 U13750 ( .A1(n11214), .A2(n13004), .ZN(n11215) );
  AOI211_X1 U13751 ( .C1(n13041), .C2(n11219), .A(n11216), .B(n11215), .ZN(
        n11229) );
  MUX2_X1 U13752 ( .A(n11218), .B(n11217), .S(n12946), .Z(n11220) );
  NAND2_X1 U13753 ( .A1(n11220), .A2(n11219), .ZN(n11545) );
  INV_X1 U13754 ( .A(n11220), .ZN(n11222) );
  NAND2_X1 U13755 ( .A1(n11222), .A2(n11221), .ZN(n11223) );
  NAND2_X1 U13756 ( .A1(n11545), .A2(n11223), .ZN(n11224) );
  AND3_X1 U13757 ( .A1(n11226), .A2(n11225), .A3(n11224), .ZN(n11227) );
  OAI21_X1 U13758 ( .B1(n11547), .B2(n11227), .A(n12916), .ZN(n11228) );
  OAI211_X1 U13759 ( .C1(n11230), .C2(n13040), .A(n11229), .B(n11228), .ZN(
        P3_U3189) );
  OAI222_X1 U13760 ( .A1(n14743), .A2(n11232), .B1(n14741), .B2(n11231), .C1(
        P3_U3151), .C2(n13033), .ZN(P3_U3276) );
  INV_X1 U13761 ( .A(n11233), .ZN(n11235) );
  OAI222_X1 U13762 ( .A1(n14635), .A2(n11234), .B1(n14638), .B2(n11235), .C1(
        n12163), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U13763 ( .A(n13545), .ZN(n15203) );
  OAI222_X1 U13764 ( .A1(n13964), .A2(n11236), .B1(n12649), .B2(n11235), .C1(
        n15203), .C2(P2_U3088), .ZN(P2_U3310) );
  INV_X1 U13765 ( .A(n11237), .ZN(n11239) );
  INV_X1 U13766 ( .A(n15169), .ZN(n13568) );
  OAI222_X1 U13767 ( .A1(n13964), .A2(n11238), .B1(n12649), .B2(n11239), .C1(
        P2_U3088), .C2(n13568), .ZN(P2_U3312) );
  INV_X1 U13768 ( .A(n11965), .ZN(n14975) );
  OAI222_X1 U13769 ( .A1(n14635), .A2(n11240), .B1(n14638), .B2(n11239), .C1(
        P1_U3086), .C2(n14975), .ZN(P1_U3340) );
  NOR2_X1 U13770 ( .A1(n11246), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11242) );
  NOR2_X1 U13771 ( .A1(n11242), .A2(n11241), .ZN(n11245) );
  MUX2_X1 U13772 ( .A(n12173), .B(P1_REG2_REG_13__SCAN_IN), .S(n11261), .Z(
        n11243) );
  INV_X1 U13773 ( .A(n11243), .ZN(n11244) );
  NAND2_X1 U13774 ( .A1(n11244), .A2(n11245), .ZN(n11262) );
  OAI211_X1 U13775 ( .C1(n11245), .C2(n11244), .A(n14232), .B(n11262), .ZN(
        n11254) );
  NAND2_X1 U13776 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n12496)
         );
  NOR2_X1 U13777 ( .A1(n11246), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11247) );
  NOR2_X1 U13778 ( .A1(n11248), .A2(n11247), .ZN(n11250) );
  XNOR2_X1 U13779 ( .A(n11261), .B(n11257), .ZN(n11249) );
  NAND2_X1 U13780 ( .A1(n11250), .A2(n11249), .ZN(n11255) );
  OAI211_X1 U13781 ( .C1(n11250), .C2(n11249), .A(n14233), .B(n11255), .ZN(
        n11251) );
  NAND2_X1 U13782 ( .A1(n12496), .A2(n11251), .ZN(n11252) );
  AOI21_X1 U13783 ( .B1(n14212), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n11252), 
        .ZN(n11253) );
  OAI211_X1 U13784 ( .C1(n14976), .C2(n11256), .A(n11254), .B(n11253), .ZN(
        P1_U3256) );
  AOI22_X1 U13785 ( .A1(n11264), .A2(n15528), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n11964), .ZN(n11259) );
  OAI21_X1 U13786 ( .B1(n11257), .B2(n11256), .A(n11255), .ZN(n11258) );
  NOR2_X1 U13787 ( .A1(n11259), .A2(n11258), .ZN(n11957) );
  AOI21_X1 U13788 ( .B1(n11259), .B2(n11258), .A(n11957), .ZN(n11270) );
  INV_X1 U13789 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14667) );
  NAND2_X1 U13790 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14867)
         );
  OAI21_X1 U13791 ( .B1(n14980), .B2(n14667), .A(n14867), .ZN(n11260) );
  AOI21_X1 U13792 ( .B1(n11264), .B2(n14206), .A(n11260), .ZN(n11269) );
  NAND2_X1 U13793 ( .A1(n11261), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11263) );
  NAND2_X1 U13794 ( .A1(n11263), .A2(n11262), .ZN(n11267) );
  MUX2_X1 U13795 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n11265), .S(n11264), .Z(
        n11266) );
  NAND2_X1 U13796 ( .A1(n11266), .A2(n11267), .ZN(n11963) );
  OAI211_X1 U13797 ( .C1(n11267), .C2(n11266), .A(n14232), .B(n11963), .ZN(
        n11268) );
  OAI211_X1 U13798 ( .C1(n11270), .C2(n14974), .A(n11269), .B(n11268), .ZN(
        P1_U3257) );
  NAND2_X1 U13799 ( .A1(n13379), .A2(n11272), .ZN(n11277) );
  OAI21_X1 U13800 ( .B1(n11687), .B2(n11274), .A(n11273), .ZN(n11275) );
  INV_X1 U13801 ( .A(n11275), .ZN(n11276) );
  NAND2_X1 U13802 ( .A1(n11277), .A2(n11276), .ZN(n11383) );
  XNOR2_X1 U13803 ( .A(n11393), .B(n11383), .ZN(n11278) );
  XNOR2_X1 U13804 ( .A(n15348), .B(n11383), .ZN(n11569) );
  XNOR2_X1 U13805 ( .A(n11569), .B(n15423), .ZN(n11280) );
  AOI21_X1 U13806 ( .B1(n11385), .B2(n11280), .A(n15432), .ZN(n11290) );
  NOR2_X1 U13807 ( .A1(n15298), .A2(n11281), .ZN(n11282) );
  NAND2_X1 U13808 ( .A1(n11283), .A2(n11282), .ZN(n12870) );
  INV_X1 U13809 ( .A(n15343), .ZN(n11284) );
  OAI22_X1 U13810 ( .A1(n11285), .A2(n12870), .B1(n11284), .B2(n12891), .ZN(
        n11288) );
  NOR2_X1 U13811 ( .A1(n11397), .A2(n11286), .ZN(n11287) );
  AOI211_X1 U13812 ( .C1(n15425), .C2(n6805), .A(n11288), .B(n11287), .ZN(
        n11289) );
  OAI21_X1 U13813 ( .B1(n11290), .B2(n15434), .A(n11289), .ZN(P3_U3177) );
  XNOR2_X1 U13814 ( .A(n11291), .B(n11294), .ZN(n11822) );
  OAI21_X1 U13815 ( .B1(n11294), .B2(n11293), .A(n11292), .ZN(n11297) );
  NAND2_X1 U13816 ( .A1(n13522), .A2(n13814), .ZN(n11296) );
  NAND2_X1 U13817 ( .A1(n13520), .A2(n13816), .ZN(n11295) );
  NAND2_X1 U13818 ( .A1(n11296), .A2(n11295), .ZN(n11368) );
  AOI21_X1 U13819 ( .B1(n11297), .B2(n13819), .A(n11368), .ZN(n11813) );
  AOI211_X1 U13820 ( .C1(n11815), .C2(n11834), .A(n8285), .B(n11848), .ZN(
        n11819) );
  AOI21_X1 U13821 ( .B1(n15251), .B2(n11815), .A(n11819), .ZN(n11298) );
  OAI211_X1 U13822 ( .C1(n15249), .C2(n11822), .A(n11813), .B(n11298), .ZN(
        n11345) );
  NAND2_X1 U13823 ( .A1(n11345), .A2(n15279), .ZN(n11299) );
  OAI21_X1 U13824 ( .B1(n15279), .B2(n10583), .A(n11299), .ZN(P2_U3505) );
  INV_X1 U13825 ( .A(n11300), .ZN(n11301) );
  NAND2_X1 U13826 ( .A1(n11302), .A2(n11301), .ZN(n14265) );
  INV_X1 U13827 ( .A(n11303), .ZN(n11304) );
  INV_X1 U13828 ( .A(n11306), .ZN(n11307) );
  INV_X1 U13829 ( .A(n11335), .ZN(n11325) );
  NAND2_X1 U13830 ( .A1(n11326), .A2(n11325), .ZN(n11328) );
  NAND2_X1 U13831 ( .A1(n11478), .A2(n11479), .ZN(n11310) );
  NAND2_X1 U13832 ( .A1(n11328), .A2(n11310), .ZN(n11584) );
  XNOR2_X1 U13833 ( .A(n11584), .B(n11318), .ZN(n15032) );
  INV_X1 U13834 ( .A(n11330), .ZN(n11312) );
  INV_X1 U13835 ( .A(n11587), .ZN(n11583) );
  AND2_X1 U13836 ( .A1(n11330), .A2(n11583), .ZN(n15011) );
  AOI211_X1 U13837 ( .C1(n11587), .C2(n11312), .A(n15014), .B(n15011), .ZN(
        n15033) );
  OAI22_X1 U13838 ( .A1(n15009), .A2(n11583), .B1(n15005), .B2(n11537), .ZN(
        n11314) );
  AOI21_X1 U13839 ( .B1(n15017), .B2(n15033), .A(n11314), .ZN(n11324) );
  NAND2_X1 U13840 ( .A1(n11338), .A2(n11440), .ZN(n11315) );
  NAND2_X1 U13841 ( .A1(n11316), .A2(n11315), .ZN(n11336) );
  NAND2_X1 U13842 ( .A1(n11336), .A2(n11335), .ZN(n11334) );
  NAND2_X1 U13843 ( .A1(n11479), .A2(n14933), .ZN(n11317) );
  XNOR2_X1 U13844 ( .A(n11586), .B(n11318), .ZN(n11319) );
  NAND2_X1 U13845 ( .A1(n11319), .A2(n15052), .ZN(n15034) );
  NAND2_X1 U13846 ( .A1(n14108), .A2(n14479), .ZN(n11320) );
  OAI21_X1 U13847 ( .B1(n11595), .B2(n14464), .A(n11320), .ZN(n11535) );
  INV_X1 U13848 ( .A(n11535), .ZN(n15036) );
  NAND2_X1 U13849 ( .A1(n15034), .A2(n15036), .ZN(n11321) );
  MUX2_X1 U13850 ( .A(n11321), .B(P1_REG2_REG_4__SCAN_IN), .S(n6550), .Z(
        n11322) );
  INV_X1 U13851 ( .A(n11322), .ZN(n11323) );
  OAI211_X1 U13852 ( .C1(n14490), .C2(n15032), .A(n11324), .B(n11323), .ZN(
        P1_U3289) );
  OR2_X1 U13853 ( .A1(n11326), .A2(n11325), .ZN(n11327) );
  NAND2_X1 U13854 ( .A1(n11328), .A2(n11327), .ZN(n11333) );
  INV_X1 U13855 ( .A(n11333), .ZN(n15026) );
  OR2_X1 U13856 ( .A1(n6550), .A2(n11329), .ZN(n14437) );
  AOI211_X1 U13857 ( .C1(n14933), .C2(n11331), .A(n15014), .B(n11330), .ZN(
        n15028) );
  OAI22_X1 U13858 ( .A1(n15009), .A2(n11478), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n15005), .ZN(n11332) );
  AOI21_X1 U13859 ( .B1(n15017), .B2(n15028), .A(n11332), .ZN(n11344) );
  NAND2_X1 U13860 ( .A1(n11333), .A2(n15059), .ZN(n11341) );
  OAI21_X1 U13861 ( .B1(n11336), .B2(n11335), .A(n11334), .ZN(n11339) );
  NAND2_X1 U13862 ( .A1(n14107), .A2(n14477), .ZN(n11337) );
  OAI21_X1 U13863 ( .B1(n11338), .B2(n14462), .A(n11337), .ZN(n14938) );
  AOI21_X1 U13864 ( .B1(n11339), .B2(n15052), .A(n14938), .ZN(n11340) );
  NAND2_X1 U13865 ( .A1(n11341), .A2(n11340), .ZN(n15029) );
  MUX2_X1 U13866 ( .A(n15029), .B(P1_REG2_REG_3__SCAN_IN), .S(n6550), .Z(
        n11342) );
  INV_X1 U13867 ( .A(n11342), .ZN(n11343) );
  OAI211_X1 U13868 ( .C1(n15026), .C2(n14437), .A(n11344), .B(n11343), .ZN(
        P1_U3290) );
  INV_X1 U13869 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n11347) );
  NAND2_X1 U13870 ( .A1(n11345), .A2(n15270), .ZN(n11346) );
  OAI21_X1 U13871 ( .B1(n15270), .B2(n11347), .A(n11346), .ZN(P2_U3448) );
  NOR2_X1 U13872 ( .A1(n11348), .A2(P2_U3088), .ZN(n11419) );
  NAND2_X1 U13873 ( .A1(n13527), .A2(n13814), .ZN(n11350) );
  NAND2_X1 U13874 ( .A1(n13525), .A2(n13816), .ZN(n11349) );
  NAND2_X1 U13875 ( .A1(n11350), .A2(n11349), .ZN(n12063) );
  AOI22_X1 U13876 ( .A1(n6553), .A2(n14848), .B1(n14845), .B2(n12063), .ZN(
        n11355) );
  XNOR2_X1 U13877 ( .A(n11352), .B(n11351), .ZN(n11353) );
  NAND2_X1 U13878 ( .A1(n15120), .A2(n11353), .ZN(n11354) );
  OAI211_X1 U13879 ( .C1(n11419), .C2(n13528), .A(n11355), .B(n11354), .ZN(
        P2_U3194) );
  INV_X1 U13880 ( .A(n11434), .ZN(n11367) );
  NAND2_X1 U13881 ( .A1(n13379), .A2(n11356), .ZN(n11357) );
  NAND2_X1 U13882 ( .A1(n11357), .A2(n11360), .ZN(n11358) );
  INV_X1 U13883 ( .A(n15368), .ZN(n11362) );
  INV_X1 U13884 ( .A(n13249), .ZN(n13209) );
  OAI22_X1 U13885 ( .A1(n15372), .A2(n10763), .B1(n15714), .B2(n15326), .ZN(
        n11364) );
  AOI21_X1 U13886 ( .B1(n13209), .B2(n11365), .A(n11364), .ZN(n11366) );
  OAI21_X1 U13887 ( .B1(n11367), .B2(n13255), .A(n11366), .ZN(P3_U3233) );
  NAND2_X1 U13888 ( .A1(n14845), .A2(n11368), .ZN(n11370) );
  OAI211_X1 U13889 ( .C1(n15124), .C2(n11816), .A(n11370), .B(n11369), .ZN(
        n11375) );
  AOI211_X1 U13890 ( .C1(n11373), .C2(n11372), .A(n13481), .B(n7165), .ZN(
        n11374) );
  AOI211_X1 U13891 ( .C1(n11815), .C2(n14848), .A(n11375), .B(n11374), .ZN(
        n11376) );
  INV_X1 U13892 ( .A(n11376), .ZN(P2_U3211) );
  XOR2_X1 U13893 ( .A(n11378), .B(n11377), .Z(n11382) );
  INV_X1 U13894 ( .A(n14845), .ZN(n13477) );
  INV_X1 U13895 ( .A(n13816), .ZN(n13423) );
  NOR2_X1 U13896 ( .A1(n13477), .A2(n13423), .ZN(n15115) );
  INV_X1 U13897 ( .A(n11419), .ZN(n11379) );
  AOI22_X1 U13898 ( .A1(n15115), .A2(n13524), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n11379), .ZN(n11381) );
  OAI211_X1 U13899 ( .C1(n11382), .C2(n13481), .A(n11381), .B(n11380), .ZN(
        P2_U3209) );
  NAND2_X1 U13900 ( .A1(n11386), .A2(n11384), .ZN(n15361) );
  OAI21_X1 U13901 ( .B1(n11386), .B2(n12640), .A(n11385), .ZN(n11387) );
  OAI21_X1 U13902 ( .B1(n15357), .B2(n11388), .A(n11387), .ZN(n11389) );
  OAI21_X1 U13903 ( .B1(n11571), .B2(n15361), .A(n11389), .ZN(n11390) );
  NAND2_X1 U13904 ( .A1(n11390), .A2(n12861), .ZN(n11395) );
  INV_X1 U13905 ( .A(n15359), .ZN(n11391) );
  OAI22_X1 U13906 ( .A1(n11391), .A2(n12870), .B1(n6804), .B2(n12891), .ZN(
        n11392) );
  AOI21_X1 U13907 ( .B1(n15425), .B2(n11393), .A(n11392), .ZN(n11394) );
  OAI211_X1 U13908 ( .C1(n11397), .C2(n11396), .A(n11395), .B(n11394), .ZN(
        P3_U3162) );
  INV_X1 U13909 ( .A(n11398), .ZN(n11524) );
  INV_X1 U13910 ( .A(n11406), .ZN(n11400) );
  INV_X1 U13911 ( .A(n11399), .ZN(n11618) );
  AOI21_X1 U13912 ( .B1(n11524), .B2(n11400), .A(n11618), .ZN(n11413) );
  INV_X1 U13913 ( .A(n15124), .ZN(n13440) );
  INV_X1 U13914 ( .A(n11770), .ZN(n11411) );
  NAND2_X1 U13915 ( .A1(n14848), .A2(n15227), .ZN(n11405) );
  NAND2_X1 U13916 ( .A1(n13524), .A2(n13814), .ZN(n11402) );
  NAND2_X1 U13917 ( .A1(n13522), .A2(n13816), .ZN(n11401) );
  NAND2_X1 U13918 ( .A1(n11402), .A2(n11401), .ZN(n11764) );
  NAND2_X1 U13919 ( .A1(n14845), .A2(n11764), .ZN(n11403) );
  NAND3_X1 U13920 ( .A1(n11405), .A2(n11404), .A3(n11403), .ZN(n11410) );
  INV_X1 U13921 ( .A(n13496), .ZN(n13488) );
  INV_X1 U13922 ( .A(n13524), .ZN(n11408) );
  NOR4_X1 U13923 ( .A1(n13488), .A2(n11408), .A3(n11407), .A4(n11406), .ZN(
        n11409) );
  AOI211_X1 U13924 ( .C1(n13440), .C2(n11411), .A(n11410), .B(n11409), .ZN(
        n11412) );
  OAI21_X1 U13925 ( .B1(n11413), .B2(n13481), .A(n11412), .ZN(P2_U3202) );
  INV_X1 U13926 ( .A(n13506), .ZN(n15117) );
  NAND2_X1 U13927 ( .A1(n13496), .A2(n13527), .ZN(n11415) );
  MUX2_X1 U13928 ( .A(n15117), .B(n11415), .S(n8105), .Z(n11416) );
  OAI211_X1 U13929 ( .C1(n11419), .C2(n11418), .A(n11417), .B(n11416), .ZN(
        P2_U3204) );
  OAI21_X1 U13930 ( .B1(n11421), .B2(n11420), .A(n11689), .ZN(n12141) );
  OAI211_X1 U13931 ( .C1(n11424), .C2(n11423), .A(n11422), .B(n10380), .ZN(
        n11426) );
  AOI22_X1 U13932 ( .A1(n15360), .A2(n15343), .B1(n11983), .B2(n15358), .ZN(
        n11425) );
  NAND2_X1 U13933 ( .A1(n11426), .A2(n11425), .ZN(n12138) );
  AOI21_X1 U13934 ( .B1(n15405), .B2(n12141), .A(n12138), .ZN(n11431) );
  INV_X1 U13935 ( .A(n15419), .ZN(n15417) );
  OAI22_X1 U13936 ( .A1(n13317), .A2(n12137), .B1(n15419), .B2(n10921), .ZN(
        n11427) );
  INV_X1 U13937 ( .A(n11427), .ZN(n11428) );
  OAI21_X1 U13938 ( .B1(n11431), .B2(n15417), .A(n11428), .ZN(P3_U3463) );
  OAI22_X1 U13939 ( .A1(n12137), .A2(n13376), .B1(n15407), .B2(n8703), .ZN(
        n11429) );
  INV_X1 U13940 ( .A(n11429), .ZN(n11430) );
  OAI21_X1 U13941 ( .B1(n11431), .B2(n15409), .A(n11430), .ZN(P3_U3402) );
  OAI22_X1 U13942 ( .A1(n13317), .A2(n11432), .B1(n15419), .B2(n10762), .ZN(
        n11433) );
  AOI21_X1 U13943 ( .B1(n11434), .B2(n15419), .A(n11433), .ZN(n11435) );
  INV_X1 U13944 ( .A(n11435), .ZN(P3_U3459) );
  MUX2_X1 U13945 ( .A(n11437), .B(n11436), .S(n14498), .Z(n11442) );
  OAI22_X1 U13946 ( .A1(n14383), .A2(n11438), .B1(n14127), .B2(n15005), .ZN(
        n11439) );
  AOI21_X1 U13947 ( .B1(n14889), .B2(n11440), .A(n11439), .ZN(n11441) );
  OAI211_X1 U13948 ( .C1(n11443), .C2(n14437), .A(n11442), .B(n11441), .ZN(
        P1_U3291) );
  INV_X1 U13949 ( .A(n11444), .ZN(n11517) );
  INV_X1 U13950 ( .A(n11452), .ZN(n11445) );
  AOI21_X1 U13951 ( .B1(n11517), .B2(n11445), .A(n6719), .ZN(n11456) );
  NAND2_X1 U13952 ( .A1(n13520), .A2(n13814), .ZN(n11447) );
  NAND2_X1 U13953 ( .A1(n13518), .A2(n13816), .ZN(n11446) );
  NAND2_X1 U13954 ( .A1(n11447), .A2(n11446), .ZN(n11606) );
  NAND2_X1 U13955 ( .A1(n14845), .A2(n11606), .ZN(n11449) );
  OAI211_X1 U13956 ( .C1(n15124), .C2(n11806), .A(n11449), .B(n11448), .ZN(
        n11454) );
  NOR4_X1 U13957 ( .A1(n11452), .A2(n13488), .A3(n11451), .A4(n11450), .ZN(
        n11453) );
  AOI211_X1 U13958 ( .C1(n11611), .C2(n13506), .A(n11454), .B(n11453), .ZN(
        n11455) );
  OAI21_X1 U13959 ( .B1(n11456), .B2(n13481), .A(n11455), .ZN(P2_U3193) );
  AOI21_X1 U13960 ( .B1(n15017), .B2(n11131), .A(n14889), .ZN(n11464) );
  OAI22_X1 U13961 ( .A1(n6550), .A2(n11458), .B1(n11457), .B2(n15005), .ZN(
        n11459) );
  AOI21_X1 U13962 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n6550), .A(n11459), .ZN(
        n11462) );
  NOR2_X1 U13963 ( .A1(n6550), .A2(n15002), .ZN(n14394) );
  OAI21_X1 U13964 ( .B1(n14394), .B2(n14898), .A(n11460), .ZN(n11461) );
  OAI211_X1 U13965 ( .C1(n11464), .C2(n11463), .A(n11462), .B(n11461), .ZN(
        P1_U3293) );
  INV_X1 U13966 ( .A(n13581), .ZN(n13561) );
  INV_X1 U13967 ( .A(n11465), .ZN(n11468) );
  OAI222_X1 U13968 ( .A1(P2_U3088), .A2(n13561), .B1(n12649), .B2(n11468), 
        .C1(n11466), .C2(n13964), .ZN(P2_U3309) );
  INV_X1 U13969 ( .A(n14222), .ZN(n11467) );
  OAI222_X1 U13970 ( .A1(n14635), .A2(n11469), .B1(n14638), .B2(n11468), .C1(
        n11467), .C2(P1_U3086), .ZN(P1_U3337) );
  INV_X1 U13971 ( .A(n11472), .ZN(n11473) );
  NAND2_X1 U13972 ( .A1(n11474), .A2(n11473), .ZN(n11475) );
  OAI22_X1 U13973 ( .A1(n11478), .A2(n11135), .B1(n12779), .B2(n11479), .ZN(
        n11477) );
  XNOR2_X1 U13974 ( .A(n11477), .B(n12777), .ZN(n11480) );
  OAI22_X1 U13975 ( .A1(n12776), .A2(n11479), .B1(n11478), .B2(n12779), .ZN(
        n11481) );
  NAND2_X1 U13976 ( .A1(n11480), .A2(n11481), .ZN(n11486) );
  INV_X1 U13977 ( .A(n11480), .ZN(n11483) );
  INV_X1 U13978 ( .A(n11481), .ZN(n11482) );
  NAND2_X1 U13979 ( .A1(n11483), .A2(n11482), .ZN(n11484) );
  NAND2_X1 U13980 ( .A1(n11486), .A2(n11484), .ZN(n14936) );
  INV_X1 U13981 ( .A(n14107), .ZN(n11588) );
  OAI22_X1 U13982 ( .A1(n12776), .A2(n11588), .B1(n11583), .B2(n12779), .ZN(
        n11491) );
  NAND2_X1 U13983 ( .A1(n11490), .A2(n11491), .ZN(n11530) );
  NAND2_X1 U13984 ( .A1(n12753), .A2(n11587), .ZN(n11488) );
  NAND2_X1 U13985 ( .A1(n12743), .A2(n14107), .ZN(n11487) );
  NAND2_X1 U13986 ( .A1(n11488), .A2(n11487), .ZN(n11489) );
  XNOR2_X1 U13987 ( .A(n11489), .B(n12746), .ZN(n11533) );
  NAND2_X1 U13988 ( .A1(n11530), .A2(n11533), .ZN(n11494) );
  NAND2_X1 U13989 ( .A1(n11494), .A2(n11531), .ZN(n11647) );
  OAI22_X1 U13990 ( .A1(n15008), .A2(n11135), .B1(n11595), .B2(n12779), .ZN(
        n11495) );
  XNOR2_X1 U13991 ( .A(n11495), .B(n12746), .ZN(n11642) );
  OR2_X1 U13992 ( .A1(n15008), .A2(n12779), .ZN(n11497) );
  INV_X2 U13993 ( .A(n12776), .ZN(n12770) );
  NAND2_X1 U13994 ( .A1(n12770), .A2(n14106), .ZN(n11496) );
  AND2_X1 U13995 ( .A1(n11497), .A2(n11496), .ZN(n11641) );
  INV_X1 U13996 ( .A(n11641), .ZN(n11643) );
  XNOR2_X1 U13997 ( .A(n11642), .B(n11643), .ZN(n11498) );
  XNOR2_X1 U13998 ( .A(n11647), .B(n11498), .ZN(n11509) );
  NAND2_X1 U13999 ( .A1(n11133), .A2(n11499), .ZN(n11500) );
  OAI21_X1 U14000 ( .B1(n11501), .B2(n11500), .A(P1_STATE_REG_SCAN_IN), .ZN(
        n11502) );
  NAND2_X1 U14001 ( .A1(n14107), .A2(n14479), .ZN(n11504) );
  NAND2_X1 U14002 ( .A1(n14105), .A2(n14477), .ZN(n11503) );
  NAND2_X1 U14003 ( .A1(n11504), .A2(n11503), .ZN(n15040) );
  AOI21_X1 U14004 ( .B1(n14960), .B2(n15040), .A(n11505), .ZN(n11507) );
  NOR2_X1 U14005 ( .A1(n15008), .A2(n14902), .ZN(n15042) );
  NAND2_X1 U14006 ( .A1(n14953), .A2(n15042), .ZN(n11506) );
  OAI211_X1 U14007 ( .C1(n14965), .C2(n15004), .A(n11507), .B(n11506), .ZN(
        n11508) );
  AOI21_X1 U14008 ( .B1(n11509), .B2(n14961), .A(n11508), .ZN(n11510) );
  INV_X1 U14009 ( .A(n11510), .ZN(P1_U3227) );
  NAND2_X1 U14010 ( .A1(n13521), .A2(n13814), .ZN(n11512) );
  NAND2_X1 U14011 ( .A1(n13519), .A2(n13816), .ZN(n11511) );
  NAND2_X1 U14012 ( .A1(n11512), .A2(n11511), .ZN(n11845) );
  NAND2_X1 U14013 ( .A1(n14845), .A2(n11845), .ZN(n11514) );
  OAI211_X1 U14014 ( .C1(n15124), .C2(n11851), .A(n11514), .B(n11513), .ZN(
        n11521) );
  NAND3_X1 U14015 ( .A1(n13496), .A2(n13521), .A3(n11515), .ZN(n11519) );
  OAI21_X1 U14016 ( .B1(n7165), .B2(n11516), .A(n15120), .ZN(n11518) );
  AOI21_X1 U14017 ( .B1(n11519), .B2(n11518), .A(n11517), .ZN(n11520) );
  AOI211_X1 U14018 ( .C1(n15245), .C2(n14848), .A(n11521), .B(n11520), .ZN(
        n11522) );
  INV_X1 U14019 ( .A(n11522), .ZN(P2_U3185) );
  INV_X1 U14020 ( .A(n15113), .ZN(n13501) );
  AOI22_X1 U14021 ( .A1(n15115), .A2(n13523), .B1(n12043), .B2(n14848), .ZN(
        n11523) );
  OAI21_X1 U14022 ( .B1(n6984), .B2(n13501), .A(n11523), .ZN(n11529) );
  AOI211_X1 U14023 ( .C1(n11526), .C2(n11525), .A(n11524), .B(n13481), .ZN(
        n11528) );
  AOI22_X1 U14024 ( .A1(n15124), .A2(n12042), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_STATE_REG_SCAN_IN), .ZN(n11527) );
  OR3_X1 U14025 ( .A1(n11529), .A2(n11528), .A3(n11527), .ZN(P2_U3190) );
  INV_X1 U14026 ( .A(n14953), .ZN(n14081) );
  NAND2_X1 U14027 ( .A1(n11587), .A2(n14951), .ZN(n15035) );
  NAND2_X1 U14028 ( .A1(n11531), .A2(n11530), .ZN(n11532) );
  XOR2_X1 U14029 ( .A(n11533), .B(n11532), .Z(n11534) );
  NAND2_X1 U14030 ( .A1(n11534), .A2(n14961), .ZN(n11540) );
  AND2_X1 U14031 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14155) );
  AOI21_X1 U14032 ( .B1(n14960), .B2(n11535), .A(n14155), .ZN(n11536) );
  OAI21_X1 U14033 ( .B1(n14965), .B2(n11537), .A(n11536), .ZN(n11538) );
  INV_X1 U14034 ( .A(n11538), .ZN(n11539) );
  OAI211_X1 U14035 ( .C1(n14081), .C2(n15035), .A(n11540), .B(n11539), .ZN(
        P1_U3230) );
  INV_X1 U14036 ( .A(n11541), .ZN(n11544) );
  OAI222_X1 U14037 ( .A1(n14743), .A2(n11544), .B1(n14741), .B2(n11543), .C1(
        P3_U3151), .C2(n11542), .ZN(P3_U3275) );
  INV_X1 U14038 ( .A(n11545), .ZN(n11546) );
  MUX2_X1 U14039 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12946), .Z(n11857) );
  XNOR2_X1 U14040 ( .A(n11857), .B(n11869), .ZN(n11548) );
  AOI21_X1 U14041 ( .B1(n11549), .B2(n11548), .A(n11858), .ZN(n11567) );
  INV_X1 U14042 ( .A(n11869), .ZN(n11860) );
  INV_X1 U14043 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11552) );
  MUX2_X1 U14044 ( .A(P3_REG2_REG_8__SCAN_IN), .B(n11552), .S(n11869), .Z(
        n11553) );
  INV_X1 U14045 ( .A(n11553), .ZN(n11554) );
  AOI21_X1 U14046 ( .B1(n11555), .B2(n11554), .A(n6730), .ZN(n11564) );
  NOR2_X1 U14047 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11556), .ZN(n12197) );
  MUX2_X1 U14048 ( .A(n11559), .B(P3_REG1_REG_8__SCAN_IN), .S(n11869), .Z(
        n11560) );
  AOI21_X1 U14049 ( .B1(n6727), .B2(n11560), .A(n11868), .ZN(n11561) );
  NOR2_X1 U14050 ( .A1(n13004), .A2(n11561), .ZN(n11562) );
  AOI211_X1 U14051 ( .C1(n15280), .C2(P3_ADDR_REG_8__SCAN_IN), .A(n12197), .B(
        n11562), .ZN(n11563) );
  OAI21_X1 U14052 ( .B1(n11564), .B2(n13040), .A(n11563), .ZN(n11565) );
  AOI21_X1 U14053 ( .B1(n11860), .B2(n13041), .A(n11565), .ZN(n11566) );
  OAI21_X1 U14054 ( .B1(n11567), .B2(n13051), .A(n11566), .ZN(P3_U3190) );
  INV_X1 U14055 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n15500) );
  NAND2_X1 U14056 ( .A1(n13104), .A2(P3_U3897), .ZN(n11568) );
  OAI21_X1 U14057 ( .B1(P3_U3897), .B2(n15500), .A(n11568), .ZN(P3_U3517) );
  NOR2_X1 U14058 ( .A1(n11569), .A2(n15423), .ZN(n15431) );
  XNOR2_X1 U14059 ( .A(n11999), .B(n11383), .ZN(n11570) );
  XNOR2_X1 U14060 ( .A(n11570), .B(n15343), .ZN(n15436) );
  AND2_X1 U14061 ( .A1(n11570), .A2(n15343), .ZN(n11574) );
  XNOR2_X1 U14062 ( .A(n12137), .B(n11571), .ZN(n11572) );
  OAI21_X1 U14063 ( .B1(n11699), .B2(n11572), .A(n11739), .ZN(n11573) );
  OAI21_X1 U14064 ( .B1(n15433), .B2(n11574), .A(n11573), .ZN(n11575) );
  INV_X1 U14065 ( .A(n11575), .ZN(n11576) );
  OAI21_X1 U14066 ( .B1(n11740), .B2(n11576), .A(n12861), .ZN(n11582) );
  INV_X1 U14067 ( .A(n11983), .ZN(n11979) );
  AOI21_X1 U14068 ( .B1(n15343), .B2(n15422), .A(n11577), .ZN(n11578) );
  OAI21_X1 U14069 ( .B1(n11979), .B2(n12891), .A(n11578), .ZN(n11579) );
  AOI21_X1 U14070 ( .B1(n11580), .B2(n15425), .A(n11579), .ZN(n11581) );
  OAI211_X1 U14071 ( .C1(n12136), .C2(n12848), .A(n11582), .B(n11581), .ZN(
        P3_U3170) );
  INV_X1 U14072 ( .A(n11717), .ZN(n11591) );
  XNOR2_X1 U14073 ( .A(n11718), .B(n11591), .ZN(n15056) );
  AND2_X1 U14074 ( .A1(n11587), .A2(n11588), .ZN(n11585) );
  OR2_X1 U14075 ( .A1(n11588), .A2(n11587), .ZN(n11589) );
  OR2_X1 U14076 ( .A1(n15008), .A2(n14106), .ZN(n11590) );
  OAI21_X1 U14077 ( .B1(n11592), .B2(n11591), .A(n11724), .ZN(n15053) );
  NAND2_X1 U14078 ( .A1(n15011), .A2(n15008), .ZN(n15012) );
  AND2_X1 U14079 ( .A1(n15012), .A2(n11719), .ZN(n11593) );
  OR3_X1 U14080 ( .A1(n11593), .A2(n14994), .A3(n15014), .ZN(n15050) );
  NOR2_X1 U14081 ( .A1(n15005), .A2(n11660), .ZN(n11597) );
  NAND2_X1 U14082 ( .A1(n14104), .A2(n14477), .ZN(n11594) );
  OAI21_X1 U14083 ( .B1(n11595), .B2(n14462), .A(n11594), .ZN(n15047) );
  MUX2_X1 U14084 ( .A(n15047), .B(P1_REG2_REG_6__SCAN_IN), .S(n6550), .Z(
        n11596) );
  AOI211_X1 U14085 ( .C1(n14889), .C2(n11719), .A(n11597), .B(n11596), .ZN(
        n11598) );
  OAI21_X1 U14086 ( .B1(n14383), .B2(n15050), .A(n11598), .ZN(n11599) );
  AOI21_X1 U14087 ( .B1(n14394), .B2(n15053), .A(n11599), .ZN(n11600) );
  OAI21_X1 U14088 ( .B1(n14490), .B2(n15056), .A(n11600), .ZN(P1_U3287) );
  OAI222_X1 U14089 ( .A1(n14743), .A2(n11602), .B1(n14741), .B2(n11601), .C1(
        P3_U3151), .C2(n11687), .ZN(P3_U3274) );
  XNOR2_X1 U14090 ( .A(n11603), .B(n7803), .ZN(n11812) );
  AOI21_X1 U14091 ( .B1(n11605), .B2(n11604), .A(n13799), .ZN(n11608) );
  AOI21_X1 U14092 ( .B1(n11608), .B2(n11607), .A(n11606), .ZN(n11804) );
  INV_X1 U14093 ( .A(n11849), .ZN(n11610) );
  INV_X1 U14094 ( .A(n12084), .ZN(n11609) );
  AOI211_X1 U14095 ( .C1(n11611), .C2(n11610), .A(n8285), .B(n11609), .ZN(
        n11809) );
  AOI21_X1 U14096 ( .B1(n15251), .B2(n11611), .A(n11809), .ZN(n11612) );
  OAI211_X1 U14097 ( .C1(n15249), .C2(n11812), .A(n11804), .B(n11612), .ZN(
        n11614) );
  NAND2_X1 U14098 ( .A1(n11614), .A2(n15279), .ZN(n11613) );
  OAI21_X1 U14099 ( .B1(n15279), .B2(n10603), .A(n11613), .ZN(P2_U3507) );
  NAND2_X1 U14100 ( .A1(n11614), .A2(n15270), .ZN(n11615) );
  OAI21_X1 U14101 ( .B1(n15270), .B2(n8241), .A(n11615), .ZN(P2_U3454) );
  AOI22_X1 U14102 ( .A1(n13496), .A2(n13523), .B1(n15120), .B2(n11616), .ZN(
        n11619) );
  NOR3_X1 U14103 ( .A1(n11619), .A2(n11618), .A3(n11617), .ZN(n11625) );
  INV_X1 U14104 ( .A(n15115), .ZN(n13503) );
  OAI22_X1 U14105 ( .A1(n13503), .A2(n11620), .B1(n15124), .B2(n11838), .ZN(
        n11624) );
  INV_X1 U14106 ( .A(n11837), .ZN(n15239) );
  NAND2_X1 U14107 ( .A1(n15113), .A2(n13523), .ZN(n11622) );
  OAI211_X1 U14108 ( .C1(n15117), .C2(n15239), .A(n11622), .B(n11621), .ZN(
        n11623) );
  NOR3_X1 U14109 ( .A1(n11625), .A2(n11624), .A3(n11623), .ZN(n11626) );
  OAI21_X1 U14110 ( .B1(n11627), .B2(n13481), .A(n11626), .ZN(P2_U3199) );
  INV_X1 U14111 ( .A(n11628), .ZN(n12648) );
  OAI222_X1 U14112 ( .A1(n14635), .A2(n15594), .B1(n14638), .B2(n12648), .C1(
        P1_U3086), .C2(n14235), .ZN(P1_U3336) );
  NAND2_X1 U14113 ( .A1(n13519), .A2(n13814), .ZN(n11630) );
  NAND2_X1 U14114 ( .A1(n13517), .A2(n13816), .ZN(n11629) );
  AND2_X1 U14115 ( .A1(n11630), .A2(n11629), .ZN(n12080) );
  INV_X1 U14116 ( .A(n12080), .ZN(n11631) );
  AOI22_X1 U14117 ( .A1(n14845), .A2(n11631), .B1(P2_REG3_REG_9__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11632) );
  OAI21_X1 U14118 ( .B1(n12082), .B2(n15124), .A(n11632), .ZN(n11637) );
  AOI22_X1 U14119 ( .A1(n13496), .A2(n13519), .B1(n15120), .B2(n11633), .ZN(
        n11635) );
  NOR3_X1 U14120 ( .A1(n6719), .A2(n11635), .A3(n11634), .ZN(n11636) );
  AOI211_X1 U14121 ( .C1(n15252), .C2(n14848), .A(n11637), .B(n11636), .ZN(
        n11638) );
  OAI21_X1 U14122 ( .B1(n11639), .B2(n13481), .A(n11638), .ZN(P2_U3203) );
  NAND2_X1 U14123 ( .A1(n12902), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n11640) );
  OAI21_X1 U14124 ( .B1(n12798), .B2(n12902), .A(n11640), .ZN(P3_U3519) );
  NAND2_X1 U14125 ( .A1(n11719), .A2(n14951), .ZN(n15048) );
  AND2_X1 U14126 ( .A1(n11642), .A2(n11641), .ZN(n11646) );
  INV_X1 U14127 ( .A(n11642), .ZN(n11644) );
  NAND2_X1 U14128 ( .A1(n11644), .A2(n11643), .ZN(n11645) );
  NAND2_X1 U14129 ( .A1(n11719), .A2(n12753), .ZN(n11649) );
  NAND2_X1 U14130 ( .A1(n12743), .A2(n14105), .ZN(n11648) );
  NAND2_X1 U14131 ( .A1(n11649), .A2(n11648), .ZN(n11650) );
  XNOR2_X1 U14132 ( .A(n11650), .B(n12777), .ZN(n11653) );
  NAND2_X1 U14133 ( .A1(n11719), .A2(n12743), .ZN(n11652) );
  NAND2_X1 U14134 ( .A1(n12770), .A2(n14105), .ZN(n11651) );
  NAND2_X1 U14135 ( .A1(n11652), .A2(n11651), .ZN(n11654) );
  INV_X1 U14136 ( .A(n11653), .ZN(n11656) );
  INV_X1 U14137 ( .A(n11654), .ZN(n11655) );
  NAND2_X1 U14138 ( .A1(n11656), .A2(n11655), .ZN(n11666) );
  NAND2_X1 U14139 ( .A1(n6736), .A2(n11666), .ZN(n11657) );
  XNOR2_X1 U14140 ( .A(n11667), .B(n11657), .ZN(n11658) );
  NAND2_X1 U14141 ( .A1(n11658), .A2(n14961), .ZN(n11663) );
  AND2_X1 U14142 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n14180) );
  AOI21_X1 U14143 ( .B1(n14960), .B2(n15047), .A(n14180), .ZN(n11659) );
  OAI21_X1 U14144 ( .B1(n14965), .B2(n11660), .A(n11659), .ZN(n11661) );
  INV_X1 U14145 ( .A(n11661), .ZN(n11662) );
  OAI211_X1 U14146 ( .C1(n14081), .C2(n15048), .A(n11663), .B(n11662), .ZN(
        P1_U3239) );
  NAND2_X1 U14147 ( .A1(n12902), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n11664) );
  OAI21_X1 U14148 ( .B1(n11665), .B2(n12902), .A(n11664), .ZN(P3_U3521) );
  NAND2_X1 U14149 ( .A1(n11734), .A2(n14951), .ZN(n15061) );
  NAND2_X1 U14150 ( .A1(n11734), .A2(n12753), .ZN(n11669) );
  NAND2_X1 U14151 ( .A1(n12743), .A2(n14104), .ZN(n11668) );
  NAND2_X1 U14152 ( .A1(n11669), .A2(n11668), .ZN(n11670) );
  XNOR2_X1 U14153 ( .A(n11670), .B(n12746), .ZN(n12287) );
  INV_X1 U14154 ( .A(n14104), .ZN(n11725) );
  NOR2_X1 U14155 ( .A1(n12776), .A2(n11725), .ZN(n11671) );
  AOI21_X1 U14156 ( .B1(n11734), .B2(n12743), .A(n11671), .ZN(n12288) );
  XNOR2_X1 U14157 ( .A(n12287), .B(n12288), .ZN(n11673) );
  AOI21_X1 U14158 ( .B1(n11672), .B2(n11673), .A(n14935), .ZN(n11675) );
  NAND2_X1 U14159 ( .A1(n11675), .A2(n12292), .ZN(n11681) );
  NAND2_X1 U14160 ( .A1(n14105), .A2(n14479), .ZN(n11677) );
  NAND2_X1 U14161 ( .A1(n14103), .A2(n14477), .ZN(n11676) );
  NAND2_X1 U14162 ( .A1(n11677), .A2(n11676), .ZN(n15060) );
  NOR2_X1 U14163 ( .A1(n11678), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14195) );
  NOR2_X1 U14164 ( .A1(n14965), .A2(n14988), .ZN(n11679) );
  AOI211_X1 U14165 ( .C1(n14960), .C2(n15060), .A(n14195), .B(n11679), .ZN(
        n11680) );
  OAI211_X1 U14166 ( .C1(n14081), .C2(n15061), .A(n11681), .B(n11680), .ZN(
        P1_U3213) );
  NOR2_X1 U14167 ( .A1(n14741), .A2(SI_22_), .ZN(n11682) );
  AOI21_X1 U14168 ( .B1(n11683), .B2(P3_STATE_REG_SCAN_IN), .A(n11682), .ZN(
        n11684) );
  OAI21_X1 U14169 ( .B1(n11685), .B2(n14743), .A(n11684), .ZN(n11686) );
  INV_X1 U14170 ( .A(n11686), .ZN(P3_U3273) );
  NOR2_X1 U14171 ( .A1(n11687), .A2(n15368), .ZN(n15349) );
  NAND2_X1 U14172 ( .A1(n15372), .A2(n15349), .ZN(n13081) );
  NAND2_X1 U14173 ( .A1(n15372), .A2(n15363), .ZN(n11688) );
  NAND2_X1 U14174 ( .A1(n11689), .A2(n11691), .ZN(n11690) );
  MUX2_X1 U14175 ( .A(n11691), .B(n11690), .S(n6801), .Z(n11693) );
  NAND2_X1 U14176 ( .A1(n11693), .A2(n11692), .ZN(n15389) );
  INV_X1 U14177 ( .A(n15389), .ZN(n11704) );
  INV_X1 U14178 ( .A(n15331), .ZN(n12003) );
  INV_X1 U14179 ( .A(n11694), .ZN(n11695) );
  AOI21_X1 U14180 ( .B1(n11697), .B2(n11696), .A(n11695), .ZN(n11698) );
  OAI222_X1 U14181 ( .A1(n15300), .A2(n12003), .B1(n15298), .B2(n11699), .C1(
        n15366), .C2(n11698), .ZN(n15387) );
  NOR2_X1 U14182 ( .A1(n15372), .A2(n10911), .ZN(n11702) );
  AND2_X1 U14183 ( .A1(n11746), .A2(n13290), .ZN(n15388) );
  NAND2_X1 U14184 ( .A1(n15336), .A2(n15388), .ZN(n11700) );
  OAI21_X1 U14185 ( .B1(n11744), .B2(n15326), .A(n11700), .ZN(n11701) );
  AOI211_X1 U14186 ( .C1(n15387), .C2(n15372), .A(n11702), .B(n11701), .ZN(
        n11703) );
  OAI21_X1 U14187 ( .B1(n13214), .B2(n11704), .A(n11703), .ZN(P3_U3228) );
  OAI21_X1 U14188 ( .B1(n11707), .B2(n11706), .A(n11705), .ZN(n12148) );
  OAI211_X1 U14189 ( .C1(n6728), .C2(n11709), .A(n11708), .B(n10380), .ZN(
        n11711) );
  AOI22_X1 U14190 ( .A1(n15360), .A2(n11983), .B1(n15310), .B2(n15358), .ZN(
        n11710) );
  NAND2_X1 U14191 ( .A1(n11711), .A2(n11710), .ZN(n12145) );
  AOI21_X1 U14192 ( .B1(n15405), .B2(n12148), .A(n12145), .ZN(n11716) );
  OAI22_X1 U14193 ( .A1(n12144), .A2(n13376), .B1(n15407), .B2(n8738), .ZN(
        n11712) );
  INV_X1 U14194 ( .A(n11712), .ZN(n11713) );
  OAI21_X1 U14195 ( .B1(n11716), .B2(n15409), .A(n11713), .ZN(P3_U3408) );
  OAI22_X1 U14196 ( .A1(n13317), .A2(n12144), .B1(n15419), .B2(n11209), .ZN(
        n11714) );
  INV_X1 U14197 ( .A(n11714), .ZN(n11715) );
  OAI21_X1 U14198 ( .B1(n11716), .B2(n15417), .A(n11715), .ZN(P3_U3465) );
  INV_X1 U14199 ( .A(n14985), .ZN(n14982) );
  NAND2_X1 U14200 ( .A1(n14983), .A2(n14982), .ZN(n11721) );
  OR2_X1 U14201 ( .A1(n11734), .A2(n14104), .ZN(n11720) );
  NAND2_X1 U14202 ( .A1(n11721), .A2(n11720), .ZN(n11880) );
  XNOR2_X1 U14203 ( .A(n11880), .B(n11722), .ZN(n15068) );
  INV_X1 U14204 ( .A(n11722), .ZN(n11879) );
  NAND2_X1 U14205 ( .A1(n11724), .A2(n11723), .ZN(n14986) );
  NAND2_X1 U14206 ( .A1(n14986), .A2(n14985), .ZN(n14984) );
  NAND2_X1 U14207 ( .A1(n11734), .A2(n11725), .ZN(n11726) );
  INV_X1 U14208 ( .A(n11729), .ZN(n11727) );
  INV_X1 U14209 ( .A(n11886), .ZN(n11728) );
  AOI211_X1 U14210 ( .C1(n11879), .C2(n11729), .A(n15002), .B(n11728), .ZN(
        n15072) );
  NAND2_X1 U14211 ( .A1(n14104), .A2(n14479), .ZN(n11731) );
  NAND2_X1 U14212 ( .A1(n14102), .A2(n14477), .ZN(n11730) );
  NAND2_X1 U14213 ( .A1(n11731), .A2(n11730), .ZN(n15069) );
  NOR2_X1 U14214 ( .A1(n15072), .A2(n15069), .ZN(n11732) );
  MUX2_X1 U14215 ( .A(n11733), .B(n11732), .S(n14498), .Z(n11738) );
  INV_X1 U14216 ( .A(n11734), .ZN(n14993) );
  NAND2_X1 U14217 ( .A1(n14994), .A2(n14993), .ZN(n14992) );
  AOI211_X1 U14218 ( .C1(n14943), .C2(n14992), .A(n15014), .B(n7331), .ZN(
        n15071) );
  INV_X1 U14219 ( .A(n14943), .ZN(n11735) );
  OAI22_X1 U14220 ( .A1(n15009), .A2(n11735), .B1(n14950), .B2(n15005), .ZN(
        n11736) );
  AOI21_X1 U14221 ( .B1(n15071), .B2(n15017), .A(n11736), .ZN(n11737) );
  OAI211_X1 U14222 ( .C1(n15068), .C2(n14490), .A(n11738), .B(n11737), .ZN(
        P1_U3285) );
  XNOR2_X1 U14223 ( .A(n11746), .B(n12640), .ZN(n11978) );
  XOR2_X1 U14224 ( .A(n11983), .B(n11978), .Z(n11741) );
  AOI21_X1 U14225 ( .B1(n11742), .B2(n11741), .A(n12011), .ZN(n11752) );
  AOI21_X1 U14226 ( .B1(n15421), .B2(n15422), .A(n11743), .ZN(n11750) );
  INV_X1 U14227 ( .A(n11744), .ZN(n11745) );
  NAND2_X1 U14228 ( .A1(n15439), .A2(n11745), .ZN(n11749) );
  NAND2_X1 U14229 ( .A1(n15425), .A2(n11746), .ZN(n11748) );
  INV_X1 U14230 ( .A(n12891), .ZN(n15420) );
  NAND2_X1 U14231 ( .A1(n15331), .A2(n15420), .ZN(n11747) );
  AND4_X1 U14232 ( .A1(n11750), .A2(n11749), .A3(n11748), .A4(n11747), .ZN(
        n11751) );
  OAI21_X1 U14233 ( .B1(n11752), .B2(n15434), .A(n11751), .ZN(P3_U3167) );
  NAND3_X1 U14234 ( .A1(n15209), .A2(n11754), .A3(n11753), .ZN(n11755) );
  OR2_X1 U14235 ( .A1(n11756), .A2(n11755), .ZN(n11757) );
  NAND2_X1 U14236 ( .A1(n15256), .A2(n11824), .ZN(n11759) );
  XNOR2_X1 U14237 ( .A(n11760), .B(n11763), .ZN(n15230) );
  OAI21_X1 U14238 ( .B1(n11763), .B2(n11762), .A(n11761), .ZN(n11765) );
  AOI21_X1 U14239 ( .B1(n11765), .B2(n13819), .A(n11764), .ZN(n15234) );
  MUX2_X1 U14240 ( .A(n11766), .B(n15234), .S(n13770), .Z(n11774) );
  OR2_X1 U14241 ( .A1(n11767), .A2(n11771), .ZN(n11768) );
  AND3_X1 U14242 ( .A1(n11768), .A2(n11836), .A3(n13690), .ZN(n15229) );
  OAI22_X1 U14243 ( .A1(n13828), .A2(n11771), .B1(n13784), .B2(n11770), .ZN(
        n11772) );
  AOI21_X1 U14244 ( .B1(n13835), .B2(n15229), .A(n11772), .ZN(n11773) );
  OAI211_X1 U14245 ( .C1(n13832), .C2(n15230), .A(n11774), .B(n11773), .ZN(
        P2_U3261) );
  INV_X1 U14246 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n15656) );
  INV_X1 U14247 ( .A(n13074), .ZN(n11775) );
  NAND2_X1 U14248 ( .A1(n11775), .A2(P3_U3897), .ZN(n11776) );
  OAI21_X1 U14249 ( .B1(P3_U3897), .B2(n15656), .A(n11776), .ZN(P3_U3520) );
  XNOR2_X1 U14250 ( .A(n11777), .B(n11786), .ZN(n13924) );
  OAI21_X1 U14251 ( .B1(n12066), .B2(n11781), .A(n13690), .ZN(n11779) );
  NOR2_X1 U14252 ( .A1(n11779), .A2(n11778), .ZN(n13921) );
  OAI22_X1 U14253 ( .A1(n13770), .A2(n10437), .B1(n11780), .B2(n13784), .ZN(
        n11783) );
  NOR2_X1 U14254 ( .A1(n13828), .A2(n11781), .ZN(n11782) );
  AOI211_X1 U14255 ( .C1(n13921), .C2(n13835), .A(n11783), .B(n11782), .ZN(
        n11791) );
  OAI21_X1 U14256 ( .B1(n11786), .B2(n11785), .A(n11784), .ZN(n11787) );
  NAND2_X1 U14257 ( .A1(n11787), .A2(n13819), .ZN(n11789) );
  NAND2_X1 U14258 ( .A1(n11789), .A2(n11788), .ZN(n13920) );
  NAND2_X1 U14259 ( .A1(n13770), .A2(n13920), .ZN(n11790) );
  OAI211_X1 U14260 ( .C1(n13924), .C2(n13832), .A(n11791), .B(n11790), .ZN(
        P2_U3263) );
  OAI21_X1 U14261 ( .B1(n11928), .B2(n11794), .A(n11792), .ZN(n11802) );
  NOR3_X1 U14262 ( .A1(n11794), .A2(n11793), .A3(n13488), .ZN(n11795) );
  OAI21_X1 U14263 ( .B1(n11795), .B2(n15113), .A(n13517), .ZN(n11800) );
  INV_X1 U14264 ( .A(n11796), .ZN(n12130) );
  OAI21_X1 U14265 ( .B1(n13503), .B2(n12121), .A(n11797), .ZN(n11798) );
  AOI21_X1 U14266 ( .B1(n12130), .B2(n13440), .A(n11798), .ZN(n11799) );
  OAI211_X1 U14267 ( .C1(n12132), .C2(n15117), .A(n11800), .B(n11799), .ZN(
        n11801) );
  AOI21_X1 U14268 ( .B1(n15120), .B2(n11802), .A(n11801), .ZN(n11803) );
  INV_X1 U14269 ( .A(n11803), .ZN(P2_U3208) );
  MUX2_X1 U14270 ( .A(n11805), .B(n11804), .S(n13770), .Z(n11811) );
  OAI22_X1 U14271 ( .A1(n13828), .A2(n11807), .B1(n11806), .B2(n13784), .ZN(
        n11808) );
  AOI21_X1 U14272 ( .B1(n11809), .B2(n13835), .A(n11808), .ZN(n11810) );
  OAI211_X1 U14273 ( .C1(n13832), .C2(n11812), .A(n11811), .B(n11810), .ZN(
        P2_U3257) );
  MUX2_X1 U14274 ( .A(n11814), .B(n11813), .S(n13770), .Z(n11821) );
  INV_X1 U14275 ( .A(n11815), .ZN(n11817) );
  OAI22_X1 U14276 ( .A1(n13828), .A2(n11817), .B1(n13784), .B2(n11816), .ZN(
        n11818) );
  AOI21_X1 U14277 ( .B1(n11819), .B2(n13835), .A(n11818), .ZN(n11820) );
  OAI211_X1 U14278 ( .C1(n11822), .C2(n13832), .A(n11821), .B(n11820), .ZN(
        P2_U3259) );
  XNOR2_X1 U14279 ( .A(n11823), .B(n11827), .ZN(n15236) );
  INV_X1 U14280 ( .A(n11824), .ZN(n11825) );
  NAND2_X1 U14281 ( .A1(n13770), .A2(n11825), .ZN(n13808) );
  AOI22_X1 U14282 ( .A1(n13814), .A2(n13523), .B1(n13521), .B2(n13816), .ZN(
        n11831) );
  OAI21_X1 U14283 ( .B1(n11828), .B2(n11827), .A(n11826), .ZN(n11829) );
  NAND2_X1 U14284 ( .A1(n11829), .A2(n13819), .ZN(n11830) );
  OAI211_X1 U14285 ( .C1(n15236), .C2(n15256), .A(n11831), .B(n11830), .ZN(
        n15240) );
  INV_X1 U14286 ( .A(n15240), .ZN(n11832) );
  MUX2_X1 U14287 ( .A(n11833), .B(n11832), .S(n13770), .Z(n11841) );
  INV_X1 U14288 ( .A(n11834), .ZN(n11835) );
  AOI211_X1 U14289 ( .C1(n11837), .C2(n11836), .A(n8285), .B(n11835), .ZN(
        n15237) );
  OAI22_X1 U14290 ( .A1(n13828), .A2(n15239), .B1(n13784), .B2(n11838), .ZN(
        n11839) );
  AOI21_X1 U14291 ( .B1(n15237), .B2(n13835), .A(n11839), .ZN(n11840) );
  OAI211_X1 U14292 ( .C1(n15236), .C2(n13808), .A(n11841), .B(n11840), .ZN(
        P2_U3260) );
  XNOR2_X1 U14293 ( .A(n11842), .B(n11843), .ZN(n15248) );
  XNOR2_X1 U14294 ( .A(n11844), .B(n11843), .ZN(n11846) );
  AOI21_X1 U14295 ( .B1(n11846), .B2(n13819), .A(n11845), .ZN(n15247) );
  MUX2_X1 U14296 ( .A(n11847), .B(n15247), .S(n13770), .Z(n11855) );
  OAI21_X1 U14297 ( .B1(n11848), .B2(n11852), .A(n13690), .ZN(n11850) );
  NOR2_X1 U14298 ( .A1(n11850), .A2(n11849), .ZN(n15244) );
  OAI22_X1 U14299 ( .A1(n13828), .A2(n11852), .B1(n13784), .B2(n11851), .ZN(
        n11853) );
  AOI21_X1 U14300 ( .B1(n15244), .B2(n13835), .A(n11853), .ZN(n11854) );
  OAI211_X1 U14301 ( .C1(n13832), .C2(n15248), .A(n11855), .B(n11854), .ZN(
        P2_U3258) );
  AOI21_X1 U14302 ( .B1(n11862), .B2(n11856), .A(n11900), .ZN(n11878) );
  INV_X1 U14303 ( .A(n11857), .ZN(n11859) );
  MUX2_X1 U14304 ( .A(n11862), .B(n11861), .S(n12946), .Z(n11863) );
  NOR2_X1 U14305 ( .A1(n11863), .A2(n11913), .ZN(n11865) );
  NOR2_X1 U14306 ( .A1(n11864), .A2(n11865), .ZN(n11905) );
  INV_X1 U14307 ( .A(n11905), .ZN(n11867) );
  AND2_X1 U14308 ( .A1(n11863), .A2(n11913), .ZN(n11904) );
  OAI21_X1 U14309 ( .B1(n11904), .B2(n11865), .A(n11864), .ZN(n11866) );
  OAI21_X1 U14310 ( .B1(n11867), .B2(n11904), .A(n11866), .ZN(n11876) );
  AOI21_X1 U14311 ( .B1(n11861), .B2(n11870), .A(n11914), .ZN(n11871) );
  NOR2_X1 U14312 ( .A1(n11871), .A2(n13004), .ZN(n11875) );
  AND2_X1 U14313 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n12014) );
  AOI21_X1 U14314 ( .B1(n15280), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n12014), .ZN(
        n11872) );
  OAI21_X1 U14315 ( .B1(n12935), .B2(n11873), .A(n11872), .ZN(n11874) );
  AOI211_X1 U14316 ( .C1(n11876), .C2(n12916), .A(n11875), .B(n11874), .ZN(
        n11877) );
  OAI21_X1 U14317 ( .B1(n11878), .B2(n13040), .A(n11877), .ZN(P3_U3191) );
  NAND2_X1 U14318 ( .A1(n11880), .A2(n11879), .ZN(n11882) );
  OR2_X1 U14319 ( .A1(n14943), .A2(n14103), .ZN(n11881) );
  NAND2_X1 U14320 ( .A1(n11882), .A2(n11881), .ZN(n11936) );
  INV_X1 U14321 ( .A(n11935), .ZN(n11941) );
  NAND2_X1 U14322 ( .A1(n11936), .A2(n11941), .ZN(n11884) );
  OR2_X1 U14323 ( .A1(n14952), .A2(n14102), .ZN(n11883) );
  NAND2_X1 U14324 ( .A1(n11884), .A2(n11883), .ZN(n12024) );
  INV_X1 U14325 ( .A(n12023), .ZN(n11887) );
  XNOR2_X1 U14326 ( .A(n12024), .B(n11887), .ZN(n15086) );
  INV_X1 U14327 ( .A(n14102), .ZN(n12302) );
  OAI211_X1 U14328 ( .C1(n11888), .C2(n11887), .A(n15052), .B(n12029), .ZN(
        n15091) );
  NAND2_X1 U14329 ( .A1(n14102), .A2(n14479), .ZN(n14877) );
  AOI21_X1 U14330 ( .B1(n15091), .B2(n14877), .A(n6550), .ZN(n11889) );
  INV_X1 U14331 ( .A(n11889), .ZN(n11895) );
  OAI22_X1 U14332 ( .A1(n14498), .A2(n11890), .B1(n14882), .B2(n15005), .ZN(
        n11893) );
  AOI21_X1 U14333 ( .B1(n14870), .B2(n11937), .A(n15014), .ZN(n11891) );
  NAND2_X1 U14334 ( .A1(n11891), .A2(n14893), .ZN(n15089) );
  NAND2_X1 U14335 ( .A1(n14100), .A2(n14477), .ZN(n14878) );
  AOI21_X1 U14336 ( .B1(n15089), .B2(n14878), .A(n14383), .ZN(n11892) );
  AOI211_X1 U14337 ( .C1(n14889), .C2(n14870), .A(n11893), .B(n11892), .ZN(
        n11894) );
  OAI211_X1 U14338 ( .C1(n15086), .C2(n14490), .A(n11895), .B(n11894), .ZN(
        P1_U3283) );
  INV_X1 U14339 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11898) );
  INV_X1 U14340 ( .A(n11896), .ZN(n11923) );
  OAI222_X1 U14341 ( .A1(n14635), .A2(n11898), .B1(n14638), .B2(n11923), .C1(
        n11897), .C2(P1_U3086), .ZN(P1_U3335) );
  NOR2_X1 U14342 ( .A1(n11913), .A2(n11899), .ZN(n11901) );
  AOI22_X1 U14343 ( .A1(n12351), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n8803), 
        .B2(n14756), .ZN(n11902) );
  AOI21_X1 U14344 ( .B1(n11903), .B2(n11902), .A(n6729), .ZN(n11922) );
  MUX2_X1 U14345 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12946), .Z(n12348) );
  XNOR2_X1 U14346 ( .A(n12348), .B(n14756), .ZN(n11906) );
  AOI21_X1 U14347 ( .B1(n11907), .B2(n11906), .A(n12349), .ZN(n11911) );
  INV_X1 U14348 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n11908) );
  NOR2_X1 U14349 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11908), .ZN(n12184) );
  NOR2_X1 U14350 ( .A1(n12935), .A2(n14756), .ZN(n11909) );
  AOI211_X1 U14351 ( .C1(n15280), .C2(P3_ADDR_REG_10__SCAN_IN), .A(n12184), 
        .B(n11909), .ZN(n11910) );
  OAI21_X1 U14352 ( .B1(n11911), .B2(n13051), .A(n11910), .ZN(n11920) );
  NOR2_X1 U14353 ( .A1(n11913), .A2(n11912), .ZN(n11915) );
  AOI22_X1 U14354 ( .A1(n12351), .A2(P3_REG1_REG_10__SCAN_IN), .B1(n8800), 
        .B2(n14756), .ZN(n11916) );
  AOI21_X1 U14355 ( .B1(n11917), .B2(n11916), .A(n6726), .ZN(n11918) );
  NOR2_X1 U14356 ( .A1(n11918), .A2(n13004), .ZN(n11919) );
  NOR2_X1 U14357 ( .A1(n11920), .A2(n11919), .ZN(n11921) );
  OAI21_X1 U14358 ( .B1(n11922), .B2(n13040), .A(n11921), .ZN(P3_U3192) );
  OAI222_X1 U14359 ( .A1(n13964), .A2(n15645), .B1(P2_U3088), .B2(n8079), .C1(
        n12649), .C2(n11923), .ZN(P2_U3307) );
  INV_X1 U14360 ( .A(n12096), .ZN(n11924) );
  AOI22_X1 U14361 ( .A1(n15113), .A2(n13518), .B1(n13440), .B2(n11924), .ZN(
        n11926) );
  OAI211_X1 U14362 ( .C1(n13503), .C2(n11927), .A(n11926), .B(n11925), .ZN(
        n11933) );
  INV_X1 U14363 ( .A(n11928), .ZN(n11929) );
  AOI211_X1 U14364 ( .C1(n11931), .C2(n11930), .A(n13481), .B(n11929), .ZN(
        n11932) );
  AOI211_X1 U14365 ( .C1(n12102), .C2(n13506), .A(n11933), .B(n11932), .ZN(
        n11934) );
  INV_X1 U14366 ( .A(n11934), .ZN(P2_U3189) );
  XNOR2_X1 U14367 ( .A(n11936), .B(n11935), .ZN(n15080) );
  INV_X1 U14368 ( .A(n14399), .ZN(n11946) );
  AOI21_X1 U14369 ( .B1(n14952), .B2(n11938), .A(n7329), .ZN(n15078) );
  AOI21_X1 U14370 ( .B1(n11941), .B2(n11940), .A(n11939), .ZN(n11945) );
  NAND2_X1 U14371 ( .A1(n14103), .A2(n14479), .ZN(n11943) );
  NAND2_X1 U14372 ( .A1(n14101), .A2(n14477), .ZN(n11942) );
  NAND2_X1 U14373 ( .A1(n11943), .A2(n11942), .ZN(n14959) );
  INV_X1 U14374 ( .A(n14959), .ZN(n11944) );
  OAI21_X1 U14375 ( .B1(n11945), .B2(n15002), .A(n11944), .ZN(n15076) );
  AOI21_X1 U14376 ( .B1(n11946), .B2(n15078), .A(n15076), .ZN(n11947) );
  MUX2_X1 U14377 ( .A(n10790), .B(n11947), .S(n14498), .Z(n11950) );
  INV_X1 U14378 ( .A(n15005), .ZN(n14888) );
  INV_X1 U14379 ( .A(n14966), .ZN(n11948) );
  AOI22_X1 U14380 ( .A1(n14889), .A2(n14952), .B1(n14888), .B2(n11948), .ZN(
        n11949) );
  OAI211_X1 U14381 ( .C1(n14490), .C2(n15080), .A(n11950), .B(n11949), .ZN(
        P1_U3284) );
  INV_X1 U14382 ( .A(n13835), .ZN(n13724) );
  INV_X1 U14383 ( .A(n13808), .ZN(n11955) );
  INV_X1 U14384 ( .A(n13784), .ZN(n13825) );
  NAND2_X1 U14385 ( .A1(n13825), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n11952) );
  NAND2_X1 U14386 ( .A1(n13799), .A2(n15256), .ZN(n11951) );
  OAI211_X1 U14387 ( .C1(n15213), .C2(n8079), .A(n11952), .B(n15214), .ZN(
        n11953) );
  MUX2_X1 U14388 ( .A(P2_REG2_REG_0__SCAN_IN), .B(n11953), .S(n13770), .Z(
        n11954) );
  AOI21_X1 U14389 ( .B1(n11955), .B2(n15217), .A(n11954), .ZN(n11956) );
  OAI21_X1 U14390 ( .B1(n15213), .B2(n13724), .A(n11956), .ZN(P2_U3265) );
  XNOR2_X1 U14391 ( .A(n12151), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n12156) );
  AOI21_X1 U14392 ( .B1(n11964), .B2(n15528), .A(n11957), .ZN(n11958) );
  NOR2_X1 U14393 ( .A1(n11965), .A2(n11958), .ZN(n11959) );
  XNOR2_X1 U14394 ( .A(n11958), .B(n11965), .ZN(n14968) );
  NOR2_X1 U14395 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n14968), .ZN(n14967) );
  NOR2_X1 U14396 ( .A1(n11959), .A2(n14967), .ZN(n12157) );
  XOR2_X1 U14397 ( .A(n12156), .B(n12157), .Z(n11960) );
  NAND2_X1 U14398 ( .A1(n11960), .A2(n14233), .ZN(n11973) );
  NAND2_X1 U14399 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14018)
         );
  INV_X1 U14400 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n14470) );
  NAND2_X1 U14401 ( .A1(n12151), .A2(n14470), .ZN(n11961) );
  OAI21_X1 U14402 ( .B1(n12151), .B2(n14470), .A(n11961), .ZN(n11962) );
  INV_X1 U14403 ( .A(n11962), .ZN(n11969) );
  OAI21_X1 U14404 ( .B1(n11265), .B2(n11964), .A(n11963), .ZN(n11966) );
  NOR2_X1 U14405 ( .A1(n11965), .A2(n11966), .ZN(n11967) );
  XOR2_X1 U14406 ( .A(n11966), .B(n14975), .Z(n14970) );
  NOR2_X1 U14407 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14970), .ZN(n14969) );
  NOR2_X1 U14408 ( .A1(n11967), .A2(n14969), .ZN(n11968) );
  NAND2_X1 U14409 ( .A1(n11968), .A2(n11969), .ZN(n12150) );
  OAI211_X1 U14410 ( .C1(n11969), .C2(n11968), .A(n14232), .B(n12150), .ZN(
        n11970) );
  NAND2_X1 U14411 ( .A1(n14018), .A2(n11970), .ZN(n11971) );
  AOI21_X1 U14412 ( .B1(n14212), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11971), 
        .ZN(n11972) );
  OAI211_X1 U14413 ( .C1(n14976), .C2(n12151), .A(n11973), .B(n11972), .ZN(
        P1_U3259) );
  NAND2_X1 U14414 ( .A1(n11974), .A2(n14762), .ZN(n11976) );
  OAI211_X1 U14415 ( .C1(n11977), .C2(n14741), .A(n11976), .B(n11975), .ZN(
        P3_U3272) );
  NAND2_X1 U14416 ( .A1(n11979), .A2(n11978), .ZN(n12005) );
  INV_X1 U14417 ( .A(n12005), .ZN(n11980) );
  NOR2_X1 U14418 ( .A1(n12011), .A2(n11980), .ZN(n11982) );
  XNOR2_X1 U14419 ( .A(n12144), .B(n12640), .ZN(n12006) );
  XNOR2_X1 U14420 ( .A(n12006), .B(n12003), .ZN(n11981) );
  NAND2_X1 U14421 ( .A1(n11982), .A2(n11981), .ZN(n12107) );
  OAI211_X1 U14422 ( .C1(n11982), .C2(n11981), .A(n12107), .B(n12861), .ZN(
        n11990) );
  NAND2_X1 U14423 ( .A1(n15310), .A2(n15420), .ZN(n11988) );
  NAND2_X1 U14424 ( .A1(n11983), .A2(n15422), .ZN(n11987) );
  NAND2_X1 U14425 ( .A1(n15425), .A2(n11984), .ZN(n11986) );
  AND4_X1 U14426 ( .A1(n11988), .A2(n11987), .A3(n11986), .A4(n11985), .ZN(
        n11989) );
  OAI211_X1 U14427 ( .C1(n12143), .C2(n12848), .A(n11990), .B(n11989), .ZN(
        P3_U3179) );
  XOR2_X1 U14428 ( .A(n11992), .B(n11991), .Z(n15383) );
  NAND2_X1 U14429 ( .A1(n11993), .A2(n11992), .ZN(n11994) );
  NAND3_X1 U14430 ( .A1(n11995), .A2(n10380), .A3(n11994), .ZN(n11997) );
  AOI22_X1 U14431 ( .A1(n15360), .A2(n15423), .B1(n15421), .B2(n15358), .ZN(
        n11996) );
  NAND2_X1 U14432 ( .A1(n11997), .A2(n11996), .ZN(n15384) );
  MUX2_X1 U14433 ( .A(n15384), .B(P3_REG2_REG_3__SCAN_IN), .S(n13255), .Z(
        n11998) );
  INV_X1 U14434 ( .A(n11998), .ZN(n12001) );
  NOR2_X1 U14435 ( .A1(n11999), .A2(n15353), .ZN(n15385) );
  AOI22_X1 U14436 ( .A1(n15336), .A2(n15385), .B1(n15369), .B2(n15440), .ZN(
        n12000) );
  OAI211_X1 U14437 ( .C1(n15383), .C2(n13214), .A(n12001), .B(n12000), .ZN(
        P3_U3230) );
  XNOR2_X1 U14438 ( .A(n15304), .B(n12640), .ZN(n12179) );
  XNOR2_X1 U14439 ( .A(n12179), .B(n15311), .ZN(n12013) );
  XNOR2_X1 U14440 ( .A(n12198), .B(n11571), .ZN(n12007) );
  XNOR2_X1 U14441 ( .A(n12007), .B(n15330), .ZN(n12195) );
  INV_X1 U14442 ( .A(n12006), .ZN(n12002) );
  NAND2_X1 U14443 ( .A1(n12003), .A2(n12002), .ZN(n12004) );
  NAND2_X1 U14444 ( .A1(n12006), .A2(n15331), .ZN(n12106) );
  OAI21_X1 U14445 ( .B1(n12195), .B2(n12106), .A(n12193), .ZN(n12009) );
  AOI22_X1 U14446 ( .A1(n12009), .A2(n12008), .B1(n12007), .B2(n15330), .ZN(
        n12010) );
  AOI21_X1 U14447 ( .B1(n12013), .B2(n12012), .A(n12181), .ZN(n12020) );
  INV_X1 U14448 ( .A(n14810), .ZN(n15299) );
  AOI21_X1 U14449 ( .B1(n15330), .B2(n15422), .A(n12014), .ZN(n12015) );
  OAI21_X1 U14450 ( .B1(n15299), .B2(n12891), .A(n12015), .ZN(n12017) );
  NOR2_X1 U14451 ( .A1(n12848), .A2(n15301), .ZN(n12016) );
  AOI211_X1 U14452 ( .C1(n15425), .C2(n12018), .A(n12017), .B(n12016), .ZN(
        n12019) );
  OAI21_X1 U14453 ( .B1(n12020), .B2(n15434), .A(n12019), .ZN(P3_U3171) );
  OAI222_X1 U14454 ( .A1(n14635), .A2(n12022), .B1(n14638), .B2(n12052), .C1(
        n12021), .C2(P1_U3086), .ZN(P1_U3334) );
  OR2_X1 U14455 ( .A1(n14870), .A2(n14101), .ZN(n12025) );
  NAND2_X1 U14456 ( .A1(n14892), .A2(n14100), .ZN(n12026) );
  AOI21_X1 U14457 ( .B1(n12032), .B2(n12027), .A(n6706), .ZN(n14782) );
  OR2_X1 U14458 ( .A1(n14870), .A2(n12321), .ZN(n12028) );
  AND2_X2 U14459 ( .A1(n12029), .A2(n12028), .ZN(n14883) );
  INV_X1 U14460 ( .A(n14100), .ZN(n12030) );
  OR2_X1 U14461 ( .A1(n14892), .A2(n12030), .ZN(n12031) );
  NOR2_X1 U14462 ( .A1(n12033), .A2(n12032), .ZN(n14778) );
  INV_X1 U14463 ( .A(n14394), .ZN(n14386) );
  NOR2_X1 U14464 ( .A1(n14778), .A2(n14386), .ZN(n12040) );
  NAND2_X1 U14465 ( .A1(n14781), .A2(n14894), .ZN(n12170) );
  OAI211_X1 U14466 ( .C1(n14781), .C2(n14894), .A(n11131), .B(n12170), .ZN(
        n14780) );
  NOR2_X1 U14467 ( .A1(n14498), .A2(n10036), .ZN(n12037) );
  NAND2_X1 U14468 ( .A1(n14100), .A2(n14479), .ZN(n12035) );
  NAND2_X1 U14469 ( .A1(n14098), .A2(n14477), .ZN(n12034) );
  AND2_X1 U14470 ( .A1(n12035), .A2(n12034), .ZN(n14779) );
  OAI22_X1 U14471 ( .A1(n6550), .A2(n14779), .B1(n12481), .B2(n15005), .ZN(
        n12036) );
  AOI211_X1 U14472 ( .C1(n12476), .C2(n14889), .A(n12037), .B(n12036), .ZN(
        n12038) );
  OAI21_X1 U14473 ( .B1(n14780), .B2(n14383), .A(n12038), .ZN(n12039) );
  AOI21_X1 U14474 ( .B1(n12040), .B2(n14785), .A(n12039), .ZN(n12041) );
  OAI21_X1 U14475 ( .B1(n14782), .B2(n14490), .A(n12041), .ZN(P1_U3281) );
  INV_X1 U14476 ( .A(n13832), .ZN(n13728) );
  AOI22_X1 U14477 ( .A1(n13734), .A2(n12043), .B1(n13825), .B2(n12042), .ZN(
        n12044) );
  OAI21_X1 U14478 ( .B1(n13724), .B2(n12045), .A(n12044), .ZN(n12046) );
  AOI21_X1 U14479 ( .B1(n13728), .B2(n12047), .A(n12046), .ZN(n12051) );
  MUX2_X1 U14480 ( .A(n12049), .B(n12048), .S(n13770), .Z(n12050) );
  NAND2_X1 U14481 ( .A1(n12051), .A2(n12050), .ZN(P2_U3262) );
  OAI222_X1 U14482 ( .A1(n13964), .A2(n12054), .B1(P2_U3088), .B2(n12053), 
        .C1(n12649), .C2(n12052), .ZN(P2_U3306) );
  XNOR2_X1 U14483 ( .A(n12055), .B(n12056), .ZN(n12062) );
  NAND2_X1 U14484 ( .A1(n13815), .A2(n13816), .ZN(n12058) );
  NAND2_X1 U14485 ( .A1(n13516), .A2(n13814), .ZN(n12057) );
  NAND2_X1 U14486 ( .A1(n12058), .A2(n12057), .ZN(n12230) );
  AOI22_X1 U14487 ( .A1(n14845), .A2(n12230), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12059) );
  OAI21_X1 U14488 ( .B1(n12233), .B2(n15124), .A(n12059), .ZN(n12060) );
  AOI21_X1 U14489 ( .B1(n12420), .B2(n13506), .A(n12060), .ZN(n12061) );
  OAI21_X1 U14490 ( .B1(n12062), .B2(n13481), .A(n12061), .ZN(P2_U3206) );
  INV_X2 U14491 ( .A(n13770), .ZN(n13812) );
  AOI21_X1 U14492 ( .B1(n12064), .B2(n13819), .A(n12063), .ZN(n15221) );
  INV_X1 U14493 ( .A(n12066), .ZN(n12067) );
  OAI211_X1 U14494 ( .C1(n15222), .C2(n8105), .A(n12067), .B(n13690), .ZN(
        n15220) );
  AOI22_X1 U14495 ( .A1(n13812), .A2(P2_REG2_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(n13825), .ZN(n12070) );
  NAND2_X1 U14496 ( .A1(n13734), .A2(n6553), .ZN(n12069) );
  OAI211_X1 U14497 ( .C1(n13724), .C2(n15220), .A(n12070), .B(n12069), .ZN(
        n12071) );
  AOI21_X1 U14498 ( .B1(n15218), .B2(n13728), .A(n12071), .ZN(n12072) );
  OAI21_X1 U14499 ( .B1(n13812), .B2(n15221), .A(n12072), .ZN(P2_U3264) );
  OR2_X1 U14500 ( .A1(n12074), .A2(n12073), .ZN(n12075) );
  NAND2_X1 U14501 ( .A1(n12076), .A2(n12075), .ZN(n15257) );
  OAI211_X1 U14502 ( .C1(n12079), .C2(n12078), .A(n12077), .B(n13819), .ZN(
        n12081) );
  NAND2_X1 U14503 ( .A1(n12081), .A2(n12080), .ZN(n15259) );
  NAND2_X1 U14504 ( .A1(n15259), .A2(n13770), .ZN(n12089) );
  OAI22_X1 U14505 ( .A1(n13770), .A2(n12083), .B1(n12082), .B2(n13784), .ZN(
        n12087) );
  AOI21_X1 U14506 ( .B1(n12084), .B2(n15252), .A(n8285), .ZN(n12085) );
  NAND2_X1 U14507 ( .A1(n12085), .A2(n12098), .ZN(n15254) );
  NOR2_X1 U14508 ( .A1(n15254), .A2(n13724), .ZN(n12086) );
  AOI211_X1 U14509 ( .C1(n13734), .C2(n15252), .A(n12087), .B(n12086), .ZN(
        n12088) );
  OAI211_X1 U14510 ( .C1(n13832), .C2(n15257), .A(n12089), .B(n12088), .ZN(
        P2_U3256) );
  XNOR2_X1 U14511 ( .A(n12090), .B(n12091), .ZN(n15267) );
  INV_X1 U14512 ( .A(n15267), .ZN(n12105) );
  XNOR2_X1 U14513 ( .A(n12092), .B(n12091), .ZN(n12095) );
  AOI22_X1 U14514 ( .A1(n13814), .A2(n13518), .B1(n15112), .B2(n13816), .ZN(
        n12094) );
  INV_X1 U14515 ( .A(n15256), .ZN(n13802) );
  NAND2_X1 U14516 ( .A1(n15267), .A2(n13802), .ZN(n12093) );
  OAI211_X1 U14517 ( .C1(n12095), .C2(n13799), .A(n12094), .B(n12093), .ZN(
        n15265) );
  NAND2_X1 U14518 ( .A1(n15265), .A2(n13770), .ZN(n12104) );
  OAI22_X1 U14519 ( .A1(n13770), .A2(n12097), .B1(n12096), .B2(n13784), .ZN(
        n12101) );
  INV_X1 U14520 ( .A(n12098), .ZN(n12099) );
  OAI211_X1 U14521 ( .C1(n15264), .C2(n12099), .A(n7494), .B(n13690), .ZN(
        n15262) );
  NOR2_X1 U14522 ( .A1(n15262), .A2(n13724), .ZN(n12100) );
  AOI211_X1 U14523 ( .C1(n13734), .C2(n12102), .A(n12101), .B(n12100), .ZN(
        n12103) );
  OAI211_X1 U14524 ( .C1(n12105), .C2(n13808), .A(n12104), .B(n12103), .ZN(
        P2_U3255) );
  NAND2_X1 U14525 ( .A1(n12107), .A2(n12106), .ZN(n12194) );
  XNOR2_X1 U14526 ( .A(n12194), .B(n12108), .ZN(n12117) );
  AOI21_X1 U14527 ( .B1(n15331), .B2(n15422), .A(n12109), .ZN(n12115) );
  INV_X1 U14528 ( .A(n15325), .ZN(n12110) );
  NAND2_X1 U14529 ( .A1(n15439), .A2(n12110), .ZN(n12114) );
  NAND2_X1 U14530 ( .A1(n15425), .A2(n12111), .ZN(n12113) );
  NAND2_X1 U14531 ( .A1(n15330), .A2(n15420), .ZN(n12112) );
  NAND4_X1 U14532 ( .A1(n12115), .A2(n12114), .A3(n12113), .A4(n12112), .ZN(
        n12116) );
  AOI21_X1 U14533 ( .B1(n12117), .B2(n12861), .A(n12116), .ZN(n12118) );
  INV_X1 U14534 ( .A(n12118), .ZN(P3_U3153) );
  OAI21_X1 U14535 ( .B1(n12120), .B2(n12123), .A(n12119), .ZN(n12128) );
  OAI22_X1 U14536 ( .A1(n12122), .A2(n13425), .B1(n12121), .B2(n13423), .ZN(
        n12127) );
  INV_X1 U14537 ( .A(n12123), .ZN(n12124) );
  XNOR2_X1 U14538 ( .A(n12125), .B(n12124), .ZN(n12217) );
  NOR2_X1 U14539 ( .A1(n12217), .A2(n15256), .ZN(n12126) );
  AOI211_X1 U14540 ( .C1(n13819), .C2(n12128), .A(n12127), .B(n12126), .ZN(
        n12216) );
  INV_X1 U14541 ( .A(n12129), .ZN(n12250) );
  AOI211_X1 U14542 ( .C1(n12214), .C2(n7494), .A(n8285), .B(n12250), .ZN(
        n12213) );
  AOI22_X1 U14543 ( .A1(n13812), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n12130), 
        .B2(n13825), .ZN(n12131) );
  OAI21_X1 U14544 ( .B1(n12132), .B2(n13828), .A(n12131), .ZN(n12134) );
  NOR2_X1 U14545 ( .A1(n12217), .A2(n13808), .ZN(n12133) );
  AOI211_X1 U14546 ( .C1(n12213), .C2(n13835), .A(n12134), .B(n12133), .ZN(
        n12135) );
  OAI21_X1 U14547 ( .B1(n12216), .B2(n13812), .A(n12135), .ZN(P2_U3254) );
  OAI22_X1 U14548 ( .A1(n13249), .A2(n12137), .B1(n12136), .B2(n15326), .ZN(
        n12140) );
  MUX2_X1 U14549 ( .A(n12138), .B(P3_REG2_REG_4__SCAN_IN), .S(n13255), .Z(
        n12139) );
  AOI211_X1 U14550 ( .C1(n15323), .C2(n12141), .A(n12140), .B(n12139), .ZN(
        n12142) );
  INV_X1 U14551 ( .A(n12142), .ZN(P3_U3229) );
  OAI22_X1 U14552 ( .A1(n13249), .A2(n12144), .B1(n12143), .B2(n15326), .ZN(
        n12147) );
  MUX2_X1 U14553 ( .A(n12145), .B(P3_REG2_REG_6__SCAN_IN), .S(n13255), .Z(
        n12146) );
  AOI211_X1 U14554 ( .C1(n15323), .C2(n12148), .A(n12147), .B(n12146), .ZN(
        n12149) );
  INV_X1 U14555 ( .A(n12149), .ZN(P3_U3227) );
  OAI21_X1 U14556 ( .B1(n12151), .B2(n14470), .A(n12150), .ZN(n12154) );
  NOR2_X1 U14557 ( .A1(n12163), .A2(n12152), .ZN(n12274) );
  AOI21_X1 U14558 ( .B1(n12152), .B2(n12163), .A(n12274), .ZN(n12153) );
  NAND2_X1 U14559 ( .A1(n12153), .A2(n12154), .ZN(n12275) );
  OAI211_X1 U14560 ( .C1(n12154), .C2(n12153), .A(n14232), .B(n12275), .ZN(
        n12162) );
  NAND2_X1 U14561 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14029)
         );
  AOI22_X1 U14562 ( .A1(n12157), .A2(n12156), .B1(P1_REG1_REG_16__SCAN_IN), 
        .B2(n12155), .ZN(n12277) );
  XNOR2_X1 U14563 ( .A(n12163), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n12279) );
  XNOR2_X1 U14564 ( .A(n12277), .B(n12279), .ZN(n12158) );
  NAND2_X1 U14565 ( .A1(n14233), .A2(n12158), .ZN(n12159) );
  NAND2_X1 U14566 ( .A1(n14029), .A2(n12159), .ZN(n12160) );
  AOI21_X1 U14567 ( .B1(n14212), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n12160), 
        .ZN(n12161) );
  OAI211_X1 U14568 ( .C1(n14976), .C2(n12163), .A(n12162), .B(n12161), .ZN(
        P1_U3260) );
  INV_X1 U14569 ( .A(n14099), .ZN(n12474) );
  OR2_X1 U14570 ( .A1(n12476), .A2(n12474), .ZN(n12165) );
  NAND3_X1 U14571 ( .A1(n14785), .A2(n7712), .A3(n12165), .ZN(n12166) );
  NAND3_X1 U14572 ( .A1(n12258), .A2(n15052), .A3(n12166), .ZN(n12168) );
  OAI22_X1 U14573 ( .A1(n12670), .A2(n14464), .B1(n12474), .B2(n14462), .ZN(
        n12494) );
  INV_X1 U14574 ( .A(n12494), .ZN(n12167) );
  NAND2_X1 U14575 ( .A1(n12168), .A2(n12167), .ZN(n12223) );
  INV_X1 U14576 ( .A(n12223), .ZN(n12178) );
  NAND2_X1 U14577 ( .A1(n12169), .A2(n7712), .ZN(n12264) );
  OAI21_X1 U14578 ( .B1(n12169), .B2(n7712), .A(n12264), .ZN(n12225) );
  INV_X1 U14579 ( .A(n12170), .ZN(n12171) );
  OR2_X2 U14580 ( .A1(n12170), .A2(n12499), .ZN(n12268) );
  OAI211_X1 U14581 ( .C1(n12171), .C2(n12492), .A(n11131), .B(n12268), .ZN(
        n12222) );
  INV_X1 U14582 ( .A(n12172), .ZN(n12497) );
  OAI22_X1 U14583 ( .A1(n14498), .A2(n12173), .B1(n12497), .B2(n15005), .ZN(
        n12174) );
  AOI21_X1 U14584 ( .B1(n12499), .B2(n14889), .A(n12174), .ZN(n12175) );
  OAI21_X1 U14585 ( .B1(n12222), .B2(n14383), .A(n12175), .ZN(n12176) );
  AOI21_X1 U14586 ( .B1(n12225), .B2(n14898), .A(n12176), .ZN(n12177) );
  OAI21_X1 U14587 ( .B1(n12178), .B2(n6550), .A(n12177), .ZN(P1_U3280) );
  XNOR2_X1 U14588 ( .A(n15287), .B(n12640), .ZN(n12327) );
  XNOR2_X1 U14589 ( .A(n12327), .B(n14810), .ZN(n12183) );
  NOR2_X1 U14590 ( .A1(n12179), .A2(n15311), .ZN(n12180) );
  OR2_X1 U14591 ( .A1(n12181), .A2(n12180), .ZN(n12182) );
  AOI211_X1 U14592 ( .C1(n12183), .C2(n12182), .A(n15434), .B(n12330), .ZN(
        n12192) );
  AOI21_X1 U14593 ( .B1(n15311), .B2(n15422), .A(n12184), .ZN(n12190) );
  NAND2_X1 U14594 ( .A1(n15425), .A2(n12185), .ZN(n12189) );
  INV_X1 U14595 ( .A(n15288), .ZN(n12186) );
  NAND2_X1 U14596 ( .A1(n15439), .A2(n12186), .ZN(n12188) );
  NAND2_X1 U14597 ( .A1(n15282), .A2(n15420), .ZN(n12187) );
  NAND4_X1 U14598 ( .A1(n12190), .A2(n12189), .A3(n12188), .A4(n12187), .ZN(
        n12191) );
  OR2_X1 U14599 ( .A1(n12192), .A2(n12191), .ZN(P3_U3157) );
  MUX2_X1 U14600 ( .A(n15310), .B(n12194), .S(n12193), .Z(n12196) );
  XNOR2_X1 U14601 ( .A(n12196), .B(n12195), .ZN(n12204) );
  AOI21_X1 U14602 ( .B1(n15310), .B2(n15422), .A(n12197), .ZN(n12202) );
  NAND2_X1 U14603 ( .A1(n15439), .A2(n15313), .ZN(n12201) );
  NAND2_X1 U14604 ( .A1(n15425), .A2(n12198), .ZN(n12200) );
  NAND2_X1 U14605 ( .A1(n15311), .A2(n15420), .ZN(n12199) );
  NAND4_X1 U14606 ( .A1(n12202), .A2(n12201), .A3(n12200), .A4(n12199), .ZN(
        n12203) );
  AOI21_X1 U14607 ( .B1(n12204), .B2(n12861), .A(n12203), .ZN(n12205) );
  INV_X1 U14608 ( .A(n12205), .ZN(P3_U3161) );
  INV_X1 U14609 ( .A(n12206), .ZN(n12208) );
  OAI222_X1 U14610 ( .A1(n12209), .A2(P3_U3151), .B1(n14743), .B2(n12208), 
        .C1(n12207), .C2(n14741), .ZN(P3_U3271) );
  OAI222_X1 U14611 ( .A1(n13964), .A2(n12212), .B1(P2_U3088), .B2(n12211), 
        .C1(n12649), .C2(n12210), .ZN(P2_U3305) );
  AOI21_X1 U14612 ( .B1(n15251), .B2(n12214), .A(n12213), .ZN(n12215) );
  OAI211_X1 U14613 ( .C1(n12217), .C2(n15255), .A(n12216), .B(n12215), .ZN(
        n12219) );
  NAND2_X1 U14614 ( .A1(n12219), .A2(n15279), .ZN(n12218) );
  OAI21_X1 U14615 ( .B1(n15279), .B2(n11041), .A(n12218), .ZN(P2_U3510) );
  INV_X1 U14616 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n12221) );
  NAND2_X1 U14617 ( .A1(n12219), .A2(n15270), .ZN(n12220) );
  OAI21_X1 U14618 ( .B1(n15270), .B2(n12221), .A(n12220), .ZN(P2_U3463) );
  OAI21_X1 U14619 ( .B1(n12492), .B2(n14902), .A(n12222), .ZN(n12224) );
  AOI211_X1 U14620 ( .C1(n15093), .C2(n12225), .A(n12224), .B(n12223), .ZN(
        n12228) );
  NAND2_X1 U14621 ( .A1(n7451), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n12226) );
  OAI21_X1 U14622 ( .B1(n12228), .B2(n7451), .A(n12226), .ZN(P1_U3498) );
  NAND2_X1 U14623 ( .A1(n15105), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n12227) );
  OAI21_X1 U14624 ( .B1(n12228), .B2(n15105), .A(n12227), .ZN(P1_U3541) );
  XNOR2_X1 U14625 ( .A(n12229), .B(n12237), .ZN(n12231) );
  AOI21_X1 U14626 ( .B1(n12231), .B2(n13819), .A(n12230), .ZN(n12422) );
  INV_X1 U14627 ( .A(n12445), .ZN(n12232) );
  AOI211_X1 U14628 ( .C1(n12420), .C2(n12249), .A(n8285), .B(n12232), .ZN(
        n12419) );
  INV_X1 U14629 ( .A(n12233), .ZN(n12234) );
  AOI22_X1 U14630 ( .A1(n13812), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n12234), 
        .B2(n13825), .ZN(n12235) );
  OAI21_X1 U14631 ( .B1(n12236), .B2(n13828), .A(n12235), .ZN(n12241) );
  INV_X1 U14632 ( .A(n12237), .ZN(n12238) );
  XNOR2_X1 U14633 ( .A(n12239), .B(n12238), .ZN(n12423) );
  NOR2_X1 U14634 ( .A1(n12423), .A2(n13832), .ZN(n12240) );
  AOI211_X1 U14635 ( .C1(n12419), .C2(n13835), .A(n12241), .B(n12240), .ZN(
        n12242) );
  OAI21_X1 U14636 ( .B1(n12422), .B2(n13812), .A(n12242), .ZN(P2_U3252) );
  XOR2_X1 U14637 ( .A(n12245), .B(n12243), .Z(n14851) );
  AOI211_X1 U14638 ( .C1(n12245), .C2(n12244), .A(n13799), .B(n6715), .ZN(
        n12246) );
  INV_X1 U14639 ( .A(n12246), .ZN(n12248) );
  AOI22_X1 U14640 ( .A1(n13814), .A2(n15112), .B1(n15114), .B2(n13816), .ZN(
        n12247) );
  OAI211_X1 U14641 ( .C1(n14851), .C2(n15256), .A(n12248), .B(n12247), .ZN(
        n14853) );
  NAND2_X1 U14642 ( .A1(n14853), .A2(n13770), .ZN(n12255) );
  OAI22_X1 U14643 ( .A1(n13770), .A2(n13550), .B1(n15123), .B2(n13784), .ZN(
        n12252) );
  OAI211_X1 U14644 ( .C1(n12250), .C2(n15118), .A(n13690), .B(n12249), .ZN(
        n14852) );
  NOR2_X1 U14645 ( .A1(n14852), .A2(n13724), .ZN(n12251) );
  AOI211_X1 U14646 ( .C1(n13734), .C2(n12253), .A(n12252), .B(n12251), .ZN(
        n12254) );
  OAI211_X1 U14647 ( .C1(n14851), .C2(n13808), .A(n12255), .B(n12254), .ZN(
        P2_U3253) );
  INV_X1 U14648 ( .A(n14869), .ZN(n12262) );
  AND2_X1 U14649 ( .A1(n14098), .A2(n14479), .ZN(n12256) );
  AOI21_X1 U14650 ( .B1(n14097), .B2(n14477), .A(n12256), .ZN(n14861) );
  INV_X1 U14651 ( .A(n14861), .ZN(n12261) );
  OR2_X1 U14652 ( .A1(n12499), .A2(n12491), .ZN(n12257) );
  NAND2_X1 U14653 ( .A1(n12258), .A2(n12257), .ZN(n12549) );
  XNOR2_X1 U14654 ( .A(n12549), .B(n7583), .ZN(n12260) );
  NOR2_X1 U14655 ( .A1(n12260), .A2(n15002), .ZN(n12375) );
  AOI211_X1 U14656 ( .C1(n14888), .C2(n12262), .A(n12261), .B(n12375), .ZN(
        n12273) );
  OR2_X1 U14657 ( .A1(n12499), .A2(n14098), .ZN(n12263) );
  INV_X1 U14658 ( .A(n12576), .ZN(n12266) );
  AOI21_X1 U14659 ( .B1(n7583), .B2(n12267), .A(n12266), .ZN(n12377) );
  INV_X1 U14660 ( .A(n12672), .ZN(n14863) );
  INV_X1 U14661 ( .A(n12268), .ZN(n12269) );
  OR2_X2 U14662 ( .A1(n12672), .A2(n12268), .ZN(n14484) );
  OAI211_X1 U14663 ( .C1(n14863), .C2(n12269), .A(n11131), .B(n14484), .ZN(
        n12374) );
  AOI22_X1 U14664 ( .A1(n12672), .A2(n14889), .B1(P1_REG2_REG_14__SCAN_IN), 
        .B2(n6550), .ZN(n12270) );
  OAI21_X1 U14665 ( .B1(n12374), .B2(n14383), .A(n12270), .ZN(n12271) );
  AOI21_X1 U14666 ( .B1(n12377), .B2(n14898), .A(n12271), .ZN(n12272) );
  OAI21_X1 U14667 ( .B1(n12273), .B2(n6550), .A(n12272), .ZN(P1_U3279) );
  INV_X1 U14668 ( .A(n12274), .ZN(n12276) );
  NAND2_X1 U14669 ( .A1(n12276), .A2(n12275), .ZN(n14223) );
  XNOR2_X1 U14670 ( .A(n14223), .B(n14222), .ZN(n14225) );
  XOR2_X1 U14671 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n14225), .Z(n12286) );
  NAND2_X1 U14672 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14065)
         );
  INV_X1 U14673 ( .A(n12277), .ZN(n12280) );
  AOI22_X1 U14674 ( .A1(n12280), .A2(n12279), .B1(P1_REG1_REG_17__SCAN_IN), 
        .B2(n12278), .ZN(n14217) );
  XNOR2_X1 U14675 ( .A(n14217), .B(n14222), .ZN(n12281) );
  NAND2_X1 U14676 ( .A1(n12281), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n14220) );
  OAI211_X1 U14677 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n12281), .A(n14233), 
        .B(n14220), .ZN(n12282) );
  NAND2_X1 U14678 ( .A1(n14065), .A2(n12282), .ZN(n12283) );
  AOI21_X1 U14679 ( .B1(n14212), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n12283), 
        .ZN(n12285) );
  NAND2_X1 U14680 ( .A1(n14206), .A2(n14222), .ZN(n12284) );
  OAI211_X1 U14681 ( .C1(n12286), .C2(n14972), .A(n12285), .B(n12284), .ZN(
        P1_U3261) );
  INV_X1 U14682 ( .A(n12287), .ZN(n12290) );
  INV_X1 U14683 ( .A(n12288), .ZN(n12289) );
  NAND2_X1 U14684 ( .A1(n12290), .A2(n12289), .ZN(n12291) );
  NAND2_X1 U14685 ( .A1(n14943), .A2(n12753), .ZN(n12294) );
  NAND2_X1 U14686 ( .A1(n12743), .A2(n14103), .ZN(n12293) );
  NAND2_X1 U14687 ( .A1(n12294), .A2(n12293), .ZN(n12295) );
  XNOR2_X1 U14688 ( .A(n12295), .B(n12777), .ZN(n12298) );
  NOR2_X1 U14689 ( .A1(n12776), .A2(n12296), .ZN(n12297) );
  AOI21_X1 U14690 ( .B1(n14943), .B2(n12743), .A(n12297), .ZN(n12299) );
  XNOR2_X1 U14691 ( .A(n12298), .B(n12299), .ZN(n14946) );
  INV_X1 U14692 ( .A(n12298), .ZN(n12300) );
  NAND2_X1 U14693 ( .A1(n12300), .A2(n12299), .ZN(n12301) );
  NOR2_X1 U14694 ( .A1(n12776), .A2(n12302), .ZN(n12303) );
  AOI21_X1 U14695 ( .B1(n14952), .B2(n12743), .A(n12303), .ZN(n12307) );
  NOR2_X1 U14696 ( .A1(n12308), .A2(n12307), .ZN(n14954) );
  NAND2_X1 U14697 ( .A1(n14952), .A2(n12753), .ZN(n12305) );
  NAND2_X1 U14698 ( .A1(n12743), .A2(n14102), .ZN(n12304) );
  NAND2_X1 U14699 ( .A1(n12305), .A2(n12304), .ZN(n12306) );
  XNOR2_X1 U14700 ( .A(n12306), .B(n12777), .ZN(n14957) );
  NAND2_X1 U14701 ( .A1(n12308), .A2(n12307), .ZN(n14955) );
  NAND2_X1 U14702 ( .A1(n14870), .A2(n12753), .ZN(n12310) );
  NAND2_X1 U14703 ( .A1(n12743), .A2(n14101), .ZN(n12309) );
  NAND2_X1 U14704 ( .A1(n12310), .A2(n12309), .ZN(n12311) );
  XNOR2_X1 U14705 ( .A(n12311), .B(n12777), .ZN(n12315) );
  NAND2_X1 U14706 ( .A1(n14870), .A2(n12743), .ZN(n12313) );
  NAND2_X1 U14707 ( .A1(n12770), .A2(n14101), .ZN(n12312) );
  NAND2_X1 U14708 ( .A1(n12313), .A2(n12312), .ZN(n12314) );
  NAND2_X1 U14709 ( .A1(n12315), .A2(n12314), .ZN(n14873) );
  NOR2_X1 U14710 ( .A1(n12315), .A2(n12314), .ZN(n14874) );
  AOI22_X1 U14711 ( .A1(n14892), .A2(n12743), .B1(n12770), .B2(n14100), .ZN(
        n12468) );
  NAND2_X1 U14712 ( .A1(n14892), .A2(n12753), .ZN(n12317) );
  NAND2_X1 U14713 ( .A1(n12743), .A2(n14100), .ZN(n12316) );
  NAND2_X1 U14714 ( .A1(n12317), .A2(n12316), .ZN(n12318) );
  XNOR2_X1 U14715 ( .A(n12318), .B(n12777), .ZN(n12470) );
  XOR2_X1 U14716 ( .A(n12468), .B(n12470), .Z(n12319) );
  AOI21_X1 U14717 ( .B1(n12320), .B2(n12319), .A(n12479), .ZN(n12326) );
  OAI22_X1 U14718 ( .A1(n12321), .A2(n14462), .B1(n12474), .B2(n14464), .ZN(
        n14884) );
  NAND2_X1 U14719 ( .A1(n14960), .A2(n14884), .ZN(n12322) );
  OAI211_X1 U14720 ( .C1(n14965), .C2(n14886), .A(n12323), .B(n12322), .ZN(
        n12324) );
  AOI21_X1 U14721 ( .B1(n14892), .B2(n14090), .A(n12324), .ZN(n12325) );
  OAI21_X1 U14722 ( .B1(n12326), .B2(n14935), .A(n12325), .ZN(P1_U3236) );
  INV_X1 U14723 ( .A(n12327), .ZN(n12328) );
  NOR2_X1 U14724 ( .A1(n15299), .A2(n12328), .ZN(n12329) );
  XNOR2_X1 U14725 ( .A(n12334), .B(n12640), .ZN(n12331) );
  NAND2_X1 U14726 ( .A1(n12332), .A2(n12331), .ZN(n12406) );
  NAND2_X1 U14727 ( .A1(n7101), .A2(n12406), .ZN(n12333) );
  XNOR2_X1 U14728 ( .A(n12333), .B(n15282), .ZN(n12341) );
  AND2_X1 U14729 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n12352) );
  AOI21_X1 U14730 ( .B1(n14810), .B2(n15422), .A(n12352), .ZN(n12339) );
  NAND2_X1 U14731 ( .A1(n12334), .A2(n15425), .ZN(n12338) );
  INV_X1 U14732 ( .A(n12335), .ZN(n14813) );
  NAND2_X1 U14733 ( .A1(n15439), .A2(n14813), .ZN(n12337) );
  NAND2_X1 U14734 ( .A1(n14809), .A2(n15420), .ZN(n12336) );
  NAND4_X1 U14735 ( .A1(n12339), .A2(n12338), .A3(n12337), .A4(n12336), .ZN(
        n12340) );
  AOI21_X1 U14736 ( .B1(n12341), .B2(n12861), .A(n12340), .ZN(n12342) );
  INV_X1 U14737 ( .A(n12342), .ZN(P3_U3176) );
  INV_X1 U14738 ( .A(n12343), .ZN(n12345) );
  OAI222_X1 U14739 ( .A1(P3_U3151), .A2(n12346), .B1(n14743), .B2(n12345), 
        .C1(n12344), .C2(n14741), .ZN(P3_U3270) );
  AOI21_X1 U14740 ( .B1(n12347), .B2(n8819), .A(n12395), .ZN(n12360) );
  INV_X1 U14741 ( .A(n12348), .ZN(n12350) );
  MUX2_X1 U14742 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12946), .Z(n12387) );
  XNOR2_X1 U14743 ( .A(n12387), .B(n14760), .ZN(n12388) );
  XNOR2_X1 U14744 ( .A(n12389), .B(n12388), .ZN(n12358) );
  AOI21_X1 U14745 ( .B1(n15280), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n12352), 
        .ZN(n12353) );
  OAI21_X1 U14746 ( .B1(n12935), .B2(n14760), .A(n12353), .ZN(n12357) );
  AOI21_X1 U14747 ( .B1(n8816), .B2(n12354), .A(n12382), .ZN(n12355) );
  NOR2_X1 U14748 ( .A1(n12355), .A2(n13004), .ZN(n12356) );
  AOI211_X1 U14749 ( .C1(n12358), .C2(n12916), .A(n12357), .B(n12356), .ZN(
        n12359) );
  OAI21_X1 U14750 ( .B1(n12360), .B2(n13040), .A(n12359), .ZN(P3_U3193) );
  XNOR2_X1 U14751 ( .A(n12361), .B(n12367), .ZN(n12364) );
  NAND2_X1 U14752 ( .A1(n15282), .A2(n15360), .ZN(n12362) );
  OAI21_X1 U14753 ( .B1(n12428), .B2(n15300), .A(n12362), .ZN(n12363) );
  AOI21_X1 U14754 ( .B1(n12364), .B2(n10380), .A(n12363), .ZN(n14829) );
  NOR2_X1 U14755 ( .A1(n12409), .A2(n15353), .ZN(n14826) );
  OAI22_X1 U14756 ( .A1(n15372), .A2(n12365), .B1(n12411), .B2(n15326), .ZN(
        n12366) );
  AOI21_X1 U14757 ( .B1(n14826), .B2(n15336), .A(n12366), .ZN(n12370) );
  XNOR2_X1 U14758 ( .A(n12368), .B(n12367), .ZN(n14827) );
  NAND2_X1 U14759 ( .A1(n14827), .A2(n15323), .ZN(n12369) );
  OAI211_X1 U14760 ( .C1(n14829), .C2(n13255), .A(n12370), .B(n12369), .ZN(
        P3_U3221) );
  INV_X1 U14761 ( .A(n12402), .ZN(n12373) );
  NAND2_X1 U14762 ( .A1(n14620), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12371) );
  OAI211_X1 U14763 ( .C1(n12373), .C2(n14638), .A(n12372), .B(n12371), .ZN(
        P1_U3332) );
  OAI211_X1 U14764 ( .C1(n14863), .C2(n14902), .A(n12374), .B(n14861), .ZN(
        n12376) );
  AOI211_X1 U14765 ( .C1(n12377), .C2(n15093), .A(n12376), .B(n12375), .ZN(
        n12380) );
  NAND2_X1 U14766 ( .A1(n7451), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n12378) );
  OAI21_X1 U14767 ( .B1(n12380), .B2(n7451), .A(n12378), .ZN(P1_U3501) );
  NAND2_X1 U14768 ( .A1(n15105), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n12379) );
  OAI21_X1 U14769 ( .B1(n12380), .B2(n15105), .A(n12379), .ZN(P1_U3542) );
  AOI22_X1 U14770 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n12396), .B1(n14765), 
        .B2(n8840), .ZN(n12383) );
  AOI21_X1 U14771 ( .B1(n12384), .B2(n12383), .A(n12910), .ZN(n12401) );
  NOR2_X1 U14772 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12385), .ZN(n12410) );
  INV_X1 U14773 ( .A(n12410), .ZN(n12386) );
  OAI21_X1 U14774 ( .B1(n13012), .B2(n15455), .A(n12386), .ZN(n12393) );
  MUX2_X1 U14775 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12946), .Z(n12905) );
  XNOR2_X1 U14776 ( .A(n12905), .B(n14765), .ZN(n12391) );
  NOR2_X1 U14777 ( .A1(n12390), .A2(n12391), .ZN(n12904) );
  AOI211_X1 U14778 ( .C1(n12391), .C2(n12390), .A(n13051), .B(n12904), .ZN(
        n12392) );
  AOI211_X1 U14779 ( .C1(n13041), .C2(n12396), .A(n12393), .B(n12392), .ZN(
        n12400) );
  AOI22_X1 U14780 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n12396), .B1(n14765), 
        .B2(n12365), .ZN(n12397) );
  OR2_X1 U14781 ( .A1(n6718), .A2(n13040), .ZN(n12399) );
  OAI211_X1 U14782 ( .C1(n12401), .C2(n13004), .A(n12400), .B(n12399), .ZN(
        P3_U3194) );
  NAND2_X1 U14783 ( .A1(n12402), .A2(n13951), .ZN(n12404) );
  OAI211_X1 U14784 ( .C1(n15676), .C2(n13964), .A(n12404), .B(n12403), .ZN(
        P2_U3304) );
  XNOR2_X1 U14785 ( .A(n12409), .B(n12640), .ZN(n12405) );
  NOR2_X1 U14786 ( .A1(n12405), .A2(n14809), .ZN(n12425) );
  AOI21_X1 U14787 ( .B1(n12405), .B2(n14809), .A(n12425), .ZN(n12408) );
  NAND2_X1 U14788 ( .A1(n12407), .A2(n12408), .ZN(n12427) );
  OAI21_X1 U14789 ( .B1(n12408), .B2(n12407), .A(n12427), .ZN(n12417) );
  NOR2_X1 U14790 ( .A1(n12409), .A2(n12882), .ZN(n12416) );
  AOI21_X1 U14791 ( .B1(n15282), .B2(n15422), .A(n12410), .ZN(n12414) );
  INV_X1 U14792 ( .A(n12411), .ZN(n12412) );
  NAND2_X1 U14793 ( .A1(n15439), .A2(n12412), .ZN(n12413) );
  OAI211_X1 U14794 ( .C1(n12428), .C2(n12891), .A(n12414), .B(n12413), .ZN(
        n12415) );
  AOI211_X1 U14795 ( .C1(n12417), .C2(n12861), .A(n12416), .B(n12415), .ZN(
        n12418) );
  INV_X1 U14796 ( .A(n12418), .ZN(P3_U3164) );
  AOI21_X1 U14797 ( .B1(n15251), .B2(n12420), .A(n12419), .ZN(n12421) );
  OAI211_X1 U14798 ( .C1(n15249), .C2(n12423), .A(n12422), .B(n12421), .ZN(
        n12439) );
  NAND2_X1 U14799 ( .A1(n12439), .A2(n15279), .ZN(n12424) );
  OAI21_X1 U14800 ( .B1(n15279), .B2(n13565), .A(n12424), .ZN(P2_U3512) );
  INV_X1 U14801 ( .A(n12425), .ZN(n12426) );
  XNOR2_X1 U14802 ( .A(n14821), .B(n11571), .ZN(n12429) );
  AND2_X1 U14803 ( .A1(n12429), .A2(n12428), .ZN(n12506) );
  INV_X1 U14804 ( .A(n12506), .ZN(n12431) );
  INV_X1 U14805 ( .A(n12429), .ZN(n12430) );
  NAND2_X1 U14806 ( .A1(n12430), .A2(n12901), .ZN(n12505) );
  NAND2_X1 U14807 ( .A1(n12431), .A2(n12505), .ZN(n12432) );
  XNOR2_X1 U14808 ( .A(n12507), .B(n12432), .ZN(n12438) );
  INV_X1 U14809 ( .A(n14821), .ZN(n12436) );
  AND2_X1 U14810 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n12908) );
  NOR2_X1 U14811 ( .A1(n13244), .A2(n12891), .ZN(n12433) );
  AOI211_X1 U14812 ( .C1(n15422), .C2(n14809), .A(n12908), .B(n12433), .ZN(
        n12434) );
  OAI21_X1 U14813 ( .B1(n12464), .B2(n12848), .A(n12434), .ZN(n12435) );
  AOI21_X1 U14814 ( .B1(n12436), .B2(n15425), .A(n12435), .ZN(n12437) );
  OAI21_X1 U14815 ( .B1(n12438), .B2(n15434), .A(n12437), .ZN(P3_U3174) );
  INV_X1 U14816 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n15622) );
  NAND2_X1 U14817 ( .A1(n12439), .A2(n15270), .ZN(n12440) );
  OAI21_X1 U14818 ( .B1(n15270), .B2(n15622), .A(n12440), .ZN(P2_U3469) );
  XNOR2_X1 U14819 ( .A(n12441), .B(n12449), .ZN(n12444) );
  OAI22_X1 U14820 ( .A1(n12443), .A2(n13425), .B1(n12442), .B2(n13423), .ZN(
        n14846) );
  AOI21_X1 U14821 ( .B1(n12444), .B2(n13819), .A(n14846), .ZN(n13918) );
  AOI211_X1 U14822 ( .C1(n14847), .C2(n12445), .A(n8285), .B(n7496), .ZN(
        n13916) );
  INV_X1 U14823 ( .A(n14847), .ZN(n12448) );
  INV_X1 U14824 ( .A(n14850), .ZN(n12446) );
  AOI22_X1 U14825 ( .A1(n13812), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n12446), 
        .B2(n13825), .ZN(n12447) );
  OAI21_X1 U14826 ( .B1(n12448), .B2(n13828), .A(n12447), .ZN(n12452) );
  XNOR2_X1 U14827 ( .A(n12450), .B(n12449), .ZN(n13919) );
  NOR2_X1 U14828 ( .A1(n13919), .A2(n13832), .ZN(n12451) );
  AOI211_X1 U14829 ( .C1(n13916), .C2(n13835), .A(n12452), .B(n12451), .ZN(
        n12453) );
  OAI21_X1 U14830 ( .B1(n13918), .B2(n13812), .A(n12453), .ZN(P2_U3251) );
  INV_X1 U14831 ( .A(n12454), .ZN(n12456) );
  OAI222_X1 U14832 ( .A1(n12457), .A2(P3_U3151), .B1(n14743), .B2(n12456), 
        .C1(n12455), .C2(n14741), .ZN(P3_U3269) );
  XNOR2_X1 U14833 ( .A(n12458), .B(n12462), .ZN(n12459) );
  NAND2_X1 U14834 ( .A1(n12459), .A2(n10380), .ZN(n12461) );
  AOI22_X1 U14835 ( .A1(n15360), .A2(n14809), .B1(n12900), .B2(n15358), .ZN(
        n12460) );
  XNOR2_X1 U14836 ( .A(n12463), .B(n12462), .ZN(n14823) );
  NOR2_X1 U14837 ( .A1(n14821), .A2(n13249), .ZN(n12466) );
  OAI22_X1 U14838 ( .A1(n15372), .A2(n8862), .B1(n12464), .B2(n15326), .ZN(
        n12465) );
  AOI211_X1 U14839 ( .C1(n14823), .C2(n15323), .A(n12466), .B(n12465), .ZN(
        n12467) );
  OAI21_X1 U14840 ( .B1(n14825), .B2(n13255), .A(n12467), .ZN(P3_U3220) );
  INV_X1 U14841 ( .A(n12468), .ZN(n12469) );
  NOR2_X1 U14842 ( .A1(n12470), .A2(n12469), .ZN(n12478) );
  NAND2_X1 U14843 ( .A1(n12476), .A2(n12753), .ZN(n12472) );
  NAND2_X1 U14844 ( .A1(n12743), .A2(n14099), .ZN(n12471) );
  NAND2_X1 U14845 ( .A1(n12472), .A2(n12471), .ZN(n12473) );
  XNOR2_X1 U14846 ( .A(n12473), .B(n12746), .ZN(n12487) );
  NOR2_X1 U14847 ( .A1(n12776), .A2(n12474), .ZN(n12475) );
  AOI21_X1 U14848 ( .B1(n12476), .B2(n12743), .A(n12475), .ZN(n12486) );
  XNOR2_X1 U14849 ( .A(n12487), .B(n12486), .ZN(n12477) );
  OAI21_X1 U14850 ( .B1(n12479), .B2(n12478), .A(n12477), .ZN(n12480) );
  NAND3_X1 U14851 ( .A1(n6724), .A2(n14961), .A3(n12480), .ZN(n12485) );
  INV_X1 U14852 ( .A(n12481), .ZN(n12483) );
  OAI22_X1 U14853 ( .A1(n14862), .A2(n14779), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10037), .ZN(n12482) );
  AOI21_X1 U14854 ( .B1(n14068), .B2(n12483), .A(n12482), .ZN(n12484) );
  OAI211_X1 U14855 ( .C1(n14781), .C2(n14864), .A(n12485), .B(n12484), .ZN(
        P1_U3224) );
  INV_X1 U14856 ( .A(n12486), .ZN(n12489) );
  INV_X1 U14857 ( .A(n12487), .ZN(n12488) );
  NOR2_X1 U14858 ( .A1(n12776), .A2(n12491), .ZN(n12490) );
  AOI21_X1 U14859 ( .B1(n12499), .B2(n12743), .A(n12490), .ZN(n12664) );
  OAI22_X1 U14860 ( .A1(n12492), .A2(n11135), .B1(n12491), .B2(n12779), .ZN(
        n12493) );
  XNOR2_X1 U14861 ( .A(n12493), .B(n12777), .ZN(n12662) );
  XOR2_X1 U14862 ( .A(n12664), .B(n12662), .Z(n12665) );
  XNOR2_X1 U14863 ( .A(n12666), .B(n12665), .ZN(n12501) );
  NAND2_X1 U14864 ( .A1(n14960), .A2(n12494), .ZN(n12495) );
  OAI211_X1 U14865 ( .C1(n14965), .C2(n12497), .A(n12496), .B(n12495), .ZN(
        n12498) );
  AOI21_X1 U14866 ( .B1(n12499), .B2(n14090), .A(n12498), .ZN(n12500) );
  OAI21_X1 U14867 ( .B1(n12501), .B2(n14935), .A(n12500), .ZN(P1_U3234) );
  INV_X1 U14868 ( .A(n12502), .ZN(n12504) );
  OAI222_X1 U14869 ( .A1(P3_U3151), .A2(n12946), .B1(n14743), .B2(n12504), 
        .C1(n12503), .C2(n14741), .ZN(P3_U3268) );
  XNOR2_X1 U14870 ( .A(n13375), .B(n12640), .ZN(n12516) );
  XNOR2_X1 U14871 ( .A(n12516), .B(n13244), .ZN(n12508) );
  OAI211_X1 U14872 ( .C1(n12509), .C2(n12508), .A(n12518), .B(n12861), .ZN(
        n12515) );
  INV_X1 U14873 ( .A(n12530), .ZN(n12513) );
  INV_X1 U14874 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n12510) );
  NOR2_X1 U14875 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12510), .ZN(n12933) );
  AOI21_X1 U14876 ( .B1(n12901), .B2(n15422), .A(n12933), .ZN(n12511) );
  OAI21_X1 U14877 ( .B1(n13231), .B2(n12891), .A(n12511), .ZN(n12512) );
  AOI21_X1 U14878 ( .B1(n12513), .B2(n15439), .A(n12512), .ZN(n12514) );
  OAI211_X1 U14879 ( .C1(n12882), .C2(n13375), .A(n12515), .B(n12514), .ZN(
        P3_U3155) );
  NAND2_X1 U14880 ( .A1(n12516), .A2(n12900), .ZN(n12517) );
  XNOR2_X1 U14881 ( .A(n12610), .B(n13231), .ZN(n12519) );
  XNOR2_X1 U14882 ( .A(n12611), .B(n12519), .ZN(n12524) );
  AND2_X1 U14883 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12943) );
  NOR2_X1 U14884 ( .A1(n13245), .A2(n12891), .ZN(n12520) );
  AOI211_X1 U14885 ( .C1(n15422), .C2(n12900), .A(n12943), .B(n12520), .ZN(
        n12521) );
  OAI21_X1 U14886 ( .B1(n13250), .B2(n12848), .A(n12521), .ZN(n12522) );
  AOI21_X1 U14887 ( .B1(n15425), .B2(n13248), .A(n12522), .ZN(n12523) );
  OAI21_X1 U14888 ( .B1(n12524), .B2(n15434), .A(n12523), .ZN(P3_U3181) );
  XNOR2_X1 U14889 ( .A(n12525), .B(n12527), .ZN(n13314) );
  INV_X1 U14890 ( .A(n13314), .ZN(n12535) );
  OAI211_X1 U14891 ( .C1(n6712), .C2(n12527), .A(n10380), .B(n12526), .ZN(
        n12529) );
  AOI22_X1 U14892 ( .A1(n12901), .A2(n15360), .B1(n15358), .B2(n12899), .ZN(
        n12528) );
  NAND2_X1 U14893 ( .A1(n12529), .A2(n12528), .ZN(n13313) );
  NOR2_X1 U14894 ( .A1(n13375), .A2(n13249), .ZN(n12533) );
  INV_X1 U14895 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12531) );
  OAI22_X1 U14896 ( .A1(n15372), .A2(n12531), .B1(n12530), .B2(n15326), .ZN(
        n12532) );
  AOI211_X1 U14897 ( .C1(n13313), .C2(n15372), .A(n12533), .B(n12532), .ZN(
        n12534) );
  OAI21_X1 U14898 ( .B1(n13214), .B2(n12535), .A(n12534), .ZN(P3_U3219) );
  INV_X1 U14899 ( .A(n12536), .ZN(n12537) );
  OAI222_X1 U14900 ( .A1(n14635), .A2(n12538), .B1(n14638), .B2(n12537), .C1(
        P1_U3086), .C2(n10373), .ZN(P1_U3327) );
  INV_X1 U14901 ( .A(n12539), .ZN(n12540) );
  AOI22_X1 U14902 ( .A1(n12540), .A2(n15120), .B1(n13496), .B2(n13684), .ZN(
        n12546) );
  NAND2_X1 U14903 ( .A1(n13669), .A2(n13816), .ZN(n12542) );
  NAND2_X1 U14904 ( .A1(n13742), .A2(n13814), .ZN(n12541) );
  NAND2_X1 U14905 ( .A1(n12542), .A2(n12541), .ZN(n13701) );
  AOI22_X1 U14906 ( .A1(n13701), .A2(n14845), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12543) );
  OAI21_X1 U14907 ( .B1(n13706), .B2(n15124), .A(n12543), .ZN(n12544) );
  AOI21_X1 U14908 ( .B1(n13875), .B2(n14848), .A(n12544), .ZN(n12545) );
  OAI21_X1 U14909 ( .B1(n12547), .B2(n12546), .A(n12545), .ZN(P2_U3207) );
  INV_X1 U14910 ( .A(n12594), .ZN(n14277) );
  INV_X1 U14911 ( .A(n14334), .ZN(n14339) );
  INV_X1 U14912 ( .A(n14352), .ZN(n14546) );
  INV_X1 U14913 ( .A(n14362), .ZN(n12564) );
  NAND2_X1 U14914 ( .A1(n12549), .A2(n12548), .ZN(n12551) );
  NAND2_X1 U14915 ( .A1(n12551), .A2(n12550), .ZN(n14476) );
  NAND2_X1 U14916 ( .A1(n14476), .A2(n14489), .ZN(n12553) );
  NAND2_X1 U14917 ( .A1(n12553), .A2(n12552), .ZN(n14458) );
  INV_X1 U14918 ( .A(n14458), .ZN(n12555) );
  INV_X1 U14919 ( .A(n14459), .ZN(n12554) );
  NAND2_X1 U14920 ( .A1(n14591), .A2(n14447), .ZN(n12556) );
  NAND2_X1 U14921 ( .A1(n14450), .A2(n12557), .ZN(n14423) );
  INV_X1 U14922 ( .A(n14422), .ZN(n14420) );
  OR2_X1 U14923 ( .A1(n14580), .A2(n14448), .ZN(n12558) );
  NAND2_X1 U14924 ( .A1(n14574), .A2(n14427), .ZN(n12560) );
  INV_X1 U14925 ( .A(n12586), .ZN(n14393) );
  NAND2_X1 U14926 ( .A1(n14401), .A2(n14409), .ZN(n12561) );
  INV_X1 U14927 ( .A(n14374), .ZN(n14371) );
  OR2_X1 U14928 ( .A1(n14381), .A2(n14396), .ZN(n12562) );
  NOR2_X1 U14929 ( .A1(n14286), .A2(n14301), .ZN(n12566) );
  NAND3_X1 U14930 ( .A1(n7370), .A2(n12595), .A3(n7369), .ZN(n12567) );
  INV_X1 U14931 ( .A(n12595), .ZN(n12597) );
  NAND2_X1 U14932 ( .A1(n14301), .A2(n14479), .ZN(n12569) );
  NAND2_X1 U14933 ( .A1(n14093), .A2(n14477), .ZN(n12568) );
  OR2_X2 U14934 ( .A1(n14595), .A2(n14484), .ZN(n14482) );
  INV_X1 U14935 ( .A(n14585), .ZN(n14444) );
  OR2_X2 U14936 ( .A1(n14551), .A2(n14376), .ZN(n14364) );
  OR2_X2 U14937 ( .A1(n14364), .A2(n14352), .ZN(n14346) );
  OR2_X2 U14938 ( .A1(n14334), .A2(n14346), .ZN(n14332) );
  INV_X1 U14939 ( .A(n14281), .ZN(n12572) );
  AOI211_X1 U14940 ( .C1(n14517), .C2(n12572), .A(n15014), .B(n14241), .ZN(
        n14516) );
  INV_X1 U14941 ( .A(n12784), .ZN(n12573) );
  AOI22_X1 U14942 ( .A1(n6550), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n12573), 
        .B2(n14888), .ZN(n12574) );
  OAI21_X1 U14943 ( .B1(n7158), .B2(n15009), .A(n12574), .ZN(n12601) );
  NAND2_X1 U14944 ( .A1(n12672), .A2(n14480), .ZN(n12575) );
  OR2_X1 U14945 ( .A1(n14591), .A2(n14478), .ZN(n12577) );
  INV_X1 U14946 ( .A(n14463), .ZN(n14425) );
  NOR2_X1 U14947 ( .A1(n14585), .A2(n14425), .ZN(n12578) );
  NAND2_X1 U14948 ( .A1(n14585), .A2(n14425), .ZN(n12579) );
  INV_X1 U14949 ( .A(n12580), .ZN(n12583) );
  INV_X1 U14950 ( .A(n12581), .ZN(n12582) );
  OR2_X1 U14951 ( .A1(n14574), .A2(n14096), .ZN(n12584) );
  NAND2_X1 U14952 ( .A1(n12585), .A2(n12584), .ZN(n14387) );
  OR2_X1 U14953 ( .A1(n14401), .A2(n13992), .ZN(n12587) );
  OR2_X1 U14954 ( .A1(n14381), .A2(n14359), .ZN(n12588) );
  NOR2_X1 U14955 ( .A1(n14352), .A2(n14358), .ZN(n12589) );
  NAND2_X1 U14956 ( .A1(n14352), .A2(n14358), .ZN(n12590) );
  OR2_X1 U14957 ( .A1(n14334), .A2(n14094), .ZN(n12591) );
  NAND2_X1 U14958 ( .A1(n12598), .A2(n12597), .ZN(n12599) );
  NAND2_X1 U14959 ( .A1(n14254), .A2(n12599), .ZN(n14520) );
  NOR2_X1 U14960 ( .A1(n14520), .A2(n14490), .ZN(n12600) );
  AOI211_X1 U14961 ( .C1(n15017), .C2(n14516), .A(n12601), .B(n12600), .ZN(
        n12602) );
  OAI21_X1 U14962 ( .B1(n14519), .B2(n6550), .A(n12602), .ZN(P1_U3265) );
  INV_X1 U14963 ( .A(n12604), .ZN(n12605) );
  AOI22_X1 U14964 ( .A1(n13812), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n12605), 
        .B2(n13825), .ZN(n12606) );
  OAI21_X1 U14965 ( .B1(n7495), .B2(n13828), .A(n12606), .ZN(n12608) );
  XNOR2_X1 U14966 ( .A(n13367), .B(n12640), .ZN(n12613) );
  INV_X1 U14967 ( .A(n12613), .ZN(n12614) );
  XNOR2_X1 U14968 ( .A(n12613), .B(n13245), .ZN(n12835) );
  XNOR2_X1 U14969 ( .A(n13363), .B(n12640), .ZN(n12615) );
  XNOR2_X1 U14970 ( .A(n12615), .B(n13232), .ZN(n12844) );
  NAND2_X1 U14971 ( .A1(n12615), .A2(n12897), .ZN(n12616) );
  XNOR2_X1 U14972 ( .A(n13359), .B(n11571), .ZN(n12878) );
  NOR2_X1 U14973 ( .A1(n12878), .A2(n13218), .ZN(n12617) );
  XNOR2_X1 U14974 ( .A(n13355), .B(n12640), .ZN(n12618) );
  XNOR2_X1 U14975 ( .A(n12618), .B(n13172), .ZN(n12811) );
  NAND2_X1 U14976 ( .A1(n12618), .A2(n13172), .ZN(n12619) );
  XNOR2_X1 U14977 ( .A(n13289), .B(n12640), .ZN(n12620) );
  XNOR2_X1 U14978 ( .A(n12620), .B(n13187), .ZN(n12863) );
  INV_X1 U14979 ( .A(n12620), .ZN(n12621) );
  NAND2_X1 U14980 ( .A1(n12621), .A2(n13187), .ZN(n12622) );
  XNOR2_X1 U14981 ( .A(n13349), .B(n12640), .ZN(n12623) );
  XNOR2_X1 U14982 ( .A(n12623), .B(n12871), .ZN(n12820) );
  XNOR2_X1 U14983 ( .A(n12808), .B(n12640), .ZN(n12628) );
  INV_X1 U14984 ( .A(n12628), .ZN(n12629) );
  OR2_X1 U14985 ( .A1(n12630), .A2(n12629), .ZN(n12631) );
  XNOR2_X1 U14986 ( .A(n13341), .B(n12640), .ZN(n12633) );
  XNOR2_X1 U14987 ( .A(n12633), .B(n13131), .ZN(n12854) );
  INV_X1 U14988 ( .A(n12633), .ZN(n12634) );
  NAND2_X1 U14989 ( .A1(n12634), .A2(n13131), .ZN(n12635) );
  XNOR2_X1 U14990 ( .A(n13337), .B(n12640), .ZN(n12636) );
  XNOR2_X1 U14991 ( .A(n12636), .B(n13089), .ZN(n12827) );
  INV_X1 U14992 ( .A(n12636), .ZN(n12637) );
  XNOR2_X1 U14993 ( .A(n13093), .B(n12640), .ZN(n12638) );
  XNOR2_X1 U14994 ( .A(n12638), .B(n13104), .ZN(n12888) );
  XNOR2_X1 U14995 ( .A(n12802), .B(n12640), .ZN(n12641) );
  INV_X1 U14996 ( .A(n13090), .ZN(n13072) );
  XNOR2_X1 U14997 ( .A(n12641), .B(n13072), .ZN(n12796) );
  NOR2_X1 U14998 ( .A1(n13074), .A2(n12891), .ZN(n12645) );
  AOI22_X1 U14999 ( .A1(n13075), .A2(n15439), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12643) );
  OAI21_X1 U15000 ( .B1(n13090), .B2(n12870), .A(n12643), .ZN(n12644) );
  AOI211_X1 U15001 ( .C1(n12646), .C2(n15425), .A(n12645), .B(n12644), .ZN(
        n12647) );
  OAI222_X1 U15002 ( .A1(n13964), .A2(n12650), .B1(n12649), .B2(n12648), .C1(
        n6555), .C2(P2_U3088), .ZN(P2_U3308) );
  INV_X1 U15003 ( .A(n12651), .ZN(n12654) );
  OAI222_X1 U15004 ( .A1(n14743), .A2(n12654), .B1(n14741), .B2(n12653), .C1(
        P3_U3151), .C2(n12652), .ZN(P3_U3267) );
  INV_X1 U15005 ( .A(n12655), .ZN(n12656) );
  OAI222_X1 U15006 ( .A1(n12657), .A2(P3_U3151), .B1(n14741), .B2(n15514), 
        .C1(n14743), .C2(n12656), .ZN(P3_U3265) );
  AND2_X1 U15007 ( .A1(n14096), .A2(n12770), .ZN(n12658) );
  AOI21_X1 U15008 ( .B1(n14574), .B2(n12743), .A(n12658), .ZN(n12709) );
  NAND2_X1 U15009 ( .A1(n14574), .A2(n12753), .ZN(n12660) );
  NAND2_X1 U15010 ( .A1(n14096), .A2(n12743), .ZN(n12659) );
  NAND2_X1 U15011 ( .A1(n12660), .A2(n12659), .ZN(n12661) );
  XNOR2_X1 U15012 ( .A(n12661), .B(n12777), .ZN(n12704) );
  INV_X1 U15013 ( .A(n12662), .ZN(n12663) );
  NAND2_X1 U15014 ( .A1(n12672), .A2(n12753), .ZN(n12668) );
  NAND2_X1 U15015 ( .A1(n12743), .A2(n14480), .ZN(n12667) );
  NAND2_X1 U15016 ( .A1(n12668), .A2(n12667), .ZN(n12669) );
  XNOR2_X1 U15017 ( .A(n12669), .B(n12746), .ZN(n12674) );
  NOR2_X1 U15018 ( .A1(n12776), .A2(n12670), .ZN(n12671) );
  AOI21_X1 U15019 ( .B1(n12672), .B2(n12743), .A(n12671), .ZN(n12673) );
  NAND2_X1 U15020 ( .A1(n12674), .A2(n12673), .ZN(n12675) );
  OAI21_X1 U15021 ( .B1(n12674), .B2(n12673), .A(n12675), .ZN(n14860) );
  NOR2_X1 U15022 ( .A1(n14859), .A2(n14860), .ZN(n14858) );
  INV_X1 U15023 ( .A(n12675), .ZN(n12676) );
  NOR2_X1 U15024 ( .A1(n14858), .A2(n12676), .ZN(n12678) );
  AOI22_X1 U15025 ( .A1(n14595), .A2(n12753), .B1(n12743), .B2(n14097), .ZN(
        n12677) );
  XOR2_X1 U15026 ( .A(n12777), .B(n12677), .Z(n12679) );
  INV_X1 U15027 ( .A(n12678), .ZN(n12682) );
  INV_X1 U15028 ( .A(n12679), .ZN(n12681) );
  INV_X1 U15029 ( .A(n12683), .ZN(n12680) );
  OAI22_X1 U15030 ( .A1(n7116), .A2(n12779), .B1(n14461), .B2(n12776), .ZN(
        n14084) );
  NAND2_X1 U15031 ( .A1(n14591), .A2(n12753), .ZN(n12685) );
  NAND2_X1 U15032 ( .A1(n14478), .A2(n12743), .ZN(n12684) );
  NAND2_X1 U15033 ( .A1(n12685), .A2(n12684), .ZN(n12686) );
  XNOR2_X1 U15034 ( .A(n12686), .B(n12746), .ZN(n12689) );
  AND2_X1 U15035 ( .A1(n14478), .A2(n12770), .ZN(n12687) );
  AOI21_X1 U15036 ( .B1(n14591), .B2(n12743), .A(n12687), .ZN(n12688) );
  NAND2_X1 U15037 ( .A1(n12689), .A2(n12688), .ZN(n12690) );
  OAI21_X1 U15038 ( .B1(n12689), .B2(n12688), .A(n12690), .ZN(n14016) );
  INV_X1 U15039 ( .A(n12690), .ZN(n14026) );
  NAND2_X1 U15040 ( .A1(n14585), .A2(n12753), .ZN(n12692) );
  NAND2_X1 U15041 ( .A1(n14425), .A2(n12743), .ZN(n12691) );
  NAND2_X1 U15042 ( .A1(n12692), .A2(n12691), .ZN(n12693) );
  XNOR2_X1 U15043 ( .A(n12693), .B(n12746), .ZN(n12695) );
  NOR2_X1 U15044 ( .A1(n14463), .A2(n12776), .ZN(n12694) );
  AOI21_X1 U15045 ( .B1(n14585), .B2(n12743), .A(n12694), .ZN(n12696) );
  NAND2_X1 U15046 ( .A1(n12695), .A2(n12696), .ZN(n12700) );
  INV_X1 U15047 ( .A(n12695), .ZN(n12698) );
  INV_X1 U15048 ( .A(n12696), .ZN(n12697) );
  NAND2_X1 U15049 ( .A1(n12698), .A2(n12697), .ZN(n12699) );
  AND2_X1 U15050 ( .A1(n12700), .A2(n12699), .ZN(n14025) );
  NAND2_X1 U15051 ( .A1(n14024), .A2(n12700), .ZN(n14062) );
  NAND2_X1 U15052 ( .A1(n14580), .A2(n12753), .ZN(n12702) );
  NAND2_X1 U15053 ( .A1(n14408), .A2(n12743), .ZN(n12701) );
  NAND2_X1 U15054 ( .A1(n12702), .A2(n12701), .ZN(n12703) );
  XNOR2_X1 U15055 ( .A(n12703), .B(n12777), .ZN(n12705) );
  AOI22_X1 U15056 ( .A1(n14580), .A2(n12743), .B1(n12770), .B2(n14408), .ZN(
        n12706) );
  XNOR2_X1 U15057 ( .A(n12705), .B(n12706), .ZN(n14063) );
  XNOR2_X1 U15058 ( .A(n12704), .B(n12709), .ZN(n13990) );
  INV_X1 U15059 ( .A(n12705), .ZN(n12707) );
  NAND2_X1 U15060 ( .A1(n12707), .A2(n12706), .ZN(n13988) );
  OR2_X1 U15061 ( .A1(n14401), .A2(n12779), .ZN(n12711) );
  NAND2_X1 U15062 ( .A1(n14409), .A2(n12770), .ZN(n12710) );
  NAND2_X1 U15063 ( .A1(n12711), .A2(n12710), .ZN(n12714) );
  OAI22_X1 U15064 ( .A1(n14401), .A2(n11135), .B1(n13992), .B2(n12779), .ZN(
        n12712) );
  XNOR2_X1 U15065 ( .A(n12712), .B(n12777), .ZN(n12713) );
  XOR2_X1 U15066 ( .A(n12714), .B(n12713), .Z(n14041) );
  NAND2_X1 U15067 ( .A1(n14381), .A2(n12753), .ZN(n12716) );
  NAND2_X1 U15068 ( .A1(n14359), .A2(n12743), .ZN(n12715) );
  NAND2_X1 U15069 ( .A1(n12716), .A2(n12715), .ZN(n12717) );
  XNOR2_X1 U15070 ( .A(n12717), .B(n12777), .ZN(n12721) );
  NAND2_X1 U15071 ( .A1(n14381), .A2(n12743), .ZN(n12719) );
  NAND2_X1 U15072 ( .A1(n14359), .A2(n12770), .ZN(n12718) );
  NAND2_X1 U15073 ( .A1(n12719), .A2(n12718), .ZN(n12720) );
  NOR2_X1 U15074 ( .A1(n12721), .A2(n12720), .ZN(n12722) );
  AOI21_X1 U15075 ( .B1(n12721), .B2(n12720), .A(n12722), .ZN(n13998) );
  INV_X1 U15076 ( .A(n12722), .ZN(n12723) );
  NAND2_X1 U15077 ( .A1(n13997), .A2(n12723), .ZN(n14051) );
  NAND2_X1 U15078 ( .A1(n14551), .A2(n12753), .ZN(n12725) );
  NAND2_X1 U15079 ( .A1(n14095), .A2(n12743), .ZN(n12724) );
  NAND2_X1 U15080 ( .A1(n12725), .A2(n12724), .ZN(n12726) );
  XNOR2_X1 U15081 ( .A(n12726), .B(n12777), .ZN(n12730) );
  NAND2_X1 U15082 ( .A1(n14551), .A2(n12743), .ZN(n12728) );
  NAND2_X1 U15083 ( .A1(n14095), .A2(n12770), .ZN(n12727) );
  NAND2_X1 U15084 ( .A1(n12728), .A2(n12727), .ZN(n12729) );
  NOR2_X1 U15085 ( .A1(n12730), .A2(n12729), .ZN(n12731) );
  AOI21_X1 U15086 ( .B1(n12730), .B2(n12729), .A(n12731), .ZN(n14052) );
  INV_X1 U15087 ( .A(n12731), .ZN(n13979) );
  NAND2_X1 U15088 ( .A1(n14352), .A2(n12753), .ZN(n12733) );
  NAND2_X1 U15089 ( .A1(n12743), .A2(n14358), .ZN(n12732) );
  NAND2_X1 U15090 ( .A1(n12733), .A2(n12732), .ZN(n12734) );
  XNOR2_X1 U15091 ( .A(n12734), .B(n12746), .ZN(n12736) );
  NOR2_X1 U15092 ( .A1(n12776), .A2(n7703), .ZN(n12735) );
  AOI21_X1 U15093 ( .B1(n14352), .B2(n12743), .A(n12735), .ZN(n12737) );
  NAND2_X1 U15094 ( .A1(n12736), .A2(n12737), .ZN(n12741) );
  INV_X1 U15095 ( .A(n12736), .ZN(n12739) );
  INV_X1 U15096 ( .A(n12737), .ZN(n12738) );
  NAND2_X1 U15097 ( .A1(n12739), .A2(n12738), .ZN(n12740) );
  NAND2_X1 U15098 ( .A1(n12741), .A2(n12740), .ZN(n13978) );
  INV_X1 U15099 ( .A(n12741), .ZN(n12742) );
  NAND2_X1 U15100 ( .A1(n14334), .A2(n12753), .ZN(n12745) );
  NAND2_X1 U15101 ( .A1(n12743), .A2(n14094), .ZN(n12744) );
  NAND2_X1 U15102 ( .A1(n12745), .A2(n12744), .ZN(n12747) );
  XNOR2_X1 U15103 ( .A(n12747), .B(n12746), .ZN(n12751) );
  NOR2_X1 U15104 ( .A1(n12776), .A2(n12748), .ZN(n12749) );
  AOI21_X1 U15105 ( .B1(n14334), .B2(n12743), .A(n12749), .ZN(n12750) );
  NAND2_X1 U15106 ( .A1(n12751), .A2(n12750), .ZN(n12752) );
  NAND2_X1 U15107 ( .A1(n14535), .A2(n12753), .ZN(n12755) );
  NAND2_X1 U15108 ( .A1(n12743), .A2(n14325), .ZN(n12754) );
  NAND2_X1 U15109 ( .A1(n12755), .A2(n12754), .ZN(n12756) );
  XNOR2_X1 U15110 ( .A(n12756), .B(n12777), .ZN(n12760) );
  NAND2_X1 U15111 ( .A1(n14535), .A2(n12743), .ZN(n12758) );
  NAND2_X1 U15112 ( .A1(n12770), .A2(n14325), .ZN(n12757) );
  NAND2_X1 U15113 ( .A1(n12758), .A2(n12757), .ZN(n12759) );
  NOR2_X1 U15114 ( .A1(n12760), .A2(n12759), .ZN(n12761) );
  AOI21_X1 U15115 ( .B1(n12760), .B2(n12759), .A(n12761), .ZN(n14008) );
  OAI22_X1 U15116 ( .A1(n14297), .A2(n11135), .B1(n14275), .B2(n12779), .ZN(
        n12762) );
  XNOR2_X1 U15117 ( .A(n12762), .B(n12777), .ZN(n12766) );
  OR2_X1 U15118 ( .A1(n14297), .A2(n12779), .ZN(n12764) );
  NAND2_X1 U15119 ( .A1(n12770), .A2(n7446), .ZN(n12763) );
  NAND2_X1 U15120 ( .A1(n12764), .A2(n12763), .ZN(n12765) );
  NOR2_X1 U15121 ( .A1(n12766), .A2(n12765), .ZN(n12767) );
  AOI21_X1 U15122 ( .B1(n12766), .B2(n12765), .A(n12767), .ZN(n14073) );
  INV_X1 U15123 ( .A(n12767), .ZN(n12768) );
  OAI22_X1 U15124 ( .A1(n14286), .A2(n11135), .B1(n14076), .B2(n12779), .ZN(
        n12769) );
  XNOR2_X1 U15125 ( .A(n12769), .B(n12777), .ZN(n12774) );
  OR2_X1 U15126 ( .A1(n14286), .A2(n12779), .ZN(n12772) );
  NAND2_X1 U15127 ( .A1(n12770), .A2(n14301), .ZN(n12771) );
  NAND2_X1 U15128 ( .A1(n12772), .A2(n12771), .ZN(n12773) );
  NOR2_X1 U15129 ( .A1(n12774), .A2(n12773), .ZN(n12775) );
  AOI21_X1 U15130 ( .B1(n12774), .B2(n12773), .A(n12775), .ZN(n13972) );
  OAI22_X1 U15131 ( .A1(n7158), .A2(n12779), .B1(n14274), .B2(n12776), .ZN(
        n12778) );
  XNOR2_X1 U15132 ( .A(n12778), .B(n12777), .ZN(n12781) );
  OAI22_X1 U15133 ( .A1(n7158), .A2(n11135), .B1(n14274), .B2(n12779), .ZN(
        n12780) );
  XNOR2_X1 U15134 ( .A(n12781), .B(n12780), .ZN(n12782) );
  XNOR2_X1 U15135 ( .A(n12783), .B(n12782), .ZN(n12790) );
  NOR2_X1 U15136 ( .A1(n14965), .A2(n12784), .ZN(n12788) );
  AOI22_X1 U15137 ( .A1(n14087), .A2(n14301), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12785) );
  OAI21_X1 U15138 ( .B1(n12786), .B2(n14085), .A(n12785), .ZN(n12787) );
  AOI211_X1 U15139 ( .C1(n14517), .C2(n14090), .A(n12788), .B(n12787), .ZN(
        n12789) );
  OAI21_X1 U15140 ( .B1(n12790), .B2(n14935), .A(n12789), .ZN(P1_U3220) );
  INV_X1 U15141 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n12793) );
  AND2_X1 U15142 ( .A1(n12791), .A2(n14634), .ZN(n12792) );
  AOI22_X1 U15143 ( .A1(n15022), .A2(n12793), .B1(n12792), .B2(n10551), .ZN(
        P1_U3446) );
  INV_X1 U15144 ( .A(n12794), .ZN(n13962) );
  OAI222_X1 U15145 ( .A1(n14635), .A2(n12795), .B1(n14638), .B2(n13962), .C1(
        P1_U3086), .C2(n10551), .ZN(P1_U3330) );
  INV_X1 U15146 ( .A(n12796), .ZN(n12797) );
  NOR2_X1 U15147 ( .A1(n12798), .A2(n12891), .ZN(n12801) );
  AOI22_X1 U15148 ( .A1(n13082), .A2(n15439), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12799) );
  OAI21_X1 U15149 ( .B1(n12830), .B2(n12870), .A(n12799), .ZN(n12800) );
  AOI211_X1 U15150 ( .C1(n12802), .C2(n15425), .A(n12801), .B(n12800), .ZN(
        n12803) );
  XNOR2_X1 U15151 ( .A(n12804), .B(n13141), .ZN(n12810) );
  AOI22_X1 U15152 ( .A1(n12896), .A2(n15422), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12806) );
  NAND2_X1 U15153 ( .A1(n13135), .A2(n15439), .ZN(n12805) );
  OAI211_X1 U15154 ( .C1(n13131), .C2(n12891), .A(n12806), .B(n12805), .ZN(
        n12807) );
  AOI21_X1 U15155 ( .B1(n12808), .B2(n15425), .A(n12807), .ZN(n12809) );
  OAI21_X1 U15156 ( .B1(n12810), .B2(n15434), .A(n12809), .ZN(P3_U3156) );
  AOI21_X1 U15157 ( .B1(n12812), .B2(n12811), .A(n15434), .ZN(n12814) );
  NAND2_X1 U15158 ( .A1(n12814), .A2(n12813), .ZN(n12818) );
  NAND2_X1 U15159 ( .A1(n13186), .A2(n15422), .ZN(n12815) );
  NAND2_X1 U15160 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13039)
         );
  OAI211_X1 U15161 ( .C1(n13156), .C2(n12891), .A(n12815), .B(n13039), .ZN(
        n12816) );
  AOI21_X1 U15162 ( .B1(n13190), .B2(n15439), .A(n12816), .ZN(n12817) );
  OAI211_X1 U15163 ( .C1(n12882), .C2(n13355), .A(n12818), .B(n12817), .ZN(
        P3_U3159) );
  AOI21_X1 U15164 ( .B1(n12820), .B2(n12819), .A(n6709), .ZN(n12825) );
  AOI22_X1 U15165 ( .A1(n13187), .A2(n15422), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12822) );
  NAND2_X1 U15166 ( .A1(n13161), .A2(n15439), .ZN(n12821) );
  OAI211_X1 U15167 ( .C1(n13157), .C2(n12891), .A(n12822), .B(n12821), .ZN(
        n12823) );
  AOI21_X1 U15168 ( .B1(n13349), .B2(n15425), .A(n12823), .ZN(n12824) );
  OAI21_X1 U15169 ( .B1(n12825), .B2(n15434), .A(n12824), .ZN(P3_U3163) );
  XOR2_X1 U15170 ( .A(n12827), .B(n12826), .Z(n12834) );
  INV_X1 U15171 ( .A(n13131), .ZN(n13103) );
  AOI22_X1 U15172 ( .A1(n13103), .A2(n15422), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12829) );
  NAND2_X1 U15173 ( .A1(n13109), .A2(n15439), .ZN(n12828) );
  OAI211_X1 U15174 ( .C1(n12830), .C2(n12891), .A(n12829), .B(n12828), .ZN(
        n12831) );
  AOI21_X1 U15175 ( .B1(n12832), .B2(n15425), .A(n12831), .ZN(n12833) );
  OAI21_X1 U15176 ( .B1(n12834), .B2(n15434), .A(n12833), .ZN(P3_U3165) );
  XNOR2_X1 U15177 ( .A(n12836), .B(n12835), .ZN(n12843) );
  INV_X1 U15178 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n12837) );
  OR2_X1 U15179 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12837), .ZN(n12966) );
  OAI21_X1 U15180 ( .B1(n13232), .B2(n12891), .A(n12966), .ZN(n12838) );
  AOI21_X1 U15181 ( .B1(n15422), .B2(n12899), .A(n12838), .ZN(n12839) );
  OAI21_X1 U15182 ( .B1(n13236), .B2(n12848), .A(n12839), .ZN(n12840) );
  AOI21_X1 U15183 ( .B1(n12841), .B2(n15425), .A(n12840), .ZN(n12842) );
  OAI21_X1 U15184 ( .B1(n12843), .B2(n15434), .A(n12842), .ZN(P3_U3166) );
  XNOR2_X1 U15185 ( .A(n12845), .B(n12844), .ZN(n12852) );
  NAND2_X1 U15186 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12996)
         );
  OAI21_X1 U15187 ( .B1(n13218), .B2(n12891), .A(n12996), .ZN(n12846) );
  AOI21_X1 U15188 ( .B1(n15422), .B2(n12898), .A(n12846), .ZN(n12847) );
  OAI21_X1 U15189 ( .B1(n13222), .B2(n12848), .A(n12847), .ZN(n12849) );
  AOI21_X1 U15190 ( .B1(n12850), .B2(n15425), .A(n12849), .ZN(n12851) );
  OAI21_X1 U15191 ( .B1(n12852), .B2(n15434), .A(n12851), .ZN(P3_U3168) );
  XOR2_X1 U15192 ( .A(n12854), .B(n12853), .Z(n12860) );
  AOI22_X1 U15193 ( .A1(n13141), .A2(n15422), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12856) );
  NAND2_X1 U15194 ( .A1(n13121), .A2(n15439), .ZN(n12855) );
  OAI211_X1 U15195 ( .C1(n13089), .C2(n12891), .A(n12856), .B(n12855), .ZN(
        n12857) );
  AOI21_X1 U15196 ( .B1(n12858), .B2(n15425), .A(n12857), .ZN(n12859) );
  OAI21_X1 U15197 ( .B1(n12860), .B2(n15434), .A(n12859), .ZN(P3_U3169) );
  INV_X1 U15198 ( .A(n13289), .ZN(n13178) );
  OAI211_X1 U15199 ( .C1(n12864), .C2(n12863), .A(n12862), .B(n12861), .ZN(
        n12868) );
  AOI22_X1 U15200 ( .A1(n13172), .A2(n15422), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12865) );
  OAI21_X1 U15201 ( .B1(n12871), .B2(n12891), .A(n12865), .ZN(n12866) );
  AOI21_X1 U15202 ( .B1(n13176), .B2(n15439), .A(n12866), .ZN(n12867) );
  OAI211_X1 U15203 ( .C1(n13178), .C2(n12882), .A(n12868), .B(n12867), .ZN(
        P3_U3173) );
  XNOR2_X1 U15204 ( .A(n12869), .B(n12896), .ZN(n12877) );
  NOR2_X1 U15205 ( .A1(n12871), .A2(n12870), .ZN(n12874) );
  INV_X1 U15206 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n15619) );
  OAI22_X1 U15207 ( .A1(n12872), .A2(n12891), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15619), .ZN(n12873) );
  AOI211_X1 U15208 ( .C1(n13145), .C2(n15439), .A(n12874), .B(n12873), .ZN(
        n12876) );
  NAND2_X1 U15209 ( .A1(n13280), .A2(n15425), .ZN(n12875) );
  OAI211_X1 U15210 ( .C1(n12877), .C2(n15434), .A(n12876), .B(n12875), .ZN(
        P3_U3175) );
  XNOR2_X1 U15211 ( .A(n12878), .B(n13186), .ZN(n12879) );
  XNOR2_X1 U15212 ( .A(n12880), .B(n12879), .ZN(n12886) );
  NAND2_X1 U15213 ( .A1(n12897), .A2(n15422), .ZN(n12881) );
  NAND2_X1 U15214 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13011)
         );
  OAI211_X1 U15215 ( .C1(n13204), .C2(n12891), .A(n12881), .B(n13011), .ZN(
        n12884) );
  NOR2_X1 U15216 ( .A1(n13359), .A2(n12882), .ZN(n12883) );
  AOI211_X1 U15217 ( .C1(n13205), .C2(n15439), .A(n12884), .B(n12883), .ZN(
        n12885) );
  OAI21_X1 U15218 ( .B1(n12886), .B2(n15434), .A(n12885), .ZN(P3_U3178) );
  XOR2_X1 U15219 ( .A(n12888), .B(n12887), .Z(n12894) );
  INV_X1 U15220 ( .A(n13089), .ZN(n13115) );
  AOI22_X1 U15221 ( .A1(n13115), .A2(n15422), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12890) );
  NAND2_X1 U15222 ( .A1(n13094), .A2(n15439), .ZN(n12889) );
  OAI211_X1 U15223 ( .C1(n13090), .C2(n12891), .A(n12890), .B(n12889), .ZN(
        n12892) );
  AOI21_X1 U15224 ( .B1(n13093), .B2(n15425), .A(n12892), .ZN(n12893) );
  OAI21_X1 U15225 ( .B1(n12894), .B2(n15434), .A(n12893), .ZN(P3_U3180) );
  MUX2_X1 U15226 ( .A(n12895), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12902), .Z(
        P3_U3522) );
  MUX2_X1 U15227 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n13072), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15228 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n13115), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U15229 ( .A(n13103), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12902), .Z(
        P3_U3515) );
  MUX2_X1 U15230 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n13141), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U15231 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12896), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15232 ( .A(n13171), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12902), .Z(
        P3_U3512) );
  MUX2_X1 U15233 ( .A(n13172), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12902), .Z(
        P3_U3510) );
  MUX2_X1 U15234 ( .A(n13186), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12902), .Z(
        P3_U3509) );
  MUX2_X1 U15235 ( .A(n12897), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12902), .Z(
        P3_U3508) );
  MUX2_X1 U15236 ( .A(n12898), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12902), .Z(
        P3_U3507) );
  MUX2_X1 U15237 ( .A(n12899), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12902), .Z(
        P3_U3506) );
  MUX2_X1 U15238 ( .A(n12900), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12902), .Z(
        P3_U3505) );
  MUX2_X1 U15239 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12901), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U15240 ( .A(n14809), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12902), .Z(
        P3_U3503) );
  MUX2_X1 U15241 ( .A(n15282), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12902), .Z(
        P3_U3502) );
  MUX2_X1 U15242 ( .A(n14810), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12902), .Z(
        P3_U3501) );
  MUX2_X1 U15243 ( .A(n15311), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12902), .Z(
        P3_U3500) );
  MUX2_X1 U15244 ( .A(n15330), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12902), .Z(
        P3_U3499) );
  MUX2_X1 U15245 ( .A(n15310), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12902), .Z(
        P3_U3498) );
  MUX2_X1 U15246 ( .A(n15331), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12902), .Z(
        P3_U3497) );
  MUX2_X1 U15247 ( .A(n15421), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12902), .Z(
        P3_U3495) );
  MUX2_X1 U15248 ( .A(n15343), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12902), .Z(
        P3_U3494) );
  MUX2_X1 U15249 ( .A(n15359), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12902), .Z(
        P3_U3491) );
  AOI21_X1 U15250 ( .B1(n12903), .B2(n8862), .A(n12920), .ZN(n12918) );
  MUX2_X1 U15251 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12946), .Z(n12925) );
  INV_X1 U15252 ( .A(n12924), .ZN(n12929) );
  XNOR2_X1 U15253 ( .A(n12925), .B(n12929), .ZN(n12906) );
  OAI21_X1 U15254 ( .B1(n12907), .B2(n12906), .A(n12923), .ZN(n12915) );
  AOI21_X1 U15255 ( .B1(n15280), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12908), 
        .ZN(n12909) );
  OAI21_X1 U15256 ( .B1(n12935), .B2(n12924), .A(n12909), .ZN(n12914) );
  AOI21_X1 U15257 ( .B1(n8863), .B2(n12911), .A(n12930), .ZN(n12912) );
  NOR2_X1 U15258 ( .A1(n12912), .A2(n13004), .ZN(n12913) );
  AOI211_X1 U15259 ( .C1(n12916), .C2(n12915), .A(n12914), .B(n12913), .ZN(
        n12917) );
  OAI21_X1 U15260 ( .B1(n12918), .B2(n13040), .A(n12917), .ZN(P3_U3195) );
  XNOR2_X1 U15261 ( .A(n12954), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n12922) );
  AOI21_X1 U15262 ( .B1(n12921), .B2(n12922), .A(n12953), .ZN(n12940) );
  XNOR2_X1 U15263 ( .A(n12954), .B(P3_REG1_REG_14__SCAN_IN), .ZN(n12931) );
  MUX2_X1 U15264 ( .A(n12922), .B(n12931), .S(n12946), .Z(n12927) );
  AOI211_X1 U15265 ( .C1(n12927), .C2(n12926), .A(n13051), .B(n12947), .ZN(
        n12938) );
  AOI21_X1 U15266 ( .B1(n6717), .B2(n12931), .A(n12941), .ZN(n12932) );
  NOR2_X1 U15267 ( .A1(n12932), .A2(n13004), .ZN(n12937) );
  AOI21_X1 U15268 ( .B1(n15280), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12933), 
        .ZN(n12934) );
  OAI21_X1 U15269 ( .B1(n12935), .B2(n12954), .A(n12934), .ZN(n12936) );
  NOR3_X1 U15270 ( .A1(n12938), .A2(n12937), .A3(n12936), .ZN(n12939) );
  OAI21_X1 U15271 ( .B1(n12940), .B2(n13040), .A(n12939), .ZN(P3_U3196) );
  AOI21_X1 U15272 ( .B1(n15480), .B2(n12942), .A(n12961), .ZN(n12959) );
  NAND2_X1 U15273 ( .A1(n15280), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n12945) );
  INV_X1 U15274 ( .A(n12943), .ZN(n12944) );
  NAND2_X1 U15275 ( .A1(n12945), .A2(n12944), .ZN(n12952) );
  MUX2_X1 U15276 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n12946), .Z(n12948) );
  MUX2_X1 U15277 ( .A(n13251), .B(n15480), .S(n12946), .Z(n12949) );
  AOI211_X1 U15278 ( .C1(n12950), .C2(n12949), .A(n13051), .B(n12969), .ZN(
        n12951) );
  AOI211_X1 U15279 ( .C1(n13041), .C2(n12977), .A(n12952), .B(n12951), .ZN(
        n12958) );
  AOI21_X1 U15280 ( .B1(n12955), .B2(n13251), .A(n12978), .ZN(n12956) );
  OR2_X1 U15281 ( .A1(n12956), .A2(n13040), .ZN(n12957) );
  OAI211_X1 U15282 ( .C1(n12959), .C2(n13004), .A(n12958), .B(n12957), .ZN(
        P3_U3197) );
  NOR2_X1 U15283 ( .A1(n12977), .A2(n12960), .ZN(n12962) );
  NAND2_X1 U15284 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12998), .ZN(n12963) );
  OAI21_X1 U15285 ( .B1(P3_REG1_REG_16__SCAN_IN), .B2(n12998), .A(n12963), 
        .ZN(n12964) );
  AOI21_X1 U15286 ( .B1(n12965), .B2(n12964), .A(n12987), .ZN(n12985) );
  NAND2_X1 U15287 ( .A1(n15280), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n12967) );
  NAND2_X1 U15288 ( .A1(n12967), .A2(n12966), .ZN(n12975) );
  MUX2_X1 U15289 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n12946), .Z(n12999) );
  XNOR2_X1 U15290 ( .A(n12999), .B(n12998), .ZN(n12973) );
  INV_X1 U15291 ( .A(n12977), .ZN(n12971) );
  INV_X1 U15292 ( .A(n12968), .ZN(n12970) );
  NOR2_X1 U15293 ( .A1(n12972), .A2(n12973), .ZN(n12997) );
  AOI211_X1 U15294 ( .C1(n12973), .C2(n12972), .A(n13051), .B(n12997), .ZN(
        n12974) );
  AOI211_X1 U15295 ( .C1(n13041), .C2(n12976), .A(n12975), .B(n12974), .ZN(
        n12984) );
  NAND2_X1 U15296 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12998), .ZN(n12980) );
  OAI21_X1 U15297 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n12998), .A(n12980), 
        .ZN(n12981) );
  AOI21_X1 U15298 ( .B1(n6687), .B2(n12981), .A(n12990), .ZN(n12982) );
  OR2_X1 U15299 ( .A1(n12982), .A2(n13040), .ZN(n12983) );
  OAI211_X1 U15300 ( .C1(n12985), .C2(n13004), .A(n12984), .B(n12983), .ZN(
        P3_U3198) );
  AND2_X1 U15301 ( .A1(n12998), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n12986) );
  INV_X1 U15302 ( .A(n13024), .ZN(n12988) );
  AOI21_X1 U15303 ( .B1(n13304), .B2(n12989), .A(n12988), .ZN(n13005) );
  INV_X1 U15304 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14730) );
  OAI21_X1 U15305 ( .B1(P3_REG2_REG_17__SCAN_IN), .B2(n12993), .A(n13017), 
        .ZN(n12994) );
  MUX2_X1 U15306 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12946), .Z(n13008) );
  XNOR2_X1 U15307 ( .A(n13008), .B(n13007), .ZN(n13001) );
  AOI211_X1 U15308 ( .C1(n13001), .C2(n13000), .A(n13051), .B(n13006), .ZN(
        n13002) );
  OAI21_X1 U15309 ( .B1(n13005), .B2(n13004), .A(n6683), .ZN(P3_U3199) );
  MUX2_X1 U15310 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12946), .Z(n13010) );
  AOI21_X1 U15311 ( .B1(n13010), .B2(n13009), .A(n13029), .ZN(n13028) );
  INV_X1 U15312 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14800) );
  OAI21_X1 U15313 ( .B1(n13012), .B2(n14800), .A(n13011), .ZN(n13020) );
  INV_X1 U15314 ( .A(n13013), .ZN(n13016) );
  OR2_X1 U15315 ( .A1(n13030), .A2(n13207), .ZN(n13036) );
  NAND2_X1 U15316 ( .A1(n13030), .A2(n13207), .ZN(n13014) );
  NAND2_X1 U15317 ( .A1(n13036), .A2(n13014), .ZN(n13015) );
  NAND3_X1 U15318 ( .A1(n13017), .A2(n13016), .A3(n13015), .ZN(n13018) );
  OR2_X1 U15319 ( .A1(n13030), .A2(n13300), .ZN(n13043) );
  NAND2_X1 U15320 ( .A1(n13030), .A2(n13300), .ZN(n13021) );
  NAND2_X1 U15321 ( .A1(n13043), .A2(n13021), .ZN(n13022) );
  AOI21_X1 U15322 ( .B1(n13024), .B2(n13023), .A(n13022), .ZN(n13045) );
  AND3_X1 U15323 ( .A1(n13024), .A2(n13023), .A3(n13022), .ZN(n13025) );
  OAI21_X1 U15324 ( .B1(n13045), .B2(n13025), .A(n13049), .ZN(n13026) );
  OAI211_X1 U15325 ( .C1(n13028), .C2(n13051), .A(n13027), .B(n13026), .ZN(
        P3_U3200) );
  XNOR2_X1 U15326 ( .A(n13033), .B(n13032), .ZN(n13038) );
  XNOR2_X1 U15327 ( .A(n13033), .B(n13296), .ZN(n13046) );
  MUX2_X1 U15328 ( .A(n13038), .B(n13046), .S(n12946), .Z(n13034) );
  INV_X1 U15329 ( .A(n13036), .ZN(n13037) );
  INV_X1 U15330 ( .A(n13043), .ZN(n13044) );
  NOR2_X1 U15331 ( .A1(n13045), .A2(n13044), .ZN(n13048) );
  INV_X1 U15332 ( .A(n13046), .ZN(n13047) );
  XNOR2_X1 U15333 ( .A(n13048), .B(n13047), .ZN(n13050) );
  NOR2_X1 U15334 ( .A1(n13054), .A2(n15326), .ZN(n13060) );
  AOI21_X1 U15335 ( .B1(n13319), .B2(n15372), .A(n13060), .ZN(n13056) );
  NAND2_X1 U15336 ( .A1(n13255), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n13055) );
  OAI211_X1 U15337 ( .C1(n13257), .C2(n13249), .A(n13056), .B(n13055), .ZN(
        P3_U3202) );
  NAND2_X1 U15338 ( .A1(n13322), .A2(n13209), .ZN(n13057) );
  OAI211_X1 U15339 ( .C1(n15372), .C2(n13058), .A(n13057), .B(n13056), .ZN(
        P3_U3203) );
  INV_X1 U15340 ( .A(n13059), .ZN(n13066) );
  AOI21_X1 U15341 ( .B1(n13255), .B2(P3_REG2_REG_29__SCAN_IN), .A(n13060), 
        .ZN(n13061) );
  OAI21_X1 U15342 ( .B1(n13062), .B2(n13249), .A(n13061), .ZN(n13063) );
  AOI21_X1 U15343 ( .B1(n13064), .B2(n15323), .A(n13063), .ZN(n13065) );
  OAI21_X1 U15344 ( .B1(n13066), .B2(n13255), .A(n13065), .ZN(P3_U3204) );
  NAND2_X1 U15345 ( .A1(n9196), .A2(n13067), .ZN(n13068) );
  XOR2_X1 U15346 ( .A(n13070), .B(n13068), .Z(n13263) );
  INV_X1 U15347 ( .A(n13263), .ZN(n13079) );
  OAI211_X1 U15348 ( .C1(n13071), .C2(n13070), .A(n13069), .B(n10380), .ZN(
        n13073) );
  AOI22_X1 U15349 ( .A1(n13075), .A2(n15369), .B1(n13255), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n13076) );
  OAI21_X1 U15350 ( .B1(n13328), .B2(n13249), .A(n13076), .ZN(n13077) );
  AOI21_X1 U15351 ( .B1(n13262), .B2(n15372), .A(n13077), .ZN(n13078) );
  OAI21_X1 U15352 ( .B1(n13214), .B2(n13079), .A(n13078), .ZN(P3_U3205) );
  INV_X1 U15353 ( .A(n13080), .ZN(n13087) );
  INV_X1 U15354 ( .A(n13081), .ZN(n15370) );
  AOI22_X1 U15355 ( .A1(n13082), .A2(n15369), .B1(n13255), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13083) );
  OAI21_X1 U15356 ( .B1(n13330), .B2(n13249), .A(n13083), .ZN(n13084) );
  AOI21_X1 U15357 ( .B1(n13085), .B2(n15370), .A(n13084), .ZN(n13086) );
  OAI21_X1 U15358 ( .B1(n13087), .B2(n13255), .A(n13086), .ZN(P3_U3206) );
  INV_X1 U15359 ( .A(n13266), .ZN(n13098) );
  XOR2_X1 U15360 ( .A(n13092), .B(n13091), .Z(n13267) );
  INV_X1 U15361 ( .A(n13093), .ZN(n13334) );
  AOI22_X1 U15362 ( .A1(n13094), .A2(n15369), .B1(n13255), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13095) );
  OAI21_X1 U15363 ( .B1(n13334), .B2(n13249), .A(n13095), .ZN(n13096) );
  AOI21_X1 U15364 ( .B1(n13267), .B2(n15323), .A(n13096), .ZN(n13097) );
  OAI21_X1 U15365 ( .B1(n13098), .B2(n13255), .A(n13097), .ZN(P3_U3207) );
  XNOR2_X1 U15366 ( .A(n13099), .B(n13101), .ZN(n13108) );
  OAI211_X1 U15367 ( .C1(n13102), .C2(n13101), .A(n13100), .B(n10380), .ZN(
        n13106) );
  AOI22_X1 U15368 ( .A1(n13104), .A2(n15358), .B1(n15360), .B2(n13103), .ZN(
        n13105) );
  OAI211_X1 U15369 ( .C1(n13107), .C2(n13108), .A(n13106), .B(n13105), .ZN(
        n13270) );
  INV_X1 U15370 ( .A(n13270), .ZN(n13113) );
  INV_X1 U15371 ( .A(n13108), .ZN(n13271) );
  AOI22_X1 U15372 ( .A1(n13109), .A2(n15369), .B1(n13255), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n13110) );
  OAI21_X1 U15373 ( .B1(n13337), .B2(n13249), .A(n13110), .ZN(n13111) );
  AOI21_X1 U15374 ( .B1(n13271), .B2(n15370), .A(n13111), .ZN(n13112) );
  OAI21_X1 U15375 ( .B1(n13113), .B2(n13255), .A(n13112), .ZN(P3_U3208) );
  AOI21_X1 U15376 ( .B1(n13117), .B2(n13114), .A(n6642), .ZN(n13120) );
  AOI22_X1 U15377 ( .A1(n13115), .A2(n15358), .B1(n15360), .B2(n13141), .ZN(
        n13119) );
  OAI21_X1 U15378 ( .B1(n6679), .B2(n13117), .A(n13116), .ZN(n13274) );
  NAND2_X1 U15379 ( .A1(n13274), .A2(n15363), .ZN(n13118) );
  OAI211_X1 U15380 ( .C1(n13120), .C2(n15366), .A(n13119), .B(n13118), .ZN(
        n13273) );
  INV_X1 U15381 ( .A(n13273), .ZN(n13125) );
  AOI22_X1 U15382 ( .A1(n13121), .A2(n15369), .B1(n13255), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n13122) );
  OAI21_X1 U15383 ( .B1(n13341), .B2(n13249), .A(n13122), .ZN(n13123) );
  AOI21_X1 U15384 ( .B1(n13274), .B2(n15370), .A(n13123), .ZN(n13124) );
  OAI21_X1 U15385 ( .B1(n13125), .B2(n13255), .A(n13124), .ZN(P3_U3209) );
  XNOR2_X1 U15386 ( .A(n13126), .B(n13127), .ZN(n13134) );
  OR2_X1 U15387 ( .A1(n13128), .A2(n13127), .ZN(n13129) );
  AND2_X1 U15388 ( .A1(n13130), .A2(n13129), .ZN(n13278) );
  OAI22_X1 U15389 ( .A1(n13131), .A2(n15300), .B1(n13157), .B2(n15298), .ZN(
        n13132) );
  AOI21_X1 U15390 ( .B1(n13278), .B2(n15363), .A(n13132), .ZN(n13133) );
  OAI21_X1 U15391 ( .B1(n15366), .B2(n13134), .A(n13133), .ZN(n13277) );
  NAND2_X1 U15392 ( .A1(n13278), .A2(n15370), .ZN(n13137) );
  AOI22_X1 U15393 ( .A1(n13135), .A2(n15369), .B1(n13255), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n13136) );
  OAI211_X1 U15394 ( .C1(n13345), .C2(n13249), .A(n13137), .B(n13136), .ZN(
        n13138) );
  AOI21_X1 U15395 ( .B1(n13277), .B2(n15372), .A(n13138), .ZN(n13139) );
  INV_X1 U15396 ( .A(n13139), .ZN(P3_U3210) );
  XNOR2_X1 U15397 ( .A(n13140), .B(n13144), .ZN(n13142) );
  AOI222_X1 U15398 ( .A1(n10380), .A2(n13142), .B1(n13141), .B2(n15358), .C1(
        n13171), .C2(n15360), .ZN(n13283) );
  XOR2_X1 U15399 ( .A(n13144), .B(n13143), .Z(n13281) );
  AOI22_X1 U15400 ( .A1(n13145), .A2(n15369), .B1(P3_REG2_REG_22__SCAN_IN), 
        .B2(n13255), .ZN(n13146) );
  OAI21_X1 U15401 ( .B1(n13147), .B2(n13249), .A(n13146), .ZN(n13148) );
  AOI21_X1 U15402 ( .B1(n13281), .B2(n15323), .A(n13148), .ZN(n13149) );
  OAI21_X1 U15403 ( .B1(n13283), .B2(n13255), .A(n13149), .ZN(P3_U3211) );
  INV_X1 U15404 ( .A(n13150), .ZN(n13154) );
  INV_X1 U15405 ( .A(n13151), .ZN(n13166) );
  OR2_X1 U15406 ( .A1(n13152), .A2(n13166), .ZN(n13153) );
  OAI211_X1 U15407 ( .C1(n13155), .C2(n13154), .A(n10380), .B(n13153), .ZN(
        n13160) );
  OAI22_X1 U15408 ( .A1(n13157), .A2(n15300), .B1(n13156), .B2(n15298), .ZN(
        n13158) );
  INV_X1 U15409 ( .A(n13158), .ZN(n13159) );
  INV_X1 U15410 ( .A(n13161), .ZN(n13163) );
  OAI22_X1 U15411 ( .A1(n13163), .A2(n15326), .B1(n13162), .B2(n15372), .ZN(
        n13164) );
  AOI21_X1 U15412 ( .B1(n13349), .B2(n13209), .A(n13164), .ZN(n13168) );
  XNOR2_X1 U15413 ( .A(n13165), .B(n13166), .ZN(n13284) );
  NAND2_X1 U15414 ( .A1(n13284), .A2(n15323), .ZN(n13167) );
  OAI211_X1 U15415 ( .C1(n13286), .C2(n13255), .A(n13168), .B(n13167), .ZN(
        P3_U3212) );
  XNOR2_X1 U15416 ( .A(n13169), .B(n13170), .ZN(n13173) );
  AOI222_X1 U15417 ( .A1(n10380), .A2(n13173), .B1(n13172), .B2(n15360), .C1(
        n13171), .C2(n15358), .ZN(n13292) );
  AOI21_X1 U15418 ( .B1(n13175), .B2(n13174), .A(n6708), .ZN(n13291) );
  AOI22_X1 U15419 ( .A1(n13255), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n13176), 
        .B2(n15369), .ZN(n13177) );
  OAI21_X1 U15420 ( .B1(n13178), .B2(n13249), .A(n13177), .ZN(n13179) );
  AOI21_X1 U15421 ( .B1(n13291), .B2(n15323), .A(n13179), .ZN(n13180) );
  OAI21_X1 U15422 ( .B1(n13292), .B2(n13255), .A(n13180), .ZN(P3_U3213) );
  XNOR2_X1 U15423 ( .A(n13181), .B(n13184), .ZN(n13295) );
  INV_X1 U15424 ( .A(n13295), .ZN(n13194) );
  INV_X1 U15425 ( .A(n13182), .ZN(n13185) );
  OAI211_X1 U15426 ( .C1(n13185), .C2(n13184), .A(n10380), .B(n13183), .ZN(
        n13189) );
  AOI22_X1 U15427 ( .A1(n13187), .A2(n15358), .B1(n15360), .B2(n13186), .ZN(
        n13188) );
  NAND2_X1 U15428 ( .A1(n13189), .A2(n13188), .ZN(n13294) );
  AOI22_X1 U15429 ( .A1(n13255), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15369), 
        .B2(n13190), .ZN(n13191) );
  OAI21_X1 U15430 ( .B1(n13355), .B2(n13249), .A(n13191), .ZN(n13192) );
  AOI21_X1 U15431 ( .B1(n13294), .B2(n15372), .A(n13192), .ZN(n13193) );
  OAI21_X1 U15432 ( .B1(n13214), .B2(n13194), .A(n13193), .ZN(P3_U3214) );
  NAND2_X1 U15433 ( .A1(n13196), .A2(n13195), .ZN(n13197) );
  INV_X1 U15434 ( .A(n13299), .ZN(n13213) );
  INV_X1 U15435 ( .A(n13199), .ZN(n13200) );
  AOI21_X1 U15436 ( .B1(n13202), .B2(n13201), .A(n13200), .ZN(n13203) );
  OAI222_X1 U15437 ( .A1(n15300), .A2(n13204), .B1(n15298), .B2(n13232), .C1(
        n15366), .C2(n13203), .ZN(n13298) );
  NAND2_X1 U15438 ( .A1(n13298), .A2(n15372), .ZN(n13212) );
  INV_X1 U15439 ( .A(n13205), .ZN(n13206) );
  OAI22_X1 U15440 ( .A1(n15372), .A2(n13207), .B1(n13206), .B2(n15326), .ZN(
        n13208) );
  AOI21_X1 U15441 ( .B1(n13210), .B2(n13209), .A(n13208), .ZN(n13211) );
  OAI211_X1 U15442 ( .C1(n13214), .C2(n13213), .A(n13212), .B(n13211), .ZN(
        P3_U3215) );
  XNOR2_X1 U15443 ( .A(n13216), .B(n13215), .ZN(n13217) );
  OAI222_X1 U15444 ( .A1(n15300), .A2(n13218), .B1(n15298), .B2(n13245), .C1(
        n13217), .C2(n15366), .ZN(n13302) );
  INV_X1 U15445 ( .A(n13302), .ZN(n13227) );
  OAI21_X1 U15446 ( .B1(n13221), .B2(n13220), .A(n13219), .ZN(n13303) );
  NOR2_X1 U15447 ( .A1(n13363), .A2(n13249), .ZN(n13225) );
  INV_X1 U15448 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13223) );
  OAI22_X1 U15449 ( .A1(n15372), .A2(n13223), .B1(n13222), .B2(n15326), .ZN(
        n13224) );
  AOI211_X1 U15450 ( .C1(n13303), .C2(n15323), .A(n13225), .B(n13224), .ZN(
        n13226) );
  OAI21_X1 U15451 ( .B1(n13227), .B2(n13255), .A(n13226), .ZN(P3_U3216) );
  XNOR2_X1 U15452 ( .A(n13228), .B(n13229), .ZN(n13230) );
  OAI222_X1 U15453 ( .A1(n15300), .A2(n13232), .B1(n15298), .B2(n13231), .C1(
        n13230), .C2(n15366), .ZN(n13306) );
  INV_X1 U15454 ( .A(n13306), .ZN(n13241) );
  OAI21_X1 U15455 ( .B1(n13235), .B2(n13234), .A(n13233), .ZN(n13307) );
  NOR2_X1 U15456 ( .A1(n13367), .A2(n13249), .ZN(n13239) );
  OAI22_X1 U15457 ( .A1(n15372), .A2(n13237), .B1(n13236), .B2(n15326), .ZN(
        n13238) );
  AOI211_X1 U15458 ( .C1(n13307), .C2(n15323), .A(n13239), .B(n13238), .ZN(
        n13240) );
  OAI21_X1 U15459 ( .B1(n13241), .B2(n13255), .A(n13240), .ZN(P3_U3217) );
  XOR2_X1 U15460 ( .A(n13242), .B(n13246), .Z(n13243) );
  OAI222_X1 U15461 ( .A1(n15300), .A2(n13245), .B1(n15298), .B2(n13244), .C1(
        n13243), .C2(n15366), .ZN(n13310) );
  INV_X1 U15462 ( .A(n13310), .ZN(n13256) );
  XNOR2_X1 U15463 ( .A(n13247), .B(n13246), .ZN(n13311) );
  INV_X1 U15464 ( .A(n13248), .ZN(n13371) );
  NOR2_X1 U15465 ( .A1(n13371), .A2(n13249), .ZN(n13253) );
  OAI22_X1 U15466 ( .A1(n15372), .A2(n13251), .B1(n13250), .B2(n15326), .ZN(
        n13252) );
  AOI211_X1 U15467 ( .C1(n13311), .C2(n15323), .A(n13253), .B(n13252), .ZN(
        n13254) );
  OAI21_X1 U15468 ( .B1(n13256), .B2(n13255), .A(n13254), .ZN(P3_U3218) );
  INV_X1 U15469 ( .A(n13257), .ZN(n13318) );
  NAND2_X1 U15470 ( .A1(n13318), .A2(n9187), .ZN(n13258) );
  NAND2_X1 U15471 ( .A1(n13319), .A2(n15419), .ZN(n13260) );
  OAI211_X1 U15472 ( .C1(n15419), .C2(n9217), .A(n13258), .B(n13260), .ZN(
        P3_U3490) );
  NAND2_X1 U15473 ( .A1(n15417), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n13259) );
  OAI211_X1 U15474 ( .C1(n13261), .C2(n13317), .A(n13260), .B(n13259), .ZN(
        P3_U3489) );
  INV_X1 U15475 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13264) );
  OAI21_X1 U15476 ( .B1(n13328), .B2(n13317), .A(n13265), .ZN(P3_U3487) );
  INV_X1 U15477 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13268) );
  AOI21_X1 U15478 ( .B1(n15405), .B2(n13267), .A(n13266), .ZN(n13331) );
  MUX2_X1 U15479 ( .A(n13268), .B(n13331), .S(n15419), .Z(n13269) );
  OAI21_X1 U15480 ( .B1(n13334), .B2(n13317), .A(n13269), .ZN(P3_U3485) );
  AOI21_X1 U15481 ( .B1(n15381), .B2(n13271), .A(n13270), .ZN(n13335) );
  MUX2_X1 U15482 ( .A(n15621), .B(n13335), .S(n15419), .Z(n13272) );
  OAI21_X1 U15483 ( .B1(n13337), .B2(n13317), .A(n13272), .ZN(P3_U3484) );
  INV_X1 U15484 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13275) );
  AOI21_X1 U15485 ( .B1(n15381), .B2(n13274), .A(n13273), .ZN(n13338) );
  MUX2_X1 U15486 ( .A(n13275), .B(n13338), .S(n15419), .Z(n13276) );
  OAI21_X1 U15487 ( .B1(n13341), .B2(n13317), .A(n13276), .ZN(P3_U3483) );
  AOI21_X1 U15488 ( .B1(n15381), .B2(n13278), .A(n13277), .ZN(n13342) );
  MUX2_X1 U15489 ( .A(n15481), .B(n13342), .S(n15419), .Z(n13279) );
  OAI21_X1 U15490 ( .B1(n13345), .B2(n13317), .A(n13279), .ZN(P3_U3482) );
  AOI22_X1 U15491 ( .A1(n13281), .A2(n15405), .B1(n13290), .B2(n13280), .ZN(
        n13282) );
  NAND2_X1 U15492 ( .A1(n13283), .A2(n13282), .ZN(n13346) );
  MUX2_X1 U15493 ( .A(P3_REG1_REG_22__SCAN_IN), .B(n13346), .S(n15419), .Z(
        P3_U3481) );
  NAND2_X1 U15494 ( .A1(n13284), .A2(n15405), .ZN(n13285) );
  NAND2_X1 U15495 ( .A1(n13286), .A2(n13285), .ZN(n13347) );
  MUX2_X1 U15496 ( .A(P3_REG1_REG_21__SCAN_IN), .B(n13347), .S(n15419), .Z(
        n13287) );
  AOI21_X1 U15497 ( .B1(n9187), .B2(n13349), .A(n13287), .ZN(n13288) );
  INV_X1 U15498 ( .A(n13288), .ZN(P3_U3480) );
  AOI22_X1 U15499 ( .A1(n13291), .A2(n15405), .B1(n13290), .B2(n13289), .ZN(
        n13293) );
  NAND2_X1 U15500 ( .A1(n13293), .A2(n13292), .ZN(n13351) );
  MUX2_X1 U15501 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n13351), .S(n15419), .Z(
        P3_U3479) );
  AOI21_X1 U15502 ( .B1(n15405), .B2(n13295), .A(n13294), .ZN(n13352) );
  MUX2_X1 U15503 ( .A(n13296), .B(n13352), .S(n15419), .Z(n13297) );
  OAI21_X1 U15504 ( .B1(n13317), .B2(n13355), .A(n13297), .ZN(P3_U3478) );
  AOI21_X1 U15505 ( .B1(n13299), .B2(n15405), .A(n13298), .ZN(n13356) );
  MUX2_X1 U15506 ( .A(n13300), .B(n13356), .S(n15419), .Z(n13301) );
  OAI21_X1 U15507 ( .B1(n13359), .B2(n13317), .A(n13301), .ZN(P3_U3477) );
  AOI21_X1 U15508 ( .B1(n15405), .B2(n13303), .A(n13302), .ZN(n13360) );
  MUX2_X1 U15509 ( .A(n13304), .B(n13360), .S(n15419), .Z(n13305) );
  OAI21_X1 U15510 ( .B1(n13363), .B2(n13317), .A(n13305), .ZN(P3_U3476) );
  INV_X1 U15511 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13308) );
  AOI21_X1 U15512 ( .B1(n15405), .B2(n13307), .A(n13306), .ZN(n13364) );
  MUX2_X1 U15513 ( .A(n13308), .B(n13364), .S(n15419), .Z(n13309) );
  OAI21_X1 U15514 ( .B1(n13367), .B2(n13317), .A(n13309), .ZN(P3_U3475) );
  AOI21_X1 U15515 ( .B1(n13311), .B2(n15405), .A(n13310), .ZN(n13368) );
  MUX2_X1 U15516 ( .A(n15480), .B(n13368), .S(n15419), .Z(n13312) );
  OAI21_X1 U15517 ( .B1(n13371), .B2(n13317), .A(n13312), .ZN(P3_U3474) );
  AOI21_X1 U15518 ( .B1(n15405), .B2(n13314), .A(n13313), .ZN(n13372) );
  MUX2_X1 U15519 ( .A(n13315), .B(n13372), .S(n15419), .Z(n13316) );
  OAI21_X1 U15520 ( .B1(n13317), .B2(n13375), .A(n13316), .ZN(P3_U3473) );
  INV_X1 U15521 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n13321) );
  NAND2_X1 U15522 ( .A1(n13318), .A2(n10411), .ZN(n13320) );
  NAND2_X1 U15523 ( .A1(n13319), .A2(n15407), .ZN(n13323) );
  OAI211_X1 U15524 ( .C1(n13321), .C2(n15407), .A(n13320), .B(n13323), .ZN(
        P3_U3458) );
  INV_X1 U15525 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n13325) );
  NAND2_X1 U15526 ( .A1(n13322), .A2(n10411), .ZN(n13324) );
  OAI211_X1 U15527 ( .C1(n13325), .C2(n15407), .A(n13324), .B(n13323), .ZN(
        P3_U3457) );
  INV_X1 U15528 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13327) );
  INV_X1 U15529 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13332) );
  MUX2_X1 U15530 ( .A(n13332), .B(n13331), .S(n15407), .Z(n13333) );
  OAI21_X1 U15531 ( .B1(n13334), .B2(n13376), .A(n13333), .ZN(P3_U3453) );
  MUX2_X1 U15532 ( .A(n15613), .B(n13335), .S(n15407), .Z(n13336) );
  OAI21_X1 U15533 ( .B1(n13337), .B2(n13376), .A(n13336), .ZN(P3_U3452) );
  INV_X1 U15534 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13339) );
  MUX2_X1 U15535 ( .A(n13339), .B(n13338), .S(n15407), .Z(n13340) );
  OAI21_X1 U15536 ( .B1(n13341), .B2(n13376), .A(n13340), .ZN(P3_U3451) );
  INV_X1 U15537 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13343) );
  MUX2_X1 U15538 ( .A(n13343), .B(n13342), .S(n15407), .Z(n13344) );
  OAI21_X1 U15539 ( .B1(n13345), .B2(n13376), .A(n13344), .ZN(P3_U3450) );
  MUX2_X1 U15540 ( .A(P3_REG0_REG_22__SCAN_IN), .B(n13346), .S(n15407), .Z(
        P3_U3449) );
  MUX2_X1 U15541 ( .A(n13347), .B(P3_REG0_REG_21__SCAN_IN), .S(n15409), .Z(
        n13348) );
  AOI21_X1 U15542 ( .B1(n10411), .B2(n13349), .A(n13348), .ZN(n13350) );
  INV_X1 U15543 ( .A(n13350), .ZN(P3_U3448) );
  MUX2_X1 U15544 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n13351), .S(n15407), .Z(
        P3_U3447) );
  MUX2_X1 U15545 ( .A(n13353), .B(n13352), .S(n15407), .Z(n13354) );
  OAI21_X1 U15546 ( .B1(n13376), .B2(n13355), .A(n13354), .ZN(P3_U3446) );
  MUX2_X1 U15547 ( .A(n13357), .B(n13356), .S(n15407), .Z(n13358) );
  OAI21_X1 U15548 ( .B1(n13359), .B2(n13376), .A(n13358), .ZN(P3_U3444) );
  MUX2_X1 U15549 ( .A(n13361), .B(n13360), .S(n15407), .Z(n13362) );
  OAI21_X1 U15550 ( .B1(n13363), .B2(n13376), .A(n13362), .ZN(P3_U3441) );
  MUX2_X1 U15551 ( .A(n13365), .B(n13364), .S(n15407), .Z(n13366) );
  OAI21_X1 U15552 ( .B1(n13367), .B2(n13376), .A(n13366), .ZN(P3_U3438) );
  INV_X1 U15553 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13369) );
  MUX2_X1 U15554 ( .A(n13369), .B(n13368), .S(n15407), .Z(n13370) );
  OAI21_X1 U15555 ( .B1(n13371), .B2(n13376), .A(n13370), .ZN(P3_U3435) );
  MUX2_X1 U15556 ( .A(n13373), .B(n13372), .S(n15407), .Z(n13374) );
  OAI21_X1 U15557 ( .B1(n13376), .B2(n13375), .A(n13374), .ZN(P3_U3432) );
  MUX2_X1 U15558 ( .A(n13377), .B(P3_D_REG_1__SCAN_IN), .S(n13378), .Z(
        P3_U3377) );
  MUX2_X1 U15559 ( .A(n13379), .B(P3_D_REG_0__SCAN_IN), .S(n13378), .Z(
        P3_U3376) );
  NAND3_X1 U15560 ( .A1(n13380), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n13384) );
  NAND2_X1 U15561 ( .A1(n13381), .A2(n14762), .ZN(n13383) );
  NAND2_X1 U15562 ( .A1(n14761), .A2(SI_31_), .ZN(n13382) );
  OAI211_X1 U15563 ( .C1(n13385), .C2(n13384), .A(n13383), .B(n13382), .ZN(
        P3_U3264) );
  INV_X1 U15564 ( .A(n13386), .ZN(n13387) );
  OAI222_X1 U15565 ( .A1(n14741), .A2(n13389), .B1(P3_U3151), .B2(n13388), 
        .C1(n14743), .C2(n13387), .ZN(P3_U3266) );
  NAND2_X1 U15566 ( .A1(n13849), .A2(n13506), .ZN(n13395) );
  OR2_X1 U15567 ( .A1(n13424), .A2(n13425), .ZN(n13393) );
  NAND2_X1 U15568 ( .A1(n13512), .A2(n13816), .ZN(n13392) );
  NAND2_X1 U15569 ( .A1(n13393), .A2(n13392), .ZN(n13623) );
  AOI22_X1 U15570 ( .A1(n14845), .A2(n13623), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13394) );
  OAI211_X1 U15571 ( .C1(n15124), .C2(n13629), .A(n13395), .B(n13394), .ZN(
        n13396) );
  INV_X1 U15572 ( .A(n13397), .ZN(n13399) );
  OAI22_X1 U15573 ( .A1(n13399), .A2(n13481), .B1(n13398), .B2(n13488), .ZN(
        n13404) );
  AOI22_X1 U15574 ( .A1(n15115), .A2(n13685), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13401) );
  AOI22_X1 U15575 ( .A1(n15113), .A2(n13684), .B1(n13440), .B2(n13694), .ZN(
        n13400) );
  OAI211_X1 U15576 ( .C1(n7784), .C2(n15117), .A(n13401), .B(n13400), .ZN(
        n13402) );
  AOI21_X1 U15577 ( .B1(n13404), .B2(n13403), .A(n13402), .ZN(n13405) );
  INV_X1 U15578 ( .A(n13405), .ZN(P2_U3188) );
  OAI21_X1 U15579 ( .B1(n13408), .B2(n13407), .A(n13406), .ZN(n13409) );
  NAND2_X1 U15580 ( .A1(n13409), .A2(n15120), .ZN(n13413) );
  INV_X1 U15581 ( .A(n13410), .ZN(n13755) );
  AOI22_X1 U15582 ( .A1(n13514), .A2(n13816), .B1(n13814), .B2(n13515), .ZN(
        n13753) );
  NAND2_X1 U15583 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13591)
         );
  OAI21_X1 U15584 ( .B1(n13477), .B2(n13753), .A(n13591), .ZN(n13411) );
  AOI21_X1 U15585 ( .B1(n13755), .B2(n13440), .A(n13411), .ZN(n13412) );
  OAI211_X1 U15586 ( .C1(n13750), .C2(n15117), .A(n13413), .B(n13412), .ZN(
        P2_U3191) );
  OAI211_X1 U15587 ( .C1(n13416), .C2(n13415), .A(n13414), .B(n15120), .ZN(
        n13422) );
  OAI22_X1 U15588 ( .A1(n13418), .A2(n13423), .B1(n13417), .B2(n13425), .ZN(
        n13716) );
  AOI22_X1 U15589 ( .A1(n13716), .A2(n14845), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13419) );
  OAI21_X1 U15590 ( .B1(n13720), .B2(n15124), .A(n13419), .ZN(n13420) );
  AOI21_X1 U15591 ( .B1(n13879), .B2(n13506), .A(n13420), .ZN(n13421) );
  NAND2_X1 U15592 ( .A1(n13422), .A2(n13421), .ZN(P2_U3195) );
  OAI22_X1 U15593 ( .A1(n13426), .A2(n13425), .B1(n13424), .B2(n13423), .ZN(
        n13655) );
  AOI22_X1 U15594 ( .A1(n14845), .A2(n13655), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13427) );
  OAI21_X1 U15595 ( .B1(n13657), .B2(n15124), .A(n13427), .ZN(n13435) );
  INV_X1 U15596 ( .A(n13428), .ZN(n13429) );
  NAND3_X1 U15597 ( .A1(n13429), .A2(n13496), .A3(n13685), .ZN(n13433) );
  OAI21_X1 U15598 ( .B1(n13453), .B2(n13430), .A(n15120), .ZN(n13432) );
  INV_X1 U15599 ( .A(n13484), .ZN(n13431) );
  AOI21_X1 U15600 ( .B1(n13433), .B2(n13432), .A(n13431), .ZN(n13434) );
  AOI211_X1 U15601 ( .C1(n13860), .C2(n13506), .A(n13435), .B(n13434), .ZN(
        n13436) );
  INV_X1 U15602 ( .A(n13436), .ZN(P2_U3197) );
  AOI21_X1 U15603 ( .B1(n13439), .B2(n13438), .A(n13437), .ZN(n13445) );
  NAND2_X1 U15604 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n15181)
         );
  AOI22_X1 U15605 ( .A1(n15113), .A2(n13796), .B1(n13440), .B2(n13804), .ZN(
        n13441) );
  OAI211_X1 U15606 ( .C1(n13503), .C2(n13442), .A(n15181), .B(n13441), .ZN(
        n13443) );
  AOI21_X1 U15607 ( .B1(n13907), .B2(n14848), .A(n13443), .ZN(n13444) );
  OAI21_X1 U15608 ( .B1(n13445), .B2(n13481), .A(n13444), .ZN(P2_U3198) );
  AOI21_X1 U15609 ( .B1(n13448), .B2(n13447), .A(n13446), .ZN(n13452) );
  NOR2_X1 U15610 ( .A1(n15124), .A2(n13785), .ZN(n13450) );
  AOI22_X1 U15611 ( .A1(n13515), .A2(n13816), .B1(n13814), .B2(n13817), .ZN(
        n13778) );
  NAND2_X1 U15612 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n15194)
         );
  OAI21_X1 U15613 ( .B1(n13477), .B2(n13778), .A(n15194), .ZN(n13449) );
  AOI211_X1 U15614 ( .C1(n13903), .C2(n14848), .A(n13450), .B(n13449), .ZN(
        n13451) );
  OAI21_X1 U15615 ( .B1(n13452), .B2(n13481), .A(n13451), .ZN(P2_U3200) );
  INV_X1 U15616 ( .A(n13453), .ZN(n13454) );
  OAI211_X1 U15617 ( .C1(n13456), .C2(n13455), .A(n13454), .B(n15120), .ZN(
        n13461) );
  NOR2_X1 U15618 ( .A1(n15124), .A2(n13674), .ZN(n13459) );
  INV_X1 U15619 ( .A(n13668), .ZN(n13457) );
  INV_X1 U15620 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n15639) );
  OAI22_X1 U15621 ( .A1(n13503), .A2(n13457), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15639), .ZN(n13458) );
  AOI211_X1 U15622 ( .C1(n15113), .C2(n13669), .A(n13459), .B(n13458), .ZN(
        n13460) );
  OAI211_X1 U15623 ( .C1(n13677), .C2(n15117), .A(n13461), .B(n13460), .ZN(
        P2_U3201) );
  INV_X1 U15624 ( .A(n13462), .ZN(n13464) );
  NAND2_X1 U15625 ( .A1(n13464), .A2(n13463), .ZN(n13465) );
  XNOR2_X1 U15626 ( .A(n13466), .B(n13465), .ZN(n13473) );
  INV_X1 U15627 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13467) );
  OAI22_X1 U15628 ( .A1(n13501), .A2(n13468), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13467), .ZN(n13471) );
  OAI22_X1 U15629 ( .A1(n13503), .A2(n13469), .B1(n15124), .B2(n13737), .ZN(
        n13470) );
  AOI211_X1 U15630 ( .C1(n13887), .C2(n14848), .A(n13471), .B(n13470), .ZN(
        n13472) );
  OAI21_X1 U15631 ( .B1(n13473), .B2(n13481), .A(n13472), .ZN(P2_U3205) );
  XNOR2_X1 U15632 ( .A(n13475), .B(n13474), .ZN(n13482) );
  NOR2_X1 U15633 ( .A1(n15124), .A2(n13768), .ZN(n13479) );
  AND2_X1 U15634 ( .A1(n13797), .A2(n13814), .ZN(n13476) );
  AOI21_X1 U15635 ( .B1(n13741), .B2(n13816), .A(n13476), .ZN(n13763) );
  NAND2_X1 U15636 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13560)
         );
  OAI21_X1 U15637 ( .B1(n13477), .B2(n13763), .A(n13560), .ZN(n13478) );
  AOI211_X1 U15638 ( .C1(n13898), .C2(n14848), .A(n13479), .B(n13478), .ZN(
        n13480) );
  OAI21_X1 U15639 ( .B1(n13482), .B2(n13481), .A(n13480), .ZN(P2_U3210) );
  OAI21_X1 U15640 ( .B1(n13490), .B2(n13484), .A(n13483), .ZN(n13485) );
  NAND2_X1 U15641 ( .A1(n13485), .A2(n15120), .ZN(n13494) );
  AOI22_X1 U15642 ( .A1(n15115), .A2(n13637), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13486) );
  OAI21_X1 U15643 ( .B1(n13641), .B2(n15124), .A(n13486), .ZN(n13487) );
  AOI21_X1 U15644 ( .B1(n13855), .B2(n14848), .A(n13487), .ZN(n13493) );
  NOR3_X1 U15645 ( .A1(n13490), .A2(n13489), .A3(n13488), .ZN(n13491) );
  OAI21_X1 U15646 ( .B1(n13491), .B2(n15113), .A(n13668), .ZN(n13492) );
  NAND3_X1 U15647 ( .A1(n13494), .A2(n13493), .A3(n13492), .ZN(P2_U3212) );
  NAND2_X1 U15648 ( .A1(n15120), .A2(n13495), .ZN(n13499) );
  NAND2_X1 U15649 ( .A1(n13496), .A2(n13796), .ZN(n13498) );
  MUX2_X1 U15650 ( .A(n13499), .B(n13498), .S(n13497), .Z(n13508) );
  OAI22_X1 U15651 ( .A1(n13501), .A2(n13500), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8375), .ZN(n13505) );
  OAI22_X1 U15652 ( .A1(n13503), .A2(n13502), .B1(n15124), .B2(n13824), .ZN(
        n13504) );
  AOI211_X1 U15653 ( .C1(n13912), .C2(n13506), .A(n13505), .B(n13504), .ZN(
        n13507) );
  NAND2_X1 U15654 ( .A1(n13508), .A2(n13507), .ZN(P2_U3213) );
  INV_X2 U15655 ( .A(P2_U3947), .ZN(n13526) );
  MUX2_X1 U15656 ( .A(n13509), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13526), .Z(
        P2_U3562) );
  MUX2_X1 U15657 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13510), .S(P2_U3947), .Z(
        P2_U3561) );
  MUX2_X1 U15658 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13511), .S(P2_U3947), .Z(
        P2_U3560) );
  MUX2_X1 U15659 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13512), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U15660 ( .A(n13637), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13526), .Z(
        P2_U3558) );
  MUX2_X1 U15661 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13513), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U15662 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13668), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U15663 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13685), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15664 ( .A(n13669), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13526), .Z(
        P2_U3554) );
  MUX2_X1 U15665 ( .A(n13684), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13526), .Z(
        P2_U3553) );
  MUX2_X1 U15666 ( .A(n13742), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13526), .Z(
        P2_U3552) );
  MUX2_X1 U15667 ( .A(n13514), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13526), .Z(
        P2_U3551) );
  MUX2_X1 U15668 ( .A(n13741), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13526), .Z(
        P2_U3550) );
  MUX2_X1 U15669 ( .A(n13515), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13526), .Z(
        P2_U3549) );
  MUX2_X1 U15670 ( .A(n13797), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13526), .Z(
        P2_U3548) );
  MUX2_X1 U15671 ( .A(n13817), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13526), .Z(
        P2_U3547) );
  MUX2_X1 U15672 ( .A(n13796), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13526), .Z(
        P2_U3546) );
  MUX2_X1 U15673 ( .A(n13815), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13526), .Z(
        P2_U3545) );
  MUX2_X1 U15674 ( .A(n13516), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13526), .Z(
        P2_U3543) );
  MUX2_X1 U15675 ( .A(n15112), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13526), .Z(
        P2_U3542) );
  MUX2_X1 U15676 ( .A(n13517), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13526), .Z(
        P2_U3541) );
  MUX2_X1 U15677 ( .A(n13518), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13526), .Z(
        P2_U3540) );
  MUX2_X1 U15678 ( .A(n13519), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13526), .Z(
        P2_U3539) );
  MUX2_X1 U15679 ( .A(n13520), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13526), .Z(
        P2_U3538) );
  MUX2_X1 U15680 ( .A(n13521), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13526), .Z(
        P2_U3537) );
  MUX2_X1 U15681 ( .A(n13522), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13526), .Z(
        P2_U3536) );
  MUX2_X1 U15682 ( .A(n13523), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13526), .Z(
        P2_U3535) );
  MUX2_X1 U15683 ( .A(n13524), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13526), .Z(
        P2_U3534) );
  MUX2_X1 U15684 ( .A(n13525), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13526), .Z(
        P2_U3533) );
  MUX2_X1 U15685 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n13527), .S(P2_U3947), .Z(
        P2_U3531) );
  INV_X1 U15686 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n13529) );
  OAI22_X1 U15687 ( .A1(n15166), .A2(n13529), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13528), .ZN(n13530) );
  AOI21_X1 U15688 ( .B1(n13531), .B2(n15168), .A(n13530), .ZN(n13544) );
  MUX2_X1 U15689 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n8117), .S(n13532), .Z(
        n13533) );
  OAI21_X1 U15690 ( .B1(n10620), .B2(n13534), .A(n13533), .ZN(n13535) );
  NAND3_X1 U15691 ( .A1(n15190), .A2(n13536), .A3(n13535), .ZN(n13543) );
  INV_X1 U15692 ( .A(n13537), .ZN(n13541) );
  AND2_X1 U15693 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n13540) );
  INV_X1 U15694 ( .A(n13538), .ZN(n13539) );
  OAI211_X1 U15695 ( .C1(n13541), .C2(n13540), .A(n15198), .B(n13539), .ZN(
        n13542) );
  NAND3_X1 U15696 ( .A1(n13544), .A2(n13543), .A3(n13542), .ZN(P2_U3215) );
  NAND2_X1 U15697 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n13545), .ZN(n13558) );
  INV_X1 U15698 ( .A(n13558), .ZN(n13546) );
  AOI21_X1 U15699 ( .B1(n13786), .B2(n15203), .A(n13546), .ZN(n15199) );
  NAND2_X1 U15700 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n13547), .ZN(n13557) );
  INV_X1 U15701 ( .A(n13557), .ZN(n13548) );
  AOI21_X1 U15702 ( .B1(n8396), .B2(n15188), .A(n13548), .ZN(n15184) );
  NAND2_X1 U15703 ( .A1(n13563), .A2(n13549), .ZN(n15126) );
  MUX2_X1 U15704 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n13550), .S(n15135), .Z(
        n15127) );
  AOI21_X1 U15705 ( .B1(n15128), .B2(n15126), .A(n15127), .ZN(n15125) );
  AOI21_X1 U15706 ( .B1(n13550), .B2(n15135), .A(n15125), .ZN(n15147) );
  MUX2_X1 U15707 ( .A(n13551), .B(P2_REG2_REG_13__SCAN_IN), .S(n15148), .Z(
        n15146) );
  NAND2_X1 U15708 ( .A1(n13552), .A2(n13553), .ZN(n13554) );
  NAND2_X1 U15709 ( .A1(n13554), .A2(n15160), .ZN(n13555) );
  NAND2_X1 U15710 ( .A1(n15169), .A2(n13555), .ZN(n13556) );
  NAND2_X1 U15711 ( .A1(n13557), .A2(n15183), .ZN(n15200) );
  NAND2_X1 U15712 ( .A1(n15199), .A2(n15200), .ZN(n15197) );
  NAND2_X1 U15713 ( .A1(n13558), .A2(n15197), .ZN(n13578) );
  AOI21_X1 U15714 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n13559), .A(n13579), 
        .ZN(n13577) );
  OAI21_X1 U15715 ( .B1(n15204), .B2(n13561), .A(n13560), .ZN(n13575) );
  XNOR2_X1 U15716 ( .A(n15203), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15192) );
  INV_X1 U15717 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n13570) );
  XNOR2_X1 U15718 ( .A(n15188), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n15178) );
  XNOR2_X1 U15719 ( .A(n15164), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n15155) );
  OAI21_X1 U15720 ( .B1(n11041), .B2(n13563), .A(n13562), .ZN(n15133) );
  MUX2_X1 U15721 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n13564), .S(n15135), .Z(
        n15134) );
  NOR2_X1 U15722 ( .A1(n15133), .A2(n15134), .ZN(n15132) );
  AOI21_X1 U15723 ( .B1(n13564), .B2(n15135), .A(n15132), .ZN(n15144) );
  MUX2_X1 U15724 ( .A(n13565), .B(P2_REG1_REG_13__SCAN_IN), .S(n15148), .Z(
        n15143) );
  NAND2_X1 U15725 ( .A1(n15144), .A2(n15143), .ZN(n15142) );
  OAI21_X1 U15726 ( .B1(n13565), .B2(n15148), .A(n15142), .ZN(n15156) );
  NAND2_X1 U15727 ( .A1(n15155), .A2(n15156), .ZN(n15154) );
  OAI21_X1 U15728 ( .B1(n15164), .B2(n13566), .A(n15154), .ZN(n13567) );
  NAND2_X1 U15729 ( .A1(n15169), .A2(n13567), .ZN(n13569) );
  XNOR2_X1 U15730 ( .A(n13568), .B(n13567), .ZN(n15173) );
  NAND2_X1 U15731 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n15173), .ZN(n15172) );
  NAND2_X1 U15732 ( .A1(n13569), .A2(n15172), .ZN(n15179) );
  NAND2_X1 U15733 ( .A1(n15178), .A2(n15179), .ZN(n15177) );
  OAI21_X1 U15734 ( .B1(n15188), .B2(n13570), .A(n15177), .ZN(n15191) );
  NAND2_X1 U15735 ( .A1(n15192), .A2(n15191), .ZN(n15189) );
  OAI21_X1 U15736 ( .B1(n15203), .B2(n13571), .A(n15189), .ZN(n13580) );
  XOR2_X1 U15737 ( .A(n13580), .B(n13581), .Z(n13572) );
  NAND2_X1 U15738 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n13572), .ZN(n13583) );
  OAI211_X1 U15739 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n13572), .A(n15190), 
        .B(n13583), .ZN(n13573) );
  INV_X1 U15740 ( .A(n13573), .ZN(n13574) );
  AOI211_X1 U15741 ( .C1(n15196), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n13575), 
        .B(n13574), .ZN(n13576) );
  OAI21_X1 U15742 ( .B1(n13577), .B2(n15129), .A(n13576), .ZN(P2_U3232) );
  INV_X1 U15743 ( .A(n13588), .ZN(n13586) );
  NAND2_X1 U15744 ( .A1(n13581), .A2(n13580), .ZN(n13582) );
  NAND2_X1 U15745 ( .A1(n13583), .A2(n13582), .ZN(n13584) );
  XOR2_X1 U15746 ( .A(n13584), .B(P2_REG1_REG_19__SCAN_IN), .Z(n13587) );
  OAI21_X1 U15747 ( .B1(n13587), .B2(n15136), .A(n15204), .ZN(n13585) );
  AOI21_X1 U15748 ( .B1(n13586), .B2(n15198), .A(n13585), .ZN(n13590) );
  AOI22_X1 U15749 ( .A1(n13588), .A2(n15198), .B1(n15190), .B2(n13587), .ZN(
        n13589) );
  MUX2_X1 U15750 ( .A(n13590), .B(n13589), .S(n6555), .Z(n13592) );
  OAI211_X1 U15751 ( .C1(n7994), .C2(n15166), .A(n13592), .B(n13591), .ZN(
        P2_U3233) );
  XOR2_X1 U15752 ( .A(n13597), .B(n13600), .Z(n13594) );
  NAND2_X1 U15753 ( .A1(n13594), .A2(n13690), .ZN(n13837) );
  OR2_X1 U15754 ( .A1(n13596), .A2(n13595), .ZN(n13839) );
  NOR2_X1 U15755 ( .A1(n13812), .A2(n13839), .ZN(n13603) );
  INV_X1 U15756 ( .A(n13597), .ZN(n13838) );
  NOR2_X1 U15757 ( .A1(n13838), .A2(n13828), .ZN(n13598) );
  AOI211_X1 U15758 ( .C1(P2_REG2_REG_31__SCAN_IN), .C2(n13812), .A(n13603), 
        .B(n13598), .ZN(n13599) );
  OAI21_X1 U15759 ( .B1(n13837), .B2(n13724), .A(n13599), .ZN(P2_U3234) );
  OAI211_X1 U15760 ( .C1(n13601), .C2(n13841), .A(n13690), .B(n13600), .ZN(
        n13840) );
  NOR2_X1 U15761 ( .A1(n13841), .A2(n13828), .ZN(n13602) );
  AOI211_X1 U15762 ( .C1(n13812), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13603), 
        .B(n13602), .ZN(n13604) );
  OAI21_X1 U15763 ( .B1(n13840), .B2(n13724), .A(n13604), .ZN(P2_U3235) );
  INV_X1 U15764 ( .A(n13605), .ZN(n13606) );
  AOI21_X1 U15765 ( .B1(n13606), .B2(n13611), .A(n13799), .ZN(n13609) );
  AOI21_X1 U15766 ( .B1(n13609), .B2(n13608), .A(n13607), .ZN(n13845) );
  OAI21_X1 U15767 ( .B1(n13612), .B2(n13611), .A(n13610), .ZN(n13846) );
  OAI22_X1 U15768 ( .A1(n13770), .A2(n13614), .B1(n13613), .B2(n13784), .ZN(
        n13615) );
  AOI21_X1 U15769 ( .B1(n13843), .B2(n13734), .A(n13615), .ZN(n13619) );
  AOI21_X1 U15770 ( .B1(n13843), .B2(n13625), .A(n8285), .ZN(n13617) );
  NAND2_X1 U15771 ( .A1(n13842), .A2(n13835), .ZN(n13618) );
  OAI211_X1 U15772 ( .C1(n13846), .C2(n13832), .A(n13619), .B(n13618), .ZN(
        n13620) );
  INV_X1 U15773 ( .A(n13620), .ZN(n13621) );
  OAI21_X1 U15774 ( .B1(n13845), .B2(n13812), .A(n13621), .ZN(P2_U3237) );
  XNOR2_X1 U15775 ( .A(n13622), .B(n13628), .ZN(n13624) );
  AOI21_X1 U15776 ( .B1(n13624), .B2(n13819), .A(n13623), .ZN(n13853) );
  AOI21_X1 U15777 ( .B1(n13849), .B2(n13646), .A(n8285), .ZN(n13626) );
  NAND2_X1 U15778 ( .A1(n13626), .A2(n13625), .ZN(n13852) );
  NAND2_X1 U15779 ( .A1(n13628), .A2(n13627), .ZN(n13847) );
  NAND3_X1 U15780 ( .A1(n13848), .A2(n13847), .A3(n13728), .ZN(n13633) );
  OAI22_X1 U15781 ( .A1(n13770), .A2(n13630), .B1(n13629), .B2(n13784), .ZN(
        n13631) );
  AOI21_X1 U15782 ( .B1(n13849), .B2(n13734), .A(n13631), .ZN(n13632) );
  OAI211_X1 U15783 ( .C1(n13852), .C2(n13724), .A(n13633), .B(n13632), .ZN(
        n13634) );
  INV_X1 U15784 ( .A(n13634), .ZN(n13635) );
  OAI21_X1 U15785 ( .B1(n13853), .B2(n13812), .A(n13635), .ZN(P2_U3238) );
  XNOR2_X1 U15786 ( .A(n13636), .B(n13639), .ZN(n13638) );
  AOI222_X1 U15787 ( .A1(n13819), .A2(n13638), .B1(n13637), .B2(n13816), .C1(
        n13668), .C2(n13814), .ZN(n13857) );
  XNOR2_X1 U15788 ( .A(n13640), .B(n13639), .ZN(n13858) );
  OAI22_X1 U15789 ( .A1(n13770), .A2(n13642), .B1(n13641), .B2(n13784), .ZN(
        n13643) );
  AOI21_X1 U15790 ( .B1(n13855), .B2(n13734), .A(n13643), .ZN(n13648) );
  OR2_X1 U15791 ( .A1(n13644), .A2(n13662), .ZN(n13645) );
  AND3_X1 U15792 ( .A1(n13646), .A2(n13645), .A3(n13690), .ZN(n13854) );
  NAND2_X1 U15793 ( .A1(n13854), .A2(n13835), .ZN(n13647) );
  OAI211_X1 U15794 ( .C1(n13858), .C2(n13832), .A(n13648), .B(n13647), .ZN(
        n13649) );
  INV_X1 U15795 ( .A(n13649), .ZN(n13650) );
  OAI21_X1 U15796 ( .B1(n13857), .B2(n13812), .A(n13650), .ZN(P2_U3239) );
  XOR2_X1 U15797 ( .A(n13651), .B(n13653), .Z(n13863) );
  OAI21_X1 U15798 ( .B1(n13654), .B2(n13653), .A(n13652), .ZN(n13656) );
  AOI21_X1 U15799 ( .B1(n13656), .B2(n13819), .A(n13655), .ZN(n13862) );
  OAI22_X1 U15800 ( .A1(n13770), .A2(n13658), .B1(n13657), .B2(n13784), .ZN(
        n13659) );
  AOI21_X1 U15801 ( .B1(n13860), .B2(n13734), .A(n13659), .ZN(n13664) );
  NAND2_X1 U15802 ( .A1(n13860), .A2(n13671), .ZN(n13660) );
  NAND2_X1 U15803 ( .A1(n13660), .A2(n13690), .ZN(n13661) );
  NOR2_X1 U15804 ( .A1(n13662), .A2(n13661), .ZN(n13859) );
  NAND2_X1 U15805 ( .A1(n13859), .A2(n13835), .ZN(n13663) );
  OAI211_X1 U15806 ( .C1(n13862), .C2(n13812), .A(n13664), .B(n13663), .ZN(
        n13665) );
  INV_X1 U15807 ( .A(n13665), .ZN(n13666) );
  OAI21_X1 U15808 ( .B1(n13863), .B2(n13832), .A(n13666), .ZN(P2_U3240) );
  XNOR2_X1 U15809 ( .A(n13667), .B(n13679), .ZN(n13670) );
  AOI222_X1 U15810 ( .A1(n13819), .A2(n13670), .B1(n13669), .B2(n13814), .C1(
        n13668), .C2(n13816), .ZN(n13867) );
  INV_X1 U15811 ( .A(n13693), .ZN(n13673) );
  INV_X1 U15812 ( .A(n13671), .ZN(n13672) );
  AOI211_X1 U15813 ( .C1(n13865), .C2(n13673), .A(n8285), .B(n13672), .ZN(
        n13864) );
  INV_X1 U15814 ( .A(n13674), .ZN(n13675) );
  AOI22_X1 U15815 ( .A1(n13812), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n13675), 
        .B2(n13825), .ZN(n13676) );
  OAI21_X1 U15816 ( .B1(n13677), .B2(n13828), .A(n13676), .ZN(n13681) );
  OAI21_X1 U15817 ( .B1(n13679), .B2(n6652), .A(n13678), .ZN(n13868) );
  NOR2_X1 U15818 ( .A1(n13868), .A2(n13832), .ZN(n13680) );
  AOI211_X1 U15819 ( .C1(n13864), .C2(n13835), .A(n13681), .B(n13680), .ZN(
        n13682) );
  OAI21_X1 U15820 ( .B1(n13867), .B2(n13812), .A(n13682), .ZN(P2_U3241) );
  XNOR2_X1 U15821 ( .A(n13683), .B(n13689), .ZN(n13686) );
  AOI222_X1 U15822 ( .A1(n13819), .A2(n13686), .B1(n13685), .B2(n13816), .C1(
        n13684), .C2(n13814), .ZN(n13872) );
  OAI21_X1 U15823 ( .B1(n13689), .B2(n13688), .A(n13687), .ZN(n13873) );
  INV_X1 U15824 ( .A(n13873), .ZN(n13698) );
  NAND2_X1 U15825 ( .A1(n13870), .A2(n13710), .ZN(n13691) );
  NAND2_X1 U15826 ( .A1(n13691), .A2(n13690), .ZN(n13692) );
  NOR2_X1 U15827 ( .A1(n13693), .A2(n13692), .ZN(n13869) );
  NAND2_X1 U15828 ( .A1(n13869), .A2(n13835), .ZN(n13696) );
  AOI22_X1 U15829 ( .A1(n13812), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n13694), 
        .B2(n13825), .ZN(n13695) );
  OAI211_X1 U15830 ( .C1(n7784), .C2(n13828), .A(n13696), .B(n13695), .ZN(
        n13697) );
  AOI21_X1 U15831 ( .B1(n13728), .B2(n13698), .A(n13697), .ZN(n13699) );
  OAI21_X1 U15832 ( .B1(n13872), .B2(n13812), .A(n13699), .ZN(P2_U3242) );
  INV_X1 U15833 ( .A(n13700), .ZN(n13705) );
  AOI21_X1 U15834 ( .B1(n6643), .B2(n13705), .A(n13799), .ZN(n13703) );
  AOI21_X1 U15835 ( .B1(n13703), .B2(n13702), .A(n13701), .ZN(n13877) );
  OAI21_X1 U15836 ( .B1(n13705), .B2(n6657), .A(n13704), .ZN(n13878) );
  OAI22_X1 U15837 ( .A1(n13770), .A2(n13707), .B1(n13706), .B2(n13784), .ZN(
        n13708) );
  AOI21_X1 U15838 ( .B1(n13875), .B2(n13734), .A(n13708), .ZN(n13712) );
  AOI21_X1 U15839 ( .B1(n13875), .B2(n13718), .A(n8285), .ZN(n13709) );
  AND2_X1 U15840 ( .A1(n13710), .A2(n13709), .ZN(n13874) );
  NAND2_X1 U15841 ( .A1(n13874), .A2(n13835), .ZN(n13711) );
  OAI211_X1 U15842 ( .C1(n13878), .C2(n13832), .A(n13712), .B(n13711), .ZN(
        n13713) );
  INV_X1 U15843 ( .A(n13713), .ZN(n13714) );
  OAI21_X1 U15844 ( .B1(n13877), .B2(n13812), .A(n13714), .ZN(P2_U3243) );
  XNOR2_X1 U15845 ( .A(n13715), .B(n13726), .ZN(n13717) );
  AOI21_X1 U15846 ( .B1(n13717), .B2(n13819), .A(n13716), .ZN(n13885) );
  AOI21_X1 U15847 ( .B1(n13879), .B2(n13732), .A(n8285), .ZN(n13719) );
  NAND2_X1 U15848 ( .A1(n13719), .A2(n13718), .ZN(n13882) );
  OAI22_X1 U15849 ( .A1(n13770), .A2(n13721), .B1(n13720), .B2(n13784), .ZN(
        n13722) );
  AOI21_X1 U15850 ( .B1(n13879), .B2(n13734), .A(n13722), .ZN(n13723) );
  OAI21_X1 U15851 ( .B1(n13882), .B2(n13724), .A(n13723), .ZN(n13725) );
  INV_X1 U15852 ( .A(n13725), .ZN(n13730) );
  NAND2_X1 U15853 ( .A1(n13727), .A2(n13726), .ZN(n13880) );
  NAND3_X1 U15854 ( .A1(n13881), .A2(n13728), .A3(n13880), .ZN(n13729) );
  OAI211_X1 U15855 ( .C1(n13885), .C2(n13812), .A(n13730), .B(n13729), .ZN(
        P2_U3244) );
  XNOR2_X1 U15856 ( .A(n13731), .B(n13740), .ZN(n13890) );
  AOI21_X1 U15857 ( .B1(n13887), .B2(n13748), .A(n8285), .ZN(n13733) );
  AND2_X1 U15858 ( .A1(n13733), .A2(n13732), .ZN(n13886) );
  NAND2_X1 U15859 ( .A1(n13887), .A2(n13734), .ZN(n13736) );
  NAND2_X1 U15860 ( .A1(n13812), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n13735) );
  OAI211_X1 U15861 ( .C1(n13784), .C2(n13737), .A(n13736), .B(n13735), .ZN(
        n13745) );
  OAI21_X1 U15862 ( .B1(n13740), .B2(n13739), .A(n13738), .ZN(n13743) );
  AOI222_X1 U15863 ( .A1(n13819), .A2(n13743), .B1(n13742), .B2(n13816), .C1(
        n13741), .C2(n13814), .ZN(n13889) );
  NOR2_X1 U15864 ( .A1(n13889), .A2(n13812), .ZN(n13744) );
  AOI211_X1 U15865 ( .C1(n13886), .C2(n13835), .A(n13745), .B(n13744), .ZN(
        n13746) );
  OAI21_X1 U15866 ( .B1(n13890), .B2(n13832), .A(n13746), .ZN(P2_U3245) );
  XNOR2_X1 U15867 ( .A(n13747), .B(n13752), .ZN(n13895) );
  AOI211_X1 U15868 ( .C1(n13893), .C2(n13765), .A(n8285), .B(n7500), .ZN(
        n13892) );
  INV_X1 U15869 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13749) );
  OAI22_X1 U15870 ( .A1(n13750), .A2(n13828), .B1(n13770), .B2(n13749), .ZN(
        n13758) );
  XOR2_X1 U15871 ( .A(n13752), .B(n13751), .Z(n13754) );
  OAI21_X1 U15872 ( .B1(n13754), .B2(n13799), .A(n13753), .ZN(n13891) );
  AOI21_X1 U15873 ( .B1(n13755), .B2(n13825), .A(n13891), .ZN(n13756) );
  NOR2_X1 U15874 ( .A1(n13756), .A2(n13812), .ZN(n13757) );
  AOI211_X1 U15875 ( .C1(n13892), .C2(n13835), .A(n13758), .B(n13757), .ZN(
        n13759) );
  OAI21_X1 U15876 ( .B1(n13832), .B2(n13895), .A(n13759), .ZN(P2_U3246) );
  XNOR2_X1 U15877 ( .A(n13761), .B(n13760), .ZN(n13900) );
  XNOR2_X1 U15878 ( .A(n6714), .B(n13762), .ZN(n13764) );
  OAI21_X1 U15879 ( .B1(n13764), .B2(n13799), .A(n13763), .ZN(n13896) );
  NAND2_X1 U15880 ( .A1(n13896), .A2(n13770), .ZN(n13774) );
  INV_X1 U15881 ( .A(n13765), .ZN(n13766) );
  AOI211_X1 U15882 ( .C1(n13898), .C2(n13780), .A(n8285), .B(n13766), .ZN(
        n13897) );
  NOR2_X1 U15883 ( .A1(n13767), .A2(n13828), .ZN(n13772) );
  INV_X1 U15884 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13769) );
  OAI22_X1 U15885 ( .A1(n13770), .A2(n13769), .B1(n13768), .B2(n13784), .ZN(
        n13771) );
  AOI211_X1 U15886 ( .C1(n13897), .C2(n13835), .A(n13772), .B(n13771), .ZN(
        n13773) );
  OAI211_X1 U15887 ( .C1(n13900), .C2(n13832), .A(n13774), .B(n13773), .ZN(
        P2_U3247) );
  XOR2_X1 U15888 ( .A(n13775), .B(n13777), .Z(n13905) );
  XOR2_X1 U15889 ( .A(n13776), .B(n13777), .Z(n13779) );
  OAI21_X1 U15890 ( .B1(n13779), .B2(n13799), .A(n13778), .ZN(n13901) );
  NAND2_X1 U15891 ( .A1(n13901), .A2(n13770), .ZN(n13790) );
  INV_X1 U15892 ( .A(n13803), .ZN(n13782) );
  INV_X1 U15893 ( .A(n13780), .ZN(n13781) );
  AOI211_X1 U15894 ( .C1(n13903), .C2(n13782), .A(n8285), .B(n13781), .ZN(
        n13902) );
  NOR2_X1 U15895 ( .A1(n13783), .A2(n13828), .ZN(n13788) );
  OAI22_X1 U15896 ( .A1(n13770), .A2(n13786), .B1(n13785), .B2(n13784), .ZN(
        n13787) );
  AOI211_X1 U15897 ( .C1(n13902), .C2(n13835), .A(n13788), .B(n13787), .ZN(
        n13789) );
  OAI211_X1 U15898 ( .C1(n13905), .C2(n13832), .A(n13790), .B(n13789), .ZN(
        P2_U3248) );
  NAND2_X1 U15899 ( .A1(n13791), .A2(n13795), .ZN(n13792) );
  XOR2_X1 U15900 ( .A(n13795), .B(n13794), .Z(n13800) );
  AOI22_X1 U15901 ( .A1(n13797), .A2(n13816), .B1(n13796), .B2(n13814), .ZN(
        n13798) );
  OAI21_X1 U15902 ( .B1(n13800), .B2(n13799), .A(n13798), .ZN(n13801) );
  AOI21_X1 U15903 ( .B1(n13802), .B2(n13807), .A(n13801), .ZN(n13909) );
  AOI211_X1 U15904 ( .C1(n13907), .C2(n13820), .A(n8285), .B(n13803), .ZN(
        n13906) );
  AOI22_X1 U15905 ( .A1(n13812), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n13804), 
        .B2(n13825), .ZN(n13805) );
  OAI21_X1 U15906 ( .B1(n13806), .B2(n13828), .A(n13805), .ZN(n13810) );
  NOR2_X1 U15907 ( .A1(n13910), .A2(n13808), .ZN(n13809) );
  AOI211_X1 U15908 ( .C1(n13906), .C2(n13835), .A(n13810), .B(n13809), .ZN(
        n13811) );
  OAI21_X1 U15909 ( .B1(n13909), .B2(n13812), .A(n13811), .ZN(P2_U3249) );
  XNOR2_X1 U15910 ( .A(n13813), .B(n13830), .ZN(n13818) );
  AOI222_X1 U15911 ( .A1(n13819), .A2(n13818), .B1(n13817), .B2(n13816), .C1(
        n13815), .C2(n13814), .ZN(n13914) );
  INV_X1 U15912 ( .A(n13820), .ZN(n13821) );
  AOI211_X1 U15913 ( .C1(n13912), .C2(n13823), .A(n8285), .B(n13821), .ZN(
        n13911) );
  INV_X1 U15914 ( .A(n13824), .ZN(n13826) );
  AOI22_X1 U15915 ( .A1(n13812), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n13826), 
        .B2(n13825), .ZN(n13827) );
  OAI21_X1 U15916 ( .B1(n13829), .B2(n13828), .A(n13827), .ZN(n13834) );
  XOR2_X1 U15917 ( .A(n13831), .B(n13830), .Z(n13915) );
  NOR2_X1 U15918 ( .A1(n13915), .A2(n13832), .ZN(n13833) );
  AOI211_X1 U15919 ( .C1(n13911), .C2(n13835), .A(n13834), .B(n13833), .ZN(
        n13836) );
  OAI21_X1 U15920 ( .B1(n13914), .B2(n13812), .A(n13836), .ZN(P2_U3250) );
  OAI211_X1 U15921 ( .C1(n13838), .C2(n15263), .A(n13837), .B(n13839), .ZN(
        n13925) );
  MUX2_X1 U15922 ( .A(n13925), .B(P2_REG1_REG_31__SCAN_IN), .S(n15277), .Z(
        P2_U3530) );
  OAI211_X1 U15923 ( .C1(n13841), .C2(n15263), .A(n13840), .B(n13839), .ZN(
        n13926) );
  MUX2_X1 U15924 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13926), .S(n15279), .Z(
        P2_U3529) );
  OAI211_X1 U15925 ( .C1(n15249), .C2(n13846), .A(n13845), .B(n13844), .ZN(
        n13927) );
  MUX2_X1 U15926 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13927), .S(n15279), .Z(
        P2_U3527) );
  NAND3_X1 U15927 ( .A1(n13848), .A2(n13847), .A3(n9794), .ZN(n13851) );
  NAND2_X1 U15928 ( .A1(n13849), .A2(n15251), .ZN(n13850) );
  NAND4_X1 U15929 ( .A1(n13853), .A2(n13852), .A3(n13851), .A4(n13850), .ZN(
        n13928) );
  MUX2_X1 U15930 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13928), .S(n15279), .Z(
        P2_U3526) );
  AOI21_X1 U15931 ( .B1(n15251), .B2(n13855), .A(n13854), .ZN(n13856) );
  OAI211_X1 U15932 ( .C1(n15249), .C2(n13858), .A(n13857), .B(n13856), .ZN(
        n13929) );
  MUX2_X1 U15933 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13929), .S(n15279), .Z(
        P2_U3525) );
  AOI21_X1 U15934 ( .B1(n15251), .B2(n13860), .A(n13859), .ZN(n13861) );
  OAI211_X1 U15935 ( .C1(n15249), .C2(n13863), .A(n13862), .B(n13861), .ZN(
        n13930) );
  MUX2_X1 U15936 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13930), .S(n15279), .Z(
        P2_U3524) );
  AOI21_X1 U15937 ( .B1(n15251), .B2(n13865), .A(n13864), .ZN(n13866) );
  OAI211_X1 U15938 ( .C1(n15249), .C2(n13868), .A(n13867), .B(n13866), .ZN(
        n13931) );
  MUX2_X1 U15939 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13931), .S(n15279), .Z(
        P2_U3523) );
  AOI21_X1 U15940 ( .B1(n15251), .B2(n13870), .A(n13869), .ZN(n13871) );
  OAI211_X1 U15941 ( .C1(n15249), .C2(n13873), .A(n13872), .B(n13871), .ZN(
        n13932) );
  MUX2_X1 U15942 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13932), .S(n15279), .Z(
        P2_U3522) );
  AOI21_X1 U15943 ( .B1(n15251), .B2(n13875), .A(n13874), .ZN(n13876) );
  OAI211_X1 U15944 ( .C1(n15249), .C2(n13878), .A(n13877), .B(n13876), .ZN(
        n13933) );
  MUX2_X1 U15945 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13933), .S(n15279), .Z(
        P2_U3521) );
  NAND2_X1 U15946 ( .A1(n13879), .A2(n15251), .ZN(n13884) );
  NAND3_X1 U15947 ( .A1(n13881), .A2(n9794), .A3(n13880), .ZN(n13883) );
  NAND4_X1 U15948 ( .A1(n13885), .A2(n13884), .A3(n13883), .A4(n13882), .ZN(
        n13934) );
  MUX2_X1 U15949 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13934), .S(n15279), .Z(
        P2_U3520) );
  AOI21_X1 U15950 ( .B1(n15251), .B2(n13887), .A(n13886), .ZN(n13888) );
  OAI211_X1 U15951 ( .C1(n15249), .C2(n13890), .A(n13889), .B(n13888), .ZN(
        n13935) );
  MUX2_X1 U15952 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13935), .S(n15279), .Z(
        P2_U3519) );
  AOI211_X1 U15953 ( .C1(n15251), .C2(n13893), .A(n13892), .B(n13891), .ZN(
        n13894) );
  OAI21_X1 U15954 ( .B1(n15249), .B2(n13895), .A(n13894), .ZN(n13936) );
  MUX2_X1 U15955 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13936), .S(n15279), .Z(
        P2_U3518) );
  AOI211_X1 U15956 ( .C1(n15251), .C2(n13898), .A(n13897), .B(n13896), .ZN(
        n13899) );
  OAI21_X1 U15957 ( .B1(n15249), .B2(n13900), .A(n13899), .ZN(n13937) );
  MUX2_X1 U15958 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13937), .S(n15279), .Z(
        P2_U3517) );
  AOI211_X1 U15959 ( .C1(n15251), .C2(n13903), .A(n13902), .B(n13901), .ZN(
        n13904) );
  OAI21_X1 U15960 ( .B1(n15249), .B2(n13905), .A(n13904), .ZN(n13938) );
  MUX2_X1 U15961 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13938), .S(n15279), .Z(
        P2_U3516) );
  AOI21_X1 U15962 ( .B1(n15251), .B2(n13907), .A(n13906), .ZN(n13908) );
  OAI211_X1 U15963 ( .C1(n15255), .C2(n13910), .A(n13909), .B(n13908), .ZN(
        n13939) );
  MUX2_X1 U15964 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13939), .S(n15279), .Z(
        P2_U3515) );
  AOI21_X1 U15965 ( .B1(n15251), .B2(n13912), .A(n13911), .ZN(n13913) );
  OAI211_X1 U15966 ( .C1(n15249), .C2(n13915), .A(n13914), .B(n13913), .ZN(
        n13940) );
  MUX2_X1 U15967 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13940), .S(n15279), .Z(
        P2_U3514) );
  AOI21_X1 U15968 ( .B1(n15251), .B2(n14847), .A(n13916), .ZN(n13917) );
  OAI211_X1 U15969 ( .C1(n15249), .C2(n13919), .A(n13918), .B(n13917), .ZN(
        n13941) );
  MUX2_X1 U15970 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13941), .S(n15279), .Z(
        P2_U3513) );
  AOI211_X1 U15971 ( .C1(n15251), .C2(n13922), .A(n13921), .B(n13920), .ZN(
        n13923) );
  OAI21_X1 U15972 ( .B1(n15249), .B2(n13924), .A(n13923), .ZN(n15225) );
  MUX2_X1 U15973 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n15225), .S(n15279), .Z(
        P2_U3501) );
  MUX2_X1 U15974 ( .A(n13925), .B(P2_REG0_REG_31__SCAN_IN), .S(n9800), .Z(
        P2_U3498) );
  MUX2_X1 U15975 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13926), .S(n15270), .Z(
        P2_U3497) );
  MUX2_X1 U15976 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13927), .S(n15270), .Z(
        P2_U3495) );
  MUX2_X1 U15977 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13928), .S(n15270), .Z(
        P2_U3494) );
  MUX2_X1 U15978 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13929), .S(n15270), .Z(
        P2_U3493) );
  MUX2_X1 U15979 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13930), .S(n15270), .Z(
        P2_U3492) );
  MUX2_X1 U15980 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13931), .S(n15270), .Z(
        P2_U3491) );
  MUX2_X1 U15981 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13932), .S(n15270), .Z(
        P2_U3490) );
  MUX2_X1 U15982 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13933), .S(n15270), .Z(
        P2_U3489) );
  MUX2_X1 U15983 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13934), .S(n15270), .Z(
        P2_U3488) );
  MUX2_X1 U15984 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13935), .S(n15270), .Z(
        P2_U3487) );
  MUX2_X1 U15985 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13936), .S(n15270), .Z(
        P2_U3486) );
  MUX2_X1 U15986 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13937), .S(n15270), .Z(
        P2_U3484) );
  MUX2_X1 U15987 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13938), .S(n15270), .Z(
        P2_U3481) );
  MUX2_X1 U15988 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13939), .S(n15270), .Z(
        P2_U3478) );
  MUX2_X1 U15989 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13940), .S(n15270), .Z(
        P2_U3475) );
  MUX2_X1 U15990 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13941), .S(n15270), .Z(
        P2_U3472) );
  INV_X1 U15991 ( .A(n13942), .ZN(n14622) );
  NOR4_X1 U15992 ( .A1(n7972), .A2(P2_IR_REG_30__SCAN_IN), .A3(n13943), .A4(
        P2_U3088), .ZN(n13944) );
  AOI21_X1 U15993 ( .B1(n13945), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13944), 
        .ZN(n13946) );
  OAI21_X1 U15994 ( .B1(n14622), .B2(n13967), .A(n13946), .ZN(P2_U3296) );
  INV_X1 U15995 ( .A(n13948), .ZN(n14627) );
  OAI222_X1 U15996 ( .A1(n13964), .A2(n13950), .B1(P2_U3088), .B2(n13949), 
        .C1(n13967), .C2(n14627), .ZN(P2_U3298) );
  NAND2_X1 U15997 ( .A1(n12536), .A2(n13951), .ZN(n13953) );
  OAI211_X1 U15998 ( .C1(n15457), .C2(n13964), .A(n13953), .B(n13952), .ZN(
        P2_U3299) );
  INV_X1 U15999 ( .A(n13954), .ZN(n14630) );
  OAI222_X1 U16000 ( .A1(n13964), .A2(n13956), .B1(n13967), .B2(n14630), .C1(
        n13955), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U16001 ( .A(n13957), .ZN(n13960) );
  INV_X1 U16002 ( .A(n13958), .ZN(n14633) );
  OAI222_X1 U16003 ( .A1(P2_U3088), .A2(n13960), .B1(n13967), .B2(n14633), 
        .C1(n13959), .C2(n13964), .ZN(P2_U3301) );
  OAI222_X1 U16004 ( .A1(n13964), .A2(n13963), .B1(n13967), .B2(n13962), .C1(
        P2_U3088), .C2(n13961), .ZN(P2_U3302) );
  INV_X1 U16005 ( .A(n13965), .ZN(n14637) );
  OAI222_X1 U16006 ( .A1(P2_U3088), .A2(n13968), .B1(n13967), .B2(n14637), 
        .C1(n13966), .C2(n13964), .ZN(P2_U3303) );
  MUX2_X1 U16007 ( .A(n6742), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OAI21_X1 U16008 ( .B1(n13972), .B2(n13971), .A(n13970), .ZN(n13973) );
  OAI22_X1 U16009 ( .A1(n14085), .A2(n14274), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13974), .ZN(n13976) );
  NOR2_X1 U16010 ( .A1(n14965), .A2(n14283), .ZN(n13975) );
  AOI211_X1 U16011 ( .C1(n14087), .C2(n7446), .A(n13976), .B(n13975), .ZN(
        n13977) );
  AND3_X1 U16012 ( .A1(n14050), .A2(n13979), .A3(n13978), .ZN(n13980) );
  OAI21_X1 U16013 ( .B1(n13981), .B2(n13980), .A(n14961), .ZN(n13987) );
  INV_X1 U16014 ( .A(n14348), .ZN(n13985) );
  AND2_X1 U16015 ( .A1(n14094), .A2(n14477), .ZN(n13982) );
  AOI21_X1 U16016 ( .B1(n14095), .B2(n14479), .A(n13982), .ZN(n14544) );
  INV_X1 U16017 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13983) );
  OAI22_X1 U16018 ( .A1(n14544), .A2(n14862), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13983), .ZN(n13984) );
  AOI21_X1 U16019 ( .B1(n13985), .B2(n14068), .A(n13984), .ZN(n13986) );
  OAI211_X1 U16020 ( .C1(n14546), .C2(n14864), .A(n13987), .B(n13986), .ZN(
        P1_U3216) );
  INV_X1 U16021 ( .A(n14574), .ZN(n14414) );
  AND2_X1 U16022 ( .A1(n14061), .A2(n13988), .ZN(n13991) );
  OAI211_X1 U16023 ( .C1(n13991), .C2(n13990), .A(n14961), .B(n13989), .ZN(
        n13996) );
  NAND2_X1 U16024 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14238)
         );
  OAI21_X1 U16025 ( .B1(n13992), .B2(n14085), .A(n14238), .ZN(n13994) );
  NOR2_X1 U16026 ( .A1(n14965), .A2(n14411), .ZN(n13993) );
  AOI211_X1 U16027 ( .C1(n14087), .C2(n14408), .A(n13994), .B(n13993), .ZN(
        n13995) );
  OAI211_X1 U16028 ( .C1(n14414), .C2(n14864), .A(n13996), .B(n13995), .ZN(
        P1_U3219) );
  INV_X1 U16029 ( .A(n14381), .ZN(n14560) );
  OAI21_X1 U16030 ( .B1(n13999), .B2(n13998), .A(n13997), .ZN(n14000) );
  NAND2_X1 U16031 ( .A1(n14000), .A2(n14961), .ZN(n14005) );
  INV_X1 U16032 ( .A(n14378), .ZN(n14003) );
  AOI22_X1 U16033 ( .A1(n14095), .A2(n14477), .B1(n14479), .B2(n14409), .ZN(
        n14558) );
  OAI22_X1 U16034 ( .A1(n14558), .A2(n14862), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14001), .ZN(n14002) );
  AOI21_X1 U16035 ( .B1(n14003), .B2(n14068), .A(n14002), .ZN(n14004) );
  OAI211_X1 U16036 ( .C1(n14560), .C2(n14864), .A(n14005), .B(n14004), .ZN(
        P1_U3223) );
  OAI21_X1 U16037 ( .B1(n14008), .B2(n14007), .A(n14006), .ZN(n14009) );
  NAND2_X1 U16038 ( .A1(n14009), .A2(n14961), .ZN(n14015) );
  INV_X1 U16039 ( .A(n14315), .ZN(n14013) );
  NAND2_X1 U16040 ( .A1(n7446), .A2(n14477), .ZN(n14011) );
  NAND2_X1 U16041 ( .A1(n14094), .A2(n14479), .ZN(n14010) );
  AND2_X1 U16042 ( .A1(n14011), .A2(n14010), .ZN(n14532) );
  INV_X1 U16043 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n15697) );
  OAI22_X1 U16044 ( .A1(n14862), .A2(n14532), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15697), .ZN(n14012) );
  AOI21_X1 U16045 ( .B1(n14068), .B2(n14013), .A(n14012), .ZN(n14014) );
  OAI211_X1 U16046 ( .C1(n7335), .C2(n14864), .A(n14015), .B(n14014), .ZN(
        P1_U3225) );
  AOI21_X1 U16047 ( .B1(n14017), .B2(n14016), .A(n6695), .ZN(n14023) );
  OAI21_X1 U16048 ( .B1(n14085), .B2(n14463), .A(n14018), .ZN(n14019) );
  AOI21_X1 U16049 ( .B1(n14087), .B2(n14097), .A(n14019), .ZN(n14020) );
  OAI21_X1 U16050 ( .B1(n14965), .B2(n14469), .A(n14020), .ZN(n14021) );
  AOI21_X1 U16051 ( .B1(n14591), .B2(n14090), .A(n14021), .ZN(n14022) );
  OAI21_X1 U16052 ( .B1(n14023), .B2(n14935), .A(n14022), .ZN(P1_U3226) );
  INV_X1 U16053 ( .A(n14024), .ZN(n14028) );
  NOR3_X1 U16054 ( .A1(n6695), .A2(n14026), .A3(n14025), .ZN(n14027) );
  OAI21_X1 U16055 ( .B1(n14028), .B2(n14027), .A(n14961), .ZN(n14033) );
  NAND2_X1 U16056 ( .A1(n14087), .A2(n14478), .ZN(n14030) );
  OAI211_X1 U16057 ( .C1(n14448), .C2(n14085), .A(n14030), .B(n14029), .ZN(
        n14031) );
  AOI21_X1 U16058 ( .B1(n14068), .B2(n14442), .A(n14031), .ZN(n14032) );
  OAI211_X1 U16059 ( .C1(n14444), .C2(n14864), .A(n14033), .B(n14032), .ZN(
        P1_U3228) );
  AOI21_X1 U16060 ( .B1(n14035), .B2(n14034), .A(n6632), .ZN(n14040) );
  AND2_X1 U16061 ( .A1(n14334), .A2(n14951), .ZN(n14540) );
  AOI22_X1 U16062 ( .A1(n14054), .A2(n14325), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14037) );
  NAND2_X1 U16063 ( .A1(n14087), .A2(n14358), .ZN(n14036) );
  OAI211_X1 U16064 ( .C1(n14965), .C2(n14335), .A(n14037), .B(n14036), .ZN(
        n14038) );
  AOI21_X1 U16065 ( .B1(n14540), .B2(n14953), .A(n14038), .ZN(n14039) );
  OAI21_X1 U16066 ( .B1(n14040), .B2(n14935), .A(n14039), .ZN(P1_U3229) );
  XNOR2_X1 U16067 ( .A(n14042), .B(n14041), .ZN(n14049) );
  OAI22_X1 U16068 ( .A1(n14396), .A2(n14085), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14043), .ZN(n14044) );
  AOI21_X1 U16069 ( .B1(n14087), .B2(n14096), .A(n14044), .ZN(n14045) );
  OAI21_X1 U16070 ( .B1(n14965), .B2(n14046), .A(n14045), .ZN(n14047) );
  AOI21_X1 U16071 ( .B1(n14566), .B2(n14090), .A(n14047), .ZN(n14048) );
  OAI21_X1 U16072 ( .B1(n14049), .B2(n14935), .A(n14048), .ZN(P1_U3233) );
  OAI21_X1 U16073 ( .B1(n14052), .B2(n14051), .A(n14050), .ZN(n14053) );
  NAND2_X1 U16074 ( .A1(n14053), .A2(n14961), .ZN(n14059) );
  INV_X1 U16075 ( .A(n14087), .ZN(n14056) );
  AOI22_X1 U16076 ( .A1(n14054), .A2(n14358), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14055) );
  OAI21_X1 U16077 ( .B1(n14396), .B2(n14056), .A(n14055), .ZN(n14057) );
  AOI21_X1 U16078 ( .B1(n14366), .B2(n14068), .A(n14057), .ZN(n14058) );
  OAI211_X1 U16079 ( .C1(n14864), .C2(n14060), .A(n14059), .B(n14058), .ZN(
        P1_U3235) );
  INV_X1 U16080 ( .A(n14580), .ZN(n14433) );
  OAI21_X1 U16081 ( .B1(n14063), .B2(n14062), .A(n14061), .ZN(n14064) );
  NAND2_X1 U16082 ( .A1(n14064), .A2(n14961), .ZN(n14070) );
  NAND2_X1 U16083 ( .A1(n14087), .A2(n14425), .ZN(n14066) );
  OAI211_X1 U16084 ( .C1(n14427), .C2(n14085), .A(n14066), .B(n14065), .ZN(
        n14067) );
  AOI21_X1 U16085 ( .B1(n14068), .B2(n14431), .A(n14067), .ZN(n14069) );
  OAI211_X1 U16086 ( .C1(n14433), .C2(n14864), .A(n14070), .B(n14069), .ZN(
        P1_U3238) );
  OAI21_X1 U16087 ( .B1(n14073), .B2(n14072), .A(n14071), .ZN(n14074) );
  NAND2_X1 U16088 ( .A1(n14074), .A2(n14961), .ZN(n14080) );
  OAI22_X1 U16089 ( .A1(n14085), .A2(n14076), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14075), .ZN(n14078) );
  NOR2_X1 U16090 ( .A1(n14965), .A2(n14294), .ZN(n14077) );
  AOI211_X1 U16091 ( .C1(n14087), .C2(n14325), .A(n14078), .B(n14077), .ZN(
        n14079) );
  OAI211_X1 U16092 ( .C1(n14528), .C2(n14081), .A(n14080), .B(n14079), .ZN(
        P1_U3240) );
  AOI21_X1 U16093 ( .B1(n14084), .B2(n14083), .A(n14082), .ZN(n14092) );
  NAND2_X1 U16094 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14978)
         );
  OAI21_X1 U16095 ( .B1(n14085), .B2(n14447), .A(n14978), .ZN(n14086) );
  AOI21_X1 U16096 ( .B1(n14087), .B2(n14480), .A(n14086), .ZN(n14088) );
  OAI21_X1 U16097 ( .B1(n14965), .B2(n14485), .A(n14088), .ZN(n14089) );
  AOI21_X1 U16098 ( .B1(n14595), .B2(n14090), .A(n14089), .ZN(n14091) );
  OAI21_X1 U16099 ( .B1(n14092), .B2(n14935), .A(n14091), .ZN(P1_U3241) );
  MUX2_X1 U16100 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14246), .S(n6551), .Z(
        P1_U3591) );
  MUX2_X1 U16101 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14262), .S(n6551), .Z(
        P1_U3590) );
  MUX2_X1 U16102 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14093), .S(n6551), .Z(
        P1_U3589) );
  MUX2_X1 U16103 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14266), .S(n6551), .Z(
        P1_U3588) );
  MUX2_X1 U16104 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14301), .S(n6551), .Z(
        P1_U3587) );
  MUX2_X1 U16105 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n7446), .S(n6551), .Z(
        P1_U3586) );
  MUX2_X1 U16106 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14325), .S(n6551), .Z(
        P1_U3585) );
  MUX2_X1 U16107 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14094), .S(n6551), .Z(
        P1_U3584) );
  MUX2_X1 U16108 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14358), .S(n6551), .Z(
        P1_U3583) );
  MUX2_X1 U16109 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14095), .S(n6551), .Z(
        P1_U3582) );
  MUX2_X1 U16110 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14359), .S(n6551), .Z(
        P1_U3581) );
  MUX2_X1 U16111 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14409), .S(n6551), .Z(
        P1_U3580) );
  MUX2_X1 U16112 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14096), .S(n6551), .Z(
        P1_U3579) );
  MUX2_X1 U16113 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14408), .S(n6551), .Z(
        P1_U3578) );
  MUX2_X1 U16114 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14425), .S(n6551), .Z(
        P1_U3577) );
  MUX2_X1 U16115 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14478), .S(n6551), .Z(
        P1_U3576) );
  MUX2_X1 U16116 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14097), .S(n6551), .Z(
        P1_U3575) );
  MUX2_X1 U16117 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14480), .S(n6551), .Z(
        P1_U3574) );
  MUX2_X1 U16118 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14098), .S(n6551), .Z(
        P1_U3573) );
  MUX2_X1 U16119 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14099), .S(n6551), .Z(
        P1_U3572) );
  MUX2_X1 U16120 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14100), .S(n6551), .Z(
        P1_U3571) );
  MUX2_X1 U16121 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14101), .S(n6551), .Z(
        P1_U3570) );
  MUX2_X1 U16122 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14102), .S(n6551), .Z(
        P1_U3569) );
  MUX2_X1 U16123 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14103), .S(n6551), .Z(
        P1_U3568) );
  MUX2_X1 U16124 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14104), .S(n6551), .Z(
        P1_U3567) );
  MUX2_X1 U16125 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14105), .S(n6551), .Z(
        P1_U3566) );
  MUX2_X1 U16126 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14106), .S(n6551), .Z(
        P1_U3565) );
  MUX2_X1 U16127 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14107), .S(n6551), .Z(
        P1_U3564) );
  MUX2_X1 U16128 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14108), .S(n6551), .Z(
        P1_U3563) );
  MUX2_X1 U16129 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14109), .S(n6551), .Z(
        P1_U3562) );
  MUX2_X1 U16130 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14110), .S(n6551), .Z(
        P1_U3561) );
  OAI22_X1 U16131 ( .A1(n14980), .A2(n15651), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14111), .ZN(n14112) );
  AOI21_X1 U16132 ( .B1(n14113), .B2(n14206), .A(n14112), .ZN(n14120) );
  OAI211_X1 U16133 ( .C1(n14115), .C2(n14114), .A(n14233), .B(n14132), .ZN(
        n14119) );
  NAND2_X1 U16134 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14122) );
  OAI211_X1 U16135 ( .C1(n14117), .C2(n10651), .A(n14232), .B(n14116), .ZN(
        n14118) );
  NAND3_X1 U16136 ( .A1(n14120), .A2(n14119), .A3(n14118), .ZN(P1_U3244) );
  MUX2_X1 U16137 ( .A(n14122), .B(n14121), .S(n14629), .Z(n14126) );
  NAND2_X1 U16138 ( .A1(n14124), .A2(n14123), .ZN(n14125) );
  OAI211_X1 U16139 ( .C1(n14126), .C2(n10373), .A(n6551), .B(n14125), .ZN(
        n14171) );
  OAI22_X1 U16140 ( .A1(n14980), .A2(n14646), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14127), .ZN(n14128) );
  AOI21_X1 U16141 ( .B1(n14129), .B2(n14206), .A(n14128), .ZN(n14138) );
  MUX2_X1 U16142 ( .A(n10631), .B(P1_REG1_REG_2__SCAN_IN), .S(n14129), .Z(
        n14130) );
  NAND3_X1 U16143 ( .A1(n14132), .A2(n14131), .A3(n14130), .ZN(n14133) );
  NAND3_X1 U16144 ( .A1(n14233), .A2(n14140), .A3(n14133), .ZN(n14137) );
  OAI211_X1 U16145 ( .C1(n14135), .C2(n14134), .A(n14232), .B(n14145), .ZN(
        n14136) );
  NAND4_X1 U16146 ( .A1(n14171), .A2(n14138), .A3(n14137), .A4(n14136), .ZN(
        P1_U3245) );
  MUX2_X1 U16147 ( .A(n10634), .B(P1_REG1_REG_3__SCAN_IN), .S(n14148), .Z(
        n14141) );
  NAND3_X1 U16148 ( .A1(n14141), .A2(n14140), .A3(n14139), .ZN(n14142) );
  NAND3_X1 U16149 ( .A1(n14233), .A2(n14158), .A3(n14142), .ZN(n14152) );
  MUX2_X1 U16150 ( .A(n14143), .B(P1_REG2_REG_3__SCAN_IN), .S(n14148), .Z(
        n14146) );
  NAND3_X1 U16151 ( .A1(n14146), .A2(n14145), .A3(n14144), .ZN(n14147) );
  NAND3_X1 U16152 ( .A1(n14232), .A2(n14165), .A3(n14147), .ZN(n14151) );
  NAND2_X1 U16153 ( .A1(n14206), .A2(n14148), .ZN(n14150) );
  AND2_X1 U16154 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n14934) );
  AOI21_X1 U16155 ( .B1(n14212), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n14934), .ZN(
        n14149) );
  NAND4_X1 U16156 ( .A1(n14152), .A2(n14151), .A3(n14150), .A4(n14149), .ZN(
        P1_U3246) );
  NOR2_X1 U16157 ( .A1(n14976), .A2(n14153), .ZN(n14154) );
  AOI211_X1 U16158 ( .C1(n14212), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n14155), .B(
        n14154), .ZN(n14170) );
  MUX2_X1 U16159 ( .A(n10637), .B(P1_REG1_REG_4__SCAN_IN), .S(n14161), .Z(
        n14156) );
  NAND3_X1 U16160 ( .A1(n14158), .A2(n14157), .A3(n14156), .ZN(n14159) );
  NAND3_X1 U16161 ( .A1(n14233), .A2(n14160), .A3(n14159), .ZN(n14169) );
  MUX2_X1 U16162 ( .A(n14162), .B(P1_REG2_REG_4__SCAN_IN), .S(n14161), .Z(
        n14163) );
  NAND3_X1 U16163 ( .A1(n14165), .A2(n14164), .A3(n14163), .ZN(n14166) );
  NAND3_X1 U16164 ( .A1(n14232), .A2(n14167), .A3(n14166), .ZN(n14168) );
  NAND4_X1 U16165 ( .A1(n14171), .A2(n14170), .A3(n14169), .A4(n14168), .ZN(
        P1_U3247) );
  OAI211_X1 U16166 ( .C1(n14173), .C2(n14172), .A(n14233), .B(n14187), .ZN(
        n14184) );
  MUX2_X1 U16167 ( .A(n14174), .B(P1_REG2_REG_6__SCAN_IN), .S(n14179), .Z(
        n14177) );
  NAND3_X1 U16168 ( .A1(n14177), .A2(n14176), .A3(n14175), .ZN(n14178) );
  NAND3_X1 U16169 ( .A1(n14232), .A2(n14192), .A3(n14178), .ZN(n14183) );
  NAND2_X1 U16170 ( .A1(n14206), .A2(n14179), .ZN(n14182) );
  AOI21_X1 U16171 ( .B1(n14212), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n14180), .ZN(
        n14181) );
  NAND4_X1 U16172 ( .A1(n14184), .A2(n14183), .A3(n14182), .A4(n14181), .ZN(
        P1_U3249) );
  MUX2_X1 U16173 ( .A(n10802), .B(P1_REG1_REG_7__SCAN_IN), .S(n14194), .Z(
        n14185) );
  NAND3_X1 U16174 ( .A1(n14187), .A2(n14186), .A3(n14185), .ZN(n14188) );
  NAND3_X1 U16175 ( .A1(n14233), .A2(n14189), .A3(n14188), .ZN(n14199) );
  MUX2_X1 U16176 ( .A(n10783), .B(P1_REG2_REG_7__SCAN_IN), .S(n14194), .Z(
        n14190) );
  NAND3_X1 U16177 ( .A1(n14192), .A2(n14191), .A3(n14190), .ZN(n14193) );
  NAND3_X1 U16178 ( .A1(n14232), .A2(n14202), .A3(n14193), .ZN(n14198) );
  NAND2_X1 U16179 ( .A1(n14206), .A2(n14194), .ZN(n14197) );
  AOI21_X1 U16180 ( .B1(n14212), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n14195), .ZN(
        n14196) );
  NAND4_X1 U16181 ( .A1(n14199), .A2(n14198), .A3(n14197), .A4(n14196), .ZN(
        P1_U3250) );
  MUX2_X1 U16182 ( .A(n11733), .B(P1_REG2_REG_8__SCAN_IN), .S(n14205), .Z(
        n14200) );
  NAND3_X1 U16183 ( .A1(n14202), .A2(n14201), .A3(n14200), .ZN(n14203) );
  NAND3_X1 U16184 ( .A1(n14232), .A2(n14204), .A3(n14203), .ZN(n14216) );
  NAND2_X1 U16185 ( .A1(n14206), .A2(n14205), .ZN(n14215) );
  OAI21_X1 U16186 ( .B1(n14209), .B2(n14208), .A(n14207), .ZN(n14210) );
  NAND2_X1 U16187 ( .A1(n14233), .A2(n14210), .ZN(n14214) );
  NOR2_X1 U16188 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9977), .ZN(n14211) );
  AOI21_X1 U16189 ( .B1(n14212), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n14211), .ZN(
        n14213) );
  NAND4_X1 U16190 ( .A1(n14216), .A2(n14215), .A3(n14214), .A4(n14213), .ZN(
        P1_U3251) );
  INV_X1 U16191 ( .A(n14217), .ZN(n14218) );
  NAND2_X1 U16192 ( .A1(n14218), .A2(n14222), .ZN(n14219) );
  NAND2_X1 U16193 ( .A1(n14220), .A2(n14219), .ZN(n14221) );
  XOR2_X1 U16194 ( .A(n14221), .B(P1_REG1_REG_19__SCAN_IN), .Z(n14234) );
  INV_X1 U16195 ( .A(n14234), .ZN(n14230) );
  NAND2_X1 U16196 ( .A1(n14223), .A2(n14222), .ZN(n14227) );
  OR2_X1 U16197 ( .A1(n14225), .A2(n14224), .ZN(n14226) );
  NAND2_X1 U16198 ( .A1(n14227), .A2(n14226), .ZN(n14228) );
  XOR2_X1 U16199 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n14228), .Z(n14231) );
  OAI21_X1 U16200 ( .B1(n14231), .B2(n14972), .A(n14976), .ZN(n14229) );
  AOI21_X1 U16201 ( .B1(n14230), .B2(n14233), .A(n14229), .ZN(n14237) );
  AOI22_X1 U16202 ( .A1(n14234), .A2(n14233), .B1(n14232), .B2(n14231), .ZN(
        n14236) );
  MUX2_X1 U16203 ( .A(n14237), .B(n14236), .S(n14235), .Z(n14239) );
  OAI211_X1 U16204 ( .C1(n14240), .C2(n14980), .A(n14239), .B(n14238), .ZN(
        P1_U3262) );
  NOR2_X2 U16205 ( .A1(n14260), .A2(n14261), .ZN(n14259) );
  NAND2_X1 U16206 ( .A1(n14259), .A2(n14507), .ZN(n14242) );
  XNOR2_X1 U16207 ( .A(n14242), .B(n14504), .ZN(n14243) );
  NAND2_X1 U16208 ( .A1(n14243), .A2(n11131), .ZN(n14503) );
  NOR2_X1 U16209 ( .A1(n14629), .A2(n14244), .ZN(n14245) );
  NOR2_X1 U16210 ( .A1(n14464), .A2(n14245), .ZN(n14263) );
  NAND2_X1 U16211 ( .A1(n14263), .A2(n14246), .ZN(n14505) );
  NOR2_X1 U16212 ( .A1(n6550), .A2(n14505), .ZN(n14252) );
  NOR2_X1 U16213 ( .A1(n14504), .A2(n15009), .ZN(n14247) );
  AOI211_X1 U16214 ( .C1(P1_REG2_REG_31__SCAN_IN), .C2(n6550), .A(n14252), .B(
        n14247), .ZN(n14248) );
  OAI21_X1 U16215 ( .B1(n14503), .B2(n14383), .A(n14248), .ZN(P1_U3263) );
  XNOR2_X1 U16216 ( .A(n14259), .B(n14249), .ZN(n14250) );
  NAND2_X1 U16217 ( .A1(n14250), .A2(n11131), .ZN(n14506) );
  NOR2_X1 U16218 ( .A1(n14507), .A2(n15009), .ZN(n14251) );
  AOI211_X1 U16219 ( .C1(n6550), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14252), .B(
        n14251), .ZN(n14253) );
  OAI21_X1 U16220 ( .B1(n14506), .B2(n14383), .A(n14253), .ZN(P1_U3264) );
  NAND2_X1 U16221 ( .A1(n14256), .A2(n14255), .ZN(n14258) );
  XNOR2_X1 U16222 ( .A(n14258), .B(n7449), .ZN(n14508) );
  INV_X1 U16223 ( .A(n14261), .ZN(n14511) );
  AOI211_X1 U16224 ( .C1(n14261), .C2(n14260), .A(n15014), .B(n14259), .ZN(
        n14513) );
  NAND2_X1 U16225 ( .A1(n14513), .A2(n15017), .ZN(n14270) );
  NAND2_X1 U16226 ( .A1(n14263), .A2(n14262), .ZN(n14510) );
  OAI22_X1 U16227 ( .A1(n14265), .A2(n14510), .B1(n14264), .B2(n15005), .ZN(
        n14268) );
  NAND2_X1 U16228 ( .A1(n14266), .A2(n14479), .ZN(n14509) );
  NOR2_X1 U16229 ( .A1(n6550), .A2(n14509), .ZN(n14267) );
  AOI211_X1 U16230 ( .C1(n6550), .C2(P1_REG2_REG_29__SCAN_IN), .A(n14268), .B(
        n14267), .ZN(n14269) );
  OAI211_X1 U16231 ( .C1(n14511), .C2(n15009), .A(n14270), .B(n14269), .ZN(
        n14271) );
  AOI21_X1 U16232 ( .B1(n14394), .B2(n14508), .A(n14271), .ZN(n14272) );
  OAI21_X1 U16233 ( .B1(n14515), .B2(n14490), .A(n14272), .ZN(P1_U3356) );
  OAI22_X1 U16234 ( .A1(n14275), .A2(n14462), .B1(n14274), .B2(n14464), .ZN(
        n14280) );
  AOI21_X1 U16235 ( .B1(n14278), .B2(n14277), .A(n14276), .ZN(n14279) );
  INV_X1 U16236 ( .A(n14293), .ZN(n14282) );
  AOI211_X1 U16237 ( .C1(n14522), .C2(n14282), .A(n15014), .B(n14281), .ZN(
        n14521) );
  INV_X1 U16238 ( .A(n14283), .ZN(n14284) );
  AOI22_X1 U16239 ( .A1(n6550), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n14284), 
        .B2(n14888), .ZN(n14285) );
  OAI21_X1 U16240 ( .B1(n14286), .B2(n15009), .A(n14285), .ZN(n14289) );
  INV_X1 U16241 ( .A(n14287), .ZN(n14525) );
  NOR2_X1 U16242 ( .A1(n14525), .A2(n14437), .ZN(n14288) );
  AOI211_X1 U16243 ( .C1(n14521), .C2(n15017), .A(n14289), .B(n14288), .ZN(
        n14290) );
  OAI21_X1 U16244 ( .B1(n14524), .B2(n6550), .A(n14290), .ZN(P1_U3266) );
  XOR2_X1 U16245 ( .A(n14291), .B(n14300), .Z(n14526) );
  INV_X1 U16246 ( .A(n14526), .ZN(n14307) );
  OAI21_X1 U16247 ( .B1(n14297), .B2(n14314), .A(n11131), .ZN(n14292) );
  OR2_X1 U16248 ( .A1(n14293), .A2(n14292), .ZN(n14527) );
  INV_X1 U16249 ( .A(n14527), .ZN(n14305) );
  NOR2_X1 U16250 ( .A1(n15005), .A2(n14294), .ZN(n14295) );
  AOI21_X1 U16251 ( .B1(n6550), .B2(P1_REG2_REG_26__SCAN_IN), .A(n14295), .ZN(
        n14296) );
  OAI21_X1 U16252 ( .B1(n14297), .B2(n15009), .A(n14296), .ZN(n14304) );
  OAI21_X1 U16253 ( .B1(n14300), .B2(n14299), .A(n14298), .ZN(n14302) );
  AOI222_X1 U16254 ( .A1(n15052), .A2(n14302), .B1(n14301), .B2(n14477), .C1(
        n14325), .C2(n14479), .ZN(n14530) );
  NOR2_X1 U16255 ( .A1(n14530), .A2(n6550), .ZN(n14303) );
  AOI211_X1 U16256 ( .C1(n14305), .C2(n15017), .A(n14304), .B(n14303), .ZN(
        n14306) );
  OAI21_X1 U16257 ( .B1(n14490), .B2(n14307), .A(n14306), .ZN(P1_U3267) );
  OAI21_X1 U16258 ( .B1(n7945), .B2(n12592), .A(n14308), .ZN(n14538) );
  OAI21_X1 U16259 ( .B1(n14311), .B2(n14310), .A(n14309), .ZN(n14531) );
  NAND2_X1 U16260 ( .A1(n14531), .A2(n14394), .ZN(n14322) );
  NAND2_X1 U16261 ( .A1(n14535), .A2(n14332), .ZN(n14312) );
  NAND2_X1 U16262 ( .A1(n14312), .A2(n11131), .ZN(n14313) );
  NOR2_X1 U16263 ( .A1(n14314), .A2(n14313), .ZN(n14533) );
  OAI21_X1 U16264 ( .B1(n15005), .B2(n14315), .A(n14532), .ZN(n14316) );
  INV_X1 U16265 ( .A(n14316), .ZN(n14319) );
  NAND2_X1 U16266 ( .A1(n14535), .A2(n14889), .ZN(n14318) );
  NAND2_X1 U16267 ( .A1(n6550), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n14317) );
  OAI211_X1 U16268 ( .C1(n6550), .C2(n14319), .A(n14318), .B(n14317), .ZN(
        n14320) );
  AOI21_X1 U16269 ( .B1(n14533), .B2(n15017), .A(n14320), .ZN(n14321) );
  OAI211_X1 U16270 ( .C1(n14538), .C2(n14490), .A(n14322), .B(n14321), .ZN(
        P1_U3268) );
  OAI21_X1 U16271 ( .B1(n14329), .B2(n14324), .A(n14323), .ZN(n14541) );
  INV_X1 U16272 ( .A(n14325), .ZN(n14326) );
  OAI22_X1 U16273 ( .A1(n7703), .A2(n14462), .B1(n14326), .B2(n14464), .ZN(
        n14331) );
  AOI211_X1 U16274 ( .C1(n14329), .C2(n14328), .A(n15002), .B(n14327), .ZN(
        n14330) );
  AOI211_X1 U16275 ( .C1(n15059), .C2(n14541), .A(n14331), .B(n14330), .ZN(
        n14543) );
  INV_X1 U16276 ( .A(n14437), .ZN(n15018) );
  INV_X1 U16277 ( .A(n14332), .ZN(n14333) );
  AOI211_X1 U16278 ( .C1(n14334), .C2(n14346), .A(n15014), .B(n14333), .ZN(
        n14539) );
  NAND2_X1 U16279 ( .A1(n14539), .A2(n15017), .ZN(n14338) );
  INV_X1 U16280 ( .A(n14335), .ZN(n14336) );
  AOI22_X1 U16281 ( .A1(n6550), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14336), 
        .B2(n14888), .ZN(n14337) );
  OAI211_X1 U16282 ( .C1(n14339), .C2(n15009), .A(n14338), .B(n14337), .ZN(
        n14340) );
  AOI21_X1 U16283 ( .B1(n15018), .B2(n14541), .A(n14340), .ZN(n14341) );
  OAI21_X1 U16284 ( .B1(n14543), .B2(n6550), .A(n14341), .ZN(P1_U3269) );
  XNOR2_X1 U16285 ( .A(n14342), .B(n14344), .ZN(n14550) );
  OAI21_X1 U16286 ( .B1(n14345), .B2(n14344), .A(n14343), .ZN(n14548) );
  AOI21_X1 U16287 ( .B1(n14352), .B2(n14364), .A(n15014), .ZN(n14347) );
  NAND2_X1 U16288 ( .A1(n14347), .A2(n14346), .ZN(n14545) );
  NOR2_X1 U16289 ( .A1(n15005), .A2(n14348), .ZN(n14349) );
  AOI21_X1 U16290 ( .B1(n6550), .B2(P1_REG2_REG_23__SCAN_IN), .A(n14349), .ZN(
        n14350) );
  OAI21_X1 U16291 ( .B1(n14544), .B2(n6550), .A(n14350), .ZN(n14351) );
  AOI21_X1 U16292 ( .B1(n14352), .B2(n14889), .A(n14351), .ZN(n14353) );
  OAI21_X1 U16293 ( .B1(n14545), .B2(n14383), .A(n14353), .ZN(n14354) );
  AOI21_X1 U16294 ( .B1(n14548), .B2(n14394), .A(n14354), .ZN(n14355) );
  OAI21_X1 U16295 ( .B1(n14490), .B2(n14550), .A(n14355), .ZN(P1_U3270) );
  XNOR2_X1 U16296 ( .A(n14362), .B(n14356), .ZN(n14357) );
  AOI22_X1 U16297 ( .A1(n14359), .A2(n14479), .B1(n14477), .B2(n14358), .ZN(
        n14360) );
  XNOR2_X1 U16298 ( .A(n14363), .B(n14362), .ZN(n14555) );
  AOI21_X1 U16299 ( .B1(n14551), .B2(n14376), .A(n15014), .ZN(n14365) );
  NAND2_X1 U16300 ( .A1(n14365), .A2(n14364), .ZN(n14553) );
  AOI22_X1 U16301 ( .A1(n6550), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n14366), 
        .B2(n14888), .ZN(n14368) );
  NAND2_X1 U16302 ( .A1(n14551), .A2(n14889), .ZN(n14367) );
  OAI211_X1 U16303 ( .C1(n14553), .C2(n14383), .A(n14368), .B(n14367), .ZN(
        n14369) );
  AOI21_X1 U16304 ( .B1(n14555), .B2(n14898), .A(n14369), .ZN(n14370) );
  OAI21_X1 U16305 ( .B1(n14556), .B2(n6550), .A(n14370), .ZN(P1_U3271) );
  XNOR2_X1 U16306 ( .A(n14372), .B(n14371), .ZN(n14564) );
  OAI21_X1 U16307 ( .B1(n14375), .B2(n14374), .A(n14373), .ZN(n14562) );
  INV_X1 U16308 ( .A(n14395), .ZN(n14377) );
  OAI211_X1 U16309 ( .C1(n14560), .C2(n14377), .A(n14376), .B(n11131), .ZN(
        n14559) );
  OAI21_X1 U16310 ( .B1(n14378), .B2(n15005), .A(n14558), .ZN(n14379) );
  MUX2_X1 U16311 ( .A(n14379), .B(P1_REG2_REG_21__SCAN_IN), .S(n6550), .Z(
        n14380) );
  AOI21_X1 U16312 ( .B1(n14381), .B2(n14889), .A(n14380), .ZN(n14382) );
  OAI21_X1 U16313 ( .B1(n14559), .B2(n14383), .A(n14382), .ZN(n14384) );
  AOI21_X1 U16314 ( .B1(n14562), .B2(n14898), .A(n14384), .ZN(n14385) );
  OAI21_X1 U16315 ( .B1(n14386), .B2(n14564), .A(n14385), .ZN(P1_U3272) );
  INV_X1 U16316 ( .A(n14387), .ZN(n14389) );
  OAI21_X1 U16317 ( .B1(n14389), .B2(n14393), .A(n14388), .ZN(n14572) );
  INV_X1 U16318 ( .A(n14390), .ZN(n14391) );
  AOI21_X1 U16319 ( .B1(n14393), .B2(n14392), .A(n14391), .ZN(n14570) );
  NAND2_X1 U16320 ( .A1(n14570), .A2(n14394), .ZN(n14405) );
  OAI21_X1 U16321 ( .B1(n14401), .B2(n6696), .A(n14395), .ZN(n14568) );
  OAI22_X1 U16322 ( .A1(n14396), .A2(n14464), .B1(n14427), .B2(n14462), .ZN(
        n14565) );
  AOI21_X1 U16323 ( .B1(n14397), .B2(n14888), .A(n14565), .ZN(n14398) );
  OAI21_X1 U16324 ( .B1(n14568), .B2(n14399), .A(n14398), .ZN(n14403) );
  INV_X1 U16325 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14400) );
  OAI22_X1 U16326 ( .A1(n14401), .A2(n15009), .B1(n14400), .B2(n14498), .ZN(
        n14402) );
  AOI21_X1 U16327 ( .B1(n14403), .B2(n14498), .A(n14402), .ZN(n14404) );
  OAI211_X1 U16328 ( .C1(n14572), .C2(n14490), .A(n14405), .B(n14404), .ZN(
        P1_U3273) );
  XNOR2_X1 U16329 ( .A(n14407), .B(n14406), .ZN(n14410) );
  AOI222_X1 U16330 ( .A1(n15052), .A2(n14410), .B1(n14409), .B2(n14477), .C1(
        n14408), .C2(n14479), .ZN(n14576) );
  AOI211_X1 U16331 ( .C1(n14574), .C2(n14429), .A(n15014), .B(n6696), .ZN(
        n14573) );
  INV_X1 U16332 ( .A(n14411), .ZN(n14412) );
  AOI22_X1 U16333 ( .A1(n6550), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14412), 
        .B2(n14888), .ZN(n14413) );
  OAI21_X1 U16334 ( .B1(n14414), .B2(n15009), .A(n14413), .ZN(n14418) );
  XNOR2_X1 U16335 ( .A(n14416), .B(n14415), .ZN(n14577) );
  NOR2_X1 U16336 ( .A1(n14577), .A2(n14490), .ZN(n14417) );
  AOI211_X1 U16337 ( .C1(n14573), .C2(n15017), .A(n14418), .B(n14417), .ZN(
        n14419) );
  OAI21_X1 U16338 ( .B1(n14576), .B2(n6550), .A(n14419), .ZN(P1_U3274) );
  XNOR2_X1 U16339 ( .A(n14421), .B(n14420), .ZN(n14426) );
  INV_X1 U16340 ( .A(n14426), .ZN(n14583) );
  XNOR2_X1 U16341 ( .A(n14423), .B(n14422), .ZN(n14424) );
  AOI222_X1 U16342 ( .A1(n14426), .A2(n15059), .B1(n14425), .B2(n14479), .C1(
        n15052), .C2(n14424), .ZN(n14582) );
  INV_X1 U16343 ( .A(n14582), .ZN(n14428) );
  NOR2_X1 U16344 ( .A1(n14427), .A2(n14464), .ZN(n14579) );
  OAI21_X1 U16345 ( .B1(n14428), .B2(n14579), .A(n14498), .ZN(n14436) );
  INV_X1 U16346 ( .A(n14429), .ZN(n14430) );
  AOI211_X1 U16347 ( .C1(n14580), .C2(n14439), .A(n15014), .B(n14430), .ZN(
        n14578) );
  AOI22_X1 U16348 ( .A1(n6550), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14431), 
        .B2(n14888), .ZN(n14432) );
  OAI21_X1 U16349 ( .B1(n14433), .B2(n15009), .A(n14432), .ZN(n14434) );
  AOI21_X1 U16350 ( .B1(n14578), .B2(n15017), .A(n14434), .ZN(n14435) );
  OAI211_X1 U16351 ( .C1(n14583), .C2(n14437), .A(n14436), .B(n14435), .ZN(
        P1_U3275) );
  XOR2_X1 U16352 ( .A(n14438), .B(n14445), .Z(n14588) );
  INV_X1 U16353 ( .A(n14467), .ZN(n14441) );
  INV_X1 U16354 ( .A(n14439), .ZN(n14440) );
  AOI211_X1 U16355 ( .C1(n14585), .C2(n14441), .A(n15014), .B(n14440), .ZN(
        n14584) );
  AOI22_X1 U16356 ( .A1(n6550), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n14442), 
        .B2(n14888), .ZN(n14443) );
  OAI21_X1 U16357 ( .B1(n14444), .B2(n15009), .A(n14443), .ZN(n14453) );
  AOI21_X1 U16358 ( .B1(n14446), .B2(n14445), .A(n15002), .ZN(n14451) );
  OAI22_X1 U16359 ( .A1(n14448), .A2(n14464), .B1(n14447), .B2(n14462), .ZN(
        n14449) );
  AOI21_X1 U16360 ( .B1(n14451), .B2(n14450), .A(n14449), .ZN(n14587) );
  NOR2_X1 U16361 ( .A1(n14587), .A2(n6550), .ZN(n14452) );
  AOI211_X1 U16362 ( .C1(n14584), .C2(n15017), .A(n14453), .B(n14452), .ZN(
        n14454) );
  OAI21_X1 U16363 ( .B1(n14490), .B2(n14588), .A(n14454), .ZN(P1_U3276) );
  XOR2_X1 U16364 ( .A(n14455), .B(n14459), .Z(n14593) );
  INV_X1 U16365 ( .A(n14456), .ZN(n14457) );
  AOI21_X1 U16366 ( .B1(n14459), .B2(n14458), .A(n14457), .ZN(n14460) );
  OAI222_X1 U16367 ( .A1(n14464), .A2(n14463), .B1(n14462), .B2(n14461), .C1(
        n15002), .C2(n14460), .ZN(n14589) );
  NAND2_X1 U16368 ( .A1(n14589), .A2(n14498), .ZN(n14474) );
  NAND2_X1 U16369 ( .A1(n14482), .A2(n14591), .ZN(n14465) );
  NAND2_X1 U16370 ( .A1(n14465), .A2(n11131), .ZN(n14466) );
  NOR2_X1 U16371 ( .A1(n14467), .A2(n14466), .ZN(n14590) );
  NOR2_X1 U16372 ( .A1(n14468), .A2(n15009), .ZN(n14472) );
  OAI22_X1 U16373 ( .A1(n14498), .A2(n14470), .B1(n14469), .B2(n15005), .ZN(
        n14471) );
  AOI211_X1 U16374 ( .C1(n14590), .C2(n15017), .A(n14472), .B(n14471), .ZN(
        n14473) );
  OAI211_X1 U16375 ( .C1(n14593), .C2(n14490), .A(n14474), .B(n14473), .ZN(
        P1_U3277) );
  XNOR2_X1 U16376 ( .A(n14476), .B(n14475), .ZN(n14481) );
  AOI222_X1 U16377 ( .A1(n15052), .A2(n14481), .B1(n14480), .B2(n14479), .C1(
        n14478), .C2(n14477), .ZN(n14597) );
  INV_X1 U16378 ( .A(n14482), .ZN(n14483) );
  AOI211_X1 U16379 ( .C1(n14595), .C2(n14484), .A(n15014), .B(n14483), .ZN(
        n14594) );
  INV_X1 U16380 ( .A(n14485), .ZN(n14486) );
  AOI22_X1 U16381 ( .A1(n6550), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n14486), 
        .B2(n14888), .ZN(n14487) );
  OAI21_X1 U16382 ( .B1(n7116), .B2(n15009), .A(n14487), .ZN(n14492) );
  AOI21_X1 U16383 ( .B1(n14489), .B2(n14488), .A(n6707), .ZN(n14598) );
  NOR2_X1 U16384 ( .A1(n14598), .A2(n14490), .ZN(n14491) );
  AOI211_X1 U16385 ( .C1(n14594), .C2(n15017), .A(n14492), .B(n14491), .ZN(
        n14493) );
  OAI21_X1 U16386 ( .B1(n6550), .B2(n14597), .A(n14493), .ZN(P1_U3278) );
  AOI22_X1 U16387 ( .A1(n15018), .A2(n14495), .B1(n14889), .B2(n14494), .ZN(
        n14502) );
  AOI22_X1 U16388 ( .A1(n15017), .A2(n14496), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n14888), .ZN(n14501) );
  NAND2_X1 U16389 ( .A1(n14498), .A2(n14497), .ZN(n14500) );
  NAND2_X1 U16390 ( .A1(n6550), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n14499) );
  NAND4_X1 U16391 ( .A1(n14502), .A2(n14501), .A3(n14500), .A4(n14499), .ZN(
        P1_U3292) );
  OAI211_X1 U16392 ( .C1(n14902), .C2(n14504), .A(n14503), .B(n14505), .ZN(
        n14600) );
  MUX2_X1 U16393 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14600), .S(n15107), .Z(
        P1_U3559) );
  OAI211_X1 U16394 ( .C1(n14902), .C2(n14507), .A(n14506), .B(n14505), .ZN(
        n14601) );
  MUX2_X1 U16395 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14601), .S(n15107), .Z(
        P1_U3558) );
  OAI211_X1 U16396 ( .C1(n14511), .C2(n14902), .A(n14510), .B(n14509), .ZN(
        n14512) );
  AOI21_X1 U16397 ( .B1(n14517), .B2(n14951), .A(n14516), .ZN(n14518) );
  OAI211_X1 U16398 ( .C1(n14599), .C2(n14520), .A(n14519), .B(n14518), .ZN(
        n14602) );
  MUX2_X1 U16399 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14602), .S(n15107), .Z(
        P1_U3556) );
  AOI21_X1 U16400 ( .B1(n14522), .B2(n14951), .A(n14521), .ZN(n14523) );
  NAND2_X1 U16401 ( .A1(n14526), .A2(n15093), .ZN(n14529) );
  NAND4_X1 U16402 ( .A1(n14530), .A2(n14529), .A3(n14528), .A4(n14527), .ZN(
        n14604) );
  MUX2_X1 U16403 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14604), .S(n15107), .Z(
        P1_U3554) );
  NAND2_X1 U16404 ( .A1(n14531), .A2(n15052), .ZN(n14537) );
  INV_X1 U16405 ( .A(n14532), .ZN(n14534) );
  AOI211_X1 U16406 ( .C1(n14535), .C2(n14951), .A(n14534), .B(n14533), .ZN(
        n14536) );
  OAI211_X1 U16407 ( .C1(n14599), .C2(n14538), .A(n14537), .B(n14536), .ZN(
        n14605) );
  MUX2_X1 U16408 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14605), .S(n15107), .Z(
        P1_U3553) );
  INV_X1 U16409 ( .A(n15055), .ZN(n15084) );
  AOI211_X1 U16410 ( .C1(n15084), .C2(n14541), .A(n14540), .B(n14539), .ZN(
        n14542) );
  NAND2_X1 U16411 ( .A1(n14543), .A2(n14542), .ZN(n14606) );
  MUX2_X1 U16412 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14606), .S(n15107), .Z(
        P1_U3552) );
  OAI211_X1 U16413 ( .C1(n14546), .C2(n14902), .A(n14545), .B(n14544), .ZN(
        n14547) );
  AOI21_X1 U16414 ( .B1(n14548), .B2(n15052), .A(n14547), .ZN(n14549) );
  OAI21_X1 U16415 ( .B1(n14599), .B2(n14550), .A(n14549), .ZN(n14607) );
  MUX2_X1 U16416 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14607), .S(n15107), .Z(
        P1_U3551) );
  NAND2_X1 U16417 ( .A1(n14551), .A2(n14951), .ZN(n14552) );
  NAND2_X1 U16418 ( .A1(n14553), .A2(n14552), .ZN(n14554) );
  AOI21_X1 U16419 ( .B1(n14555), .B2(n15093), .A(n14554), .ZN(n14557) );
  NAND2_X1 U16420 ( .A1(n14557), .A2(n14556), .ZN(n14608) );
  MUX2_X1 U16421 ( .A(n14608), .B(P1_REG1_REG_22__SCAN_IN), .S(n15105), .Z(
        P1_U3550) );
  OAI211_X1 U16422 ( .C1(n14560), .C2(n14902), .A(n14559), .B(n14558), .ZN(
        n14561) );
  AOI21_X1 U16423 ( .B1(n14562), .B2(n15093), .A(n14561), .ZN(n14563) );
  OAI21_X1 U16424 ( .B1(n15002), .B2(n14564), .A(n14563), .ZN(n14609) );
  MUX2_X1 U16425 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14609), .S(n15107), .Z(
        P1_U3549) );
  AOI21_X1 U16426 ( .B1(n14566), .B2(n14951), .A(n14565), .ZN(n14567) );
  OAI21_X1 U16427 ( .B1(n14568), .B2(n15014), .A(n14567), .ZN(n14569) );
  AOI21_X1 U16428 ( .B1(n14570), .B2(n15052), .A(n14569), .ZN(n14571) );
  OAI21_X1 U16429 ( .B1(n14599), .B2(n14572), .A(n14571), .ZN(n14610) );
  MUX2_X1 U16430 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14610), .S(n15107), .Z(
        P1_U3548) );
  AOI21_X1 U16431 ( .B1(n14574), .B2(n14951), .A(n14573), .ZN(n14575) );
  OAI211_X1 U16432 ( .C1(n14599), .C2(n14577), .A(n14576), .B(n14575), .ZN(
        n14611) );
  MUX2_X1 U16433 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14611), .S(n15107), .Z(
        P1_U3547) );
  AOI211_X1 U16434 ( .C1(n14580), .C2(n14951), .A(n14579), .B(n14578), .ZN(
        n14581) );
  OAI211_X1 U16435 ( .C1(n14583), .C2(n15055), .A(n14582), .B(n14581), .ZN(
        n14612) );
  MUX2_X1 U16436 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14612), .S(n15107), .Z(
        P1_U3546) );
  AOI21_X1 U16437 ( .B1(n14585), .B2(n14951), .A(n14584), .ZN(n14586) );
  OAI211_X1 U16438 ( .C1(n14588), .C2(n14599), .A(n14587), .B(n14586), .ZN(
        n14613) );
  MUX2_X1 U16439 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14613), .S(n15107), .Z(
        P1_U3545) );
  AOI211_X1 U16440 ( .C1(n14591), .C2(n14951), .A(n14590), .B(n14589), .ZN(
        n14592) );
  OAI21_X1 U16441 ( .B1(n14599), .B2(n14593), .A(n14592), .ZN(n14614) );
  MUX2_X1 U16442 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14614), .S(n15107), .Z(
        P1_U3544) );
  AOI21_X1 U16443 ( .B1(n14595), .B2(n14951), .A(n14594), .ZN(n14596) );
  OAI211_X1 U16444 ( .C1(n14599), .C2(n14598), .A(n14597), .B(n14596), .ZN(
        n14615) );
  MUX2_X1 U16445 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n14615), .S(n15107), .Z(
        P1_U3543) );
  MUX2_X1 U16446 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14600), .S(n15096), .Z(
        P1_U3527) );
  MUX2_X1 U16447 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14601), .S(n15096), .Z(
        P1_U3526) );
  MUX2_X1 U16448 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14602), .S(n15096), .Z(
        P1_U3524) );
  MUX2_X1 U16449 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14603), .S(n15096), .Z(
        P1_U3523) );
  MUX2_X1 U16450 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14604), .S(n15096), .Z(
        P1_U3522) );
  MUX2_X1 U16451 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14605), .S(n15096), .Z(
        P1_U3521) );
  MUX2_X1 U16452 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14606), .S(n15096), .Z(
        P1_U3520) );
  MUX2_X1 U16453 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14607), .S(n15096), .Z(
        P1_U3519) );
  MUX2_X1 U16454 ( .A(n14608), .B(P1_REG0_REG_22__SCAN_IN), .S(n7451), .Z(
        P1_U3518) );
  MUX2_X1 U16455 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14609), .S(n15096), .Z(
        P1_U3517) );
  MUX2_X1 U16456 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14610), .S(n15096), .Z(
        P1_U3516) );
  MUX2_X1 U16457 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14611), .S(n15096), .Z(
        P1_U3515) );
  MUX2_X1 U16458 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14612), .S(n15096), .Z(
        P1_U3513) );
  MUX2_X1 U16459 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14613), .S(n15096), .Z(
        P1_U3510) );
  MUX2_X1 U16460 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14614), .S(n15096), .Z(
        P1_U3507) );
  MUX2_X1 U16461 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n14615), .S(n15096), .Z(
        P1_U3504) );
  INV_X1 U16462 ( .A(n14616), .ZN(n14618) );
  NOR4_X1 U16463 ( .A1(n14618), .A2(P1_IR_REG_30__SCAN_IN), .A3(n14617), .A4(
        P1_U3086), .ZN(n14619) );
  AOI21_X1 U16464 ( .B1(n14620), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14619), 
        .ZN(n14621) );
  OAI21_X1 U16465 ( .B1(n14622), .B2(n14638), .A(n14621), .ZN(P1_U3324) );
  OAI222_X1 U16466 ( .A1(n14638), .A2(n14624), .B1(P1_U3086), .B2(n14623), 
        .C1(n15515), .C2(n14635), .ZN(P1_U3325) );
  OAI222_X1 U16467 ( .A1(n14635), .A2(n14628), .B1(n14638), .B2(n14627), .C1(
        n14626), .C2(P1_U3086), .ZN(P1_U3326) );
  INV_X1 U16468 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14631) );
  OAI222_X1 U16469 ( .A1(n14635), .A2(n14631), .B1(n14638), .B2(n14630), .C1(
        P1_U3086), .C2(n14629), .ZN(P1_U3328) );
  OAI222_X1 U16470 ( .A1(P1_U3086), .A2(n14634), .B1(n14638), .B2(n14633), 
        .C1(n14632), .C2(n14635), .ZN(P1_U3329) );
  OAI222_X1 U16471 ( .A1(P1_U3086), .A2(n14639), .B1(n14638), .B2(n14637), 
        .C1(n14636), .C2(n14635), .ZN(P1_U3331) );
  MUX2_X1 U16472 ( .A(n14641), .B(n14640), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16473 ( .A(n14642), .ZN(n14643) );
  MUX2_X1 U16474 ( .A(n14643), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16475 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14671) );
  INV_X1 U16476 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14644) );
  NOR2_X1 U16477 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14644), .ZN(n14670) );
  INV_X1 U16478 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14981) );
  NOR2_X1 U16479 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14981), .ZN(n14669) );
  XOR2_X1 U16480 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(n14667), .Z(n14677) );
  INV_X1 U16481 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14665) );
  XOR2_X1 U16482 ( .A(n15455), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n14678) );
  INV_X1 U16483 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14662) );
  INV_X1 U16484 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14658) );
  INV_X1 U16485 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14656) );
  XOR2_X1 U16486 ( .A(n14656), .B(P1_ADDR_REG_9__SCAN_IN), .Z(n14680) );
  XOR2_X1 U16487 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), .Z(
        n14689) );
  NOR2_X1 U16488 ( .A1(n14648), .A2(n10920), .ZN(n14650) );
  NOR2_X1 U16489 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14652), .ZN(n14653) );
  XOR2_X1 U16490 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n14652), .Z(n14705) );
  XNOR2_X1 U16491 ( .A(n15566), .B(P1_ADDR_REG_8__SCAN_IN), .ZN(n14708) );
  NOR2_X1 U16492 ( .A1(n14658), .A2(n14657), .ZN(n14660) );
  XNOR2_X1 U16493 ( .A(n14662), .B(P1_ADDR_REG_11__SCAN_IN), .ZN(n14716) );
  NAND2_X1 U16494 ( .A1(n14678), .A2(n14679), .ZN(n14663) );
  INV_X1 U16495 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14719) );
  NAND2_X1 U16496 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14719), .ZN(n14664) );
  NAND2_X1 U16497 ( .A1(n14677), .A2(n14676), .ZN(n14666) );
  INV_X1 U16498 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14668) );
  OAI22_X1 U16499 ( .A1(n14669), .A2(n14674), .B1(P1_ADDR_REG_15__SCAN_IN), 
        .B2(n14668), .ZN(n14673) );
  OAI22_X1 U16500 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n14671), .B1(n14670), 
        .B2(n14673), .ZN(n14728) );
  XNOR2_X1 U16501 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14728), .ZN(n14729) );
  XOR2_X1 U16502 ( .A(n14730), .B(n14729), .Z(n14791) );
  XNOR2_X1 U16503 ( .A(n14671), .B(P3_ADDR_REG_16__SCAN_IN), .ZN(n14672) );
  XNOR2_X1 U16504 ( .A(n14673), .B(n14672), .ZN(n14931) );
  XOR2_X1 U16505 ( .A(n14981), .B(P3_ADDR_REG_15__SCAN_IN), .Z(n14675) );
  XOR2_X1 U16506 ( .A(n14675), .B(n14674), .Z(n14725) );
  XNOR2_X1 U16507 ( .A(n14677), .B(n14676), .ZN(n14923) );
  XOR2_X1 U16508 ( .A(n14679), .B(n14678), .Z(n14916) );
  XOR2_X1 U16509 ( .A(n14681), .B(n14680), .Z(n14713) );
  NOR2_X1 U16510 ( .A1(n14683), .A2(n10442), .ZN(n14695) );
  NOR2_X1 U16511 ( .A1(n14687), .A2(n13529), .ZN(n14688) );
  AOI21_X1 U16512 ( .B1(n14685), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n14684), .ZN(
        n15740) );
  INV_X1 U16513 ( .A(n15740), .ZN(n14686) );
  NAND2_X1 U16514 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n14686), .ZN(n15748) );
  NOR2_X1 U16515 ( .A1(n15748), .A2(n15747), .ZN(n15746) );
  XOR2_X1 U16516 ( .A(n14690), .B(n14689), .Z(n14738) );
  XOR2_X1 U16517 ( .A(n14691), .B(P1_ADDR_REG_3__SCAN_IN), .Z(n14692) );
  NAND2_X1 U16518 ( .A1(n14693), .A2(n14692), .ZN(n14694) );
  NAND2_X1 U16519 ( .A1(n15745), .A2(n10459), .ZN(n15744) );
  NAND2_X1 U16520 ( .A1(n14694), .A2(n15744), .ZN(n15735) );
  NAND2_X1 U16521 ( .A1(n14697), .A2(n14698), .ZN(n14699) );
  INV_X1 U16522 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15738) );
  NOR2_X1 U16523 ( .A1(n14700), .A2(n7247), .ZN(n14703) );
  XOR2_X1 U16524 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n11071), .Z(n14702) );
  XNOR2_X1 U16525 ( .A(n14702), .B(n14701), .ZN(n14767) );
  NOR2_X1 U16526 ( .A1(n14706), .A2(n14704), .ZN(n14707) );
  XNOR2_X1 U16527 ( .A(n14705), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15743) );
  XNOR2_X1 U16528 ( .A(n14709), .B(n14708), .ZN(n14711) );
  NAND2_X1 U16529 ( .A1(n14710), .A2(n14711), .ZN(n14712) );
  INV_X1 U16530 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14773) );
  XNOR2_X1 U16531 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n14715), .ZN(n14775) );
  XNOR2_X1 U16532 ( .A(n14717), .B(n14716), .ZN(n14912) );
  NAND2_X1 U16533 ( .A1(n6581), .A2(n14912), .ZN(n14718) );
  XNOR2_X1 U16534 ( .A(n14719), .B(P1_ADDR_REG_13__SCAN_IN), .ZN(n14720) );
  XNOR2_X1 U16535 ( .A(n14721), .B(n14720), .ZN(n14723) );
  NAND2_X1 U16536 ( .A1(n14722), .A2(n14723), .ZN(n14724) );
  INV_X1 U16537 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14919) );
  INV_X1 U16538 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15165) );
  NAND2_X1 U16539 ( .A1(n14726), .A2(n14725), .ZN(n14928) );
  NAND2_X1 U16540 ( .A1(n14931), .A2(n14930), .ZN(n14929) );
  NOR2_X1 U16541 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14728), .ZN(n14732) );
  NOR2_X1 U16542 ( .A1(n14730), .A2(n14729), .ZN(n14731) );
  NOR2_X1 U16543 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n14800), .ZN(n14733) );
  AOI21_X1 U16544 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n14800), .A(n14733), 
        .ZN(n14798) );
  XOR2_X1 U16545 ( .A(n14797), .B(n14798), .Z(n14793) );
  INV_X1 U16546 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n15674) );
  NAND2_X1 U16547 ( .A1(n14734), .A2(n15674), .ZN(n14796) );
  OAI21_X1 U16548 ( .B1(n14734), .B2(n15674), .A(n14796), .ZN(SUB_1596_U62) );
  AOI21_X1 U16549 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14735) );
  OAI21_X1 U16550 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n14735), 
        .ZN(U28) );
  AOI21_X1 U16551 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14736) );
  OAI21_X1 U16552 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14736), 
        .ZN(U29) );
  AOI21_X1 U16553 ( .B1(n14739), .B2(n14738), .A(n14737), .ZN(n14740) );
  XOR2_X1 U16554 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n14740), .Z(SUB_1596_U61) );
  OAI22_X1 U16555 ( .A1(n14744), .A2(n14743), .B1(n14742), .B2(n14741), .ZN(
        n14745) );
  INV_X1 U16556 ( .A(n14745), .ZN(n14746) );
  OAI21_X1 U16557 ( .B1(P3_U3151), .B2(n14747), .A(n14746), .ZN(P3_U3289) );
  AOI22_X1 U16558 ( .A1(n14748), .A2(n14762), .B1(SI_3_), .B2(n14761), .ZN(
        n14749) );
  OAI21_X1 U16559 ( .B1(P3_U3151), .B2(n14750), .A(n14749), .ZN(P3_U3292) );
  AOI22_X1 U16560 ( .A1(n14751), .A2(n14762), .B1(n14761), .B2(SI_2_), .ZN(
        n14752) );
  OAI21_X1 U16561 ( .B1(P3_U3151), .B2(n6548), .A(n14752), .ZN(P3_U3293) );
  AOI22_X1 U16562 ( .A1(n14754), .A2(n14762), .B1(SI_10_), .B2(n14761), .ZN(
        n14755) );
  OAI21_X1 U16563 ( .B1(P3_U3151), .B2(n14756), .A(n14755), .ZN(P3_U3285) );
  INV_X1 U16564 ( .A(n14757), .ZN(n14758) );
  AOI22_X1 U16565 ( .A1(n14758), .A2(n14762), .B1(SI_11_), .B2(n14761), .ZN(
        n14759) );
  OAI21_X1 U16566 ( .B1(P3_U3151), .B2(n14760), .A(n14759), .ZN(P3_U3284) );
  AOI22_X1 U16567 ( .A1(n14763), .A2(n14762), .B1(SI_12_), .B2(n14761), .ZN(
        n14764) );
  OAI21_X1 U16568 ( .B1(P3_U3151), .B2(n14765), .A(n14764), .ZN(P3_U3283) );
  AOI21_X1 U16569 ( .B1(n14768), .B2(n14767), .A(n14766), .ZN(SUB_1596_U57) );
  OAI21_X1 U16570 ( .B1(n14770), .B2(n10601), .A(n14769), .ZN(SUB_1596_U55) );
  AOI21_X1 U16571 ( .B1(n14773), .B2(n14772), .A(n14771), .ZN(SUB_1596_U54) );
  AOI21_X1 U16572 ( .B1(n14776), .B2(n14775), .A(n14774), .ZN(n14777) );
  XOR2_X1 U16573 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14777), .Z(SUB_1596_U70)
         );
  NOR2_X1 U16574 ( .A1(n14778), .A2(n15002), .ZN(n14786) );
  OAI211_X1 U16575 ( .C1(n14781), .C2(n14902), .A(n14780), .B(n14779), .ZN(
        n14784) );
  AOI21_X1 U16576 ( .B1(n15081), .B2(n15055), .A(n14782), .ZN(n14783) );
  AOI211_X1 U16577 ( .C1(n14786), .C2(n14785), .A(n14784), .B(n14783), .ZN(
        n14788) );
  INV_X1 U16578 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n15554) );
  AOI22_X1 U16579 ( .A1(n15096), .A2(n14788), .B1(n15554), .B2(n7451), .ZN(
        P1_U3495) );
  AOI22_X1 U16580 ( .A1(n15107), .A2(n14788), .B1(n14787), .B2(n15105), .ZN(
        P1_U3540) );
  AOI21_X1 U16581 ( .B1(n14791), .B2(n14790), .A(n14789), .ZN(n14792) );
  XOR2_X1 U16582 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n14792), .Z(SUB_1596_U63)
         );
  NAND2_X1 U16583 ( .A1(n14794), .A2(n14793), .ZN(n14795) );
  NAND2_X1 U16584 ( .A1(n14796), .A2(n14795), .ZN(n14806) );
  NAND2_X1 U16585 ( .A1(n14798), .A2(n14797), .ZN(n14799) );
  OAI21_X1 U16586 ( .B1(n14800), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n14799), 
        .ZN(n14804) );
  XNOR2_X1 U16587 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n14802) );
  XNOR2_X1 U16588 ( .A(n14801), .B(n14802), .ZN(n14803) );
  XNOR2_X1 U16589 ( .A(n14804), .B(n14803), .ZN(n14805) );
  XNOR2_X1 U16590 ( .A(n14806), .B(n14805), .ZN(SUB_1596_U4) );
  XNOR2_X1 U16591 ( .A(n14807), .B(n8831), .ZN(n14808) );
  NAND2_X1 U16592 ( .A1(n14808), .A2(n10380), .ZN(n14812) );
  AOI22_X1 U16593 ( .A1(n15360), .A2(n14810), .B1(n14809), .B2(n15358), .ZN(
        n14811) );
  NAND2_X1 U16594 ( .A1(n14812), .A2(n14811), .ZN(n14832) );
  AOI21_X1 U16595 ( .B1(n15369), .B2(n14813), .A(n14832), .ZN(n14820) );
  NAND2_X1 U16596 ( .A1(n14815), .A2(n14814), .ZN(n14816) );
  NAND2_X1 U16597 ( .A1(n14817), .A2(n14816), .ZN(n14830) );
  NOR2_X1 U16598 ( .A1(n14818), .A2(n15353), .ZN(n14831) );
  AOI22_X1 U16599 ( .A1(n14830), .A2(n15323), .B1(n14831), .B2(n15336), .ZN(
        n14819) );
  OAI221_X1 U16600 ( .B1(n13255), .B2(n14820), .C1(n15372), .C2(n8819), .A(
        n14819), .ZN(P3_U3222) );
  NOR2_X1 U16601 ( .A1(n14821), .A2(n15353), .ZN(n14822) );
  AOI21_X1 U16602 ( .B1(n14823), .B2(n15405), .A(n14822), .ZN(n14824) );
  AND2_X1 U16603 ( .A1(n14825), .A2(n14824), .ZN(n14834) );
  AOI22_X1 U16604 ( .A1(n15419), .A2(n14834), .B1(n8863), .B2(n15417), .ZN(
        P3_U3472) );
  AOI21_X1 U16605 ( .B1(n14827), .B2(n15405), .A(n14826), .ZN(n14828) );
  AND2_X1 U16606 ( .A1(n14829), .A2(n14828), .ZN(n14836) );
  AOI22_X1 U16607 ( .A1(n15419), .A2(n14836), .B1(n8840), .B2(n15417), .ZN(
        P3_U3471) );
  AND2_X1 U16608 ( .A1(n14830), .A2(n15405), .ZN(n14833) );
  NOR3_X1 U16609 ( .A1(n14833), .A2(n14832), .A3(n14831), .ZN(n14838) );
  AOI22_X1 U16610 ( .A1(n15419), .A2(n14838), .B1(n8816), .B2(n15417), .ZN(
        P3_U3470) );
  INV_X1 U16611 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14835) );
  AOI22_X1 U16612 ( .A1(n15409), .A2(n14835), .B1(n14834), .B2(n15407), .ZN(
        P3_U3429) );
  INV_X1 U16613 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14837) );
  AOI22_X1 U16614 ( .A1(n15409), .A2(n14837), .B1(n14836), .B2(n15407), .ZN(
        P3_U3426) );
  INV_X1 U16615 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14839) );
  AOI22_X1 U16616 ( .A1(n15409), .A2(n14839), .B1(n14838), .B2(n15407), .ZN(
        P3_U3423) );
  NAND2_X1 U16617 ( .A1(n14841), .A2(n14840), .ZN(n14842) );
  NAND2_X1 U16618 ( .A1(n14843), .A2(n14842), .ZN(n14844) );
  AOI222_X1 U16619 ( .A1(n14848), .A2(n14847), .B1(n14846), .B2(n14845), .C1(
        n14844), .C2(n15120), .ZN(n14849) );
  NAND2_X1 U16620 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n15158)
         );
  OAI211_X1 U16621 ( .C1(n15124), .C2(n14850), .A(n14849), .B(n15158), .ZN(
        P2_U3187) );
  INV_X1 U16622 ( .A(n15255), .ZN(n15268) );
  INV_X1 U16623 ( .A(n14851), .ZN(n14855) );
  OAI21_X1 U16624 ( .B1(n15118), .B2(n15263), .A(n14852), .ZN(n14854) );
  AOI211_X1 U16625 ( .C1(n15268), .C2(n14855), .A(n14854), .B(n14853), .ZN(
        n14857) );
  AOI22_X1 U16626 ( .A1(n15279), .A2(n14857), .B1(n13564), .B2(n15277), .ZN(
        P2_U3511) );
  INV_X1 U16627 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14856) );
  AOI22_X1 U16628 ( .A1(n15270), .A2(n14857), .B1(n14856), .B2(n9800), .ZN(
        P2_U3466) );
  AOI21_X1 U16629 ( .B1(n14860), .B2(n14859), .A(n14858), .ZN(n14865) );
  OAI222_X1 U16630 ( .A1(n14935), .A2(n14865), .B1(n14864), .B2(n14863), .C1(
        n14862), .C2(n14861), .ZN(n14866) );
  INV_X1 U16631 ( .A(n14866), .ZN(n14868) );
  OAI211_X1 U16632 ( .C1(n14965), .C2(n14869), .A(n14868), .B(n14867), .ZN(
        P1_U3215) );
  NAND2_X1 U16633 ( .A1(n14870), .A2(n14951), .ZN(n15088) );
  INV_X1 U16634 ( .A(n15088), .ZN(n14872) );
  AOI21_X1 U16635 ( .B1(n14872), .B2(n14953), .A(n14871), .ZN(n14881) );
  NOR2_X1 U16636 ( .A1(n14874), .A2(n7848), .ZN(n14875) );
  XNOR2_X1 U16637 ( .A(n14876), .B(n14875), .ZN(n14879) );
  NAND2_X1 U16638 ( .A1(n14878), .A2(n14877), .ZN(n15087) );
  AOI22_X1 U16639 ( .A1(n14879), .A2(n14961), .B1(n14960), .B2(n15087), .ZN(
        n14880) );
  OAI211_X1 U16640 ( .C1(n14882), .C2(n14965), .A(n14881), .B(n14880), .ZN(
        P1_U3217) );
  XNOR2_X1 U16641 ( .A(n14883), .B(n14891), .ZN(n14885) );
  AOI21_X1 U16642 ( .B1(n14885), .B2(n15052), .A(n14884), .ZN(n14904) );
  INV_X1 U16643 ( .A(n14886), .ZN(n14887) );
  AOI222_X1 U16644 ( .A1(n14892), .A2(n14889), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n6550), .C1(n14888), .C2(n14887), .ZN(n14900) );
  XOR2_X1 U16645 ( .A(n14891), .B(n14890), .Z(n14907) );
  INV_X1 U16646 ( .A(n14892), .ZN(n14903) );
  INV_X1 U16647 ( .A(n14893), .ZN(n14896) );
  INV_X1 U16648 ( .A(n14894), .ZN(n14895) );
  OAI211_X1 U16649 ( .C1(n14903), .C2(n14896), .A(n14895), .B(n11131), .ZN(
        n14901) );
  INV_X1 U16650 ( .A(n14901), .ZN(n14897) );
  AOI22_X1 U16651 ( .A1(n14907), .A2(n14898), .B1(n15017), .B2(n14897), .ZN(
        n14899) );
  OAI211_X1 U16652 ( .C1(n6550), .C2(n14904), .A(n14900), .B(n14899), .ZN(
        P1_U3282) );
  OAI21_X1 U16653 ( .B1(n14903), .B2(n14902), .A(n14901), .ZN(n14906) );
  INV_X1 U16654 ( .A(n14904), .ZN(n14905) );
  AOI211_X1 U16655 ( .C1(n14907), .C2(n15093), .A(n14906), .B(n14905), .ZN(
        n14910) );
  AOI22_X1 U16656 ( .A1(n15107), .A2(n14910), .B1(n14908), .B2(n15105), .ZN(
        P1_U3539) );
  INV_X1 U16657 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14909) );
  AOI22_X1 U16658 ( .A1(n15096), .A2(n14910), .B1(n14909), .B2(n7451), .ZN(
        P1_U3492) );
  AOI21_X1 U16659 ( .B1(n6581), .B2(n14912), .A(n14911), .ZN(n14913) );
  XOR2_X1 U16660 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n14913), .Z(SUB_1596_U69)
         );
  AOI21_X1 U16661 ( .B1(n14916), .B2(n14915), .A(n14914), .ZN(n14917) );
  XNOR2_X1 U16662 ( .A(n7653), .B(n14917), .ZN(SUB_1596_U68) );
  OAI21_X1 U16663 ( .B1(n14920), .B2(n14919), .A(n14918), .ZN(SUB_1596_U67) );
  OAI21_X1 U16664 ( .B1(n14923), .B2(n14922), .A(n14921), .ZN(n14924) );
  XNOR2_X1 U16665 ( .A(n14924), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI222_X1 U16666 ( .A1(n15165), .A2(n14928), .B1(n15165), .B2(n14927), .C1(
        n14926), .C2(n14925), .ZN(SUB_1596_U65) );
  OAI21_X1 U16667 ( .B1(n14931), .B2(n14930), .A(n14929), .ZN(n14932) );
  XNOR2_X1 U16668 ( .A(n14932), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  AND2_X1 U16669 ( .A1(n14951), .A2(n14933), .ZN(n15027) );
  AOI21_X1 U16670 ( .B1(n14953), .B2(n15027), .A(n14934), .ZN(n14942) );
  AOI21_X1 U16671 ( .B1(n14937), .B2(n14936), .A(n14935), .ZN(n14940) );
  AOI22_X1 U16672 ( .A1(n14940), .A2(n14939), .B1(n14960), .B2(n14938), .ZN(
        n14941) );
  OAI211_X1 U16673 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n14965), .A(n14942), .B(
        n14941), .ZN(P1_U3218) );
  AND2_X1 U16674 ( .A1(n14943), .A2(n14951), .ZN(n15070) );
  AOI22_X1 U16675 ( .A1(n15070), .A2(n14953), .B1(P1_REG3_REG_8__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14949) );
  OAI21_X1 U16676 ( .B1(n14946), .B2(n14945), .A(n14944), .ZN(n14947) );
  AOI22_X1 U16677 ( .A1(n14947), .A2(n14961), .B1(n14960), .B2(n15069), .ZN(
        n14948) );
  OAI211_X1 U16678 ( .C1(n14950), .C2(n14965), .A(n14949), .B(n14948), .ZN(
        P1_U3221) );
  AND2_X1 U16679 ( .A1(n14952), .A2(n14951), .ZN(n15077) );
  AOI22_X1 U16680 ( .A1(n15077), .A2(n14953), .B1(P1_REG3_REG_9__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14964) );
  INV_X1 U16681 ( .A(n14954), .ZN(n14956) );
  NAND2_X1 U16682 ( .A1(n14956), .A2(n14955), .ZN(n14958) );
  XNOR2_X1 U16683 ( .A(n14958), .B(n14957), .ZN(n14962) );
  AOI22_X1 U16684 ( .A1(n14962), .A2(n14961), .B1(n14960), .B2(n14959), .ZN(
        n14963) );
  OAI211_X1 U16685 ( .C1(n14966), .C2(n14965), .A(n14964), .B(n14963), .ZN(
        P1_U3231) );
  AOI21_X1 U16686 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n14968), .A(n14967), 
        .ZN(n14973) );
  AOI21_X1 U16687 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14970), .A(n14969), 
        .ZN(n14971) );
  OAI222_X1 U16688 ( .A1(n14976), .A2(n14975), .B1(n14974), .B2(n14973), .C1(
        n14972), .C2(n14971), .ZN(n14977) );
  INV_X1 U16689 ( .A(n14977), .ZN(n14979) );
  OAI211_X1 U16690 ( .C1(n14981), .C2(n14980), .A(n14979), .B(n14978), .ZN(
        P1_U3258) );
  XNOR2_X1 U16691 ( .A(n14983), .B(n14982), .ZN(n15066) );
  OAI21_X1 U16692 ( .B1(n14986), .B2(n14985), .A(n14984), .ZN(n14987) );
  AND2_X1 U16693 ( .A1(n14987), .A2(n15052), .ZN(n15064) );
  AOI211_X1 U16694 ( .C1(n15059), .C2(n15066), .A(n15060), .B(n15064), .ZN(
        n14998) );
  NOR2_X1 U16695 ( .A1(n15005), .A2(n14988), .ZN(n14989) );
  AOI21_X1 U16696 ( .B1(n6550), .B2(P1_REG2_REG_7__SCAN_IN), .A(n14989), .ZN(
        n14990) );
  OAI21_X1 U16697 ( .B1(n15009), .B2(n14993), .A(n14990), .ZN(n14991) );
  INV_X1 U16698 ( .A(n14991), .ZN(n14997) );
  OAI211_X1 U16699 ( .C1(n14994), .C2(n14993), .A(n14992), .B(n11131), .ZN(
        n15063) );
  INV_X1 U16700 ( .A(n15063), .ZN(n14995) );
  AOI22_X1 U16701 ( .A1(n15066), .A2(n15018), .B1(n15017), .B2(n14995), .ZN(
        n14996) );
  OAI211_X1 U16702 ( .C1(n6550), .C2(n14998), .A(n14997), .B(n14996), .ZN(
        P1_U3286) );
  XNOR2_X1 U16703 ( .A(n14999), .B(n15001), .ZN(n15045) );
  XOR2_X1 U16704 ( .A(n15001), .B(n15000), .Z(n15003) );
  NOR2_X1 U16705 ( .A1(n15003), .A2(n15002), .ZN(n15043) );
  AOI211_X1 U16706 ( .C1(n15059), .C2(n15045), .A(n15040), .B(n15043), .ZN(
        n15021) );
  NOR2_X1 U16707 ( .A1(n15005), .A2(n15004), .ZN(n15006) );
  AOI21_X1 U16708 ( .B1(n6550), .B2(P1_REG2_REG_5__SCAN_IN), .A(n15006), .ZN(
        n15007) );
  OAI21_X1 U16709 ( .B1(n15009), .B2(n15008), .A(n15007), .ZN(n15010) );
  INV_X1 U16710 ( .A(n15010), .ZN(n15020) );
  INV_X1 U16711 ( .A(n15011), .ZN(n15015) );
  INV_X1 U16712 ( .A(n15012), .ZN(n15013) );
  AOI211_X1 U16713 ( .C1(n15016), .C2(n15015), .A(n15014), .B(n15013), .ZN(
        n15041) );
  AOI22_X1 U16714 ( .A1(n15045), .A2(n15018), .B1(n15017), .B2(n15041), .ZN(
        n15019) );
  OAI211_X1 U16715 ( .C1(n6550), .C2(n15021), .A(n15020), .B(n15019), .ZN(
        P1_U3288) );
  INV_X1 U16716 ( .A(n15022), .ZN(n15023) );
  INV_X1 U16717 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15538) );
  NOR2_X1 U16718 ( .A1(n15023), .A2(n15538), .ZN(P1_U3294) );
  AND2_X1 U16719 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15022), .ZN(P1_U3295) );
  AND2_X1 U16720 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15022), .ZN(P1_U3296) );
  AND2_X1 U16721 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15022), .ZN(P1_U3297) );
  AND2_X1 U16722 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15022), .ZN(P1_U3298) );
  AND2_X1 U16723 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15022), .ZN(P1_U3299) );
  AND2_X1 U16724 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15022), .ZN(P1_U3300) );
  AND2_X1 U16725 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15022), .ZN(P1_U3301) );
  AND2_X1 U16726 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15022), .ZN(P1_U3302) );
  AND2_X1 U16727 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15022), .ZN(P1_U3303) );
  AND2_X1 U16728 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15022), .ZN(P1_U3304) );
  AND2_X1 U16729 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15022), .ZN(P1_U3305) );
  AND2_X1 U16730 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15022), .ZN(P1_U3306) );
  AND2_X1 U16731 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15022), .ZN(P1_U3307) );
  AND2_X1 U16732 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15022), .ZN(P1_U3308) );
  INV_X1 U16733 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n15469) );
  NOR2_X1 U16734 ( .A1(n15023), .A2(n15469), .ZN(P1_U3309) );
  AND2_X1 U16735 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15022), .ZN(P1_U3310) );
  INV_X1 U16736 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n15581) );
  NOR2_X1 U16737 ( .A1(n15023), .A2(n15581), .ZN(P1_U3311) );
  AND2_X1 U16738 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15022), .ZN(P1_U3312) );
  AND2_X1 U16739 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15022), .ZN(P1_U3313) );
  AND2_X1 U16740 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15022), .ZN(P1_U3314) );
  AND2_X1 U16741 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15022), .ZN(P1_U3315) );
  AND2_X1 U16742 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15022), .ZN(P1_U3316) );
  AND2_X1 U16743 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15022), .ZN(P1_U3317) );
  AND2_X1 U16744 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15022), .ZN(P1_U3318) );
  AND2_X1 U16745 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15022), .ZN(P1_U3319) );
  AND2_X1 U16746 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15022), .ZN(P1_U3320) );
  AND2_X1 U16747 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15022), .ZN(P1_U3321) );
  AND2_X1 U16748 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15022), .ZN(P1_U3322) );
  INV_X1 U16749 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n15497) );
  NOR2_X1 U16750 ( .A1(n15023), .A2(n15497), .ZN(P1_U3323) );
  INV_X1 U16751 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15024) );
  AOI22_X1 U16752 ( .A1(n15096), .A2(n15025), .B1(n15024), .B2(n7451), .ZN(
        P1_U3459) );
  NOR2_X1 U16753 ( .A1(n15026), .A2(n15055), .ZN(n15030) );
  NOR4_X1 U16754 ( .A1(n15030), .A2(n15029), .A3(n15028), .A4(n15027), .ZN(
        n15097) );
  INV_X1 U16755 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n15031) );
  AOI22_X1 U16756 ( .A1(n15096), .A2(n15097), .B1(n15031), .B2(n7451), .ZN(
        P1_U3468) );
  INV_X1 U16757 ( .A(n15032), .ZN(n15039) );
  INV_X1 U16758 ( .A(n15033), .ZN(n15037) );
  NAND4_X1 U16759 ( .A1(n15037), .A2(n15036), .A3(n15035), .A4(n15034), .ZN(
        n15038) );
  AOI21_X1 U16760 ( .B1(n15039), .B2(n15093), .A(n15038), .ZN(n15098) );
  INV_X1 U16761 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n15580) );
  AOI22_X1 U16762 ( .A1(n15096), .A2(n15098), .B1(n15580), .B2(n7451), .ZN(
        P1_U3471) );
  OR4_X1 U16763 ( .A1(n15043), .A2(n15042), .A3(n15041), .A4(n15040), .ZN(
        n15044) );
  AOI21_X1 U16764 ( .B1(n15045), .B2(n15093), .A(n15044), .ZN(n15099) );
  INV_X1 U16765 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15046) );
  AOI22_X1 U16766 ( .A1(n15096), .A2(n15099), .B1(n15046), .B2(n7451), .ZN(
        P1_U3474) );
  INV_X1 U16767 ( .A(n15056), .ZN(n15058) );
  INV_X1 U16768 ( .A(n15047), .ZN(n15049) );
  NAND3_X1 U16769 ( .A1(n15050), .A2(n15049), .A3(n15048), .ZN(n15051) );
  AOI21_X1 U16770 ( .B1(n15053), .B2(n15052), .A(n15051), .ZN(n15054) );
  OAI21_X1 U16771 ( .B1(n15056), .B2(n15055), .A(n15054), .ZN(n15057) );
  AOI21_X1 U16772 ( .B1(n15059), .B2(n15058), .A(n15057), .ZN(n15100) );
  INV_X1 U16773 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n15567) );
  AOI22_X1 U16774 ( .A1(n15096), .A2(n15100), .B1(n15567), .B2(n7451), .ZN(
        P1_U3477) );
  INV_X1 U16775 ( .A(n15060), .ZN(n15062) );
  NAND3_X1 U16776 ( .A1(n15063), .A2(n15062), .A3(n15061), .ZN(n15065) );
  AOI211_X1 U16777 ( .C1(n15066), .C2(n15093), .A(n15065), .B(n15064), .ZN(
        n15101) );
  INV_X1 U16778 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15067) );
  AOI22_X1 U16779 ( .A1(n15096), .A2(n15101), .B1(n15067), .B2(n7451), .ZN(
        P1_U3480) );
  INV_X1 U16780 ( .A(n15068), .ZN(n15074) );
  OR4_X1 U16781 ( .A1(n15072), .A2(n15071), .A3(n15070), .A4(n15069), .ZN(
        n15073) );
  AOI21_X1 U16782 ( .B1(n15093), .B2(n15074), .A(n15073), .ZN(n15103) );
  INV_X1 U16783 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15075) );
  AOI22_X1 U16784 ( .A1(n15096), .A2(n15103), .B1(n15075), .B2(n7451), .ZN(
        P1_U3483) );
  INV_X1 U16785 ( .A(n15080), .ZN(n15083) );
  AOI211_X1 U16786 ( .C1(n15078), .C2(n11131), .A(n15077), .B(n15076), .ZN(
        n15079) );
  OAI21_X1 U16787 ( .B1(n15081), .B2(n15080), .A(n15079), .ZN(n15082) );
  AOI21_X1 U16788 ( .B1(n15084), .B2(n15083), .A(n15082), .ZN(n15104) );
  INV_X1 U16789 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15085) );
  AOI22_X1 U16790 ( .A1(n15096), .A2(n15104), .B1(n15085), .B2(n7451), .ZN(
        P1_U3486) );
  INV_X1 U16791 ( .A(n15086), .ZN(n15094) );
  INV_X1 U16792 ( .A(n15087), .ZN(n15090) );
  NAND4_X1 U16793 ( .A1(n15091), .A2(n15090), .A3(n15089), .A4(n15088), .ZN(
        n15092) );
  AOI21_X1 U16794 ( .B1(n15094), .B2(n15093), .A(n15092), .ZN(n15106) );
  INV_X1 U16795 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n15095) );
  AOI22_X1 U16796 ( .A1(n15096), .A2(n15106), .B1(n15095), .B2(n7451), .ZN(
        P1_U3489) );
  AOI22_X1 U16797 ( .A1(n15107), .A2(n15097), .B1(n10634), .B2(n15105), .ZN(
        P1_U3531) );
  AOI22_X1 U16798 ( .A1(n15107), .A2(n15098), .B1(n10637), .B2(n15105), .ZN(
        P1_U3532) );
  AOI22_X1 U16799 ( .A1(n15107), .A2(n15099), .B1(n10629), .B2(n15105), .ZN(
        P1_U3533) );
  AOI22_X1 U16800 ( .A1(n15107), .A2(n15100), .B1(n10801), .B2(n15105), .ZN(
        P1_U3534) );
  AOI22_X1 U16801 ( .A1(n15107), .A2(n15101), .B1(n10802), .B2(n15105), .ZN(
        P1_U3535) );
  AOI22_X1 U16802 ( .A1(n15107), .A2(n15103), .B1(n15102), .B2(n15105), .ZN(
        P1_U3536) );
  AOI22_X1 U16803 ( .A1(n15107), .A2(n15104), .B1(n9993), .B2(n15105), .ZN(
        P1_U3537) );
  AOI22_X1 U16804 ( .A1(n15107), .A2(n15106), .B1(n15536), .B2(n15105), .ZN(
        P1_U3538) );
  NOR2_X1 U16805 ( .A1(n15196), .A2(P2_U3947), .ZN(P2_U3087) );
  NAND2_X1 U16806 ( .A1(n15109), .A2(n15108), .ZN(n15110) );
  XNOR2_X1 U16807 ( .A(n15111), .B(n15110), .ZN(n15121) );
  AOI22_X1 U16808 ( .A1(n15115), .A2(n15114), .B1(n15113), .B2(n15112), .ZN(
        n15116) );
  OAI21_X1 U16809 ( .B1(n15118), .B2(n15117), .A(n15116), .ZN(n15119) );
  AOI21_X1 U16810 ( .B1(n15121), .B2(n15120), .A(n15119), .ZN(n15122) );
  NAND2_X1 U16811 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n15140)
         );
  OAI211_X1 U16812 ( .C1(n15124), .C2(n15123), .A(n15122), .B(n15140), .ZN(
        P2_U3196) );
  INV_X1 U16813 ( .A(n15125), .ZN(n15131) );
  NAND3_X1 U16814 ( .A1(n15128), .A2(n15127), .A3(n15126), .ZN(n15130) );
  AOI21_X1 U16815 ( .B1(n15131), .B2(n15130), .A(n15129), .ZN(n15139) );
  AOI21_X1 U16816 ( .B1(n15134), .B2(n15133), .A(n15132), .ZN(n15137) );
  OAI22_X1 U16817 ( .A1(n15137), .A2(n15136), .B1(n15135), .B2(n15204), .ZN(
        n15138) );
  NOR2_X1 U16818 ( .A1(n15139), .A2(n15138), .ZN(n15141) );
  OAI211_X1 U16819 ( .C1(n7653), .C2(n15166), .A(n15141), .B(n15140), .ZN(
        P2_U3226) );
  AOI22_X1 U16820 ( .A1(n15196), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3088), .ZN(n15153) );
  OAI211_X1 U16821 ( .C1(n15144), .C2(n15143), .A(n15142), .B(n15190), .ZN(
        n15152) );
  OAI211_X1 U16822 ( .C1(n15147), .C2(n15146), .A(n15145), .B(n15198), .ZN(
        n15151) );
  INV_X1 U16823 ( .A(n15148), .ZN(n15149) );
  NAND2_X1 U16824 ( .A1(n15168), .A2(n15149), .ZN(n15150) );
  NAND4_X1 U16825 ( .A1(n15153), .A2(n15152), .A3(n15151), .A4(n15150), .ZN(
        P2_U3227) );
  OAI211_X1 U16826 ( .C1(n15156), .C2(n15155), .A(n15190), .B(n15154), .ZN(
        n15157) );
  NAND2_X1 U16827 ( .A1(n15158), .A2(n15157), .ZN(n15159) );
  AOI21_X1 U16828 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(n15196), .A(n15159), 
        .ZN(n15163) );
  OAI211_X1 U16829 ( .C1(P2_REG2_REG_14__SCAN_IN), .C2(n15161), .A(n15198), 
        .B(n15160), .ZN(n15162) );
  OAI211_X1 U16830 ( .C1(n15204), .C2(n15164), .A(n15163), .B(n15162), .ZN(
        P2_U3228) );
  OAI22_X1 U16831 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8375), .B1(n15166), .B2(
        n15165), .ZN(n15167) );
  AOI21_X1 U16832 ( .B1(n15169), .B2(n15168), .A(n15167), .ZN(n15176) );
  OAI211_X1 U16833 ( .C1(n15171), .C2(P2_REG2_REG_15__SCAN_IN), .A(n15198), 
        .B(n15170), .ZN(n15175) );
  OAI211_X1 U16834 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n15173), .A(n15190), 
        .B(n15172), .ZN(n15174) );
  NAND3_X1 U16835 ( .A1(n15176), .A2(n15175), .A3(n15174), .ZN(P2_U3229) );
  OAI211_X1 U16836 ( .C1(n15179), .C2(n15178), .A(n15190), .B(n15177), .ZN(
        n15180) );
  NAND2_X1 U16837 ( .A1(n15181), .A2(n15180), .ZN(n15182) );
  AOI21_X1 U16838 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(n15196), .A(n15182), 
        .ZN(n15187) );
  OAI211_X1 U16839 ( .C1(n15185), .C2(n15184), .A(n15198), .B(n15183), .ZN(
        n15186) );
  OAI211_X1 U16840 ( .C1(n15204), .C2(n15188), .A(n15187), .B(n15186), .ZN(
        P2_U3230) );
  OAI211_X1 U16841 ( .C1(n15192), .C2(n15191), .A(n15190), .B(n15189), .ZN(
        n15193) );
  NAND2_X1 U16842 ( .A1(n15194), .A2(n15193), .ZN(n15195) );
  AOI21_X1 U16843 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(n15196), .A(n15195), 
        .ZN(n15202) );
  OAI211_X1 U16844 ( .C1(n15200), .C2(n15199), .A(n15198), .B(n15197), .ZN(
        n15201) );
  OAI211_X1 U16845 ( .C1(n15204), .C2(n15203), .A(n15202), .B(n15201), .ZN(
        P2_U3231) );
  INV_X1 U16846 ( .A(n15210), .ZN(n15212) );
  AND2_X1 U16847 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15206), .ZN(P2_U3266) );
  AND2_X1 U16848 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15206), .ZN(P2_U3267) );
  AND2_X1 U16849 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15206), .ZN(P2_U3268) );
  AND2_X1 U16850 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15206), .ZN(P2_U3269) );
  AND2_X1 U16851 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15206), .ZN(P2_U3270) );
  AND2_X1 U16852 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15206), .ZN(P2_U3271) );
  AND2_X1 U16853 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15206), .ZN(P2_U3272) );
  AND2_X1 U16854 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15206), .ZN(P2_U3273) );
  AND2_X1 U16855 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15206), .ZN(P2_U3274) );
  AND2_X1 U16856 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15206), .ZN(P2_U3275) );
  AND2_X1 U16857 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15206), .ZN(P2_U3276) );
  AND2_X1 U16858 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15206), .ZN(P2_U3277) );
  INV_X1 U16859 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n15504) );
  NOR2_X1 U16860 ( .A1(n15207), .A2(n15504), .ZN(P2_U3278) );
  AND2_X1 U16861 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15206), .ZN(P2_U3279) );
  INV_X1 U16862 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n15557) );
  NOR2_X1 U16863 ( .A1(n15207), .A2(n15557), .ZN(P2_U3280) );
  INV_X1 U16864 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15616) );
  NOR2_X1 U16865 ( .A1(n15207), .A2(n15616), .ZN(P2_U3281) );
  AND2_X1 U16866 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15206), .ZN(P2_U3282) );
  AND2_X1 U16867 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15206), .ZN(P2_U3283) );
  INV_X1 U16868 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n15570) );
  NOR2_X1 U16869 ( .A1(n15207), .A2(n15570), .ZN(P2_U3284) );
  AND2_X1 U16870 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15206), .ZN(P2_U3285) );
  AND2_X1 U16871 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15206), .ZN(P2_U3286) );
  AND2_X1 U16872 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15206), .ZN(P2_U3287) );
  AND2_X1 U16873 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15206), .ZN(P2_U3288) );
  AND2_X1 U16874 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15206), .ZN(P2_U3289) );
  AND2_X1 U16875 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15206), .ZN(P2_U3290) );
  AND2_X1 U16876 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15206), .ZN(P2_U3291) );
  INV_X1 U16877 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n15442) );
  NOR2_X1 U16878 ( .A1(n15207), .A2(n15442), .ZN(P2_U3292) );
  AND2_X1 U16879 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15206), .ZN(P2_U3293) );
  INV_X1 U16880 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n15614) );
  NOR2_X1 U16881 ( .A1(n15207), .A2(n15614), .ZN(P2_U3294) );
  INV_X1 U16882 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n15501) );
  NOR2_X1 U16883 ( .A1(n15207), .A2(n15501), .ZN(P2_U3295) );
  AOI22_X1 U16884 ( .A1(n15210), .A2(n15209), .B1(n15208), .B2(n15212), .ZN(
        P2_U3416) );
  AOI21_X1 U16885 ( .B1(n15489), .B2(n15212), .A(n15211), .ZN(P2_U3417) );
  INV_X1 U16886 ( .A(n15213), .ZN(n15216) );
  INV_X1 U16887 ( .A(n15214), .ZN(n15215) );
  AOI211_X1 U16888 ( .C1(n15268), .C2(n15217), .A(n15216), .B(n15215), .ZN(
        n15271) );
  AOI22_X1 U16889 ( .A1(n15270), .A2(n15271), .B1(n8098), .B2(n9800), .ZN(
        P2_U3430) );
  INV_X1 U16890 ( .A(n15218), .ZN(n15219) );
  AOI21_X1 U16891 ( .B1(n15256), .B2(n15255), .A(n15219), .ZN(n15224) );
  OAI211_X1 U16892 ( .C1(n15222), .C2(n15263), .A(n15221), .B(n15220), .ZN(
        n15223) );
  NOR2_X1 U16893 ( .A1(n15224), .A2(n15223), .ZN(n15272) );
  AOI22_X1 U16894 ( .A1(n15270), .A2(n15272), .B1(n7608), .B2(n9800), .ZN(
        P2_U3433) );
  INV_X1 U16895 ( .A(n15225), .ZN(n15226) );
  AOI22_X1 U16896 ( .A1(n15270), .A2(n15226), .B1(n8135), .B2(n9800), .ZN(
        P2_U3436) );
  AND2_X1 U16897 ( .A1(n15227), .A2(n15251), .ZN(n15228) );
  NOR2_X1 U16898 ( .A1(n15229), .A2(n15228), .ZN(n15233) );
  OR2_X1 U16899 ( .A1(n15230), .A2(n15255), .ZN(n15232) );
  OR2_X1 U16900 ( .A1(n15230), .A2(n15256), .ZN(n15231) );
  INV_X1 U16901 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15235) );
  AOI22_X1 U16902 ( .A1(n15270), .A2(n15273), .B1(n15235), .B2(n9800), .ZN(
        P2_U3442) );
  INV_X1 U16903 ( .A(n15236), .ZN(n15242) );
  INV_X1 U16904 ( .A(n15237), .ZN(n15238) );
  OAI21_X1 U16905 ( .B1(n15239), .B2(n15263), .A(n15238), .ZN(n15241) );
  AOI211_X1 U16906 ( .C1(n15268), .C2(n15242), .A(n15241), .B(n15240), .ZN(
        n15274) );
  INV_X1 U16907 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15243) );
  AOI22_X1 U16908 ( .A1(n15270), .A2(n15274), .B1(n15243), .B2(n9800), .ZN(
        P2_U3445) );
  AOI21_X1 U16909 ( .B1(n15251), .B2(n15245), .A(n15244), .ZN(n15246) );
  OAI211_X1 U16910 ( .C1(n15249), .C2(n15248), .A(n15247), .B(n15246), .ZN(
        n15250) );
  INV_X1 U16911 ( .A(n15250), .ZN(n15275) );
  AOI22_X1 U16912 ( .A1(n15270), .A2(n15275), .B1(n8223), .B2(n9800), .ZN(
        P2_U3451) );
  NAND2_X1 U16913 ( .A1(n15252), .A2(n15251), .ZN(n15253) );
  OAI211_X1 U16914 ( .C1(n15257), .C2(n15255), .A(n15254), .B(n15253), .ZN(
        n15260) );
  NOR2_X1 U16915 ( .A1(n15257), .A2(n15256), .ZN(n15258) );
  NOR3_X1 U16916 ( .A1(n15260), .A2(n15259), .A3(n15258), .ZN(n15276) );
  INV_X1 U16917 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n15261) );
  AOI22_X1 U16918 ( .A1(n15270), .A2(n15276), .B1(n15261), .B2(n9800), .ZN(
        P2_U3457) );
  OAI21_X1 U16919 ( .B1(n15264), .B2(n15263), .A(n15262), .ZN(n15266) );
  AOI211_X1 U16920 ( .C1(n15268), .C2(n15267), .A(n15266), .B(n15265), .ZN(
        n15278) );
  INV_X1 U16921 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15269) );
  AOI22_X1 U16922 ( .A1(n15270), .A2(n15278), .B1(n15269), .B2(n9800), .ZN(
        P2_U3460) );
  AOI22_X1 U16923 ( .A1(n15279), .A2(n15271), .B1(n10620), .B2(n15277), .ZN(
        P2_U3499) );
  AOI22_X1 U16924 ( .A1(n15279), .A2(n15272), .B1(n8117), .B2(n15277), .ZN(
        P2_U3500) );
  AOI22_X1 U16925 ( .A1(n15279), .A2(n15273), .B1(n10577), .B2(n15277), .ZN(
        P2_U3503) );
  AOI22_X1 U16926 ( .A1(n15279), .A2(n15274), .B1(n10579), .B2(n15277), .ZN(
        P2_U3504) );
  AOI22_X1 U16927 ( .A1(n15279), .A2(n15275), .B1(n10586), .B2(n15277), .ZN(
        P2_U3506) );
  AOI22_X1 U16928 ( .A1(n15279), .A2(n15276), .B1(n10673), .B2(n15277), .ZN(
        P2_U3508) );
  AOI22_X1 U16929 ( .A1(n15279), .A2(n15278), .B1(n8277), .B2(n15277), .ZN(
        P2_U3509) );
  NOR2_X1 U16930 ( .A1(P3_U3897), .A2(n15280), .ZN(P3_U3150) );
  XOR2_X1 U16931 ( .A(n15281), .B(n15283), .Z(n15406) );
  NAND2_X1 U16932 ( .A1(n15406), .A2(n15323), .ZN(n15293) );
  INV_X1 U16933 ( .A(n15311), .ZN(n15286) );
  XNOR2_X1 U16934 ( .A(n15284), .B(n15283), .ZN(n15285) );
  OAI222_X1 U16935 ( .A1(n15300), .A2(n7100), .B1(n15298), .B2(n15286), .C1(
        n15285), .C2(n15366), .ZN(n15403) );
  INV_X1 U16936 ( .A(n15336), .ZN(n15290) );
  NOR2_X1 U16937 ( .A1(n15287), .A2(n15353), .ZN(n15404) );
  INV_X1 U16938 ( .A(n15404), .ZN(n15289) );
  OAI22_X1 U16939 ( .A1(n15290), .A2(n15289), .B1(n15288), .B2(n15326), .ZN(
        n15291) );
  AOI221_X1 U16940 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n13255), .C1(n15403), 
        .C2(n15372), .A(n15291), .ZN(n15292) );
  NAND2_X1 U16941 ( .A1(n15293), .A2(n15292), .ZN(P3_U3223) );
  INV_X1 U16942 ( .A(n15330), .ZN(n15297) );
  XNOR2_X1 U16943 ( .A(n15294), .B(n15295), .ZN(n15296) );
  OAI222_X1 U16944 ( .A1(n15300), .A2(n15299), .B1(n15298), .B2(n15297), .C1(
        n15296), .C2(n15366), .ZN(n15399) );
  OAI22_X1 U16945 ( .A1(n11862), .A2(n15372), .B1(n15326), .B2(n15301), .ZN(
        n15307) );
  XNOR2_X1 U16946 ( .A(n15303), .B(n15302), .ZN(n15401) );
  NOR2_X1 U16947 ( .A1(n15304), .A2(n15353), .ZN(n15400) );
  AOI22_X1 U16948 ( .A1(n15401), .A2(n15323), .B1(n15400), .B2(n15336), .ZN(
        n15305) );
  INV_X1 U16949 ( .A(n15305), .ZN(n15306) );
  AOI211_X1 U16950 ( .C1(n15372), .C2(n15399), .A(n15307), .B(n15306), .ZN(
        n15308) );
  INV_X1 U16951 ( .A(n15308), .ZN(P3_U3224) );
  XNOR2_X1 U16952 ( .A(n15309), .B(n15315), .ZN(n15312) );
  AOI222_X1 U16953 ( .A1(n10380), .A2(n15312), .B1(n15311), .B2(n15358), .C1(
        n15310), .C2(n15360), .ZN(n15395) );
  AOI22_X1 U16954 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n13255), .B1(n15369), 
        .B2(n15313), .ZN(n15319) );
  OAI21_X1 U16955 ( .B1(n15316), .B2(n15315), .A(n15314), .ZN(n15398) );
  NOR2_X1 U16956 ( .A1(n15317), .A2(n15353), .ZN(n15397) );
  AOI22_X1 U16957 ( .A1(n15398), .A2(n15323), .B1(n15397), .B2(n15336), .ZN(
        n15318) );
  OAI211_X1 U16958 ( .C1(n13255), .C2(n15395), .A(n15319), .B(n15318), .ZN(
        P3_U3225) );
  OAI21_X1 U16959 ( .B1(n15322), .B2(n15321), .A(n15320), .ZN(n15393) );
  NAND2_X1 U16960 ( .A1(n15393), .A2(n15323), .ZN(n15338) );
  NOR2_X1 U16961 ( .A1(n15324), .A2(n15353), .ZN(n15392) );
  NOR2_X1 U16962 ( .A1(n15326), .A2(n15325), .ZN(n15335) );
  OAI211_X1 U16963 ( .C1(n15329), .C2(n15328), .A(n15327), .B(n10380), .ZN(
        n15333) );
  AOI22_X1 U16964 ( .A1(n15360), .A2(n15331), .B1(n15330), .B2(n15358), .ZN(
        n15332) );
  NAND2_X1 U16965 ( .A1(n15333), .A2(n15332), .ZN(n15391) );
  MUX2_X1 U16966 ( .A(P3_REG2_REG_7__SCAN_IN), .B(n15391), .S(n15372), .Z(
        n15334) );
  AOI211_X1 U16967 ( .C1(n15336), .C2(n15392), .A(n15335), .B(n15334), .ZN(
        n15337) );
  NAND2_X1 U16968 ( .A1(n15338), .A2(n15337), .ZN(P3_U3226) );
  XNOR2_X1 U16969 ( .A(n15339), .B(n15341), .ZN(n15347) );
  OAI21_X1 U16970 ( .B1(n15342), .B2(n15341), .A(n15340), .ZN(n15380) );
  NAND2_X1 U16971 ( .A1(n15380), .A2(n15363), .ZN(n15346) );
  AOI22_X1 U16972 ( .A1(n15360), .A2(n15344), .B1(n15343), .B2(n15358), .ZN(
        n15345) );
  OAI211_X1 U16973 ( .C1(n15366), .C2(n15347), .A(n15346), .B(n15345), .ZN(
        n15378) );
  NOR2_X1 U16974 ( .A1(n15348), .A2(n15353), .ZN(n15379) );
  AOI22_X1 U16975 ( .A1(n15380), .A2(n15349), .B1(n15379), .B2(n15368), .ZN(
        n15350) );
  INV_X1 U16976 ( .A(n15350), .ZN(n15351) );
  AOI211_X1 U16977 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15369), .A(n15378), .B(
        n15351), .ZN(n15352) );
  AOI22_X1 U16978 ( .A1(n13255), .A2(n10766), .B1(n15352), .B2(n15372), .ZN(
        P3_U3231) );
  NOR2_X1 U16979 ( .A1(n15354), .A2(n15353), .ZN(n15375) );
  AOI21_X1 U16980 ( .B1(n15357), .B2(n15356), .A(n15355), .ZN(n15367) );
  AOI22_X1 U16981 ( .A1(n15360), .A2(n15359), .B1(n15423), .B2(n15358), .ZN(
        n15365) );
  NAND2_X1 U16982 ( .A1(n15362), .A2(n15361), .ZN(n15376) );
  NAND2_X1 U16983 ( .A1(n15376), .A2(n15363), .ZN(n15364) );
  OAI211_X1 U16984 ( .C1(n15367), .C2(n15366), .A(n15365), .B(n15364), .ZN(
        n15374) );
  AOI21_X1 U16985 ( .B1(n15375), .B2(n15368), .A(n15374), .ZN(n15373) );
  AOI22_X1 U16986 ( .A1(n15376), .A2(n15370), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15369), .ZN(n15371) );
  OAI221_X1 U16987 ( .B1(n13255), .B2(n15373), .C1(n15372), .C2(n10757), .A(
        n15371), .ZN(P3_U3232) );
  INV_X1 U16988 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15377) );
  AOI211_X1 U16989 ( .C1(n15381), .C2(n15376), .A(n15375), .B(n15374), .ZN(
        n15410) );
  AOI22_X1 U16990 ( .A1(n15409), .A2(n15377), .B1(n15410), .B2(n15407), .ZN(
        P3_U3393) );
  INV_X1 U16991 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15382) );
  AOI211_X1 U16992 ( .C1(n15381), .C2(n15380), .A(n15379), .B(n15378), .ZN(
        n15411) );
  AOI22_X1 U16993 ( .A1(n15409), .A2(n15382), .B1(n15411), .B2(n15407), .ZN(
        P3_U3396) );
  INV_X1 U16994 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15713) );
  INV_X1 U16995 ( .A(n15383), .ZN(n15386) );
  AOI211_X1 U16996 ( .C1(n15386), .C2(n15405), .A(n15385), .B(n15384), .ZN(
        n15412) );
  AOI22_X1 U16997 ( .A1(n15409), .A2(n15713), .B1(n15412), .B2(n15407), .ZN(
        P3_U3399) );
  INV_X1 U16998 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15390) );
  AOI211_X1 U16999 ( .C1(n15405), .C2(n15389), .A(n15388), .B(n15387), .ZN(
        n15413) );
  AOI22_X1 U17000 ( .A1(n15409), .A2(n15390), .B1(n15413), .B2(n15407), .ZN(
        P3_U3405) );
  INV_X1 U17001 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15394) );
  AOI211_X1 U17002 ( .C1(n15405), .C2(n15393), .A(n15392), .B(n15391), .ZN(
        n15414) );
  AOI22_X1 U17003 ( .A1(n15409), .A2(n15394), .B1(n15414), .B2(n15407), .ZN(
        P3_U3411) );
  INV_X1 U17004 ( .A(n15395), .ZN(n15396) );
  AOI211_X1 U17005 ( .C1(n15405), .C2(n15398), .A(n15397), .B(n15396), .ZN(
        n15415) );
  AOI22_X1 U17006 ( .A1(n15409), .A2(n8767), .B1(n15415), .B2(n15407), .ZN(
        P3_U3414) );
  INV_X1 U17007 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15402) );
  AOI211_X1 U17008 ( .C1(n15401), .C2(n15405), .A(n15400), .B(n15399), .ZN(
        n15416) );
  AOI22_X1 U17009 ( .A1(n15409), .A2(n15402), .B1(n15416), .B2(n15407), .ZN(
        P3_U3417) );
  INV_X1 U17010 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15408) );
  AOI211_X1 U17011 ( .C1(n15406), .C2(n15405), .A(n15404), .B(n15403), .ZN(
        n15418) );
  AOI22_X1 U17012 ( .A1(n15409), .A2(n15408), .B1(n15418), .B2(n15407), .ZN(
        P3_U3420) );
  AOI22_X1 U17013 ( .A1(n15419), .A2(n15410), .B1(n10756), .B2(n15417), .ZN(
        P3_U3460) );
  AOI22_X1 U17014 ( .A1(n15419), .A2(n15411), .B1(n10765), .B2(n15417), .ZN(
        P3_U3461) );
  AOI22_X1 U17015 ( .A1(n15419), .A2(n15412), .B1(n10875), .B2(n15417), .ZN(
        P3_U3462) );
  AOI22_X1 U17016 ( .A1(n15419), .A2(n15413), .B1(n10910), .B2(n15417), .ZN(
        P3_U3464) );
  AOI22_X1 U17017 ( .A1(n15419), .A2(n15414), .B1(n11217), .B2(n15417), .ZN(
        P3_U3466) );
  AOI22_X1 U17018 ( .A1(n15419), .A2(n15415), .B1(n11559), .B2(n15417), .ZN(
        P3_U3467) );
  AOI22_X1 U17019 ( .A1(n15419), .A2(n15416), .B1(n11861), .B2(n15417), .ZN(
        P3_U3468) );
  AOI22_X1 U17020 ( .A1(n15419), .A2(n15418), .B1(n8800), .B2(n15417), .ZN(
        P3_U3469) );
  NAND2_X1 U17021 ( .A1(n15421), .A2(n15420), .ZN(n15430) );
  NAND2_X1 U17022 ( .A1(n15423), .A2(n15422), .ZN(n15429) );
  NAND2_X1 U17023 ( .A1(n15425), .A2(n15424), .ZN(n15428) );
  INV_X1 U17024 ( .A(n15426), .ZN(n15427) );
  NAND4_X1 U17025 ( .A1(n15430), .A2(n15429), .A3(n15428), .A4(n15427), .ZN(
        n15438) );
  OR2_X1 U17026 ( .A1(n15432), .A2(n15431), .ZN(n15435) );
  AOI211_X1 U17027 ( .C1(n15436), .C2(n15435), .A(n15434), .B(n15433), .ZN(
        n15437) );
  AOI211_X1 U17028 ( .C1(n15440), .C2(n15439), .A(n15438), .B(n15437), .ZN(
        n15673) );
  AOI22_X1 U17029 ( .A1(n15442), .A2(keyinput127), .B1(keyinput89), .B2(n13707), .ZN(n15441) );
  OAI221_X1 U17030 ( .B1(n15442), .B2(keyinput127), .C1(n13707), .C2(
        keyinput89), .A(n15441), .ZN(n15453) );
  INV_X1 U17031 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n15444) );
  AOI22_X1 U17032 ( .A1(n15445), .A2(keyinput9), .B1(n15444), .B2(keyinput104), 
        .ZN(n15443) );
  OAI221_X1 U17033 ( .B1(n15445), .B2(keyinput9), .C1(n15444), .C2(keyinput104), .A(n15443), .ZN(n15452) );
  INV_X1 U17034 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n15716) );
  AOI22_X1 U17035 ( .A1(n15447), .A2(keyinput22), .B1(n15716), .B2(keyinput32), 
        .ZN(n15446) );
  OAI221_X1 U17036 ( .B1(n15447), .B2(keyinput22), .C1(n15716), .C2(keyinput32), .A(n15446), .ZN(n15451) );
  XNOR2_X1 U17037 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput45), .ZN(n15449) );
  XNOR2_X1 U17038 ( .A(SI_13_), .B(keyinput60), .ZN(n15448) );
  NAND2_X1 U17039 ( .A1(n15449), .A2(n15448), .ZN(n15450) );
  NOR4_X1 U17040 ( .A1(n15453), .A2(n15452), .A3(n15451), .A4(n15450), .ZN(
        n15495) );
  AOI22_X1 U17041 ( .A1(n15455), .A2(keyinput88), .B1(n10802), .B2(keyinput42), 
        .ZN(n15454) );
  OAI221_X1 U17042 ( .B1(n15455), .B2(keyinput88), .C1(n10802), .C2(keyinput42), .A(n15454), .ZN(n15467) );
  AOI22_X1 U17043 ( .A1(n15458), .A2(keyinput7), .B1(n15457), .B2(keyinput66), 
        .ZN(n15456) );
  OAI221_X1 U17044 ( .B1(n15458), .B2(keyinput7), .C1(n15457), .C2(keyinput66), 
        .A(n15456), .ZN(n15466) );
  INV_X1 U17045 ( .A(P3_B_REG_SCAN_IN), .ZN(n15460) );
  AOI22_X1 U17046 ( .A1(n15461), .A2(keyinput77), .B1(keyinput110), .B2(n15460), .ZN(n15459) );
  OAI221_X1 U17047 ( .B1(n15461), .B2(keyinput77), .C1(n15460), .C2(
        keyinput110), .A(n15459), .ZN(n15465) );
  XOR2_X1 U17048 ( .A(n11202), .B(keyinput1), .Z(n15463) );
  XNOR2_X1 U17049 ( .A(P1_REG3_REG_5__SCAN_IN), .B(keyinput5), .ZN(n15462) );
  NAND2_X1 U17050 ( .A1(n15463), .A2(n15462), .ZN(n15464) );
  NOR4_X1 U17051 ( .A1(n15467), .A2(n15466), .A3(n15465), .A4(n15464), .ZN(
        n15494) );
  AOI22_X1 U17052 ( .A1(n15469), .A2(keyinput17), .B1(keyinput122), .B2(n10631), .ZN(n15468) );
  OAI221_X1 U17053 ( .B1(n15469), .B2(keyinput17), .C1(n10631), .C2(
        keyinput122), .A(n15468), .ZN(n15478) );
  AOI22_X1 U17054 ( .A1(n11861), .A2(keyinput6), .B1(keyinput65), .B2(n13529), 
        .ZN(n15470) );
  OAI221_X1 U17055 ( .B1(n11861), .B2(keyinput6), .C1(n13529), .C2(keyinput65), 
        .A(n15470), .ZN(n15477) );
  AOI22_X1 U17056 ( .A1(n15472), .A2(keyinput36), .B1(n15710), .B2(keyinput123), .ZN(n15471) );
  OAI221_X1 U17057 ( .B1(n15472), .B2(keyinput36), .C1(n15710), .C2(
        keyinput123), .A(n15471), .ZN(n15476) );
  XNOR2_X1 U17058 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput62), .ZN(n15474)
         );
  XNOR2_X1 U17059 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput106), .ZN(n15473)
         );
  NAND2_X1 U17060 ( .A1(n15474), .A2(n15473), .ZN(n15475) );
  NOR4_X1 U17061 ( .A1(n15478), .A2(n15477), .A3(n15476), .A4(n15475), .ZN(
        n15493) );
  AOI22_X1 U17062 ( .A1(n15481), .A2(keyinput41), .B1(keyinput126), .B2(n15480), .ZN(n15479) );
  OAI221_X1 U17063 ( .B1(n15481), .B2(keyinput41), .C1(n15480), .C2(
        keyinput126), .A(n15479), .ZN(n15484) );
  XOR2_X1 U17064 ( .A(P1_REG0_REG_24__SCAN_IN), .B(keyinput26), .Z(n15483) );
  XOR2_X1 U17065 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(keyinput73), .Z(n15482) );
  NOR3_X1 U17066 ( .A1(n15484), .A2(n15483), .A3(n15482), .ZN(n15488) );
  XNOR2_X1 U17067 ( .A(P3_IR_REG_7__SCAN_IN), .B(keyinput94), .ZN(n15487) );
  XNOR2_X1 U17068 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput71), .ZN(n15486)
         );
  XNOR2_X1 U17069 ( .A(P2_REG1_REG_15__SCAN_IN), .B(keyinput18), .ZN(n15485)
         );
  NAND4_X1 U17070 ( .A1(n15488), .A2(n15487), .A3(n15486), .A4(n15485), .ZN(
        n15491) );
  XNOR2_X1 U17071 ( .A(n15489), .B(keyinput16), .ZN(n15490) );
  NOR2_X1 U17072 ( .A1(n15491), .A2(n15490), .ZN(n15492) );
  NAND4_X1 U17073 ( .A1(n15495), .A2(n15494), .A3(n15493), .A4(n15492), .ZN(
        n15671) );
  INV_X1 U17074 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n15498) );
  AOI22_X1 U17075 ( .A1(n15498), .A2(keyinput28), .B1(keyinput112), .B2(n15497), .ZN(n15496) );
  OAI221_X1 U17076 ( .B1(n15498), .B2(keyinput28), .C1(n15497), .C2(
        keyinput112), .A(n15496), .ZN(n15510) );
  AOI22_X1 U17077 ( .A1(n15501), .A2(keyinput14), .B1(keyinput81), .B2(n15500), 
        .ZN(n15499) );
  OAI221_X1 U17078 ( .B1(n15501), .B2(keyinput14), .C1(n15500), .C2(keyinput81), .A(n15499), .ZN(n15509) );
  AOI22_X1 U17079 ( .A1(n15504), .A2(keyinput38), .B1(keyinput90), .B2(n15503), 
        .ZN(n15502) );
  OAI221_X1 U17080 ( .B1(n15504), .B2(keyinput38), .C1(n15503), .C2(keyinput90), .A(n15502), .ZN(n15508) );
  XNOR2_X1 U17081 ( .A(P3_IR_REG_4__SCAN_IN), .B(keyinput61), .ZN(n15506) );
  XNOR2_X1 U17082 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput12), .ZN(n15505)
         );
  NAND2_X1 U17083 ( .A1(n15506), .A2(n15505), .ZN(n15507) );
  NOR4_X1 U17084 ( .A1(n15510), .A2(n15509), .A3(n15508), .A4(n15507), .ZN(
        n15552) );
  AOI22_X1 U17085 ( .A1(n15512), .A2(keyinput24), .B1(keyinput72), .B2(n10657), 
        .ZN(n15511) );
  OAI221_X1 U17086 ( .B1(n15512), .B2(keyinput24), .C1(n10657), .C2(keyinput72), .A(n15511), .ZN(n15522) );
  AOI22_X1 U17087 ( .A1(n15515), .A2(keyinput0), .B1(keyinput93), .B2(n15514), 
        .ZN(n15513) );
  OAI221_X1 U17088 ( .B1(n15515), .B2(keyinput0), .C1(n15514), .C2(keyinput93), 
        .A(n15513), .ZN(n15521) );
  XOR2_X1 U17089 ( .A(n10765), .B(keyinput102), .Z(n15519) );
  XNOR2_X1 U17090 ( .A(P3_IR_REG_18__SCAN_IN), .B(keyinput2), .ZN(n15518) );
  XNOR2_X1 U17091 ( .A(SI_5_), .B(keyinput82), .ZN(n15517) );
  XNOR2_X1 U17092 ( .A(P1_REG0_REG_23__SCAN_IN), .B(keyinput108), .ZN(n15516)
         );
  NAND4_X1 U17093 ( .A1(n15519), .A2(n15518), .A3(n15517), .A4(n15516), .ZN(
        n15520) );
  NOR3_X1 U17094 ( .A1(n15522), .A2(n15521), .A3(n15520), .ZN(n15551) );
  AOI22_X1 U17095 ( .A1(n8223), .A2(keyinput31), .B1(keyinput87), .B2(n15696), 
        .ZN(n15523) );
  OAI221_X1 U17096 ( .B1(n8223), .B2(keyinput31), .C1(n15696), .C2(keyinput87), 
        .A(n15523), .ZN(n15534) );
  INV_X1 U17097 ( .A(P1_WR_REG_SCAN_IN), .ZN(n15525) );
  AOI22_X1 U17098 ( .A1(n15715), .A2(keyinput78), .B1(keyinput105), .B2(n15525), .ZN(n15524) );
  OAI221_X1 U17099 ( .B1(n15715), .B2(keyinput78), .C1(n15525), .C2(
        keyinput105), .A(n15524), .ZN(n15533) );
  AOI22_X1 U17100 ( .A1(n15528), .A2(keyinput114), .B1(n15527), .B2(keyinput80), .ZN(n15526) );
  OAI221_X1 U17101 ( .B1(n15528), .B2(keyinput114), .C1(n15527), .C2(
        keyinput80), .A(n15526), .ZN(n15532) );
  XNOR2_X1 U17102 ( .A(P1_REG3_REG_2__SCAN_IN), .B(keyinput13), .ZN(n15530) );
  XNOR2_X1 U17103 ( .A(SI_9_), .B(keyinput63), .ZN(n15529) );
  NAND2_X1 U17104 ( .A1(n15530), .A2(n15529), .ZN(n15531) );
  NOR4_X1 U17105 ( .A1(n15534), .A2(n15533), .A3(n15532), .A4(n15531), .ZN(
        n15550) );
  AOI22_X1 U17106 ( .A1(n15536), .A2(keyinput95), .B1(n13721), .B2(keyinput8), 
        .ZN(n15535) );
  OAI221_X1 U17107 ( .B1(n15536), .B2(keyinput95), .C1(n13721), .C2(keyinput8), 
        .A(n15535), .ZN(n15548) );
  AOI22_X1 U17108 ( .A1(n15538), .A2(keyinput39), .B1(keyinput59), .B2(n10442), 
        .ZN(n15537) );
  OAI221_X1 U17109 ( .B1(n15538), .B2(keyinput39), .C1(n10442), .C2(keyinput59), .A(n15537), .ZN(n15547) );
  AOI22_X1 U17110 ( .A1(n15541), .A2(keyinput92), .B1(n15540), .B2(keyinput51), 
        .ZN(n15539) );
  OAI221_X1 U17111 ( .B1(n15541), .B2(keyinput92), .C1(n15540), .C2(keyinput51), .A(n15539), .ZN(n15546) );
  AOI22_X1 U17112 ( .A1(n15544), .A2(keyinput44), .B1(keyinput40), .B2(n15543), 
        .ZN(n15542) );
  OAI221_X1 U17113 ( .B1(n15544), .B2(keyinput44), .C1(n15543), .C2(keyinput40), .A(n15542), .ZN(n15545) );
  NOR4_X1 U17114 ( .A1(n15548), .A2(n15547), .A3(n15546), .A4(n15545), .ZN(
        n15549) );
  NAND4_X1 U17115 ( .A1(n15552), .A2(n15551), .A3(n15550), .A4(n15549), .ZN(
        n15670) );
  AOI22_X1 U17116 ( .A1(n15555), .A2(keyinput84), .B1(keyinput30), .B2(n15554), 
        .ZN(n15553) );
  OAI221_X1 U17117 ( .B1(n15555), .B2(keyinput84), .C1(n15554), .C2(keyinput30), .A(n15553), .ZN(n15564) );
  AOI22_X1 U17118 ( .A1(n15557), .A2(keyinput109), .B1(keyinput120), .B2(
        n13786), .ZN(n15556) );
  OAI221_X1 U17119 ( .B1(n15557), .B2(keyinput109), .C1(n13786), .C2(
        keyinput120), .A(n15556), .ZN(n15563) );
  AOI22_X1 U17120 ( .A1(n15559), .A2(keyinput111), .B1(keyinput124), .B2(
        n10169), .ZN(n15558) );
  OAI221_X1 U17121 ( .B1(n15559), .B2(keyinput111), .C1(n10169), .C2(
        keyinput124), .A(n15558), .ZN(n15562) );
  AOI22_X1 U17122 ( .A1(n15676), .A2(keyinput100), .B1(keyinput74), .B2(n9083), 
        .ZN(n15560) );
  OAI221_X1 U17123 ( .B1(n15676), .B2(keyinput100), .C1(n9083), .C2(keyinput74), .A(n15560), .ZN(n15561) );
  NOR4_X1 U17124 ( .A1(n15564), .A2(n15563), .A3(n15562), .A4(n15561), .ZN(
        n15611) );
  AOI22_X1 U17125 ( .A1(n15567), .A2(keyinput4), .B1(keyinput35), .B2(n15566), 
        .ZN(n15565) );
  OAI221_X1 U17126 ( .B1(n15567), .B2(keyinput4), .C1(n15566), .C2(keyinput35), 
        .A(n15565), .ZN(n15578) );
  INV_X1 U17127 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n15569) );
  AOI22_X1 U17128 ( .A1(n15570), .A2(keyinput33), .B1(keyinput119), .B2(n15569), .ZN(n15568) );
  OAI221_X1 U17129 ( .B1(n15570), .B2(keyinput33), .C1(n15569), .C2(
        keyinput119), .A(n15568), .ZN(n15577) );
  INV_X1 U17130 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n15572) );
  AOI22_X1 U17131 ( .A1(n9039), .A2(keyinput56), .B1(n15572), .B2(keyinput64), 
        .ZN(n15571) );
  OAI221_X1 U17132 ( .B1(n9039), .B2(keyinput56), .C1(n15572), .C2(keyinput64), 
        .A(n15571), .ZN(n15576) );
  XOR2_X1 U17133 ( .A(n15674), .B(keyinput70), .Z(n15574) );
  XNOR2_X1 U17134 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput91), .ZN(n15573) );
  NAND2_X1 U17135 ( .A1(n15574), .A2(n15573), .ZN(n15575) );
  NOR4_X1 U17136 ( .A1(n15578), .A2(n15577), .A3(n15576), .A4(n15575), .ZN(
        n15610) );
  AOI22_X1 U17137 ( .A1(n15581), .A2(keyinput19), .B1(keyinput101), .B2(n15580), .ZN(n15579) );
  OAI221_X1 U17138 ( .B1(n15581), .B2(keyinput19), .C1(n15580), .C2(
        keyinput101), .A(n15579), .ZN(n15592) );
  INV_X1 U17139 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n15583) );
  AOI22_X1 U17140 ( .A1(n15584), .A2(keyinput118), .B1(keyinput49), .B2(n15583), .ZN(n15582) );
  OAI221_X1 U17141 ( .B1(n15584), .B2(keyinput118), .C1(n15583), .C2(
        keyinput49), .A(n15582), .ZN(n15591) );
  AOI22_X1 U17142 ( .A1(n15586), .A2(keyinput99), .B1(n15713), .B2(keyinput79), 
        .ZN(n15585) );
  OAI221_X1 U17143 ( .B1(n15586), .B2(keyinput99), .C1(n15713), .C2(keyinput79), .A(n15585), .ZN(n15590) );
  XNOR2_X1 U17144 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput52), .ZN(n15588) );
  XNOR2_X1 U17145 ( .A(keyinput67), .B(P3_REG2_REG_1__SCAN_IN), .ZN(n15587) );
  NAND2_X1 U17146 ( .A1(n15588), .A2(n15587), .ZN(n15589) );
  NOR4_X1 U17147 ( .A1(n15592), .A2(n15591), .A3(n15590), .A4(n15589), .ZN(
        n15609) );
  AOI22_X1 U17148 ( .A1(n15595), .A2(keyinput11), .B1(n15594), .B2(keyinput75), 
        .ZN(n15593) );
  OAI221_X1 U17149 ( .B1(n15595), .B2(keyinput11), .C1(n15594), .C2(keyinput75), .A(n15593), .ZN(n15607) );
  AOI22_X1 U17150 ( .A1(n15598), .A2(keyinput113), .B1(keyinput115), .B2(
        n15597), .ZN(n15596) );
  OAI221_X1 U17151 ( .B1(n15598), .B2(keyinput113), .C1(n15597), .C2(
        keyinput115), .A(n15596), .ZN(n15606) );
  INV_X1 U17152 ( .A(P2_WR_REG_SCAN_IN), .ZN(n15600) );
  AOI22_X1 U17153 ( .A1(n7739), .A2(keyinput69), .B1(keyinput48), .B2(n15600), 
        .ZN(n15599) );
  OAI221_X1 U17154 ( .B1(n7739), .B2(keyinput69), .C1(n15600), .C2(keyinput48), 
        .A(n15599), .ZN(n15605) );
  AOI22_X1 U17155 ( .A1(n15603), .A2(keyinput25), .B1(keyinput46), .B2(n15602), 
        .ZN(n15601) );
  OAI221_X1 U17156 ( .B1(n15603), .B2(keyinput25), .C1(n15602), .C2(keyinput46), .A(n15601), .ZN(n15604) );
  NOR4_X1 U17157 ( .A1(n15607), .A2(n15606), .A3(n15605), .A4(n15604), .ZN(
        n15608) );
  NAND4_X1 U17158 ( .A1(n15611), .A2(n15610), .A3(n15609), .A4(n15608), .ZN(
        n15669) );
  AOI22_X1 U17159 ( .A1(n15614), .A2(keyinput117), .B1(keyinput53), .B2(n15613), .ZN(n15612) );
  OAI221_X1 U17160 ( .B1(n15614), .B2(keyinput117), .C1(n15613), .C2(
        keyinput53), .A(n15612), .ZN(n15626) );
  AOI22_X1 U17161 ( .A1(n15617), .A2(keyinput10), .B1(n15616), .B2(keyinput116), .ZN(n15615) );
  OAI221_X1 U17162 ( .B1(n15617), .B2(keyinput10), .C1(n15616), .C2(
        keyinput116), .A(n15615), .ZN(n15625) );
  AOI22_X1 U17163 ( .A1(n15714), .A2(keyinput50), .B1(n15619), .B2(keyinput107), .ZN(n15618) );
  OAI221_X1 U17164 ( .B1(n15714), .B2(keyinput50), .C1(n15619), .C2(
        keyinput107), .A(n15618), .ZN(n15624) );
  AOI22_X1 U17165 ( .A1(n15622), .A2(keyinput47), .B1(keyinput3), .B2(n15621), 
        .ZN(n15620) );
  OAI221_X1 U17166 ( .B1(n15622), .B2(keyinput47), .C1(n15621), .C2(keyinput3), 
        .A(n15620), .ZN(n15623) );
  NOR4_X1 U17167 ( .A1(n15626), .A2(n15625), .A3(n15624), .A4(n15623), .ZN(
        n15667) );
  AOI22_X1 U17168 ( .A1(n15628), .A2(keyinput98), .B1(keyinput76), .B2(n8495), 
        .ZN(n15627) );
  OAI221_X1 U17169 ( .B1(n15628), .B2(keyinput98), .C1(n8495), .C2(keyinput76), 
        .A(n15627), .ZN(n15637) );
  AOI22_X1 U17170 ( .A1(n15630), .A2(keyinput125), .B1(n9977), .B2(keyinput55), 
        .ZN(n15629) );
  OAI221_X1 U17171 ( .B1(n15630), .B2(keyinput125), .C1(n9977), .C2(keyinput55), .A(n15629), .ZN(n15636) );
  XOR2_X1 U17172 ( .A(n9993), .B(keyinput58), .Z(n15634) );
  XOR2_X1 U17173 ( .A(n11418), .B(keyinput85), .Z(n15633) );
  XNOR2_X1 U17174 ( .A(P3_IR_REG_8__SCAN_IN), .B(keyinput34), .ZN(n15632) );
  XNOR2_X1 U17175 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput54), .ZN(n15631) );
  NAND4_X1 U17176 ( .A1(n15634), .A2(n15633), .A3(n15632), .A4(n15631), .ZN(
        n15635) );
  NOR3_X1 U17177 ( .A1(n15637), .A2(n15636), .A3(n15635), .ZN(n15666) );
  AOI22_X1 U17178 ( .A1(n15639), .A2(keyinput37), .B1(keyinput57), .B2(n8396), 
        .ZN(n15638) );
  OAI221_X1 U17179 ( .B1(n15639), .B2(keyinput37), .C1(n8396), .C2(keyinput57), 
        .A(n15638), .ZN(n15649) );
  AOI22_X1 U17180 ( .A1(n15675), .A2(keyinput103), .B1(n15641), .B2(keyinput97), .ZN(n15640) );
  OAI221_X1 U17181 ( .B1(n15675), .B2(keyinput103), .C1(n15641), .C2(
        keyinput97), .A(n15640), .ZN(n15648) );
  AOI22_X1 U17182 ( .A1(n15738), .A2(keyinput21), .B1(keyinput68), .B2(n15643), 
        .ZN(n15642) );
  OAI221_X1 U17183 ( .B1(n15738), .B2(keyinput21), .C1(n15643), .C2(keyinput68), .A(n15642), .ZN(n15647) );
  AOI22_X1 U17184 ( .A1(n15697), .A2(keyinput83), .B1(n15645), .B2(keyinput29), 
        .ZN(n15644) );
  OAI221_X1 U17185 ( .B1(n15697), .B2(keyinput83), .C1(n15645), .C2(keyinput29), .A(n15644), .ZN(n15646) );
  NOR4_X1 U17186 ( .A1(n15649), .A2(n15648), .A3(n15647), .A4(n15646), .ZN(
        n15665) );
  AOI22_X1 U17187 ( .A1(n15652), .A2(keyinput27), .B1(keyinput15), .B2(n15651), 
        .ZN(n15650) );
  OAI221_X1 U17188 ( .B1(n15652), .B2(keyinput27), .C1(n15651), .C2(keyinput15), .A(n15650), .ZN(n15663) );
  AOI22_X1 U17189 ( .A1(n15654), .A2(keyinput23), .B1(keyinput96), .B2(n11890), 
        .ZN(n15653) );
  OAI221_X1 U17190 ( .B1(n15654), .B2(keyinput23), .C1(n11890), .C2(keyinput96), .A(n15653), .ZN(n15662) );
  AOI22_X1 U17191 ( .A1(n15657), .A2(keyinput86), .B1(keyinput20), .B2(n15656), 
        .ZN(n15655) );
  OAI221_X1 U17192 ( .B1(n15657), .B2(keyinput86), .C1(n15656), .C2(keyinput20), .A(n15655), .ZN(n15661) );
  XNOR2_X1 U17193 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(keyinput43), .ZN(n15659)
         );
  XNOR2_X1 U17194 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput121), .ZN(n15658) );
  NAND2_X1 U17195 ( .A1(n15659), .A2(n15658), .ZN(n15660) );
  NOR4_X1 U17196 ( .A1(n15663), .A2(n15662), .A3(n15661), .A4(n15660), .ZN(
        n15664) );
  NAND4_X1 U17197 ( .A1(n15667), .A2(n15666), .A3(n15665), .A4(n15664), .ZN(
        n15668) );
  NOR4_X1 U17198 ( .A1(n15671), .A2(n15670), .A3(n15669), .A4(n15668), .ZN(
        n15672) );
  XNOR2_X1 U17199 ( .A(n15673), .B(n15672), .ZN(n15733) );
  NOR4_X1 U17200 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_REG0_REG_6__SCAN_IN), 
        .A3(P1_REG2_REG_5__SCAN_IN), .A4(P1_REG0_REG_4__SCAN_IN), .ZN(n15731)
         );
  NOR4_X1 U17201 ( .A1(P2_REG0_REG_13__SCAN_IN), .A2(P2_REG3_REG_0__SCAN_IN), 
        .A3(P2_REG0_REG_7__SCAN_IN), .A4(P1_REG0_REG_24__SCAN_IN), .ZN(n15730)
         );
  NAND4_X1 U17202 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .A3(P2_REG3_REG_16__SCAN_IN), .A4(P1_IR_REG_9__SCAN_IN), .ZN(n15683)
         );
  NAND4_X1 U17203 ( .A1(P3_DATAO_REG_2__SCAN_IN), .A2(n15676), .A3(n15675), 
        .A4(n15674), .ZN(n15682) );
  NOR4_X1 U17204 ( .A1(P2_REG2_REG_21__SCAN_IN), .A2(P2_REG1_REG_15__SCAN_IN), 
        .A3(P1_REG2_REG_15__SCAN_IN), .A4(P1_REG1_REG_15__SCAN_IN), .ZN(n15680) );
  NOR4_X1 U17205 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG1_REG_14__SCAN_IN), 
        .A3(P1_REG3_REG_2__SCAN_IN), .A4(P3_ADDR_REG_8__SCAN_IN), .ZN(n15679)
         );
  NOR4_X1 U17206 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(P1_DATAO_REG_14__SCAN_IN), .A3(P3_REG1_REG_23__SCAN_IN), .A4(P3_REG1_REG_15__SCAN_IN), .ZN(n15678) );
  NOR4_X1 U17207 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(P1_DATAO_REG_26__SCAN_IN), 
        .A3(P1_DATAO_REG_13__SCAN_IN), .A4(P2_REG2_REG_22__SCAN_IN), .ZN(
        n15677) );
  NAND4_X1 U17208 ( .A1(n15680), .A2(n15679), .A3(n15678), .A4(n15677), .ZN(
        n15681) );
  NOR3_X1 U17209 ( .A1(n15683), .A2(n15682), .A3(n15681), .ZN(n15729) );
  OR4_X1 U17210 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_1__SCAN_IN), 
        .A3(P2_ADDR_REG_5__SCAN_IN), .A4(n10442), .ZN(n15727) );
  NAND4_X1 U17211 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_REG3_REG_5__SCAN_IN), 
        .A3(SI_13_), .A4(P1_IR_REG_18__SCAN_IN), .ZN(n15687) );
  NAND4_X1 U17212 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_REG1_REG_30__SCAN_IN), 
        .A3(P3_REG1_REG_25__SCAN_IN), .A4(P3_DATAO_REG_5__SCAN_IN), .ZN(n15686) );
  NAND4_X1 U17213 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_REG0_REG_23__SCAN_IN), 
        .A3(P1_REG2_REG_21__SCAN_IN), .A4(P1_REG0_REG_21__SCAN_IN), .ZN(n15685) );
  NAND4_X1 U17214 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_REG1_REG_29__SCAN_IN), 
        .A3(P1_REG1_REG_31__SCAN_IN), .A4(P1_REG0_REG_31__SCAN_IN), .ZN(n15684) );
  NOR4_X1 U17215 ( .A1(n15687), .A2(n15686), .A3(n15685), .A4(n15684), .ZN(
        n15705) );
  NAND4_X1 U17216 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG2_REG_23__SCAN_IN), 
        .A3(P2_REG2_REG_16__SCAN_IN), .A4(P1_REG0_REG_16__SCAN_IN), .ZN(n15691) );
  NAND4_X1 U17217 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(P1_REG0_REG_17__SCAN_IN), 
        .A3(P1_REG0_REG_12__SCAN_IN), .A4(P1_REG1_REG_10__SCAN_IN), .ZN(n15690) );
  NAND4_X1 U17218 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(P3_REG2_REG_26__SCAN_IN), .A3(P1_REG3_REG_8__SCAN_IN), .A4(P3_DATAO_REG_1__SCAN_IN), .ZN(n15689) );
  NAND4_X1 U17219 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(
        P1_DATAO_REG_12__SCAN_IN), .A3(P2_DATAO_REG_22__SCAN_IN), .A4(
        P2_REG2_REG_17__SCAN_IN), .ZN(n15688) );
  NOR4_X1 U17220 ( .A1(n15691), .A2(n15690), .A3(n15689), .A4(n15688), .ZN(
        n15704) );
  NOR4_X1 U17221 ( .A1(P2_D_REG_1__SCAN_IN), .A2(P2_REG3_REG_13__SCAN_IN), 
        .A3(P2_REG3_REG_10__SCAN_IN), .A4(P3_DATAO_REG_26__SCAN_IN), .ZN(
        n15695) );
  NOR4_X1 U17222 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), 
        .A3(P3_DATAO_REG_29__SCAN_IN), .A4(P3_DATAO_REG_20__SCAN_IN), .ZN(
        n15694) );
  NOR4_X1 U17223 ( .A1(P2_D_REG_13__SCAN_IN), .A2(SI_9_), .A3(SI_5_), .A4(
        P2_REG1_REG_27__SCAN_IN), .ZN(n15693) );
  NOR4_X1 U17224 ( .A1(P3_REG0_REG_27__SCAN_IN), .A2(P3_REG0_REG_25__SCAN_IN), 
        .A3(P3_REG2_REG_6__SCAN_IN), .A4(P3_REG1_REG_9__SCAN_IN), .ZN(n15692)
         );
  AND4_X1 U17225 ( .A1(n15695), .A2(n15694), .A3(n15693), .A4(n15692), .ZN(
        n15703) );
  NAND4_X1 U17226 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(
        P2_DATAO_REG_30__SCAN_IN), .A3(P1_REG2_REG_10__SCAN_IN), .A4(
        P1_REG1_REG_7__SCAN_IN), .ZN(n15701) );
  NAND4_X1 U17227 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_REG3_REG_5__SCAN_IN), 
        .A3(P1_REG0_REG_20__SCAN_IN), .A4(P1_REG1_REG_9__SCAN_IN), .ZN(n15700)
         );
  NAND4_X1 U17228 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(P3_REG3_REG_27__SCAN_IN), 
        .A3(n15697), .A4(n15696), .ZN(n15699) );
  NAND4_X1 U17229 ( .A1(SI_30_), .A2(P3_REG2_REG_27__SCAN_IN), .A3(
        P3_REG2_REG_24__SCAN_IN), .A4(P3_REG0_REG_22__SCAN_IN), .ZN(n15698) );
  NOR4_X1 U17230 ( .A1(n15701), .A2(n15700), .A3(n15699), .A4(n15698), .ZN(
        n15702) );
  NAND4_X1 U17231 ( .A1(n15705), .A2(n15704), .A3(n15703), .A4(n15702), .ZN(
        n15726) );
  NOR3_X1 U17232 ( .A1(n15707), .A2(n15706), .A3(P3_IR_REG_7__SCAN_IN), .ZN(
        n15709) );
  NOR2_X1 U17233 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n15708) );
  NAND4_X1 U17234 ( .A1(n15709), .A2(n15708), .A3(P1_WR_REG_SCAN_IN), .A4(
        P2_WR_REG_SCAN_IN), .ZN(n15712) );
  NAND4_X1 U17235 ( .A1(P3_B_REG_SCAN_IN), .A2(P3_REG1_REG_2__SCAN_IN), .A3(
        P3_D_REG_30__SCAN_IN), .A4(n15710), .ZN(n15711) );
  NOR2_X1 U17236 ( .A1(n15712), .A2(n15711), .ZN(n15724) );
  NAND4_X1 U17237 ( .A1(P2_RD_REG_SCAN_IN), .A2(P3_D_REG_4__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(n15713), .ZN(n15720) );
  NAND4_X1 U17238 ( .A1(P3_REG2_REG_1__SCAN_IN), .A2(P1_REG1_REG_2__SCAN_IN), 
        .A3(P3_ADDR_REG_12__SCAN_IN), .A4(n15714), .ZN(n15719) );
  NAND4_X1 U17239 ( .A1(n15717), .A2(n15716), .A3(n15715), .A4(
        P3_IR_REG_8__SCAN_IN), .ZN(n15718) );
  NOR3_X1 U17240 ( .A1(n15720), .A2(n15719), .A3(n15718), .ZN(n15722) );
  NAND4_X1 U17241 ( .A1(n15724), .A2(n15723), .A3(n15722), .A4(n15721), .ZN(
        n15725) );
  NOR3_X1 U17242 ( .A1(n15727), .A2(n15726), .A3(n15725), .ZN(n15728) );
  NAND4_X1 U17243 ( .A1(n15731), .A2(n15730), .A3(n15729), .A4(n15728), .ZN(
        n15732) );
  XNOR2_X1 U17244 ( .A(n15733), .B(n15732), .ZN(P3_U3158) );
  AOI21_X1 U17245 ( .B1(n15736), .B2(n15735), .A(n15734), .ZN(SUB_1596_U59) );
  OAI21_X1 U17246 ( .B1(n15739), .B2(n15738), .A(n15737), .ZN(SUB_1596_U58) );
  XNOR2_X1 U17247 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15740), .ZN(SUB_1596_U53)
         );
  AOI21_X1 U17248 ( .B1(n15743), .B2(n15742), .A(n15741), .ZN(SUB_1596_U56) );
  OAI21_X1 U17249 ( .B1(n15745), .B2(n10459), .A(n15744), .ZN(SUB_1596_U60) );
  AOI21_X1 U17250 ( .B1(n15748), .B2(n15747), .A(n15746), .ZN(SUB_1596_U5) );
  AND2_X2 U7356 ( .A1(n7342), .A2(n7341), .ZN(n8004) );
  AND3_X1 U9610 ( .A1(n6802), .A2(n6803), .A3(n6678), .ZN(n8643) );
  AND2_X1 U7368 ( .A1(n12032), .A2(n6621), .ZN(n7718) );
  AOI21_X1 U7364 ( .B1(n7464), .B2(n7583), .A(n6646), .ZN(n7462) );
  NAND3_X2 U7449 ( .A1(n8119), .A2(n8120), .A3(n8118), .ZN(n7609) );
  NAND2_X1 U9679 ( .A1(n6975), .A2(n7951), .ZN(n12441) );
  NOR2_X1 U7317 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n9804) );
  CLKBUF_X1 U7348 ( .A(n9566), .Z(n9655) );
  AND2_X1 U7354 ( .A1(n6837), .A2(n6836), .ZN(n13006) );
  INV_X1 U7472 ( .A(n12946), .ZN(n10764) );
  NAND2_X2 U7473 ( .A1(n12652), .A2(n12946), .ZN(n8675) );
  CLKBUF_X1 U8015 ( .A(n8888), .Z(n7223) );
  CLKBUF_X1 U9628 ( .A(n14753), .Z(n6548) );
endmodule

