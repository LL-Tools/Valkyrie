

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9628, n9629, n9630, n9631, n9632, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,
         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,
         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,
         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,
         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,
         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
         n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
         n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,
         n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,
         n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
         n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
         n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312,
         n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
         n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
         n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,
         n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,
         n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
         n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368,
         n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,
         n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,
         n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
         n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400,
         n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
         n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,
         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
         n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440,
         n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
         n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456,
         n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,
         n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472,
         n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
         n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,
         n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
         n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
         n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,
         n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
         n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,
         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,
         n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600,
         n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
         n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,
         n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
         n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,
         n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
         n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,
         n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
         n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,
         n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
         n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064,
         n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072,
         n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080,
         n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088,
         n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,
         n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,
         n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,
         n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
         n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
         n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,
         n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144,
         n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
         n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,
         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
         n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
         n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,
         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,
         n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
         n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,
         n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
         n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,
         n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,
         n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
         n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
         n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
         n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,
         n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,
         n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
         n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
         n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,
         n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360,
         n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
         n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,
         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,
         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496,
         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
         n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
         n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536,
         n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,
         n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
         n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
         n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
         n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
         n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608,
         n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,
         n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
         n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
         n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
         n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
         n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
         n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664,
         n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
         n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680,
         n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688,
         n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,
         n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
         n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712,
         n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,
         n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
         n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736,
         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,
         n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
         n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808,
         n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
         n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824,
         n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
         n20833, n20834, n20835, n20836, n20837, n20838, n20839;

  AOI21_X1 U11029 ( .B1(n15653), .B2(n15652), .A(n15651), .ZN(n15663) );
  AND2_X1 U11030 ( .A1(n12127), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20020)
         );
  NOR2_X1 U11031 ( .A1(n17280), .A2(n17457), .ZN(n17276) );
  NAND2_X1 U11032 ( .A1(n11002), .A2(n13968), .ZN(n9818) );
  INV_X2 U11033 ( .A(n14841), .ZN(n14844) );
  NAND2_X1 U11034 ( .A1(n13777), .A2(n13778), .ZN(n13917) );
  NAND2_X1 U11035 ( .A1(n11594), .A2(n11593), .ZN(n13610) );
  NAND2_X1 U11036 ( .A1(n13961), .A2(n12733), .ZN(n13777) );
  INV_X2 U11037 ( .A(n12874), .ZN(n14841) );
  INV_X2 U11038 ( .A(n16531), .ZN(n16837) );
  NAND3_X2 U11039 ( .A1(n10297), .A2(n10296), .A3(n10295), .ZN(n18204) );
  AOI211_X1 U11040 ( .C1(n14285), .C2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n10294), .B(n10293), .ZN(n10295) );
  OR2_X1 U11041 ( .A1(n9610), .A2(n10619), .ZN(n9609) );
  AND2_X1 U11043 ( .A1(n10515), .A2(n10430), .ZN(n12460) );
  AND2_X1 U11044 ( .A1(n10672), .A2(n12429), .ZN(n10673) );
  CLKBUF_X1 U11045 ( .A(n10675), .Z(n12625) );
  CLKBUF_X1 U11046 ( .A(n10153), .Z(n17140) );
  INV_X1 U11047 ( .A(n16952), .ZN(n10280) );
  CLKBUF_X1 U11048 ( .A(n10279), .Z(n17124) );
  CLKBUF_X2 U11049 ( .A(n10153), .Z(n17018) );
  INV_X2 U11050 ( .A(n17155), .ZN(n10141) );
  INV_X1 U11051 ( .A(n16983), .ZN(n17158) );
  CLKBUF_X2 U11053 ( .A(n11250), .Z(n12026) );
  CLKBUF_X2 U11054 ( .A(n11530), .Z(n9592) );
  CLKBUF_X2 U11055 ( .A(n11305), .Z(n12020) );
  CLKBUF_X2 U11056 ( .A(n10551), .Z(n19765) );
  NAND2_X1 U11057 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10103) );
  AND2_X1 U11058 ( .A1(n11370), .A2(n13570), .ZN(n11397) );
  CLKBUF_X1 U11059 ( .A(n11379), .Z(n20044) );
  AND4_X1 U11060 ( .A1(n11332), .A2(n11331), .A3(n11330), .A4(n11329), .ZN(
        n11338) );
  AND2_X1 U11061 ( .A1(n13564), .A2(n11234), .ZN(n11273) );
  AND2_X2 U11062 ( .A1(n10671), .A2(n13699), .ZN(n10677) );
  AND2_X1 U11063 ( .A1(n13590), .A2(n13575), .ZN(n11305) );
  AND2_X1 U11064 ( .A1(n9763), .A2(n11233), .ZN(n11283) );
  AND2_X1 U11065 ( .A1(n11235), .A2(n11233), .ZN(n11300) );
  AND2_X2 U11066 ( .A1(n13575), .A2(n13564), .ZN(n11496) );
  AND2_X2 U11067 ( .A1(n13590), .A2(n11234), .ZN(n11266) );
  AND2_X1 U11068 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11234) );
  AND2_X2 U11069 ( .A1(n11554), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11232) );
  NAND2_X2 U11070 ( .A1(n18613), .A2(n18130), .ZN(n18028) );
  AND2_X1 U11071 ( .A1(n10663), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12392) );
  CLKBUF_X2 U11073 ( .A(n11300), .Z(n12028) );
  AND2_X2 U11074 ( .A1(n11225), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11235) );
  NOR2_X1 U11075 ( .A1(n11586), .A2(n9767), .ZN(n9766) );
  BUF_X2 U11076 ( .A(n11255), .Z(n12018) );
  AND4_X1 U11077 ( .A1(n11291), .A2(n11290), .A3(n11289), .A4(n11288), .ZN(
        n11292) );
  XNOR2_X1 U11078 ( .A(n11586), .B(n11585), .ZN(n12838) );
  AND2_X1 U11081 ( .A1(n12596), .A2(n10430), .ZN(n12464) );
  AND2_X1 U11082 ( .A1(n9587), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12380) );
  AND2_X2 U11083 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10674) );
  NOR2_X1 U11084 ( .A1(n18195), .A2(n10319), .ZN(n10391) );
  INV_X1 U11085 ( .A(n17037), .ZN(n16900) );
  NAND2_X1 U11086 ( .A1(n12921), .A2(n12946), .ZN(n13025) );
  INV_X1 U11087 ( .A(n13285), .ZN(n13630) );
  OR2_X1 U11088 ( .A1(n11380), .A2(n11381), .ZN(n14302) );
  XNOR2_X1 U11089 ( .A(n9602), .B(n20154), .ZN(n20642) );
  AND2_X1 U11091 ( .A1(n12596), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10714) );
  INV_X1 U11092 ( .A(n19835), .ZN(n19812) );
  OR2_X1 U11093 ( .A1(n13461), .A2(n13460), .ZN(n13535) );
  AOI211_X1 U11095 ( .C1(n13412), .C2(n13731), .A(n13712), .B(n13711), .ZN(
        n15767) );
  NOR2_X2 U11096 ( .A1(n17312), .A2(n10176), .ZN(n17722) );
  INV_X1 U11097 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10070) );
  INV_X1 U11098 ( .A(n17723), .ZN(n17632) );
  INV_X1 U11099 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18771) );
  AND2_X1 U11100 ( .A1(n9605), .A2(n9764), .ZN(n9585) );
  NOR2_X4 U11101 ( .A1(n12680), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12770) );
  INV_X2 U11102 ( .A(n12530), .ZN(n9630) );
  INV_X2 U11103 ( .A(n12530), .ZN(n9629) );
  NOR2_X2 U11104 ( .A1(n15068), .A2(n15070), .ZN(n15069) );
  INV_X1 U11105 ( .A(n9600), .ZN(n15384) );
  AND2_X2 U11106 ( .A1(n16264), .A2(n9740), .ZN(n9600) );
  NOR2_X2 U11107 ( .A1(n14013), .A2(n9708), .ZN(n11704) );
  NOR2_X2 U11108 ( .A1(n17761), .A2(n17775), .ZN(n16798) );
  AND2_X1 U11109 ( .A1(n11235), .A2(n11233), .ZN(n9586) );
  AOI21_X2 U11110 ( .B1(n15347), .B2(n15334), .A(n15333), .ZN(n15338) );
  NOR2_X2 U11111 ( .A1(n15078), .A2(n12547), .ZN(n12569) );
  NOR2_X2 U11112 ( .A1(n15077), .A2(n15079), .ZN(n15078) );
  NAND2_X2 U11113 ( .A1(n14095), .A2(n10885), .ZN(n14157) );
  INV_X2 U11114 ( .A(n18161), .ZN(n10392) );
  AND2_X1 U11115 ( .A1(n10663), .A2(n10430), .ZN(n12379) );
  NAND2_X2 U11116 ( .A1(n13299), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13298) );
  AND2_X2 U11117 ( .A1(n13672), .A2(n9718), .ZN(n13895) );
  INV_X4 U11118 ( .A(n10166), .ZN(n17151) );
  INV_X2 U11119 ( .A(n10099), .ZN(n10166) );
  AND2_X2 U11120 ( .A1(n10671), .A2(n13699), .ZN(n9587) );
  NAND2_X2 U11121 ( .A1(n15093), .A2(n10091), .ZN(n15085) );
  AOI21_X2 U11122 ( .B1(n15373), .B2(n15371), .A(n15360), .ZN(n15361) );
  AND2_X1 U11123 ( .A1(n11232), .A2(n13590), .ZN(n11977) );
  XNOR2_X2 U11124 ( .A(n10784), .B(n10785), .ZN(n13819) );
  NAND2_X2 U11125 ( .A1(n10766), .A2(n10765), .ZN(n10784) );
  AND2_X2 U11126 ( .A1(n10671), .A2(n10596), .ZN(n9588) );
  AND2_X2 U11127 ( .A1(n10671), .A2(n10596), .ZN(n10663) );
  INV_X4 U11128 ( .A(n10089), .ZN(n17123) );
  INV_X2 U11129 ( .A(n12678), .ZN(n15217) );
  NOR2_X1 U11130 ( .A1(n15065), .A2(n11207), .ZN(n15044) );
  NOR2_X1 U11131 ( .A1(n16552), .A2(n16553), .ZN(n16551) );
  NOR2_X2 U11132 ( .A1(n17422), .A2(n17227), .ZN(n17223) );
  NAND2_X1 U11133 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17228), .ZN(n17227) );
  INV_X2 U11134 ( .A(n17811), .ZN(n17798) );
  XNOR2_X1 U11135 ( .A(n12843), .B(n12936), .ZN(n19964) );
  AOI21_X1 U11136 ( .B1(n11086), .B2(n11094), .A(n11085), .ZN(n11084) );
  NAND2_X1 U11137 ( .A1(n11504), .A2(n11503), .ZN(n20154) );
  NOR2_X1 U11138 ( .A1(n13440), .A2(n12711), .ZN(n13804) );
  NAND2_X1 U11139 ( .A1(n10621), .A2(n9816), .ZN(n10594) );
  NOR2_X2 U11140 ( .A1(n13535), .A2(n13536), .ZN(n13615) );
  NAND3_X1 U11141 ( .A1(n9821), .A2(n10578), .A3(n9822), .ZN(n10595) );
  CLKBUF_X2 U11142 ( .A(n12714), .Z(n12757) );
  INV_X2 U11143 ( .A(n10549), .ZN(n10553) );
  NAND2_X2 U11144 ( .A1(n20024), .A2(n11366), .ZN(n13163) );
  NAND2_X2 U11145 ( .A1(n10433), .A2(n10432), .ZN(n9622) );
  INV_X1 U11146 ( .A(n12911), .ZN(n13544) );
  INV_X2 U11147 ( .A(n11367), .ZN(n11366) );
  AND4_X1 U11148 ( .A1(n11324), .A2(n11323), .A3(n11322), .A4(n11321), .ZN(
        n11340) );
  INV_X1 U11149 ( .A(n12623), .ZN(n9589) );
  BUF_X2 U11150 ( .A(n11410), .Z(n12027) );
  CLKBUF_X3 U11151 ( .A(n10665), .Z(n12596) );
  BUF_X2 U11152 ( .A(n11278), .Z(n12019) );
  CLKBUF_X2 U11153 ( .A(n11995), .Z(n11643) );
  CLKBUF_X2 U11154 ( .A(n11283), .Z(n12025) );
  CLKBUF_X2 U11155 ( .A(n11273), .Z(n11825) );
  INV_X1 U11156 ( .A(n9863), .ZN(n14755) );
  NAND2_X1 U11157 ( .A1(n10019), .A2(n10017), .ZN(n10020) );
  NAND2_X1 U11158 ( .A1(n9743), .A2(n9697), .ZN(n10019) );
  NOR2_X1 U11159 ( .A1(n15284), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15547) );
  OAI21_X1 U11160 ( .B1(n14603), .B2(n20022), .A(n9783), .ZN(n9782) );
  OAI21_X1 U11161 ( .B1(n14374), .B2(n14360), .A(n14361), .ZN(n14603) );
  AND2_X1 U11162 ( .A1(n15289), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15342) );
  NAND2_X1 U11163 ( .A1(n14649), .A2(n14844), .ZN(n14625) );
  OAI21_X1 U11164 ( .B1(n15418), .B2(n9994), .A(n9992), .ZN(n15308) );
  NOR2_X1 U11165 ( .A1(n15322), .A2(n15321), .ZN(n15325) );
  NAND2_X1 U11166 ( .A1(n9833), .A2(n9830), .ZN(n15418) );
  INV_X1 U11167 ( .A(n16265), .ZN(n11017) );
  NAND2_X1 U11168 ( .A1(n9867), .A2(n9866), .ZN(n14674) );
  NAND2_X1 U11169 ( .A1(n11013), .A2(n11012), .ZN(n16265) );
  OR2_X1 U11170 ( .A1(n14934), .A2(n14933), .ZN(n15499) );
  AND2_X1 U11171 ( .A1(n11003), .A2(n9711), .ZN(n9817) );
  OR2_X1 U11172 ( .A1(n12477), .A2(n12498), .ZN(n10091) );
  XNOR2_X1 U11173 ( .A(n15044), .B(n15043), .ZN(n15235) );
  NAND2_X1 U11174 ( .A1(n12882), .A2(n10023), .ZN(n14729) );
  NAND2_X1 U11175 ( .A1(n14087), .A2(n12880), .ZN(n12882) );
  AOI211_X1 U11176 ( .C1(n16548), .C2(n16894), .A(n16538), .B(n16537), .ZN(
        n16539) );
  OR2_X1 U11177 ( .A1(n15063), .A2(n15062), .ZN(n15065) );
  OAI21_X1 U11178 ( .B1(n13818), .B2(n13817), .A(n10995), .ZN(n14029) );
  NOR2_X1 U11179 ( .A1(n16551), .A2(n16837), .ZN(n16543) );
  NAND2_X1 U11180 ( .A1(n10875), .A2(n10874), .ZN(n10906) );
  AND2_X1 U11181 ( .A1(n17590), .A2(n10405), .ZN(n17521) );
  XNOR2_X1 U11182 ( .A(n10877), .B(n10873), .ZN(n10972) );
  NOR2_X1 U11183 ( .A1(n10029), .A2(n10027), .ZN(n10026) );
  NAND2_X1 U11184 ( .A1(n9703), .A2(n12891), .ZN(n10037) );
  AOI21_X1 U11185 ( .B1(n12891), .B2(n10036), .A(n10035), .ZN(n10034) );
  INV_X1 U11186 ( .A(n10873), .ZN(n10876) );
  NAND2_X1 U11187 ( .A1(n10872), .A2(n10871), .ZN(n10879) );
  INV_X1 U11188 ( .A(n14696), .ZN(n10035) );
  AND2_X1 U11189 ( .A1(n12881), .A2(n9868), .ZN(n10023) );
  NAND2_X1 U11190 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17702), .ZN(n17663) );
  OR2_X1 U11191 ( .A1(n12873), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16045) );
  AND2_X1 U11192 ( .A1(n12861), .A2(n12860), .ZN(n16050) );
  AND2_X1 U11193 ( .A1(n14864), .A2(n14865), .ZN(n14696) );
  OR2_X1 U11194 ( .A1(n10852), .A2(n10851), .ZN(n10872) );
  AND2_X1 U11195 ( .A1(n10832), .A2(n10831), .ZN(n10873) );
  OR2_X1 U11196 ( .A1(n10813), .A2(n10812), .ZN(n10832) );
  NAND2_X1 U11197 ( .A1(n14419), .A2(n14401), .ZN(n14403) );
  INV_X1 U11198 ( .A(n19964), .ZN(n9590) );
  NAND2_X1 U11199 ( .A1(n12842), .A2(n12841), .ZN(n12843) );
  NAND2_X1 U11200 ( .A1(n10377), .A2(n17710), .ZN(n18013) );
  NAND2_X1 U11201 ( .A1(n11517), .A2(n9657), .ZN(n12803) );
  NAND2_X1 U11202 ( .A1(n13457), .A2(n11578), .ZN(n13532) );
  NOR2_X1 U11203 ( .A1(n10653), .A2(n10652), .ZN(n10661) );
  NAND2_X1 U11204 ( .A1(n12155), .A2(n12154), .ZN(n13410) );
  NAND2_X1 U11205 ( .A1(n17276), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17275) );
  AOI211_X1 U11206 ( .C1(n19089), .C2(n19737), .A(n19131), .B(n19520), .ZN(
        n19084) );
  AND2_X1 U11207 ( .A1(n13194), .A2(n12145), .ZN(n13257) );
  XNOR2_X1 U11208 ( .A(n12164), .B(n12165), .ZN(n13411) );
  NAND2_X1 U11209 ( .A1(n12163), .A2(n12162), .ZN(n12164) );
  NAND2_X1 U11210 ( .A1(n13270), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20005) );
  CLKBUF_X1 U11211 ( .A(n12822), .Z(n20268) );
  AND2_X1 U11212 ( .A1(n10657), .A2(n10654), .ZN(n19409) );
  NAND2_X1 U11213 ( .A1(n9948), .A2(n9815), .ZN(n10634) );
  NOR2_X2 U11214 ( .A1(n11069), .A2(n10961), .ZN(n11054) );
  NAND2_X1 U11215 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n10214), .ZN(
        n17995) );
  CLKBUF_X1 U11216 ( .A(n14534), .Z(n16010) );
  CLKBUF_X1 U11217 ( .A(n12128), .Z(n16011) );
  NAND2_X1 U11218 ( .A1(n11024), .A2(n11034), .ZN(n11069) );
  NOR2_X1 U11219 ( .A1(n16633), .A2(n16837), .ZN(n16627) );
  XNOR2_X1 U11220 ( .A(n11482), .B(n11481), .ZN(n9764) );
  NOR2_X1 U11221 ( .A1(n17555), .A2(n16634), .ZN(n16633) );
  NOR2_X2 U11222 ( .A1(n19098), .A2(n19523), .ZN(n19099) );
  OAI22_X1 U11223 ( .A1(n13568), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n12830), 
        .B2(n11490), .ZN(n11482) );
  NOR2_X2 U11224 ( .A1(n19086), .A2(n19523), .ZN(n19087) );
  NOR2_X2 U11225 ( .A1(n19110), .A2(n19523), .ZN(n19111) );
  NAND2_X1 U11226 ( .A1(n20272), .A2(n20556), .ZN(n11504) );
  NOR2_X1 U11227 ( .A1(n16641), .A2(n16837), .ZN(n16634) );
  INV_X1 U11228 ( .A(n9815), .ZN(n19079) );
  NAND2_X1 U11229 ( .A1(n10594), .A2(n10593), .ZN(n10620) );
  NAND2_X1 U11230 ( .A1(n11483), .A2(n9780), .ZN(n13568) );
  INV_X1 U11231 ( .A(n12141), .ZN(n13728) );
  NAND2_X1 U11232 ( .A1(n11455), .A2(n11454), .ZN(n11565) );
  OAI211_X2 U11233 ( .C1(n9781), .C2(n9779), .A(n11466), .B(n9778), .ZN(n11483) );
  NAND2_X1 U11234 ( .A1(n13615), .A2(n13614), .ZN(n13682) );
  INV_X2 U11235 ( .A(n17430), .ZN(n17454) );
  NOR2_X2 U11236 ( .A1(n10974), .A2(n10973), .ZN(n11000) );
  NAND2_X1 U11237 ( .A1(n11392), .A2(n11391), .ZN(n11438) );
  NAND2_X1 U11238 ( .A1(n10993), .A2(n10992), .ZN(n10974) );
  AND2_X1 U11239 ( .A1(n13378), .A2(n13377), .ZN(n13380) );
  AOI211_X1 U11240 ( .C1(n10389), .C2(n10388), .A(n10387), .B(n10386), .ZN(
        n10398) );
  OR2_X1 U11241 ( .A1(n15046), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10586) );
  NAND2_X1 U11242 ( .A1(n11407), .A2(n11406), .ZN(n11436) );
  NOR2_X1 U11243 ( .A1(n16684), .A2(n16837), .ZN(n16673) );
  NOR2_X1 U11244 ( .A1(n13683), .A2(n14004), .ZN(n9918) );
  OR2_X1 U11245 ( .A1(n10393), .A2(n16485), .ZN(n10396) );
  NAND2_X1 U11246 ( .A1(n10600), .A2(n13196), .ZN(n10585) );
  NAND2_X1 U11247 ( .A1(n9826), .A2(n9825), .ZN(n10571) );
  CLKBUF_X1 U11248 ( .A(n9615), .Z(n12694) );
  AND2_X1 U11249 ( .A1(n10565), .A2(n13330), .ZN(n13196) );
  NAND2_X1 U11250 ( .A1(n10542), .A2(n12657), .ZN(n10561) );
  AND2_X1 U11251 ( .A1(n10565), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10583) );
  NAND2_X1 U11252 ( .A1(n10525), .A2(n9621), .ZN(n12657) );
  OR2_X1 U11253 ( .A1(n13565), .A2(n9776), .ZN(n9775) );
  INV_X1 U11255 ( .A(n12652), .ZN(n10537) );
  NAND2_X1 U11256 ( .A1(n13630), .A2(n12949), .ZN(n13016) );
  NAND2_X1 U11257 ( .A1(n12943), .A2(n11374), .ZN(n13036) );
  NOR2_X1 U11258 ( .A1(n10524), .A2(n10540), .ZN(n10525) );
  AND2_X1 U11259 ( .A1(n13334), .A2(n19765), .ZN(n9621) );
  AND2_X1 U11260 ( .A1(n13330), .A2(n10539), .ZN(n12660) );
  OR2_X1 U11261 ( .A1(n12946), .A2(n13009), .ZN(n12990) );
  AND2_X1 U11262 ( .A1(n11361), .A2(n9768), .ZN(n13028) );
  AND2_X1 U11263 ( .A1(n11377), .A2(n13290), .ZN(n11398) );
  AND2_X1 U11264 ( .A1(n10530), .A2(n10553), .ZN(n10534) );
  NAND2_X4 U11265 ( .A1(n12922), .A2(n12949), .ZN(n12943) );
  INV_X1 U11266 ( .A(n13163), .ZN(n13627) );
  AND2_X1 U11267 ( .A1(n10584), .A2(n10529), .ZN(n13334) );
  INV_X1 U11268 ( .A(n10551), .ZN(n13691) );
  OR2_X1 U11269 ( .A1(n12917), .A2(n20556), .ZN(n11490) );
  NAND2_X4 U11270 ( .A1(n12070), .A2(n11379), .ZN(n11368) );
  INV_X1 U11272 ( .A(n12909), .ZN(n13033) );
  AND2_X1 U11273 ( .A1(n17487), .A2(n9940), .ZN(n16364) );
  NAND2_X1 U11274 ( .A1(n10458), .A2(n10457), .ZN(n10529) );
  INV_X1 U11275 ( .A(n10538), .ZN(n12677) );
  INV_X4 U11276 ( .A(n11372), .ZN(n20024) );
  INV_X1 U11277 ( .A(n11371), .ZN(n20040) );
  NAND2_X1 U11278 ( .A1(n10077), .A2(n10518), .ZN(n10519) );
  NAND2_X1 U11279 ( .A1(n10431), .A2(n10430), .ZN(n10432) );
  NAND4_X1 U11280 ( .A1(n10494), .A2(n10493), .A3(n10492), .A4(n10491), .ZN(
        n10495) );
  OR2_X2 U11281 ( .A1(n11271), .A2(n11272), .ZN(n13290) );
  NAND4_X2 U11282 ( .A1(n11295), .A2(n11294), .A3(n11293), .A4(n11292), .ZN(
        n11376) );
  OR2_X1 U11283 ( .A1(n11431), .A2(n11430), .ZN(n12876) );
  INV_X2 U11284 ( .A(U212), .ZN(n16440) );
  OR2_X2 U11285 ( .A1(n11261), .A2(n11260), .ZN(n11371) );
  OR2_X2 U11286 ( .A1(n16441), .A2(n16384), .ZN(n16443) );
  AND4_X2 U11287 ( .A1(n11317), .A2(n11316), .A3(n11315), .A4(n11314), .ZN(
        n12911) );
  NAND2_X1 U11288 ( .A1(n16526), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17574) );
  AND4_X1 U11289 ( .A1(n11299), .A2(n11298), .A3(n11297), .A4(n11296), .ZN(
        n11317) );
  AND4_X1 U11290 ( .A1(n11304), .A2(n11303), .A3(n11302), .A4(n11301), .ZN(
        n11316) );
  AND4_X1 U11291 ( .A1(n11282), .A2(n11281), .A3(n11280), .A4(n11279), .ZN(
        n11294) );
  AND4_X1 U11292 ( .A1(n10486), .A2(n10485), .A3(n10484), .A4(n10483), .ZN(
        n10487) );
  AND3_X1 U11293 ( .A1(n10517), .A2(n10516), .A3(n10430), .ZN(n10518) );
  AND2_X1 U11294 ( .A1(n10452), .A2(n10451), .ZN(n10456) );
  AND4_X1 U11295 ( .A1(n10479), .A2(n10478), .A3(n10477), .A4(n10476), .ZN(
        n10480) );
  AND4_X1 U11296 ( .A1(n11344), .A2(n11343), .A3(n11342), .A4(n11341), .ZN(
        n11360) );
  AND4_X1 U11297 ( .A1(n11356), .A2(n11355), .A3(n11354), .A4(n11353), .ZN(
        n11357) );
  AND4_X1 U11298 ( .A1(n11352), .A2(n11351), .A3(n11350), .A4(n11349), .ZN(
        n11358) );
  AND4_X1 U11299 ( .A1(n11277), .A2(n11276), .A3(n11275), .A4(n11274), .ZN(
        n11295) );
  AND4_X1 U11300 ( .A1(n11287), .A2(n11286), .A3(n11285), .A4(n11284), .ZN(
        n11293) );
  AND4_X1 U11301 ( .A1(n11348), .A2(n11347), .A3(n11346), .A4(n11345), .ZN(
        n11359) );
  AND4_X1 U11302 ( .A1(n11328), .A2(n11327), .A3(n11326), .A4(n11325), .ZN(
        n11339) );
  AND4_X1 U11303 ( .A1(n11336), .A2(n11335), .A3(n11334), .A4(n11333), .ZN(
        n11337) );
  AND4_X1 U11304 ( .A1(n11313), .A2(n11312), .A3(n11311), .A4(n11310), .ZN(
        n11314) );
  AND3_X1 U11305 ( .A1(n10454), .A2(n10453), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10455) );
  AND2_X1 U11306 ( .A1(n10446), .A2(n10430), .ZN(n10450) );
  AND4_X1 U11307 ( .A1(n11309), .A2(n11308), .A3(n11307), .A4(n11306), .ZN(
        n11315) );
  CLKBUF_X3 U11308 ( .A(n10154), .Z(n17157) );
  INV_X2 U11309 ( .A(n18094), .ZN(n9846) );
  CLKBUF_X1 U11310 ( .A(n13129), .Z(n13850) );
  INV_X2 U11311 ( .A(n16481), .ZN(n16483) );
  BUF_X4 U11312 ( .A(n10152), .Z(n9591) );
  INV_X2 U11313 ( .A(n10137), .ZN(n9593) );
  BUF_X4 U11315 ( .A(n10140), .Z(n9595) );
  INV_X1 U11316 ( .A(n12619), .ZN(n9641) );
  OR2_X1 U11317 ( .A1(n10101), .A2(n10103), .ZN(n10089) );
  OAI21_X1 U11318 ( .B1(n12670), .B2(n12669), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13129) );
  AND2_X2 U11319 ( .A1(n9989), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10670) );
  AND2_X1 U11320 ( .A1(n18627), .A2(n18210), .ZN(n18261) );
  NAND2_X1 U11321 ( .A1(n20789), .A2(n18784), .ZN(n10104) );
  INV_X2 U11322 ( .A(n15782), .ZN(n18612) );
  NAND2_X1 U11323 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18771), .ZN(
        n18633) );
  NAND2_X1 U11324 ( .A1(n18778), .A2(n18771), .ZN(n10101) );
  AND2_X2 U11325 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13153) );
  AND2_X2 U11326 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13564) );
  INV_X1 U11327 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11554) );
  BUF_X4 U11328 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n10596) );
  INV_X2 U11329 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n20789) );
  AND2_X1 U11330 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15782) );
  OR2_X2 U11331 ( .A1(n20124), .A2(n11408), .ZN(n9750) );
  NAND2_X1 U11332 ( .A1(n12138), .A2(n12137), .ZN(n12142) );
  INV_X1 U11333 ( .A(n15385), .ZN(n9596) );
  NAND2_X2 U11334 ( .A1(n9626), .A2(n11372), .ZN(n11399) );
  NOR2_X2 U11335 ( .A1(n17426), .A2(n17218), .ZN(n17214) );
  NOR4_X2 U11336 ( .A1(n17309), .A2(n17286), .A3(n20748), .A4(n17453), .ZN(
        n17199) );
  CLKBUF_X1 U11337 ( .A(n14096), .Z(n9597) );
  OAI21_X1 U11338 ( .B1(n15379), .B2(n15380), .A(n15331), .ZN(n9598) );
  OAI21_X1 U11339 ( .B1(n15379), .B2(n15380), .A(n15331), .ZN(n9599) );
  OAI21_X1 U11340 ( .B1(n15379), .B2(n15380), .A(n15331), .ZN(n15373) );
  OAI21_X4 U11341 ( .B1(n15389), .B2(n15388), .A(n15329), .ZN(n15379) );
  NOR2_X1 U11342 ( .A1(n10972), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14031) );
  NAND2_X1 U11343 ( .A1(n10976), .A2(n18937), .ZN(n10996) );
  OR2_X1 U11344 ( .A1(n10647), .A2(n10645), .ZN(n10624) );
  AND2_X1 U11345 ( .A1(n11233), .A2(n13590), .ZN(n11409) );
  AND3_X2 U11346 ( .A1(n11393), .A2(n11318), .A3(n11366), .ZN(n9771) );
  NOR2_X2 U11347 ( .A1(n13947), .A2(n13937), .ZN(n13936) );
  NOR2_X2 U11348 ( .A1(n13805), .A2(n13833), .ZN(n13834) );
  AND2_X2 U11349 ( .A1(n13415), .A2(n10059), .ZN(n13665) );
  INV_X1 U11350 ( .A(n14661), .ZN(n9601) );
  NAND2_X1 U11351 ( .A1(n9605), .A2(n9764), .ZN(n9602) );
  NAND3_X1 U11353 ( .A1(n9746), .A2(n10024), .A3(n9744), .ZN(n9604) );
  AND2_X1 U11354 ( .A1(n9811), .A2(n11461), .ZN(n9605) );
  NAND3_X1 U11355 ( .A1(n9746), .A2(n10024), .A3(n9744), .ZN(n14087) );
  NOR2_X4 U11356 ( .A1(n15283), .A2(n10914), .ZN(n15265) );
  INV_X1 U11357 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9989) );
  OR2_X2 U11358 ( .A1(n10585), .A2(n10574), .ZN(n9687) );
  OR2_X4 U11359 ( .A1(n11249), .A2(n11248), .ZN(n12070) );
  INV_X2 U11360 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11227) );
  NAND2_X1 U11361 ( .A1(n12803), .A2(n12806), .ZN(n12874) );
  XNOR2_X1 U11362 ( .A(n12803), .B(n11544), .ZN(n12866) );
  NAND2_X1 U11363 ( .A1(n13290), .A2(n12045), .ZN(n12909) );
  INV_X1 U11364 ( .A(n10790), .ZN(n9606) );
  OAI21_X1 U11365 ( .B1(n10020), .B2(n14746), .A(n9864), .ZN(n9863) );
  INV_X1 U11366 ( .A(n13502), .ZN(n9748) );
  NAND2_X2 U11367 ( .A1(n13540), .A2(n13539), .ZN(n13538) );
  NAND2_X1 U11369 ( .A1(n10594), .A2(n9611), .ZN(n9608) );
  AND2_X2 U11370 ( .A1(n9608), .A2(n9609), .ZN(n11113) );
  INV_X1 U11371 ( .A(n10607), .ZN(n9610) );
  AND2_X1 U11372 ( .A1(n10593), .A2(n10607), .ZN(n9611) );
  NAND2_X2 U11373 ( .A1(n13243), .A2(n10067), .ZN(n13371) );
  NOR2_X4 U11374 ( .A1(n13371), .A2(n12617), .ZN(n13415) );
  AND2_X1 U11375 ( .A1(n9638), .A2(n10430), .ZN(n13712) );
  NOR2_X2 U11377 ( .A1(n9759), .A2(n13610), .ZN(n14000) );
  NAND2_X1 U11378 ( .A1(n11365), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11389) );
  NOR2_X2 U11379 ( .A1(n14143), .A2(n14132), .ZN(n14527) );
  NOR2_X2 U11380 ( .A1(n14403), .A2(n14393), .ZN(n9912) );
  NOR2_X1 U11381 ( .A1(n10647), .A2(n10645), .ZN(n9613) );
  OAI211_X1 U11382 ( .C1(n10882), .C2(n10998), .A(n10881), .B(n10880), .ZN(
        n14094) );
  NAND2_X1 U11383 ( .A1(n10882), .A2(n10084), .ZN(n10881) );
  NAND2_X2 U11384 ( .A1(n11627), .A2(n11626), .ZN(n14013) );
  INV_X1 U11385 ( .A(n10554), .ZN(n9614) );
  INV_X1 U11386 ( .A(n9614), .ZN(n9615) );
  INV_X1 U11387 ( .A(n10550), .ZN(n10508) );
  NAND2_X1 U11388 ( .A1(n9757), .A2(n11721), .ZN(n14497) );
  NOR2_X2 U11389 ( .A1(n17743), .A2(n17747), .ZN(n17714) );
  INV_X1 U11391 ( .A(n10551), .ZN(n9618) );
  CLKBUF_X1 U11392 ( .A(n10565), .Z(n9628) );
  AND4_X1 U11393 ( .A1(n9687), .A2(n10579), .A3(n10578), .A4(n10577), .ZN(
        n10580) );
  NAND2_X2 U11394 ( .A1(n10674), .A2(n13699), .ZN(n12619) );
  INV_X1 U11395 ( .A(n9989), .ZN(n9619) );
  INV_X1 U11396 ( .A(n9619), .ZN(n9620) );
  NAND2_X1 U11397 ( .A1(n9824), .A2(n10537), .ZN(n10578) );
  INV_X1 U11398 ( .A(n10528), .ZN(n12678) );
  INV_X1 U11399 ( .A(n10585), .ZN(n15046) );
  OR2_X1 U11400 ( .A1(n14373), .A2(n9987), .ZN(n14361) );
  OR2_X1 U11401 ( .A1(n11389), .A2(n11463), .ZN(n11468) );
  NAND2_X2 U11402 ( .A1(n11389), .A2(n11385), .ZN(n11464) );
  NAND2_X1 U11403 ( .A1(n10563), .A2(n10562), .ZN(n10599) );
  INV_X2 U11404 ( .A(n10529), .ZN(n10548) );
  NAND2_X1 U11405 ( .A1(n10768), .A2(n10767), .ZN(n10788) );
  AOI211_X1 U11406 ( .C1(n13412), .C2(n19078), .A(n13873), .B(n13872), .ZN(
        n13874) );
  NAND2_X1 U11407 ( .A1(n13412), .A2(n10636), .ZN(n19571) );
  NAND2_X1 U11408 ( .A1(n13412), .A2(n10649), .ZN(n19487) );
  AND2_X1 U11409 ( .A1(n19103), .A2(n10529), .ZN(n10530) );
  NAND2_X1 U11410 ( .A1(n10433), .A2(n10432), .ZN(n10533) );
  NAND2_X2 U11411 ( .A1(n10531), .A2(n10534), .ZN(n10929) );
  INV_X2 U11412 ( .A(n14704), .ZN(n14717) );
  INV_X1 U11413 ( .A(n13208), .ZN(n13306) );
  NAND2_X1 U11414 ( .A1(n10535), .A2(n10534), .ZN(n13208) );
  NAND2_X1 U11415 ( .A1(n10563), .A2(n10562), .ZN(n9623) );
  NAND2_X1 U11416 ( .A1(n10563), .A2(n10562), .ZN(n9624) );
  INV_X1 U11417 ( .A(n12596), .ZN(n9625) );
  AND2_X1 U11418 ( .A1(n12429), .A2(n10671), .ZN(n12452) );
  AND2_X2 U11419 ( .A1(n10033), .A2(n10031), .ZN(n12894) );
  NAND2_X1 U11420 ( .A1(n11363), .A2(n12911), .ZN(n13032) );
  INV_X1 U11421 ( .A(n11367), .ZN(n9626) );
  NAND2_X4 U11422 ( .A1(n10445), .A2(n10444), .ZN(n10550) );
  NAND2_X4 U11423 ( .A1(n9675), .A2(n9648), .ZN(n12045) );
  AND4_X2 U11424 ( .A1(n11239), .A2(n11238), .A3(n11237), .A4(n11236), .ZN(
        n9648) );
  INV_X1 U11425 ( .A(n10546), .ZN(n10565) );
  INV_X2 U11426 ( .A(n9622), .ZN(n12685) );
  NAND2_X2 U11427 ( .A1(n10547), .A2(n10546), .ZN(n12658) );
  NAND2_X2 U11428 ( .A1(n15288), .A2(n15465), .ZN(n15283) );
  NAND2_X1 U11429 ( .A1(n11388), .A2(n11387), .ZN(n9796) );
  NOR2_X2 U11430 ( .A1(n10622), .A2(n13728), .ZN(n19526) );
  OAI21_X2 U11431 ( .B1(n15069), .B2(n15059), .A(n12607), .ZN(n15053) );
  XNOR2_X2 U11432 ( .A(n10620), .B(n9607), .ZN(n12146) );
  INV_X2 U11433 ( .A(n12045), .ZN(n11566) );
  OR2_X1 U11434 ( .A1(n10727), .A2(n10625), .ZN(n10626) );
  INV_X4 U11435 ( .A(n10523), .ZN(n10528) );
  OAI21_X2 U11437 ( .B1(n15396), .B2(n15327), .A(n15395), .ZN(n15389) );
  OAI21_X2 U11438 ( .B1(n15407), .B2(n15326), .A(n15405), .ZN(n15396) );
  NOR2_X4 U11439 ( .A1(n14181), .A2(n14192), .ZN(n14191) );
  AOI211_X2 U11440 ( .C1(n19078), .C2(n15595), .A(n15344), .B(n15343), .ZN(
        n15345) );
  AOI211_X2 U11441 ( .C1(n15605), .C2(n15604), .A(n15603), .B(n15602), .ZN(
        n15606) );
  NAND2_X2 U11443 ( .A1(n12150), .A2(n12149), .ZN(n12151) );
  NAND2_X2 U11444 ( .A1(n11566), .A2(n12070), .ZN(n11380) );
  NAND2_X1 U11445 ( .A1(n12813), .A2(n12812), .ZN(n12819) );
  NAND2_X2 U11446 ( .A1(n13819), .A2(n16300), .ZN(n13820) );
  NOR2_X2 U11447 ( .A1(n14683), .A2(n14682), .ZN(n14477) );
  XNOR2_X2 U11448 ( .A(n12827), .B(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13504) );
  OR2_X2 U11449 ( .A1(n13412), .A2(n10648), .ZN(n10800) );
  NAND2_X2 U11450 ( .A1(n9585), .A2(n20154), .ZN(n11586) );
  NAND3_X2 U11451 ( .A1(n9949), .A2(n10787), .A3(n13820), .ZN(n10882) );
  AOI21_X2 U11452 ( .B1(n12520), .B2(n10064), .A(n10063), .ZN(n12546) );
  XNOR2_X2 U11453 ( .A(n11438), .B(n11437), .ZN(n11568) );
  OAI21_X4 U11454 ( .B1(n13646), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11421), 
        .ZN(n12807) );
  NAND2_X4 U11455 ( .A1(n20064), .A2(n9750), .ZN(n13646) );
  AND2_X1 U11456 ( .A1(n11232), .A2(n13590), .ZN(n9631) );
  AND2_X1 U11457 ( .A1(n11232), .A2(n13590), .ZN(n9632) );
  NOR2_X4 U11458 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10671) );
  NAND3_X2 U11459 ( .A1(n9651), .A2(n9772), .A3(n9771), .ZN(n12048) );
  AND2_X1 U11460 ( .A1(n11232), .A2(n11235), .ZN(n9634) );
  AND2_X1 U11461 ( .A1(n11232), .A2(n11235), .ZN(n9635) );
  AND2_X1 U11462 ( .A1(n11232), .A2(n11235), .ZN(n11250) );
  AND2_X1 U11463 ( .A1(n11235), .A2(n13575), .ZN(n9636) );
  AND2_X2 U11464 ( .A1(n11235), .A2(n13575), .ZN(n9637) );
  AND2_X2 U11465 ( .A1(n10674), .A2(n10596), .ZN(n9638) );
  AND2_X1 U11466 ( .A1(n11232), .A2(n13590), .ZN(n9639) );
  AND2_X1 U11467 ( .A1(n11232), .A2(n13590), .ZN(n9640) );
  INV_X1 U11468 ( .A(n12587), .ZN(n9642) );
  BUF_X4 U11470 ( .A(n11255), .Z(n9644) );
  AND2_X4 U11471 ( .A1(n9763), .A2(n13575), .ZN(n11255) );
  NAND3_X2 U11472 ( .A1(n9814), .A2(n10007), .A3(n10006), .ZN(n14594) );
  OAI21_X2 U11473 ( .B1(n10722), .B2(n10721), .A(n10720), .ZN(n10723) );
  AOI21_X2 U11474 ( .B1(n9623), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n10570), .ZN(n10591) );
  XNOR2_X2 U11475 ( .A(n11565), .B(n11564), .ZN(n12818) );
  NAND2_X2 U11476 ( .A1(n14389), .A2(n11950), .ZN(n14373) );
  NOR2_X4 U11477 ( .A1(n14404), .A2(n14407), .ZN(n14389) );
  AND2_X1 U11478 ( .A1(n13564), .A2(n11234), .ZN(n9645) );
  XNOR2_X2 U11479 ( .A(n9646), .B(n9762), .ZN(n14586) );
  BUF_X1 U11480 ( .A(n14350), .Z(n9646) );
  AND2_X1 U11481 ( .A1(n12546), .A2(n10074), .ZN(n12547) );
  NAND2_X1 U11482 ( .A1(n19109), .A2(n10564), .ZN(n9825) );
  NAND2_X1 U11483 ( .A1(n13331), .A2(n10553), .ZN(n9826) );
  XNOR2_X1 U11484 ( .A(n10178), .B(n9841), .ZN(n10195) );
  INV_X1 U11485 ( .A(n10008), .ZN(n10007) );
  NAND2_X1 U11486 ( .A1(n14674), .A2(n14841), .ZN(n10006) );
  NAND2_X1 U11487 ( .A1(n12894), .A2(n9665), .ZN(n9814) );
  AOI21_X1 U11488 ( .B1(n10339), .B2(n10345), .A(n10344), .ZN(n18601) );
  NAND2_X1 U11489 ( .A1(n20024), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11491) );
  NOR2_X1 U11490 ( .A1(n10596), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12429) );
  AND2_X1 U11491 ( .A1(n12677), .A2(n19737), .ZN(n12683) );
  NAND2_X1 U11492 ( .A1(n9756), .A2(n9726), .ZN(n14484) );
  INV_X1 U11493 ( .A(n14497), .ZN(n9756) );
  INV_X1 U11494 ( .A(n15935), .ZN(n9972) );
  CLKBUF_X1 U11495 ( .A(n11574), .Z(n13621) );
  INV_X1 U11496 ( .A(n14311), .ZN(n9743) );
  NAND2_X1 U11497 ( .A1(n20048), .A2(n13033), .ZN(n9776) );
  NAND3_X1 U11498 ( .A1(n12917), .A2(n11372), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12071) );
  NAND2_X1 U11499 ( .A1(n9811), .A2(n11461), .ZN(n11551) );
  NAND2_X1 U11500 ( .A1(n11558), .A2(n11557), .ZN(n9811) );
  NAND2_X1 U11501 ( .A1(n9685), .A2(n12911), .ZN(n11319) );
  INV_X1 U11502 ( .A(n11376), .ZN(n11379) );
  NAND2_X1 U11503 ( .A1(n10066), .A2(n10065), .ZN(n10064) );
  AND2_X1 U11504 ( .A1(n12519), .A2(n15083), .ZN(n10063) );
  INV_X1 U11505 ( .A(n15083), .ZN(n10065) );
  AND2_X1 U11506 ( .A1(n19764), .A2(n10508), .ZN(n12517) );
  INV_X1 U11507 ( .A(n15118), .ZN(n10062) );
  OR2_X1 U11508 ( .A1(n9897), .A2(n13992), .ZN(n9896) );
  AND2_X1 U11509 ( .A1(n10901), .A2(n10900), .ZN(n10902) );
  NAND2_X1 U11510 ( .A1(n15309), .A2(n9681), .ZN(n9828) );
  INV_X1 U11511 ( .A(n11092), .ZN(n9829) );
  NOR2_X1 U11512 ( .A1(n10879), .A2(n10876), .ZN(n10874) );
  CLKBUF_X2 U11513 ( .A(n12705), .Z(n12795) );
  NAND2_X1 U11514 ( .A1(n10556), .A2(n10555), .ZN(n10557) );
  NAND2_X1 U11515 ( .A1(n10554), .A2(n10553), .ZN(n10555) );
  INV_X1 U11516 ( .A(n10647), .ZN(n9947) );
  NAND2_X1 U11517 ( .A1(n10657), .A2(n10647), .ZN(n10622) );
  OR2_X1 U11518 ( .A1(n18635), .A2(n10098), .ZN(n14284) );
  NOR2_X1 U11519 ( .A1(n10223), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10044) );
  NAND2_X1 U11520 ( .A1(n17721), .A2(n10048), .ZN(n17619) );
  AND2_X1 U11521 ( .A1(n10216), .A2(n17975), .ZN(n10048) );
  NOR2_X1 U11522 ( .A1(n14205), .A2(n14204), .ZN(n15780) );
  OR2_X1 U11523 ( .A1(n10103), .A2(n18635), .ZN(n9674) );
  AND2_X1 U11524 ( .A1(n20417), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12041) );
  NOR2_X1 U11525 ( .A1(n13599), .A2(n19780), .ZN(n13264) );
  AOI21_X1 U11526 ( .B1(n10037), .B2(n10034), .A(n10032), .ZN(n10031) );
  INV_X1 U11527 ( .A(n14688), .ZN(n10032) );
  OR2_X1 U11529 ( .A1(n11217), .A2(n14936), .ZN(n15237) );
  AND2_X1 U11530 ( .A1(n13416), .A2(n9655), .ZN(n10060) );
  AND2_X1 U11531 ( .A1(n9998), .A2(n15211), .ZN(n9997) );
  NAND2_X1 U11532 ( .A1(n9999), .A2(n10001), .ZN(n9998) );
  INV_X1 U11533 ( .A(n13348), .ZN(n13344) );
  XNOR2_X1 U11534 ( .A(n12142), .B(n12143), .ZN(n13192) );
  NAND2_X1 U11535 ( .A1(n13192), .A2(n13191), .ZN(n13194) );
  NOR2_X1 U11536 ( .A1(n10634), .A2(n10655), .ZN(n19089) );
  NAND2_X1 U11537 ( .A1(n10438), .A2(n10430), .ZN(n10445) );
  NAND2_X1 U11538 ( .A1(n10443), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10444) );
  AND2_X1 U11539 ( .A1(n19747), .A2(n10940), .ZN(n13687) );
  NOR2_X1 U11540 ( .A1(n10335), .A2(n10334), .ZN(n10345) );
  OAI21_X1 U11541 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n16821), .A(
        n10338), .ZN(n10344) );
  NAND2_X1 U11542 ( .A1(n10201), .A2(n17316), .ZN(n10176) );
  OR2_X1 U11543 ( .A1(n17781), .A2(n9650), .ZN(n9788) );
  OR2_X1 U11544 ( .A1(n15235), .A2(n16272), .ZN(n9956) );
  NAND2_X1 U11545 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n9804) );
  NAND2_X1 U11546 ( .A1(n12018), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n9803) );
  AOI22_X1 U11547 ( .A1(n10675), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10478) );
  NAND2_X1 U11548 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n9810) );
  NAND2_X1 U11549 ( .A1(n9643), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n9809) );
  CLKBUF_X1 U11550 ( .A(n11266), .Z(n11920) );
  NAND2_X1 U11551 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n9806) );
  NAND2_X1 U11552 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n9805) );
  NAND2_X1 U11553 ( .A1(n11378), .A2(n11398), .ZN(n9755) );
  NOR2_X1 U11554 ( .A1(n13290), .A2(n20417), .ZN(n11569) );
  OR2_X1 U11555 ( .A1(n11420), .A2(n11419), .ZN(n12809) );
  NOR2_X1 U11556 ( .A1(n11368), .A2(n11372), .ZN(n13038) );
  AND4_X1 U11557 ( .A1(n10739), .A2(n10738), .A3(n10737), .A4(n10736), .ZN(
        n10740) );
  NOR2_X1 U11558 ( .A1(n12070), .A2(n11376), .ZN(n12047) );
  NAND2_X1 U11559 ( .A1(n14875), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12011) );
  INV_X1 U11560 ( .A(n14444), .ZN(n9757) );
  INV_X1 U11561 ( .A(n14013), .ZN(n9976) );
  AND2_X1 U11562 ( .A1(n9800), .A2(n9799), .ZN(n11614) );
  NAND2_X1 U11563 ( .A1(n11517), .A2(n9862), .ZN(n11603) );
  INV_X1 U11564 ( .A(n11569), .ZN(n11905) );
  INV_X1 U11565 ( .A(n11574), .ZN(n12014) );
  NOR2_X1 U11566 ( .A1(n9926), .A2(n14472), .ZN(n9925) );
  INV_X1 U11567 ( .A(n9927), .ZN(n9926) );
  NOR2_X1 U11568 ( .A1(n9929), .A2(n9928), .ZN(n9927) );
  INV_X1 U11569 ( .A(n14480), .ZN(n9928) );
  INV_X1 U11570 ( .A(n14824), .ZN(n9929) );
  INV_X1 U11571 ( .A(n12862), .ZN(n10029) );
  AND2_X1 U11572 ( .A1(n12855), .A2(n12865), .ZN(n9861) );
  INV_X1 U11573 ( .A(n13682), .ZN(n9919) );
  AND2_X1 U11574 ( .A1(n13053), .A2(n13045), .ZN(n13399) );
  OAI21_X1 U11575 ( .B1(n20671), .B2(n16168), .A(n20633), .ZN(n20023) );
  OR2_X1 U11576 ( .A1(n13589), .A2(n13588), .ZN(n15832) );
  NOR2_X1 U11577 ( .A1(n11049), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11038) );
  NAND2_X1 U11578 ( .A1(n11054), .A2(n9876), .ZN(n11059) );
  INV_X1 U11579 ( .A(n12343), .ZN(n12453) );
  NAND2_X1 U11580 ( .A1(n10583), .A2(n10571), .ZN(n9821) );
  NAND2_X1 U11581 ( .A1(n10573), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9822) );
  INV_X1 U11582 ( .A(n13195), .ZN(n9824) );
  INV_X1 U11583 ( .A(n15146), .ZN(n9891) );
  AND2_X1 U11584 ( .A1(n9659), .A2(n14050), .ZN(n10069) );
  INV_X1 U11585 ( .A(n15695), .ZN(n12761) );
  INV_X1 U11586 ( .A(n15213), .ZN(n9840) );
  INV_X1 U11587 ( .A(n9839), .ZN(n9838) );
  OAI21_X1 U11588 ( .B1(n9997), .B2(n9840), .A(n15232), .ZN(n9839) );
  NOR2_X1 U11589 ( .A1(n15282), .A2(n9910), .ZN(n9909) );
  INV_X1 U11590 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n9910) );
  NAND2_X1 U11591 ( .A1(n10561), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10562) );
  AND2_X1 U11592 ( .A1(n15075), .A2(n14959), .ZN(n9968) );
  INV_X1 U11593 ( .A(n14178), .ZN(n9964) );
  INV_X1 U11594 ( .A(n13667), .ZN(n9960) );
  INV_X1 U11595 ( .A(n10003), .ZN(n9832) );
  AND2_X1 U11596 ( .A1(n10004), .A2(n16246), .ZN(n10003) );
  INV_X1 U11597 ( .A(n15220), .ZN(n15240) );
  INV_X1 U11598 ( .A(n15046), .ZN(n11204) );
  INV_X1 U11599 ( .A(n14031), .ZN(n9949) );
  OR2_X1 U11600 ( .A1(n10782), .A2(n10781), .ZN(n12721) );
  NAND2_X1 U11601 ( .A1(n13842), .A2(n10753), .ZN(n13317) );
  OR2_X1 U11602 ( .A1(n10647), .A2(n12141), .ZN(n10655) );
  NOR2_X1 U11603 ( .A1(n10647), .A2(n13728), .ZN(n10654) );
  AOI22_X1 U11604 ( .A1(n9630), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10510) );
  NAND2_X1 U11605 ( .A1(n20827), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10937) );
  AND2_X1 U11606 ( .A1(n10131), .A2(n10053), .ZN(n10052) );
  NAND2_X1 U11607 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10051) );
  INV_X1 U11608 ( .A(n10132), .ZN(n10054) );
  OR2_X1 U11609 ( .A1(n10102), .A2(n18612), .ZN(n16983) );
  NOR2_X1 U11610 ( .A1(n18633), .A2(n10104), .ZN(n10154) );
  NOR2_X1 U11611 ( .A1(n9942), .A2(n17472), .ZN(n9941) );
  INV_X1 U11612 ( .A(n9943), .ZN(n9942) );
  AND3_X1 U11613 ( .A1(n17712), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17673) );
  NOR2_X1 U11614 ( .A1(n17320), .A2(n10177), .ZN(n10201) );
  NOR2_X1 U11615 ( .A1(n17619), .A2(n16341), .ZN(n10218) );
  NAND2_X1 U11616 ( .A1(n10212), .A2(n10223), .ZN(n10217) );
  NAND2_X1 U11617 ( .A1(n10211), .A2(n10210), .ZN(n10212) );
  NAND2_X1 U11618 ( .A1(n10217), .A2(n9843), .ZN(n9842) );
  INV_X1 U11619 ( .A(n10218), .ZN(n9843) );
  NAND2_X1 U11620 ( .A1(n17767), .A2(n10196), .ZN(n10199) );
  NAND2_X1 U11621 ( .A1(n17339), .A2(n10353), .ZN(n10179) );
  INV_X1 U11622 ( .A(n18191), .ZN(n10319) );
  NAND2_X1 U11623 ( .A1(n18191), .A2(n10382), .ZN(n10394) );
  NOR2_X1 U11624 ( .A1(n13047), .A2(n13048), .ZN(n13563) );
  OR2_X1 U11625 ( .A1(n20667), .A2(n13623), .ZN(n19831) );
  AND2_X1 U11626 ( .A1(n19831), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13639) );
  OR2_X1 U11627 ( .A1(n12048), .A2(n12906), .ZN(n13546) );
  INV_X2 U11628 ( .A(n11905), .ZN(n12042) );
  NAND2_X1 U11629 ( .A1(n14360), .A2(n9988), .ZN(n9987) );
  INV_X1 U11630 ( .A(n14375), .ZN(n9988) );
  INV_X1 U11631 ( .A(n14391), .ZN(n11950) );
  NAND2_X1 U11632 ( .A1(n11911), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11951) );
  CLKBUF_X1 U11633 ( .A(n14497), .Z(n14498) );
  AOI21_X1 U11634 ( .B1(n11556), .B2(n9971), .A(n9970), .ZN(n9969) );
  INV_X1 U11635 ( .A(n11578), .ZN(n9970) );
  NAND2_X1 U11636 ( .A1(n14362), .A2(n13026), .ZN(n14327) );
  NAND2_X1 U11637 ( .A1(n10022), .A2(n10018), .ZN(n10017) );
  AND2_X1 U11638 ( .A1(n10021), .A2(n14750), .ZN(n10018) );
  NAND2_X1 U11639 ( .A1(n9912), .A2(n9911), .ZN(n14378) );
  INV_X1 U11640 ( .A(n14376), .ZN(n9911) );
  NAND2_X1 U11641 ( .A1(n10005), .A2(n14841), .ZN(n14652) );
  OR2_X1 U11642 ( .A1(n14674), .A2(n10010), .ZN(n10005) );
  INV_X1 U11643 ( .A(n12889), .ZN(n10036) );
  NOR2_X1 U11644 ( .A1(n10037), .A2(n14842), .ZN(n9865) );
  NAND2_X1 U11645 ( .A1(n14503), .A2(n9706), .ZN(n14834) );
  INV_X1 U11646 ( .A(n14487), .ZN(n9921) );
  NAND2_X1 U11647 ( .A1(n14503), .A2(n9922), .ZN(n14857) );
  NAND2_X1 U11648 ( .A1(n14503), .A2(n14493), .ZN(n14859) );
  AND2_X1 U11649 ( .A1(n13053), .A2(n14877), .ZN(n13403) );
  NOR2_X1 U11650 ( .A1(n9774), .A2(n11368), .ZN(n9773) );
  AND2_X1 U11651 ( .A1(n15843), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n14301) );
  INV_X1 U11652 ( .A(n20127), .ZN(n20122) );
  OR2_X1 U11653 ( .A1(n13601), .A2(n20383), .ZN(n20156) );
  AND2_X1 U11654 ( .A1(n20330), .A2(n20162), .ZN(n20450) );
  AND2_X1 U11655 ( .A1(n12113), .A2(n12112), .ZN(n13599) );
  AND2_X1 U11656 ( .A1(n20555), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15843) );
  AND2_X1 U11657 ( .A1(n13685), .A2(n13687), .ZN(n13694) );
  AND2_X1 U11658 ( .A1(n12655), .A2(n12656), .ZN(n13705) );
  AND2_X1 U11659 ( .A1(n10956), .A2(n10952), .ZN(n12648) );
  NOR2_X1 U11660 ( .A1(n11045), .A2(n9877), .ZN(n9875) );
  NOR2_X1 U11661 ( .A1(n13842), .A2(n13706), .ZN(n13218) );
  XOR2_X1 U11662 ( .A(n12609), .B(n12608), .Z(n15054) );
  NOR2_X1 U11663 ( .A1(n12569), .A2(n12570), .ZN(n15059) );
  NOR2_X1 U11664 ( .A1(n14962), .A2(n9893), .ZN(n9892) );
  INV_X1 U11665 ( .A(n14980), .ZN(n9893) );
  AOI21_X1 U11666 ( .B1(n15085), .B2(n15088), .A(n12499), .ZN(n12520) );
  INV_X1 U11667 ( .A(n15105), .ZN(n10061) );
  AND2_X1 U11668 ( .A1(n12778), .A2(n12777), .ZN(n14994) );
  AND3_X1 U11669 ( .A1(n12765), .A2(n12764), .A3(n12763), .ZN(n15033) );
  AND3_X1 U11670 ( .A1(n12752), .A2(n12751), .A3(n12750), .ZN(n13937) );
  INV_X1 U11671 ( .A(n9896), .ZN(n9895) );
  AOI22_X1 U11672 ( .A1(n13842), .A2(n13705), .B1(n13694), .B2(n13695), .ZN(
        n13220) );
  AND2_X1 U11673 ( .A1(n19014), .A2(n12661), .ZN(n13515) );
  NOR2_X1 U11674 ( .A1(n15237), .A2(n15236), .ZN(n13768) );
  AND3_X1 U11675 ( .A1(n10892), .A2(n10891), .A3(n10890), .ZN(n10904) );
  AND4_X1 U11676 ( .A1(n10898), .A2(n10897), .A3(n10896), .A4(n10895), .ZN(
        n10903) );
  AND4_X1 U11677 ( .A1(n10889), .A2(n10888), .A3(n10887), .A4(n10886), .ZN(
        n10905) );
  NAND2_X1 U11678 ( .A1(n9996), .A2(n9838), .ZN(n9836) );
  AOI21_X1 U11679 ( .B1(n9838), .B2(n9840), .A(n9835), .ZN(n9834) );
  INV_X1 U11680 ( .A(n15233), .ZN(n9835) );
  INV_X1 U11681 ( .A(n9993), .ZN(n9992) );
  INV_X1 U11682 ( .A(n9991), .ZN(n9994) );
  OAI21_X1 U11683 ( .B1(n11082), .B2(n9995), .A(n15315), .ZN(n9993) );
  NOR2_X2 U11684 ( .A1(n14899), .A2(n15409), .ZN(n14901) );
  CLKBUF_X1 U11685 ( .A(n14899), .Z(n14900) );
  INV_X1 U11686 ( .A(n15019), .ZN(n9901) );
  OAI21_X1 U11687 ( .B1(n14157), .B2(n9952), .A(n9950), .ZN(n15441) );
  NAND2_X1 U11688 ( .A1(n14158), .A2(n9951), .ZN(n9950) );
  NOR2_X1 U11689 ( .A1(n14158), .A2(n9951), .ZN(n9952) );
  AND2_X1 U11690 ( .A1(n9958), .A2(n9678), .ZN(n13251) );
  XNOR2_X1 U11691 ( .A(n11116), .B(n11114), .ZN(n11117) );
  NOR2_X1 U11692 ( .A1(n13348), .A2(n10929), .ZN(n13349) );
  AND2_X1 U11693 ( .A1(n19762), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12156) );
  NAND2_X1 U11694 ( .A1(n12135), .A2(n19737), .ZN(n12161) );
  OR2_X1 U11695 ( .A1(n12142), .A2(n12144), .ZN(n12145) );
  NOR2_X2 U11696 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19520) );
  OR2_X1 U11697 ( .A1(n19721), .A2(n14073), .ZN(n19493) );
  OR2_X1 U11698 ( .A1(n19721), .A2(n19732), .ZN(n19568) );
  NAND2_X1 U11699 ( .A1(n13844), .A2(n13843), .ZN(n13845) );
  NAND2_X1 U11700 ( .A1(n10425), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10433) );
  OR2_X1 U11701 ( .A1(n16585), .A2(n16837), .ZN(n9946) );
  OR2_X1 U11702 ( .A1(n10394), .A2(n14208), .ZN(n17397) );
  INV_X1 U11703 ( .A(n18652), .ZN(n17399) );
  NAND2_X1 U11704 ( .A1(n17538), .A2(n9933), .ZN(n9932) );
  NOR2_X1 U11705 ( .A1(n9935), .A2(n9934), .ZN(n9933) );
  INV_X1 U11706 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n9934) );
  NOR2_X1 U11707 ( .A1(n9663), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9794) );
  NAND2_X1 U11708 ( .A1(n17477), .A2(n10225), .ZN(n15795) );
  AND2_X1 U11709 ( .A1(n17722), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10225) );
  OAI21_X1 U11710 ( .B1(n17465), .B2(n9854), .A(n16375), .ZN(n9853) );
  NAND2_X1 U11711 ( .A1(n9850), .A2(n16376), .ZN(n9849) );
  OR2_X1 U11712 ( .A1(n16377), .A2(n18794), .ZN(n9850) );
  NOR2_X1 U11713 ( .A1(n9852), .A2(n18796), .ZN(n9851) );
  NOR2_X1 U11714 ( .A1(n16374), .A2(n16375), .ZN(n9852) );
  NAND2_X1 U11715 ( .A1(n10045), .A2(n17521), .ZN(n10224) );
  INV_X1 U11716 ( .A(n10044), .ZN(n10039) );
  OAI211_X1 U11717 ( .C1(n17521), .C2(n17845), .A(n10041), .B(n10040), .ZN(
        n17492) );
  AOI21_X1 U11718 ( .B1(n10038), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n9658), .ZN(n10041) );
  INV_X1 U11719 ( .A(n17722), .ZN(n10223) );
  NOR2_X1 U11720 ( .A1(n17722), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9859) );
  NOR2_X1 U11721 ( .A1(n9786), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9785) );
  INV_X1 U11722 ( .A(n10207), .ZN(n9786) );
  NAND2_X1 U11723 ( .A1(n17728), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17727) );
  NAND2_X1 U11724 ( .A1(n10194), .A2(n17791), .ZN(n17781) );
  NAND3_X1 U11725 ( .A1(n10254), .A2(n10253), .A3(n10252), .ZN(n18172) );
  NOR2_X1 U11726 ( .A1(n15780), .A2(n15779), .ZN(n18626) );
  NOR2_X1 U11727 ( .A1(n10395), .A2(n10394), .ZN(n18652) );
  NAND2_X1 U11728 ( .A1(n14571), .A2(n12130), .ZN(n16015) );
  INV_X2 U11729 ( .A(n14571), .ZN(n16008) );
  OR2_X1 U11730 ( .A1(n19968), .A2(n13267), .ZN(n14723) );
  AND2_X1 U11731 ( .A1(n14723), .A2(n13300), .ZN(n16032) );
  INV_X1 U11732 ( .A(n19968), .ZN(n16035) );
  INV_X1 U11733 ( .A(n19981), .ZN(n20017) );
  NAND2_X1 U11734 ( .A1(n13053), .A2(n12920), .ZN(n16126) );
  NAND2_X1 U11735 ( .A1(n20268), .A2(n20155), .ZN(n20639) );
  AND2_X1 U11736 ( .A1(n13694), .A2(n13318), .ZN(n19758) );
  OR2_X1 U11737 ( .A1(n10931), .A2(n10930), .ZN(n10933) );
  NAND2_X1 U11738 ( .A1(n15029), .A2(n18893), .ZN(n18888) );
  AND2_X1 U11739 ( .A1(n9698), .A2(n9661), .ZN(n10059) );
  NAND2_X1 U11740 ( .A1(n10617), .A2(n10616), .ZN(n10618) );
  OR2_X1 U11741 ( .A1(n14934), .A2(n12798), .ZN(n12799) );
  AOI21_X2 U11742 ( .B1(n13220), .B2(n13336), .A(n18832), .ZN(n19014) );
  INV_X1 U11743 ( .A(n19072), .ZN(n16250) );
  AND2_X1 U11744 ( .A1(n19067), .A2(n11211), .ZN(n19078) );
  OR2_X1 U11745 ( .A1(n18834), .A2(n10753), .ZN(n19075) );
  NAND2_X1 U11746 ( .A1(n15485), .A2(n15484), .ZN(n15486) );
  NAND2_X1 U11747 ( .A1(n9837), .A2(n15213), .ZN(n15231) );
  XNOR2_X1 U11748 ( .A(n15230), .B(n15480), .ZN(n15492) );
  NAND2_X1 U11749 ( .A1(n13344), .A2(n13323), .ZN(n16315) );
  INV_X1 U11750 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20827) );
  OR2_X1 U11751 ( .A1(n12142), .A2(n13202), .ZN(n19739) );
  INV_X1 U11752 ( .A(n19520), .ZN(n19714) );
  CLKBUF_X1 U11753 ( .A(n10538), .Z(n10753) );
  NOR2_X1 U11754 ( .A1(n18602), .A2(n17398), .ZN(n18823) );
  XNOR2_X1 U11755 ( .A(n16543), .B(n9939), .ZN(n9938) );
  INV_X1 U11756 ( .A(n16544), .ZN(n9939) );
  INV_X1 U11757 ( .A(n16845), .ZN(n16874) );
  INV_X1 U11758 ( .A(n18204), .ZN(n17120) );
  NOR3_X1 U11759 ( .A1(n18204), .A2(n17275), .A3(n17243), .ZN(n17263) );
  NOR2_X1 U11760 ( .A1(n10110), .A2(n10109), .ZN(n17312) );
  NOR2_X1 U11761 ( .A1(n10130), .A2(n10129), .ZN(n17328) );
  NOR2_X1 U11762 ( .A1(n16335), .A2(n16334), .ZN(n16336) );
  INV_X2 U11763 ( .A(n17663), .ZN(n17609) );
  NOR2_X2 U11764 ( .A1(n17312), .A2(n17815), .ZN(n17723) );
  NOR2_X2 U11765 ( .A1(n18804), .A2(n16494), .ZN(n17803) );
  INV_X1 U11766 ( .A(n17803), .ZN(n17816) );
  AOI21_X1 U11767 ( .B1(n16333), .B2(n18058), .A(n10416), .ZN(n10417) );
  XNOR2_X1 U11768 ( .A(n10057), .B(n16343), .ZN(n16349) );
  NAND2_X1 U11769 ( .A1(n9791), .A2(n10058), .ZN(n10057) );
  INV_X1 U11770 ( .A(n15851), .ZN(n10058) );
  INV_X1 U11771 ( .A(n18142), .ZN(n18125) );
  NOR2_X1 U11772 ( .A1(n18794), .A2(n18143), .ZN(n18142) );
  INV_X1 U11773 ( .A(n16839), .ZN(n18661) );
  NOR2_X1 U11774 ( .A1(n10735), .A2(n10734), .ZN(n10739) );
  AND2_X1 U11775 ( .A1(n9802), .A2(n9801), .ZN(n11798) );
  NAND2_X1 U11776 ( .A1(n9643), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n9802) );
  NAND2_X1 U11777 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n9801) );
  AND2_X1 U11778 ( .A1(n9804), .A2(n9803), .ZN(n11631) );
  NAND2_X1 U11779 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n9799) );
  NAND2_X1 U11780 ( .A1(n12018), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n9800) );
  AND2_X1 U11781 ( .A1(n11585), .A2(n11595), .ZN(n9862) );
  OR2_X1 U11782 ( .A1(n11514), .A2(n11513), .ZN(n12846) );
  INV_X1 U11783 ( .A(n12823), .ZN(n12830) );
  NOR2_X1 U11784 ( .A1(n11371), .A2(n11372), .ZN(n11363) );
  AOI22_X1 U11785 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11688), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11230) );
  AND2_X1 U11786 ( .A1(n11007), .A2(n10999), .ZN(n9874) );
  INV_X1 U11787 ( .A(n12519), .ZN(n10066) );
  OR2_X1 U11788 ( .A1(n10752), .A2(n10751), .ZN(n12715) );
  NAND4_X1 U11789 ( .A1(n12685), .A2(n10550), .A3(n10529), .A4(n10528), .ZN(
        n10564) );
  NAND2_X1 U11790 ( .A1(n10508), .A2(n10523), .ZN(n10554) );
  AOI22_X1 U11791 ( .A1(n10675), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10446) );
  NOR2_X1 U11792 ( .A1(n10086), .A2(n10490), .ZN(n10494) );
  NAND2_X1 U11793 ( .A1(n10489), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10490) );
  AND3_X1 U11794 ( .A1(n13216), .A2(n13215), .A3(n13332), .ZN(n13312) );
  NAND2_X1 U11795 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10053) );
  INV_X1 U11796 ( .A(n10400), .ZN(n10381) );
  NOR2_X1 U11797 ( .A1(n10384), .A2(n10381), .ZN(n10382) );
  OR2_X1 U11798 ( .A1(n11380), .A2(n11366), .ZN(n13048) );
  AOI22_X1 U11799 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11266), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11245) );
  NAND2_X1 U11800 ( .A1(n11361), .A2(n13290), .ZN(n12068) );
  NAND2_X1 U11801 ( .A1(n14478), .A2(n9705), .ZN(n14404) );
  NOR2_X1 U11802 ( .A1(n14431), .A2(n9983), .ZN(n9982) );
  INV_X1 U11803 ( .A(n9984), .ZN(n9983) );
  NOR2_X1 U11804 ( .A1(n14470), .A2(n14668), .ZN(n9984) );
  AOI22_X1 U11805 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11828) );
  AOI21_X1 U11806 ( .B1(n9632), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A(n9733), .ZN(n11814) );
  AND2_X1 U11807 ( .A1(n9810), .A2(n9809), .ZN(n11774) );
  AND2_X1 U11808 ( .A1(n9808), .A2(n9807), .ZN(n11762) );
  NAND2_X1 U11809 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n9807) );
  NAND2_X1 U11810 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n9808) );
  INV_X1 U11811 ( .A(n12011), .ZN(n12037) );
  NAND2_X1 U11812 ( .A1(n11739), .A2(n9975), .ZN(n9974) );
  INV_X1 U11813 ( .A(n14492), .ZN(n9975) );
  NOR2_X1 U11814 ( .A1(n9981), .A2(n9980), .ZN(n9979) );
  INV_X1 U11815 ( .A(n14442), .ZN(n9980) );
  NOR2_X1 U11816 ( .A1(n9981), .A2(n9978), .ZN(n9977) );
  AND2_X1 U11817 ( .A1(n9798), .A2(n9797), .ZN(n11663) );
  NAND2_X1 U11818 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n9798) );
  NAND2_X1 U11819 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n9797) );
  AND2_X1 U11820 ( .A1(n9806), .A2(n9805), .ZN(n11651) );
  NAND2_X1 U11821 ( .A1(n11642), .A2(n14129), .ZN(n9981) );
  XNOR2_X1 U11822 ( .A(n9766), .B(n9765), .ZN(n12845) );
  INV_X1 U11823 ( .A(n11595), .ZN(n9765) );
  INV_X1 U11824 ( .A(n11585), .ZN(n9767) );
  NAND2_X1 U11825 ( .A1(n12067), .A2(n9754), .ZN(n13166) );
  OAI21_X1 U11826 ( .B1(n14844), .B2(n14653), .A(n10009), .ZN(n10008) );
  NAND2_X1 U11827 ( .A1(n14841), .A2(n10010), .ZN(n10009) );
  NAND2_X1 U11828 ( .A1(n12896), .A2(n15867), .ZN(n10010) );
  NOR2_X1 U11829 ( .A1(n14860), .A2(n9923), .ZN(n9922) );
  INV_X1 U11830 ( .A(n14493), .ZN(n9923) );
  NAND2_X1 U11831 ( .A1(n14717), .A2(n12888), .ZN(n14693) );
  INV_X1 U11832 ( .A(n12854), .ZN(n9745) );
  INV_X1 U11833 ( .A(n12864), .ZN(n10025) );
  INV_X1 U11834 ( .A(n16044), .ZN(n10028) );
  NOR2_X1 U11835 ( .A1(n20024), .A2(n9769), .ZN(n9768) );
  AND3_X1 U11836 ( .A1(n11440), .A2(n11435), .A3(n11434), .ZN(n11459) );
  OR2_X1 U11837 ( .A1(n11502), .A2(n11501), .ZN(n12847) );
  INV_X1 U11838 ( .A(n12071), .ZN(n12105) );
  NAND2_X1 U11839 ( .A1(n11255), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11341) );
  NAND2_X1 U11840 ( .A1(n11364), .A2(n11366), .ZN(n13565) );
  INV_X1 U11841 ( .A(n13032), .ZN(n11364) );
  NAND2_X1 U11842 ( .A1(n13035), .A2(n9753), .ZN(n13040) );
  NAND2_X1 U11843 ( .A1(n11369), .A2(n9772), .ZN(n13570) );
  AND2_X1 U11844 ( .A1(n13560), .A2(n13559), .ZN(n13592) );
  INV_X1 U11845 ( .A(n12818), .ZN(n20383) );
  NAND2_X1 U11846 ( .A1(n11491), .A2(n11490), .ZN(n12092) );
  AND2_X1 U11847 ( .A1(n12057), .A2(n12056), .ZN(n12072) );
  OR2_X1 U11848 ( .A1(n12058), .A2(n12055), .ZN(n12057) );
  NOR2_X1 U11849 ( .A1(n12671), .A2(n10550), .ZN(n10535) );
  OR2_X1 U11850 ( .A1(n14949), .A2(n11109), .ZN(n10968) );
  AND2_X1 U11851 ( .A1(n15090), .A2(n9879), .ZN(n9878) );
  AND2_X1 U11852 ( .A1(n11054), .A2(n10964), .ZN(n11062) );
  NOR2_X1 U11853 ( .A1(n9869), .A2(n9870), .ZN(n11019) );
  NAND2_X1 U11854 ( .A1(n9872), .A2(n9871), .ZN(n9870) );
  OR2_X1 U11855 ( .A1(n11005), .A2(n15217), .ZN(n11094) );
  AND2_X1 U11856 ( .A1(n9874), .A2(n11004), .ZN(n9872) );
  NAND2_X1 U11857 ( .A1(n11000), .A2(n9874), .ZN(n11005) );
  NOR2_X1 U11858 ( .A1(n9869), .A2(n9873), .ZN(n11009) );
  INV_X1 U11859 ( .A(n10999), .ZN(n9873) );
  AND2_X1 U11860 ( .A1(n10982), .A2(n10953), .ZN(n10993) );
  NAND2_X1 U11861 ( .A1(n10610), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10569) );
  NAND2_X1 U11862 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10678), .ZN(
        n12343) );
  INV_X1 U11863 ( .A(n10547), .ZN(n10539) );
  INV_X1 U11864 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15236) );
  AOI21_X1 U11865 ( .B1(n11082), .B2(n11083), .A(n9995), .ZN(n9991) );
  NAND2_X1 U11866 ( .A1(n14895), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14896) );
  NOR2_X1 U11867 ( .A1(n14896), .A2(n11216), .ZN(n14911) );
  AND2_X1 U11868 ( .A1(n9963), .A2(n9962), .ZN(n9961) );
  INV_X1 U11869 ( .A(n14988), .ZN(n9962) );
  AND2_X1 U11870 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11215) );
  NOR2_X1 U11871 ( .A1(n9649), .A2(n9906), .ZN(n9905) );
  NOR2_X1 U11872 ( .A1(n14106), .A2(n9908), .ZN(n9907) );
  NAND2_X1 U11873 ( .A1(n13153), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13772) );
  AOI22_X1 U11874 ( .A1(n13320), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n13749), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10544) );
  NOR2_X1 U11875 ( .A1(n14187), .A2(n14196), .ZN(n11171) );
  AND2_X1 U11876 ( .A1(n12761), .A2(n9900), .ZN(n9899) );
  INV_X1 U11877 ( .A(n15033), .ZN(n9900) );
  INV_X1 U11878 ( .A(n14058), .ZN(n9965) );
  NOR2_X1 U11879 ( .A1(n16275), .A2(n11029), .ZN(n9953) );
  OR2_X1 U11880 ( .A1(n13918), .A2(n9898), .ZN(n9897) );
  INV_X1 U11881 ( .A(n16288), .ZN(n9898) );
  AND2_X1 U11882 ( .A1(n15220), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11006) );
  NAND2_X1 U11883 ( .A1(n14096), .A2(n14097), .ZN(n9990) );
  AND2_X1 U11884 ( .A1(n10830), .A2(n10072), .ZN(n12725) );
  AOI21_X1 U11885 ( .B1(n10599), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n10603), .ZN(n10605) );
  AOI21_X1 U11886 ( .B1(n10599), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10613), .ZN(n11114) );
  AND2_X1 U11887 ( .A1(n10719), .A2(n10087), .ZN(n12703) );
  NAND2_X1 U11888 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12152) );
  NAND2_X1 U11889 ( .A1(n10482), .A2(n10481), .ZN(n10549) );
  NAND2_X1 U11890 ( .A1(n10079), .A2(n10083), .ZN(n10482) );
  NAND2_X1 U11891 ( .A1(n10480), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10481) );
  NAND2_X1 U11892 ( .A1(n19728), .A2(n19573), .ZN(n13851) );
  NAND2_X1 U11893 ( .A1(n18784), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10098) );
  NAND2_X1 U11894 ( .A1(n9844), .A2(n15782), .ZN(n17155) );
  NOR2_X1 U11895 ( .A1(n20789), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9844) );
  NAND2_X1 U11896 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20789), .ZN(
        n10102) );
  NOR2_X1 U11897 ( .A1(n10101), .A2(n10098), .ZN(n10093) );
  NOR2_X1 U11898 ( .A1(n17804), .A2(n9944), .ZN(n9943) );
  NOR2_X1 U11899 ( .A1(n17120), .A2(n18179), .ZN(n10400) );
  NAND2_X1 U11900 ( .A1(n17738), .A2(n10203), .ZN(n10206) );
  INV_X1 U11901 ( .A(n17339), .ZN(n10352) );
  NAND2_X1 U11902 ( .A1(n17397), .A2(n15783), .ZN(n15776) );
  NAND2_X1 U11903 ( .A1(n10396), .A2(n17399), .ZN(n15775) );
  AOI21_X1 U11904 ( .B1(n18147), .B2(n18807), .A(n18779), .ZN(n18159) );
  CLKBUF_X1 U11905 ( .A(n13028), .Z(n13029) );
  NOR2_X1 U11906 ( .A1(n11654), .A2(n19809), .ZN(n11658) );
  NAND2_X1 U11907 ( .A1(n13639), .A2(n13638), .ZN(n19835) );
  AND2_X1 U11908 ( .A1(n12990), .A2(n12923), .ZN(n12924) );
  INV_X1 U11909 ( .A(n20020), .ZN(n20021) );
  INV_X1 U11910 ( .A(n13394), .ZN(n19944) );
  NAND2_X1 U11911 ( .A1(n9986), .A2(n14320), .ZN(n9985) );
  INV_X1 U11912 ( .A(n14351), .ZN(n9986) );
  NOR2_X1 U11913 ( .A1(n11989), .A2(n14602), .ZN(n11990) );
  NAND2_X1 U11914 ( .A1(n11990), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13624) );
  OR2_X1 U11915 ( .A1(n11951), .A2(n14621), .ZN(n11952) );
  OR2_X1 U11916 ( .A1(n14630), .A2(n12014), .ZN(n11932) );
  AND2_X1 U11917 ( .A1(n11859), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11860) );
  NOR2_X1 U11918 ( .A1(n11822), .A2(n15903), .ZN(n11823) );
  NAND2_X1 U11919 ( .A1(n11790), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11822) );
  INV_X1 U11920 ( .A(n14484), .ZN(n11788) );
  OR2_X1 U11921 ( .A1(n11771), .A2(n15933), .ZN(n11789) );
  INV_X1 U11922 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15933) );
  CLKBUF_X1 U11923 ( .A(n14484), .Z(n14485) );
  AND2_X1 U11924 ( .A1(n11722), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11740) );
  INV_X1 U11925 ( .A(n14497), .ZN(n9973) );
  NOR2_X1 U11926 ( .A1(n11705), .A2(n14455), .ZN(n11722) );
  NAND2_X1 U11927 ( .A1(n11687), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11705) );
  INV_X1 U11928 ( .A(n11673), .ZN(n11687) );
  AND2_X1 U11929 ( .A1(n11658), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11659) );
  NAND2_X1 U11930 ( .A1(n11659), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11673) );
  AND4_X1 U11931 ( .A1(n11625), .A2(n11624), .A3(n11623), .A4(n11622), .ZN(
        n14014) );
  AND2_X1 U11932 ( .A1(n11606), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11628) );
  NAND2_X1 U11933 ( .A1(n11550), .A2(n11549), .ZN(n14009) );
  OAI21_X1 U11934 ( .B1(n11905), .B2(n14011), .A(n11547), .ZN(n11548) );
  CLKBUF_X1 U11935 ( .A(n14007), .Z(n14008) );
  AND2_X1 U11936 ( .A1(n11604), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11606) );
  INV_X1 U11937 ( .A(n14001), .ZN(n9760) );
  INV_X1 U11938 ( .A(n13610), .ZN(n9758) );
  AND2_X1 U11939 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11579) );
  XNOR2_X1 U11940 ( .A(n12819), .B(n13298), .ZN(n13270) );
  NOR2_X1 U11941 ( .A1(n13166), .A2(n11368), .ZN(n13265) );
  INV_X1 U11942 ( .A(n10019), .ZN(n14312) );
  NAND2_X1 U11943 ( .A1(n14607), .A2(n13065), .ZN(n14311) );
  NOR2_X1 U11944 ( .A1(n14844), .A2(n14757), .ZN(n10021) );
  AND2_X1 U11945 ( .A1(n13022), .A2(n13021), .ZN(n14363) );
  NAND2_X1 U11946 ( .A1(n14608), .A2(n14617), .ZN(n14607) );
  AND2_X1 U11947 ( .A1(n13013), .A2(n13012), .ZN(n14401) );
  AND2_X1 U11948 ( .A1(n14833), .A2(n9714), .ZN(n14432) );
  INV_X1 U11949 ( .A(n14433), .ZN(n9924) );
  NAND2_X1 U11950 ( .A1(n14833), .A2(n9925), .ZN(n14474) );
  NAND2_X1 U11951 ( .A1(n9749), .A2(n14844), .ZN(n14651) );
  NAND2_X1 U11952 ( .A1(n12894), .A2(n9664), .ZN(n9749) );
  NAND2_X1 U11953 ( .A1(n14651), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14649) );
  AND2_X1 U11954 ( .A1(n13003), .A2(n13002), .ZN(n14824) );
  NAND2_X1 U11955 ( .A1(n14833), .A2(n9927), .ZN(n14823) );
  AND2_X1 U11956 ( .A1(n14833), .A2(n14480), .ZN(n14825) );
  AND2_X1 U11957 ( .A1(n10034), .A2(n12895), .ZN(n9866) );
  XNOR2_X1 U11958 ( .A(n14841), .B(n16076), .ZN(n14697) );
  NOR2_X1 U11959 ( .A1(n14509), .A2(n12981), .ZN(n14503) );
  CLKBUF_X1 U11960 ( .A(n14693), .Z(n14694) );
  OR2_X1 U11961 ( .A1(n14451), .A2(n14452), .ZN(n14509) );
  NAND2_X1 U11962 ( .A1(n13053), .A2(n13563), .ZN(n16095) );
  AND2_X1 U11963 ( .A1(n12967), .A2(n12966), .ZN(n14526) );
  AND2_X1 U11964 ( .A1(n14527), .A2(n14526), .ZN(n14528) );
  NAND2_X1 U11965 ( .A1(n12961), .A2(n12960), .ZN(n14143) );
  INV_X1 U11966 ( .A(n14146), .ZN(n12960) );
  INV_X1 U11967 ( .A(n14145), .ZN(n12961) );
  NAND2_X1 U11968 ( .A1(n9918), .A2(n9917), .ZN(n9916) );
  INV_X1 U11969 ( .A(n9734), .ZN(n9917) );
  NAND2_X1 U11970 ( .A1(n9861), .A2(n12803), .ZN(n12861) );
  AND3_X1 U11971 ( .A1(n12948), .A2(n12990), .A3(n12947), .ZN(n14004) );
  NAND2_X1 U11972 ( .A1(n9590), .A2(n12844), .ZN(n10012) );
  NOR2_X1 U11973 ( .A1(n10015), .A2(n10016), .ZN(n10011) );
  NAND2_X1 U11974 ( .A1(n9919), .A2(n12945), .ZN(n14003) );
  INV_X1 U11975 ( .A(n16095), .ZN(n19994) );
  AND2_X1 U11976 ( .A1(n13055), .A2(n13054), .ZN(n19989) );
  INV_X1 U11977 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11458) );
  AOI21_X1 U11978 ( .B1(n11565), .B2(n11564), .A(n12804), .ZN(n11557) );
  INV_X1 U11979 ( .A(n14302), .ZN(n14875) );
  INV_X1 U11980 ( .A(n11468), .ZN(n9779) );
  NAND2_X1 U11981 ( .A1(n11408), .A2(n11468), .ZN(n9778) );
  INV_X1 U11982 ( .A(n13592), .ZN(n15814) );
  OR2_X1 U11983 ( .A1(n13601), .A2(n12818), .ZN(n20303) );
  INV_X1 U11984 ( .A(n20210), .ZN(n20445) );
  NAND2_X1 U11985 ( .A1(n20269), .A2(n20642), .ZN(n20647) );
  INV_X1 U11986 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20493) );
  INV_X1 U11987 ( .A(n12070), .ZN(n20048) );
  NAND2_X1 U11988 ( .A1(n13601), .A2(n20383), .ZN(n20354) );
  NAND2_X1 U11989 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20489) );
  NAND2_X1 U11990 ( .A1(n20268), .A2(n20154), .ZN(n20498) );
  AOI21_X1 U11991 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20415), .A(n20066), 
        .ZN(n20501) );
  OR2_X1 U11992 ( .A1(n20498), .A2(n20445), .ZN(n20452) );
  NAND3_X1 U11993 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20556), .A3(n20023), 
        .ZN(n20055) );
  NOR2_X2 U11994 ( .A1(n20020), .A2(n20022), .ZN(n20057) );
  NOR2_X2 U11995 ( .A1(n20022), .A2(n20021), .ZN(n20056) );
  NAND2_X1 U11996 ( .A1(n12677), .A2(n10551), .ZN(n10547) );
  AOI21_X1 U11997 ( .B1(n10927), .B2(n10925), .A(n10924), .ZN(n10931) );
  OR2_X1 U11998 ( .A1(n10968), .A2(n10967), .ZN(n15216) );
  AND2_X1 U11999 ( .A1(n11084), .A2(n11089), .ZN(n11093) );
  NAND2_X1 U12000 ( .A1(n11054), .A2(n9656), .ZN(n11049) );
  OR2_X1 U12001 ( .A1(n11055), .A2(n11063), .ZN(n18897) );
  AND2_X1 U12002 ( .A1(n11019), .A2(n13528), .ZN(n11023) );
  AND2_X1 U12003 ( .A1(n14974), .A2(n14959), .ZN(n15076) );
  AOI211_X1 U12004 ( .C1(n12497), .C2(n12495), .A(n12564), .B(n12500), .ZN(
        n15088) );
  AND4_X1 U12005 ( .A1(n12391), .A2(n12390), .A3(n12389), .A4(n12388), .ZN(
        n15118) );
  AOI22_X1 U12006 ( .A1(n13321), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n13749), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10588) );
  INV_X1 U12007 ( .A(n18832), .ZN(n13318) );
  AND2_X1 U12008 ( .A1(n9722), .A2(n9890), .ZN(n9889) );
  INV_X1 U12009 ( .A(n14950), .ZN(n9890) );
  NAND2_X1 U12010 ( .A1(n14978), .A2(n9722), .ZN(n15148) );
  AND2_X1 U12011 ( .A1(n12786), .A2(n12785), .ZN(n14962) );
  NAND2_X1 U12012 ( .A1(n14978), .A2(n14980), .ZN(n14979) );
  INV_X1 U12013 ( .A(n14994), .ZN(n9888) );
  AND2_X1 U12014 ( .A1(n12358), .A2(n12357), .ZN(n14192) );
  CLKBUF_X1 U12015 ( .A(n14181), .Z(n14182) );
  OR2_X1 U12016 ( .A1(n12319), .A2(n12318), .ZN(n14050) );
  CLKBUF_X1 U12017 ( .A(n14048), .Z(n14049) );
  AND3_X1 U12018 ( .A1(n12760), .A2(n12759), .A3(n12758), .ZN(n15695) );
  AND3_X1 U12019 ( .A1(n12745), .A2(n12744), .A3(n12743), .ZN(n13992) );
  NOR2_X1 U12020 ( .A1(n13917), .A2(n9896), .ZN(n13991) );
  AOI21_X1 U12021 ( .B1(n13079), .B2(n13140), .A(n19766), .ZN(n19023) );
  INV_X1 U12022 ( .A(n13129), .ZN(n13852) );
  AND2_X1 U12023 ( .A1(n9968), .A2(n9967), .ZN(n9966) );
  INV_X1 U12024 ( .A(n14943), .ZN(n9967) );
  AND2_X1 U12025 ( .A1(n14917), .A2(n9662), .ZN(n14928) );
  NAND2_X1 U12026 ( .A1(n14917), .A2(n9909), .ZN(n14923) );
  NAND2_X1 U12027 ( .A1(n14917), .A2(n9652), .ZN(n14925) );
  CLKBUF_X1 U12028 ( .A(n14917), .Z(n14919) );
  CLKBUF_X1 U12029 ( .A(n14896), .Z(n14913) );
  CLKBUF_X1 U12030 ( .A(n14911), .Z(n14912) );
  NAND2_X1 U12031 ( .A1(n14901), .A2(n9653), .ZN(n14908) );
  AND2_X1 U12032 ( .A1(n14901), .A2(n9701), .ZN(n14907) );
  AND2_X1 U12033 ( .A1(n14901), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14906) );
  NAND2_X1 U12034 ( .A1(n13672), .A2(n9693), .ZN(n13896) );
  CLKBUF_X1 U12035 ( .A(n13925), .Z(n13928) );
  INV_X1 U12036 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n14106) );
  NOR2_X1 U12037 ( .A1(n13771), .A2(n14106), .ZN(n13775) );
  NOR2_X1 U12038 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13749) );
  INV_X1 U12039 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13976) );
  XNOR2_X1 U12040 ( .A(n10605), .B(n10604), .ZN(n10619) );
  INV_X1 U12041 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15480) );
  NOR2_X1 U12042 ( .A1(n11111), .A2(n10002), .ZN(n10001) );
  INV_X1 U12043 ( .A(n15468), .ZN(n10002) );
  AND2_X1 U12044 ( .A1(n10000), .A2(n15242), .ZN(n9999) );
  NAND2_X1 U12045 ( .A1(n11111), .A2(n9739), .ZN(n10000) );
  NAND2_X1 U12046 ( .A1(n9828), .A2(n9827), .ZN(n15243) );
  AND2_X1 U12047 ( .A1(n10085), .A2(n15292), .ZN(n9827) );
  NAND2_X1 U12048 ( .A1(n14974), .A2(n9968), .ZN(n15074) );
  AND4_X1 U12049 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15465) );
  OR3_X1 U12050 ( .A1(n14961), .A2(n15240), .A3(n10914), .ZN(n15275) );
  NOR2_X1 U12051 ( .A1(n9668), .A2(n14973), .ZN(n14974) );
  NAND2_X1 U12052 ( .A1(n11171), .A2(n9963), .ZN(n15117) );
  AND2_X1 U12053 ( .A1(n14040), .A2(n9700), .ZN(n14189) );
  OR3_X1 U12054 ( .A1(n11080), .A2(n15240), .A3(n15610), .ZN(n15371) );
  NAND2_X1 U12055 ( .A1(n12762), .A2(n9695), .ZN(n15020) );
  AND2_X1 U12056 ( .A1(n12762), .A2(n9899), .ZN(n15034) );
  NAND2_X1 U12057 ( .A1(n14040), .A2(n9694), .ZN(n14179) );
  AND2_X1 U12058 ( .A1(n15692), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15656) );
  OR2_X1 U12059 ( .A1(n16293), .A2(n15464), .ZN(n15719) );
  INV_X1 U12060 ( .A(n13897), .ZN(n9959) );
  AND2_X1 U12061 ( .A1(n13895), .A2(n13907), .ZN(n14040) );
  AND2_X1 U12062 ( .A1(n9831), .A2(n15423), .ZN(n9830) );
  NAND2_X1 U12063 ( .A1(n16265), .A2(n9704), .ZN(n9833) );
  NAND2_X1 U12064 ( .A1(n11017), .A2(n10003), .ZN(n15322) );
  NOR2_X1 U12065 ( .A1(n15736), .A2(n16267), .ZN(n10004) );
  NOR2_X1 U12066 ( .A1(n13526), .A2(n13525), .ZN(n13672) );
  NAND2_X1 U12067 ( .A1(n13672), .A2(n13671), .ZN(n13674) );
  NAND2_X1 U12068 ( .A1(n11017), .A2(n11016), .ZN(n15734) );
  NOR2_X1 U12069 ( .A1(n13917), .A2(n13918), .ZN(n16287) );
  OR2_X1 U12070 ( .A1(n13519), .A2(n13520), .ZN(n13526) );
  INV_X1 U12071 ( .A(n13374), .ZN(n9957) );
  XNOR2_X1 U12072 ( .A(n9818), .B(n14166), .ZN(n14097) );
  NAND2_X1 U12073 ( .A1(n13820), .A2(n10787), .ZN(n14030) );
  AND2_X1 U12074 ( .A1(n13825), .A2(n15611), .ZN(n14167) );
  AND3_X1 U12075 ( .A1(n12724), .A2(n12723), .A3(n12722), .ZN(n13833) );
  NAND2_X1 U12076 ( .A1(n13831), .A2(n15659), .ZN(n15611) );
  AOI21_X1 U12077 ( .B1(n12141), .B2(n12156), .A(n12140), .ZN(n13191) );
  AND2_X1 U12078 ( .A1(n19520), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19728) );
  AND2_X1 U12079 ( .A1(n19721), .A2(n19732), .ZN(n19143) );
  NOR2_X2 U12080 ( .A1(n10634), .A2(n10633), .ZN(n19169) );
  INV_X1 U12081 ( .A(n19143), .ZN(n19380) );
  NAND2_X1 U12082 ( .A1(n19721), .A2(n14073), .ZN(n19707) );
  OR2_X1 U12083 ( .A1(n19145), .A2(n19739), .ZN(n19494) );
  NAND2_X2 U12084 ( .A1(n10520), .A2(n10519), .ZN(n19103) );
  NAND2_X1 U12085 ( .A1(n10088), .A2(n9680), .ZN(n10520) );
  NAND2_X1 U12086 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19573), .ZN(n19108) );
  INV_X1 U12087 ( .A(n19126), .ZN(n19116) );
  INV_X1 U12088 ( .A(n19127), .ZN(n19117) );
  NOR2_X2 U12089 ( .A1(n13852), .A2(n13851), .ZN(n19126) );
  NOR2_X2 U12090 ( .A1(n13850), .A2(n13851), .ZN(n19127) );
  OR2_X1 U12091 ( .A1(n19145), .A2(n19144), .ZN(n19519) );
  OR2_X1 U12092 ( .A1(n19494), .A2(n19568), .ZN(n19085) );
  INV_X1 U12093 ( .A(n19108), .ZN(n19124) );
  NAND2_X1 U12094 ( .A1(n13304), .A2(n12654), .ZN(n13842) );
  NAND2_X1 U12095 ( .A1(n10537), .A2(n12653), .ZN(n12654) );
  NOR2_X1 U12096 ( .A1(n16564), .A2(n17461), .ZN(n16563) );
  NAND2_X1 U12097 ( .A1(n17673), .A2(n17714), .ZN(n16738) );
  NOR2_X1 U12098 ( .A1(n10054), .A2(n10050), .ZN(n10049) );
  INV_X1 U12099 ( .A(n10139), .ZN(n10055) );
  INV_X1 U12100 ( .A(n18617), .ZN(n15879) );
  NOR2_X1 U12101 ( .A1(n17398), .A2(n17348), .ZN(n17368) );
  NAND2_X1 U12102 ( .A1(n17487), .A2(n9941), .ZN(n16365) );
  AND2_X1 U12103 ( .A1(n9941), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9940) );
  NAND2_X1 U12104 ( .A1(n17487), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17471) );
  NAND2_X1 U12105 ( .A1(n9936), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9935) );
  INV_X1 U12106 ( .A(n17575), .ZN(n9936) );
  INV_X1 U12107 ( .A(n17612), .ZN(n9945) );
  NOR2_X1 U12108 ( .A1(n17798), .A2(n17762), .ZN(n17702) );
  NOR2_X1 U12109 ( .A1(n16325), .A2(n18658), .ZN(n16332) );
  NOR2_X1 U12110 ( .A1(n9793), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9792) );
  INV_X1 U12111 ( .A(n9794), .ZN(n9793) );
  NOR2_X1 U12112 ( .A1(n17560), .A2(n10222), .ZN(n17516) );
  AND2_X1 U12113 ( .A1(n10221), .A2(n10220), .ZN(n10222) );
  NAND2_X1 U12114 ( .A1(n9842), .A2(n10402), .ZN(n10221) );
  NOR2_X1 U12115 ( .A1(n17594), .A2(n17722), .ZN(n17560) );
  OAI211_X1 U12116 ( .C1(n10218), .C2(n17957), .A(n10217), .B(n9707), .ZN(
        n17595) );
  NOR2_X1 U12117 ( .A1(n17595), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17594) );
  INV_X1 U12118 ( .A(n9842), .ZN(n17605) );
  NOR2_X1 U12119 ( .A1(n17640), .A2(n10208), .ZN(n17929) );
  NOR2_X1 U12120 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17667), .ZN(
        n17642) );
  INV_X1 U12121 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17979) );
  INV_X1 U12122 ( .A(n18014), .ZN(n17990) );
  NAND2_X1 U12123 ( .A1(n10215), .A2(n9855), .ZN(n17667) );
  NOR2_X1 U12124 ( .A1(n9856), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9855) );
  INV_X1 U12125 ( .A(n9857), .ZN(n9856) );
  INV_X1 U12126 ( .A(n18631), .ZN(n10401) );
  NOR2_X1 U12127 ( .A1(n9858), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9857) );
  INV_X1 U12128 ( .A(n9859), .ZN(n9858) );
  NAND2_X1 U12129 ( .A1(n18059), .A2(n17722), .ZN(n17721) );
  XNOR2_X1 U12130 ( .A(n10206), .B(n10205), .ZN(n17728) );
  INV_X1 U12131 ( .A(n10204), .ZN(n10205) );
  XNOR2_X1 U12132 ( .A(n10199), .B(n10198), .ZN(n17751) );
  NAND2_X1 U12133 ( .A1(n17751), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17750) );
  XNOR2_X1 U12134 ( .A(n17339), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17801) );
  NAND2_X1 U12135 ( .A1(n17809), .A2(n17801), .ZN(n17800) );
  OR3_X1 U12136 ( .A1(n17120), .A2(n14203), .A3(n15876), .ZN(n10397) );
  NOR2_X1 U12137 ( .A1(n18822), .A2(n14204), .ZN(n18639) );
  NAND2_X1 U12138 ( .A1(n18778), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n18635) );
  INV_X1 U12139 ( .A(n18639), .ZN(n18613) );
  NOR2_X1 U12140 ( .A1(n10244), .A2(n10243), .ZN(n18167) );
  INV_X1 U12141 ( .A(n10390), .ZN(n18179) );
  NOR2_X1 U12142 ( .A1(n10286), .A2(n10285), .ZN(n18191) );
  INV_X1 U12143 ( .A(n17201), .ZN(n18195) );
  NAND3_X1 U12144 ( .A1(n10317), .A2(n10316), .A3(n10315), .ZN(n18161) );
  NOR2_X1 U12145 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18159), .ZN(n18414) );
  INV_X1 U12146 ( .A(n18414), .ZN(n18509) );
  NOR3_X1 U12147 ( .A1(n18808), .A2(n18820), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n18812) );
  INV_X1 U12148 ( .A(n14301), .ZN(n19780) );
  NAND2_X1 U12149 ( .A1(n14324), .A2(n14325), .ZN(n20667) );
  INV_X1 U12150 ( .A(n19875), .ZN(n19821) );
  INV_X1 U12151 ( .A(n19884), .ZN(n19862) );
  INV_X1 U12152 ( .A(n19864), .ZN(n19879) );
  XNOR2_X1 U12153 ( .A(n11483), .B(n20157), .ZN(n20272) );
  AND2_X1 U12154 ( .A1(n13639), .A2(n13633), .ZN(n19884) );
  INV_X1 U12155 ( .A(n11436), .ZN(n11437) );
  AND2_X1 U12156 ( .A1(n14317), .A2(n13628), .ZN(n19852) );
  AND2_X1 U12157 ( .A1(n19831), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19876) );
  INV_X1 U12158 ( .A(n14515), .ZN(n19895) );
  INV_X1 U12159 ( .A(n14532), .ZN(n19894) );
  AND2_X2 U12160 ( .A1(n13278), .A2(n14301), .ZN(n19899) );
  INV_X1 U12161 ( .A(n16015), .ZN(n14566) );
  OR2_X1 U12162 ( .A1(n14519), .A2(n14518), .ZN(n15976) );
  NAND2_X1 U12163 ( .A1(n12115), .A2(n12114), .ZN(n14571) );
  INV_X1 U12164 ( .A(n14580), .ZN(n14573) );
  AND2_X1 U12165 ( .A1(n13229), .A2(n13264), .ZN(n19903) );
  AND2_X1 U12166 ( .A1(n11399), .A2(n20567), .ZN(n13295) );
  XNOR2_X1 U12167 ( .A(n13625), .B(n14336), .ZN(n14317) );
  OR2_X1 U12168 ( .A1(n13624), .A2(n14584), .ZN(n13625) );
  INV_X1 U12169 ( .A(n14320), .ZN(n9762) );
  INV_X1 U12170 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15926) );
  AND2_X1 U12171 ( .A1(n14498), .A2(n14507), .ZN(n15964) );
  NAND2_X1 U12172 ( .A1(n9752), .A2(n13458), .ZN(n13459) );
  INV_X1 U12173 ( .A(n14723), .ZN(n19962) );
  XNOR2_X1 U12174 ( .A(n14323), .B(n14328), .ZN(n14745) );
  NAND2_X1 U12175 ( .A1(n10020), .A2(n14746), .ZN(n9864) );
  OR2_X1 U12176 ( .A1(n14829), .A2(n13060), .ZN(n14810) );
  NAND2_X1 U12177 ( .A1(n9867), .A2(n10034), .ZN(n14689) );
  NAND2_X1 U12178 ( .A1(n13538), .A2(n12837), .ZN(n19965) );
  AND2_X1 U12179 ( .A1(n16093), .A2(n13046), .ZN(n19988) );
  AND2_X1 U12180 ( .A1(n13053), .A2(n13031), .ZN(n19981) );
  INV_X1 U12181 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20415) );
  INV_X1 U12182 ( .A(n14873), .ZN(n20499) );
  INV_X1 U12183 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20019) );
  NAND2_X1 U12184 ( .A1(n13600), .A2(n20066), .ZN(n20653) );
  AND2_X1 U12185 ( .A1(n12899), .A2(n11367), .ZN(n14877) );
  NOR2_X1 U12186 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n14880) );
  INV_X1 U12187 ( .A(n20553), .ZN(n20058) );
  INV_X1 U12188 ( .A(n20114), .ZN(n20116) );
  INV_X1 U12189 ( .A(n20153), .ZN(n20145) );
  OAI21_X1 U12190 ( .B1(n9737), .B2(n20163), .A(n20450), .ZN(n20181) );
  INV_X1 U12191 ( .A(n20178), .ZN(n20180) );
  INV_X1 U12192 ( .A(n20208), .ZN(n20200) );
  OR2_X1 U12193 ( .A1(n20639), .A2(n20445), .ZN(n20267) );
  OAI211_X1 U12194 ( .C1(n10080), .C2(n20389), .A(n20328), .B(n20279), .ZN(
        n20296) );
  INV_X1 U12195 ( .A(n20353), .ZN(n20345) );
  OAI22_X1 U12196 ( .A1(n20332), .A2(n20331), .B1(n20330), .B2(n20443), .ZN(
        n20349) );
  INV_X1 U12197 ( .A(n20376), .ZN(n20379) );
  NOR2_X1 U12198 ( .A1(n20389), .A2(n13599), .ZN(n15846) );
  INV_X1 U12199 ( .A(n16170), .ZN(n16168) );
  INV_X1 U12200 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20555) );
  INV_X1 U12201 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20389) );
  NOR2_X1 U12202 ( .A1(n10528), .A2(n10540), .ZN(n10531) );
  NAND2_X1 U12203 ( .A1(n15804), .A2(n18893), .ZN(n16222) );
  NAND2_X1 U12204 ( .A1(n15002), .A2(n18893), .ZN(n18862) );
  OR2_X1 U12205 ( .A1(n16172), .A2(n13792), .ZN(n18922) );
  NAND2_X1 U12206 ( .A1(n11054), .A2(n9875), .ZN(n11044) );
  NOR2_X1 U12207 ( .A1(n9903), .A2(n9682), .ZN(n9902) );
  NAND2_X1 U12208 ( .A1(n15030), .A2(n15400), .ZN(n15029) );
  INV_X1 U12209 ( .A(n18947), .ZN(n18901) );
  INV_X1 U12210 ( .A(n18935), .ZN(n18931) );
  INV_X1 U12211 ( .A(n18922), .ZN(n18954) );
  INV_X1 U12212 ( .A(n19628), .ZN(n18949) );
  NAND2_X1 U12213 ( .A1(n19758), .A2(n13786), .ZN(n18936) );
  NOR2_X2 U12214 ( .A1(n19758), .A2(n13784), .ZN(n18940) );
  OR2_X1 U12215 ( .A1(n12305), .A2(n12304), .ZN(n14045) );
  CLKBUF_X1 U12216 ( .A(n13899), .Z(n13900) );
  OR2_X1 U12217 ( .A1(n12258), .A2(n12257), .ZN(n13666) );
  AND4_X1 U12218 ( .A1(n12220), .A2(n12219), .A3(n12218), .A4(n12217), .ZN(
        n12221) );
  OR2_X1 U12219 ( .A1(n12183), .A2(n12182), .ZN(n13416) );
  NOR2_X1 U12220 ( .A1(n10068), .A2(n9725), .ZN(n10067) );
  INV_X1 U12221 ( .A(n13242), .ZN(n10068) );
  INV_X1 U12222 ( .A(n15114), .ZN(n15119) );
  INV_X1 U12223 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n14115) );
  INV_X1 U12224 ( .A(n13198), .ZN(n15110) );
  NAND2_X1 U12225 ( .A1(n15110), .A2(n9622), .ZN(n15114) );
  OAI21_X1 U12226 ( .B1(n15053), .B2(n15054), .A(n9721), .ZN(n12634) );
  AOI21_X1 U12227 ( .B1(n15068), .B2(n15070), .A(n15069), .ZN(n15071) );
  XNOR2_X1 U12228 ( .A(n12520), .B(n12519), .ZN(n15082) );
  AND2_X1 U12229 ( .A1(n15006), .A2(n15004), .ZN(n15190) );
  AND2_X1 U12230 ( .A1(n13515), .A2(n13850), .ZN(n18955) );
  AND2_X1 U12231 ( .A1(n19014), .A2(n12684), .ZN(n16235) );
  NAND2_X1 U12232 ( .A1(n15156), .A2(n13516), .ZN(n19012) );
  INV_X1 U12233 ( .A(n19014), .ZN(n19015) );
  INV_X1 U12234 ( .A(n15206), .ZN(n19016) );
  INV_X1 U12235 ( .A(n15185), .ZN(n19017) );
  INV_X1 U12236 ( .A(n19012), .ZN(n19022) );
  AND2_X2 U12237 ( .A1(n13791), .A2(n12687), .ZN(n13788) );
  NAND2_X1 U12238 ( .A1(n9836), .A2(n9834), .ZN(n15223) );
  INV_X1 U12239 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15303) );
  INV_X1 U12240 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15409) );
  INV_X1 U12241 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15425) );
  INV_X1 U12242 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19068) );
  NAND2_X1 U12243 ( .A1(n18834), .A2(n11210), .ZN(n19067) );
  INV_X1 U12244 ( .A(n19059), .ZN(n16262) );
  INV_X1 U12245 ( .A(n19067), .ZN(n19069) );
  XNOR2_X1 U12246 ( .A(n15050), .B(n15049), .ZN(n16175) );
  INV_X1 U12247 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15682) );
  INV_X1 U12248 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16275) );
  INV_X1 U12249 ( .A(n15440), .ZN(n10909) );
  AND2_X1 U12250 ( .A1(n9958), .A2(n9647), .ZN(n13246) );
  INV_X1 U12251 ( .A(n16308), .ZN(n16282) );
  NOR2_X1 U12252 ( .A1(n19350), .A2(n19726), .ZN(n19742) );
  AND2_X1 U12253 ( .A1(n13194), .A2(n13193), .ZN(n19732) );
  OR2_X1 U12254 ( .A1(n13192), .A2(n13191), .ZN(n13193) );
  INV_X1 U12255 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15875) );
  NAND2_X1 U12256 ( .A1(n19079), .A2(n12156), .ZN(n12138) );
  INV_X1 U12257 ( .A(n19732), .ZN(n14073) );
  AOI21_X1 U12258 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19762), .A(n13222), 
        .ZN(n15768) );
  OAI21_X1 U12259 ( .B1(n19092), .B2(n19091), .A(n19090), .ZN(n19132) );
  AOI211_X2 U12260 ( .C1(n19088), .C2(n19091), .A(n19523), .B(n19084), .ZN(
        n19135) );
  INV_X1 U12261 ( .A(n19166), .ZN(n19156) );
  NOR2_X1 U12262 ( .A1(n19380), .A2(n19327), .ZN(n19188) );
  INV_X1 U12263 ( .A(n19233), .ZN(n19251) );
  INV_X1 U12264 ( .A(n19266), .ZN(n19283) );
  NOR2_X2 U12265 ( .A1(n19288), .A2(n19493), .ZN(n19281) );
  INV_X1 U12266 ( .A(n19294), .ZN(n19312) );
  NOR2_X1 U12267 ( .A1(n19568), .A2(n19288), .ZN(n19344) );
  INV_X1 U12268 ( .A(n19326), .ZN(n19345) );
  INV_X1 U12269 ( .A(n19379), .ZN(n19371) );
  INV_X1 U12270 ( .A(n19401), .ZN(n19404) );
  NOR2_X1 U12271 ( .A1(n19494), .A2(n19380), .ZN(n19428) );
  OAI22_X1 U12272 ( .A1(n20707), .A2(n19117), .B1(n19102), .B2(n19116), .ZN(
        n19499) );
  OAI22_X1 U12273 ( .A1(n20785), .A2(n19116), .B1(n19107), .B2(n19117), .ZN(
        n19538) );
  OR3_X1 U12274 ( .A1(n19524), .A2(n19523), .A3(n19522), .ZN(n19558) );
  OAI21_X1 U12275 ( .B1(n19529), .B2(n19528), .A(n19527), .ZN(n19557) );
  INV_X1 U12276 ( .A(n19545), .ZN(n19555) );
  OAI22_X1 U12277 ( .A1(n16385), .A2(n19117), .B1(n18200), .B2(n19116), .ZN(
        n19556) );
  INV_X1 U12278 ( .A(n19535), .ZN(n19580) );
  INV_X1 U12279 ( .A(n19502), .ZN(n19586) );
  INV_X1 U12280 ( .A(n19499), .ZN(n19589) );
  INV_X1 U12281 ( .A(n19541), .ZN(n19591) );
  INV_X1 U12282 ( .A(n19538), .ZN(n19594) );
  AOI22_X1 U12283 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19127), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19126), .ZN(n19600) );
  AND2_X1 U12284 ( .A1(n10548), .A2(n19124), .ZN(n19595) );
  AOI22_X1 U12285 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19126), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19127), .ZN(n19606) );
  INV_X1 U12286 ( .A(n19549), .ZN(n19603) );
  AND2_X1 U12287 ( .A1(n12678), .A2(n19124), .ZN(n19601) );
  AND2_X1 U12288 ( .A1(n10550), .A2(n19124), .ZN(n19607) );
  INV_X1 U12289 ( .A(n19085), .ZN(n19618) );
  INV_X1 U12290 ( .A(n19561), .ZN(n19617) );
  OR2_X1 U12291 ( .A1(n19631), .A2(n19350), .ZN(n18832) );
  AND2_X1 U12292 ( .A1(n19741), .A2(n10943), .ZN(n16319) );
  NAND2_X1 U12293 ( .A1(n13842), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16320) );
  INV_X1 U12294 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18820) );
  INV_X1 U12295 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18808) );
  INV_X1 U12296 ( .A(n17875), .ZN(n18794) );
  INV_X1 U12297 ( .A(n16332), .ZN(n16494) );
  AND2_X1 U12298 ( .A1(n9946), .A2(n17479), .ZN(n16571) );
  NOR2_X1 U12299 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16721), .ZN(n16704) );
  NOR2_X1 U12300 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16743), .ZN(n16730) );
  OAI211_X1 U12301 ( .C1(n16510), .C2(n18435), .A(n16776), .B(n18810), .ZN(
        n16855) );
  INV_X1 U12302 ( .A(n16833), .ZN(n16868) );
  INV_X1 U12303 ( .A(n16843), .ZN(n16875) );
  AND2_X1 U12304 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16991), .ZN(n16977) );
  NAND2_X1 U12305 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17045), .ZN(n17029) );
  AND2_X1 U12306 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17031), .ZN(n17045) );
  NOR3_X1 U12307 ( .A1(n15877), .A2(n14208), .A3(n18658), .ZN(n17195) );
  NAND2_X1 U12308 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17223), .ZN(n17218) );
  INV_X1 U12309 ( .A(n17233), .ZN(n17228) );
  NAND2_X1 U12310 ( .A1(n17234), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n17233) );
  INV_X1 U12311 ( .A(n17249), .ZN(n17273) );
  INV_X1 U12312 ( .A(n17237), .ZN(n17274) );
  AOI22_X1 U12313 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10296) );
  NAND2_X1 U12314 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17307), .ZN(n17302) );
  AND3_X1 U12315 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(n17314), .ZN(n17307) );
  NAND2_X1 U12316 ( .A1(n17196), .A2(n18204), .ZN(n17327) );
  INV_X1 U12317 ( .A(n10353), .ZN(n17334) );
  NAND2_X1 U12318 ( .A1(n15879), .A2(n17196), .ZN(n17335) );
  INV_X1 U12319 ( .A(n17341), .ZN(n17338) );
  NAND2_X1 U12320 ( .A1(n17196), .A2(P3_EAX_REG_1__SCAN_IN), .ZN(n17343) );
  NOR2_X1 U12321 ( .A1(n17327), .A2(n15879), .ZN(n17341) );
  INV_X1 U12322 ( .A(n17335), .ZN(n17340) );
  AOI21_X1 U12323 ( .B1(n17400), .B2(n17399), .A(n17398), .ZN(n17430) );
  NOR2_X2 U12324 ( .A1(n18804), .A2(n17454), .ZN(n17449) );
  INV_X1 U12325 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17457) );
  NOR2_X2 U12326 ( .A1(n17454), .A2(n18167), .ZN(n17455) );
  INV_X1 U12327 ( .A(n17449), .ZN(n20803) );
  NOR2_X1 U12328 ( .A1(n17574), .A2(n9930), .ZN(n17524) );
  NAND2_X1 U12329 ( .A1(n17538), .A2(n9931), .ZN(n9930) );
  INV_X1 U12330 ( .A(n9935), .ZN(n9931) );
  INV_X1 U12331 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17544) );
  NOR2_X1 U12332 ( .A1(n16341), .A2(n17709), .ZN(n17601) );
  NAND2_X1 U12333 ( .A1(n16798), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17743) );
  INV_X1 U12334 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17747) );
  NOR2_X2 U12335 ( .A1(n18509), .A2(n18411), .ZN(n18545) );
  INV_X1 U12336 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17804) );
  INV_X1 U12337 ( .A(n17795), .ZN(n17805) );
  NAND2_X1 U12338 ( .A1(n18808), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17812) );
  NAND2_X1 U12339 ( .A1(n10226), .A2(n9794), .ZN(n15794) );
  NOR2_X1 U12340 ( .A1(n9846), .A2(n17463), .ZN(n9845) );
  AND2_X1 U12341 ( .A1(n10043), .A2(n9715), .ZN(n17493) );
  NAND2_X1 U12342 ( .A1(n10224), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10043) );
  OR2_X1 U12343 ( .A1(n17886), .A2(n17885), .ZN(n17868) );
  INV_X1 U12344 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17957) );
  NAND2_X1 U12345 ( .A1(n10215), .A2(n9859), .ZN(n17689) );
  NOR2_X1 U12346 ( .A1(n10216), .A2(n17722), .ZN(n17698) );
  INV_X1 U12347 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n20725) );
  AND2_X1 U12348 ( .A1(n10046), .A2(n10047), .ZN(n17768) );
  NAND2_X1 U12349 ( .A1(n17779), .A2(n18110), .ZN(n10046) );
  AOI21_X2 U12350 ( .B1(n15777), .B2(n10351), .A(n18658), .ZN(n18127) );
  INV_X1 U12351 ( .A(n18127), .ZN(n18143) );
  INV_X1 U12352 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18156) );
  OAI211_X1 U12353 ( .C1(n18658), .C2(n18626), .A(n18160), .B(n15781), .ZN(
        n18782) );
  INV_X1 U12354 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18176) );
  INV_X1 U12355 ( .A(n18812), .ZN(n18658) );
  INV_X1 U12356 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18752) );
  OAI211_X1 U12357 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18677), .B(n18743), .ZN(n18674) );
  CLKBUF_X1 U12358 ( .A(n16468), .Z(n16477) );
  INV_X1 U12359 ( .A(n9782), .ZN(n14606) );
  AOI21_X1 U12360 ( .B1(n16032), .B2(n14605), .A(n14604), .ZN(n9783) );
  NOR4_X1 U12361 ( .A1(n14742), .A2(n14741), .A3(n14740), .A4(n14739), .ZN(
        n14743) );
  OAI211_X1 U12362 ( .C1(n14755), .C2(n16126), .A(n9914), .B(n9913), .ZN(
        P1_U3001) );
  NOR2_X1 U12363 ( .A1(n9915), .A2(n14754), .ZN(n9914) );
  OR2_X1 U12364 ( .A1(n14745), .A2(n20017), .ZN(n9913) );
  OR2_X1 U12365 ( .A1(n14752), .A2(n14753), .ZN(n9915) );
  AND2_X1 U12366 ( .A1(n13069), .A2(n9691), .ZN(n9812) );
  OAI21_X1 U12367 ( .B1(n15492), .B2(n19075), .A(n9954), .ZN(P2_U2984) );
  NAND2_X1 U12368 ( .A1(n9956), .A2(n9955), .ZN(n9880) );
  INV_X1 U12369 ( .A(n15239), .ZN(n9955) );
  AOI21_X1 U12370 ( .B1(n11221), .B2(n19078), .A(n11220), .ZN(n11222) );
  AOI21_X1 U12371 ( .B1(n15490), .B2(n16281), .A(n15489), .ZN(n15491) );
  AOI21_X1 U12372 ( .B1(n15487), .B2(n15739), .A(n15486), .ZN(n15488) );
  AOI21_X1 U12373 ( .B1(n9938), .B2(n18661), .A(n9937), .ZN(n16550) );
  OR2_X1 U12374 ( .A1(n16546), .A2(n16547), .ZN(n9937) );
  AOI21_X1 U12375 ( .B1(n16337), .B2(n17723), .A(n16336), .ZN(n16338) );
  OAI21_X1 U12376 ( .B1(n16340), .B2(n18125), .A(n10417), .ZN(n10418) );
  AOI21_X1 U12377 ( .B1(n16349), .B2(n18057), .A(n10056), .ZN(n15854) );
  OR2_X1 U12378 ( .A1(n15853), .A2(n16348), .ZN(n10056) );
  INV_X2 U12379 ( .A(n9593), .ZN(n17153) );
  INV_X1 U12380 ( .A(n10093), .ZN(n16952) );
  INV_X1 U12381 ( .A(n9674), .ZN(n17080) );
  OR2_X1 U12382 ( .A1(n11116), .A2(n11115), .ZN(n9647) );
  NAND2_X1 U12383 ( .A1(n17516), .A2(n17520), .ZN(n17515) );
  INV_X1 U12384 ( .A(n17515), .ZN(n10038) );
  INV_X1 U12385 ( .A(n12894), .ZN(n14661) );
  NAND2_X1 U12386 ( .A1(n9973), .A2(n11739), .ZN(n14490) );
  AND2_X1 U12387 ( .A1(n12911), .A2(n11371), .ZN(n11373) );
  AND2_X1 U12388 ( .A1(n14478), .A2(n9982), .ZN(n14416) );
  NAND2_X1 U12389 ( .A1(n9976), .A2(n9979), .ZN(n14441) );
  INV_X1 U12390 ( .A(n10599), .ZN(n11121) );
  NAND2_X1 U12391 ( .A1(n17727), .A2(n9785), .ZN(n10216) );
  NAND2_X1 U12392 ( .A1(n9907), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9649) );
  AND2_X1 U12393 ( .A1(n17780), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9650) );
  AND2_X1 U12394 ( .A1(n12683), .A2(n12678), .ZN(n12714) );
  INV_X2 U12395 ( .A(n11126), .ZN(n11148) );
  NAND2_X1 U12396 ( .A1(n15006), .A2(n9720), .ZN(n14993) );
  AND3_X1 U12397 ( .A1(n11320), .A2(n11319), .A3(n20024), .ZN(n9651) );
  NAND2_X1 U12398 ( .A1(n11113), .A2(n11117), .ZN(n9958) );
  NAND2_X1 U12399 ( .A1(n9904), .A2(n9907), .ZN(n13774) );
  NAND2_X1 U12400 ( .A1(n9958), .A2(n9724), .ZN(n13252) );
  AND2_X1 U12401 ( .A1(n14191), .A2(n9723), .ZN(n15108) );
  AND2_X1 U12402 ( .A1(n9909), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9652) );
  NAND2_X1 U12403 ( .A1(n9758), .A2(n9784), .ZN(n13678) );
  AND2_X1 U12404 ( .A1(n9701), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9653) );
  AND2_X1 U12405 ( .A1(n9763), .A2(n11234), .ZN(n11530) );
  NAND2_X1 U12406 ( .A1(n13415), .A2(n10060), .ZN(n9654) );
  NAND2_X1 U12407 ( .A1(n12204), .A2(n12203), .ZN(n9655) );
  AND2_X1 U12408 ( .A1(n9875), .A2(n11043), .ZN(n9656) );
  AND2_X1 U12409 ( .A1(n9862), .A2(n11541), .ZN(n9657) );
  OR2_X1 U12410 ( .A1(n10044), .A2(n10042), .ZN(n9658) );
  AND2_X1 U12411 ( .A1(n12291), .A2(n14045), .ZN(n9659) );
  AND2_X1 U12412 ( .A1(n9723), .A2(n15109), .ZN(n9660) );
  NAND2_X1 U12413 ( .A1(n12244), .A2(n12243), .ZN(n9661) );
  AND2_X1 U12414 ( .A1(n9652), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9662) );
  XNOR2_X2 U12415 ( .A(n16326), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16531) );
  NOR2_X1 U12416 ( .A1(n13682), .A2(n9916), .ZN(n14016) );
  OR2_X1 U12417 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17722), .ZN(
        n9663) );
  AND2_X1 U12418 ( .A1(n12893), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9664) );
  AND2_X1 U12419 ( .A1(n9664), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9665) );
  AND2_X1 U12420 ( .A1(n10913), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9666) );
  AND2_X1 U12421 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9667) );
  CLKBUF_X3 U12422 ( .A(n12922), .Z(n13009) );
  AND2_X1 U12423 ( .A1(n11372), .A2(n11367), .ZN(n12946) );
  INV_X1 U12424 ( .A(n12946), .ZN(n13285) );
  INV_X1 U12425 ( .A(n10673), .ZN(n12394) );
  OR2_X1 U12426 ( .A1(n15096), .A2(n15097), .ZN(n9668) );
  OR2_X1 U12427 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10936), .ZN(
        n9669) );
  INV_X1 U12428 ( .A(n18893), .ZN(n18942) );
  OR2_X1 U12429 ( .A1(n17574), .A2(n9932), .ZN(n9670) );
  CLKBUF_X3 U12430 ( .A(n10180), .Z(n17159) );
  INV_X1 U12431 ( .A(n10166), .ZN(n14282) );
  NOR2_X2 U12432 ( .A1(n18633), .A2(n10098), .ZN(n10099) );
  NAND2_X2 U12433 ( .A1(n13196), .A2(n10600), .ZN(n9671) );
  NOR2_X1 U12434 ( .A1(n17812), .A2(n17798), .ZN(n17596) );
  NAND2_X1 U12435 ( .A1(n9828), .A2(n15292), .ZN(n15267) );
  OR3_X1 U12436 ( .A1(n14373), .A2(n9987), .A3(n9985), .ZN(n9672) );
  NAND2_X1 U12437 ( .A1(n15265), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15258) );
  NAND2_X1 U12438 ( .A1(n16264), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15731) );
  NOR2_X1 U12439 ( .A1(n14497), .A2(n9974), .ZN(n14491) );
  NAND2_X1 U12440 ( .A1(n14478), .A2(n11840), .ZN(n14469) );
  NAND2_X1 U12441 ( .A1(n9600), .A2(n10913), .ZN(n15369) );
  NAND2_X1 U12442 ( .A1(n16264), .A2(n9953), .ZN(n9673) );
  INV_X2 U12443 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10430) );
  NAND2_X1 U12444 ( .A1(n15308), .A2(n15307), .ZN(n15309) );
  INV_X1 U12445 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17674) );
  INV_X1 U12446 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13145) );
  INV_X1 U12447 ( .A(n11368), .ZN(n9772) );
  AND4_X1 U12448 ( .A1(n11231), .A2(n11230), .A3(n11229), .A4(n11228), .ZN(
        n9675) );
  AND2_X1 U12449 ( .A1(n10226), .A2(n17818), .ZN(n9676) );
  NAND2_X1 U12450 ( .A1(n14478), .A2(n9984), .ZN(n9677) );
  OAI21_X1 U12451 ( .B1(n15243), .B2(n10001), .A(n9999), .ZN(n15212) );
  AND2_X1 U12452 ( .A1(n9647), .A2(n13245), .ZN(n9678) );
  NAND2_X1 U12453 ( .A1(n15309), .A2(n11092), .ZN(n15290) );
  NAND2_X1 U12454 ( .A1(n12882), .A2(n12881), .ZN(n14149) );
  NAND2_X1 U12455 ( .A1(n15322), .A2(n15323), .ZN(n15422) );
  NOR2_X1 U12456 ( .A1(n14013), .A2(n9981), .ZN(n14127) );
  NAND2_X1 U12457 ( .A1(n14729), .A2(n12883), .ZN(n14704) );
  NAND2_X1 U12458 ( .A1(n9600), .A2(n9666), .ZN(n15352) );
  AND3_X1 U12459 ( .A1(n9957), .A2(n9678), .A3(n13250), .ZN(n9679) );
  NAND2_X1 U12460 ( .A1(n13338), .A2(n10527), .ZN(n10573) );
  AND2_X1 U12461 ( .A1(n10512), .A2(n10511), .ZN(n9680) );
  NAND2_X1 U12462 ( .A1(n9628), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9823) );
  INV_X1 U12463 ( .A(n13683), .ZN(n12945) );
  AND2_X1 U12464 ( .A1(n15162), .A2(n15163), .ZN(n14978) );
  NOR2_X1 U12465 ( .A1(n15291), .A2(n9829), .ZN(n9681) );
  NOR2_X1 U12466 ( .A1(n18892), .A2(n18895), .ZN(n9682) );
  NAND2_X1 U12467 ( .A1(n10022), .A2(n10021), .ZN(n9683) );
  AND2_X1 U12468 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n9945), .ZN(
        n9684) );
  INV_X1 U12469 ( .A(n12844), .ZN(n10015) );
  INV_X1 U12470 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15442) );
  AND2_X1 U12471 ( .A1(n12070), .A2(n12045), .ZN(n9685) );
  NAND2_X1 U12472 ( .A1(n11017), .A2(n10004), .ZN(n9686) );
  OR2_X1 U12473 ( .A1(n15850), .A2(n17722), .ZN(n9795) );
  NAND2_X1 U12474 ( .A1(n15265), .A2(n9667), .ZN(n15249) );
  AND3_X1 U12475 ( .A1(n11469), .A2(n11468), .A3(n11467), .ZN(n9688) );
  BUF_X1 U12476 ( .A(n10549), .Z(n19109) );
  AND2_X1 U12477 ( .A1(n16694), .A2(n9684), .ZN(n9689) );
  INV_X1 U12478 ( .A(n9791), .ZN(n15850) );
  NAND2_X1 U12479 ( .A1(n10226), .A2(n9792), .ZN(n9791) );
  OR2_X1 U12480 ( .A1(n9823), .A2(n10584), .ZN(n9690) );
  NOR2_X1 U12481 ( .A1(n12700), .A2(n12699), .ZN(n12709) );
  AND2_X1 U12482 ( .A1(n10075), .A2(n13070), .ZN(n9691) );
  AND2_X1 U12483 ( .A1(n11108), .A2(n15275), .ZN(n15242) );
  OR2_X1 U12484 ( .A1(n11224), .A2(n11223), .ZN(P2_U2985) );
  INV_X1 U12485 ( .A(n12706), .ZN(n12712) );
  NOR2_X1 U12486 ( .A1(n17574), .A2(n17575), .ZN(n16524) );
  NAND2_X1 U12487 ( .A1(n9990), .A2(n11003), .ZN(n14160) );
  NOR2_X1 U12488 ( .A1(n14013), .A2(n14140), .ZN(n14128) );
  NAND2_X1 U12489 ( .A1(n14191), .A2(n9660), .ZN(n15103) );
  AND2_X1 U12490 ( .A1(n13899), .A2(n9659), .ZN(n14043) );
  OR2_X1 U12491 ( .A1(n13917), .A2(n9897), .ZN(n13990) );
  NOR2_X1 U12492 ( .A1(n13929), .A2(n15425), .ZN(n13924) );
  NOR2_X1 U12493 ( .A1(n13772), .A2(n19068), .ZN(n13773) );
  NOR2_X1 U12494 ( .A1(n13925), .A2(n16261), .ZN(n13926) );
  NOR2_X1 U12495 ( .A1(n13771), .A2(n9649), .ZN(n13911) );
  AND2_X1 U12496 ( .A1(n13671), .A2(n9960), .ZN(n9693) );
  AND2_X1 U12497 ( .A1(n14039), .A2(n9965), .ZN(n9694) );
  INV_X1 U12498 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19762) );
  AND2_X1 U12499 ( .A1(n9899), .A2(n14051), .ZN(n9695) );
  NAND2_X1 U12500 ( .A1(n14191), .A2(n14199), .ZN(n14198) );
  NAND2_X1 U12501 ( .A1(n12762), .A2(n12761), .ZN(n15032) );
  AND2_X1 U12502 ( .A1(n11171), .A2(n9961), .ZN(n9696) );
  NAND2_X1 U12503 ( .A1(n14040), .A2(n14039), .ZN(n14038) );
  AND2_X1 U12504 ( .A1(n14844), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9697) );
  NAND2_X1 U12505 ( .A1(n9819), .A2(n10997), .ZN(n14096) );
  AND2_X1 U12506 ( .A1(n10060), .A2(n12223), .ZN(n9698) );
  OR2_X1 U12507 ( .A1(n13932), .A2(n11036), .ZN(n9699) );
  AND2_X1 U12508 ( .A1(n9651), .A2(n9773), .ZN(n12899) );
  AND2_X1 U12509 ( .A1(n9694), .A2(n9964), .ZN(n9700) );
  AND2_X1 U12510 ( .A1(n11215), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9701) );
  INV_X1 U12511 ( .A(n12921), .ZN(n12939) );
  INV_X1 U12512 ( .A(n12949), .ZN(n12921) );
  AND3_X1 U12513 ( .A1(n9689), .A2(n17673), .A3(n17714), .ZN(n16526) );
  NOR2_X1 U12514 ( .A1(n15174), .A2(n15173), .ZN(n15162) );
  OR2_X1 U12515 ( .A1(n17574), .A2(n9935), .ZN(n9702) );
  AND2_X1 U12516 ( .A1(n14863), .A2(n14697), .ZN(n9703) );
  AND2_X1 U12517 ( .A1(n15323), .A2(n9699), .ZN(n9704) );
  AND2_X1 U12518 ( .A1(n9982), .A2(n14417), .ZN(n9705) );
  AND2_X1 U12519 ( .A1(n9922), .A2(n9921), .ZN(n9706) );
  AND2_X1 U12520 ( .A1(n12222), .A2(n12221), .ZN(n13524) );
  OR2_X1 U12521 ( .A1(n10223), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9707) );
  INV_X1 U12522 ( .A(n9912), .ZN(n14392) );
  NOR2_X1 U12523 ( .A1(n9979), .A2(n9977), .ZN(n9708) );
  AND2_X1 U12524 ( .A1(n10215), .A2(n9857), .ZN(n9709) );
  AND2_X1 U12525 ( .A1(n9695), .A2(n9901), .ZN(n9710) );
  INV_X1 U12526 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15364) );
  INV_X1 U12527 ( .A(n11602), .ZN(n11541) );
  INV_X1 U12528 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19735) );
  AND2_X1 U12529 ( .A1(n15435), .A2(n15433), .ZN(n9711) );
  INV_X1 U12530 ( .A(n9877), .ZN(n9876) );
  NAND2_X1 U12531 ( .A1(n10965), .A2(n10964), .ZN(n9877) );
  NAND2_X1 U12532 ( .A1(n14978), .A2(n9892), .ZN(n9712) );
  AND2_X1 U12533 ( .A1(n14841), .A2(n14746), .ZN(n9713) );
  AND2_X1 U12534 ( .A1(n9925), .A2(n9924), .ZN(n9714) );
  AND2_X1 U12535 ( .A1(n10040), .A2(n10039), .ZN(n9715) );
  AND2_X1 U12536 ( .A1(n9895), .A2(n13946), .ZN(n9716) );
  AND2_X1 U12537 ( .A1(n9700), .A2(n14188), .ZN(n9717) );
  AND2_X1 U12538 ( .A1(n9693), .A2(n9959), .ZN(n9718) );
  AND2_X1 U12539 ( .A1(n9653), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9719) );
  INV_X1 U12540 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n20747) );
  INV_X1 U12541 ( .A(n13481), .ZN(n19934) );
  INV_X1 U12542 ( .A(n11731), .ZN(n9971) );
  NAND2_X1 U12543 ( .A1(n13243), .A2(n13242), .ZN(n13241) );
  AND2_X1 U12544 ( .A1(n14901), .A2(n9719), .ZN(n14895) );
  NAND2_X1 U12545 ( .A1(n14917), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14918) );
  AND2_X1 U12546 ( .A1(n15189), .A2(n15004), .ZN(n9720) );
  OR2_X1 U12547 ( .A1(n12610), .A2(n12609), .ZN(n9721) );
  AND2_X1 U12548 ( .A1(n9958), .A2(n9679), .ZN(n13373) );
  AND2_X1 U12549 ( .A1(n9892), .A2(n9891), .ZN(n9722) );
  INV_X1 U12550 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11226) );
  AND2_X1 U12551 ( .A1(n14199), .A2(n10062), .ZN(n9723) );
  NAND2_X1 U12552 ( .A1(n14911), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14916) );
  AND2_X1 U12553 ( .A1(n9678), .A2(n13250), .ZN(n9724) );
  AND2_X1 U12554 ( .A1(n13899), .A2(n12291), .ZN(n14042) );
  OR2_X1 U12555 ( .A1(n19130), .A2(n13370), .ZN(n9725) );
  NOR2_X1 U12556 ( .A1(n13418), .A2(n13417), .ZN(n11136) );
  NAND2_X1 U12557 ( .A1(n9919), .A2(n9918), .ZN(n9920) );
  NOR2_X1 U12558 ( .A1(n9974), .A2(n9972), .ZN(n9726) );
  AND2_X1 U12559 ( .A1(n13415), .A2(n9698), .ZN(n9727) );
  AND2_X1 U12560 ( .A1(n13415), .A2(n13416), .ZN(n9728) );
  AND2_X1 U12561 ( .A1(n9660), .A2(n10061), .ZN(n9729) );
  AND2_X1 U12562 ( .A1(n9961), .A2(n15101), .ZN(n9730) );
  AND2_X1 U12563 ( .A1(n9720), .A2(n9888), .ZN(n9731) );
  INV_X1 U12564 ( .A(n13290), .ZN(n9769) );
  AND2_X1 U12565 ( .A1(n17487), .A2(n9943), .ZN(n9732) );
  INV_X1 U12566 ( .A(n9775), .ZN(n12916) );
  INV_X2 U12567 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13699) );
  NOR2_X1 U12568 ( .A1(n10326), .A2(n10325), .ZN(n18600) );
  AND2_X1 U12569 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n9733)
         );
  NAND2_X1 U12570 ( .A1(n12953), .A2(n12952), .ZN(n9734) );
  INV_X1 U12571 ( .A(n14524), .ZN(n9978) );
  INV_X1 U12572 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n9871) );
  INV_X1 U12573 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17679) );
  AND2_X1 U12574 ( .A1(n9885), .A2(n9884), .ZN(n9735) );
  AND2_X1 U12575 ( .A1(n9878), .A2(n16204), .ZN(n9736) );
  INV_X1 U12576 ( .A(n9886), .ZN(n9885) );
  NAND2_X1 U12577 ( .A1(n14932), .A2(n12798), .ZN(n9886) );
  NOR2_X1 U12578 ( .A1(n20384), .A2(n20209), .ZN(n9737) );
  NOR2_X1 U12579 ( .A1(n20384), .A2(n20492), .ZN(n9738) );
  INV_X1 U12580 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n9879) );
  INV_X1 U12581 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9944) );
  INV_X1 U12582 ( .A(n17324), .ZN(n9841) );
  AND3_X1 U12583 ( .A1(n17673), .A2(n17714), .A3(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17634) );
  INV_X2 U12584 ( .A(n12619), .ZN(n10488) );
  INV_X1 U12585 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17818) );
  OR2_X1 U12586 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9739) );
  INV_X1 U12587 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n9951) );
  AND2_X1 U12588 ( .A1(n9953), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9740) );
  AND2_X1 U12589 ( .A1(n9666), .A2(n15608), .ZN(n9741) );
  INV_X1 U12590 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n9906) );
  INV_X1 U12591 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n9908) );
  INV_X1 U12592 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12617) );
  AND2_X1 U12593 ( .A1(n9667), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9742) );
  NOR2_X4 U12594 ( .A1(n20575), .A2(n20676), .ZN(n20621) );
  NOR2_X4 U12595 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13590) );
  NAND2_X1 U12596 ( .A1(n16054), .A2(n12854), .ZN(n16049) );
  NAND2_X1 U12597 ( .A1(n10026), .A2(n9745), .ZN(n9744) );
  NAND2_X1 U12598 ( .A1(n9747), .A2(n10026), .ZN(n9746) );
  INV_X1 U12599 ( .A(n16054), .ZN(n9747) );
  NAND3_X1 U12600 ( .A1(n10013), .A2(n10012), .A3(n16055), .ZN(n16054) );
  NAND2_X2 U12601 ( .A1(n9748), .A2(n12828), .ZN(n12836) );
  NOR2_X2 U12602 ( .A1(n13503), .A2(n13504), .ZN(n13502) );
  NAND2_X1 U12603 ( .A1(n9688), .A2(n9750), .ZN(n9780) );
  OR2_X1 U12604 ( .A1(n11576), .A2(n9751), .ZN(n13654) );
  NOR2_X1 U12605 ( .A1(n13262), .A2(n13261), .ZN(n9751) );
  INV_X1 U12606 ( .A(n11576), .ZN(n9752) );
  AND2_X2 U12607 ( .A1(n13262), .A2(n13261), .ZN(n11576) );
  NAND3_X1 U12608 ( .A1(n11378), .A2(n11398), .A3(n20044), .ZN(n11403) );
  NAND2_X1 U12609 ( .A1(n12921), .A2(n9755), .ZN(n9753) );
  NOR2_X1 U12610 ( .A1(n9755), .A2(n11374), .ZN(n9754) );
  NAND2_X1 U12611 ( .A1(n9784), .A2(n9760), .ZN(n9759) );
  NAND2_X1 U12612 ( .A1(n14000), .A2(n14009), .ZN(n14007) );
  OAI21_X1 U12613 ( .B1(n14755), .B2(n16035), .A(n9761), .ZN(P1_U2969) );
  AOI21_X1 U12614 ( .B1(n14586), .B2(n14671), .A(n14585), .ZN(n9761) );
  AND2_X2 U12615 ( .A1(n14477), .A2(n14479), .ZN(n14478) );
  XNOR2_X2 U12616 ( .A(n12807), .B(n11459), .ZN(n11558) );
  AND2_X2 U12617 ( .A1(n11232), .A2(n9763), .ZN(n11995) );
  AND2_X2 U12618 ( .A1(n11226), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9763) );
  XNOR2_X1 U12619 ( .A(n11551), .B(n9764), .ZN(n12822) );
  INV_X1 U12620 ( .A(n11586), .ZN(n11517) );
  INV_X1 U12621 ( .A(n9770), .ZN(n11394) );
  NAND4_X1 U12622 ( .A1(n11320), .A2(n11319), .A3(n11318), .A4(n11393), .ZN(
        n9770) );
  NAND2_X1 U12623 ( .A1(n11393), .A2(n11318), .ZN(n9774) );
  NAND4_X1 U12624 ( .A1(n12915), .A2(n9777), .A3(n9775), .A4(n12048), .ZN(
        n11365) );
  NAND2_X1 U12625 ( .A1(n13028), .A2(n12897), .ZN(n9777) );
  NAND2_X1 U12626 ( .A1(n13028), .A2(n11367), .ZN(n12915) );
  INV_X1 U12627 ( .A(n20124), .ZN(n9781) );
  INV_X1 U12628 ( .A(n13679), .ZN(n9784) );
  NAND2_X1 U12629 ( .A1(n17727), .A2(n10207), .ZN(n10214) );
  AND2_X1 U12630 ( .A1(n17769), .A2(n9789), .ZN(n9787) );
  NAND2_X1 U12631 ( .A1(n9788), .A2(n9787), .ZN(n17767) );
  OR2_X1 U12632 ( .A1(n17781), .A2(n17780), .ZN(n10047) );
  NAND2_X1 U12633 ( .A1(n9790), .A2(n18110), .ZN(n9789) );
  INV_X1 U12634 ( .A(n17780), .ZN(n9790) );
  NAND2_X1 U12635 ( .A1(n17781), .A2(n17780), .ZN(n17779) );
  OR2_X2 U12636 ( .A1(n10150), .A2(n10151), .ZN(n17339) );
  INV_X1 U12637 ( .A(n9795), .ZN(n10227) );
  NAND2_X1 U12638 ( .A1(n20124), .A2(n11408), .ZN(n20064) );
  XNOR2_X2 U12639 ( .A(n9796), .B(n11390), .ZN(n20124) );
  OAI21_X1 U12640 ( .B1(n14593), .B2(n16126), .A(n9812), .ZN(P1_U3002) );
  XNOR2_X1 U12641 ( .A(n9813), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14593) );
  OAI21_X1 U12642 ( .B1(n14841), .B2(n14311), .A(n9683), .ZN(n9813) );
  NAND2_X2 U12643 ( .A1(n10615), .A2(n10614), .ZN(n9816) );
  NAND2_X1 U12644 ( .A1(n10618), .A2(n9816), .ZN(n9815) );
  XNOR2_X2 U12645 ( .A(n10621), .B(n9816), .ZN(n12141) );
  NAND2_X1 U12646 ( .A1(n9990), .A2(n9817), .ZN(n11013) );
  NAND2_X1 U12647 ( .A1(n9818), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11003) );
  NAND2_X1 U12648 ( .A1(n14028), .A2(n14029), .ZN(n9819) );
  NAND2_X1 U12649 ( .A1(n10586), .A2(n9820), .ZN(n10589) );
  NAND4_X1 U12650 ( .A1(n9821), .A2(n9690), .A3(n10578), .A4(n9822), .ZN(n9820) );
  NAND3_X1 U12651 ( .A1(n9832), .A2(n15323), .A3(n9699), .ZN(n9831) );
  NAND2_X1 U12652 ( .A1(n9996), .A2(n9997), .ZN(n9837) );
  NOR2_X2 U12653 ( .A1(n10179), .A2(n17328), .ZN(n10178) );
  INV_X2 U12654 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18784) );
  NAND2_X1 U12655 ( .A1(n9847), .A2(n9845), .ZN(n16380) );
  INV_X1 U12656 ( .A(n9848), .ZN(n9847) );
  AOI21_X1 U12657 ( .B1(n9853), .B2(n9851), .A(n9849), .ZN(n9848) );
  AND2_X1 U12658 ( .A1(n17477), .A2(n17722), .ZN(n9854) );
  OAI21_X1 U12659 ( .B1(n14594), .B2(n14596), .A(n14841), .ZN(n14617) );
  NAND3_X1 U12660 ( .A1(n14625), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n9860), .ZN(n14608) );
  NAND2_X1 U12661 ( .A1(n14594), .A2(n14595), .ZN(n9860) );
  NAND2_X1 U12662 ( .A1(n14717), .A2(n9865), .ZN(n9867) );
  NAND2_X1 U12663 ( .A1(n14841), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9868) );
  INV_X1 U12664 ( .A(n11000), .ZN(n9869) );
  NAND2_X1 U12665 ( .A1(n11000), .A2(n9872), .ZN(n11015) );
  NAND2_X1 U12666 ( .A1(n11093), .A2(n9878), .ZN(n11105) );
  NAND2_X1 U12667 ( .A1(n11093), .A2(n9736), .ZN(n10966) );
  NAND2_X1 U12668 ( .A1(n11093), .A2(n15090), .ZN(n11104) );
  INV_X1 U12669 ( .A(n10966), .ZN(n14946) );
  AOI21_X1 U12670 ( .B1(n15490), .B2(n16250), .A(n9880), .ZN(n9954) );
  XNOR2_X1 U12671 ( .A(n15234), .B(n15231), .ZN(n15490) );
  AND2_X1 U12672 ( .A1(n15136), .A2(n14932), .ZN(n14934) );
  NAND2_X1 U12673 ( .A1(n15136), .A2(n9885), .ZN(n15449) );
  NAND3_X1 U12674 ( .A1(n9883), .A2(n9882), .A3(n9881), .ZN(n16174) );
  NAND2_X1 U12675 ( .A1(n9886), .A2(n15448), .ZN(n9881) );
  NAND2_X1 U12676 ( .A1(n15136), .A2(n9735), .ZN(n9882) );
  OR2_X1 U12677 ( .A1(n15136), .A2(n9884), .ZN(n9883) );
  INV_X1 U12678 ( .A(n15448), .ZN(n9884) );
  NAND2_X1 U12679 ( .A1(n9887), .A2(n15454), .ZN(n15473) );
  OR2_X1 U12680 ( .A1(n16174), .A2(n16305), .ZN(n9887) );
  NAND2_X1 U12681 ( .A1(n15006), .A2(n9731), .ZN(n15174) );
  AND2_X2 U12682 ( .A1(n14978), .A2(n9889), .ZN(n15134) );
  INV_X1 U12683 ( .A(n13917), .ZN(n9894) );
  NAND2_X1 U12684 ( .A1(n9894), .A2(n9716), .ZN(n13947) );
  NAND2_X2 U12685 ( .A1(n12762), .A2(n9710), .ZN(n15197) );
  AND2_X4 U12686 ( .A1(n13770), .A2(n13769), .ZN(n18893) );
  NAND2_X1 U12687 ( .A1(n13770), .A2(n9902), .ZN(n15030) );
  INV_X1 U12688 ( .A(n13769), .ZN(n9903) );
  INV_X1 U12689 ( .A(n13771), .ZN(n9904) );
  NAND2_X1 U12690 ( .A1(n9905), .A2(n9904), .ZN(n13925) );
  NOR2_X2 U12691 ( .A1(n14378), .A2(n14363), .ZN(n14362) );
  INV_X1 U12692 ( .A(n9920), .ZN(n16139) );
  NAND4_X1 U12693 ( .A1(n17673), .A2(n17714), .A3(n16694), .A4(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17610) );
  AOI21_X1 U12694 ( .B1(n16585), .B2(n17479), .A(n16837), .ZN(n16564) );
  INV_X1 U12695 ( .A(n9946), .ZN(n16572) );
  NOR2_X2 U12696 ( .A1(n10658), .A2(n13728), .ZN(n19290) );
  OR2_X2 U12697 ( .A1(n10634), .A2(n9947), .ZN(n10658) );
  INV_X1 U12698 ( .A(n12157), .ZN(n9948) );
  AND2_X2 U12699 ( .A1(n9600), .A2(n9741), .ZN(n15288) );
  AND2_X2 U12700 ( .A1(n15265), .A2(n9742), .ZN(n15250) );
  NAND2_X2 U12701 ( .A1(n15439), .A2(n10911), .ZN(n16264) );
  NAND2_X2 U12702 ( .A1(n15250), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15230) );
  NAND2_X1 U12703 ( .A1(n11171), .A2(n9730), .ZN(n15096) );
  INV_X1 U12704 ( .A(n11171), .ZN(n14195) );
  INV_X1 U12705 ( .A(n15115), .ZN(n9963) );
  NAND2_X1 U12706 ( .A1(n14040), .A2(n9717), .ZN(n14187) );
  NAND2_X1 U12707 ( .A1(n14974), .A2(n9966), .ZN(n15063) );
  OAI21_X1 U12708 ( .B1(n12822), .B2(n11555), .A(n9969), .ZN(n13458) );
  NOR2_X1 U12709 ( .A1(n14373), .A2(n14375), .ZN(n14374) );
  NOR3_X1 U12710 ( .A1(n14373), .A2(n14351), .A3(n9987), .ZN(n14350) );
  NAND2_X2 U12711 ( .A1(n10670), .A2(n13699), .ZN(n12530) );
  OAI21_X1 U12712 ( .B1(n15418), .B2(n11083), .A(n11082), .ZN(n15313) );
  INV_X1 U12713 ( .A(n15314), .ZN(n9995) );
  NAND2_X1 U12714 ( .A1(n15243), .A2(n9999), .ZN(n9996) );
  NOR2_X4 U12715 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13575) );
  NAND2_X1 U12716 ( .A1(n13538), .A2(n10011), .ZN(n10013) );
  INV_X1 U12717 ( .A(n12837), .ZN(n10016) );
  OAI21_X1 U12718 ( .B1(n13538), .B2(n9590), .A(n10014), .ZN(n16056) );
  AOI21_X1 U12719 ( .B1(n10016), .B2(n19964), .A(n10015), .ZN(n10014) );
  NAND2_X1 U12720 ( .A1(n19965), .A2(n19964), .ZN(n19963) );
  NAND2_X1 U12721 ( .A1(n10020), .A2(n9713), .ZN(n14314) );
  INV_X1 U12722 ( .A(n14607), .ZN(n10022) );
  INV_X1 U12723 ( .A(n16045), .ZN(n10027) );
  AOI21_X1 U12724 ( .B1(n10025), .B2(n16045), .A(n10028), .ZN(n10024) );
  NAND2_X1 U12725 ( .A1(n10030), .A2(n12864), .ZN(n16043) );
  NAND2_X1 U12726 ( .A1(n16049), .A2(n12862), .ZN(n10030) );
  NAND2_X1 U12727 ( .A1(n14693), .A2(n10034), .ZN(n10033) );
  AND2_X1 U12728 ( .A1(n17515), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10045) );
  NAND2_X1 U12729 ( .A1(n17515), .A2(n10223), .ZN(n10040) );
  OAI21_X1 U12730 ( .B1(n17845), .B2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n17833), .ZN(n10042) );
  NOR2_X2 U12731 ( .A1(n18015), .A2(n10215), .ZN(n18059) );
  NAND3_X1 U12732 ( .A1(n10055), .A2(n10073), .A3(n10049), .ZN(n10353) );
  NAND3_X1 U12733 ( .A1(n10133), .A2(n10052), .A3(n10051), .ZN(n10050) );
  NOR2_X2 U12734 ( .A1(n15795), .A2(n16359), .ZN(n15851) );
  INV_X2 U12735 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18778) );
  AND2_X2 U12736 ( .A1(n14191), .A2(n9729), .ZN(n15104) );
  XNOR2_X1 U12737 ( .A(n12546), .B(n10074), .ZN(n15077) );
  NAND2_X2 U12738 ( .A1(n12168), .A2(n12167), .ZN(n13243) );
  NAND2_X1 U12739 ( .A1(n13899), .A2(n10069), .ZN(n14048) );
  INV_X1 U12740 ( .A(n14048), .ZN(n12335) );
  AND2_X2 U12741 ( .A1(n10070), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10672) );
  INV_X1 U12742 ( .A(n13611), .ZN(n11593) );
  NAND2_X1 U12743 ( .A1(n13924), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14899) );
  AOI21_X1 U12744 ( .B1(n12822), .B2(n12865), .A(n12826), .ZN(n13503) );
  OR2_X2 U12745 ( .A1(n10624), .A2(n13412), .ZN(n19136) );
  INV_X1 U12746 ( .A(n13612), .ZN(n11594) );
  INV_X1 U12747 ( .A(n15441), .ZN(n10910) );
  NAND2_X1 U12748 ( .A1(n15092), .A2(n15095), .ZN(n15093) );
  XNOR2_X1 U12749 ( .A(n15104), .B(n12498), .ZN(n15092) );
  XNOR2_X2 U12750 ( .A(n12836), .B(n12829), .ZN(n13540) );
  INV_X1 U12751 ( .A(n12949), .ZN(n11369) );
  OR2_X1 U12752 ( .A1(n11380), .A2(n12917), .ZN(n11378) );
  NAND2_X1 U12753 ( .A1(n11380), .A2(n11371), .ZN(n11393) );
  NAND2_X2 U12754 ( .A1(n11371), .A2(n11367), .ZN(n12949) );
  NAND2_X1 U12755 ( .A1(n13864), .A2(n15240), .ZN(n10981) );
  NAND2_X1 U12756 ( .A1(n14331), .A2(n12116), .ZN(n12134) );
  AOI22_X1 U12757 ( .A1(n9629), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10435) );
  NAND2_X1 U12758 ( .A1(n10463), .A2(n10430), .ZN(n10470) );
  INV_X1 U12759 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n19726) );
  INV_X1 U12760 ( .A(n14389), .ZN(n14406) );
  NOR2_X1 U12761 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11574) );
  NAND2_X2 U12762 ( .A1(n14571), .A2(n13291), .ZN(n15997) );
  OR2_X1 U12763 ( .A1(n15877), .A2(n15876), .ZN(n10071) );
  AND4_X1 U12764 ( .A1(n10829), .A2(n10828), .A3(n10827), .A4(n10826), .ZN(
        n10072) );
  AND3_X1 U12765 ( .A1(n10136), .A2(n10135), .A3(n10134), .ZN(n10073) );
  AND2_X1 U12766 ( .A1(n12565), .A2(n12544), .ZN(n10074) );
  INV_X1 U12767 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19097) );
  OR2_X1 U12768 ( .A1(n14460), .A2(n20017), .ZN(n10075) );
  NOR2_X1 U12769 ( .A1(n14684), .A2(n14477), .ZN(n10076) );
  AND2_X1 U12770 ( .A1(n10514), .A2(n10513), .ZN(n10077) );
  AND4_X1 U12771 ( .A1(n10688), .A2(n10687), .A3(n10686), .A4(n10685), .ZN(
        n10078) );
  INV_X1 U12772 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15523) );
  INV_X1 U12773 ( .A(n10610), .ZN(n11126) );
  NAND2_X1 U12774 ( .A1(n9618), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12652) );
  AND2_X1 U12775 ( .A1(n10473), .A2(n10472), .ZN(n10079) );
  INV_X1 U12776 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14455) );
  NOR2_X1 U12777 ( .A1(n20384), .A2(n20355), .ZN(n10080) );
  NOR2_X1 U12778 ( .A1(n20384), .A2(n20123), .ZN(n10081) );
  AND2_X2 U12779 ( .A1(n13263), .A2(n20503), .ZN(n14671) );
  INV_X2 U12780 ( .A(n19901), .ZN(n19930) );
  INV_X1 U12781 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16541) );
  AND2_X1 U12782 ( .A1(n19290), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10082) );
  AND3_X1 U12783 ( .A1(n10475), .A2(n10430), .A3(n10474), .ZN(n10083) );
  INV_X1 U12784 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13370) );
  INV_X2 U12785 ( .A(n17352), .ZN(n17394) );
  INV_X1 U12786 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19633) );
  INV_X1 U12787 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11216) );
  AND2_X1 U12788 ( .A1(n10883), .A2(n10998), .ZN(n10084) );
  AND2_X1 U12789 ( .A1(n15270), .A2(n15276), .ZN(n10085) );
  NAND2_X1 U12790 ( .A1(n20556), .A2(n20023), .ZN(n20066) );
  AND2_X1 U12791 ( .A1(n10675), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10086) );
  AND4_X1 U12792 ( .A1(n10718), .A2(n10717), .A3(n10716), .A4(n10715), .ZN(
        n10087) );
  AND3_X1 U12793 ( .A1(n10510), .A2(n10509), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10088) );
  NAND2_X1 U12794 ( .A1(n13344), .A2(n13327), .ZN(n16305) );
  INV_X1 U12795 ( .A(n16305), .ZN(n15739) );
  INV_X1 U12796 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n18896) );
  INV_X1 U12797 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19725) );
  INV_X1 U12798 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n15112) );
  INV_X1 U12799 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10914) );
  INV_X2 U12800 ( .A(n18818), .ZN(n18817) );
  NOR2_X1 U12801 ( .A1(n18612), .A2(n10103), .ZN(n10137) );
  INV_X1 U12802 ( .A(n15636), .ZN(n10913) );
  INV_X2 U12803 ( .A(n19777), .ZN(n19776) );
  AND2_X1 U12804 ( .A1(n20564), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20666) );
  INV_X1 U12805 ( .A(n20666), .ZN(n20676) );
  INV_X1 U12806 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n11362) );
  INV_X1 U12807 ( .A(n15479), .ZN(n15487) );
  NAND2_X1 U12808 ( .A1(n15449), .A2(n12799), .ZN(n15479) );
  INV_X1 U12809 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20417) );
  INV_X1 U12810 ( .A(n10100), .ZN(n10287) );
  NOR2_X2 U12811 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20641) );
  AND4_X1 U12812 ( .A1(n15497), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n15470), .ZN(n10090) );
  NOR2_X1 U12813 ( .A1(n10102), .A2(n18635), .ZN(n10279) );
  INV_X1 U12814 ( .A(n10676), .ZN(n12412) );
  INV_X1 U12815 ( .A(n10714), .ZN(n10899) );
  INV_X1 U12816 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19737) );
  INV_X1 U12817 ( .A(n13328), .ZN(n18925) );
  AND2_X1 U12818 ( .A1(n13749), .A2(n19520), .ZN(n13328) );
  NAND4_X1 U12819 ( .A1(n15335), .A2(n11078), .A3(n15348), .A4(n15405), .ZN(
        n10092) );
  OR2_X1 U12820 ( .A1(n12078), .A2(n12077), .ZN(n12085) );
  AND2_X1 U12821 ( .A1(n19169), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10638) );
  AOI211_X1 U12822 ( .C1(n12090), .C2(n12089), .A(n12088), .B(n12087), .ZN(
        n12102) );
  AOI22_X1 U12823 ( .A1(n10675), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9629), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10467) );
  AOI22_X1 U12824 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19409), .B1(
        n19356), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10660) );
  BUF_X1 U12825 ( .A(n11688), .Z(n11994) );
  OR2_X1 U12826 ( .A1(n11527), .A2(n11526), .ZN(n12857) );
  AND2_X1 U12827 ( .A1(n10538), .A2(n19103), .ZN(n10532) );
  OAI21_X1 U12828 ( .B1(n10523), .B2(n10553), .A(n10554), .ZN(n10522) );
  AOI22_X1 U12829 ( .A1(n9630), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10441) );
  INV_X1 U12830 ( .A(n12073), .ZN(n12063) );
  INV_X1 U12831 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11225) );
  INV_X1 U12832 ( .A(n12876), .ZN(n11439) );
  OR2_X1 U12833 ( .A1(n11540), .A2(n11539), .ZN(n12868) );
  AOI22_X1 U12834 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11239) );
  OR2_X1 U12835 ( .A1(n12807), .A2(n11460), .ZN(n11461) );
  AOI22_X1 U12836 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10422) );
  INV_X1 U12837 ( .A(n15332), .ZN(n11081) );
  NAND2_X1 U12838 ( .A1(n10691), .A2(n10690), .ZN(n10692) );
  AOI22_X1 U12839 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10515), .B1(
        n9630), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10447) );
  AOI21_X1 U12840 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n18156), .A(
        n10330), .ZN(n10331) );
  OR2_X1 U12841 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20019), .ZN(
        n12056) );
  INV_X1 U12842 ( .A(n14486), .ZN(n11787) );
  INV_X1 U12843 ( .A(n14506), .ZN(n11721) );
  INV_X1 U12844 ( .A(n14014), .ZN(n11626) );
  NOR2_X1 U12845 ( .A1(n11439), .A2(n11490), .ZN(n12804) );
  OR2_X1 U12846 ( .A1(n11479), .A2(n11478), .ZN(n12823) );
  INV_X1 U12847 ( .A(n13524), .ZN(n12223) );
  INV_X1 U12848 ( .A(n14184), .ZN(n12334) );
  NAND2_X1 U12849 ( .A1(n12684), .A2(n12683), .ZN(n12706) );
  NOR2_X1 U12850 ( .A1(n10092), .A2(n11081), .ZN(n11082) );
  INV_X1 U12851 ( .A(n10723), .ZN(n10768) );
  NAND2_X1 U12852 ( .A1(n9613), .A2(n13412), .ZN(n10727) );
  NAND2_X1 U12853 ( .A1(n10456), .A2(n10455), .ZN(n10457) );
  AOI21_X1 U12854 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18623), .A(
        n10327), .ZN(n10329) );
  NAND2_X1 U12855 ( .A1(n18762), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10228) );
  NOR2_X1 U12856 ( .A1(n12071), .A2(n12817), .ZN(n12100) );
  INV_X1 U12857 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14380) );
  AND2_X1 U12858 ( .A1(n11910), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11911) );
  INV_X1 U12859 ( .A(n11548), .ZN(n11549) );
  INV_X1 U12860 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n12008) );
  NOR2_X1 U12861 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12895) );
  OR2_X1 U12862 ( .A1(n11451), .A2(n11450), .ZN(n12814) );
  INV_X1 U12863 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13977) );
  AND2_X1 U12864 ( .A1(n12473), .A2(n12472), .ZN(n12494) );
  INV_X1 U12865 ( .A(n10777), .ZN(n12424) );
  AOI21_X1 U12866 ( .B1(n15483), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n15482), .ZN(n15484) );
  AND2_X1 U12867 ( .A1(n12788), .A2(n12787), .ZN(n15146) );
  NAND2_X1 U12868 ( .A1(n12655), .A2(n13330), .ZN(n10587) );
  NOR2_X2 U12869 ( .A1(n10622), .A2(n12141), .ZN(n10807) );
  NOR2_X1 U12870 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18784), .ZN(
        n10333) );
  INV_X1 U12871 ( .A(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n20713) );
  INV_X1 U12872 ( .A(n10414), .ZN(n10229) );
  OR2_X1 U12873 ( .A1(n11952), .A2(n14380), .ZN(n11989) );
  OR2_X1 U12874 ( .A1(n14645), .A2(n12014), .ZN(n11889) );
  NOR2_X1 U12875 ( .A1(n11789), .A2(n15926), .ZN(n11790) );
  NOR2_X2 U12876 ( .A1(n12045), .A2(n12008), .ZN(n11731) );
  OAI211_X1 U12877 ( .C1(n12071), .C2(n11458), .A(n11457), .B(n11456), .ZN(
        n11564) );
  NOR2_X1 U12878 ( .A1(n20645), .A2(n20273), .ZN(n20356) );
  NOR2_X1 U12879 ( .A1(n13568), .A2(n20387), .ZN(n20491) );
  AND2_X1 U12880 ( .A1(n10538), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19764) );
  INV_X1 U12881 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14952) );
  INV_X1 U12882 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14922) );
  OR2_X1 U12883 ( .A1(n12372), .A2(n12371), .ZN(n14199) );
  NOR2_X2 U12884 ( .A1(n14916), .A2(n15303), .ZN(n14917) );
  AND2_X1 U12885 ( .A1(n12772), .A2(n12771), .ZN(n15196) );
  INV_X1 U12886 ( .A(n10615), .ZN(n10616) );
  INV_X1 U12887 ( .A(n18674), .ZN(n18803) );
  INV_X1 U12888 ( .A(n10415), .ZN(n10416) );
  NOR4_X1 U12889 ( .A1(n18185), .A2(n10390), .A3(n10320), .A4(n10389), .ZN(
        n18607) );
  INV_X1 U12890 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14336) );
  AND2_X1 U12891 ( .A1(n13007), .A2(n13006), .ZN(n14472) );
  AND2_X1 U12892 ( .A1(n11740), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11758) );
  INV_X1 U12893 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19809) );
  INV_X1 U12894 ( .A(n19876), .ZN(n19867) );
  NAND2_X1 U12895 ( .A1(n11489), .A2(n11488), .ZN(n20157) );
  NAND2_X1 U12896 ( .A1(n11860), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11909) );
  INV_X1 U12897 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15903) );
  NAND2_X1 U12898 ( .A1(n11758), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11771) );
  AND2_X1 U12899 ( .A1(n11731), .A2(n11672), .ZN(n14524) );
  AND3_X1 U12900 ( .A1(n12963), .A2(n12990), .A3(n12962), .ZN(n14132) );
  NOR2_X1 U12901 ( .A1(n16093), .A2(n19994), .ZN(n20008) );
  OR2_X1 U12902 ( .A1(n13403), .A2(n13399), .ZN(n16093) );
  INV_X1 U12903 ( .A(n20066), .ZN(n20162) );
  OR2_X1 U12904 ( .A1(n20642), .A2(n20268), .ZN(n20127) );
  INV_X1 U12905 ( .A(n20154), .ZN(n20155) );
  AND2_X1 U12906 ( .A1(n20444), .A2(n20162), .ZN(n20328) );
  OR2_X1 U12907 ( .A1(n20648), .A2(n20383), .ZN(n20385) );
  INV_X1 U12908 ( .A(n20641), .ZN(n20646) );
  AND2_X1 U12909 ( .A1(n20669), .A2(n20640), .ZN(n15835) );
  NOR2_X1 U12910 ( .A1(n19766), .A2(n19768), .ZN(n13779) );
  INV_X1 U12911 ( .A(n16184), .ZN(n16185) );
  INV_X1 U12912 ( .A(n14907), .ZN(n14897) );
  NAND2_X1 U12913 ( .A1(n15470), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13769) );
  AND2_X1 U12914 ( .A1(n10933), .A2(n10932), .ZN(n19747) );
  AND3_X1 U12915 ( .A1(n12739), .A2(n12738), .A3(n12737), .ZN(n13918) );
  INV_X1 U12916 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15282) );
  NOR2_X1 U12917 ( .A1(n10090), .A2(n15453), .ZN(n15454) );
  OR2_X1 U12918 ( .A1(n14935), .A2(n10971), .ZN(n15213) );
  AND2_X1 U12919 ( .A1(n15467), .A2(n15560), .ZN(n15536) );
  OR2_X1 U12920 ( .A1(n15690), .A2(n15451), .ZN(n15631) );
  INV_X1 U12921 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15610) );
  AND2_X1 U12922 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15692) );
  NAND2_X1 U12923 ( .A1(n12680), .A2(n9618), .ZN(n19761) );
  INV_X1 U12924 ( .A(n19228), .ZN(n19288) );
  OAI21_X2 U12925 ( .B1(n16320), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n13845), 
        .ZN(n19573) );
  AOI211_X1 U12926 ( .C1(n10347), .C2(n10346), .A(n10345), .B(n10344), .ZN(
        n18795) );
  NOR2_X1 U12927 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16654), .ZN(n16643) );
  NOR2_X1 U12928 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16678), .ZN(n16663) );
  NAND2_X1 U12929 ( .A1(n18823), .A2(n18161), .ZN(n16514) );
  INV_X1 U12930 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17056) );
  NAND2_X1 U12931 ( .A1(n18803), .A2(n15775), .ZN(n17348) );
  INV_X1 U12932 ( .A(n17724), .ZN(n16334) );
  INV_X1 U12933 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n20720) );
  INV_X1 U12934 ( .A(n17929), .ZN(n16341) );
  INV_X1 U12935 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17636) );
  NOR2_X1 U12936 ( .A1(n17596), .A2(n17609), .ZN(n17795) );
  NOR2_X1 U12937 ( .A1(n17605), .A2(n17897), .ZN(n17549) );
  INV_X1 U12938 ( .A(n17884), .ZN(n17962) );
  INV_X1 U12939 ( .A(n10216), .ZN(n10215) );
  INV_X1 U12940 ( .A(n18210), .ZN(n18253) );
  INV_X1 U12941 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18623) );
  INV_X1 U12942 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n20785) );
  AOI22_X1 U12943 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10297) );
  NAND2_X1 U12944 ( .A1(n11823), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11858) );
  NOR2_X1 U12945 ( .A1(n15904), .A2(n15986), .ZN(n15943) );
  AND2_X1 U12946 ( .A1(n19831), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13628) );
  AND2_X1 U12947 ( .A1(n13639), .A2(n13631), .ZN(n19875) );
  INV_X1 U12948 ( .A(n15982), .ZN(n19857) );
  INV_X1 U12949 ( .A(n19899), .ZN(n14510) );
  AND2_X1 U12950 ( .A1(n14571), .A2(n13292), .ZN(n14580) );
  INV_X1 U12951 ( .A(n13481), .ZN(n19954) );
  INV_X2 U12952 ( .A(n13466), .ZN(n19959) );
  AND2_X1 U12953 ( .A1(n9677), .A2(n14471), .ZN(n15889) );
  AND2_X1 U12954 ( .A1(n13610), .A2(n13613), .ZN(n19967) );
  AND2_X1 U12955 ( .A1(n13265), .A2(n13264), .ZN(n19968) );
  NAND2_X1 U12956 ( .A1(n14880), .A2(n20556), .ZN(n13266) );
  INV_X1 U12957 ( .A(n16126), .ZN(n20004) );
  NAND2_X1 U12958 ( .A1(n12914), .A2(n12913), .ZN(n13053) );
  INV_X1 U12959 ( .A(n15846), .ZN(n20633) );
  OAI22_X1 U12960 ( .A1(n20031), .A2(n20030), .B1(n20330), .B2(n20159), .ZN(
        n20060) );
  OAI22_X1 U12961 ( .A1(n20099), .A2(n20098), .B1(n20330), .B2(n20216), .ZN(
        n20117) );
  AND2_X1 U12962 ( .A1(n13601), .A2(n12818), .ZN(n20210) );
  INV_X1 U12963 ( .A(n20212), .ZN(n20234) );
  INV_X1 U12964 ( .A(n20267), .ZN(n20258) );
  INV_X1 U12965 ( .A(n20261), .ZN(n20295) );
  INV_X1 U12966 ( .A(n20156), .ZN(n20270) );
  INV_X1 U12967 ( .A(n20325), .ZN(n20348) );
  OAI22_X1 U12968 ( .A1(n20393), .A2(n20392), .B1(n20444), .B2(n20391), .ZN(
        n20408) );
  INV_X1 U12969 ( .A(n20385), .ZN(n20438) );
  OAI211_X1 U12970 ( .C1(n20481), .C2(n20451), .A(n20450), .B(n20449), .ZN(
        n20484) );
  INV_X1 U12971 ( .A(n20452), .ZN(n20549) );
  OR2_X1 U12972 ( .A1(n13227), .A2(n15859), .ZN(n15840) );
  INV_X1 U12973 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20564) );
  INV_X1 U12974 ( .A(n20623), .ZN(n20617) );
  NAND2_X1 U12975 ( .A1(n16186), .A2(n16185), .ZN(n16187) );
  NAND2_X1 U12976 ( .A1(n18861), .A2(n18893), .ZN(n14991) );
  NAND2_X1 U12977 ( .A1(n18886), .A2(n18893), .ZN(n15017) );
  INV_X1 U12978 ( .A(n18936), .ZN(n18923) );
  INV_X1 U12979 ( .A(n18940), .ZN(n18927) );
  AND2_X1 U12980 ( .A1(n11026), .A2(n11025), .ZN(n13943) );
  INV_X1 U12981 ( .A(n18925), .ZN(n18939) );
  INV_X1 U12982 ( .A(n18946), .ZN(n18902) );
  AND2_X1 U12983 ( .A1(n12290), .A2(n12289), .ZN(n13905) );
  CLKBUF_X1 U12984 ( .A(n15093), .Z(n15094) );
  AND2_X1 U12985 ( .A1(n13515), .A2(n13852), .ZN(n18957) );
  INV_X1 U12986 ( .A(n19739), .ZN(n19144) );
  OAI21_X1 U12987 ( .B1(n12687), .B2(n19756), .A(n13791), .ZN(n13094) );
  NOR2_X1 U12988 ( .A1(n13078), .A2(n13077), .ZN(n13791) );
  AND2_X1 U12989 ( .A1(n14195), .A2(n14197), .ZN(n15628) );
  INV_X1 U12990 ( .A(n19075), .ZN(n16251) );
  AND2_X1 U12991 ( .A1(n19067), .A2(n19070), .ZN(n19059) );
  AND2_X1 U12992 ( .A1(n14179), .A2(n14059), .ZN(n18885) );
  INV_X1 U12993 ( .A(n16306), .ZN(n16281) );
  INV_X1 U12994 ( .A(n16315), .ZN(n15757) );
  XNOR2_X1 U12995 ( .A(n13410), .B(n13411), .ZN(n19145) );
  INV_X1 U12996 ( .A(n19573), .ZN(n19523) );
  AND2_X1 U12997 ( .A1(n19145), .A2(n19739), .ZN(n19228) );
  AND2_X1 U12998 ( .A1(n19228), .A2(n19171), .ZN(n19221) );
  INV_X1 U12999 ( .A(n19254), .ZN(n19246) );
  OAI21_X1 U13000 ( .B1(n19262), .B2(n19261), .A(n19260), .ZN(n19282) );
  INV_X1 U13001 ( .A(n19315), .ZN(n19307) );
  INV_X1 U13002 ( .A(n19352), .ZN(n19355) );
  NAND2_X1 U13003 ( .A1(n19145), .A2(n19144), .ZN(n19327) );
  NOR2_X1 U13004 ( .A1(n19519), .A2(n19707), .ZN(n19433) );
  OAI21_X1 U13005 ( .B1(n13856), .B2(n13855), .A(n13854), .ZN(n19480) );
  NOR2_X2 U13006 ( .A1(n19519), .A2(n19493), .ZN(n19515) );
  INV_X1 U13007 ( .A(n19612), .ZN(n19550) );
  AND2_X1 U13008 ( .A1(n9622), .A2(n19124), .ZN(n19613) );
  OR3_X1 U13009 ( .A1(n13751), .A2(n13750), .A3(n19755), .ZN(n19625) );
  INV_X1 U13010 ( .A(n19756), .ZN(n19768) );
  INV_X1 U13011 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19649) );
  NOR2_X1 U13012 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16635), .ZN(n16623) );
  INV_X1 U13013 ( .A(n16687), .ZN(n16696) );
  NOR2_X1 U13014 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16700), .ZN(n16686) );
  INV_X1 U13015 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n20697) );
  NOR2_X1 U13016 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16760), .ZN(n16748) );
  NOR2_X2 U13017 ( .A1(n16511), .A2(n16514), .ZN(n16833) );
  NOR2_X2 U13018 ( .A1(n18752), .A2(n16877), .ZN(n16824) );
  INV_X1 U13019 ( .A(n16855), .ZN(n16877) );
  INV_X1 U13020 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16883) );
  INV_X1 U13021 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n20688) );
  NOR2_X1 U13022 ( .A1(n17056), .A2(n17170), .ZN(n17121) );
  AND2_X1 U13023 ( .A1(n14219), .A2(n17177), .ZN(n17171) );
  AOI21_X1 U13024 ( .B1(n14207), .B2(n14206), .A(n15780), .ZN(n15877) );
  INV_X1 U13025 ( .A(n17259), .ZN(n17255) );
  NAND2_X1 U13026 ( .A1(n18812), .A2(n18601), .ZN(n17398) );
  OR2_X1 U13027 ( .A1(n18805), .A2(n17397), .ZN(n17400) );
  NAND2_X1 U13028 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17472) );
  INV_X1 U13029 ( .A(n18167), .ZN(n18804) );
  AND2_X1 U13030 ( .A1(n17824), .A2(n15787), .ZN(n16377) );
  INV_X1 U13031 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17878) );
  INV_X1 U13032 ( .A(n17312), .ZN(n16375) );
  INV_X1 U13033 ( .A(n17947), .ZN(n18057) );
  NOR2_X1 U13034 ( .A1(n9846), .A2(n18127), .ZN(n18121) );
  NOR2_X1 U13035 ( .A1(n18796), .A2(n18143), .ZN(n18140) );
  INV_X1 U13036 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18781) );
  INV_X1 U13037 ( .A(n18765), .ZN(n18779) );
  INV_X2 U13038 ( .A(n18545), .ZN(n18507) );
  INV_X1 U13039 ( .A(n18343), .ZN(n18335) );
  INV_X1 U13040 ( .A(n18296), .ZN(n18363) );
  INV_X1 U13041 ( .A(n18383), .ZN(n18452) );
  NOR2_X1 U13042 ( .A1(n18623), .A2(n18410), .ZN(n18483) );
  INV_X1 U13043 ( .A(n18456), .ZN(n18533) );
  NOR2_X1 U13044 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18627) );
  INV_X1 U13045 ( .A(n18667), .ZN(n18807) );
  INV_X1 U13046 ( .A(n18814), .ZN(n18805) );
  INV_X1 U13047 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18677) );
  NOR2_X1 U13048 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13075), .ZN(n16468)
         );
  NAND2_X1 U13049 ( .A1(n13264), .A2(n13029), .ZN(n14325) );
  INV_X1 U13050 ( .A(n20666), .ZN(n20664) );
  NAND2_X1 U13051 ( .A1(n13626), .A2(n13628), .ZN(n15982) );
  INV_X1 U13052 ( .A(n19852), .ZN(n19892) );
  NAND2_X1 U13053 ( .A1(n19899), .A2(n9769), .ZN(n14532) );
  INV_X1 U13054 ( .A(n15889), .ZN(n14562) );
  INV_X1 U13055 ( .A(n15964), .ZN(n14576) );
  AND2_X1 U13056 ( .A1(n13486), .A2(n13485), .ZN(n20059) );
  AND2_X1 U13057 ( .A1(n13456), .A2(n13455), .ZN(n20027) );
  NAND2_X1 U13058 ( .A1(n19903), .A2(n11372), .ZN(n13436) );
  INV_X1 U13059 ( .A(n19903), .ZN(n19932) );
  NOR2_X1 U13060 ( .A1(n14325), .A2(n13295), .ZN(n13481) );
  AOI21_X1 U13061 ( .B1(n14331), .B2(n14671), .A(n14318), .ZN(n14319) );
  INV_X1 U13062 ( .A(n16032), .ZN(n19972) );
  INV_X1 U13063 ( .A(n14671), .ZN(n20022) );
  OR2_X1 U13064 ( .A1(n13266), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16122) );
  INV_X1 U13065 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20762) );
  INV_X1 U13066 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20274) );
  INV_X1 U13067 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16158) );
  NAND2_X1 U13068 ( .A1(n20122), .A2(n20270), .ZN(n20084) );
  NAND2_X1 U13069 ( .A1(n20122), .A2(n20413), .ZN(n20114) );
  NAND2_X1 U13070 ( .A1(n20122), .A2(n20210), .ZN(n20153) );
  NAND2_X1 U13071 ( .A1(n20122), .A2(n20121), .ZN(n20178) );
  OR2_X1 U13072 ( .A1(n20639), .A2(n20156), .ZN(n20208) );
  OR2_X1 U13073 ( .A1(n20639), .A2(n20303), .ZN(n20239) );
  OR2_X1 U13074 ( .A1(n20639), .A2(n20354), .ZN(n20261) );
  NAND2_X1 U13075 ( .A1(n20271), .A2(n20270), .ZN(n20323) );
  OR2_X1 U13076 ( .A1(n20647), .A2(n20303), .ZN(n20353) );
  OR2_X1 U13077 ( .A1(n20647), .A2(n20445), .ZN(n20376) );
  OR2_X1 U13078 ( .A1(n20647), .A2(n20354), .ZN(n20412) );
  NAND2_X1 U13079 ( .A1(n20414), .A2(n20413), .ZN(n20487) );
  OR2_X1 U13080 ( .A1(n20498), .A2(n20354), .ZN(n20553) );
  INV_X2 U13081 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20556) );
  INV_X1 U13082 ( .A(n20632), .ZN(n20560) );
  NAND2_X1 U13083 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20669) );
  INV_X1 U13084 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20586) );
  INV_X1 U13085 ( .A(n20621), .ZN(n20619) );
  INV_X1 U13086 ( .A(n15872), .ZN(n18829) );
  NAND2_X1 U13087 ( .A1(n10945), .A2(n13318), .ZN(n18834) );
  NAND2_X1 U13088 ( .A1(n19758), .A2(n13781), .ZN(n18946) );
  NAND2_X1 U13089 ( .A1(n18927), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18935) );
  NAND2_X1 U13090 ( .A1(n19758), .A2(n13780), .ZN(n18947) );
  INV_X1 U13091 ( .A(n15628), .ZN(n15015) );
  INV_X1 U13092 ( .A(n15677), .ZN(n15042) );
  INV_X1 U13093 ( .A(n15110), .ZN(n15122) );
  XNOR2_X1 U13094 ( .A(n13257), .B(n13258), .ZN(n19721) );
  NAND2_X1 U13095 ( .A1(n19014), .A2(n13204), .ZN(n15185) );
  NOR2_X1 U13096 ( .A1(n19017), .A2(n19016), .ZN(n18994) );
  NAND2_X1 U13097 ( .A1(n12685), .A2(n19014), .ZN(n15206) );
  NAND2_X1 U13098 ( .A1(n19023), .A2(n10537), .ZN(n13368) );
  INV_X1 U13099 ( .A(n19023), .ZN(n19056) );
  INV_X1 U13100 ( .A(n13788), .ZN(n13140) );
  INV_X1 U13101 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16261) );
  OR2_X1 U13102 ( .A1(n18834), .A2(n12687), .ZN(n19072) );
  INV_X1 U13103 ( .A(n19078), .ZN(n16272) );
  NAND2_X1 U13104 ( .A1(n13349), .A2(n9628), .ZN(n16306) );
  NAND2_X1 U13105 ( .A1(n13349), .A2(n10559), .ZN(n16308) );
  INV_X1 U13106 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19718) );
  INV_X1 U13107 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13226) );
  INV_X1 U13108 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19130) );
  NAND2_X1 U13109 ( .A1(n19143), .A2(n19228), .ZN(n19166) );
  INV_X1 U13110 ( .A(n19188), .ZN(n19196) );
  INV_X1 U13111 ( .A(n19221), .ZN(n19219) );
  OR2_X1 U13112 ( .A1(n19327), .A2(n19707), .ZN(n19254) );
  INV_X1 U13113 ( .A(n19281), .ZN(n19275) );
  OR2_X1 U13114 ( .A1(n19327), .A2(n19493), .ZN(n19315) );
  INV_X1 U13115 ( .A(n19344), .ZN(n19342) );
  OR2_X1 U13116 ( .A1(n19327), .A2(n19568), .ZN(n19379) );
  OR2_X1 U13117 ( .A1(n19519), .A2(n19380), .ZN(n19401) );
  INV_X1 U13118 ( .A(n19428), .ZN(n19437) );
  INV_X1 U13119 ( .A(n19433), .ZN(n19465) );
  AOI21_X1 U13120 ( .B1(n13849), .B2(n13848), .A(n13847), .ZN(n19484) );
  INV_X1 U13121 ( .A(n19515), .ZN(n19513) );
  OR2_X1 U13122 ( .A1(n19494), .A2(n19493), .ZN(n19545) );
  AOI22_X1 U13123 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19126), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19127), .ZN(n19583) );
  OR2_X1 U13124 ( .A1(n19519), .A2(n19568), .ZN(n19622) );
  NOR2_X1 U13125 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n15872) );
  INV_X1 U13126 ( .A(n19705), .ZN(n19632) );
  NAND2_X1 U13127 ( .A1(n19633), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19777) );
  INV_X1 U13128 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16515) );
  NOR2_X1 U13129 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16619), .ZN(n16612) );
  INV_X1 U13130 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17070) );
  NAND2_X1 U13131 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18666), .ZN(n16839) );
  INV_X1 U13132 ( .A(n16824), .ZN(n16865) );
  NOR3_X1 U13133 ( .A1(n16884), .A2(n16883), .A3(n16950), .ZN(n16945) );
  NOR2_X1 U13134 ( .A1(n20688), .A2(n17029), .ZN(n17017) );
  AND2_X1 U13135 ( .A1(n17195), .A2(n18204), .ZN(n17193) );
  INV_X2 U13136 ( .A(n17193), .ZN(n17188) );
  INV_X1 U13137 ( .A(n17327), .ZN(n17332) );
  NOR2_X1 U13138 ( .A1(n10120), .A2(n10119), .ZN(n17320) );
  NOR2_X1 U13139 ( .A1(n17391), .A2(n17331), .ZN(n17337) );
  NAND2_X1 U13140 ( .A1(n18161), .A2(n17368), .ZN(n17367) );
  INV_X1 U13141 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n20748) );
  INV_X1 U13142 ( .A(n17368), .ZN(n17396) );
  INV_X1 U13143 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17422) );
  INV_X1 U13144 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18190) );
  INV_X1 U13145 ( .A(n17455), .ZN(n20805) );
  INV_X1 U13146 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17453) );
  INV_X1 U13147 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17520) );
  INV_X1 U13148 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17867) );
  INV_X1 U13149 ( .A(n17601), .ZN(n17618) );
  AOI22_X1 U13150 ( .A1(n18013), .A2(n17803), .B1(n17724), .B2(n18015), .ZN(
        n17709) );
  INV_X1 U13151 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17775) );
  NAND2_X1 U13152 ( .A1(n16332), .A2(n18804), .ZN(n17815) );
  NAND2_X1 U13153 ( .A1(n16375), .A2(n18140), .ZN(n17947) );
  INV_X1 U13154 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18045) );
  INV_X1 U13155 ( .A(n18121), .ZN(n18128) );
  INV_X1 U13156 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18622) );
  INV_X1 U13157 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18644) );
  INV_X1 U13158 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16821) );
  INV_X1 U13159 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n20823) );
  INV_X1 U13160 ( .A(n18292), .ZN(n18282) );
  NAND2_X1 U13161 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18297), .ZN(
        n18343) );
  INV_X1 U13162 ( .A(n18380), .ZN(n18388) );
  INV_X1 U13163 ( .A(n18431), .ZN(n18425) );
  INV_X1 U13164 ( .A(n18475), .ZN(n18469) );
  INV_X1 U13165 ( .A(n18213), .ZN(n18555) );
  INV_X1 U13166 ( .A(n18223), .ZN(n18581) );
  NOR2_X1 U13167 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18667) );
  INV_X1 U13168 ( .A(n18750), .ZN(n18668) );
  NAND2_X1 U13169 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18814) );
  INV_X1 U13170 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18703) );
  NAND2_X1 U13171 ( .A1(n18677), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18818) );
  INV_X1 U13172 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18200) );
  INV_X1 U13173 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16480) );
  INV_X1 U13174 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19653) );
  NAND2_X1 U13175 ( .A1(n12134), .A2(n12133), .ZN(P1_U2873) );
  NAND2_X1 U13176 ( .A1(n10420), .A2(n10419), .ZN(P3_U2831) );
  INV_X1 U13177 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16359) );
  NAND2_X1 U13178 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17821) );
  INV_X1 U13179 ( .A(n17821), .ZN(n10403) );
  INV_X2 U13180 ( .A(n9674), .ZN(n17156) );
  AOI22_X1 U13181 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10097) );
  INV_X2 U13182 ( .A(n14284), .ZN(n14241) );
  NOR2_X2 U13183 ( .A1(n18612), .A2(n10104), .ZN(n10152) );
  AOI22_X1 U13184 ( .A1(n14241), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10096) );
  INV_X2 U13185 ( .A(n16952), .ZN(n17152) );
  NOR2_X2 U13186 ( .A1(n10102), .A2(n18633), .ZN(n10180) );
  AOI22_X1 U13187 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10095) );
  AOI22_X1 U13188 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10094) );
  NAND4_X1 U13189 ( .A1(n10097), .A2(n10096), .A3(n10095), .A4(n10094), .ZN(
        n10110) );
  NOR2_X2 U13190 ( .A1(n10104), .A2(n10101), .ZN(n17037) );
  AOI22_X1 U13191 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10108) );
  NOR2_X2 U13192 ( .A1(n18633), .A2(n10103), .ZN(n10100) );
  NOR2_X2 U13193 ( .A1(n10102), .A2(n10101), .ZN(n10153) );
  AOI22_X1 U13194 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17018), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10107) );
  BUF_X2 U13195 ( .A(n10279), .Z(n17079) );
  AOI22_X1 U13196 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17079), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10106) );
  NOR2_X2 U13197 ( .A1(n10104), .A2(n18635), .ZN(n10140) );
  AOI22_X1 U13198 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10105) );
  NAND4_X1 U13199 ( .A1(n10108), .A2(n10107), .A3(n10106), .A4(n10105), .ZN(
        n10109) );
  AOI22_X1 U13200 ( .A1(n14241), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10114) );
  AOI22_X1 U13201 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10113) );
  INV_X2 U13202 ( .A(n9593), .ZN(n17036) );
  AOI22_X1 U13203 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10112) );
  AOI22_X1 U13204 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10111) );
  NAND4_X1 U13205 ( .A1(n10114), .A2(n10113), .A3(n10112), .A4(n10111), .ZN(
        n10120) );
  AOI22_X1 U13206 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10118) );
  AOI22_X1 U13207 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10117) );
  AOI22_X1 U13208 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10116) );
  AOI22_X1 U13209 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10115) );
  NAND4_X1 U13210 ( .A1(n10118), .A2(n10117), .A3(n10116), .A4(n10115), .ZN(
        n10119) );
  AOI22_X1 U13211 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10124) );
  AOI22_X1 U13212 ( .A1(n10100), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10123) );
  AOI22_X1 U13213 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10122) );
  AOI22_X1 U13214 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10121) );
  NAND4_X1 U13215 ( .A1(n10124), .A2(n10123), .A3(n10122), .A4(n10121), .ZN(
        n10130) );
  AOI22_X1 U13216 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10128) );
  AOI22_X1 U13217 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10180), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10127) );
  INV_X2 U13218 ( .A(n14284), .ZN(n17150) );
  AOI22_X1 U13219 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10126) );
  AOI22_X1 U13220 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10140), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10125) );
  NAND4_X1 U13221 ( .A1(n10128), .A2(n10127), .A3(n10126), .A4(n10125), .ZN(
        n10129) );
  AOI22_X1 U13222 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17018), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10133) );
  AOI22_X1 U13223 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10132) );
  AOI22_X1 U13224 ( .A1(n10100), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10180), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10131) );
  AOI22_X1 U13225 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10136) );
  AOI22_X1 U13226 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10135) );
  NAND2_X1 U13227 ( .A1(n10154), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n10134) );
  AOI22_X1 U13228 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10140), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10138) );
  OAI21_X1 U13229 ( .B1(n9593), .B2(n18176), .A(n10138), .ZN(n10139) );
  AOI22_X1 U13230 ( .A1(n10100), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n10140), .ZN(n10145) );
  AOI22_X1 U13231 ( .A1(n10154), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n10093), .ZN(n10144) );
  AOI22_X1 U13232 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17018), .B1(
        n14241), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10143) );
  AOI22_X1 U13233 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n10141), .ZN(n10142) );
  NAND4_X1 U13234 ( .A1(n10145), .A2(n10144), .A3(n10143), .A4(n10142), .ZN(
        n10151) );
  AOI22_X1 U13235 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17153), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10149) );
  AOI22_X1 U13236 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n17151), .ZN(n10148) );
  AOI22_X1 U13237 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n9591), .B1(
        n10180), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10147) );
  AOI22_X1 U13238 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10146) );
  NAND4_X1 U13239 ( .A1(n10149), .A2(n10148), .A3(n10147), .A4(n10146), .ZN(
        n10150) );
  AOI22_X1 U13240 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10164) );
  AOI22_X1 U13241 ( .A1(n17018), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10163) );
  INV_X1 U13242 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18188) );
  AOI22_X1 U13243 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10155) );
  OAI21_X1 U13244 ( .B1(n9593), .B2(n18188), .A(n10155), .ZN(n10161) );
  AOI22_X1 U13245 ( .A1(n10100), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10180), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10159) );
  AOI22_X1 U13246 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10158) );
  AOI22_X1 U13247 ( .A1(n10280), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10140), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10157) );
  AOI22_X1 U13248 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10156) );
  NAND4_X1 U13249 ( .A1(n10159), .A2(n10158), .A3(n10157), .A4(n10156), .ZN(
        n10160) );
  AOI211_X1 U13250 ( .C1(n17157), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n10161), .B(n10160), .ZN(n10162) );
  NAND3_X1 U13251 ( .A1(n10164), .A2(n10163), .A3(n10162), .ZN(n17324) );
  NAND2_X1 U13252 ( .A1(n10178), .A2(n17324), .ZN(n10177) );
  AOI22_X1 U13253 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10175) );
  AOI22_X1 U13254 ( .A1(n14241), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U13255 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10165) );
  OAI21_X1 U13256 ( .B1(n10166), .B2(n20713), .A(n10165), .ZN(n10172) );
  AOI22_X1 U13257 ( .A1(n10280), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10170) );
  AOI22_X1 U13258 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10169) );
  AOI22_X1 U13259 ( .A1(n17018), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17079), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10168) );
  AOI22_X1 U13260 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10167) );
  NAND4_X1 U13261 ( .A1(n10170), .A2(n10169), .A3(n10168), .A4(n10167), .ZN(
        n10171) );
  AOI211_X1 U13262 ( .C1(n17166), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n10172), .B(n10171), .ZN(n10173) );
  NAND3_X1 U13263 ( .A1(n10175), .A2(n10174), .A3(n10173), .ZN(n17316) );
  INV_X1 U13264 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17845) );
  AOI21_X1 U13265 ( .B1(n17312), .B2(n10176), .A(n17722), .ZN(n10204) );
  XOR2_X1 U13266 ( .A(n17320), .B(n10177), .Z(n10197) );
  NAND2_X1 U13267 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n10195), .ZN(
        n10196) );
  INV_X1 U13268 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18110) );
  XOR2_X1 U13269 ( .A(n17328), .B(n10179), .Z(n17780) );
  XNOR2_X1 U13270 ( .A(n17334), .B(n17339), .ZN(n10193) );
  NAND2_X1 U13271 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10193), .ZN(
        n10194) );
  NAND2_X1 U13272 ( .A1(n10352), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10191) );
  AOI22_X1 U13273 ( .A1(n10154), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17018), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10184) );
  AOI22_X1 U13274 ( .A1(n10180), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10183) );
  AOI22_X1 U13275 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10182) );
  AOI22_X1 U13276 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10181) );
  NAND4_X1 U13277 ( .A1(n10184), .A2(n10183), .A3(n10182), .A4(n10181), .ZN(
        n10190) );
  AOI22_X1 U13278 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10188) );
  AOI22_X1 U13279 ( .A1(n10100), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10187) );
  AOI22_X1 U13280 ( .A1(n14241), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10186) );
  AOI22_X1 U13281 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10185) );
  NAND4_X1 U13282 ( .A1(n10188), .A2(n10187), .A3(n10186), .A4(n10185), .ZN(
        n10189) );
  NOR2_X1 U13283 ( .A1(n10190), .A2(n10189), .ZN(n17810) );
  NOR2_X1 U13284 ( .A1(n17810), .A2(n18781), .ZN(n17809) );
  NAND2_X1 U13285 ( .A1(n10191), .A2(n17800), .ZN(n17792) );
  INV_X1 U13286 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10192) );
  XNOR2_X1 U13287 ( .A(n10193), .B(n10192), .ZN(n17793) );
  NAND2_X1 U13288 ( .A1(n17792), .A2(n17793), .ZN(n17791) );
  XOR2_X1 U13289 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n10195), .Z(
        n17769) );
  NAND2_X1 U13290 ( .A1(n10197), .A2(n10199), .ZN(n10200) );
  INV_X1 U13291 ( .A(n10197), .ZN(n10198) );
  NAND2_X1 U13292 ( .A1(n10200), .A2(n17750), .ZN(n17739) );
  XOR2_X1 U13293 ( .A(n17316), .B(n10201), .Z(n10202) );
  XOR2_X1 U13294 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n10202), .Z(
        n17740) );
  NAND2_X1 U13295 ( .A1(n17739), .A2(n17740), .ZN(n17738) );
  NAND2_X1 U13296 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n10202), .ZN(
        n10203) );
  NAND2_X1 U13297 ( .A1(n10204), .A2(n10206), .ZN(n10207) );
  NAND2_X1 U13298 ( .A1(n17642), .A2(n17979), .ZN(n17620) );
  INV_X1 U13299 ( .A(n17620), .ZN(n10211) );
  INV_X1 U13300 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10209) );
  INV_X1 U13301 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10208) );
  AND2_X1 U13302 ( .A1(n10209), .A2(n10208), .ZN(n10210) );
  NAND2_X1 U13303 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17680) );
  NOR2_X1 U13304 ( .A1(n17680), .A2(n17679), .ZN(n18021) );
  NAND2_X1 U13305 ( .A1(n18021), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10213) );
  INV_X1 U13306 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17660) );
  NOR2_X1 U13307 ( .A1(n10213), .A2(n17660), .ZN(n17974) );
  NAND2_X1 U13308 ( .A1(n17974), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17640) );
  INV_X1 U13309 ( .A(n10213), .ZN(n17975) );
  INV_X2 U13310 ( .A(n17995), .ZN(n18015) );
  NAND2_X1 U13311 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17897) );
  INV_X1 U13312 ( .A(n17897), .ZN(n17932) );
  NAND2_X1 U13313 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17893) );
  INV_X1 U13314 ( .A(n17893), .ZN(n17874) );
  NAND3_X1 U13315 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n17874), .ZN(n17533) );
  INV_X1 U13316 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17886) );
  NOR2_X1 U13317 ( .A1(n17533), .A2(n17886), .ZN(n10405) );
  NAND2_X1 U13318 ( .A1(n17932), .A2(n10405), .ZN(n16342) );
  NOR2_X1 U13319 ( .A1(n17867), .A2(n16342), .ZN(n10402) );
  INV_X1 U13320 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17898) );
  NAND2_X1 U13321 ( .A1(n17898), .A2(n10223), .ZN(n17589) );
  NOR2_X1 U13322 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17589), .ZN(
        n10219) );
  NAND2_X1 U13323 ( .A1(n10219), .A2(n17878), .ZN(n17550) );
  NOR2_X1 U13324 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17550), .ZN(
        n17536) );
  NAND3_X1 U13325 ( .A1(n17536), .A2(n17867), .A3(n17886), .ZN(n10220) );
  OR2_X2 U13326 ( .A1(n17560), .A2(n17549), .ZN(n17590) );
  INV_X1 U13327 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17833) );
  NAND2_X1 U13328 ( .A1(n17722), .A2(n10224), .ZN(n17502) );
  OAI211_X2 U13329 ( .C1(n10403), .C2(n10223), .A(n17492), .B(n17502), .ZN(
        n10226) );
  NOR2_X2 U13330 ( .A1(n10226), .A2(n17818), .ZN(n17477) );
  AOI221_X1 U13331 ( .B1(n15851), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), 
        .C1(n10223), .C2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(n10227), .ZN(
        n10234) );
  INV_X1 U13332 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18762) );
  AOI22_X1 U13333 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n10223), .B1(
        n17722), .B2(n18762), .ZN(n10233) );
  NAND2_X1 U13334 ( .A1(n9795), .A2(n10228), .ZN(n10230) );
  NOR2_X1 U13335 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18762), .ZN(
        n10414) );
  OAI21_X1 U13336 ( .B1(n10230), .B2(n15851), .A(n10229), .ZN(n10231) );
  NAND2_X1 U13337 ( .A1(n10231), .A2(n10233), .ZN(n10232) );
  OAI21_X1 U13338 ( .B1(n10234), .B2(n10233), .A(n10232), .ZN(n16337) );
  AOI22_X1 U13339 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10238) );
  AOI22_X1 U13340 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10237) );
  AOI22_X1 U13341 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9591), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10236) );
  AOI22_X1 U13342 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10235) );
  NAND4_X1 U13343 ( .A1(n10238), .A2(n10237), .A3(n10236), .A4(n10235), .ZN(
        n10244) );
  INV_X2 U13344 ( .A(n10287), .ZN(n17081) );
  AOI22_X1 U13345 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10242) );
  INV_X2 U13346 ( .A(n16983), .ZN(n14285) );
  AOI22_X1 U13347 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10241) );
  AOI22_X1 U13348 ( .A1(n14241), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17079), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10240) );
  AOI22_X1 U13349 ( .A1(n17018), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10239) );
  NAND4_X1 U13350 ( .A1(n10242), .A2(n10241), .A3(n10240), .A4(n10239), .ZN(
        n10243) );
  AOI22_X1 U13351 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10254) );
  AOI22_X1 U13352 ( .A1(n14241), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10280), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10253) );
  AOI22_X1 U13353 ( .A1(n17079), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10245) );
  OAI21_X1 U13354 ( .B1(n16900), .B2(n18176), .A(n10245), .ZN(n10251) );
  AOI22_X1 U13355 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10249) );
  AOI22_X1 U13356 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10248) );
  AOI22_X1 U13357 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10247) );
  AOI22_X1 U13358 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10246) );
  NAND4_X1 U13359 ( .A1(n10249), .A2(n10248), .A3(n10247), .A4(n10246), .ZN(
        n10250) );
  AOI211_X1 U13360 ( .C1(n17123), .C2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n10251), .B(n10250), .ZN(n10252) );
  NOR2_X1 U13361 ( .A1(n18167), .A2(n18172), .ZN(n10343) );
  AOI22_X1 U13362 ( .A1(n17079), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10264) );
  AOI22_X1 U13363 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10263) );
  AOI22_X1 U13364 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10255) );
  OAI21_X1 U13365 ( .B1(n10287), .B2(n20713), .A(n10255), .ZN(n10261) );
  AOI22_X1 U13366 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10259) );
  AOI22_X1 U13367 ( .A1(n17018), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10180), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10258) );
  AOI22_X1 U13368 ( .A1(n10137), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10257) );
  AOI22_X1 U13369 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10280), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10256) );
  NAND4_X1 U13370 ( .A1(n10259), .A2(n10258), .A3(n10257), .A4(n10256), .ZN(
        n10260) );
  AOI211_X1 U13371 ( .C1(n17123), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n10261), .B(n10260), .ZN(n10262) );
  NAND3_X1 U13372 ( .A1(n10264), .A2(n10263), .A3(n10262), .ZN(n17201) );
  NAND2_X1 U13373 ( .A1(n10343), .A2(n17201), .ZN(n10326) );
  AOI22_X1 U13374 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10268) );
  AOI22_X1 U13375 ( .A1(n17018), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10267) );
  AOI22_X1 U13376 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10266) );
  AOI22_X1 U13377 ( .A1(n17079), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10265) );
  NAND4_X1 U13378 ( .A1(n10268), .A2(n10267), .A3(n10266), .A4(n10265), .ZN(
        n10274) );
  AOI22_X1 U13379 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10272) );
  AOI22_X1 U13380 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10271) );
  AOI22_X1 U13381 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10270) );
  AOI22_X1 U13382 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10269) );
  NAND4_X1 U13383 ( .A1(n10272), .A2(n10271), .A3(n10270), .A4(n10269), .ZN(
        n10273) );
  NOR2_X1 U13384 ( .A1(n10274), .A2(n10273), .ZN(n14207) );
  AOI22_X1 U13385 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10278) );
  AOI22_X1 U13386 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10180), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10277) );
  AOI22_X1 U13387 ( .A1(n14241), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10276) );
  AOI22_X1 U13388 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10275) );
  NAND4_X1 U13389 ( .A1(n10278), .A2(n10277), .A3(n10276), .A4(n10275), .ZN(
        n10286) );
  AOI22_X1 U13390 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10284) );
  AOI22_X1 U13391 ( .A1(n17018), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17079), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10283) );
  AOI22_X1 U13392 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10280), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10282) );
  AOI22_X1 U13393 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10281) );
  NAND4_X1 U13394 ( .A1(n10284), .A2(n10283), .A3(n10282), .A4(n10281), .ZN(
        n10285) );
  NAND2_X1 U13395 ( .A1(n10319), .A2(n18195), .ZN(n18617) );
  AOI22_X1 U13396 ( .A1(n17018), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10288) );
  OAI21_X1 U13397 ( .B1(n16900), .B2(n20823), .A(n10288), .ZN(n10294) );
  AOI22_X1 U13398 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10280), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10292) );
  AOI22_X1 U13399 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10291) );
  AOI22_X1 U13400 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10290) );
  AOI22_X1 U13401 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10289) );
  NAND4_X1 U13402 ( .A1(n10292), .A2(n10291), .A3(n10290), .A4(n10289), .ZN(
        n10293) );
  AOI22_X1 U13403 ( .A1(n14241), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10307) );
  AOI22_X1 U13404 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10306) );
  INV_X1 U13405 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18182) );
  AOI22_X1 U13406 ( .A1(n17079), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10298) );
  OAI21_X1 U13407 ( .B1(n16900), .B2(n18182), .A(n10298), .ZN(n10304) );
  AOI22_X1 U13408 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10302) );
  AOI22_X1 U13409 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10301) );
  AOI22_X1 U13410 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10300) );
  AOI22_X1 U13411 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10180), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10299) );
  NAND4_X1 U13412 ( .A1(n10302), .A2(n10301), .A3(n10300), .A4(n10299), .ZN(
        n10303) );
  AOI211_X1 U13413 ( .C1(n17123), .C2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A(
        n10304), .B(n10303), .ZN(n10305) );
  NAND3_X1 U13414 ( .A1(n10307), .A2(n10306), .A3(n10305), .ZN(n10390) );
  AOI22_X1 U13415 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U13416 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10316) );
  INV_X1 U13417 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18164) );
  AOI22_X1 U13418 ( .A1(n14241), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10308) );
  OAI21_X1 U13419 ( .B1(n16900), .B2(n18164), .A(n10308), .ZN(n10314) );
  AOI22_X1 U13420 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10312) );
  AOI22_X1 U13421 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10311) );
  AOI22_X1 U13422 ( .A1(n17079), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10137), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10310) );
  AOI22_X1 U13423 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10309) );
  NAND4_X1 U13424 ( .A1(n10312), .A2(n10311), .A3(n10310), .A4(n10309), .ZN(
        n10313) );
  AOI211_X1 U13425 ( .C1(n17123), .C2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n10314), .B(n10313), .ZN(n10315) );
  NAND2_X1 U13426 ( .A1(n10392), .A2(n18804), .ZN(n10393) );
  INV_X1 U13427 ( .A(n18172), .ZN(n10341) );
  NAND2_X1 U13428 ( .A1(n10393), .A2(n10341), .ZN(n10388) );
  NOR3_X1 U13429 ( .A1(n10391), .A2(n10381), .A3(n10388), .ZN(n10318) );
  OAI21_X1 U13430 ( .B1(n14207), .B2(n15879), .A(n10318), .ZN(n10325) );
  INV_X1 U13431 ( .A(n18600), .ZN(n18796) );
  INV_X1 U13432 ( .A(n14207), .ZN(n18185) );
  NAND2_X1 U13433 ( .A1(n18204), .A2(n10392), .ZN(n10320) );
  NAND2_X1 U13434 ( .A1(n17201), .A2(n10319), .ZN(n10389) );
  NAND2_X1 U13435 ( .A1(n18607), .A2(n18172), .ZN(n16485) );
  AND2_X1 U13436 ( .A1(n18204), .A2(n10389), .ZN(n10322) );
  NOR2_X1 U13437 ( .A1(n14207), .A2(n17201), .ZN(n18606) );
  NOR3_X1 U13438 ( .A1(n18606), .A2(n10391), .A3(n18172), .ZN(n10379) );
  AOI22_X1 U13439 ( .A1(n10392), .A2(n10379), .B1(n18179), .B2(n10320), .ZN(
        n10321) );
  OAI21_X1 U13440 ( .B1(n10322), .B2(n14207), .A(n10321), .ZN(n10323) );
  AOI21_X1 U13441 ( .B1(n14207), .B2(n15879), .A(n10323), .ZN(n10324) );
  INV_X1 U13442 ( .A(n10324), .ZN(n10387) );
  NAND2_X1 U13443 ( .A1(n18167), .A2(n18161), .ZN(n10395) );
  AOI21_X1 U13444 ( .B1(n18204), .B2(n18617), .A(n10395), .ZN(n10383) );
  AOI211_X1 U13445 ( .C1(n16485), .C2(n10325), .A(n10387), .B(n10383), .ZN(
        n15777) );
  INV_X1 U13446 ( .A(n10326), .ZN(n10350) );
  AOI22_X1 U13447 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18623), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18778), .ZN(n10347) );
  AND2_X1 U13448 ( .A1(n10347), .A2(n10333), .ZN(n10327) );
  AOI22_X1 U13449 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n18156), .B2(n18771), .ZN(
        n10328) );
  XNOR2_X1 U13450 ( .A(n10329), .B(n10328), .ZN(n10334) );
  INV_X1 U13451 ( .A(n10334), .ZN(n10340) );
  NOR2_X1 U13452 ( .A1(n10329), .A2(n10328), .ZN(n10330) );
  AOI22_X1 U13453 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16821), .B1(
        n10331), .B2(n20789), .ZN(n10336) );
  NOR2_X1 U13454 ( .A1(n10331), .A2(n20789), .ZN(n10337) );
  NAND2_X1 U13455 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16821), .ZN(
        n10332) );
  OAI22_X1 U13456 ( .A1(n10336), .A2(n18644), .B1(n10337), .B2(n10332), .ZN(
        n10335) );
  AOI211_X1 U13457 ( .C1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .C2(n18784), .A(
        n10333), .B(n10335), .ZN(n10346) );
  XOR2_X1 U13458 ( .A(n10347), .B(n10333), .Z(n10339) );
  OAI21_X1 U13459 ( .B1(n10337), .B2(n18644), .A(n10336), .ZN(n10338) );
  INV_X1 U13460 ( .A(n18601), .ZN(n16491) );
  AOI21_X1 U13461 ( .B1(n10340), .B2(n10346), .A(n16491), .ZN(n18797) );
  NOR2_X1 U13462 ( .A1(n18191), .A2(n18172), .ZN(n10380) );
  NAND2_X2 U13463 ( .A1(n18817), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18743) );
  OAI21_X1 U13464 ( .B1(n10341), .B2(n18804), .A(n18674), .ZN(n10342) );
  OAI21_X1 U13465 ( .B1(n10343), .B2(n10342), .A(n18814), .ZN(n16490) );
  NOR3_X1 U13466 ( .A1(n10380), .A2(n16491), .A3(n16490), .ZN(n10349) );
  INV_X1 U13467 ( .A(n18795), .ZN(n14205) );
  AOI211_X1 U13468 ( .C1(n14207), .C2(n10389), .A(n18172), .B(n14205), .ZN(
        n10348) );
  AOI211_X1 U13469 ( .C1(n10350), .C2(n18797), .A(n10349), .B(n10348), .ZN(
        n10351) );
  NAND2_X1 U13470 ( .A1(n16337), .A2(n18057), .ZN(n10420) );
  INV_X1 U13471 ( .A(n17640), .ZN(n17959) );
  NOR2_X1 U13472 ( .A1(n17810), .A2(n10352), .ZN(n10360) );
  NOR2_X1 U13473 ( .A1(n10360), .A2(n10353), .ZN(n10358) );
  NOR2_X1 U13474 ( .A1(n10358), .A2(n17328), .ZN(n10357) );
  NAND2_X1 U13475 ( .A1(n10357), .A2(n17324), .ZN(n10356) );
  NOR2_X1 U13476 ( .A1(n17320), .A2(n10356), .ZN(n10355) );
  NAND2_X1 U13477 ( .A1(n10355), .A2(n17316), .ZN(n10354) );
  NOR2_X1 U13478 ( .A1(n17312), .A2(n10354), .ZN(n10376) );
  XNOR2_X1 U13479 ( .A(n10354), .B(n16375), .ZN(n10372) );
  XOR2_X1 U13480 ( .A(n10355), .B(n17316), .Z(n10368) );
  XOR2_X1 U13481 ( .A(n10356), .B(n17320), .Z(n17754) );
  INV_X1 U13482 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18097) );
  XOR2_X1 U13483 ( .A(n10357), .B(n17324), .Z(n17764) );
  XOR2_X1 U13484 ( .A(n17328), .B(n10358), .Z(n10359) );
  NAND2_X1 U13485 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n10359), .ZN(
        n10365) );
  XOR2_X1 U13486 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n10359), .Z(
        n17778) );
  XOR2_X1 U13487 ( .A(n17334), .B(n10360), .Z(n10361) );
  NAND2_X1 U13488 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10361), .ZN(
        n10364) );
  XOR2_X1 U13489 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n10361), .Z(
        n17790) );
  INV_X1 U13490 ( .A(n17810), .ZN(n15880) );
  AOI21_X1 U13491 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17339), .A(
        n15880), .ZN(n10363) );
  NOR2_X1 U13492 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17339), .ZN(
        n10362) );
  AOI221_X1 U13493 ( .B1(n15880), .B2(n17339), .C1(n10363), .C2(n18781), .A(
        n10362), .ZN(n17789) );
  NAND2_X1 U13494 ( .A1(n17790), .A2(n17789), .ZN(n17788) );
  NAND2_X1 U13495 ( .A1(n10364), .A2(n17788), .ZN(n17777) );
  NAND2_X1 U13496 ( .A1(n17778), .A2(n17777), .ZN(n17776) );
  NAND2_X1 U13497 ( .A1(n10365), .A2(n17776), .ZN(n17765) );
  NAND2_X1 U13498 ( .A1(n17764), .A2(n17765), .ZN(n17763) );
  NOR2_X1 U13499 ( .A1(n17764), .A2(n17765), .ZN(n10366) );
  AOI21_X1 U13500 ( .B1(n18097), .B2(n17763), .A(n10366), .ZN(n17753) );
  NOR2_X1 U13501 ( .A1(n17754), .A2(n17753), .ZN(n10367) );
  INV_X1 U13502 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18085) );
  NAND2_X1 U13503 ( .A1(n17754), .A2(n17753), .ZN(n17752) );
  OAI21_X1 U13504 ( .B1(n10367), .B2(n18085), .A(n17752), .ZN(n10369) );
  NAND2_X1 U13505 ( .A1(n10368), .A2(n10369), .ZN(n10370) );
  XOR2_X1 U13506 ( .A(n10369), .B(n10368), .Z(n17742) );
  NAND2_X1 U13507 ( .A1(n17742), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17741) );
  NAND2_X1 U13508 ( .A1(n10370), .A2(n17741), .ZN(n10373) );
  NOR2_X1 U13509 ( .A1(n10372), .A2(n10373), .ZN(n17732) );
  NOR2_X1 U13510 ( .A1(n17732), .A2(n20725), .ZN(n10371) );
  NAND2_X1 U13511 ( .A1(n10376), .A2(n10371), .ZN(n10377) );
  INV_X1 U13512 ( .A(n10371), .ZN(n10375) );
  AND2_X1 U13513 ( .A1(n10373), .A2(n10372), .ZN(n17733) );
  AOI21_X1 U13514 ( .B1(n10376), .B2(n10375), .A(n17733), .ZN(n10374) );
  OAI21_X1 U13515 ( .B1(n10376), .B2(n10375), .A(n10374), .ZN(n17711) );
  NAND2_X1 U13516 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17711), .ZN(
        n17710) );
  NAND2_X1 U13517 ( .A1(n17959), .A2(n18013), .ZN(n17633) );
  NOR2_X2 U13518 ( .A1(n17633), .A2(n10208), .ZN(n17883) );
  NAND2_X1 U13519 ( .A1(n17883), .A2(n10402), .ZN(n17859) );
  NOR2_X1 U13520 ( .A1(n17859), .A2(n17520), .ZN(n17501) );
  NAND2_X1 U13521 ( .A1(n17501), .A2(n10403), .ZN(n15786) );
  INV_X1 U13522 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17463) );
  NOR2_X1 U13523 ( .A1(n17818), .A2(n17463), .ZN(n15787) );
  NAND2_X1 U13524 ( .A1(n15787), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16354) );
  NOR2_X1 U13525 ( .A1(n15786), .A2(n16354), .ZN(n16362) );
  NAND2_X1 U13526 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16362), .ZN(
        n10378) );
  XNOR2_X1 U13527 ( .A(n18762), .B(n10378), .ZN(n16340) );
  NAND2_X1 U13528 ( .A1(n10395), .A2(n10393), .ZN(n18822) );
  NOR2_X1 U13529 ( .A1(n10380), .A2(n10379), .ZN(n10384) );
  NAND2_X1 U13530 ( .A1(n18606), .A2(n10382), .ZN(n14204) );
  NAND2_X1 U13531 ( .A1(n18804), .A2(n18161), .ZN(n14208) );
  OAI21_X1 U13532 ( .B1(n10384), .B2(n10383), .A(n10390), .ZN(n10385) );
  INV_X1 U13533 ( .A(n10385), .ZN(n10386) );
  AND2_X1 U13534 ( .A1(n18607), .A2(n10398), .ZN(n18632) );
  NOR2_X1 U13535 ( .A1(n18172), .A2(n10390), .ZN(n18605) );
  NAND2_X1 U13536 ( .A1(n10391), .A2(n18605), .ZN(n14203) );
  NAND2_X1 U13537 ( .A1(n18167), .A2(n10392), .ZN(n15876) );
  OR2_X1 U13538 ( .A1(n10392), .A2(n10394), .ZN(n16486) );
  NAND3_X2 U13539 ( .A1(n10397), .A2(n16486), .A3(n10396), .ZN(n18631) );
  NAND2_X1 U13540 ( .A1(n18632), .A2(n10401), .ZN(n15783) );
  NOR2_X2 U13541 ( .A1(n15776), .A2(n15775), .ZN(n18602) );
  NAND2_X2 U13542 ( .A1(n18602), .A2(n10397), .ZN(n18621) );
  INV_X2 U13543 ( .A(n18621), .ZN(n18130) );
  INV_X2 U13544 ( .A(n18028), .ZN(n18022) );
  NAND2_X1 U13545 ( .A1(n18804), .A2(n10401), .ZN(n10399) );
  OAI21_X1 U13546 ( .B1(n10400), .B2(n10399), .A(n10398), .ZN(n18604) );
  AOI21_X2 U13547 ( .B1(n18605), .B2(n10401), .A(n18604), .ZN(n18618) );
  NAND2_X2 U13548 ( .A1(n18022), .A2(n18618), .ZN(n18051) );
  NOR2_X4 U13549 ( .A1(n18804), .A2(n18051), .ZN(n17875) );
  NAND2_X1 U13550 ( .A1(n18015), .A2(n17929), .ZN(n17884) );
  NAND2_X1 U13551 ( .A1(n10402), .A2(n17962), .ZN(n17858) );
  NOR2_X1 U13552 ( .A1(n17520), .A2(n17858), .ZN(n17500) );
  NAND2_X1 U13553 ( .A1(n10403), .A2(n17500), .ZN(n17826) );
  NOR2_X1 U13554 ( .A1(n16354), .A2(n17826), .ZN(n16358) );
  NAND2_X1 U13555 ( .A1(n16358), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10404) );
  XOR2_X1 U13556 ( .A(n10404), .B(n18762), .Z(n16333) );
  NAND2_X1 U13557 ( .A1(n17312), .A2(n18140), .ZN(n17996) );
  INV_X1 U13558 ( .A(n17996), .ZN(n18058) );
  NAND2_X1 U13559 ( .A1(n18051), .A2(n18127), .ZN(n18129) );
  INV_X1 U13560 ( .A(n18129), .ZN(n15793) );
  INV_X1 U13561 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18740) );
  INV_X1 U13562 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18763) );
  NAND2_X1 U13563 ( .A1(n18763), .A2(n18752), .ZN(n18766) );
  OR3_X2 U13564 ( .A1(n18766), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18094) );
  NOR2_X1 U13565 ( .A1(n18740), .A2(n18094), .ZN(n16331) );
  NAND2_X1 U13566 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17841) );
  NOR2_X1 U13567 ( .A1(n17821), .A2(n17841), .ZN(n16344) );
  INV_X1 U13568 ( .A(n16344), .ZN(n17817) );
  AOI21_X1 U13569 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18048) );
  NAND3_X1 U13570 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18072) );
  INV_X1 U13571 ( .A(n18072), .ZN(n18063) );
  NAND4_X1 U13572 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A4(n18063), .ZN(n17961) );
  NOR2_X1 U13573 ( .A1(n18048), .A2(n17961), .ZN(n17949) );
  NAND2_X1 U13574 ( .A1(n17929), .A2(n17949), .ZN(n17876) );
  NOR2_X1 U13575 ( .A1(n17897), .A2(n17876), .ZN(n17931) );
  NAND2_X1 U13576 ( .A1(n10405), .A2(n17931), .ZN(n17862) );
  OAI21_X1 U13577 ( .B1(n17817), .B2(n17862), .A(n18639), .ZN(n17822) );
  INV_X1 U13578 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18054) );
  NAND2_X1 U13579 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18091) );
  NOR2_X1 U13580 ( .A1(n18072), .A2(n18091), .ZN(n18050) );
  NAND3_X1 U13581 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n18050), .ZN(n18039) );
  OR2_X1 U13582 ( .A1(n18054), .A2(n18039), .ZN(n17950) );
  NOR2_X1 U13583 ( .A1(n16341), .A2(n17950), .ZN(n17930) );
  NOR2_X1 U13584 ( .A1(n17897), .A2(n17533), .ZN(n17880) );
  NAND2_X1 U13585 ( .A1(n17930), .A2(n17880), .ZN(n17820) );
  OR2_X1 U13586 ( .A1(n17886), .A2(n17820), .ZN(n10406) );
  OAI21_X1 U13587 ( .B1(n17817), .B2(n10406), .A(n18621), .ZN(n10409) );
  NOR2_X1 U13588 ( .A1(n18781), .A2(n10406), .ZN(n17819) );
  INV_X1 U13589 ( .A(n17819), .ZN(n10407) );
  NAND2_X1 U13590 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n16344), .ZN(
        n16372) );
  INV_X1 U13591 ( .A(n18618), .ZN(n18611) );
  OAI21_X1 U13592 ( .B1(n10407), .B2(n16372), .A(n18611), .ZN(n10408) );
  NAND4_X1 U13593 ( .A1(n18128), .A2(n17822), .A3(n10409), .A4(n10408), .ZN(
        n15790) );
  AOI22_X1 U13594 ( .A1(n15793), .A2(n16354), .B1(n18094), .B2(n15790), .ZN(
        n15856) );
  INV_X1 U13595 ( .A(n17876), .ZN(n10411) );
  AOI21_X1 U13596 ( .B1(n18611), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18621), .ZN(n18114) );
  INV_X1 U13597 ( .A(n18114), .ZN(n10410) );
  AOI22_X1 U13598 ( .A1(n18639), .A2(n10411), .B1(n10410), .B2(n17930), .ZN(
        n16371) );
  NOR2_X1 U13599 ( .A1(n16371), .A2(n16342), .ZN(n17842) );
  NAND4_X1 U13600 ( .A1(n15787), .A2(n18127), .A3(n17842), .A4(n16344), .ZN(
        n15788) );
  NAND3_X1 U13601 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n18762), .ZN(n10412) );
  OAI22_X1 U13602 ( .A1(n15856), .A2(n18762), .B1(n15788), .B2(n10412), .ZN(
        n10413) );
  AOI211_X1 U13603 ( .C1(n10414), .C2(n15793), .A(n16331), .B(n10413), .ZN(
        n10415) );
  INV_X1 U13604 ( .A(n10418), .ZN(n10419) );
  AND2_X4 U13605 ( .A1(n10674), .A2(n10596), .ZN(n10664) );
  AOI22_X1 U13606 ( .A1(n9630), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10424) );
  AOI22_X1 U13607 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10423) );
  AND2_X4 U13608 ( .A1(n10670), .A2(n10596), .ZN(n10665) );
  AND2_X4 U13609 ( .A1(n10672), .A2(n13699), .ZN(n10675) );
  AND2_X4 U13610 ( .A1(n10672), .A2(n10596), .ZN(n10515) );
  AOI22_X1 U13611 ( .A1(n10675), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10421) );
  NAND4_X1 U13612 ( .A1(n10424), .A2(n10423), .A3(n10422), .A4(n10421), .ZN(
        n10425) );
  AOI22_X1 U13613 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9587), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10429) );
  AOI22_X1 U13614 ( .A1(n9629), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10428) );
  AOI22_X1 U13615 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10427) );
  AOI22_X1 U13616 ( .A1(n10675), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10426) );
  NAND4_X1 U13617 ( .A1(n10429), .A2(n10428), .A3(n10427), .A4(n10426), .ZN(
        n10431) );
  AOI22_X1 U13618 ( .A1(n10675), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9641), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10437) );
  AOI22_X1 U13619 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10436) );
  AOI22_X1 U13620 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10434) );
  NAND4_X1 U13621 ( .A1(n10437), .A2(n10436), .A3(n10435), .A4(n10434), .ZN(
        n10438) );
  AOI22_X1 U13622 ( .A1(n10675), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9641), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10442) );
  AOI22_X1 U13623 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9587), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10440) );
  AOI22_X1 U13624 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10439) );
  NAND4_X1 U13625 ( .A1(n10439), .A2(n10441), .A3(n10440), .A4(n10442), .ZN(
        n10443) );
  AOI22_X1 U13626 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10449) );
  AOI22_X1 U13627 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10448) );
  NAND4_X1 U13628 ( .A1(n10450), .A2(n10449), .A3(n10448), .A4(n10447), .ZN(
        n10458) );
  AOI22_X1 U13629 ( .A1(n9629), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__4__SCAN_IN), .B2(n10515), .ZN(n10452) );
  AOI22_X1 U13630 ( .A1(n10675), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9641), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10451) );
  AOI22_X1 U13631 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10454) );
  AOI22_X1 U13632 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9587), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10453) );
  AOI22_X1 U13633 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9587), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10462) );
  AOI22_X1 U13634 ( .A1(n9630), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10461) );
  AOI22_X1 U13635 ( .A1(n10675), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9641), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10460) );
  AOI22_X1 U13636 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10459) );
  NAND4_X1 U13637 ( .A1(n10462), .A2(n10461), .A3(n10460), .A4(n10459), .ZN(
        n10463) );
  AOI22_X1 U13638 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9641), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10466) );
  AOI22_X1 U13639 ( .A1(n10515), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10465) );
  AOI22_X1 U13640 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10464) );
  NAND4_X1 U13641 ( .A1(n10467), .A2(n10466), .A3(n10465), .A4(n10464), .ZN(
        n10468) );
  NAND2_X1 U13642 ( .A1(n10468), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10469) );
  NAND2_X2 U13643 ( .A1(n10469), .A2(n10470), .ZN(n10523) );
  XNOR2_X1 U13644 ( .A(n10550), .B(n10523), .ZN(n13205) );
  OAI21_X1 U13645 ( .B1(n10528), .B2(n10550), .A(n10548), .ZN(n10471) );
  OAI211_X1 U13646 ( .C1(n13205), .C2(n10548), .A(n10471), .B(n9622), .ZN(
        n13331) );
  AOI22_X1 U13647 ( .A1(n10675), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10473) );
  AOI22_X1 U13648 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9638), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U13649 ( .A1(n9629), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10475) );
  AOI22_X1 U13650 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10474) );
  AOI22_X1 U13651 ( .A1(n9629), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10479) );
  AOI22_X1 U13652 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10477) );
  AOI22_X1 U13653 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10476) );
  AOI22_X1 U13654 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13655 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U13656 ( .A1(n10675), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10484) );
  AOI22_X1 U13657 ( .A1(n9630), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10483) );
  NAND2_X1 U13658 ( .A1(n10487), .A2(n10430), .ZN(n10496) );
  NAND2_X1 U13659 ( .A1(n10488), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10489) );
  AOI22_X1 U13660 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10493) );
  AOI22_X1 U13661 ( .A1(n9630), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U13662 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10491) );
  NAND2_X2 U13663 ( .A1(n10496), .A2(n10495), .ZN(n10551) );
  AOI22_X1 U13664 ( .A1(n10675), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10500) );
  AOI22_X1 U13665 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9587), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U13666 ( .A1(n9630), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10498) );
  AOI22_X1 U13667 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10497) );
  NAND4_X1 U13668 ( .A1(n10500), .A2(n10499), .A3(n10498), .A4(n10497), .ZN(
        n10506) );
  AOI22_X1 U13669 ( .A1(n10675), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10504) );
  AOI22_X1 U13670 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10503) );
  AOI22_X1 U13671 ( .A1(n9629), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10502) );
  AOI22_X1 U13672 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10501) );
  NAND4_X1 U13673 ( .A1(n10504), .A2(n10503), .A3(n10502), .A4(n10501), .ZN(
        n10505) );
  MUX2_X2 U13674 ( .A(n10506), .B(n10505), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10538) );
  INV_X1 U13675 ( .A(n10538), .ZN(n12680) );
  NAND3_X1 U13676 ( .A1(n10564), .A2(n12680), .A3(n9615), .ZN(n10572) );
  NAND2_X1 U13677 ( .A1(n10572), .A2(n19765), .ZN(n10527) );
  NAND2_X1 U13678 ( .A1(n10548), .A2(n9622), .ZN(n10507) );
  OAI21_X1 U13679 ( .B1(n10548), .B2(n10508), .A(n10507), .ZN(n10521) );
  AOI22_X1 U13680 ( .A1(n10675), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9641), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10509) );
  AOI22_X1 U13681 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10512) );
  AOI22_X1 U13682 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9587), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10511) );
  AOI22_X1 U13683 ( .A1(n10675), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9641), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10514) );
  AOI22_X1 U13684 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10513) );
  AOI22_X1 U13685 ( .A1(n9629), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10515), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10517) );
  AOI22_X1 U13686 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n9587), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10516) );
  NAND3_X1 U13687 ( .A1(n10522), .A2(n10521), .A3(n19103), .ZN(n10526) );
  NAND2_X1 U13688 ( .A1(n10549), .A2(n10523), .ZN(n10524) );
  NAND2_X1 U13689 ( .A1(n10550), .A2(n10533), .ZN(n10540) );
  NAND2_X1 U13690 ( .A1(n19103), .A2(n10549), .ZN(n10584) );
  NAND2_X1 U13691 ( .A1(n10525), .A2(n13334), .ZN(n10541) );
  NAND3_X1 U13692 ( .A1(n10526), .A2(n10541), .A3(n19765), .ZN(n13338) );
  NAND2_X1 U13693 ( .A1(n10532), .A2(n10929), .ZN(n10536) );
  NAND2_X1 U13694 ( .A1(n10528), .A2(n9622), .ZN(n12671) );
  NAND2_X1 U13695 ( .A1(n10536), .A2(n13208), .ZN(n13195) );
  NAND2_X1 U13696 ( .A1(n10595), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10545) );
  INV_X1 U13697 ( .A(n10584), .ZN(n13330) );
  INV_X1 U13698 ( .A(n10540), .ZN(n12661) );
  NAND3_X1 U13699 ( .A1(n12660), .A2(n10528), .A3(n12661), .ZN(n10542) );
  INV_X1 U13700 ( .A(n10561), .ZN(n10543) );
  OR2_X2 U13701 ( .A1(n13208), .A2(n19765), .ZN(n13078) );
  NAND2_X2 U13702 ( .A1(n10543), .A2(n13078), .ZN(n13320) );
  NAND2_X1 U13703 ( .A1(n10545), .A2(n10544), .ZN(n10590) );
  NAND3_X1 U13704 ( .A1(n12658), .A2(n10548), .A3(n9622), .ZN(n10558) );
  NAND3_X1 U13705 ( .A1(n10508), .A2(n10528), .A3(n10551), .ZN(n10552) );
  NAND2_X1 U13706 ( .A1(n19109), .A2(n10552), .ZN(n10556) );
  NOR2_X2 U13707 ( .A1(n10558), .A2(n10557), .ZN(n12655) );
  INV_X1 U13708 ( .A(n19761), .ZN(n10559) );
  NAND2_X1 U13709 ( .A1(n10559), .A2(n13306), .ZN(n13748) );
  NAND2_X1 U13710 ( .A1(n10587), .A2(n13748), .ZN(n10560) );
  NAND2_X1 U13711 ( .A1(n10560), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10563) );
  INV_X1 U13713 ( .A(n10564), .ZN(n12659) );
  AND2_X2 U13714 ( .A1(n12659), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10600) );
  NAND2_X1 U13715 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10566) );
  OAI21_X1 U13716 ( .B1(n10585), .B2(n14115), .A(n10566), .ZN(n10567) );
  INV_X1 U13717 ( .A(n10567), .ZN(n10568) );
  NAND2_X1 U13718 ( .A1(n10568), .A2(n10569), .ZN(n10570) );
  XNOR2_X2 U13719 ( .A(n10590), .B(n10591), .ZN(n10621) );
  AOI21_X1 U13720 ( .B1(n10571), .B2(n10572), .A(n10573), .ZN(n10582) );
  NAND2_X1 U13721 ( .A1(n9624), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10581) );
  INV_X1 U13722 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n10574) );
  INV_X1 U13723 ( .A(n13749), .ZN(n10576) );
  NAND2_X1 U13724 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10575) );
  AND2_X1 U13725 ( .A1(n10576), .A2(n10575), .ZN(n10579) );
  NAND2_X1 U13726 ( .A1(n10610), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10577) );
  OAI211_X2 U13727 ( .C1(n10582), .C2(n19762), .A(n10581), .B(n10580), .ZN(
        n10615) );
  INV_X1 U13728 ( .A(n9617), .ZN(n13321) );
  NAND2_X1 U13729 ( .A1(n10589), .A2(n10588), .ZN(n10614) );
  INV_X1 U13730 ( .A(n10590), .ZN(n10592) );
  NAND2_X1 U13731 ( .A1(n10592), .A2(n10591), .ZN(n10593) );
  NAND2_X1 U13732 ( .A1(n10595), .A2(n10596), .ZN(n10598) );
  AOI21_X1 U13733 ( .B1(n19762), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10597) );
  NAND2_X1 U13734 ( .A1(n10598), .A2(n10597), .ZN(n10604) );
  NAND2_X1 U13735 ( .A1(n10610), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10602) );
  NAND2_X1 U13736 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10601) );
  OAI211_X1 U13737 ( .C1(n13977), .C2(n9671), .A(n10602), .B(n10601), .ZN(
        n10603) );
  INV_X1 U13738 ( .A(n10604), .ZN(n10606) );
  NAND2_X1 U13739 ( .A1(n10606), .A2(n10605), .ZN(n10607) );
  NAND2_X1 U13740 ( .A1(n10595), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10609) );
  NAND2_X1 U13741 ( .A1(n13749), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10608) );
  NAND2_X1 U13742 ( .A1(n10609), .A2(n10608), .ZN(n11116) );
  INV_X1 U13743 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10949) );
  NAND2_X1 U13744 ( .A1(n10610), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10612) );
  NAND2_X1 U13745 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10611) );
  OAI211_X1 U13746 ( .C1(n10949), .C2(n9671), .A(n10612), .B(n10611), .ZN(
        n10613) );
  XNOR2_X2 U13747 ( .A(n11113), .B(n11117), .ZN(n12157) );
  INV_X1 U13748 ( .A(n10614), .ZN(n10617) );
  AND2_X1 U13749 ( .A1(n12157), .A2(n9815), .ZN(n10657) );
  BUF_X4 U13750 ( .A(n12146), .Z(n10647) );
  NAND2_X1 U13751 ( .A1(n19526), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10632) );
  NOR2_X4 U13752 ( .A1(n10658), .A2(n12141), .ZN(n19229) );
  NAND2_X1 U13753 ( .A1(n19229), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10631) );
  NAND2_X1 U13754 ( .A1(n10807), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10630) );
  INV_X1 U13755 ( .A(n19089), .ZN(n10833) );
  INV_X1 U13756 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12486) );
  NOR2_X1 U13757 ( .A1(n10833), .A2(n12486), .ZN(n10628) );
  INV_X1 U13758 ( .A(n10621), .ZN(n10623) );
  NAND2_X1 U13759 ( .A1(n19079), .A2(n10623), .ZN(n10645) );
  BUF_X4 U13760 ( .A(n12157), .Z(n13412) );
  INV_X1 U13761 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12189) );
  INV_X1 U13762 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10625) );
  OAI211_X1 U13763 ( .C1(n19136), .C2(n12189), .A(n10626), .B(n10753), .ZN(
        n10627) );
  NOR2_X1 U13764 ( .A1(n10628), .A2(n10627), .ZN(n10629) );
  NAND4_X1 U13765 ( .A1(n10632), .A2(n10631), .A3(n10630), .A4(n10629), .ZN(
        n10722) );
  INV_X1 U13766 ( .A(n10654), .ZN(n10633) );
  INV_X1 U13767 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12198) );
  AND2_X1 U13768 ( .A1(n10621), .A2(n19079), .ZN(n10639) );
  NAND2_X1 U13769 ( .A1(n10647), .A2(n10639), .ZN(n10635) );
  OR2_X2 U13770 ( .A1(n13412), .A2(n10635), .ZN(n19319) );
  INV_X1 U13771 ( .A(n10635), .ZN(n10636) );
  INV_X1 U13772 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12197) );
  OAI22_X1 U13773 ( .A1(n12198), .A2(n19319), .B1(n19571), .B2(n12197), .ZN(
        n10637) );
  NOR2_X1 U13774 ( .A1(n10638), .A2(n10637), .ZN(n10662) );
  INV_X1 U13775 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10644) );
  INV_X1 U13776 ( .A(n10639), .ZN(n10640) );
  OR2_X1 U13777 ( .A1(n10647), .A2(n10640), .ZN(n10642) );
  INV_X1 U13778 ( .A(n10642), .ZN(n10641) );
  NAND2_X2 U13779 ( .A1(n10641), .A2(n13412), .ZN(n19442) );
  OR2_X2 U13780 ( .A1(n10642), .A2(n13412), .ZN(n10792) );
  INV_X1 U13781 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10643) );
  OAI22_X1 U13782 ( .A1(n10644), .A2(n19442), .B1(n10792), .B2(n10643), .ZN(
        n10653) );
  INV_X1 U13783 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10651) );
  INV_X1 U13784 ( .A(n10645), .ZN(n10646) );
  NAND2_X1 U13785 ( .A1(n10647), .A2(n10646), .ZN(n10648) );
  INV_X1 U13786 ( .A(n10648), .ZN(n10649) );
  INV_X1 U13787 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10650) );
  OAI22_X1 U13788 ( .A1(n10651), .A2(n10800), .B1(n19487), .B2(n10650), .ZN(
        n10652) );
  INV_X1 U13789 ( .A(n10655), .ZN(n10656) );
  AND2_X2 U13790 ( .A1(n10657), .A2(n10656), .ZN(n19356) );
  NAND2_X1 U13791 ( .A1(n19290), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10659) );
  NAND4_X1 U13792 ( .A1(n10661), .A2(n10662), .A3(n10660), .A4(n10659), .ZN(
        n10721) );
  AND2_X2 U13793 ( .A1(n12623), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12377) );
  NAND3_X1 U13794 ( .A1(n10596), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10936) );
  AOI22_X1 U13795 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n12340), .ZN(n10669) );
  INV_X1 U13796 ( .A(n10515), .ZN(n12598) );
  AOI22_X1 U13797 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12392), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10668) );
  AND2_X2 U13798 ( .A1(n12587), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10777) );
  AOI22_X1 U13799 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10777), .B1(
        n13712), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10667) );
  AOI22_X1 U13800 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12464), .B1(
        n10714), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10666) );
  NAND4_X1 U13801 ( .A1(n10669), .A2(n10668), .A3(n10667), .A4(n10666), .ZN(
        n10684) );
  AND2_X2 U13802 ( .A1(n10670), .A2(n12429), .ZN(n12451) );
  AOI22_X1 U13803 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12452), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10682) );
  AND2_X1 U13804 ( .A1(n12429), .A2(n10674), .ZN(n10704) );
  AOI22_X1 U13805 ( .A1(n10673), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10681) );
  AND2_X2 U13806 ( .A1(n12625), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10676) );
  AOI22_X1 U13807 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12380), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10680) );
  INV_X1 U13808 ( .A(n10936), .ZN(n10678) );
  AOI22_X1 U13809 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n12453), .ZN(n10679) );
  NAND4_X1 U13810 ( .A1(n10682), .A2(n10681), .A3(n10680), .A4(n10679), .ZN(
        n10683) );
  NOR2_X1 U13811 ( .A1(n10684), .A2(n10683), .ZN(n12693) );
  INV_X1 U13812 ( .A(n10538), .ZN(n12687) );
  AOI22_X1 U13813 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10688) );
  NAND2_X1 U13814 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10687) );
  NAND2_X1 U13815 ( .A1(n12464), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10686) );
  NAND2_X1 U13816 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10685) );
  AOI22_X1 U13817 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13712), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10689) );
  INV_X1 U13818 ( .A(n10689), .ZN(n10693) );
  INV_X1 U13819 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n19265) );
  AOI22_X1 U13820 ( .A1(n12380), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10691) );
  AOI22_X1 U13821 ( .A1(n10714), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10777), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10690) );
  NOR2_X1 U13822 ( .A1(n10693), .A2(n10692), .ZN(n10699) );
  NAND2_X1 U13823 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10697) );
  NAND2_X1 U13824 ( .A1(n10673), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10696) );
  INV_X1 U13825 ( .A(n9669), .ZN(n12340) );
  AOI22_X1 U13826 ( .A1(n12453), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10695) );
  NAND2_X1 U13827 ( .A1(n12452), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10694) );
  AND4_X1 U13828 ( .A1(n10697), .A2(n10696), .A3(n10695), .A4(n10694), .ZN(
        n10698) );
  NAND3_X1 U13829 ( .A1(n10078), .A2(n10699), .A3(n10698), .ZN(n12679) );
  NAND2_X1 U13830 ( .A1(n12687), .A2(n12679), .ZN(n13383) );
  OR2_X1 U13831 ( .A1(n12693), .A2(n13383), .ZN(n10761) );
  NAND2_X1 U13832 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n10703) );
  NAND2_X1 U13833 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10702) );
  NAND2_X1 U13834 ( .A1(n10777), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10701) );
  NAND2_X1 U13835 ( .A1(n13712), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10700) );
  NAND4_X1 U13836 ( .A1(n10703), .A2(n10702), .A3(n10701), .A4(n10700), .ZN(
        n10713) );
  AOI22_X1 U13837 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n12451), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10711) );
  NAND2_X1 U13838 ( .A1(n12380), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10710) );
  NAND2_X1 U13839 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10709) );
  INV_X1 U13840 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10706) );
  NAND2_X1 U13841 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n12340), .ZN(
        n10705) );
  OAI21_X1 U13842 ( .B1(n12343), .B2(n10706), .A(n10705), .ZN(n10707) );
  AOI21_X1 U13843 ( .B1(n12452), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n10707), .ZN(n10708) );
  NAND4_X1 U13844 ( .A1(n10711), .A2(n10710), .A3(n10709), .A4(n10708), .ZN(
        n10712) );
  NOR2_X1 U13845 ( .A1(n10713), .A2(n10712), .ZN(n10719) );
  AOI22_X1 U13846 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__2__SCAN_IN), .B2(n10673), .ZN(n10718) );
  NAND2_X1 U13847 ( .A1(n12464), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10717) );
  NAND2_X1 U13848 ( .A1(n10714), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10716) );
  NAND2_X1 U13849 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10715) );
  NAND2_X1 U13850 ( .A1(n10761), .A2(n12703), .ZN(n10720) );
  NAND2_X1 U13851 ( .A1(n19526), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10725) );
  NAND2_X1 U13852 ( .A1(n10807), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10724) );
  NAND2_X1 U13853 ( .A1(n10725), .A2(n10724), .ZN(n10726) );
  NOR2_X1 U13854 ( .A1(n10082), .A2(n10726), .ZN(n10742) );
  INV_X1 U13855 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10728) );
  INV_X1 U13856 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12240) );
  OAI22_X1 U13857 ( .A1(n10728), .A2(n10727), .B1(n19319), .B2(n12240), .ZN(
        n10731) );
  INV_X1 U13858 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10729) );
  INV_X1 U13859 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12239) );
  OAI22_X1 U13860 ( .A1(n10729), .A2(n10792), .B1(n19571), .B2(n12239), .ZN(
        n10730) );
  NOR2_X1 U13861 ( .A1(n10731), .A2(n10730), .ZN(n10741) );
  INV_X1 U13862 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10733) );
  INV_X1 U13863 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10732) );
  OAI22_X1 U13864 ( .A1(n10733), .A2(n19442), .B1(n10800), .B2(n10732), .ZN(
        n10735) );
  INV_X1 U13865 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12229) );
  INV_X1 U13866 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12533) );
  OAI22_X1 U13867 ( .A1(n12229), .A2(n19136), .B1(n19487), .B2(n12533), .ZN(
        n10734) );
  NAND2_X1 U13868 ( .A1(n19229), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10738) );
  AOI22_X1 U13869 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19169), .B1(
        n19356), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10737) );
  AOI22_X1 U13870 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19089), .B1(
        n19409), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10736) );
  NAND3_X1 U13871 ( .A1(n10742), .A2(n10740), .A3(n10741), .ZN(n10755) );
  AOI22_X1 U13872 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12460), .B1(
        n12377), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10746) );
  AOI22_X1 U13873 ( .A1(n12380), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__3__SCAN_IN), .B2(n10704), .ZN(n10745) );
  AOI22_X1 U13874 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__3__SCAN_IN), .B2(n12340), .ZN(n10744) );
  AOI22_X1 U13875 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10673), .B1(
        n12452), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10743) );
  NAND4_X1 U13876 ( .A1(n10746), .A2(n10745), .A3(n10744), .A4(n10743), .ZN(
        n10752) );
  AOI22_X1 U13877 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12464), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10750) );
  AOI22_X1 U13878 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n12453), .ZN(n10749) );
  AOI22_X1 U13879 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13712), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10748) );
  AOI22_X1 U13880 ( .A1(n10714), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10777), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10747) );
  NAND4_X1 U13881 ( .A1(n10750), .A2(n10749), .A3(n10748), .A4(n10747), .ZN(
        n10751) );
  INV_X1 U13882 ( .A(n12715), .ZN(n10948) );
  NAND2_X1 U13883 ( .A1(n10948), .A2(n12687), .ZN(n10754) );
  AND2_X2 U13884 ( .A1(n10755), .A2(n10754), .ZN(n10767) );
  XNOR2_X2 U13885 ( .A(n10723), .B(n10767), .ZN(n13864) );
  INV_X1 U13886 ( .A(n13383), .ZN(n10756) );
  INV_X1 U13887 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13345) );
  NOR2_X1 U13888 ( .A1(n10756), .A2(n13345), .ZN(n13381) );
  INV_X1 U13889 ( .A(n12693), .ZN(n10758) );
  INV_X1 U13890 ( .A(n12679), .ZN(n10757) );
  XNOR2_X1 U13891 ( .A(n10758), .B(n10757), .ZN(n10759) );
  NAND2_X1 U13892 ( .A1(n13381), .A2(n10759), .ZN(n10760) );
  XOR2_X1 U13893 ( .A(n13381), .B(n10759), .Z(n13143) );
  NAND2_X1 U13894 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13143), .ZN(
        n13142) );
  NAND2_X1 U13895 ( .A1(n10760), .A2(n13142), .ZN(n10762) );
  XOR2_X1 U13896 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n10762), .Z(
        n13152) );
  XNOR2_X1 U13897 ( .A(n12703), .B(n10761), .ZN(n13151) );
  NAND2_X1 U13898 ( .A1(n13152), .A2(n13151), .ZN(n13150) );
  NAND2_X1 U13899 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10762), .ZN(
        n10763) );
  NAND2_X1 U13900 ( .A1(n13150), .A2(n10763), .ZN(n10764) );
  INV_X1 U13901 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13877) );
  XNOR2_X1 U13902 ( .A(n10764), .B(n13877), .ZN(n13865) );
  NAND2_X1 U13903 ( .A1(n13864), .A2(n13865), .ZN(n10766) );
  NAND2_X1 U13904 ( .A1(n10764), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10765) );
  AOI22_X1 U13905 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12460), .B1(
        n12377), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10776) );
  AOI22_X1 U13906 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12464), .B1(
        n10714), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10775) );
  AOI22_X1 U13907 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12379), .B1(
        n12380), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10774) );
  NAND2_X1 U13908 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10772) );
  NAND2_X1 U13909 ( .A1(n12452), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10771) );
  NAND2_X1 U13910 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10770) );
  AOI22_X1 U13911 ( .A1(n12453), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__4__SCAN_IN), .B2(n12340), .ZN(n10769) );
  AND4_X1 U13912 ( .A1(n10772), .A2(n10771), .A3(n10770), .A4(n10769), .ZN(
        n10773) );
  NAND4_X1 U13913 ( .A1(n10776), .A2(n10775), .A3(n10774), .A4(n10773), .ZN(
        n10782) );
  AOI22_X1 U13914 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n13712), .B1(
        n10777), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10780) );
  AOI22_X1 U13915 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__4__SCAN_IN), .B2(n10673), .ZN(n10779) );
  NAND2_X1 U13916 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10778) );
  NAND3_X1 U13917 ( .A1(n10780), .A2(n10779), .A3(n10778), .ZN(n10781) );
  INV_X1 U13918 ( .A(n12721), .ZN(n10783) );
  XNOR2_X1 U13919 ( .A(n10788), .B(n10783), .ZN(n10785) );
  INV_X1 U13920 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n16300) );
  INV_X1 U13921 ( .A(n10784), .ZN(n10786) );
  NAND2_X1 U13922 ( .A1(n10786), .A2(n10785), .ZN(n10787) );
  INV_X1 U13923 ( .A(n10788), .ZN(n10789) );
  NAND2_X2 U13924 ( .A1(n10789), .A2(n12721), .ZN(n10877) );
  AOI22_X1 U13925 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19169), .B1(
        n19409), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10806) );
  INV_X1 U13926 ( .A(n19356), .ZN(n10790) );
  INV_X1 U13927 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12397) );
  OAI22_X1 U13928 ( .A1(n10833), .A2(n13370), .B1(n10790), .B2(n12397), .ZN(
        n10791) );
  INV_X1 U13929 ( .A(n10791), .ZN(n10805) );
  INV_X1 U13930 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10794) );
  INV_X1 U13931 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10793) );
  OAI22_X1 U13932 ( .A1(n10794), .A2(n19136), .B1(n10792), .B2(n10793), .ZN(
        n10797) );
  INV_X1 U13933 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10795) );
  INV_X1 U13934 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12395) );
  OAI22_X1 U13935 ( .A1(n10795), .A2(n10727), .B1(n19571), .B2(n12395), .ZN(
        n10796) );
  NOR2_X1 U13936 ( .A1(n10797), .A2(n10796), .ZN(n10804) );
  INV_X1 U13937 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10799) );
  INV_X1 U13938 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10798) );
  OAI22_X1 U13939 ( .A1(n10799), .A2(n19442), .B1(n19319), .B2(n10798), .ZN(
        n10802) );
  INV_X1 U13940 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12393) );
  INV_X1 U13941 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12579) );
  OAI22_X1 U13942 ( .A1(n12393), .A2(n10800), .B1(n19487), .B2(n12579), .ZN(
        n10801) );
  NOR2_X1 U13943 ( .A1(n10802), .A2(n10801), .ZN(n10803) );
  NAND4_X1 U13944 ( .A1(n10806), .A2(n10805), .A3(n10804), .A4(n10803), .ZN(
        n10813) );
  NAND2_X1 U13945 ( .A1(n19229), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10811) );
  NAND2_X1 U13946 ( .A1(n19290), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10810) );
  NAND2_X1 U13947 ( .A1(n19526), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10809) );
  NAND2_X1 U13948 ( .A1(n10807), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10808) );
  NAND4_X1 U13949 ( .A1(n10811), .A2(n10810), .A3(n10809), .A4(n10808), .ZN(
        n10812) );
  NAND2_X1 U13950 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10817) );
  NAND2_X1 U13951 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10816) );
  NAND2_X1 U13952 ( .A1(n10777), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10815) );
  NAND2_X1 U13953 ( .A1(n13712), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10814) );
  NAND4_X1 U13954 ( .A1(n10817), .A2(n10816), .A3(n10815), .A4(n10814), .ZN(
        n10825) );
  AOI22_X1 U13955 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10823) );
  NAND2_X1 U13956 ( .A1(n12380), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10822) );
  NAND2_X1 U13957 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10821) );
  NAND2_X1 U13958 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n12340), .ZN(
        n10818) );
  OAI21_X1 U13959 ( .B1(n12343), .B2(n13370), .A(n10818), .ZN(n10819) );
  AOI21_X1 U13960 ( .B1(n12452), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n10819), .ZN(n10820) );
  NAND4_X1 U13961 ( .A1(n10823), .A2(n10822), .A3(n10821), .A4(n10820), .ZN(
        n10824) );
  NOR2_X1 U13962 ( .A1(n10825), .A2(n10824), .ZN(n10830) );
  AOI22_X1 U13963 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10829) );
  NAND2_X1 U13964 ( .A1(n12464), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10828) );
  NAND2_X1 U13965 ( .A1(n10714), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10827) );
  NAND2_X1 U13966 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10826) );
  NAND2_X1 U13967 ( .A1(n12687), .A2(n12725), .ZN(n10831) );
  INV_X1 U13968 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16303) );
  INV_X1 U13969 ( .A(n10877), .ZN(n10875) );
  AOI22_X1 U13970 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19169), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10846) );
  INV_X1 U13971 ( .A(n19409), .ZN(n19414) );
  INV_X1 U13972 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12421) );
  OAI22_X1 U13973 ( .A1(n19130), .A2(n10833), .B1(n19414), .B2(n12421), .ZN(
        n10834) );
  INV_X1 U13974 ( .A(n10834), .ZN(n10845) );
  INV_X1 U13975 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10836) );
  INV_X1 U13976 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10835) );
  OAI22_X1 U13977 ( .A1(n10836), .A2(n19319), .B1(n10800), .B2(n10835), .ZN(
        n10838) );
  INV_X1 U13978 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12592) );
  INV_X1 U13979 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12411) );
  OAI22_X1 U13980 ( .A1(n12592), .A2(n19442), .B1(n19487), .B2(n12411), .ZN(
        n10837) );
  NOR2_X1 U13981 ( .A1(n10838), .A2(n10837), .ZN(n10844) );
  INV_X1 U13982 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12595) );
  INV_X1 U13983 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10839) );
  OAI22_X1 U13984 ( .A1(n12595), .A2(n19136), .B1(n10792), .B2(n10839), .ZN(
        n10842) );
  INV_X1 U13985 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12417) );
  INV_X1 U13986 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10840) );
  OAI22_X1 U13987 ( .A1(n12417), .A2(n10727), .B1(n19571), .B2(n10840), .ZN(
        n10841) );
  NOR2_X1 U13988 ( .A1(n10842), .A2(n10841), .ZN(n10843) );
  NAND4_X1 U13989 ( .A1(n10846), .A2(n10845), .A3(n10844), .A4(n10843), .ZN(
        n10852) );
  NAND2_X1 U13990 ( .A1(n19229), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10850) );
  NAND2_X1 U13991 ( .A1(n19290), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10849) );
  NAND2_X1 U13992 ( .A1(n19526), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10848) );
  NAND2_X1 U13993 ( .A1(n10807), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10847) );
  NAND4_X1 U13994 ( .A1(n10850), .A2(n10849), .A3(n10848), .A4(n10847), .ZN(
        n10851) );
  NAND2_X1 U13995 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n10856) );
  NAND2_X1 U13996 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n10855) );
  NAND2_X1 U13997 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10854) );
  NAND2_X1 U13998 ( .A1(n10777), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10853) );
  AND4_X1 U13999 ( .A1(n10856), .A2(n10855), .A3(n10854), .A4(n10853), .ZN(
        n10869) );
  AOI22_X1 U14000 ( .A1(n12464), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13712), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10868) );
  NAND2_X1 U14001 ( .A1(n10714), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10859) );
  NAND2_X1 U14002 ( .A1(n10673), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n10858) );
  NAND2_X1 U14003 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n10857) );
  AND3_X1 U14004 ( .A1(n10859), .A2(n10858), .A3(n10857), .ZN(n10867) );
  AOI22_X1 U14005 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10865) );
  NAND2_X1 U14006 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10864) );
  NAND2_X1 U14007 ( .A1(n12380), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10863) );
  NAND2_X1 U14008 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n12340), .ZN(
        n10860) );
  OAI21_X1 U14009 ( .B1(n19130), .B2(n12343), .A(n10860), .ZN(n10861) );
  AOI21_X1 U14010 ( .B1(n12452), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n10861), .ZN(n10862) );
  AND4_X1 U14011 ( .A1(n10865), .A2(n10864), .A3(n10863), .A4(n10862), .ZN(
        n10866) );
  NAND4_X1 U14012 ( .A1(n10869), .A2(n10868), .A3(n10867), .A4(n10866), .ZN(
        n12729) );
  INV_X1 U14013 ( .A(n12729), .ZN(n10870) );
  NAND2_X1 U14014 ( .A1(n10870), .A2(n12687), .ZN(n10871) );
  OAI21_X1 U14015 ( .B1(n10877), .B2(n10876), .A(n10879), .ZN(n10878) );
  AND2_X2 U14016 ( .A1(n10906), .A2(n10878), .ZN(n10998) );
  NAND2_X1 U14017 ( .A1(n10972), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10883) );
  INV_X1 U14018 ( .A(n10883), .ZN(n14033) );
  NAND2_X1 U14019 ( .A1(n14033), .A2(n10879), .ZN(n10880) );
  NAND2_X1 U14020 ( .A1(n14094), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14095) );
  NAND2_X1 U14021 ( .A1(n10882), .A2(n10883), .ZN(n10884) );
  NAND2_X1 U14022 ( .A1(n10884), .A2(n10998), .ZN(n10885) );
  NAND2_X1 U14023 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10889) );
  NAND2_X1 U14024 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10888) );
  NAND2_X1 U14025 ( .A1(n10777), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10887) );
  NAND2_X1 U14026 ( .A1(n13712), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10886) );
  NAND2_X1 U14027 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10892) );
  NAND2_X1 U14028 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10891) );
  NAND2_X1 U14029 ( .A1(n10673), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10890) );
  AOI22_X1 U14030 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n12451), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10898) );
  NAND2_X1 U14031 ( .A1(n12380), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10897) );
  NAND2_X1 U14032 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10896) );
  NAND2_X1 U14033 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n12340), .ZN(
        n10893) );
  OAI21_X1 U14034 ( .B1(n12343), .B2(n12617), .A(n10893), .ZN(n10894) );
  AOI21_X1 U14035 ( .B1(n12452), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n10894), .ZN(n10895) );
  NAND2_X1 U14036 ( .A1(n12464), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10901) );
  NAND2_X1 U14037 ( .A1(n10714), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10900) );
  XNOR2_X1 U14038 ( .A(n10906), .B(n15240), .ZN(n14158) );
  INV_X1 U14039 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15753) );
  OAI21_X1 U14040 ( .B1(n10906), .B2(n15240), .A(n15753), .ZN(n10908) );
  INV_X1 U14041 ( .A(n10906), .ZN(n10907) );
  NAND2_X1 U14042 ( .A1(n10907), .A2(n11006), .ZN(n10911) );
  NAND2_X1 U14043 ( .A1(n10908), .A2(n10911), .ZN(n15440) );
  NAND2_X1 U14044 ( .A1(n10910), .A2(n10909), .ZN(n15439) );
  NAND2_X1 U14045 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15646) );
  INV_X1 U14046 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15652) );
  NOR2_X1 U14047 ( .A1(n15646), .A2(n15652), .ZN(n10912) );
  NAND2_X1 U14048 ( .A1(n15656), .A2(n10912), .ZN(n15636) );
  NAND2_X1 U14049 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15458) );
  INV_X1 U14050 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15517) );
  OAI21_X1 U14051 ( .B1(n15250), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15230), .ZN(n15507) );
  MUX2_X1 U14052 ( .A(n19735), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n10938) );
  INV_X1 U14053 ( .A(n10937), .ZN(n10915) );
  NAND2_X1 U14054 ( .A1(n10938), .A2(n10915), .ZN(n10917) );
  NAND2_X1 U14055 ( .A1(n19735), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10916) );
  NAND2_X1 U14056 ( .A1(n10917), .A2(n10916), .ZN(n10921) );
  MUX2_X1 U14057 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n19725), .S(
        n10596), .Z(n10919) );
  XNOR2_X1 U14058 ( .A(n10921), .B(n10919), .ZN(n12638) );
  INV_X1 U14059 ( .A(n12703), .ZN(n10918) );
  MUX2_X1 U14060 ( .A(n12638), .B(n10918), .S(n9628), .Z(n10946) );
  INV_X1 U14061 ( .A(n10938), .ZN(n12642) );
  OAI21_X1 U14062 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20827), .A(
        n10937), .ZN(n12643) );
  NOR2_X1 U14063 ( .A1(n12642), .A2(n12643), .ZN(n10928) );
  INV_X1 U14064 ( .A(n10919), .ZN(n10920) );
  NAND2_X1 U14065 ( .A1(n10921), .A2(n10920), .ZN(n10923) );
  NAND2_X1 U14066 ( .A1(n19725), .A2(n10596), .ZN(n10922) );
  NAND2_X1 U14067 ( .A1(n10923), .A2(n10922), .ZN(n10927) );
  XNOR2_X1 U14068 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10925) );
  NOR2_X1 U14069 ( .A1(n10430), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10924) );
  NOR2_X1 U14070 ( .A1(n15875), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10930) );
  NAND2_X1 U14071 ( .A1(n10931), .A2(n10930), .ZN(n10956) );
  INV_X1 U14072 ( .A(n10925), .ZN(n10926) );
  XNOR2_X1 U14073 ( .A(n10927), .B(n10926), .ZN(n10952) );
  OAI21_X1 U14074 ( .B1(n10946), .B2(n10928), .A(n12648), .ZN(n19748) );
  NAND2_X1 U14075 ( .A1(n15875), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10932) );
  NAND2_X1 U14076 ( .A1(n10559), .A2(n19747), .ZN(n10934) );
  NOR2_X1 U14077 ( .A1(n10929), .A2(n10934), .ZN(n10935) );
  NAND2_X1 U14078 ( .A1(n19748), .A2(n10935), .ZN(n13311) );
  NAND2_X1 U14079 ( .A1(n13226), .A2(n10936), .ZN(n13223) );
  INV_X1 U14080 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n18835) );
  OAI211_X1 U14081 ( .C1(n10714), .C2(n13223), .A(P2_STATE2_REG_1__SCAN_IN), 
        .B(n18835), .ZN(n19741) );
  NAND2_X1 U14082 ( .A1(n12648), .A2(n12638), .ZN(n10941) );
  XNOR2_X1 U14083 ( .A(n10938), .B(n10937), .ZN(n12636) );
  INV_X1 U14084 ( .A(n10941), .ZN(n10939) );
  NAND2_X1 U14085 ( .A1(n12636), .A2(n10939), .ZN(n10940) );
  OAI21_X1 U14086 ( .B1(n12643), .B2(n10941), .A(n13687), .ZN(n10942) );
  NAND2_X1 U14087 ( .A1(n19726), .A2(n10942), .ZN(n10943) );
  INV_X1 U14088 ( .A(n16319), .ZN(n19750) );
  NOR2_X1 U14089 ( .A1(n10929), .A2(n19750), .ZN(n13305) );
  NAND2_X1 U14090 ( .A1(n13305), .A2(n9628), .ZN(n10944) );
  NAND2_X1 U14091 ( .A1(n13311), .A2(n10944), .ZN(n10945) );
  NAND2_X1 U14092 ( .A1(n19726), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19631) );
  NOR2_X1 U14093 ( .A1(n15507), .A2(n19075), .ZN(n11224) );
  MUX2_X1 U14094 ( .A(n10946), .B(n13977), .S(n15217), .Z(n10982) );
  NAND2_X1 U14095 ( .A1(n14115), .A2(n10574), .ZN(n10947) );
  MUX2_X1 U14096 ( .A(n12693), .B(n10947), .S(n15217), .Z(n10985) );
  NAND2_X1 U14097 ( .A1(n10546), .A2(n12678), .ZN(n10955) );
  NAND2_X1 U14098 ( .A1(n9628), .A2(n10948), .ZN(n10950) );
  MUX2_X1 U14099 ( .A(n10950), .B(n10949), .S(n15217), .Z(n10951) );
  OAI21_X1 U14100 ( .B1(n10952), .B2(n10955), .A(n10951), .ZN(n10977) );
  NOR2_X1 U14101 ( .A1(n10985), .A2(n10977), .ZN(n10953) );
  NAND2_X1 U14102 ( .A1(n9628), .A2(n12721), .ZN(n10954) );
  MUX2_X1 U14103 ( .A(n10954), .B(P2_EBX_REG_4__SCAN_IN), .S(n15217), .Z(
        n10959) );
  INV_X1 U14104 ( .A(n10955), .ZN(n10957) );
  NAND2_X1 U14105 ( .A1(n10957), .A2(n10956), .ZN(n10958) );
  NAND2_X1 U14106 ( .A1(n10959), .A2(n10958), .ZN(n10992) );
  MUX2_X1 U14107 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n12725), .S(n12678), .Z(
        n10973) );
  INV_X1 U14108 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13967) );
  MUX2_X1 U14109 ( .A(n13967), .B(n12729), .S(n12678), .Z(n10999) );
  INV_X1 U14110 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13391) );
  MUX2_X1 U14111 ( .A(n13391), .B(n15220), .S(n12678), .Z(n11007) );
  NAND2_X1 U14112 ( .A1(n15217), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11004) );
  INV_X1 U14113 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n13528) );
  INV_X1 U14114 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n10960) );
  NAND2_X1 U14115 ( .A1(n11023), .A2(n10960), .ZN(n11032) );
  NAND2_X1 U14116 ( .A1(n11094), .A2(n11032), .ZN(n11024) );
  NAND2_X1 U14117 ( .A1(n15217), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11034) );
  NAND2_X1 U14118 ( .A1(n15217), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11068) );
  INV_X1 U14119 ( .A(n11068), .ZN(n10961) );
  INV_X1 U14120 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n10962) );
  NAND2_X1 U14121 ( .A1(n18896), .A2(n10962), .ZN(n10963) );
  NAND2_X1 U14122 ( .A1(n15217), .A2(n10963), .ZN(n10964) );
  OAI21_X1 U14123 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(P2_EBX_REG_16__SCAN_IN), 
        .A(n15217), .ZN(n10965) );
  INV_X1 U14124 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n11166) );
  NOR2_X1 U14125 ( .A1(n12678), .A2(n11166), .ZN(n11045) );
  NAND2_X1 U14126 ( .A1(n10528), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11043) );
  NAND2_X1 U14127 ( .A1(n11038), .A2(n15112), .ZN(n11086) );
  INV_X1 U14128 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15799) );
  NOR2_X1 U14129 ( .A1(n12678), .A2(n15799), .ZN(n11085) );
  NAND2_X1 U14130 ( .A1(n10528), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11089) );
  INV_X1 U14131 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n15090) );
  NAND2_X1 U14132 ( .A1(n11094), .A2(n10966), .ZN(n11099) );
  NAND2_X1 U14133 ( .A1(n15217), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14947) );
  NAND2_X1 U14134 ( .A1(n11099), .A2(n14947), .ZN(n14949) );
  INV_X1 U14135 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n11200) );
  NOR2_X1 U14136 ( .A1(n12678), .A2(n11200), .ZN(n11109) );
  INV_X1 U14137 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n11205) );
  NOR2_X1 U14138 ( .A1(n12678), .A2(n11205), .ZN(n10967) );
  NAND2_X1 U14139 ( .A1(n10968), .A2(n10967), .ZN(n10969) );
  NAND2_X1 U14140 ( .A1(n15216), .A2(n10969), .ZN(n14935) );
  OR2_X1 U14141 ( .A1(n14935), .A2(n15240), .ZN(n10970) );
  INV_X1 U14142 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15496) );
  NAND2_X1 U14143 ( .A1(n10970), .A2(n15496), .ZN(n15211) );
  NAND2_X1 U14144 ( .A1(n15220), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10971) );
  NAND2_X1 U14145 ( .A1(n15211), .A2(n15213), .ZN(n11112) );
  NAND2_X1 U14146 ( .A1(n10972), .A2(n15240), .ZN(n10976) );
  AND2_X1 U14147 ( .A1(n10974), .A2(n10973), .ZN(n10975) );
  OR2_X1 U14148 ( .A1(n10975), .A2(n11000), .ZN(n18937) );
  XNOR2_X1 U14149 ( .A(n10996), .B(n16303), .ZN(n14028) );
  INV_X1 U14150 ( .A(n10993), .ZN(n10980) );
  INV_X1 U14151 ( .A(n10982), .ZN(n10978) );
  OAI21_X1 U14152 ( .B1(n10978), .B2(n10985), .A(n10977), .ZN(n10979) );
  NAND2_X1 U14153 ( .A1(n10980), .A2(n10979), .ZN(n13808) );
  NAND2_X1 U14154 ( .A1(n10981), .A2(n13808), .ZN(n10989) );
  NAND2_X1 U14155 ( .A1(n10989), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13866) );
  XNOR2_X1 U14156 ( .A(n10982), .B(n10985), .ZN(n13980) );
  INV_X1 U14157 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13823) );
  XNOR2_X1 U14158 ( .A(n13980), .B(n13823), .ZN(n13156) );
  AND2_X1 U14159 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n10983) );
  NAND2_X1 U14160 ( .A1(n15217), .A2(n10983), .ZN(n10984) );
  NAND2_X1 U14161 ( .A1(n10985), .A2(n10984), .ZN(n14121) );
  INV_X1 U14162 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14067) );
  MUX2_X1 U14163 ( .A(P2_EBX_REG_0__SCAN_IN), .B(n12679), .S(n12678), .Z(
        n14076) );
  NAND2_X1 U14164 ( .A1(n14076), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13384) );
  OAI21_X1 U14165 ( .B1(n14121), .B2(n14067), .A(n13384), .ZN(n10987) );
  NAND2_X1 U14166 ( .A1(n14121), .A2(n14067), .ZN(n10986) );
  AND2_X1 U14167 ( .A1(n10987), .A2(n10986), .ZN(n13155) );
  NAND2_X1 U14168 ( .A1(n13156), .A2(n13155), .ZN(n13443) );
  NAND2_X1 U14169 ( .A1(n13980), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10988) );
  AND2_X1 U14170 ( .A1(n13443), .A2(n10988), .ZN(n13869) );
  NAND2_X1 U14171 ( .A1(n13866), .A2(n13869), .ZN(n10991) );
  INV_X1 U14172 ( .A(n10989), .ZN(n10990) );
  NAND2_X1 U14173 ( .A1(n10990), .A2(n13877), .ZN(n13867) );
  NAND2_X1 U14174 ( .A1(n10991), .A2(n13867), .ZN(n13818) );
  XNOR2_X1 U14175 ( .A(n10993), .B(n10992), .ZN(n13891) );
  XNOR2_X1 U14176 ( .A(n13891), .B(n16300), .ZN(n13817) );
  INV_X1 U14177 ( .A(n13891), .ZN(n10994) );
  NAND2_X1 U14178 ( .A1(n10994), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10995) );
  NAND2_X1 U14179 ( .A1(n10996), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10997) );
  NAND2_X1 U14180 ( .A1(n10998), .A2(n15240), .ZN(n11002) );
  NOR2_X1 U14181 ( .A1(n11000), .A2(n10999), .ZN(n11001) );
  OR2_X1 U14182 ( .A1(n11009), .A2(n11001), .ZN(n13968) );
  INV_X1 U14183 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14166) );
  XNOR2_X1 U14184 ( .A(n11005), .B(n11004), .ZN(n13914) );
  NAND2_X1 U14185 ( .A1(n13914), .A2(n11006), .ZN(n15435) );
  INV_X1 U14186 ( .A(n11007), .ZN(n11008) );
  XNOR2_X1 U14187 ( .A(n11009), .B(n11008), .ZN(n13793) );
  NAND2_X1 U14188 ( .A1(n13793), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15433) );
  NAND2_X1 U14189 ( .A1(n13914), .A2(n15220), .ZN(n11010) );
  NAND2_X1 U14190 ( .A1(n11010), .A2(n15753), .ZN(n15436) );
  INV_X1 U14191 ( .A(n13793), .ZN(n11011) );
  NAND2_X1 U14192 ( .A1(n11011), .A2(n9951), .ZN(n15432) );
  AND2_X1 U14193 ( .A1(n15436), .A2(n15432), .ZN(n11012) );
  NAND2_X1 U14194 ( .A1(n15217), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11014) );
  XNOR2_X1 U14195 ( .A(n11015), .B(n11014), .ZN(n18924) );
  NAND2_X1 U14196 ( .A1(n18924), .A2(n15220), .ZN(n11030) );
  INV_X1 U14197 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11029) );
  AND2_X1 U14198 ( .A1(n11030), .A2(n11029), .ZN(n16267) );
  INV_X1 U14199 ( .A(n16267), .ZN(n11016) );
  NAND2_X1 U14200 ( .A1(n10528), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11018) );
  OAI21_X1 U14201 ( .B1(n11019), .B2(n11018), .A(n11094), .ZN(n11020) );
  OR2_X1 U14202 ( .A1(n11023), .A2(n11020), .ZN(n13987) );
  INV_X1 U14203 ( .A(n13987), .ZN(n11021) );
  NAND2_X1 U14204 ( .A1(n11021), .A2(n15220), .ZN(n11031) );
  AND2_X1 U14205 ( .A1(n11031), .A2(n16275), .ZN(n15736) );
  NAND2_X1 U14206 ( .A1(n10528), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11022) );
  OR2_X1 U14207 ( .A1(n11023), .A2(n11022), .ZN(n11026) );
  INV_X1 U14208 ( .A(n11024), .ZN(n11025) );
  NAND2_X1 U14209 ( .A1(n13943), .A2(n15220), .ZN(n11027) );
  INV_X1 U14210 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16276) );
  NAND2_X1 U14211 ( .A1(n11027), .A2(n16276), .ZN(n16246) );
  INV_X1 U14212 ( .A(n11027), .ZN(n11028) );
  NAND2_X1 U14213 ( .A1(n11028), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16247) );
  NOR2_X1 U14214 ( .A1(n11030), .A2(n11029), .ZN(n16266) );
  NOR2_X1 U14215 ( .A1(n16275), .A2(n11031), .ZN(n15735) );
  NOR2_X1 U14216 ( .A1(n16266), .A2(n15735), .ZN(n16245) );
  AND2_X1 U14217 ( .A1(n16247), .A2(n16245), .ZN(n15323) );
  INV_X1 U14218 ( .A(n11032), .ZN(n11033) );
  OR2_X1 U14219 ( .A1(n11034), .A2(n11033), .ZN(n11035) );
  NAND2_X1 U14220 ( .A1(n11069), .A2(n11035), .ZN(n13932) );
  NAND2_X1 U14221 ( .A1(n15220), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11036) );
  OR2_X1 U14222 ( .A1(n13932), .A2(n15240), .ZN(n11037) );
  INV_X1 U14223 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15726) );
  NAND2_X1 U14224 ( .A1(n11037), .A2(n15726), .ZN(n15423) );
  INV_X1 U14225 ( .A(n11038), .ZN(n11040) );
  NOR2_X1 U14226 ( .A1(n12678), .A2(n15112), .ZN(n11039) );
  INV_X1 U14227 ( .A(n11094), .ZN(n11102) );
  AOI21_X1 U14228 ( .B1(n11040), .B2(n11039), .A(n11102), .ZN(n11041) );
  NAND2_X1 U14229 ( .A1(n11041), .A2(n11086), .ZN(n14992) );
  OR2_X1 U14230 ( .A1(n14992), .A2(n15240), .ZN(n11042) );
  INV_X1 U14231 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15604) );
  NAND2_X1 U14232 ( .A1(n11042), .A2(n15604), .ZN(n15336) );
  XNOR2_X1 U14233 ( .A(n11044), .B(n11043), .ZN(n15012) );
  NAND2_X1 U14234 ( .A1(n15012), .A2(n15220), .ZN(n11079) );
  INV_X1 U14235 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n20778) );
  NAND2_X1 U14236 ( .A1(n11079), .A2(n20778), .ZN(n15358) );
  INV_X1 U14237 ( .A(n11045), .ZN(n11046) );
  XNOR2_X1 U14238 ( .A(n11059), .B(n11046), .ZN(n18868) );
  NAND2_X1 U14239 ( .A1(n18868), .A2(n15220), .ZN(n11047) );
  NAND2_X1 U14240 ( .A1(n11047), .A2(n15610), .ZN(n15372) );
  AND2_X1 U14241 ( .A1(n15358), .A2(n15372), .ZN(n15346) );
  NAND2_X1 U14242 ( .A1(n15217), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11048) );
  XNOR2_X1 U14243 ( .A(n11049), .B(n11048), .ZN(n18856) );
  NAND2_X1 U14244 ( .A1(n18856), .A2(n15220), .ZN(n11050) );
  INV_X1 U14245 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15612) );
  NAND2_X1 U14246 ( .A1(n11050), .A2(n15612), .ZN(n15349) );
  AND2_X1 U14247 ( .A1(n15346), .A2(n15349), .ZN(n15334) );
  NAND2_X1 U14248 ( .A1(n15217), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11051) );
  INV_X1 U14249 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n14060) );
  NAND2_X1 U14250 ( .A1(n11062), .A2(n14060), .ZN(n11058) );
  OAI211_X1 U14251 ( .C1(n11062), .C2(n11051), .A(n11094), .B(n11058), .ZN(
        n18881) );
  OR2_X1 U14252 ( .A1(n18881), .A2(n15240), .ZN(n11052) );
  XNOR2_X1 U14253 ( .A(n11052), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15328) );
  NOR2_X1 U14254 ( .A1(n11054), .A2(n18896), .ZN(n11053) );
  MUX2_X1 U14255 ( .A(n11054), .B(n11053), .S(n15217), .Z(n11055) );
  AND2_X1 U14256 ( .A1(n11054), .A2(n18896), .ZN(n11063) );
  INV_X1 U14257 ( .A(n18897), .ZN(n11056) );
  NAND2_X1 U14258 ( .A1(n11056), .A2(n15220), .ZN(n11076) );
  INV_X1 U14259 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15691) );
  NAND2_X1 U14260 ( .A1(n11076), .A2(n15691), .ZN(n15404) );
  INV_X1 U14261 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n11162) );
  NOR2_X1 U14262 ( .A1(n12678), .A2(n11162), .ZN(n11057) );
  NAND2_X1 U14263 ( .A1(n11058), .A2(n11057), .ZN(n11060) );
  NAND2_X1 U14264 ( .A1(n11060), .A2(n11059), .ZN(n15018) );
  OR2_X1 U14265 ( .A1(n15018), .A2(n15240), .ZN(n11061) );
  NAND2_X1 U14266 ( .A1(n11061), .A2(n15652), .ZN(n15331) );
  INV_X1 U14267 ( .A(n11062), .ZN(n11066) );
  INV_X1 U14268 ( .A(n11063), .ZN(n11064) );
  NAND3_X1 U14269 ( .A1(n11064), .A2(P2_EBX_REG_15__SCAN_IN), .A3(n15217), 
        .ZN(n11065) );
  NAND2_X1 U14270 ( .A1(n11066), .A2(n11065), .ZN(n15031) );
  OR2_X1 U14271 ( .A1(n15031), .A2(n15240), .ZN(n11067) );
  NAND2_X1 U14272 ( .A1(n11067), .A2(n15682), .ZN(n15395) );
  XNOR2_X1 U14273 ( .A(n11069), .B(n11068), .ZN(n18907) );
  NAND2_X1 U14274 ( .A1(n18907), .A2(n15220), .ZN(n11071) );
  INV_X1 U14275 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11070) );
  NAND2_X1 U14276 ( .A1(n11071), .A2(n11070), .ZN(n15417) );
  AND4_X1 U14277 ( .A1(n15404), .A2(n15331), .A3(n15395), .A4(n15417), .ZN(
        n11072) );
  NAND4_X1 U14278 ( .A1(n15336), .A2(n15334), .A3(n15328), .A4(n11072), .ZN(
        n11083) );
  OR3_X1 U14279 ( .A1(n14992), .A2(n15240), .A3(n15604), .ZN(n15335) );
  OR3_X1 U14280 ( .A1(n15018), .A2(n15240), .A3(n15652), .ZN(n15330) );
  INV_X1 U14281 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11073) );
  OR3_X1 U14282 ( .A1(n18881), .A2(n15240), .A3(n11073), .ZN(n15329) );
  OR3_X1 U14283 ( .A1(n15031), .A2(n15240), .A3(n15682), .ZN(n15394) );
  AND2_X1 U14284 ( .A1(n15220), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11074) );
  NAND2_X1 U14285 ( .A1(n18907), .A2(n11074), .ZN(n15416) );
  AND4_X1 U14286 ( .A1(n15330), .A2(n15329), .A3(n15394), .A4(n15416), .ZN(
        n11078) );
  AND2_X1 U14287 ( .A1(n15220), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11075) );
  NAND2_X1 U14288 ( .A1(n18856), .A2(n11075), .ZN(n15348) );
  INV_X1 U14289 ( .A(n11076), .ZN(n11077) );
  NAND2_X1 U14290 ( .A1(n11077), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15405) );
  OR2_X1 U14291 ( .A1(n11079), .A2(n20778), .ZN(n15359) );
  INV_X1 U14292 ( .A(n18868), .ZN(n11080) );
  AND2_X1 U14293 ( .A1(n15359), .A2(n15371), .ZN(n15332) );
  INV_X1 U14294 ( .A(n11084), .ZN(n11090) );
  NAND2_X1 U14295 ( .A1(n11086), .A2(n11085), .ZN(n11087) );
  NAND2_X1 U14296 ( .A1(n11090), .A2(n11087), .ZN(n15800) );
  OR2_X1 U14297 ( .A1(n15800), .A2(n15240), .ZN(n11088) );
  INV_X1 U14298 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15587) );
  NAND2_X1 U14299 ( .A1(n11088), .A2(n15587), .ZN(n15314) );
  OR2_X1 U14300 ( .A1(n11088), .A2(n15587), .ZN(n15315) );
  XNOR2_X1 U14301 ( .A(n11090), .B(n11089), .ZN(n16217) );
  NAND2_X1 U14302 ( .A1(n16217), .A2(n15220), .ZN(n11091) );
  XNOR2_X1 U14303 ( .A(n11091), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15307) );
  INV_X1 U14304 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15574) );
  OR2_X1 U14305 ( .A1(n11091), .A2(n15574), .ZN(n11092) );
  INV_X1 U14306 ( .A(n11093), .ZN(n11096) );
  NAND3_X1 U14307 ( .A1(n11096), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n15217), 
        .ZN(n11095) );
  OAI211_X1 U14308 ( .C1(n11096), .C2(P2_EBX_REG_24__SCAN_IN), .A(n11095), .B(
        n11094), .ZN(n14983) );
  OR2_X1 U14309 ( .A1(n14983), .A2(n15240), .ZN(n11097) );
  INV_X1 U14310 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15559) );
  NOR2_X1 U14311 ( .A1(n11097), .A2(n15559), .ZN(n15291) );
  NAND2_X1 U14312 ( .A1(n11097), .A2(n15559), .ZN(n15292) );
  INV_X1 U14313 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n16204) );
  NOR2_X1 U14314 ( .A1(n12678), .A2(n16204), .ZN(n11098) );
  NAND2_X1 U14315 ( .A1(n11105), .A2(n11098), .ZN(n11100) );
  INV_X1 U14316 ( .A(n11099), .ZN(n15219) );
  NAND2_X1 U14317 ( .A1(n11100), .A2(n15219), .ZN(n16205) );
  OR2_X1 U14318 ( .A1(n16205), .A2(n15240), .ZN(n11101) );
  XNOR2_X1 U14319 ( .A(n11101), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15270) );
  NOR2_X1 U14320 ( .A1(n12678), .A2(n9879), .ZN(n11103) );
  AOI21_X1 U14321 ( .B1(n11104), .B2(n11103), .A(n11102), .ZN(n11106) );
  NAND2_X1 U14322 ( .A1(n11106), .A2(n11105), .ZN(n14961) );
  OR2_X1 U14323 ( .A1(n14961), .A2(n15240), .ZN(n11107) );
  NAND2_X1 U14324 ( .A1(n11107), .A2(n10914), .ZN(n15276) );
  NAND2_X1 U14325 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15468) );
  INV_X1 U14326 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15537) );
  OR3_X1 U14327 ( .A1(n16205), .A2(n15240), .A3(n15537), .ZN(n11108) );
  INV_X1 U14328 ( .A(n11109), .ZN(n11110) );
  XNOR2_X1 U14329 ( .A(n14949), .B(n11110), .ZN(n16193) );
  NAND2_X1 U14330 ( .A1(n16193), .A2(n15220), .ZN(n15246) );
  INV_X1 U14331 ( .A(n15246), .ZN(n11111) );
  XOR2_X1 U14332 ( .A(n11112), .B(n15212), .Z(n15510) );
  INV_X1 U14333 ( .A(n11114), .ZN(n11115) );
  INV_X1 U14334 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n11120) );
  NAND2_X1 U14335 ( .A1(n15045), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11119) );
  AOI22_X1 U14336 ( .A1(n11148), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11118) );
  OAI211_X1 U14337 ( .C1(n11120), .C2(n9671), .A(n11119), .B(n11118), .ZN(
        n13245) );
  INV_X1 U14338 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n18953) );
  INV_X4 U14339 ( .A(n11121), .ZN(n15045) );
  NAND2_X1 U14340 ( .A1(n15045), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11123) );
  AOI22_X1 U14341 ( .A1(n11148), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11122) );
  OAI211_X1 U14342 ( .C1(n11204), .C2(n18953), .A(n11123), .B(n11122), .ZN(
        n13250) );
  AOI22_X1 U14343 ( .A1(n11148), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11124) );
  OAI21_X1 U14344 ( .B1(n9671), .B2(n13967), .A(n11124), .ZN(n11125) );
  AOI21_X1 U14345 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15045), .A(
        n11125), .ZN(n13374) );
  NAND2_X1 U14346 ( .A1(n15045), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11131) );
  NAND2_X1 U14347 ( .A1(n11148), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11128) );
  NAND2_X1 U14348 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11127) );
  OAI211_X1 U14349 ( .C1(n13391), .C2(n9671), .A(n11128), .B(n11127), .ZN(
        n11129) );
  INV_X1 U14350 ( .A(n11129), .ZN(n11130) );
  NAND2_X1 U14351 ( .A1(n11131), .A2(n11130), .ZN(n13389) );
  NAND2_X1 U14352 ( .A1(n13373), .A2(n13389), .ZN(n13418) );
  INV_X1 U14353 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n11134) );
  NAND2_X1 U14354 ( .A1(n11148), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11133) );
  NAND2_X1 U14355 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11132) );
  OAI211_X1 U14356 ( .C1(n11134), .C2(n9671), .A(n11133), .B(n11132), .ZN(
        n11135) );
  AOI21_X1 U14357 ( .B1(n15045), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n11135), .ZN(n13417) );
  INV_X1 U14358 ( .A(n11136), .ZN(n13519) );
  NAND2_X1 U14359 ( .A1(n11148), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11138) );
  NAND2_X1 U14360 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11137) );
  OAI211_X1 U14361 ( .C1(n9871), .C2(n9671), .A(n11138), .B(n11137), .ZN(
        n11139) );
  AOI21_X1 U14362 ( .B1(n15045), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n11139), .ZN(n13520) );
  NAND2_X1 U14363 ( .A1(n11148), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11141) );
  NAND2_X1 U14364 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11140) );
  OAI211_X1 U14365 ( .C1(n13528), .C2(n9671), .A(n11141), .B(n11140), .ZN(
        n11142) );
  AOI21_X1 U14366 ( .B1(n15045), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n11142), .ZN(n13525) );
  NAND2_X1 U14367 ( .A1(n15045), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11144) );
  AOI22_X1 U14368 ( .A1(n11148), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11143) );
  OAI211_X1 U14369 ( .C1(n9671), .C2(n10960), .A(n11144), .B(n11143), .ZN(
        n13671) );
  INV_X1 U14370 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n13931) );
  NAND2_X1 U14371 ( .A1(n11148), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11146) );
  NAND2_X1 U14372 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11145) );
  OAI211_X1 U14373 ( .C1(n13931), .C2(n9671), .A(n11146), .B(n11145), .ZN(
        n11147) );
  AOI21_X1 U14374 ( .B1(n15045), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n11147), .ZN(n13667) );
  INV_X1 U14375 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11151) );
  NAND2_X1 U14376 ( .A1(n11148), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11150) );
  NAND2_X1 U14377 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11149) );
  OAI211_X1 U14378 ( .C1(n11151), .C2(n11204), .A(n11150), .B(n11149), .ZN(
        n11152) );
  AOI21_X1 U14379 ( .B1(n15045), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n11152), .ZN(n13897) );
  NAND2_X1 U14380 ( .A1(n15045), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11154) );
  AOI22_X1 U14381 ( .A1(n11148), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11153) );
  OAI211_X1 U14382 ( .C1(n11204), .C2(n18896), .A(n11154), .B(n11153), .ZN(
        n13907) );
  NAND2_X1 U14383 ( .A1(n15045), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11156) );
  AOI22_X1 U14384 ( .A1(n11148), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11155) );
  OAI211_X1 U14385 ( .C1(n11204), .C2(n10962), .A(n11156), .B(n11155), .ZN(
        n14039) );
  NAND2_X1 U14386 ( .A1(n11148), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11158) );
  NAND2_X1 U14387 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11157) );
  OAI211_X1 U14388 ( .C1(n14060), .C2(n11204), .A(n11158), .B(n11157), .ZN(
        n11159) );
  AOI21_X1 U14389 ( .B1(n15045), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11159), .ZN(n14058) );
  NAND2_X1 U14390 ( .A1(n11148), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11161) );
  NAND2_X1 U14391 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11160) );
  OAI211_X1 U14392 ( .C1(n11162), .C2(n11204), .A(n11161), .B(n11160), .ZN(
        n11163) );
  AOI21_X1 U14393 ( .B1(n15045), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11163), .ZN(n14178) );
  NAND2_X1 U14394 ( .A1(n15045), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11165) );
  AOI22_X1 U14395 ( .A1(n11148), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11164) );
  OAI211_X1 U14396 ( .C1(n9671), .C2(n11166), .A(n11165), .B(n11164), .ZN(
        n14188) );
  INV_X1 U14397 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n11169) );
  NAND2_X1 U14398 ( .A1(n11148), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11168) );
  NAND2_X1 U14399 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11167) );
  OAI211_X1 U14400 ( .C1(n11169), .C2(n11204), .A(n11168), .B(n11167), .ZN(
        n11170) );
  AOI21_X1 U14401 ( .B1(n15045), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n11170), .ZN(n14196) );
  INV_X1 U14402 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n11174) );
  NAND2_X1 U14403 ( .A1(n11148), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11173) );
  NAND2_X1 U14404 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11172) );
  OAI211_X1 U14405 ( .C1(n11174), .C2(n11204), .A(n11173), .B(n11172), .ZN(
        n11175) );
  AOI21_X1 U14406 ( .B1(n15045), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11175), .ZN(n15115) );
  NAND2_X1 U14407 ( .A1(n11148), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11177) );
  NAND2_X1 U14408 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11176) );
  OAI211_X1 U14409 ( .C1(n15112), .C2(n11204), .A(n11177), .B(n11176), .ZN(
        n11178) );
  AOI21_X1 U14410 ( .B1(n15045), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11178), .ZN(n14988) );
  NAND2_X1 U14411 ( .A1(n15045), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11180) );
  AOI22_X1 U14412 ( .A1(n11148), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11179) );
  OAI211_X1 U14413 ( .C1(n11204), .C2(n15799), .A(n11180), .B(n11179), .ZN(
        n15101) );
  INV_X1 U14414 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n11183) );
  NAND2_X1 U14415 ( .A1(n11148), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11182) );
  NAND2_X1 U14416 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11181) );
  OAI211_X1 U14417 ( .C1(n11183), .C2(n11204), .A(n11182), .B(n11181), .ZN(
        n11184) );
  AOI21_X1 U14418 ( .B1(n15045), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n11184), .ZN(n15097) );
  NAND2_X1 U14419 ( .A1(n11148), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11186) );
  NAND2_X1 U14420 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11185) );
  OAI211_X1 U14421 ( .C1(n15090), .C2(n11204), .A(n11186), .B(n11185), .ZN(
        n11187) );
  AOI21_X1 U14422 ( .B1(n15045), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11187), .ZN(n14973) );
  NAND2_X1 U14423 ( .A1(n15045), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11191) );
  NOR2_X1 U14424 ( .A1(n9671), .A2(n9879), .ZN(n11189) );
  INV_X1 U14425 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19686) );
  OAI22_X1 U14426 ( .A1(n11126), .A2(n19686), .B1(n19726), .B2(n15282), .ZN(
        n11188) );
  NOR2_X1 U14427 ( .A1(n11189), .A2(n11188), .ZN(n11190) );
  NAND2_X1 U14428 ( .A1(n11191), .A2(n11190), .ZN(n14959) );
  NAND2_X1 U14429 ( .A1(n15045), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11193) );
  AOI22_X1 U14430 ( .A1(n11148), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11192) );
  OAI211_X1 U14431 ( .C1(n11204), .C2(n16204), .A(n11193), .B(n11192), .ZN(
        n15075) );
  INV_X1 U14432 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n11196) );
  NAND2_X1 U14433 ( .A1(n11148), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11195) );
  NAND2_X1 U14434 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11194) );
  OAI211_X1 U14435 ( .C1(n11196), .C2(n11204), .A(n11195), .B(n11194), .ZN(
        n11197) );
  AOI21_X1 U14436 ( .B1(n15045), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11197), .ZN(n14943) );
  NAND2_X1 U14437 ( .A1(n11148), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11199) );
  NAND2_X1 U14438 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11198) );
  OAI211_X1 U14439 ( .C1(n11200), .C2(n11204), .A(n11199), .B(n11198), .ZN(
        n11201) );
  AOI21_X1 U14440 ( .B1(n15045), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11201), .ZN(n15062) );
  NAND2_X1 U14441 ( .A1(n11148), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11203) );
  NAND2_X1 U14442 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11202) );
  OAI211_X1 U14443 ( .C1(n11205), .C2(n11204), .A(n11203), .B(n11202), .ZN(
        n11206) );
  AOI21_X1 U14444 ( .B1(n15045), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11206), .ZN(n11207) );
  INV_X1 U14445 ( .A(n15044), .ZN(n11209) );
  NAND2_X1 U14446 ( .A1(n15065), .A2(n11207), .ZN(n11208) );
  NAND2_X1 U14447 ( .A1(n11209), .A2(n11208), .ZN(n15503) );
  INV_X1 U14448 ( .A(n15503), .ZN(n11221) );
  NAND2_X1 U14449 ( .A1(n19726), .A2(n19737), .ZN(n19708) );
  INV_X1 U14450 ( .A(n19708), .ZN(n14070) );
  OR2_X1 U14451 ( .A1(n19520), .A2(n14070), .ZN(n19736) );
  NAND2_X1 U14452 ( .A1(n19736), .A2(n19762), .ZN(n11210) );
  AND2_X1 U14453 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n11211) );
  INV_X1 U14454 ( .A(n12156), .ZN(n11214) );
  INV_X1 U14455 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n11212) );
  NAND2_X1 U14456 ( .A1(n11212), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11213) );
  NAND2_X1 U14457 ( .A1(n11214), .A2(n11213), .ZN(n19070) );
  NAND2_X1 U14458 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n13773), .ZN(
        n13771) );
  NAND2_X1 U14459 ( .A1(n13926), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13929) );
  NAND2_X1 U14460 ( .A1(n14928), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11217) );
  INV_X1 U14461 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14936) );
  NAND2_X1 U14462 ( .A1(n11217), .A2(n14936), .ZN(n11218) );
  NAND2_X1 U14463 ( .A1(n15237), .A2(n11218), .ZN(n14930) );
  NAND2_X1 U14464 ( .A1(n13328), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15498) );
  NAND2_X1 U14465 ( .A1(n19069), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11219) );
  OAI211_X1 U14466 ( .C1(n16262), .C2(n14930), .A(n15498), .B(n11219), .ZN(
        n11220) );
  OAI21_X1 U14467 ( .B1(n15510), .B2(n19072), .A(n11222), .ZN(n11223) );
  AOI22_X1 U14468 ( .A1(n9635), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11231) );
  AND2_X4 U14469 ( .A1(n11235), .A2(n13575), .ZN(n11960) );
  AND2_X2 U14470 ( .A1(n11232), .A2(n13564), .ZN(n11688) );
  AND2_X2 U14471 ( .A1(n11227), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11233) );
  AND2_X2 U14472 ( .A1(n11233), .A2(n13564), .ZN(n11278) );
  AOI22_X1 U14473 ( .A1(n11530), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11278), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11229) );
  AOI22_X1 U14474 ( .A1(n9586), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11273), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11228) );
  AOI22_X1 U14475 ( .A1(n9632), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11266), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11238) );
  AOI22_X1 U14476 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11237) );
  AND2_X2 U14477 ( .A1(n11235), .A2(n11234), .ZN(n11410) );
  AOI22_X1 U14478 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11236) );
  AOI22_X1 U14479 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11243) );
  AOI22_X1 U14480 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11242) );
  AOI22_X1 U14481 ( .A1(n11250), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11688), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11241) );
  AOI22_X1 U14482 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11240) );
  NAND4_X1 U14483 ( .A1(n11243), .A2(n11242), .A3(n11241), .A4(n11240), .ZN(
        n11249) );
  AOI22_X1 U14484 ( .A1(n11960), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11247) );
  AOI22_X1 U14485 ( .A1(n11530), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11278), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11246) );
  AOI22_X1 U14486 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9645), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11244) );
  NAND4_X1 U14487 ( .A1(n11247), .A2(n11246), .A3(n11245), .A4(n11244), .ZN(
        n11248) );
  AOI22_X1 U14488 ( .A1(n11250), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11300), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11254) );
  AOI22_X1 U14489 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11977), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11253) );
  AOI22_X1 U14490 ( .A1(n11530), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11278), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11252) );
  AOI22_X1 U14491 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11266), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11251) );
  NAND4_X1 U14492 ( .A1(n11254), .A2(n11253), .A3(n11252), .A4(n11251), .ZN(
        n11261) );
  AOI22_X1 U14493 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11259) );
  AOI22_X1 U14494 ( .A1(n11960), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11688), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11258) );
  AOI22_X1 U14495 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11257) );
  AOI22_X1 U14496 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11273), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11256) );
  NAND4_X1 U14497 ( .A1(n11259), .A2(n11258), .A3(n11257), .A4(n11256), .ZN(
        n11260) );
  AOI22_X1 U14498 ( .A1(n11250), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9643), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11265) );
  AOI22_X1 U14499 ( .A1(n11960), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11688), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11264) );
  AOI22_X1 U14500 ( .A1(n11530), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11278), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11263) );
  AOI22_X1 U14501 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9645), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11262) );
  NAND4_X1 U14502 ( .A1(n11265), .A2(n11264), .A3(n11263), .A4(n11262), .ZN(
        n11272) );
  AOI22_X1 U14503 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11270) );
  AOI22_X1 U14504 ( .A1(n9640), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11266), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11269) );
  AOI22_X1 U14505 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11268) );
  AOI22_X1 U14506 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11267) );
  NAND4_X1 U14507 ( .A1(n11270), .A2(n11269), .A3(n11268), .A4(n11267), .ZN(
        n11271) );
  NAND2_X1 U14508 ( .A1(n11960), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11277) );
  NAND2_X1 U14509 ( .A1(n11250), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11276) );
  NAND2_X1 U14510 ( .A1(n11688), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11275) );
  NAND2_X1 U14511 ( .A1(n9645), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11274) );
  NAND2_X1 U14512 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11282) );
  NAND2_X1 U14513 ( .A1(n11706), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11281) );
  NAND2_X1 U14514 ( .A1(n11530), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11280) );
  NAND2_X1 U14515 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11279) );
  NAND2_X1 U14516 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11287) );
  NAND2_X1 U14517 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11286) );
  NAND2_X1 U14518 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11285) );
  NAND2_X1 U14519 ( .A1(n11305), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11284) );
  NAND2_X1 U14520 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11291) );
  NAND2_X1 U14521 ( .A1(n9640), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11290) );
  NAND2_X1 U14522 ( .A1(n11496), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11289) );
  NAND2_X1 U14523 ( .A1(n11266), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11288) );
  NAND2_X1 U14524 ( .A1(n13290), .A2(n11376), .ZN(n11381) );
  NAND2_X1 U14525 ( .A1(n12909), .A2(n11381), .ZN(n11320) );
  NAND2_X1 U14526 ( .A1(n9635), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11299) );
  NAND2_X1 U14527 ( .A1(n11960), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11298) );
  NAND2_X1 U14528 ( .A1(n12018), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11297) );
  NAND2_X1 U14529 ( .A1(n9645), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11296) );
  NAND2_X1 U14530 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n11304) );
  NAND2_X1 U14531 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11303) );
  NAND2_X1 U14532 ( .A1(n11530), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11302) );
  NAND2_X1 U14533 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11301) );
  NAND2_X1 U14534 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11309) );
  NAND2_X1 U14535 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11308) );
  NAND2_X1 U14536 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11307) );
  NAND2_X1 U14537 ( .A1(n11305), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11306) );
  NAND2_X1 U14538 ( .A1(n9632), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11313) );
  NAND2_X1 U14539 ( .A1(n11688), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11312) );
  NAND2_X1 U14540 ( .A1(n11266), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11311) );
  NAND2_X1 U14541 ( .A1(n11496), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11310) );
  NAND2_X1 U14542 ( .A1(n13544), .A2(n11368), .ZN(n11318) );
  NAND2_X1 U14543 ( .A1(n11960), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11324) );
  NAND2_X1 U14544 ( .A1(n11688), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11323) );
  NAND2_X1 U14545 ( .A1(n11250), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11322) );
  NAND2_X1 U14546 ( .A1(n9643), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11321) );
  NAND2_X1 U14547 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11328) );
  NAND2_X1 U14548 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11327) );
  NAND2_X1 U14549 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11326) );
  NAND2_X1 U14550 ( .A1(n11266), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11325) );
  NAND2_X1 U14551 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11332) );
  NAND2_X1 U14552 ( .A1(n11530), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11331) );
  NAND2_X1 U14553 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11330) );
  NAND2_X1 U14554 ( .A1(n9645), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11329) );
  NAND2_X1 U14555 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11336) );
  NAND2_X1 U14556 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11335) );
  NAND2_X1 U14557 ( .A1(n11305), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11334) );
  NAND2_X1 U14558 ( .A1(n11496), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11333) );
  NAND4_X4 U14559 ( .A1(n11340), .A2(n11339), .A3(n11338), .A4(n11337), .ZN(
        n11372) );
  NAND2_X1 U14560 ( .A1(n9637), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11344) );
  NAND2_X1 U14561 ( .A1(n11688), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11343) );
  NAND2_X1 U14562 ( .A1(n9634), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11342) );
  NAND2_X1 U14563 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11348) );
  NAND2_X1 U14564 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11347) );
  NAND2_X1 U14565 ( .A1(n9639), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11346) );
  NAND2_X1 U14566 ( .A1(n11266), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11345) );
  NAND2_X1 U14567 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11352) );
  NAND2_X1 U14568 ( .A1(n11530), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11351) );
  NAND2_X1 U14569 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11350) );
  NAND2_X1 U14570 ( .A1(n11273), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11349) );
  NAND2_X1 U14571 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11356) );
  NAND2_X1 U14572 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11355) );
  NAND2_X1 U14573 ( .A1(n11305), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11354) );
  NAND2_X1 U14574 ( .A1(n11496), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11353) );
  NAND4_X4 U14575 ( .A1(n11360), .A2(n11359), .A3(n11358), .A4(n11357), .ZN(
        n11367) );
  NAND3_X1 U14576 ( .A1(n11373), .A2(n11566), .A3(n12047), .ZN(n13164) );
  INV_X1 U14577 ( .A(n13164), .ZN(n11361) );
  XNOR2_X1 U14578 ( .A(n11362), .B(P1_STATE_REG_2__SCAN_IN), .ZN(n12897) );
  OR2_X1 U14579 ( .A1(n11399), .A2(n11379), .ZN(n11370) );
  NAND2_X1 U14580 ( .A1(n20040), .A2(n11372), .ZN(n12922) );
  INV_X1 U14581 ( .A(n11373), .ZN(n11374) );
  NAND2_X1 U14582 ( .A1(n12911), .A2(n11372), .ZN(n11375) );
  NAND2_X1 U14583 ( .A1(n13163), .A2(n11375), .ZN(n13037) );
  AND4_X2 U14584 ( .A1(n11397), .A2(n13032), .A3(n13036), .A4(n13037), .ZN(
        n11384) );
  NAND2_X1 U14585 ( .A1(n20048), .A2(n12045), .ZN(n11377) );
  NAND2_X1 U14586 ( .A1(n11403), .A2(n14302), .ZN(n11383) );
  NAND2_X1 U14587 ( .A1(n9770), .A2(n20024), .ZN(n11382) );
  NAND3_X1 U14588 ( .A1(n11384), .A2(n11383), .A3(n11382), .ZN(n13047) );
  NAND2_X1 U14589 ( .A1(n13047), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11385) );
  NAND2_X1 U14590 ( .A1(n11464), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11388) );
  NAND2_X1 U14591 ( .A1(n20493), .A2(n20415), .ZN(n20384) );
  NAND2_X1 U14592 ( .A1(n20384), .A2(n20489), .ZN(n20326) );
  OR2_X1 U14593 ( .A1(n15843), .A2(n20493), .ZN(n11462) );
  OAI21_X1 U14594 ( .B1(n13266), .B2(n20326), .A(n11462), .ZN(n11386) );
  INV_X1 U14595 ( .A(n11386), .ZN(n11387) );
  INV_X1 U14596 ( .A(n11389), .ZN(n11390) );
  NAND2_X1 U14597 ( .A1(n11464), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11392) );
  MUX2_X1 U14598 ( .A(n15843), .B(n13266), .S(n20415), .Z(n11391) );
  NAND2_X1 U14599 ( .A1(n11393), .A2(n12949), .ZN(n11395) );
  MUX2_X1 U14600 ( .A(n11395), .B(n11394), .S(n13627), .Z(n11407) );
  OR2_X1 U14601 ( .A1(n13032), .A2(n12045), .ZN(n11396) );
  NAND2_X1 U14602 ( .A1(n11397), .A2(n11396), .ZN(n13043) );
  INV_X1 U14603 ( .A(n11398), .ZN(n11400) );
  INV_X1 U14604 ( .A(n11399), .ZN(n12877) );
  NAND2_X1 U14605 ( .A1(n11400), .A2(n12877), .ZN(n11401) );
  NAND4_X1 U14606 ( .A1(n11401), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n14880), 
        .A4(n13037), .ZN(n11402) );
  NOR2_X1 U14607 ( .A1(n13043), .A2(n11402), .ZN(n11405) );
  NAND3_X1 U14608 ( .A1(n11403), .A2(n11367), .A3(n14302), .ZN(n11404) );
  AND2_X1 U14609 ( .A1(n11405), .A2(n11404), .ZN(n11406) );
  NAND2_X1 U14610 ( .A1(n11438), .A2(n11436), .ZN(n11408) );
  INV_X1 U14611 ( .A(n11490), .ZN(n11432) );
  AOI22_X1 U14612 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(n9594), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11414) );
  AOI22_X1 U14613 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11413) );
  AOI22_X1 U14614 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11412) );
  AOI22_X1 U14615 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11411) );
  NAND4_X1 U14616 ( .A1(n11414), .A2(n11413), .A3(n11412), .A4(n11411), .ZN(
        n11420) );
  AOI22_X1 U14617 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11418) );
  AOI22_X1 U14618 ( .A1(n11960), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11994), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11417) );
  AOI22_X1 U14619 ( .A1(n12020), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11266), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11416) );
  AOI22_X1 U14620 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11415) );
  NAND4_X1 U14621 ( .A1(n11418), .A2(n11417), .A3(n11416), .A4(n11415), .ZN(
        n11419) );
  NAND2_X1 U14622 ( .A1(n11432), .A2(n12809), .ZN(n11421) );
  AOI22_X1 U14623 ( .A1(n11960), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11994), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11425) );
  AOI22_X1 U14624 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11424) );
  AOI22_X1 U14625 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14626 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11273), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11422) );
  NAND4_X1 U14627 ( .A1(n11425), .A2(n11424), .A3(n11423), .A4(n11422), .ZN(
        n11431) );
  AOI22_X1 U14628 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11429) );
  AOI22_X1 U14629 ( .A1(n9639), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11266), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11428) );
  AOI22_X1 U14630 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U14631 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11426) );
  NAND4_X1 U14632 ( .A1(n11429), .A2(n11428), .A3(n11427), .A4(n11426), .ZN(
        n11430) );
  NAND2_X1 U14633 ( .A1(n11432), .A2(n11439), .ZN(n11440) );
  NAND2_X1 U14634 ( .A1(n12105), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11435) );
  INV_X1 U14635 ( .A(n12809), .ZN(n11433) );
  OR2_X1 U14636 ( .A1(n11491), .A2(n11433), .ZN(n11434) );
  NAND2_X1 U14637 ( .A1(n11568), .A2(n20556), .ZN(n11455) );
  INV_X1 U14638 ( .A(n11440), .ZN(n11452) );
  AOI22_X1 U14639 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11445) );
  AOI22_X1 U14640 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12028), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11444) );
  AOI22_X1 U14641 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11443) );
  AOI22_X1 U14642 ( .A1(n11994), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11442) );
  NAND4_X1 U14643 ( .A1(n11445), .A2(n11444), .A3(n11443), .A4(n11442), .ZN(
        n11451) );
  AOI22_X1 U14644 ( .A1(n11960), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11449) );
  AOI22_X1 U14645 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11448) );
  AOI22_X1 U14646 ( .A1(n11977), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11266), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11447) );
  AOI22_X1 U14647 ( .A1(n12018), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11446) );
  NAND4_X1 U14648 ( .A1(n11449), .A2(n11448), .A3(n11447), .A4(n11446), .ZN(
        n11450) );
  MUX2_X1 U14649 ( .A(n12804), .B(n11452), .S(n12814), .Z(n11453) );
  INV_X1 U14650 ( .A(n11453), .ZN(n11454) );
  AOI21_X1 U14651 ( .B1(n20044), .B2(n12876), .A(n20556), .ZN(n11457) );
  NAND2_X1 U14652 ( .A1(n20024), .A2(n12814), .ZN(n11456) );
  INV_X1 U14653 ( .A(n11459), .ZN(n11460) );
  AND2_X1 U14654 ( .A1(n11462), .A2(n11225), .ZN(n11463) );
  NOR2_X1 U14655 ( .A1(n15843), .A2(n20274), .ZN(n11465) );
  AOI21_X1 U14656 ( .B1(n11464), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11465), .ZN(n11469) );
  INV_X1 U14657 ( .A(n13266), .ZN(n11487) );
  XNOR2_X1 U14658 ( .A(n20489), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20029) );
  NAND2_X1 U14659 ( .A1(n11487), .A2(n20029), .ZN(n11467) );
  NAND2_X1 U14660 ( .A1(n11469), .A2(n11467), .ZN(n11466) );
  AOI22_X1 U14661 ( .A1(n11960), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11688), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11473) );
  AOI22_X1 U14662 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11472) );
  AOI22_X1 U14663 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11471) );
  AOI22_X1 U14664 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11470) );
  NAND4_X1 U14665 ( .A1(n11473), .A2(n11472), .A3(n11471), .A4(n11470), .ZN(
        n11479) );
  AOI22_X1 U14666 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11477) );
  AOI22_X1 U14667 ( .A1(n9632), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11266), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11476) );
  INV_X1 U14668 ( .A(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n20742) );
  AOI22_X1 U14669 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11475) );
  AOI22_X1 U14670 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11474) );
  NAND4_X1 U14671 ( .A1(n11477), .A2(n11476), .A3(n11475), .A4(n11474), .ZN(
        n11478) );
  INV_X1 U14672 ( .A(n11491), .ZN(n11480) );
  AOI22_X1 U14673 ( .A1(n11480), .A2(n12823), .B1(n12105), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11481) );
  NAND2_X1 U14674 ( .A1(n11464), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11489) );
  INV_X1 U14675 ( .A(n20489), .ZN(n11485) );
  INV_X1 U14676 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20655) );
  NAND2_X1 U14677 ( .A1(n20655), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20209) );
  INV_X1 U14678 ( .A(n20209), .ZN(n11484) );
  NAND2_X1 U14679 ( .A1(n11485), .A2(n11484), .ZN(n20240) );
  OAI21_X1 U14680 ( .B1(n20489), .B2(n20274), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11486) );
  NAND2_X1 U14681 ( .A1(n20240), .A2(n11486), .ZN(n20275) );
  INV_X1 U14682 ( .A(n15843), .ZN(n15836) );
  AOI22_X1 U14683 ( .A1(n20275), .A2(n11487), .B1(n15836), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11488) );
  AOI22_X1 U14684 ( .A1(n11960), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11688), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11495) );
  AOI22_X1 U14685 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9644), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11494) );
  AOI22_X1 U14686 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11493) );
  AOI22_X1 U14687 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11492) );
  NAND4_X1 U14688 ( .A1(n11495), .A2(n11494), .A3(n11493), .A4(n11492), .ZN(
        n11502) );
  AOI22_X1 U14689 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11500) );
  AOI22_X1 U14690 ( .A1(n9640), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11499) );
  AOI22_X1 U14691 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11498) );
  AOI22_X1 U14692 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11497) );
  NAND4_X1 U14693 ( .A1(n11500), .A2(n11499), .A3(n11498), .A4(n11497), .ZN(
        n11501) );
  AOI22_X1 U14694 ( .A1(n12092), .A2(n12847), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n12105), .ZN(n11503) );
  AOI22_X1 U14695 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11688), .B1(
        n11960), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11508) );
  AOI22_X1 U14696 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12026), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U14697 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n9592), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11506) );
  AOI22_X1 U14698 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11505) );
  NAND4_X1 U14699 ( .A1(n11508), .A2(n11507), .A3(n11506), .A4(n11505), .ZN(
        n11514) );
  AOI22_X1 U14700 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U14701 ( .A1(n9639), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11511) );
  AOI22_X1 U14702 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11510) );
  AOI22_X1 U14703 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11509) );
  NAND4_X1 U14704 ( .A1(n11512), .A2(n11511), .A3(n11510), .A4(n11509), .ZN(
        n11513) );
  NAND2_X1 U14705 ( .A1(n12092), .A2(n12846), .ZN(n11516) );
  NAND2_X1 U14706 ( .A1(n12105), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11515) );
  NAND2_X1 U14707 ( .A1(n11516), .A2(n11515), .ZN(n11585) );
  AOI22_X1 U14708 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11521) );
  AOI22_X1 U14709 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11960), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U14710 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11519) );
  AOI22_X1 U14711 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11518) );
  NAND4_X1 U14712 ( .A1(n11521), .A2(n11520), .A3(n11519), .A4(n11518), .ZN(
        n11527) );
  AOI22_X1 U14713 ( .A1(n11994), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12028), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11525) );
  AOI22_X1 U14714 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11524) );
  AOI22_X1 U14715 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U14716 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11522) );
  NAND4_X1 U14717 ( .A1(n11525), .A2(n11524), .A3(n11523), .A4(n11522), .ZN(
        n11526) );
  NAND2_X1 U14718 ( .A1(n12092), .A2(n12857), .ZN(n11529) );
  NAND2_X1 U14719 ( .A1(n12105), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11528) );
  NAND2_X1 U14720 ( .A1(n11529), .A2(n11528), .ZN(n11595) );
  AOI22_X1 U14721 ( .A1(n11960), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11688), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11534) );
  AOI22_X1 U14722 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9644), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11533) );
  INV_X1 U14723 ( .A(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n20739) );
  AOI22_X1 U14724 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11532) );
  AOI22_X1 U14725 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11531) );
  NAND4_X1 U14726 ( .A1(n11534), .A2(n11533), .A3(n11532), .A4(n11531), .ZN(
        n11540) );
  AOI22_X1 U14727 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U14728 ( .A1(n11977), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11537) );
  AOI22_X1 U14729 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U14730 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11535) );
  NAND4_X1 U14731 ( .A1(n11538), .A2(n11537), .A3(n11536), .A4(n11535), .ZN(
        n11539) );
  AOI22_X1 U14732 ( .A1(n12092), .A2(n12868), .B1(n12105), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11602) );
  NAND2_X1 U14733 ( .A1(n12092), .A2(n12876), .ZN(n11543) );
  NAND2_X1 U14734 ( .A1(n12105), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11542) );
  NAND2_X1 U14735 ( .A1(n11543), .A2(n11542), .ZN(n11544) );
  NAND2_X1 U14736 ( .A1(n12866), .A2(n11731), .ZN(n11550) );
  INV_X1 U14737 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n14011) );
  NAND2_X1 U14738 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11579), .ZN(
        n11596) );
  NAND2_X1 U14739 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11545) );
  NOR2_X1 U14740 ( .A1(n11596), .A2(n11545), .ZN(n11604) );
  NOR2_X1 U14741 ( .A1(n11606), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11546) );
  OR2_X1 U14742 ( .A1(n11628), .A2(n11546), .ZN(n19839) );
  AOI22_X1 U14743 ( .A1(n19839), .A2(n13621), .B1(n12041), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11547) );
  NAND2_X1 U14744 ( .A1(n13033), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11590) );
  XNOR2_X1 U14745 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13660) );
  AOI21_X1 U14746 ( .B1(n11574), .B2(n13660), .A(n12041), .ZN(n11553) );
  NAND2_X1 U14747 ( .A1(n12042), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11552) );
  OAI211_X1 U14748 ( .C1(n11590), .C2(n11554), .A(n11553), .B(n11552), .ZN(
        n11555) );
  INV_X1 U14749 ( .A(n11555), .ZN(n11556) );
  NAND2_X1 U14750 ( .A1(n12041), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11578) );
  INV_X1 U14751 ( .A(n13458), .ZN(n11577) );
  XNOR2_X2 U14752 ( .A(n11558), .B(n11557), .ZN(n13601) );
  NAND2_X1 U14753 ( .A1(n13601), .A2(n11731), .ZN(n11563) );
  NAND2_X1 U14754 ( .A1(n12042), .A2(P1_EAX_REG_1__SCAN_IN), .ZN(n11560) );
  NAND2_X1 U14755 ( .A1(n20417), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11559) );
  OAI211_X1 U14756 ( .C1(n11590), .C2(n11225), .A(n11560), .B(n11559), .ZN(
        n11561) );
  INV_X1 U14757 ( .A(n11561), .ZN(n11562) );
  NAND2_X1 U14758 ( .A1(n11563), .A2(n11562), .ZN(n13262) );
  NAND2_X1 U14759 ( .A1(n12818), .A2(n11566), .ZN(n11567) );
  NAND2_X1 U14760 ( .A1(n11567), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13279) );
  NAND2_X1 U14761 ( .A1(n11569), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11571) );
  NAND2_X1 U14762 ( .A1(n20417), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11570) );
  OAI211_X1 U14763 ( .C1(n11590), .C2(n11226), .A(n11571), .B(n11570), .ZN(
        n11572) );
  AOI21_X1 U14764 ( .B1(n11568), .B2(n11731), .A(n11572), .ZN(n11573) );
  OR2_X1 U14765 ( .A1(n13279), .A2(n11573), .ZN(n13280) );
  INV_X1 U14766 ( .A(n11573), .ZN(n13281) );
  OR2_X1 U14767 ( .A1(n13281), .A2(n12014), .ZN(n11575) );
  NAND2_X1 U14768 ( .A1(n13280), .A2(n11575), .ZN(n13261) );
  NAND2_X1 U14769 ( .A1(n11577), .A2(n11576), .ZN(n13457) );
  NAND2_X1 U14770 ( .A1(n20642), .A2(n11731), .ZN(n11584) );
  OAI21_X1 U14771 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11579), .A(
        n11596), .ZN(n13767) );
  AOI22_X1 U14772 ( .A1(n13621), .A2(n13767), .B1(n12041), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11581) );
  NAND2_X1 U14773 ( .A1(n12042), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11580) );
  OAI211_X1 U14774 ( .C1(n11590), .C2(n11227), .A(n11581), .B(n11580), .ZN(
        n11582) );
  INV_X1 U14775 ( .A(n11582), .ZN(n11583) );
  NAND2_X1 U14776 ( .A1(n11584), .A2(n11583), .ZN(n13533) );
  NAND2_X1 U14777 ( .A1(n13532), .A2(n13533), .ZN(n13612) );
  INV_X1 U14778 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11587) );
  XNOR2_X1 U14779 ( .A(n11587), .B(n11596), .ZN(n19971) );
  NAND2_X1 U14780 ( .A1(n20417), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11589) );
  NAND2_X1 U14781 ( .A1(n12042), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11588) );
  OAI211_X1 U14782 ( .C1(n11590), .C2(n16158), .A(n11589), .B(n11588), .ZN(
        n11591) );
  MUX2_X1 U14783 ( .A(n19971), .B(n11591), .S(n12014), .Z(n11592) );
  AOI21_X1 U14784 ( .B1(n12838), .B2(n11731), .A(n11592), .ZN(n13611) );
  INV_X1 U14785 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n11600) );
  INV_X1 U14786 ( .A(n11596), .ZN(n11597) );
  AOI21_X1 U14787 ( .B1(n11597), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11598) );
  OR2_X1 U14788 ( .A1(n11598), .A2(n11604), .ZN(n19874) );
  AOI22_X1 U14789 ( .A1(n19874), .A2(n13621), .B1(n12041), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11599) );
  OAI21_X1 U14790 ( .B1(n11905), .B2(n11600), .A(n11599), .ZN(n11601) );
  AOI21_X1 U14791 ( .B1(n12845), .B2(n11731), .A(n11601), .ZN(n13679) );
  NAND2_X1 U14792 ( .A1(n11603), .A2(n11602), .ZN(n12855) );
  INV_X1 U14793 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11610) );
  NOR2_X1 U14794 ( .A1(n11604), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11605) );
  OR2_X1 U14795 ( .A1(n11606), .A2(n11605), .ZN(n19850) );
  INV_X1 U14796 ( .A(n12041), .ZN(n11607) );
  INV_X1 U14797 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19848) );
  NOR2_X1 U14798 ( .A1(n11607), .A2(n19848), .ZN(n11608) );
  AOI21_X1 U14799 ( .B1(n19850), .B2(n13621), .A(n11608), .ZN(n11609) );
  OAI21_X1 U14800 ( .B1(n11905), .B2(n11610), .A(n11609), .ZN(n11611) );
  AOI21_X1 U14801 ( .B1(n12855), .B2(n11731), .A(n11611), .ZN(n14001) );
  INV_X1 U14802 ( .A(n14007), .ZN(n11627) );
  AOI22_X1 U14803 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9637), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11615) );
  AOI22_X1 U14804 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11613) );
  AOI22_X1 U14805 ( .A1(n11994), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11612) );
  NAND4_X1 U14806 ( .A1(n11615), .A2(n11614), .A3(n11613), .A4(n11612), .ZN(
        n11621) );
  AOI22_X1 U14807 ( .A1(n9640), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11619) );
  AOI22_X1 U14808 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14809 ( .A1(n12020), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U14810 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11616) );
  NAND4_X1 U14811 ( .A1(n11619), .A2(n11618), .A3(n11617), .A4(n11616), .ZN(
        n11620) );
  OAI21_X1 U14812 ( .B1(n11621), .B2(n11620), .A(n11731), .ZN(n11625) );
  NAND2_X1 U14813 ( .A1(n12042), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11624) );
  XNOR2_X1 U14814 ( .A(n11628), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n19824) );
  NAND2_X1 U14815 ( .A1(n19824), .A2(n13621), .ZN(n11623) );
  NAND2_X1 U14816 ( .A1(n12041), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11622) );
  NAND2_X1 U14817 ( .A1(n11628), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11654) );
  XOR2_X1 U14818 ( .A(n19809), .B(n11654), .Z(n19813) );
  AOI22_X1 U14819 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11632) );
  AOI22_X1 U14820 ( .A1(n9632), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U14821 ( .A1(n11994), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11629) );
  NAND4_X1 U14822 ( .A1(n11632), .A2(n11631), .A3(n11630), .A4(n11629), .ZN(
        n11638) );
  AOI22_X1 U14823 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11636) );
  AOI22_X1 U14824 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U14825 ( .A1(n9637), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11634) );
  AOI22_X1 U14826 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11633) );
  NAND4_X1 U14827 ( .A1(n11636), .A2(n11635), .A3(n11634), .A4(n11633), .ZN(
        n11637) );
  OR2_X1 U14828 ( .A1(n11638), .A2(n11637), .ZN(n11639) );
  AOI22_X1 U14829 ( .A1(n11731), .A2(n11639), .B1(n12041), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11641) );
  NAND2_X1 U14830 ( .A1(n12042), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11640) );
  OAI211_X1 U14831 ( .C1(n19813), .C2(n12014), .A(n11641), .B(n11640), .ZN(
        n11642) );
  INV_X1 U14832 ( .A(n11642), .ZN(n14140) );
  AOI22_X1 U14833 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U14834 ( .A1(n11960), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11688), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14835 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14836 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11644) );
  NAND4_X1 U14837 ( .A1(n11647), .A2(n11646), .A3(n11645), .A4(n11644), .ZN(
        n11653) );
  AOI22_X1 U14838 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11650) );
  AOI22_X1 U14839 ( .A1(n9640), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11649) );
  AOI22_X1 U14840 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11648) );
  NAND4_X1 U14841 ( .A1(n11651), .A2(n11650), .A3(n11649), .A4(n11648), .ZN(
        n11652) );
  NOR2_X1 U14842 ( .A1(n11653), .A2(n11652), .ZN(n11657) );
  XNOR2_X1 U14843 ( .A(n11658), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14731) );
  NAND2_X1 U14844 ( .A1(n14731), .A2(n13621), .ZN(n11656) );
  AOI22_X1 U14845 ( .A1(n12042), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n12041), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11655) );
  OAI211_X1 U14846 ( .C1(n11657), .C2(n9971), .A(n11656), .B(n11655), .ZN(
        n14129) );
  NAND2_X1 U14847 ( .A1(n12042), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n11661) );
  OAI21_X1 U14848 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11659), .A(
        n11673), .ZN(n16042) );
  AOI22_X1 U14849 ( .A1(n13621), .A2(n16042), .B1(n12041), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11660) );
  NAND2_X1 U14850 ( .A1(n11661), .A2(n11660), .ZN(n14442) );
  AOI22_X1 U14851 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11665) );
  AOI22_X1 U14852 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11664) );
  AOI22_X1 U14853 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11662) );
  NAND4_X1 U14854 ( .A1(n11665), .A2(n11664), .A3(n11663), .A4(n11662), .ZN(
        n11671) );
  AOI22_X1 U14855 ( .A1(n9637), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11688), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11669) );
  AOI22_X1 U14856 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11668) );
  AOI22_X1 U14857 ( .A1(n12020), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U14858 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11666) );
  NAND4_X1 U14859 ( .A1(n11669), .A2(n11668), .A3(n11667), .A4(n11666), .ZN(
        n11670) );
  OR2_X1 U14860 ( .A1(n11671), .A2(n11670), .ZN(n11672) );
  XOR2_X1 U14861 ( .A(n14455), .B(n11705), .Z(n14725) );
  AOI22_X1 U14862 ( .A1(n11977), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11677) );
  AOI22_X1 U14863 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9637), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14864 ( .A1(n11994), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11675) );
  AOI22_X1 U14865 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11674) );
  NAND4_X1 U14866 ( .A1(n11677), .A2(n11676), .A3(n11675), .A4(n11674), .ZN(
        n11683) );
  AOI22_X1 U14867 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11681) );
  AOI22_X1 U14868 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U14869 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U14870 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11678) );
  NAND4_X1 U14871 ( .A1(n11681), .A2(n11680), .A3(n11679), .A4(n11678), .ZN(
        n11682) );
  OR2_X1 U14872 ( .A1(n11683), .A2(n11682), .ZN(n11684) );
  AOI22_X1 U14873 ( .A1(n11731), .A2(n11684), .B1(n12041), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11686) );
  NAND2_X1 U14874 ( .A1(n12042), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11685) );
  OAI211_X1 U14875 ( .C1(n14725), .C2(n12014), .A(n11686), .B(n11685), .ZN(
        n14445) );
  XOR2_X1 U14876 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11687), .Z(
        n16031) );
  AOI22_X1 U14877 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9639), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U14878 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11960), .B1(
        n11994), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11691) );
  AOI22_X1 U14879 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12027), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11690) );
  AOI22_X1 U14880 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11689) );
  NAND4_X1 U14881 ( .A1(n11692), .A2(n11691), .A3(n11690), .A4(n11689), .ZN(
        n11698) );
  AOI22_X1 U14882 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12026), .B1(
        n12028), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U14883 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n9592), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14884 ( .A1(n12025), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14885 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11693) );
  NAND4_X1 U14886 ( .A1(n11696), .A2(n11695), .A3(n11694), .A4(n11693), .ZN(
        n11697) );
  OAI21_X1 U14887 ( .B1(n11698), .B2(n11697), .A(n11731), .ZN(n11701) );
  NAND2_X1 U14888 ( .A1(n12042), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11700) );
  NAND2_X1 U14889 ( .A1(n12041), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11699) );
  AND3_X1 U14890 ( .A1(n11701), .A2(n11700), .A3(n11699), .ZN(n11702) );
  OAI21_X1 U14891 ( .B1(n16031), .B2(n12014), .A(n11702), .ZN(n14516) );
  AND2_X1 U14892 ( .A1(n14445), .A2(n14516), .ZN(n11703) );
  NAND2_X1 U14893 ( .A1(n11704), .A2(n11703), .ZN(n14444) );
  XNOR2_X1 U14894 ( .A(n11722), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15962) );
  AOI22_X1 U14895 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11710) );
  AOI22_X1 U14896 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U14897 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11708) );
  AOI22_X1 U14898 ( .A1(n12018), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11707) );
  NAND4_X1 U14899 ( .A1(n11710), .A2(n11709), .A3(n11708), .A4(n11707), .ZN(
        n11716) );
  AOI22_X1 U14900 ( .A1(n11994), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11714) );
  AOI22_X1 U14901 ( .A1(n9637), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12028), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U14902 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U14903 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11711) );
  NAND4_X1 U14904 ( .A1(n11714), .A2(n11713), .A3(n11712), .A4(n11711), .ZN(
        n11715) );
  OAI21_X1 U14905 ( .B1(n11716), .B2(n11715), .A(n11731), .ZN(n11719) );
  NAND2_X1 U14906 ( .A1(n12042), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11718) );
  NAND2_X1 U14907 ( .A1(n12041), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11717) );
  NAND3_X1 U14908 ( .A1(n11719), .A2(n11718), .A3(n11717), .ZN(n11720) );
  AOI21_X1 U14909 ( .B1(n15962), .B2(n13621), .A(n11720), .ZN(n14506) );
  XOR2_X1 U14910 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n11740), .Z(
        n16021) );
  INV_X1 U14911 ( .A(n16021), .ZN(n11738) );
  AOI22_X1 U14912 ( .A1(n9632), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11726) );
  AOI22_X1 U14913 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11960), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11725) );
  AOI22_X1 U14914 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11724) );
  AOI22_X1 U14915 ( .A1(n11994), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11723) );
  NAND4_X1 U14916 ( .A1(n11726), .A2(n11725), .A3(n11724), .A4(n11723), .ZN(
        n11733) );
  AOI22_X1 U14917 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11730) );
  AOI22_X1 U14918 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11729) );
  AOI22_X1 U14919 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11728) );
  AOI22_X1 U14920 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11727) );
  NAND4_X1 U14921 ( .A1(n11730), .A2(n11729), .A3(n11728), .A4(n11727), .ZN(
        n11732) );
  OAI21_X1 U14922 ( .B1(n11733), .B2(n11732), .A(n11731), .ZN(n11736) );
  NAND2_X1 U14923 ( .A1(n12042), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11735) );
  NAND2_X1 U14924 ( .A1(n12041), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11734) );
  NAND3_X1 U14925 ( .A1(n11736), .A2(n11735), .A3(n11734), .ZN(n11737) );
  AOI21_X1 U14926 ( .B1(n11738), .B2(n13621), .A(n11737), .ZN(n14500) );
  INV_X1 U14927 ( .A(n14500), .ZN(n11739) );
  INV_X1 U14928 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11741) );
  XNOR2_X1 U14929 ( .A(n11758), .B(n11741), .ZN(n15950) );
  NAND2_X1 U14930 ( .A1(n15950), .A2(n13621), .ZN(n11757) );
  AOI22_X1 U14931 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12028), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11745) );
  AOI22_X1 U14932 ( .A1(n11994), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11744) );
  AOI22_X1 U14933 ( .A1(n9643), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11743) );
  AOI22_X1 U14934 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11742) );
  NAND4_X1 U14935 ( .A1(n11745), .A2(n11744), .A3(n11743), .A4(n11742), .ZN(
        n11753) );
  AOI22_X1 U14936 ( .A1(n9639), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9637), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11751) );
  NAND2_X1 U14937 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11747) );
  NAND2_X1 U14938 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11746) );
  AND3_X1 U14939 ( .A1(n11747), .A2(n11746), .A3(n12014), .ZN(n11750) );
  AOI22_X1 U14940 ( .A1(n12025), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11749) );
  AOI22_X1 U14941 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11748) );
  NAND4_X1 U14942 ( .A1(n11751), .A2(n11750), .A3(n11749), .A4(n11748), .ZN(
        n11752) );
  NAND2_X1 U14943 ( .A1(n12011), .A2(n12014), .ZN(n11851) );
  OAI21_X1 U14944 ( .B1(n11753), .B2(n11752), .A(n11851), .ZN(n11755) );
  AOI22_X1 U14945 ( .A1(n12042), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20417), .ZN(n11754) );
  NAND2_X1 U14946 ( .A1(n11755), .A2(n11754), .ZN(n11756) );
  NAND2_X1 U14947 ( .A1(n11757), .A2(n11756), .ZN(n14492) );
  XOR2_X1 U14948 ( .A(n15933), .B(n11771), .Z(n16016) );
  AOI22_X1 U14949 ( .A1(n12042), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n12041), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11770) );
  AOI22_X1 U14950 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11761) );
  AOI22_X1 U14951 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U14952 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11759) );
  NAND4_X1 U14953 ( .A1(n11762), .A2(n11761), .A3(n11760), .A4(n11759), .ZN(
        n11768) );
  AOI22_X1 U14954 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11766) );
  AOI22_X1 U14955 ( .A1(n11688), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11765) );
  AOI22_X1 U14956 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U14957 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11763) );
  NAND4_X1 U14958 ( .A1(n11766), .A2(n11765), .A3(n11764), .A4(n11763), .ZN(
        n11767) );
  OAI21_X1 U14959 ( .B1(n11768), .B2(n11767), .A(n12037), .ZN(n11769) );
  OAI211_X1 U14960 ( .C1(n16016), .C2(n12014), .A(n11770), .B(n11769), .ZN(
        n15935) );
  XNOR2_X1 U14961 ( .A(n11789), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15929) );
  NAND2_X1 U14962 ( .A1(n15929), .A2(n13621), .ZN(n11786) );
  AOI22_X1 U14963 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U14964 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11278), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U14965 ( .A1(n11994), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11772) );
  NAND4_X1 U14966 ( .A1(n11775), .A2(n11774), .A3(n11773), .A4(n11772), .ZN(
        n11781) );
  AOI22_X1 U14967 ( .A1(n11960), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11779) );
  AOI22_X1 U14968 ( .A1(n11977), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11778) );
  AOI22_X1 U14969 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11777) );
  AOI22_X1 U14970 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11776) );
  NAND4_X1 U14971 ( .A1(n11779), .A2(n11778), .A3(n11777), .A4(n11776), .ZN(
        n11780) );
  NOR2_X1 U14972 ( .A1(n11781), .A2(n11780), .ZN(n11784) );
  AOI21_X1 U14973 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15926), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11782) );
  AOI21_X1 U14974 ( .B1(n12042), .B2(P1_EAX_REG_18__SCAN_IN), .A(n11782), .ZN(
        n11783) );
  OAI21_X1 U14975 ( .B1(n12011), .B2(n11784), .A(n11783), .ZN(n11785) );
  NAND2_X1 U14976 ( .A1(n11786), .A2(n11785), .ZN(n14486) );
  NAND2_X1 U14977 ( .A1(n11788), .A2(n11787), .ZN(n14683) );
  OAI21_X1 U14978 ( .B1(n11790), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n11822), .ZN(n15915) );
  OR2_X1 U14979 ( .A1(n15915), .A2(n12014), .ZN(n11805) );
  AOI22_X1 U14980 ( .A1(n9640), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11794) );
  AOI22_X1 U14981 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11793) );
  AOI22_X1 U14982 ( .A1(n11994), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11792) );
  AOI22_X1 U14983 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11791) );
  NAND4_X1 U14984 ( .A1(n11794), .A2(n11793), .A3(n11792), .A4(n11791), .ZN(
        n11800) );
  AOI22_X1 U14985 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11278), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11797) );
  AOI22_X1 U14986 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11796) );
  AOI22_X1 U14987 ( .A1(n9637), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11795) );
  NAND4_X1 U14988 ( .A1(n11798), .A2(n11797), .A3(n11796), .A4(n11795), .ZN(
        n11799) );
  NOR2_X1 U14989 ( .A1(n11800), .A2(n11799), .ZN(n11803) );
  INV_X1 U14990 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20640) );
  OAI21_X1 U14991 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n20640), .A(
        n20417), .ZN(n11802) );
  NAND2_X1 U14992 ( .A1(n12042), .A2(P1_EAX_REG_19__SCAN_IN), .ZN(n11801) );
  OAI211_X1 U14993 ( .C1(n12011), .C2(n11803), .A(n11802), .B(n11801), .ZN(
        n11804) );
  NAND2_X1 U14994 ( .A1(n11805), .A2(n11804), .ZN(n14682) );
  XNOR2_X1 U14995 ( .A(n11822), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15912) );
  AOI22_X1 U14996 ( .A1(n9637), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11278), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11811) );
  NAND2_X1 U14997 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11807) );
  NAND2_X1 U14998 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11806) );
  AND3_X1 U14999 ( .A1(n11807), .A2(n11806), .A3(n12014), .ZN(n11810) );
  AOI22_X1 U15000 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12025), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11809) );
  AOI22_X1 U15001 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12028), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11808) );
  NAND4_X1 U15002 ( .A1(n11811), .A2(n11810), .A3(n11809), .A4(n11808), .ZN(
        n11817) );
  AOI22_X1 U15003 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12026), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11815) );
  AOI22_X1 U15004 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11813) );
  AOI22_X1 U15005 ( .A1(n11994), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11273), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11812) );
  NAND4_X1 U15006 ( .A1(n11815), .A2(n11814), .A3(n11813), .A4(n11812), .ZN(
        n11816) );
  OR2_X1 U15007 ( .A1(n11817), .A2(n11816), .ZN(n11820) );
  INV_X1 U15008 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n11818) );
  OAI22_X1 U15009 ( .A1(n11905), .A2(n11818), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15903), .ZN(n11819) );
  AOI21_X1 U15010 ( .B1(n11851), .B2(n11820), .A(n11819), .ZN(n11821) );
  AOI21_X1 U15011 ( .B1(n15912), .B2(n13621), .A(n11821), .ZN(n14479) );
  OR2_X1 U15012 ( .A1(n11823), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11824) );
  NAND2_X1 U15013 ( .A1(n11858), .A2(n11824), .ZN(n15901) );
  AOI22_X1 U15014 ( .A1(n9632), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U15015 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11278), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11827) );
  AOI22_X1 U15016 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11826) );
  NAND4_X1 U15017 ( .A1(n11829), .A2(n11828), .A3(n11827), .A4(n11826), .ZN(
        n11835) );
  AOI22_X1 U15018 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9637), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U15019 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11832) );
  AOI22_X1 U15020 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11831) );
  AOI22_X1 U15021 ( .A1(n11994), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11830) );
  NAND4_X1 U15022 ( .A1(n11833), .A2(n11832), .A3(n11831), .A4(n11830), .ZN(
        n11834) );
  NOR2_X1 U15023 ( .A1(n11835), .A2(n11834), .ZN(n11838) );
  OAI21_X1 U15024 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20640), .A(
        n20417), .ZN(n11837) );
  NAND2_X1 U15025 ( .A1(n12042), .A2(P1_EAX_REG_21__SCAN_IN), .ZN(n11836) );
  OAI211_X1 U15026 ( .C1(n12011), .C2(n11838), .A(n11837), .B(n11836), .ZN(
        n11839) );
  OAI21_X1 U15027 ( .B1(n15901), .B2(n12014), .A(n11839), .ZN(n14668) );
  INV_X1 U15028 ( .A(n14668), .ZN(n11840) );
  XNOR2_X1 U15029 ( .A(n11858), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15882) );
  NAND2_X1 U15030 ( .A1(n15882), .A2(n13621), .ZN(n11857) );
  AOI22_X1 U15031 ( .A1(n11994), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U15032 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11843) );
  AOI22_X1 U15033 ( .A1(n11441), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11842) );
  AOI22_X1 U15034 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11841) );
  NAND4_X1 U15035 ( .A1(n11844), .A2(n11843), .A3(n11842), .A4(n11841), .ZN(
        n11853) );
  AOI22_X1 U15036 ( .A1(n12025), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U15037 ( .A1(n11960), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12028), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11849) );
  NAND2_X1 U15038 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11846) );
  NAND2_X1 U15039 ( .A1(n9639), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11845) );
  AND3_X1 U15040 ( .A1(n11846), .A2(n11845), .A3(n12014), .ZN(n11848) );
  AOI22_X1 U15041 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11847) );
  NAND4_X1 U15042 ( .A1(n11850), .A2(n11849), .A3(n11848), .A4(n11847), .ZN(
        n11852) );
  OAI21_X1 U15043 ( .B1(n11853), .B2(n11852), .A(n11851), .ZN(n11855) );
  AOI22_X1 U15044 ( .A1(n12042), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20417), .ZN(n11854) );
  NAND2_X1 U15045 ( .A1(n11855), .A2(n11854), .ZN(n11856) );
  NAND2_X1 U15046 ( .A1(n11857), .A2(n11856), .ZN(n14470) );
  INV_X1 U15047 ( .A(n11858), .ZN(n11859) );
  INV_X1 U15048 ( .A(n11860), .ZN(n11862) );
  INV_X1 U15049 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11861) );
  NAND2_X1 U15050 ( .A1(n11862), .A2(n11861), .ZN(n11863) );
  NAND2_X1 U15051 ( .A1(n11909), .A2(n11863), .ZN(n14645) );
  AOI22_X1 U15052 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11867) );
  AOI22_X1 U15053 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11866) );
  AOI22_X1 U15054 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11865) );
  AOI22_X1 U15055 ( .A1(n9639), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11864) );
  NAND4_X1 U15056 ( .A1(n11867), .A2(n11866), .A3(n11865), .A4(n11864), .ZN(
        n11873) );
  AOI22_X1 U15057 ( .A1(n11960), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11994), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U15058 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U15059 ( .A1(n12020), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11869) );
  AOI22_X1 U15060 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11868) );
  NAND4_X1 U15061 ( .A1(n11871), .A2(n11870), .A3(n11869), .A4(n11868), .ZN(
        n11872) );
  NOR2_X1 U15062 ( .A1(n11873), .A2(n11872), .ZN(n11890) );
  AOI22_X1 U15063 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U15064 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11876) );
  AOI22_X1 U15065 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U15066 ( .A1(n11688), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11874) );
  NAND4_X1 U15067 ( .A1(n11877), .A2(n11876), .A3(n11875), .A4(n11874), .ZN(
        n11883) );
  AOI22_X1 U15068 ( .A1(n12025), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9632), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11881) );
  AOI22_X1 U15069 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9637), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U15070 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9644), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11879) );
  AOI22_X1 U15071 ( .A1(n12020), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11878) );
  NAND4_X1 U15072 ( .A1(n11881), .A2(n11880), .A3(n11879), .A4(n11878), .ZN(
        n11882) );
  NOR2_X1 U15073 ( .A1(n11883), .A2(n11882), .ZN(n11891) );
  XNOR2_X1 U15074 ( .A(n11890), .B(n11891), .ZN(n11887) );
  NAND2_X1 U15075 ( .A1(n12008), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11884) );
  NAND2_X1 U15076 ( .A1(n12014), .A2(n11884), .ZN(n11885) );
  AOI21_X1 U15077 ( .B1(n12042), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11885), .ZN(
        n11886) );
  OAI21_X1 U15078 ( .B1(n12011), .B2(n11887), .A(n11886), .ZN(n11888) );
  NAND2_X1 U15079 ( .A1(n11889), .A2(n11888), .ZN(n14431) );
  XNOR2_X1 U15080 ( .A(n11909), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14641) );
  NOR2_X1 U15081 ( .A1(n11891), .A2(n11890), .ZN(n11915) );
  AOI22_X1 U15082 ( .A1(n9637), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11994), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U15083 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9644), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11894) );
  AOI22_X1 U15084 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U15085 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11892) );
  NAND4_X1 U15086 ( .A1(n11895), .A2(n11894), .A3(n11893), .A4(n11892), .ZN(
        n11901) );
  AOI22_X1 U15087 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11899) );
  AOI22_X1 U15088 ( .A1(n11977), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11898) );
  AOI22_X1 U15089 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11897) );
  AOI22_X1 U15090 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11896) );
  NAND4_X1 U15091 ( .A1(n11899), .A2(n11898), .A3(n11897), .A4(n11896), .ZN(
        n11900) );
  OR2_X1 U15092 ( .A1(n11901), .A2(n11900), .ZN(n11914) );
  INV_X1 U15093 ( .A(n11914), .ZN(n11902) );
  XNOR2_X1 U15094 ( .A(n11915), .B(n11902), .ZN(n11907) );
  INV_X1 U15095 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n11904) );
  NAND2_X1 U15096 ( .A1(n12008), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11903) );
  OAI211_X1 U15097 ( .C1(n11905), .C2(n11904), .A(n12014), .B(n11903), .ZN(
        n11906) );
  AOI21_X1 U15098 ( .B1(n11907), .B2(n12037), .A(n11906), .ZN(n11908) );
  AOI21_X1 U15099 ( .B1(n14641), .B2(n13621), .A(n11908), .ZN(n14417) );
  INV_X1 U15100 ( .A(n11909), .ZN(n11910) );
  INV_X1 U15101 ( .A(n11911), .ZN(n11912) );
  INV_X1 U15102 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11927) );
  NAND2_X1 U15103 ( .A1(n11912), .A2(n11927), .ZN(n11913) );
  NAND2_X1 U15104 ( .A1(n11951), .A2(n11913), .ZN(n14630) );
  NAND2_X1 U15105 ( .A1(n11915), .A2(n11914), .ZN(n11933) );
  AOI22_X1 U15106 ( .A1(n9640), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11919) );
  AOI22_X1 U15107 ( .A1(n9637), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11918) );
  AOI22_X1 U15108 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12028), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11917) );
  AOI22_X1 U15109 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11916) );
  NAND4_X1 U15110 ( .A1(n11919), .A2(n11918), .A3(n11917), .A4(n11916), .ZN(
        n11926) );
  AOI22_X1 U15111 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U15112 ( .A1(n12020), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11920), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11923) );
  AOI22_X1 U15113 ( .A1(n11994), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11922) );
  AOI22_X1 U15114 ( .A1(n12018), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11921) );
  NAND4_X1 U15115 ( .A1(n11924), .A2(n11923), .A3(n11922), .A4(n11921), .ZN(
        n11925) );
  NOR2_X1 U15116 ( .A1(n11926), .A2(n11925), .ZN(n11934) );
  XNOR2_X1 U15117 ( .A(n11933), .B(n11934), .ZN(n11930) );
  AOI21_X1 U15118 ( .B1(n11927), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11928) );
  AOI21_X1 U15119 ( .B1(n12042), .B2(P1_EAX_REG_25__SCAN_IN), .A(n11928), .ZN(
        n11929) );
  OAI21_X1 U15120 ( .B1(n11930), .B2(n12011), .A(n11929), .ZN(n11931) );
  NAND2_X1 U15121 ( .A1(n11932), .A2(n11931), .ZN(n14407) );
  XNOR2_X1 U15122 ( .A(n11951), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14619) );
  NAND2_X1 U15123 ( .A1(n14619), .A2(n13621), .ZN(n11949) );
  NOR2_X1 U15124 ( .A1(n11934), .A2(n11933), .ZN(n11955) );
  AOI22_X1 U15125 ( .A1(n9637), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11994), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11938) );
  AOI22_X1 U15126 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9644), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11937) );
  AOI22_X1 U15127 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11936) );
  AOI22_X1 U15128 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11273), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11935) );
  NAND4_X1 U15129 ( .A1(n11938), .A2(n11937), .A3(n11936), .A4(n11935), .ZN(
        n11944) );
  AOI22_X1 U15130 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11942) );
  AOI22_X1 U15131 ( .A1(n11977), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11266), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11941) );
  AOI22_X1 U15132 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11940) );
  AOI22_X1 U15133 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11939) );
  NAND4_X1 U15134 ( .A1(n11942), .A2(n11941), .A3(n11940), .A4(n11939), .ZN(
        n11943) );
  OR2_X1 U15135 ( .A1(n11944), .A2(n11943), .ZN(n11954) );
  XNOR2_X1 U15136 ( .A(n11955), .B(n11954), .ZN(n11947) );
  INV_X1 U15137 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14621) );
  AOI21_X1 U15138 ( .B1(n14621), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11945) );
  AOI21_X1 U15139 ( .B1(n12042), .B2(P1_EAX_REG_26__SCAN_IN), .A(n11945), .ZN(
        n11946) );
  OAI21_X1 U15140 ( .B1(n11947), .B2(n12011), .A(n11946), .ZN(n11948) );
  NAND2_X1 U15141 ( .A1(n11949), .A2(n11948), .ZN(n14391) );
  NAND2_X1 U15142 ( .A1(n11952), .A2(n14380), .ZN(n11953) );
  NAND2_X1 U15143 ( .A1(n11989), .A2(n11953), .ZN(n14612) );
  NAND2_X1 U15144 ( .A1(n11955), .A2(n11954), .ZN(n11984) );
  AOI22_X1 U15145 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11994), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11959) );
  AOI22_X1 U15146 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n9592), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U15147 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U15148 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11956) );
  NAND4_X1 U15149 ( .A1(n11959), .A2(n11958), .A3(n11957), .A4(n11956), .ZN(
        n11966) );
  AOI22_X1 U15150 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12025), .B1(
        n9640), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11964) );
  AOI22_X1 U15151 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n9644), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11963) );
  AOI22_X1 U15152 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n9594), .B1(
        n11266), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U15153 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11961) );
  NAND4_X1 U15154 ( .A1(n11964), .A2(n11963), .A3(n11962), .A4(n11961), .ZN(
        n11965) );
  NOR2_X1 U15155 ( .A1(n11966), .A2(n11965), .ZN(n11985) );
  XNOR2_X1 U15156 ( .A(n11984), .B(n11985), .ZN(n11969) );
  AOI21_X1 U15157 ( .B1(n14380), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11967) );
  AOI21_X1 U15158 ( .B1(n12042), .B2(P1_EAX_REG_27__SCAN_IN), .A(n11967), .ZN(
        n11968) );
  OAI21_X1 U15159 ( .B1(n11969), .B2(n12011), .A(n11968), .ZN(n11970) );
  OAI21_X1 U15160 ( .B1(n14612), .B2(n12014), .A(n11970), .ZN(n14375) );
  INV_X1 U15161 ( .A(n11989), .ZN(n11971) );
  XOR2_X1 U15162 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B(n11971), .Z(
        n14605) );
  INV_X1 U15163 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14602) );
  NOR2_X1 U15164 ( .A1(n14602), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11972) );
  AOI211_X1 U15165 ( .C1(n12042), .C2(P1_EAX_REG_28__SCAN_IN), .A(n13621), .B(
        n11972), .ZN(n11988) );
  AOI22_X1 U15166 ( .A1(n9637), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11994), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U15167 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9644), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11975) );
  AOI22_X1 U15168 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U15169 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11273), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11973) );
  NAND4_X1 U15170 ( .A1(n11976), .A2(n11975), .A3(n11974), .A4(n11973), .ZN(
        n11983) );
  AOI22_X1 U15171 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11981) );
  AOI22_X1 U15172 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11266), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11980) );
  AOI22_X1 U15173 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12020), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11979) );
  AOI22_X1 U15174 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11441), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11978) );
  NAND4_X1 U15175 ( .A1(n11981), .A2(n11980), .A3(n11979), .A4(n11978), .ZN(
        n11982) );
  OR2_X1 U15176 ( .A1(n11983), .A2(n11982), .ZN(n12006) );
  NOR2_X1 U15177 ( .A1(n11985), .A2(n11984), .ZN(n12007) );
  XOR2_X1 U15178 ( .A(n12006), .B(n12007), .Z(n11986) );
  NAND2_X1 U15179 ( .A1(n11986), .A2(n12037), .ZN(n11987) );
  AOI22_X1 U15180 ( .A1(n14605), .A2(n13621), .B1(n11988), .B2(n11987), .ZN(
        n14360) );
  INV_X1 U15181 ( .A(n11990), .ZN(n11992) );
  INV_X1 U15182 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11991) );
  NAND2_X1 U15183 ( .A1(n11992), .A2(n11991), .ZN(n11993) );
  NAND2_X1 U15184 ( .A1(n13624), .A2(n11993), .ZN(n14589) );
  AOI22_X1 U15185 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11994), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U15186 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11998) );
  AOI22_X1 U15187 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11266), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11997) );
  AOI22_X1 U15188 ( .A1(n12020), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11996) );
  NAND4_X1 U15189 ( .A1(n11999), .A2(n11998), .A3(n11997), .A4(n11996), .ZN(
        n12005) );
  AOI22_X1 U15190 ( .A1(n12025), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9639), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12003) );
  AOI22_X1 U15191 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9636), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U15192 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U15193 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11273), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12000) );
  NAND4_X1 U15194 ( .A1(n12003), .A2(n12002), .A3(n12001), .A4(n12000), .ZN(
        n12004) );
  NOR2_X1 U15195 ( .A1(n12005), .A2(n12004), .ZN(n12017) );
  NAND2_X1 U15196 ( .A1(n12007), .A2(n12006), .ZN(n12016) );
  XNOR2_X1 U15197 ( .A(n12017), .B(n12016), .ZN(n12012) );
  AOI21_X1 U15198 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n12008), .A(
        n13621), .ZN(n12010) );
  NAND2_X1 U15199 ( .A1(n12042), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12009) );
  OAI211_X1 U15200 ( .C1(n12012), .C2(n12011), .A(n12010), .B(n12009), .ZN(
        n12013) );
  OAI21_X1 U15201 ( .B1(n14589), .B2(n12014), .A(n12013), .ZN(n14351) );
  XNOR2_X1 U15202 ( .A(n13624), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14582) );
  INV_X1 U15203 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14584) );
  NOR2_X1 U15204 ( .A1(n14584), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12015) );
  AOI211_X1 U15205 ( .C1(n12042), .C2(P1_EAX_REG_30__SCAN_IN), .A(n12015), .B(
        n13621), .ZN(n12040) );
  NOR2_X1 U15206 ( .A1(n12017), .A2(n12016), .ZN(n12036) );
  AOI22_X1 U15207 ( .A1(n11977), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12024) );
  AOI22_X1 U15208 ( .A1(n11994), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9643), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12023) );
  AOI22_X1 U15209 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12019), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12022) );
  AOI22_X1 U15210 ( .A1(n12020), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12021) );
  NAND4_X1 U15211 ( .A1(n12024), .A2(n12023), .A3(n12022), .A4(n12021), .ZN(
        n12034) );
  AOI22_X1 U15212 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U15213 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11960), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12031) );
  AOI22_X1 U15214 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11266), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12030) );
  AOI22_X1 U15215 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12029) );
  NAND4_X1 U15216 ( .A1(n12032), .A2(n12031), .A3(n12030), .A4(n12029), .ZN(
        n12033) );
  NOR2_X1 U15217 ( .A1(n12034), .A2(n12033), .ZN(n12035) );
  XNOR2_X1 U15218 ( .A(n12036), .B(n12035), .ZN(n12038) );
  NAND2_X1 U15219 ( .A1(n12038), .A2(n12037), .ZN(n12039) );
  AOI22_X1 U15220 ( .A1(n14582), .A2(n13621), .B1(n12040), .B2(n12039), .ZN(
        n14320) );
  AOI22_X1 U15221 ( .A1(n12042), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n12041), .ZN(n12043) );
  INV_X1 U15222 ( .A(n12043), .ZN(n12044) );
  XNOR2_X2 U15223 ( .A(n9672), .B(n12044), .ZN(n14331) );
  AND2_X1 U15224 ( .A1(n20040), .A2(n12911), .ZN(n12046) );
  NAND4_X1 U15225 ( .A1(n12047), .A2(n12046), .A3(n9769), .A4(n12045), .ZN(
        n13275) );
  XNOR2_X1 U15226 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12064) );
  NAND2_X1 U15227 ( .A1(n20415), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12073) );
  NAND2_X1 U15228 ( .A1(n12064), .A2(n12063), .ZN(n12050) );
  NAND2_X1 U15229 ( .A1(n20493), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12049) );
  NAND2_X1 U15230 ( .A1(n12050), .A2(n12049), .ZN(n12060) );
  XNOR2_X1 U15231 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12059) );
  NAND2_X1 U15232 ( .A1(n12060), .A2(n12059), .ZN(n12052) );
  NAND2_X1 U15233 ( .A1(n20274), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12051) );
  NAND2_X1 U15234 ( .A1(n12052), .A2(n12051), .ZN(n12062) );
  MUX2_X1 U15235 ( .A(n20655), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12061) );
  NAND2_X1 U15236 ( .A1(n12062), .A2(n12061), .ZN(n12054) );
  NAND2_X1 U15237 ( .A1(n20655), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12053) );
  NAND2_X1 U15238 ( .A1(n12054), .A2(n12053), .ZN(n12058) );
  NOR2_X1 U15239 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16158), .ZN(
        n12055) );
  NOR3_X1 U15240 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20019), .A3(
        n12058), .ZN(n12095) );
  XNOR2_X1 U15241 ( .A(n12060), .B(n12059), .ZN(n12104) );
  XNOR2_X1 U15242 ( .A(n12062), .B(n12061), .ZN(n12099) );
  XNOR2_X1 U15243 ( .A(n12064), .B(n12063), .ZN(n12082) );
  NOR4_X1 U15244 ( .A1(n12095), .A2(n12104), .A3(n12099), .A4(n12082), .ZN(
        n12065) );
  NOR2_X1 U15245 ( .A1(n12072), .A2(n12065), .ZN(n13167) );
  NAND2_X1 U15246 ( .A1(n13167), .A2(n20669), .ZN(n12906) );
  OAI21_X1 U15247 ( .B1(n13163), .B2(n13275), .A(n13546), .ZN(n12066) );
  NAND2_X1 U15248 ( .A1(n12066), .A2(n14301), .ZN(n12115) );
  NAND2_X1 U15249 ( .A1(n14302), .A2(n20024), .ZN(n12067) );
  INV_X1 U15250 ( .A(n13166), .ZN(n12901) );
  NAND2_X1 U15251 ( .A1(n12901), .A2(n13627), .ZN(n13561) );
  INV_X1 U15252 ( .A(n20669), .ZN(n20567) );
  NOR2_X1 U15253 ( .A1(n12068), .A2(n20567), .ZN(n13549) );
  NAND2_X1 U15254 ( .A1(n13549), .A2(n13630), .ZN(n12069) );
  NAND2_X1 U15255 ( .A1(n13561), .A2(n12069), .ZN(n13554) );
  NAND2_X1 U15256 ( .A1(n12070), .A2(n11367), .ZN(n12817) );
  NAND2_X1 U15257 ( .A1(n12100), .A2(n12072), .ZN(n12113) );
  NAND2_X1 U15258 ( .A1(n12072), .A2(n12092), .ZN(n12111) );
  NOR2_X1 U15259 ( .A1(n20024), .A2(n11368), .ZN(n12074) );
  OAI21_X1 U15260 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20415), .A(
        n12073), .ZN(n12075) );
  AOI21_X1 U15261 ( .B1(n20048), .B2(n11372), .A(n11367), .ZN(n12091) );
  NOR3_X1 U15262 ( .A1(n12074), .A2(n12075), .A3(n12091), .ZN(n12078) );
  INV_X1 U15263 ( .A(n12075), .ZN(n12076) );
  AOI21_X1 U15264 ( .B1(n12076), .B2(n12092), .A(n12100), .ZN(n12077) );
  INV_X1 U15265 ( .A(n12085), .ZN(n12090) );
  INV_X1 U15266 ( .A(n12817), .ZN(n12865) );
  INV_X1 U15267 ( .A(n12092), .ZN(n12081) );
  INV_X1 U15268 ( .A(n12082), .ZN(n12079) );
  AOI21_X1 U15269 ( .B1(n12865), .B2(n12081), .A(n12079), .ZN(n12086) );
  INV_X1 U15270 ( .A(n12086), .ZN(n12089) );
  INV_X1 U15271 ( .A(n12091), .ZN(n12080) );
  NOR3_X1 U15272 ( .A1(n12081), .A2(n12080), .A3(n12104), .ZN(n12088) );
  NOR2_X1 U15273 ( .A1(n20556), .A2(n12070), .ZN(n12096) );
  AOI21_X1 U15274 ( .B1(n12092), .B2(n11367), .A(n12096), .ZN(n12084) );
  NAND2_X1 U15275 ( .A1(n12105), .A2(n12082), .ZN(n12083) );
  AOI22_X1 U15276 ( .A1(n12086), .A2(n12085), .B1(n12084), .B2(n12083), .ZN(
        n12087) );
  INV_X1 U15277 ( .A(n12104), .ZN(n12093) );
  AOI21_X1 U15278 ( .B1(n12093), .B2(n12092), .A(n12091), .ZN(n12094) );
  NOR3_X1 U15279 ( .A1(n12102), .A2(n12094), .A3(n12099), .ZN(n12098) );
  INV_X1 U15280 ( .A(n12095), .ZN(n12101) );
  NOR3_X1 U15281 ( .A1(n11366), .A2(n12096), .A3(n12101), .ZN(n12097) );
  AOI211_X1 U15282 ( .C1(n12100), .C2(n12099), .A(n12098), .B(n12097), .ZN(
        n12108) );
  NOR2_X1 U15283 ( .A1(n12105), .A2(n12101), .ZN(n12107) );
  INV_X1 U15284 ( .A(n12102), .ZN(n12103) );
  NAND3_X1 U15285 ( .A1(n12105), .A2(n12104), .A3(n12103), .ZN(n12106) );
  OAI21_X1 U15286 ( .B1(n12108), .B2(n12107), .A(n12106), .ZN(n12109) );
  AOI21_X1 U15287 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20556), .A(
        n12109), .ZN(n12110) );
  NAND2_X1 U15288 ( .A1(n12111), .A2(n12110), .ZN(n12112) );
  NAND2_X1 U15289 ( .A1(n13554), .A2(n13264), .ZN(n12114) );
  AND2_X1 U15290 ( .A1(n14571), .A2(n9769), .ZN(n12116) );
  NOR4_X1 U15291 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12120) );
  NOR4_X1 U15292 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12119) );
  NOR4_X1 U15293 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12118) );
  NOR4_X1 U15294 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12117) );
  AND4_X1 U15295 ( .A1(n12120), .A2(n12119), .A3(n12118), .A4(n12117), .ZN(
        n12126) );
  NOR4_X1 U15296 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12124) );
  NOR4_X1 U15297 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12123) );
  NOR4_X1 U15298 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12122) );
  INV_X1 U15299 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n12121) );
  AND4_X1 U15300 ( .A1(n12124), .A2(n12123), .A3(n12122), .A4(n12121), .ZN(
        n12125) );
  NAND2_X1 U15301 ( .A1(n12126), .A2(n12125), .ZN(n12127) );
  NOR3_X1 U15302 ( .A1(n16008), .A2(n20020), .A3(n12909), .ZN(n12128) );
  AOI22_X1 U15303 ( .A1(n16011), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n16008), .ZN(n12129) );
  INV_X1 U15304 ( .A(n12129), .ZN(n12132) );
  AND2_X1 U15305 ( .A1(n13033), .A2(n20020), .ZN(n12130) );
  INV_X1 U15306 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16385) );
  NOR2_X1 U15307 ( .A1(n16015), .A2(n16385), .ZN(n12131) );
  NOR2_X1 U15308 ( .A1(n12132), .A2(n12131), .ZN(n12133) );
  NAND2_X1 U15309 ( .A1(n10550), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12135) );
  NOR2_X1 U15310 ( .A1(n19714), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12136) );
  AOI21_X1 U15311 ( .B1(n12161), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n12136), .ZN(n12137) );
  NAND2_X1 U15312 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12143) );
  NAND2_X1 U15313 ( .A1(n12161), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12139) );
  NAND2_X1 U15314 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19438) );
  NAND2_X1 U15315 ( .A1(n19735), .A2(n20827), .ZN(n19348) );
  AND2_X1 U15316 ( .A1(n19438), .A2(n19348), .ZN(n19289) );
  NAND2_X1 U15317 ( .A1(n19289), .A2(n19520), .ZN(n19411) );
  NAND2_X1 U15318 ( .A1(n12139), .A2(n19411), .ZN(n12140) );
  INV_X1 U15319 ( .A(n12143), .ZN(n12144) );
  NAND2_X1 U15320 ( .A1(n12146), .A2(n12156), .ZN(n12150) );
  NAND2_X1 U15321 ( .A1(n19438), .A2(n19725), .ZN(n12147) );
  NOR2_X1 U15322 ( .A1(n19725), .A2(n19735), .ZN(n19562) );
  AND2_X1 U15323 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19562), .ZN(
        n12158) );
  INV_X1 U15324 ( .A(n12158), .ZN(n12159) );
  NAND2_X1 U15325 ( .A1(n12147), .A2(n12159), .ZN(n13840) );
  NOR2_X1 U15326 ( .A1(n13840), .A2(n19714), .ZN(n12148) );
  AOI21_X1 U15327 ( .B1(n12161), .B2(n10596), .A(n12148), .ZN(n12149) );
  NAND2_X1 U15328 ( .A1(n13257), .A2(n13258), .ZN(n12155) );
  INV_X1 U15329 ( .A(n12152), .ZN(n12153) );
  NAND2_X1 U15330 ( .A1(n12151), .A2(n12153), .ZN(n12154) );
  NAND2_X1 U15331 ( .A1(n12157), .A2(n12156), .ZN(n12163) );
  NAND2_X1 U15332 ( .A1(n12158), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19570) );
  NAND2_X1 U15333 ( .A1(n19718), .A2(n12159), .ZN(n12160) );
  AND3_X1 U15334 ( .A1(n19570), .A2(n19520), .A3(n12160), .ZN(n13853) );
  AOI21_X1 U15335 ( .B1(n12161), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13853), .ZN(n12162) );
  NAND2_X1 U15336 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12165) );
  NAND2_X1 U15337 ( .A1(n13410), .A2(n13411), .ZN(n12168) );
  INV_X1 U15338 ( .A(n12165), .ZN(n12166) );
  AOI22_X1 U15339 ( .A1(n12164), .A2(n12166), .B1(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n10550), .ZN(n12167) );
  INV_X1 U15340 ( .A(n12517), .ZN(n12564) );
  INV_X1 U15341 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19121) );
  NOR2_X1 U15342 ( .A1(n12564), .A2(n19121), .ZN(n13242) );
  AOI22_X1 U15343 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12460), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12177) );
  AOI22_X1 U15344 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12174) );
  NAND2_X1 U15345 ( .A1(n12380), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12173) );
  NAND2_X1 U15346 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12172) );
  INV_X1 U15347 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12169) );
  OAI22_X1 U15348 ( .A1(n12343), .A2(n12169), .B1(n19097), .B2(n9669), .ZN(
        n12170) );
  AOI21_X1 U15349 ( .B1(n12452), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n12170), .ZN(n12171) );
  AND4_X1 U15350 ( .A1(n12174), .A2(n12173), .A3(n12172), .A4(n12171), .ZN(
        n12176) );
  AOI22_X1 U15351 ( .A1(n10777), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13712), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12175) );
  NAND3_X1 U15352 ( .A1(n12177), .A2(n12176), .A3(n12175), .ZN(n12183) );
  AOI22_X1 U15353 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12181) );
  NAND2_X1 U15354 ( .A1(n12464), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12180) );
  NAND2_X1 U15355 ( .A1(n10714), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12179) );
  NAND2_X1 U15356 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12178) );
  NAND4_X1 U15357 ( .A1(n12181), .A2(n12180), .A3(n12179), .A4(n12178), .ZN(
        n12182) );
  NAND2_X1 U15358 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12187) );
  NAND2_X1 U15359 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12186) );
  NAND2_X1 U15360 ( .A1(n10777), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12185) );
  NAND2_X1 U15361 ( .A1(n13712), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12184) );
  NAND4_X1 U15362 ( .A1(n12187), .A2(n12186), .A3(n12185), .A4(n12184), .ZN(
        n12196) );
  AOI22_X1 U15363 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12451), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12194) );
  NAND2_X1 U15364 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12193) );
  NAND2_X1 U15365 ( .A1(n12380), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12192) );
  NAND2_X1 U15366 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12340), .ZN(
        n12188) );
  OAI21_X1 U15367 ( .B1(n12343), .B2(n12189), .A(n12188), .ZN(n12190) );
  AOI21_X1 U15368 ( .B1(n12452), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n12190), .ZN(n12191) );
  NAND4_X1 U15369 ( .A1(n12194), .A2(n12193), .A3(n12192), .A4(n12191), .ZN(
        n12195) );
  NOR2_X1 U15370 ( .A1(n12196), .A2(n12195), .ZN(n12204) );
  INV_X1 U15371 ( .A(n12464), .ZN(n12398) );
  OAI22_X1 U15372 ( .A1(n12198), .A2(n12398), .B1(n10899), .B2(n12197), .ZN(
        n12202) );
  INV_X1 U15373 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n19471) );
  NAND2_X1 U15374 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12200) );
  NAND2_X1 U15375 ( .A1(n10673), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12199) );
  OAI211_X1 U15376 ( .C1(n12412), .C2(n19471), .A(n12200), .B(n12199), .ZN(
        n12201) );
  NOR2_X1 U15377 ( .A1(n12202), .A2(n12201), .ZN(n12203) );
  NAND2_X1 U15378 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12208) );
  NAND2_X1 U15379 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12207) );
  NAND2_X1 U15380 ( .A1(n10777), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n12206) );
  NAND2_X1 U15381 ( .A1(n13712), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12205) );
  NAND4_X1 U15382 ( .A1(n12208), .A2(n12207), .A3(n12206), .A4(n12205), .ZN(
        n12216) );
  AOI22_X1 U15383 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12451), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12214) );
  NAND2_X1 U15384 ( .A1(n12380), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12213) );
  NAND2_X1 U15385 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n12212) );
  INV_X1 U15386 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12209) );
  OAI22_X1 U15387 ( .A1(n12343), .A2(n12209), .B1(n10706), .B2(n9669), .ZN(
        n12210) );
  AOI21_X1 U15388 ( .B1(n12452), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n12210), .ZN(n12211) );
  NAND4_X1 U15389 ( .A1(n12214), .A2(n12213), .A3(n12212), .A4(n12211), .ZN(
        n12215) );
  NOR2_X1 U15390 ( .A1(n12216), .A2(n12215), .ZN(n12222) );
  AOI22_X1 U15391 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__2__SCAN_IN), .B2(n10673), .ZN(n12220) );
  NAND2_X1 U15392 ( .A1(n12464), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12219) );
  NAND2_X1 U15393 ( .A1(n10714), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12218) );
  NAND2_X1 U15394 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n12217) );
  NAND2_X1 U15395 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12227) );
  NAND2_X1 U15396 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12226) );
  NAND2_X1 U15397 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12225) );
  NAND2_X1 U15398 ( .A1(n13712), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12224) );
  NAND4_X1 U15399 ( .A1(n12227), .A2(n12226), .A3(n12225), .A4(n12224), .ZN(
        n12236) );
  AOI22_X1 U15400 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12451), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12234) );
  NAND2_X1 U15401 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12233) );
  NAND2_X1 U15402 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12232) );
  NAND2_X1 U15403 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12340), .ZN(
        n12228) );
  OAI21_X1 U15404 ( .B1(n12343), .B2(n12229), .A(n12228), .ZN(n12230) );
  AOI21_X1 U15405 ( .B1(n12452), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n12230), .ZN(n12231) );
  NAND4_X1 U15406 ( .A1(n12234), .A2(n12233), .A3(n12232), .A4(n12231), .ZN(
        n12235) );
  NOR2_X1 U15407 ( .A1(n12236), .A2(n12235), .ZN(n12244) );
  NAND2_X1 U15408 ( .A1(n12380), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12238) );
  NAND2_X1 U15409 ( .A1(n10673), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n12237) );
  OAI211_X1 U15410 ( .C1(n10899), .C2(n12239), .A(n12238), .B(n12237), .ZN(
        n12242) );
  OAI22_X1 U15411 ( .A1(n12398), .A2(n12240), .B1(n12424), .B2(n12533), .ZN(
        n12241) );
  NOR2_X1 U15412 ( .A1(n12242), .A2(n12241), .ZN(n12243) );
  AOI22_X1 U15413 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12460), .B1(
        n12377), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15414 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12379), .B1(
        n12380), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12251) );
  NAND2_X1 U15415 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12248) );
  NAND2_X1 U15416 ( .A1(n12452), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12247) );
  NAND2_X1 U15417 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12246) );
  AOI22_X1 U15418 ( .A1(n12453), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n12340), .ZN(n12245) );
  AND4_X1 U15419 ( .A1(n12248), .A2(n12247), .A3(n12246), .A4(n12245), .ZN(
        n12250) );
  AOI22_X1 U15420 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10777), .B1(
        n13712), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12249) );
  NAND4_X1 U15421 ( .A1(n12252), .A2(n12251), .A3(n12250), .A4(n12249), .ZN(
        n12258) );
  AOI22_X1 U15422 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__4__SCAN_IN), .B2(n10673), .ZN(n12256) );
  INV_X1 U15423 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n20792) );
  NAND2_X1 U15424 ( .A1(n12464), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12255) );
  NAND2_X1 U15425 ( .A1(n10714), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12254) );
  NAND2_X1 U15426 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12253) );
  NAND4_X1 U15427 ( .A1(n12256), .A2(n12255), .A3(n12254), .A4(n12253), .ZN(
        n12257) );
  NAND2_X1 U15428 ( .A1(n13665), .A2(n13666), .ZN(n13898) );
  AOI22_X1 U15429 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12380), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12266) );
  AOI22_X1 U15430 ( .A1(n12464), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13712), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15431 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10777), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12264) );
  NAND2_X1 U15432 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12262) );
  NAND2_X1 U15433 ( .A1(n10673), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n12261) );
  AOI22_X1 U15434 ( .A1(n12453), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12260) );
  NAND2_X1 U15435 ( .A1(n12452), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12259) );
  AND4_X1 U15436 ( .A1(n12262), .A2(n12261), .A3(n12260), .A4(n12259), .ZN(
        n12263) );
  NAND4_X1 U15437 ( .A1(n12266), .A2(n12265), .A3(n12264), .A4(n12263), .ZN(
        n12272) );
  AOI22_X1 U15438 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12270) );
  NAND2_X1 U15439 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12269) );
  NAND2_X1 U15440 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n12268) );
  NAND2_X1 U15441 ( .A1(n10714), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12267) );
  NAND4_X1 U15442 ( .A1(n12270), .A2(n12269), .A3(n12268), .A4(n12267), .ZN(
        n12271) );
  NOR2_X1 U15443 ( .A1(n12272), .A2(n12271), .ZN(n12753) );
  NOR2_X2 U15444 ( .A1(n13898), .A2(n12753), .ZN(n13899) );
  NAND2_X1 U15445 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12276) );
  NAND2_X1 U15446 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12275) );
  NAND2_X1 U15447 ( .A1(n10777), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12274) );
  NAND2_X1 U15448 ( .A1(n13712), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12273) );
  NAND4_X1 U15449 ( .A1(n12276), .A2(n12275), .A3(n12274), .A4(n12273), .ZN(
        n12284) );
  AOI22_X1 U15450 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12282) );
  NAND2_X1 U15451 ( .A1(n12380), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12281) );
  NAND2_X1 U15452 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12280) );
  NAND2_X1 U15453 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12340), .ZN(
        n12277) );
  OAI21_X1 U15454 ( .B1(n12343), .B2(n12595), .A(n12277), .ZN(n12278) );
  AOI21_X1 U15455 ( .B1(n12452), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n12278), .ZN(n12279) );
  NAND4_X1 U15456 ( .A1(n12282), .A2(n12281), .A3(n12280), .A4(n12279), .ZN(
        n12283) );
  NOR2_X1 U15457 ( .A1(n12284), .A2(n12283), .ZN(n12290) );
  AOI22_X1 U15458 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12288) );
  NAND2_X1 U15459 ( .A1(n12464), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12287) );
  NAND2_X1 U15460 ( .A1(n10714), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12286) );
  NAND2_X1 U15461 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12285) );
  AND4_X1 U15462 ( .A1(n12288), .A2(n12287), .A3(n12286), .A4(n12285), .ZN(
        n12289) );
  INV_X1 U15463 ( .A(n13905), .ZN(n12291) );
  AOI22_X1 U15464 ( .A1(n12380), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12299) );
  AOI22_X1 U15465 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10777), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15466 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13712), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12297) );
  NAND2_X1 U15467 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12295) );
  NAND2_X1 U15468 ( .A1(n12452), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12294) );
  NAND2_X1 U15469 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12293) );
  AOI22_X1 U15470 ( .A1(n12453), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n12340), .ZN(n12292) );
  AND4_X1 U15471 ( .A1(n12295), .A2(n12294), .A3(n12293), .A4(n12292), .ZN(
        n12296) );
  NAND4_X1 U15472 ( .A1(n12299), .A2(n12298), .A3(n12297), .A4(n12296), .ZN(
        n12305) );
  AOI22_X1 U15473 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12303) );
  NAND2_X1 U15474 ( .A1(n12464), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12302) );
  NAND2_X1 U15475 ( .A1(n10714), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12301) );
  NAND2_X1 U15476 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12300) );
  NAND4_X1 U15477 ( .A1(n12303), .A2(n12302), .A3(n12301), .A4(n12300), .ZN(
        n12304) );
  AOI22_X1 U15478 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12460), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12313) );
  AOI22_X1 U15479 ( .A1(n12380), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12312) );
  NAND2_X1 U15480 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12309) );
  NAND2_X1 U15481 ( .A1(n12452), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12308) );
  NAND2_X1 U15482 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12307) );
  AOI22_X1 U15483 ( .A1(n12453), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12306) );
  AND4_X1 U15484 ( .A1(n12309), .A2(n12308), .A3(n12307), .A4(n12306), .ZN(
        n12311) );
  AOI22_X1 U15485 ( .A1(n10777), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13712), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12310) );
  NAND4_X1 U15486 ( .A1(n12313), .A2(n12312), .A3(n12311), .A4(n12310), .ZN(
        n12319) );
  AOI22_X1 U15487 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12317) );
  NAND2_X1 U15488 ( .A1(n12464), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12316) );
  NAND2_X1 U15489 ( .A1(n10714), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12315) );
  NAND2_X1 U15490 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12314) );
  NAND4_X1 U15491 ( .A1(n12317), .A2(n12316), .A3(n12315), .A4(n12314), .ZN(
        n12318) );
  AOI22_X1 U15492 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n12377), .B1(
        n12460), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12327) );
  AOI22_X1 U15493 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12379), .B1(
        n12380), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12326) );
  NAND2_X1 U15494 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12323) );
  NAND2_X1 U15495 ( .A1(n12452), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12322) );
  NAND2_X1 U15496 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12321) );
  AOI22_X1 U15497 ( .A1(n12453), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n12340), .ZN(n12320) );
  AND4_X1 U15498 ( .A1(n12323), .A2(n12322), .A3(n12321), .A4(n12320), .ZN(
        n12325) );
  AOI22_X1 U15499 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n10777), .B1(
        n13712), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12324) );
  NAND4_X1 U15500 ( .A1(n12327), .A2(n12326), .A3(n12325), .A4(n12324), .ZN(
        n12333) );
  AOI22_X1 U15501 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n10673), .ZN(n12331) );
  NAND2_X1 U15502 ( .A1(n12464), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12330) );
  NAND2_X1 U15503 ( .A1(n10714), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12329) );
  NAND2_X1 U15504 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12328) );
  NAND4_X1 U15505 ( .A1(n12331), .A2(n12330), .A3(n12329), .A4(n12328), .ZN(
        n12332) );
  NOR2_X1 U15506 ( .A1(n12333), .A2(n12332), .ZN(n14184) );
  NAND2_X1 U15507 ( .A1(n12335), .A2(n12334), .ZN(n14181) );
  NAND2_X1 U15508 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n12339) );
  NAND2_X1 U15509 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12338) );
  NAND2_X1 U15510 ( .A1(n10777), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12337) );
  NAND2_X1 U15511 ( .A1(n13712), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12336) );
  NAND4_X1 U15512 ( .A1(n12339), .A2(n12338), .A3(n12337), .A4(n12336), .ZN(
        n12350) );
  AOI22_X1 U15513 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12451), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12348) );
  NAND2_X1 U15514 ( .A1(n12380), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12347) );
  NAND2_X1 U15515 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12346) );
  INV_X1 U15516 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12342) );
  NAND2_X1 U15517 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n12340), .ZN(
        n12341) );
  OAI21_X1 U15518 ( .B1(n12343), .B2(n12342), .A(n12341), .ZN(n12344) );
  AOI21_X1 U15519 ( .B1(n12452), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n12344), .ZN(n12345) );
  NAND4_X1 U15520 ( .A1(n12348), .A2(n12347), .A3(n12346), .A4(n12345), .ZN(
        n12349) );
  NOR2_X1 U15521 ( .A1(n12350), .A2(n12349), .ZN(n12358) );
  INV_X1 U15522 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12351) );
  OAI22_X1 U15523 ( .A1(n10706), .A2(n10899), .B1(n12398), .B2(n12351), .ZN(
        n12356) );
  INV_X1 U15524 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12354) );
  NAND2_X1 U15525 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12353) );
  NAND2_X1 U15526 ( .A1(n10673), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12352) );
  OAI211_X1 U15527 ( .C1(n12412), .C2(n12354), .A(n12353), .B(n12352), .ZN(
        n12355) );
  NOR2_X1 U15528 ( .A1(n12356), .A2(n12355), .ZN(n12357) );
  AOI22_X1 U15529 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n12377), .B1(
        n12460), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12366) );
  AOI22_X1 U15530 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12379), .B1(
        n12380), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12365) );
  NAND2_X1 U15531 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n12362) );
  NAND2_X1 U15532 ( .A1(n12452), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n12361) );
  NAND2_X1 U15533 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12360) );
  AOI22_X1 U15534 ( .A1(n12453), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n12340), .ZN(n12359) );
  AND4_X1 U15535 ( .A1(n12362), .A2(n12361), .A3(n12360), .A4(n12359), .ZN(
        n12364) );
  AOI22_X1 U15536 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n10777), .B1(
        n13712), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12363) );
  NAND4_X1 U15537 ( .A1(n12366), .A2(n12365), .A3(n12364), .A4(n12363), .ZN(
        n12372) );
  AOI22_X1 U15538 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__3__SCAN_IN), .B2(n10673), .ZN(n12370) );
  NAND2_X1 U15539 ( .A1(n12464), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12369) );
  NAND2_X1 U15540 ( .A1(n10714), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12368) );
  NAND2_X1 U15541 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n12367) );
  NAND4_X1 U15542 ( .A1(n12370), .A2(n12369), .A3(n12368), .A4(n12367), .ZN(
        n12371) );
  INV_X1 U15543 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12376) );
  INV_X1 U15544 ( .A(n12452), .ZN(n12375) );
  AOI22_X1 U15545 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12374) );
  AOI22_X1 U15546 ( .A1(n12453), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n12340), .ZN(n12373) );
  OAI211_X1 U15547 ( .C1(n12376), .C2(n12375), .A(n12374), .B(n12373), .ZN(
        n12387) );
  INV_X1 U15548 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12378) );
  INV_X1 U15549 ( .A(n12460), .ZN(n12418) );
  INV_X1 U15550 ( .A(n12377), .ZN(n12420) );
  INV_X1 U15551 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12556) );
  OAI22_X1 U15552 ( .A1(n12378), .A2(n12418), .B1(n12420), .B2(n12556), .ZN(
        n12386) );
  INV_X1 U15553 ( .A(n12379), .ZN(n12450) );
  INV_X1 U15554 ( .A(n12380), .ZN(n12449) );
  INV_X1 U15555 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12381) );
  OAI22_X1 U15556 ( .A1(n20792), .A2(n12450), .B1(n12449), .B2(n12381), .ZN(
        n12385) );
  INV_X1 U15557 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12383) );
  INV_X1 U15558 ( .A(n13712), .ZN(n12422) );
  INV_X1 U15559 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12382) );
  OAI22_X1 U15560 ( .A1(n12383), .A2(n12424), .B1(n12422), .B2(n12382), .ZN(
        n12384) );
  NOR4_X1 U15561 ( .A1(n12387), .A2(n12386), .A3(n12385), .A4(n12384), .ZN(
        n12391) );
  AOI22_X1 U15562 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10714), .B1(
        n12464), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12390) );
  AOI22_X1 U15563 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__4__SCAN_IN), .B2(n10673), .ZN(n12389) );
  NAND2_X1 U15564 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12388) );
  INV_X1 U15565 ( .A(n12392), .ZN(n12396) );
  OAI22_X1 U15566 ( .A1(n12396), .A2(n12395), .B1(n12394), .B2(n12393), .ZN(
        n12400) );
  OAI22_X1 U15567 ( .A1(n12398), .A2(n12397), .B1(n10899), .B2(n13370), .ZN(
        n12399) );
  AOI211_X1 U15568 ( .C1(n10676), .C2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n12400), .B(n12399), .ZN(n12408) );
  AOI22_X1 U15569 ( .A1(n12380), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12404) );
  AOI22_X1 U15570 ( .A1(n12453), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12403) );
  AOI22_X1 U15571 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12402) );
  NAND2_X1 U15572 ( .A1(n12452), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12401) );
  AND4_X1 U15573 ( .A1(n12404), .A2(n12403), .A3(n12402), .A4(n12401), .ZN(
        n12407) );
  AOI22_X1 U15574 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12460), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12406) );
  AOI22_X1 U15575 ( .A1(n10777), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13712), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12405) );
  NAND4_X1 U15576 ( .A1(n12408), .A2(n12407), .A3(n12406), .A4(n12405), .ZN(
        n15109) );
  AOI22_X1 U15577 ( .A1(n12464), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10714), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12410) );
  AOI22_X1 U15578 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10673), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12409) );
  OAI211_X1 U15579 ( .C1(n12412), .C2(n12411), .A(n12410), .B(n12409), .ZN(
        n12428) );
  AOI22_X1 U15580 ( .A1(n12380), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12416) );
  AOI22_X1 U15581 ( .A1(n12453), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12415) );
  AOI22_X1 U15582 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12414) );
  NAND2_X1 U15583 ( .A1(n12452), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n12413) );
  NAND4_X1 U15584 ( .A1(n12416), .A2(n12415), .A3(n12414), .A4(n12413), .ZN(
        n12427) );
  INV_X1 U15585 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12419) );
  OAI22_X1 U15586 ( .A1(n12420), .A2(n12419), .B1(n12418), .B2(n12417), .ZN(
        n12426) );
  INV_X1 U15587 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12423) );
  OAI22_X1 U15588 ( .A1(n12424), .A2(n12423), .B1(n12422), .B2(n12421), .ZN(
        n12425) );
  NOR4_X1 U15589 ( .A1(n12428), .A2(n12427), .A3(n12426), .A4(n12425), .ZN(
        n15105) );
  INV_X1 U15590 ( .A(n12598), .ZN(n12624) );
  AOI22_X1 U15591 ( .A1(n12624), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12596), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U15592 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9588), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12437) );
  AOI22_X1 U15593 ( .A1(n12623), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12436) );
  INV_X1 U15594 ( .A(n10677), .ZN(n12594) );
  INV_X1 U15595 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12433) );
  NAND2_X1 U15596 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12432) );
  INV_X1 U15597 ( .A(n12429), .ZN(n12431) );
  NAND2_X1 U15598 ( .A1(n10596), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12430) );
  NAND2_X1 U15599 ( .A1(n12431), .A2(n12430), .ZN(n12616) );
  OAI211_X1 U15600 ( .C1(n12594), .C2(n12433), .A(n12432), .B(n12616), .ZN(
        n12434) );
  INV_X1 U15601 ( .A(n12434), .ZN(n12435) );
  NAND4_X1 U15602 ( .A1(n12438), .A2(n12437), .A3(n12436), .A4(n12435), .ZN(
        n12447) );
  AOI22_X1 U15603 ( .A1(n12624), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12596), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12445) );
  AOI22_X1 U15604 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9588), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12444) );
  AOI22_X1 U15605 ( .A1(n12623), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12443) );
  INV_X1 U15606 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12440) );
  NAND2_X1 U15607 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12439) );
  INV_X1 U15608 ( .A(n12616), .ZN(n12578) );
  OAI211_X1 U15609 ( .C1(n12594), .C2(n12440), .A(n12439), .B(n12578), .ZN(
        n12441) );
  INV_X1 U15610 ( .A(n12441), .ZN(n12442) );
  NAND4_X1 U15611 ( .A1(n12445), .A2(n12444), .A3(n12443), .A4(n12442), .ZN(
        n12446) );
  NAND2_X1 U15612 ( .A1(n12447), .A2(n12446), .ZN(n12476) );
  INV_X1 U15613 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n20770) );
  INV_X1 U15614 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12448) );
  OAI22_X1 U15615 ( .A1(n20770), .A2(n12450), .B1(n12449), .B2(n12448), .ZN(
        n12459) );
  NAND2_X1 U15616 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12457) );
  NAND2_X1 U15617 ( .A1(n12452), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12456) );
  NAND2_X1 U15618 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12455) );
  AOI22_X1 U15619 ( .A1(n12453), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n12340), .ZN(n12454) );
  NAND4_X1 U15620 ( .A1(n12457), .A2(n12456), .A3(n12455), .A4(n12454), .ZN(
        n12458) );
  NOR2_X1 U15621 ( .A1(n12459), .A2(n12458), .ZN(n12463) );
  AOI22_X1 U15622 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n12377), .B1(
        n12460), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12462) );
  AOI22_X1 U15623 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n10777), .B1(
        n13712), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12461) );
  NAND3_X1 U15624 ( .A1(n12463), .A2(n12462), .A3(n12461), .ZN(n12470) );
  AOI22_X1 U15625 ( .A1(n12392), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n10673), .ZN(n12468) );
  NAND2_X1 U15626 ( .A1(n12464), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12467) );
  NAND2_X1 U15627 ( .A1(n10714), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12466) );
  NAND2_X1 U15628 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12465) );
  NAND4_X1 U15629 ( .A1(n12468), .A2(n12467), .A3(n12466), .A4(n12465), .ZN(
        n12469) );
  NOR2_X1 U15630 ( .A1(n12470), .A2(n12469), .ZN(n12471) );
  OAI21_X1 U15631 ( .B1(n12687), .B2(n12476), .A(n12471), .ZN(n12475) );
  INV_X1 U15632 ( .A(n12471), .ZN(n12473) );
  INV_X1 U15633 ( .A(n12476), .ZN(n12472) );
  NAND2_X1 U15634 ( .A1(n12494), .A2(n10753), .ZN(n12474) );
  NAND2_X1 U15635 ( .A1(n12475), .A2(n12474), .ZN(n12498) );
  NOR2_X1 U15636 ( .A1(n10753), .A2(n12476), .ZN(n15095) );
  INV_X1 U15637 ( .A(n15104), .ZN(n12477) );
  AOI22_X1 U15638 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12623), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12484) );
  AOI22_X1 U15639 ( .A1(n12624), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12596), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12483) );
  AOI22_X1 U15640 ( .A1(n9587), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12482) );
  INV_X1 U15641 ( .A(n10663), .ZN(n12618) );
  INV_X1 U15642 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12479) );
  NAND2_X1 U15643 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12478) );
  OAI211_X1 U15644 ( .C1(n12618), .C2(n12479), .A(n12478), .B(n12578), .ZN(
        n12480) );
  INV_X1 U15645 ( .A(n12480), .ZN(n12481) );
  NAND4_X1 U15646 ( .A1(n12484), .A2(n12483), .A3(n12482), .A4(n12481), .ZN(
        n12493) );
  AOI22_X1 U15647 ( .A1(n12623), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12624), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12491) );
  AOI22_X1 U15648 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12490) );
  AOI22_X1 U15649 ( .A1(n12596), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9638), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12489) );
  NAND2_X1 U15650 ( .A1(n12587), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12485) );
  OAI211_X1 U15651 ( .C1(n12618), .C2(n12486), .A(n12485), .B(n12616), .ZN(
        n12487) );
  INV_X1 U15652 ( .A(n12487), .ZN(n12488) );
  NAND4_X1 U15653 ( .A1(n12491), .A2(n12490), .A3(n12489), .A4(n12488), .ZN(
        n12492) );
  AND2_X1 U15654 ( .A1(n12493), .A2(n12492), .ZN(n15086) );
  INV_X1 U15655 ( .A(n15086), .ZN(n12497) );
  INV_X1 U15656 ( .A(n12494), .ZN(n12495) );
  AND2_X1 U15657 ( .A1(n12494), .A2(n15086), .ZN(n12500) );
  INV_X1 U15658 ( .A(n15095), .ZN(n12496) );
  NOR3_X1 U15659 ( .A1(n12498), .A2(n12497), .A3(n12496), .ZN(n12499) );
  INV_X1 U15660 ( .A(n12500), .ZN(n12523) );
  AOI22_X1 U15661 ( .A1(n12624), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12596), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12507) );
  AOI22_X1 U15662 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12506) );
  AOI22_X1 U15663 ( .A1(n12623), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12505) );
  INV_X1 U15664 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12502) );
  NAND2_X1 U15665 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n12501) );
  OAI211_X1 U15666 ( .C1(n12594), .C2(n12502), .A(n12501), .B(n12616), .ZN(
        n12503) );
  INV_X1 U15667 ( .A(n12503), .ZN(n12504) );
  NAND4_X1 U15668 ( .A1(n12507), .A2(n12506), .A3(n12505), .A4(n12504), .ZN(
        n12516) );
  AOI22_X1 U15669 ( .A1(n12624), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12596), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12514) );
  AOI22_X1 U15670 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9588), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12513) );
  AOI22_X1 U15671 ( .A1(n12623), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12512) );
  INV_X1 U15672 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12509) );
  NAND2_X1 U15673 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12508) );
  OAI211_X1 U15674 ( .C1(n12594), .C2(n12509), .A(n12508), .B(n12578), .ZN(
        n12510) );
  INV_X1 U15675 ( .A(n12510), .ZN(n12511) );
  NAND4_X1 U15676 ( .A1(n12514), .A2(n12513), .A3(n12512), .A4(n12511), .ZN(
        n12515) );
  AND2_X1 U15677 ( .A1(n12516), .A2(n12515), .ZN(n12521) );
  XNOR2_X1 U15678 ( .A(n12523), .B(n12521), .ZN(n12518) );
  NAND2_X1 U15679 ( .A1(n12518), .A2(n12517), .ZN(n12519) );
  NAND2_X1 U15680 ( .A1(n12687), .A2(n12521), .ZN(n15083) );
  INV_X1 U15681 ( .A(n12521), .ZN(n12522) );
  NOR2_X1 U15682 ( .A1(n12523), .A2(n12522), .ZN(n12541) );
  AOI22_X1 U15683 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12623), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12529) );
  AOI22_X1 U15684 ( .A1(n12624), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9587), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12528) );
  AOI22_X1 U15685 ( .A1(n12596), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12527) );
  INV_X1 U15686 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19114) );
  NAND2_X1 U15687 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n12524) );
  OAI211_X1 U15688 ( .C1(n12618), .C2(n19114), .A(n12524), .B(n12616), .ZN(
        n12525) );
  INV_X1 U15689 ( .A(n12525), .ZN(n12526) );
  NAND4_X1 U15690 ( .A1(n12529), .A2(n12528), .A3(n12527), .A4(n12526), .ZN(
        n12540) );
  AOI22_X1 U15691 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12624), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12538) );
  AOI22_X1 U15692 ( .A1(n10677), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9638), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12537) );
  AOI22_X1 U15693 ( .A1(n12596), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12536) );
  INV_X1 U15694 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12531) );
  OR2_X1 U15695 ( .A1(n12618), .A2(n12531), .ZN(n12532) );
  OAI211_X1 U15696 ( .C1(n12530), .C2(n12533), .A(n12578), .B(n12532), .ZN(
        n12534) );
  INV_X1 U15697 ( .A(n12534), .ZN(n12535) );
  NAND4_X1 U15698 ( .A1(n12538), .A2(n12537), .A3(n12536), .A4(n12535), .ZN(
        n12539) );
  AND2_X1 U15699 ( .A1(n12540), .A2(n12539), .ZN(n12545) );
  NAND2_X1 U15700 ( .A1(n12541), .A2(n12545), .ZN(n12565) );
  INV_X1 U15701 ( .A(n12541), .ZN(n12543) );
  INV_X1 U15702 ( .A(n12545), .ZN(n12542) );
  AOI21_X1 U15703 ( .B1(n12543), .B2(n12542), .A(n12564), .ZN(n12544) );
  NAND2_X1 U15704 ( .A1(n12687), .A2(n12545), .ZN(n15079) );
  AOI22_X1 U15705 ( .A1(n12624), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12596), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12554) );
  AOI22_X1 U15706 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12553) );
  AOI22_X1 U15707 ( .A1(n12623), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12552) );
  INV_X1 U15708 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12549) );
  NAND2_X1 U15709 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12548) );
  OAI211_X1 U15710 ( .C1(n12594), .C2(n12549), .A(n12548), .B(n12616), .ZN(
        n12550) );
  INV_X1 U15711 ( .A(n12550), .ZN(n12551) );
  NAND4_X1 U15712 ( .A1(n12554), .A2(n12553), .A3(n12552), .A4(n12551), .ZN(
        n12563) );
  AOI22_X1 U15713 ( .A1(n12624), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12596), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12561) );
  AOI22_X1 U15714 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9588), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12560) );
  AOI22_X1 U15715 ( .A1(n12623), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12559) );
  NAND2_X1 U15716 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12555) );
  OAI211_X1 U15717 ( .C1(n12594), .C2(n12556), .A(n12555), .B(n12578), .ZN(
        n12557) );
  INV_X1 U15718 ( .A(n12557), .ZN(n12558) );
  NAND4_X1 U15719 ( .A1(n12561), .A2(n12560), .A3(n12559), .A4(n12558), .ZN(
        n12562) );
  NAND2_X1 U15720 ( .A1(n12563), .A2(n12562), .ZN(n12567) );
  AOI21_X1 U15721 ( .B1(n12565), .B2(n12567), .A(n12564), .ZN(n12566) );
  OR2_X1 U15722 ( .A1(n12565), .A2(n12567), .ZN(n15057) );
  NAND2_X1 U15723 ( .A1(n12566), .A2(n15057), .ZN(n12570) );
  XNOR2_X1 U15724 ( .A(n12569), .B(n12570), .ZN(n15068) );
  INV_X1 U15725 ( .A(n12567), .ZN(n12568) );
  NAND2_X1 U15726 ( .A1(n12687), .A2(n12568), .ZN(n15070) );
  AOI22_X1 U15727 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12624), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12576) );
  AOI22_X1 U15728 ( .A1(n12623), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9587), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12575) );
  AOI22_X1 U15729 ( .A1(n12596), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12574) );
  NAND2_X1 U15730 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12571) );
  OAI211_X1 U15731 ( .C1(n12618), .C2(n13370), .A(n12571), .B(n12616), .ZN(
        n12572) );
  INV_X1 U15732 ( .A(n12572), .ZN(n12573) );
  NAND4_X1 U15733 ( .A1(n12576), .A2(n12575), .A3(n12574), .A4(n12573), .ZN(
        n12586) );
  AOI22_X1 U15734 ( .A1(n12624), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12596), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12584) );
  AOI22_X1 U15735 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12583) );
  AOI22_X1 U15736 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9638), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12582) );
  INV_X1 U15737 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13860) );
  OR2_X1 U15738 ( .A1(n12594), .A2(n13860), .ZN(n12577) );
  OAI211_X1 U15739 ( .C1(n9589), .C2(n12579), .A(n12578), .B(n12577), .ZN(
        n12580) );
  INV_X1 U15740 ( .A(n12580), .ZN(n12581) );
  NAND4_X1 U15741 ( .A1(n12584), .A2(n12583), .A3(n12582), .A4(n12581), .ZN(
        n12585) );
  AND2_X1 U15742 ( .A1(n12586), .A2(n12585), .ZN(n12607) );
  AOI22_X1 U15743 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12589) );
  AOI22_X1 U15744 ( .A1(n12623), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12588) );
  NAND2_X1 U15745 ( .A1(n12589), .A2(n12588), .ZN(n12606) );
  INV_X1 U15746 ( .A(n10664), .ZN(n13701) );
  AOI22_X1 U15747 ( .A1(n12624), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12596), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12591) );
  AOI21_X1 U15748 ( .B1(n10677), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n12616), .ZN(n12590) );
  OAI211_X1 U15749 ( .C1(n13701), .C2(n12592), .A(n12591), .B(n12590), .ZN(
        n12605) );
  INV_X1 U15750 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12593) );
  OAI21_X1 U15751 ( .B1(n12594), .B2(n12593), .A(n12616), .ZN(n12600) );
  INV_X1 U15752 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12597) );
  OAI22_X1 U15753 ( .A1(n12598), .A2(n12597), .B1(n9625), .B2(n12595), .ZN(
        n12599) );
  AOI211_X1 U15754 ( .C1(n9638), .C2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n12600), .B(n12599), .ZN(n12603) );
  AOI22_X1 U15755 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9588), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12602) );
  AOI22_X1 U15756 ( .A1(n12623), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12601) );
  NAND3_X1 U15757 ( .A1(n12603), .A2(n12602), .A3(n12601), .ZN(n12604) );
  OAI21_X1 U15758 ( .B1(n12606), .B2(n12605), .A(n12604), .ZN(n12609) );
  INV_X1 U15759 ( .A(n12607), .ZN(n15060) );
  NOR3_X1 U15760 ( .A1(n15057), .A2(n12687), .A3(n15060), .ZN(n12608) );
  INV_X1 U15761 ( .A(n12608), .ZN(n12610) );
  AOI22_X1 U15762 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12624), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12612) );
  AOI22_X1 U15763 ( .A1(n10677), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9638), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12611) );
  NAND2_X1 U15764 ( .A1(n12612), .A2(n12611), .ZN(n12631) );
  INV_X1 U15765 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12615) );
  AOI22_X1 U15766 ( .A1(n12596), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12614) );
  AOI21_X1 U15767 ( .B1(n10663), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n12616), .ZN(n12613) );
  OAI211_X1 U15768 ( .C1(n9589), .C2(n12615), .A(n12614), .B(n12613), .ZN(
        n12630) );
  OAI21_X1 U15769 ( .B1(n12618), .B2(n12617), .A(n12616), .ZN(n12622) );
  INV_X1 U15770 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12620) );
  OAI22_X1 U15771 ( .A1(n9642), .A2(n20770), .B1(n13701), .B2(n12620), .ZN(
        n12621) );
  AOI211_X1 U15772 ( .C1(n12623), .C2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A(
        n12622), .B(n12621), .ZN(n12628) );
  AOI22_X1 U15773 ( .A1(n12596), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9587), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12627) );
  AOI22_X1 U15774 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12624), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12626) );
  NAND3_X1 U15775 ( .A1(n12628), .A2(n12627), .A3(n12626), .ZN(n12629) );
  OAI21_X1 U15776 ( .B1(n12631), .B2(n12630), .A(n12629), .ZN(n12632) );
  INV_X1 U15777 ( .A(n12632), .ZN(n12633) );
  XNOR2_X1 U15778 ( .A(n12634), .B(n12633), .ZN(n14310) );
  NAND2_X1 U15779 ( .A1(n12652), .A2(n10753), .ZN(n12635) );
  MUX2_X1 U15780 ( .A(n12635), .B(n10546), .S(n12638), .Z(n12647) );
  INV_X1 U15781 ( .A(n12643), .ZN(n12637) );
  OAI21_X1 U15782 ( .B1(n10753), .B2(n12637), .A(n12636), .ZN(n12640) );
  NAND2_X1 U15783 ( .A1(n12687), .A2(n12638), .ZN(n12639) );
  NAND2_X1 U15784 ( .A1(n12640), .A2(n12639), .ZN(n12641) );
  NAND2_X1 U15785 ( .A1(n12641), .A2(n19765), .ZN(n12645) );
  OAI21_X1 U15786 ( .B1(n12643), .B2(n12642), .A(n9628), .ZN(n12644) );
  NAND2_X1 U15787 ( .A1(n12645), .A2(n12644), .ZN(n12646) );
  NAND2_X1 U15788 ( .A1(n12647), .A2(n12646), .ZN(n12649) );
  MUX2_X1 U15789 ( .A(n10546), .B(n12649), .S(n12648), .Z(n12650) );
  NAND2_X1 U15790 ( .A1(n12650), .A2(n19747), .ZN(n12651) );
  MUX2_X1 U15791 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n12651), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n13304) );
  INV_X1 U15792 ( .A(n19747), .ZN(n12653) );
  AND3_X1 U15793 ( .A1(n19103), .A2(n12687), .A3(n12678), .ZN(n12656) );
  NAND2_X1 U15794 ( .A1(n9616), .A2(n13078), .ZN(n13685) );
  NAND2_X1 U15795 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19756) );
  AND2_X1 U15796 ( .A1(n12658), .A2(n19756), .ZN(n13695) );
  NAND2_X1 U15797 ( .A1(n12660), .A2(n12659), .ZN(n13336) );
  INV_X1 U15798 ( .A(n12694), .ZN(n13204) );
  NOR4_X1 U15799 ( .A1(P2_ADDRESS_REG_16__SCAN_IN), .A2(
        P2_ADDRESS_REG_15__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n12665) );
  NOR4_X1 U15800 ( .A1(P2_ADDRESS_REG_20__SCAN_IN), .A2(
        P2_ADDRESS_REG_19__SCAN_IN), .A3(P2_ADDRESS_REG_18__SCAN_IN), .A4(
        P2_ADDRESS_REG_17__SCAN_IN), .ZN(n12664) );
  NOR4_X1 U15801 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12663) );
  NOR4_X1 U15802 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12662) );
  NAND4_X1 U15803 ( .A1(n12665), .A2(n12664), .A3(n12663), .A4(n12662), .ZN(
        n12670) );
  NOR4_X1 U15804 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_10__SCAN_IN), .A4(
        P2_ADDRESS_REG_25__SCAN_IN), .ZN(n12668) );
  NOR4_X1 U15805 ( .A1(P2_ADDRESS_REG_24__SCAN_IN), .A2(
        P2_ADDRESS_REG_23__SCAN_IN), .A3(P2_ADDRESS_REG_22__SCAN_IN), .A4(
        P2_ADDRESS_REG_21__SCAN_IN), .ZN(n12667) );
  NOR4_X1 U15806 ( .A1(P2_ADDRESS_REG_13__SCAN_IN), .A2(
        P2_ADDRESS_REG_28__SCAN_IN), .A3(P2_ADDRESS_REG_27__SCAN_IN), .A4(
        P2_ADDRESS_REG_26__SCAN_IN), .ZN(n12666) );
  NAND4_X1 U15807 ( .A1(n12668), .A2(n12667), .A3(n12666), .A4(n19653), .ZN(
        n12669) );
  INV_X1 U15808 ( .A(n18955), .ZN(n15132) );
  INV_X1 U15809 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n12676) );
  INV_X1 U15810 ( .A(n12671), .ZN(n12684) );
  NAND2_X1 U15811 ( .A1(n13850), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12674) );
  INV_X1 U15812 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n12672) );
  OR2_X1 U15813 ( .A1(n13850), .A2(n12672), .ZN(n12673) );
  NAND2_X1 U15814 ( .A1(n12674), .A2(n12673), .ZN(n18963) );
  AOI22_X1 U15815 ( .A1(n16235), .A2(n18963), .B1(n19015), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n12675) );
  OAI21_X1 U15816 ( .B1(n15132), .B2(n12676), .A(n12675), .ZN(n12801) );
  NAND2_X1 U15817 ( .A1(n12714), .A2(n12679), .ZN(n12682) );
  NAND2_X1 U15818 ( .A1(n12770), .A2(n13204), .ZN(n12702) );
  MUX2_X1 U15819 ( .A(n9622), .B(n20827), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12681) );
  NAND3_X1 U15820 ( .A1(n12682), .A2(n12702), .A3(n12681), .ZN(n13378) );
  INV_X1 U15821 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18848) );
  OR2_X1 U15822 ( .A1(n12706), .A2(n18848), .ZN(n12690) );
  NAND2_X1 U15823 ( .A1(n12685), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n12686) );
  OAI211_X1 U15824 ( .C1(n12687), .C2(n13345), .A(n12686), .B(n19737), .ZN(
        n12688) );
  INV_X1 U15825 ( .A(n12688), .ZN(n12689) );
  NAND2_X1 U15826 ( .A1(n12690), .A2(n12689), .ZN(n13377) );
  NOR2_X1 U15827 ( .A1(n9622), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12705) );
  AOI22_X1 U15828 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n12705), .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n12692) );
  INV_X1 U15829 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20772) );
  OR2_X1 U15830 ( .A1(n12706), .A2(n20772), .ZN(n12691) );
  NAND2_X1 U15831 ( .A1(n12692), .A2(n12691), .ZN(n12698) );
  XNOR2_X1 U15832 ( .A(n13380), .B(n12698), .ZN(n13324) );
  INV_X1 U15833 ( .A(n12757), .ZN(n12704) );
  OR2_X1 U15834 ( .A1(n12693), .A2(n12704), .ZN(n12697) );
  NAND2_X1 U15835 ( .A1(n12694), .A2(n9622), .ZN(n12695) );
  MUX2_X1 U15836 ( .A(n12695), .B(n19735), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12696) );
  NAND2_X1 U15837 ( .A1(n12697), .A2(n12696), .ZN(n13325) );
  NOR2_X1 U15838 ( .A1(n13324), .A2(n13325), .ZN(n12700) );
  NOR2_X1 U15839 ( .A1(n13380), .A2(n12698), .ZN(n12699) );
  NAND2_X1 U15840 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12701) );
  OAI211_X1 U15841 ( .C1(n12704), .C2(n12703), .A(n12702), .B(n12701), .ZN(
        n12710) );
  XNOR2_X1 U15842 ( .A(n12709), .B(n12710), .ZN(n13439) );
  AOI22_X1 U15843 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n12708) );
  INV_X1 U15844 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19652) );
  OR2_X1 U15845 ( .A1(n12706), .A2(n19652), .ZN(n12707) );
  NAND2_X1 U15846 ( .A1(n12708), .A2(n12707), .ZN(n13438) );
  NOR2_X1 U15847 ( .A1(n13439), .A2(n13438), .ZN(n13440) );
  NOR2_X1 U15848 ( .A1(n12709), .A2(n12710), .ZN(n12711) );
  INV_X1 U15849 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n12713) );
  OR2_X1 U15850 ( .A1(n12706), .A2(n12713), .ZN(n12719) );
  AOI22_X1 U15851 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12718) );
  NAND2_X1 U15852 ( .A1(n12795), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12717) );
  NAND2_X1 U15853 ( .A1(n12757), .A2(n12715), .ZN(n12716) );
  NAND4_X1 U15854 ( .A1(n12719), .A2(n12718), .A3(n12717), .A4(n12716), .ZN(
        n13803) );
  NAND2_X1 U15855 ( .A1(n13804), .A2(n13803), .ZN(n13805) );
  AOI22_X1 U15856 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n12724) );
  INV_X1 U15857 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12720) );
  OR2_X1 U15858 ( .A1(n12706), .A2(n12720), .ZN(n12723) );
  NAND2_X1 U15859 ( .A1(n12757), .A2(n12721), .ZN(n12722) );
  AOI22_X1 U15860 ( .A1(n12712), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n12770), 
        .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12728) );
  INV_X1 U15861 ( .A(n12725), .ZN(n12726) );
  AOI22_X1 U15862 ( .A1(n12757), .A2(n12726), .B1(n12795), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n12727) );
  NAND2_X1 U15863 ( .A1(n12728), .A2(n12727), .ZN(n16302) );
  NAND2_X1 U15864 ( .A1(n13834), .A2(n16302), .ZN(n16301) );
  NAND2_X1 U15865 ( .A1(n12757), .A2(n12729), .ZN(n13958) );
  NAND2_X1 U15866 ( .A1(n16301), .A2(n13958), .ZN(n12732) );
  AOI22_X1 U15867 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n12731) );
  INV_X1 U15868 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19657) );
  OR2_X1 U15869 ( .A1(n12706), .A2(n19657), .ZN(n12730) );
  NAND2_X1 U15870 ( .A1(n12731), .A2(n12730), .ZN(n13957) );
  NAND2_X1 U15871 ( .A1(n12732), .A2(n13957), .ZN(n13961) );
  NAND2_X1 U15872 ( .A1(n12757), .A2(n15220), .ZN(n12733) );
  AOI22_X1 U15873 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n12735) );
  INV_X1 U15874 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19659) );
  OR2_X1 U15875 ( .A1(n12706), .A2(n19659), .ZN(n12734) );
  NAND2_X1 U15876 ( .A1(n12735), .A2(n12734), .ZN(n13778) );
  AOI22_X1 U15877 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n12739) );
  INV_X1 U15878 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n12736) );
  OR2_X1 U15879 ( .A1(n12706), .A2(n12736), .ZN(n12738) );
  NAND2_X1 U15880 ( .A1(n12757), .A2(n13416), .ZN(n12737) );
  INV_X1 U15881 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n12742) );
  AOI22_X1 U15882 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n12741) );
  NAND2_X1 U15883 ( .A1(n12757), .A2(n9655), .ZN(n12740) );
  OAI211_X1 U15884 ( .C1(n12706), .C2(n12742), .A(n12741), .B(n12740), .ZN(
        n16288) );
  AOI22_X1 U15885 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n12745) );
  INV_X1 U15886 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n13995) );
  OR2_X1 U15887 ( .A1(n12706), .A2(n13995), .ZN(n12744) );
  NAND2_X1 U15888 ( .A1(n12757), .A2(n12223), .ZN(n12743) );
  INV_X1 U15889 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n12748) );
  AOI22_X1 U15890 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n12747) );
  NAND2_X1 U15891 ( .A1(n12757), .A2(n9661), .ZN(n12746) );
  OAI211_X1 U15892 ( .C1(n12706), .C2(n12748), .A(n12747), .B(n12746), .ZN(
        n13946) );
  AOI22_X1 U15893 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n12752) );
  INV_X1 U15894 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n12749) );
  OR2_X1 U15895 ( .A1(n12706), .A2(n12749), .ZN(n12751) );
  NAND2_X1 U15896 ( .A1(n12757), .A2(n13666), .ZN(n12750) );
  INV_X1 U15897 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n12756) );
  AOI22_X1 U15898 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n12755) );
  INV_X1 U15899 ( .A(n12753), .ZN(n13901) );
  NAND2_X1 U15900 ( .A1(n12714), .A2(n13901), .ZN(n12754) );
  OAI211_X1 U15901 ( .C1(n12706), .C2(n12756), .A(n12755), .B(n12754), .ZN(
        n15703) );
  NAND2_X1 U15902 ( .A1(n13936), .A2(n15703), .ZN(n15693) );
  INV_X2 U15903 ( .A(n15693), .ZN(n12762) );
  NAND2_X1 U15904 ( .A1(n12712), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n12760) );
  AOI22_X1 U15905 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n12759) );
  NAND2_X1 U15906 ( .A1(n12757), .A2(n12291), .ZN(n12758) );
  AOI22_X1 U15907 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n12765) );
  INV_X1 U15908 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19667) );
  OR2_X1 U15909 ( .A1(n12706), .A2(n19667), .ZN(n12764) );
  NAND2_X1 U15910 ( .A1(n12757), .A2(n14045), .ZN(n12763) );
  AOI22_X1 U15911 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n12767) );
  INV_X1 U15912 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19669) );
  OR2_X1 U15913 ( .A1(n12706), .A2(n19669), .ZN(n12766) );
  NAND2_X1 U15914 ( .A1(n12767), .A2(n12766), .ZN(n14051) );
  INV_X1 U15915 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19671) );
  OR2_X1 U15916 ( .A1(n12706), .A2(n19671), .ZN(n12769) );
  AOI22_X1 U15917 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n12768) );
  AND2_X1 U15918 ( .A1(n12769), .A2(n12768), .ZN(n15019) );
  NAND2_X1 U15919 ( .A1(n12712), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n12772) );
  AOI22_X1 U15920 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n12771) );
  NOR2_X4 U15921 ( .A1(n15197), .A2(n15196), .ZN(n15006) );
  AOI22_X1 U15922 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12774) );
  INV_X1 U15923 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19675) );
  OR2_X1 U15924 ( .A1(n12706), .A2(n19675), .ZN(n12773) );
  NAND2_X1 U15925 ( .A1(n12774), .A2(n12773), .ZN(n15004) );
  AOI22_X1 U15926 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n12776) );
  INV_X1 U15927 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19677) );
  OR2_X1 U15928 ( .A1(n12706), .A2(n19677), .ZN(n12775) );
  NAND2_X1 U15929 ( .A1(n12776), .A2(n12775), .ZN(n15189) );
  INV_X1 U15930 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20763) );
  OR2_X1 U15931 ( .A1(n12706), .A2(n20763), .ZN(n12778) );
  AOI22_X1 U15932 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n12777) );
  NAND2_X1 U15933 ( .A1(n12712), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12780) );
  AOI22_X1 U15934 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n12779) );
  AND2_X1 U15935 ( .A1(n12780), .A2(n12779), .ZN(n15173) );
  AOI22_X1 U15936 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n12782) );
  INV_X1 U15937 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19682) );
  OR2_X1 U15938 ( .A1(n12706), .A2(n19682), .ZN(n12781) );
  NAND2_X1 U15939 ( .A1(n12782), .A2(n12781), .ZN(n15163) );
  AOI22_X1 U15940 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n12784) );
  INV_X1 U15941 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19684) );
  OR2_X1 U15942 ( .A1(n12706), .A2(n19684), .ZN(n12783) );
  NAND2_X1 U15943 ( .A1(n12784), .A2(n12783), .ZN(n14980) );
  OR2_X1 U15944 ( .A1(n12706), .A2(n19686), .ZN(n12786) );
  AOI22_X1 U15945 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n12785) );
  NAND2_X1 U15946 ( .A1(n12712), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12788) );
  AOI22_X1 U15947 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n12787) );
  NAND2_X1 U15948 ( .A1(n12712), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12790) );
  AOI22_X1 U15949 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n12789) );
  AND2_X1 U15950 ( .A1(n12790), .A2(n12789), .ZN(n14950) );
  AOI22_X1 U15951 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n12792) );
  INV_X1 U15952 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19691) );
  OR2_X1 U15953 ( .A1(n12706), .A2(n19691), .ZN(n12791) );
  NAND2_X1 U15954 ( .A1(n12792), .A2(n12791), .ZN(n15133) );
  AND2_X2 U15955 ( .A1(n15134), .A2(n15133), .ZN(n15136) );
  AOI22_X1 U15956 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n12794) );
  INV_X1 U15957 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19693) );
  OR2_X1 U15958 ( .A1(n12706), .A2(n19693), .ZN(n12793) );
  NAND2_X1 U15959 ( .A1(n12794), .A2(n12793), .ZN(n14932) );
  NAND2_X1 U15960 ( .A1(n12712), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12797) );
  AOI22_X1 U15961 ( .A1(n12770), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n12795), .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n12796) );
  NAND2_X1 U15962 ( .A1(n12797), .A2(n12796), .ZN(n12798) );
  NOR2_X1 U15963 ( .A1(n15479), .A2(n15206), .ZN(n12800) );
  AOI211_X1 U15964 ( .C1(BUF1_REG_30__SCAN_IN), .C2(n18957), .A(n12801), .B(
        n12800), .ZN(n12802) );
  OAI21_X1 U15965 ( .B1(n14310), .B2(n15185), .A(n12802), .ZN(P2_U2889) );
  INV_X1 U15966 ( .A(n12804), .ZN(n12805) );
  NOR2_X1 U15967 ( .A1(n12805), .A2(n12817), .ZN(n12806) );
  INV_X1 U15968 ( .A(n12807), .ZN(n12808) );
  NAND2_X1 U15969 ( .A1(n12808), .A2(n11367), .ZN(n12813) );
  NAND2_X1 U15970 ( .A1(n12809), .A2(n12814), .ZN(n12831) );
  OAI21_X1 U15971 ( .B1(n12814), .B2(n12809), .A(n12831), .ZN(n12810) );
  OAI211_X1 U15972 ( .C1(n12810), .C2(n11399), .A(n11373), .B(n12070), .ZN(
        n12811) );
  INV_X1 U15973 ( .A(n12811), .ZN(n12812) );
  NAND2_X1 U15974 ( .A1(n20024), .A2(n11371), .ZN(n12824) );
  OAI21_X1 U15975 ( .B1(n11399), .B2(n12814), .A(n12824), .ZN(n12815) );
  INV_X1 U15976 ( .A(n12815), .ZN(n12816) );
  OAI21_X2 U15977 ( .B1(n12818), .B2(n12817), .A(n12816), .ZN(n13299) );
  INV_X1 U15978 ( .A(n12819), .ZN(n12820) );
  OR2_X1 U15979 ( .A1(n13298), .A2(n12820), .ZN(n12821) );
  NAND2_X2 U15980 ( .A1(n20005), .A2(n12821), .ZN(n12827) );
  XNOR2_X1 U15981 ( .A(n12831), .B(n12823), .ZN(n12825) );
  OAI21_X1 U15982 ( .B1(n12825), .B2(n11399), .A(n12824), .ZN(n12826) );
  NAND2_X1 U15983 ( .A1(n12827), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12828) );
  INV_X1 U15984 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12829) );
  NAND2_X1 U15985 ( .A1(n20642), .A2(n12865), .ZN(n12835) );
  NAND2_X1 U15986 ( .A1(n12831), .A2(n12830), .ZN(n12849) );
  INV_X1 U15987 ( .A(n12847), .ZN(n12832) );
  XNOR2_X1 U15988 ( .A(n12849), .B(n12832), .ZN(n12833) );
  NAND2_X1 U15989 ( .A1(n12833), .A2(n12877), .ZN(n12834) );
  NAND2_X1 U15990 ( .A1(n12835), .A2(n12834), .ZN(n13539) );
  NAND2_X1 U15991 ( .A1(n12836), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12837) );
  NAND2_X1 U15992 ( .A1(n12838), .A2(n12865), .ZN(n12842) );
  NAND2_X1 U15993 ( .A1(n12849), .A2(n12847), .ZN(n12839) );
  XNOR2_X1 U15994 ( .A(n12839), .B(n12846), .ZN(n12840) );
  NAND2_X1 U15995 ( .A1(n12840), .A2(n12877), .ZN(n12841) );
  INV_X1 U15996 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12936) );
  NAND2_X1 U15997 ( .A1(n12843), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12844) );
  NAND2_X1 U15998 ( .A1(n12845), .A2(n12865), .ZN(n12852) );
  AND2_X1 U15999 ( .A1(n12847), .A2(n12846), .ZN(n12848) );
  NAND2_X1 U16000 ( .A1(n12849), .A2(n12848), .ZN(n12856) );
  XNOR2_X1 U16001 ( .A(n12856), .B(n12857), .ZN(n12850) );
  NAND2_X1 U16002 ( .A1(n12850), .A2(n12877), .ZN(n12851) );
  NAND2_X1 U16003 ( .A1(n12852), .A2(n12851), .ZN(n12853) );
  INV_X1 U16004 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16155) );
  XNOR2_X1 U16005 ( .A(n12853), .B(n16155), .ZN(n16055) );
  NAND2_X1 U16006 ( .A1(n12853), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12854) );
  INV_X1 U16007 ( .A(n12856), .ZN(n12858) );
  NAND2_X1 U16008 ( .A1(n12858), .A2(n12857), .ZN(n12867) );
  XNOR2_X1 U16009 ( .A(n12867), .B(n12868), .ZN(n12859) );
  NAND2_X1 U16010 ( .A1(n12859), .A2(n12877), .ZN(n12860) );
  INV_X1 U16011 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16149) );
  NAND2_X1 U16012 ( .A1(n16050), .A2(n16149), .ZN(n12862) );
  INV_X1 U16013 ( .A(n16050), .ZN(n12863) );
  NAND2_X1 U16014 ( .A1(n12863), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12864) );
  NAND2_X1 U16015 ( .A1(n12866), .A2(n12865), .ZN(n12872) );
  INV_X1 U16016 ( .A(n12867), .ZN(n12869) );
  NAND2_X1 U16017 ( .A1(n12869), .A2(n12868), .ZN(n12875) );
  XNOR2_X1 U16018 ( .A(n12875), .B(n12876), .ZN(n12870) );
  NAND2_X1 U16019 ( .A1(n12870), .A2(n12877), .ZN(n12871) );
  NAND2_X1 U16020 ( .A1(n12872), .A2(n12871), .ZN(n12873) );
  NAND2_X1 U16021 ( .A1(n12873), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16044) );
  INV_X1 U16022 ( .A(n12875), .ZN(n12878) );
  NAND3_X1 U16023 ( .A1(n12878), .A2(n12877), .A3(n12876), .ZN(n12879) );
  NAND2_X1 U16024 ( .A1(n12874), .A2(n12879), .ZN(n14088) );
  OR2_X1 U16025 ( .A1(n14088), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12880) );
  NAND2_X1 U16026 ( .A1(n14088), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12881) );
  INV_X1 U16027 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n14150) );
  NAND2_X1 U16028 ( .A1(n14844), .A2(n14150), .ZN(n12883) );
  NAND2_X1 U16029 ( .A1(n14841), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14707) );
  INV_X1 U16030 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14855) );
  NAND2_X1 U16031 ( .A1(n12874), .A2(n14855), .ZN(n12884) );
  NAND2_X1 U16032 ( .A1(n14707), .A2(n12884), .ZN(n14722) );
  INV_X1 U16033 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16098) );
  NAND2_X1 U16034 ( .A1(n12874), .A2(n16098), .ZN(n14720) );
  NAND2_X1 U16035 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12885) );
  NAND2_X1 U16036 ( .A1(n12874), .A2(n12885), .ZN(n14716) );
  NAND2_X1 U16037 ( .A1(n14720), .A2(n14716), .ZN(n12886) );
  NOR2_X1 U16038 ( .A1(n14722), .A2(n12886), .ZN(n14706) );
  INV_X1 U16039 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16081) );
  NAND2_X1 U16040 ( .A1(n14844), .A2(n16081), .ZN(n12887) );
  NAND2_X1 U16041 ( .A1(n14706), .A2(n12887), .ZN(n14842) );
  INV_X1 U16042 ( .A(n14842), .ZN(n12888) );
  INV_X1 U16043 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14869) );
  NAND2_X1 U16044 ( .A1(n14844), .A2(n14869), .ZN(n14863) );
  OAI21_X1 U16045 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(n14841), .ZN(n12889) );
  INV_X1 U16046 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12890) );
  NAND2_X1 U16047 ( .A1(n14844), .A2(n12890), .ZN(n12891) );
  NAND2_X1 U16048 ( .A1(n14841), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14864) );
  NOR2_X1 U16049 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14845) );
  NOR2_X1 U16050 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14705) );
  NAND3_X1 U16051 ( .A1(n14845), .A2(n14705), .A3(n16098), .ZN(n12892) );
  NAND2_X1 U16052 ( .A1(n14841), .A2(n12892), .ZN(n14865) );
  XNOR2_X1 U16053 ( .A(n14844), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14688) );
  NAND2_X1 U16054 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14662) );
  INV_X1 U16055 ( .A(n14662), .ZN(n12893) );
  INV_X1 U16056 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12896) );
  NAND3_X1 U16057 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14595) );
  INV_X1 U16058 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14797) );
  INV_X1 U16059 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14775) );
  INV_X1 U16060 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14801) );
  NAND3_X1 U16061 ( .A1(n14797), .A2(n14775), .A3(n14801), .ZN(n14596) );
  AND2_X1 U16062 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13065) );
  INV_X1 U16063 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14600) );
  INV_X1 U16064 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14609) );
  NAND2_X1 U16065 ( .A1(n14600), .A2(n14609), .ZN(n14757) );
  NAND2_X1 U16066 ( .A1(n12897), .A2(n20564), .ZN(n15859) );
  NAND2_X1 U16067 ( .A1(n11367), .A2(n15859), .ZN(n12898) );
  NAND2_X1 U16068 ( .A1(n13544), .A2(n12898), .ZN(n12907) );
  INV_X1 U16069 ( .A(n12899), .ZN(n12903) );
  AND2_X1 U16070 ( .A1(n13048), .A2(n11372), .ZN(n12900) );
  NAND2_X1 U16071 ( .A1(n11403), .A2(n12900), .ZN(n13041) );
  NAND2_X1 U16072 ( .A1(n12901), .A2(n13041), .ZN(n12902) );
  NAND2_X1 U16073 ( .A1(n12903), .A2(n12902), .ZN(n13547) );
  INV_X1 U16074 ( .A(n13048), .ZN(n12904) );
  NAND2_X1 U16075 ( .A1(n13599), .A2(n12904), .ZN(n12905) );
  OAI211_X1 U16076 ( .C1(n12907), .C2(n12906), .A(n13547), .B(n12905), .ZN(
        n12908) );
  NAND2_X1 U16077 ( .A1(n12908), .A2(n14301), .ZN(n12914) );
  NAND2_X1 U16078 ( .A1(n11366), .A2(n15859), .ZN(n13629) );
  NAND2_X1 U16079 ( .A1(n13549), .A2(n13629), .ZN(n12910) );
  NAND3_X1 U16080 ( .A1(n12910), .A2(n11372), .A3(n12909), .ZN(n12912) );
  NAND3_X1 U16081 ( .A1(n12912), .A2(n13264), .A3(n12911), .ZN(n12913) );
  AND2_X1 U16082 ( .A1(n12915), .A2(n13561), .ZN(n12919) );
  INV_X1 U16083 ( .A(n13265), .ZN(n15827) );
  NAND2_X1 U16084 ( .A1(n12916), .A2(n12917), .ZN(n12918) );
  NAND4_X1 U16085 ( .A1(n12919), .A2(n15827), .A3(n12048), .A4(n12918), .ZN(
        n12920) );
  MUX2_X1 U16086 ( .A(n13025), .B(n13009), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n12925) );
  NAND2_X1 U16087 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13285), .ZN(
        n12923) );
  NAND2_X1 U16088 ( .A1(n12925), .A2(n12924), .ZN(n12929) );
  NAND2_X1 U16089 ( .A1(n13009), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12928) );
  INV_X1 U16090 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n12926) );
  NAND2_X1 U16091 ( .A1(n12949), .A2(n12926), .ZN(n12927) );
  NAND2_X1 U16092 ( .A1(n12928), .A2(n12927), .ZN(n13273) );
  XNOR2_X1 U16093 ( .A(n12929), .B(n13273), .ZN(n13284) );
  NAND2_X1 U16094 ( .A1(n13284), .A2(n13630), .ZN(n13288) );
  NAND2_X1 U16095 ( .A1(n13288), .A2(n12929), .ZN(n13461) );
  MUX2_X1 U16096 ( .A(n13025), .B(n13009), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n12931) );
  NAND2_X1 U16097 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13285), .ZN(
        n12930) );
  AND3_X1 U16098 ( .A1(n12931), .A2(n12990), .A3(n12930), .ZN(n13460) );
  INV_X1 U16099 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n12932) );
  NAND2_X1 U16100 ( .A1(n13630), .A2(n12932), .ZN(n12934) );
  NAND2_X1 U16101 ( .A1(n12939), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12933) );
  NAND3_X1 U16102 ( .A1(n12934), .A2(n13009), .A3(n12933), .ZN(n12935) );
  OAI21_X1 U16103 ( .B1(n13016), .B2(P1_EBX_REG_3__SCAN_IN), .A(n12935), .ZN(
        n13536) );
  OR2_X1 U16104 ( .A1(n13025), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n12942) );
  NAND2_X1 U16105 ( .A1(n13009), .A2(n12936), .ZN(n12940) );
  INV_X1 U16106 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n12937) );
  NAND2_X1 U16107 ( .A1(n13630), .A2(n12937), .ZN(n12938) );
  NAND3_X1 U16108 ( .A1(n12940), .A2(n12939), .A3(n12938), .ZN(n12941) );
  NAND2_X1 U16109 ( .A1(n12942), .A2(n12941), .ZN(n13614) );
  MUX2_X1 U16110 ( .A(n13016), .B(n12939), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n12944) );
  OAI21_X1 U16111 ( .B1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n12943), .A(
        n12944), .ZN(n13683) );
  MUX2_X1 U16112 ( .A(n13025), .B(n13009), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12948) );
  NAND2_X1 U16113 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13285), .ZN(
        n12947) );
  INV_X1 U16114 ( .A(n13016), .ZN(n12999) );
  INV_X1 U16115 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n19898) );
  NAND2_X1 U16116 ( .A1(n12999), .A2(n19898), .ZN(n12953) );
  NAND2_X1 U16117 ( .A1(n13630), .A2(n19898), .ZN(n12951) );
  NAND2_X1 U16118 ( .A1(n12939), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12950) );
  NAND3_X1 U16119 ( .A1(n12951), .A2(n13009), .A3(n12950), .ZN(n12952) );
  OR2_X1 U16120 ( .A1(n13025), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n12958) );
  INV_X1 U16121 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12954) );
  NAND2_X1 U16122 ( .A1(n13009), .A2(n12954), .ZN(n12956) );
  INV_X1 U16123 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n19822) );
  NAND2_X1 U16124 ( .A1(n13630), .A2(n19822), .ZN(n12955) );
  NAND3_X1 U16125 ( .A1(n12956), .A2(n12939), .A3(n12955), .ZN(n12957) );
  NAND2_X1 U16126 ( .A1(n12958), .A2(n12957), .ZN(n14017) );
  NAND2_X1 U16127 ( .A1(n14016), .A2(n14017), .ZN(n14145) );
  MUX2_X1 U16128 ( .A(n13016), .B(n12939), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n12959) );
  OAI21_X1 U16129 ( .B1(n12943), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n12959), .ZN(n14146) );
  MUX2_X1 U16130 ( .A(n13025), .B(n13009), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n12963) );
  NAND2_X1 U16131 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n13285), .ZN(
        n12962) );
  INV_X1 U16132 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14533) );
  NAND2_X1 U16133 ( .A1(n12999), .A2(n14533), .ZN(n12967) );
  NAND2_X1 U16134 ( .A1(n13630), .A2(n14533), .ZN(n12965) );
  NAND2_X1 U16135 ( .A1(n12939), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12964) );
  NAND3_X1 U16136 ( .A1(n12965), .A2(n13009), .A3(n12964), .ZN(n12966) );
  OR2_X1 U16137 ( .A1(n13025), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n12971) );
  NAND2_X1 U16138 ( .A1(n13009), .A2(n16098), .ZN(n12969) );
  INV_X1 U16139 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15969) );
  NAND2_X1 U16140 ( .A1(n13630), .A2(n15969), .ZN(n12968) );
  NAND3_X1 U16141 ( .A1(n12969), .A2(n12939), .A3(n12968), .ZN(n12970) );
  NAND2_X1 U16142 ( .A1(n12971), .A2(n12970), .ZN(n14520) );
  NAND2_X1 U16143 ( .A1(n14528), .A2(n14520), .ZN(n14451) );
  INV_X1 U16144 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14512) );
  NAND2_X1 U16145 ( .A1(n13630), .A2(n14512), .ZN(n12973) );
  NAND2_X1 U16146 ( .A1(n12939), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12972) );
  NAND3_X1 U16147 ( .A1(n12973), .A2(n13009), .A3(n12972), .ZN(n12974) );
  OAI21_X1 U16148 ( .B1(n13016), .B2(P1_EBX_REG_13__SCAN_IN), .A(n12974), .ZN(
        n14452) );
  MUX2_X1 U16149 ( .A(n13016), .B(n12939), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12975) );
  OAI21_X1 U16150 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n12943), .A(
        n12975), .ZN(n12976) );
  INV_X1 U16151 ( .A(n12976), .ZN(n14501) );
  OR2_X1 U16152 ( .A1(n13025), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n12980) );
  NAND2_X1 U16153 ( .A1(n13009), .A2(n16081), .ZN(n12978) );
  INV_X1 U16154 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15959) );
  NAND2_X1 U16155 ( .A1(n13630), .A2(n15959), .ZN(n12977) );
  NAND3_X1 U16156 ( .A1(n12978), .A2(n12939), .A3(n12977), .ZN(n12979) );
  NAND2_X1 U16157 ( .A1(n12980), .A2(n12979), .ZN(n14508) );
  NAND2_X1 U16158 ( .A1(n14501), .A2(n14508), .ZN(n12981) );
  OR2_X1 U16159 ( .A1(n13025), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n12985) );
  INV_X1 U16160 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16076) );
  NAND2_X1 U16161 ( .A1(n13009), .A2(n16076), .ZN(n12983) );
  INV_X1 U16162 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15946) );
  NAND2_X1 U16163 ( .A1(n13630), .A2(n15946), .ZN(n12982) );
  NAND3_X1 U16164 ( .A1(n12983), .A2(n12939), .A3(n12982), .ZN(n12984) );
  NAND2_X1 U16165 ( .A1(n12985), .A2(n12984), .ZN(n14493) );
  INV_X1 U16166 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n15995) );
  NAND2_X1 U16167 ( .A1(n13630), .A2(n15995), .ZN(n12987) );
  NAND2_X1 U16168 ( .A1(n12939), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12986) );
  NAND3_X1 U16169 ( .A1(n12987), .A2(n13009), .A3(n12986), .ZN(n12988) );
  OAI21_X1 U16170 ( .B1(n13016), .B2(P1_EBX_REG_17__SCAN_IN), .A(n12988), .ZN(
        n14860) );
  MUX2_X1 U16171 ( .A(n13025), .B(n13009), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n12991) );
  NAND2_X1 U16172 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n13285), .ZN(
        n12989) );
  AND3_X1 U16173 ( .A1(n12991), .A2(n12990), .A3(n12989), .ZN(n14487) );
  INV_X1 U16174 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n15992) );
  NAND2_X1 U16175 ( .A1(n13630), .A2(n15992), .ZN(n12993) );
  NAND2_X1 U16176 ( .A1(n12939), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12992) );
  NAND3_X1 U16177 ( .A1(n12993), .A2(n13009), .A3(n12992), .ZN(n12994) );
  OAI21_X1 U16178 ( .B1(n13016), .B2(P1_EBX_REG_19__SCAN_IN), .A(n12994), .ZN(
        n14835) );
  NOR2_X4 U16179 ( .A1(n14834), .A2(n14835), .ZN(n14833) );
  OR2_X1 U16180 ( .A1(n13025), .A2(P1_EBX_REG_20__SCAN_IN), .ZN(n12998) );
  INV_X1 U16181 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15867) );
  NAND2_X1 U16182 ( .A1(n13009), .A2(n15867), .ZN(n12996) );
  INV_X1 U16183 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15902) );
  NAND2_X1 U16184 ( .A1(n13630), .A2(n15902), .ZN(n12995) );
  NAND3_X1 U16185 ( .A1(n12996), .A2(n12939), .A3(n12995), .ZN(n12997) );
  NAND2_X1 U16186 ( .A1(n12998), .A2(n12997), .ZN(n14480) );
  INV_X1 U16187 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15989) );
  NAND2_X1 U16188 ( .A1(n12999), .A2(n15989), .ZN(n13003) );
  NAND2_X1 U16189 ( .A1(n13630), .A2(n15989), .ZN(n13001) );
  NAND2_X1 U16190 ( .A1(n12939), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13000) );
  NAND3_X1 U16191 ( .A1(n13001), .A2(n13009), .A3(n13000), .ZN(n13002) );
  OR2_X1 U16192 ( .A1(n13025), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n13007) );
  INV_X1 U16193 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14653) );
  NAND2_X1 U16194 ( .A1(n13009), .A2(n14653), .ZN(n13005) );
  INV_X1 U16195 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15887) );
  NAND2_X1 U16196 ( .A1(n13630), .A2(n15887), .ZN(n13004) );
  NAND3_X1 U16197 ( .A1(n13005), .A2(n12939), .A3(n13004), .ZN(n13006) );
  MUX2_X1 U16198 ( .A(n13016), .B(n12939), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n13008) );
  OAI21_X1 U16199 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n12943), .A(
        n13008), .ZN(n14433) );
  MUX2_X1 U16200 ( .A(n13025), .B(n13009), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n13011) );
  NAND2_X1 U16201 ( .A1(n13285), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13010) );
  NAND2_X1 U16202 ( .A1(n13011), .A2(n13010), .ZN(n14418) );
  AND2_X2 U16203 ( .A1(n14432), .A2(n14418), .ZN(n14419) );
  MUX2_X1 U16204 ( .A(n13016), .B(n12939), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n13013) );
  OR2_X1 U16205 ( .A1(n12943), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13012) );
  MUX2_X1 U16206 ( .A(n13025), .B(n13009), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n13015) );
  NAND2_X1 U16207 ( .A1(n13285), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13014) );
  AND2_X1 U16208 ( .A1(n13015), .A2(n13014), .ZN(n14393) );
  MUX2_X1 U16209 ( .A(n13016), .B(n12939), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n13017) );
  OAI21_X1 U16210 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n12943), .A(
        n13017), .ZN(n14376) );
  OR2_X1 U16211 ( .A1(n13025), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n13022) );
  NAND2_X1 U16212 ( .A1(n13009), .A2(n14600), .ZN(n13020) );
  INV_X1 U16213 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n13018) );
  NAND2_X1 U16214 ( .A1(n13630), .A2(n13018), .ZN(n13019) );
  NAND3_X1 U16215 ( .A1(n13020), .A2(n12939), .A3(n13019), .ZN(n13021) );
  OR2_X1 U16216 ( .A1(n12943), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13024) );
  INV_X1 U16217 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14461) );
  NAND2_X1 U16218 ( .A1(n13630), .A2(n14461), .ZN(n13023) );
  NAND2_X1 U16219 ( .A1(n13024), .A2(n13023), .ZN(n14321) );
  OAI22_X1 U16220 ( .A1(n14321), .A2(n12921), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n13025), .ZN(n13026) );
  OR2_X1 U16221 ( .A1(n14362), .A2(n13026), .ZN(n13027) );
  NAND2_X1 U16222 ( .A1(n14327), .A2(n13027), .ZN(n14460) );
  NAND2_X1 U16223 ( .A1(n13029), .A2(n11366), .ZN(n13227) );
  NAND2_X1 U16224 ( .A1(n12916), .A2(n20044), .ZN(n13030) );
  NAND2_X1 U16225 ( .A1(n13227), .A2(n13030), .ZN(n13031) );
  INV_X1 U16226 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20620) );
  NOR2_X1 U16227 ( .A1(n16122), .A2(n20620), .ZN(n14587) );
  INV_X1 U16228 ( .A(n14587), .ZN(n13070) );
  INV_X1 U16229 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14750) );
  OAI21_X1 U16230 ( .B1(n12911), .B2(n13033), .A(n13032), .ZN(n13034) );
  NAND2_X1 U16231 ( .A1(n13034), .A2(n11367), .ZN(n13035) );
  OAI21_X1 U16232 ( .B1(n13038), .B2(n13037), .A(n13036), .ZN(n13039) );
  NOR2_X1 U16233 ( .A1(n13040), .A2(n13039), .ZN(n13042) );
  OAI211_X1 U16234 ( .C1(n11394), .C2(n13163), .A(n13042), .B(n13041), .ZN(
        n13569) );
  AND2_X1 U16235 ( .A1(n13043), .A2(n20024), .ZN(n13044) );
  OR2_X1 U16236 ( .A1(n13569), .A2(n13044), .ZN(n13045) );
  NOR2_X1 U16237 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13403), .ZN(
        n20007) );
  INV_X1 U16238 ( .A(n20007), .ZN(n13046) );
  INV_X1 U16239 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20011) );
  NOR2_X1 U16240 ( .A1(n20762), .A2(n20011), .ZN(n19993) );
  INV_X1 U16241 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16132) );
  NAND2_X1 U16242 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19975) );
  NOR2_X1 U16243 ( .A1(n16155), .A2(n19975), .ZN(n16145) );
  INV_X1 U16244 ( .A(n16145), .ZN(n16133) );
  NOR4_X1 U16245 ( .A1(n12954), .A2(n16132), .A3(n16149), .A4(n16133), .ZN(
        n13049) );
  INV_X1 U16246 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16114) );
  NOR2_X1 U16247 ( .A1(n16114), .A2(n14150), .ZN(n16116) );
  NAND2_X1 U16248 ( .A1(n13049), .A2(n16116), .ZN(n16092) );
  INV_X1 U16249 ( .A(n16092), .ZN(n16096) );
  NAND4_X1 U16250 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n19993), .A4(n16096), .ZN(
        n14854) );
  INV_X1 U16251 ( .A(n14854), .ZN(n13051) );
  INV_X1 U16252 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14882) );
  OAI21_X1 U16253 ( .B1(n14882), .B2(n20011), .A(n20762), .ZN(n16094) );
  NAND2_X1 U16254 ( .A1(n16094), .A2(n13049), .ZN(n16113) );
  INV_X1 U16255 ( .A(n16113), .ZN(n16124) );
  NAND4_X1 U16256 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n16116), .A4(n16124), .ZN(
        n14853) );
  NOR2_X1 U16257 ( .A1(n16095), .A2(n14853), .ZN(n13050) );
  AOI21_X1 U16258 ( .B1(n19988), .B2(n13051), .A(n13050), .ZN(n16091) );
  INV_X1 U16259 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16064) );
  NAND2_X1 U16260 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14851) );
  NOR2_X1 U16261 ( .A1(n14869), .A2(n16076), .ZN(n16070) );
  NAND2_X1 U16262 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n16070), .ZN(
        n14852) );
  OR3_X1 U16263 ( .A1(n16064), .A2(n14851), .A3(n14852), .ZN(n13056) );
  OR2_X1 U16264 ( .A1(n16091), .A2(n13056), .ZN(n15861) );
  INV_X1 U16265 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15864) );
  NOR2_X1 U16266 ( .A1(n15861), .A2(n15864), .ZN(n15868) );
  NAND2_X1 U16267 ( .A1(n15868), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14829) );
  NAND2_X1 U16268 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13060) );
  INV_X1 U16269 ( .A(n14595), .ZN(n14778) );
  NAND2_X1 U16270 ( .A1(n14778), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13052) );
  NOR2_X1 U16271 ( .A1(n14810), .A2(n13052), .ZN(n14765) );
  NAND2_X1 U16272 ( .A1(n14765), .A2(n13065), .ZN(n14751) );
  NOR2_X1 U16273 ( .A1(n13056), .A2(n14853), .ZN(n13058) );
  INV_X2 U16274 ( .A(n16122), .ZN(n20014) );
  NOR2_X1 U16275 ( .A1(n13053), .A2(n20014), .ZN(n13401) );
  INV_X1 U16276 ( .A(n13401), .ZN(n13055) );
  NAND2_X1 U16277 ( .A1(n13399), .A2(n14882), .ZN(n13054) );
  OAI21_X1 U16278 ( .B1(n13056), .B2(n14854), .A(n16093), .ZN(n13057) );
  OAI211_X1 U16279 ( .C1(n13058), .C2(n16095), .A(n19989), .B(n13057), .ZN(
        n15862) );
  OR2_X1 U16280 ( .A1(n15862), .A2(n14662), .ZN(n13059) );
  NAND2_X1 U16281 ( .A1(n20008), .A2(n19989), .ZN(n16112) );
  NAND2_X1 U16282 ( .A1(n13059), .A2(n16112), .ZN(n14828) );
  INV_X1 U16283 ( .A(n13060), .ZN(n13061) );
  OR2_X1 U16284 ( .A1(n20008), .A2(n13061), .ZN(n13062) );
  NAND2_X1 U16285 ( .A1(n14828), .A2(n13062), .ZN(n14808) );
  AOI21_X1 U16286 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(n20008), .ZN(n13063) );
  NOR2_X1 U16287 ( .A1(n14808), .A2(n13063), .ZN(n14786) );
  AND2_X1 U16288 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13064) );
  NAND2_X1 U16289 ( .A1(n14786), .A2(n13064), .ZN(n14767) );
  INV_X1 U16290 ( .A(n13065), .ZN(n14756) );
  NOR2_X1 U16291 ( .A1(n16095), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13066) );
  NOR2_X1 U16292 ( .A1(n14808), .A2(n13066), .ZN(n14795) );
  NAND2_X1 U16293 ( .A1(n14795), .A2(n20008), .ZN(n14766) );
  OAI21_X1 U16294 ( .B1(n14767), .B2(n14756), .A(n14766), .ZN(n13067) );
  AND2_X1 U16295 ( .A1(n13067), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14748) );
  AOI21_X1 U16296 ( .B1(n14750), .B2(n14751), .A(n14748), .ZN(n13068) );
  INV_X1 U16297 ( .A(n13068), .ZN(n13069) );
  NOR2_X1 U16298 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13072) );
  NOR4_X1 U16299 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13071) );
  NAND4_X1 U16300 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13072), .A4(n13071), .ZN(n13075) );
  INV_X1 U16301 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20665) );
  NOR3_X1 U16302 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20665), .ZN(n13074) );
  NOR4_X1 U16303 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13073) );
  NAND4_X1 U16304 ( .A1(n20020), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13074), .A4(
        n13073), .ZN(U214) );
  NOR2_X1 U16305 ( .A1(n13129), .A2(n13075), .ZN(n16384) );
  NAND2_X1 U16306 ( .A1(n16384), .A2(U214), .ZN(U212) );
  INV_X1 U16307 ( .A(n13317), .ZN(n13076) );
  NOR2_X1 U16308 ( .A1(n9616), .A2(n18832), .ZN(n13080) );
  NAND2_X1 U16309 ( .A1(n13076), .A2(n13080), .ZN(n13079) );
  NAND2_X1 U16310 ( .A1(n13687), .A2(n13318), .ZN(n13077) );
  NOR2_X1 U16311 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19641) );
  AOI211_X1 U16312 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(P2_STATE_REG_0__SCAN_IN), .B(n19641), .ZN(n19763) );
  INV_X1 U16313 ( .A(n19763), .ZN(n19766) );
  AND2_X2 U16314 ( .A1(n19762), .A2(n19742), .ZN(n19757) );
  NOR2_X4 U16315 ( .A1(n19023), .A2(n19757), .ZN(n19054) );
  AND2_X1 U16316 ( .A1(n19054), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NAND2_X1 U16317 ( .A1(n13080), .A2(n13687), .ZN(n14122) );
  INV_X1 U16318 ( .A(n14122), .ZN(n13083) );
  INV_X1 U16319 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13082) );
  INV_X1 U16320 ( .A(n13791), .ZN(n13081) );
  NAND2_X1 U16321 ( .A1(n19520), .A2(n19726), .ZN(n13085) );
  OAI211_X1 U16322 ( .C1(n13083), .C2(n13082), .A(n13081), .B(n13085), .ZN(
        P2_U2814) );
  NOR2_X1 U16323 ( .A1(n19758), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n13086)
         );
  INV_X1 U16324 ( .A(n12658), .ZN(n13084) );
  AOI22_X1 U16325 ( .A1(n13086), .A2(n13085), .B1(n13084), .B2(n19758), .ZN(
        P2_U3612) );
  AOI22_X1 U16326 ( .A1(n13788), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n13094), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n13087) );
  NAND3_X1 U16327 ( .A1(n13791), .A2(n10753), .A3(n19756), .ZN(n13131) );
  INV_X1 U16328 ( .A(n13131), .ZN(n13135) );
  AOI22_X1 U16329 ( .A1(n13852), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13850), .ZN(n19125) );
  INV_X1 U16330 ( .A(n19125), .ZN(n15172) );
  NAND2_X1 U16331 ( .A1(n13135), .A2(n15172), .ZN(n13097) );
  NAND2_X1 U16332 ( .A1(n13087), .A2(n13097), .ZN(P2_U2973) );
  AOI22_X1 U16333 ( .A1(n13788), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n13094), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13088) );
  AOI22_X1 U16334 ( .A1(n13852), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n13129), .ZN(n18969) );
  INV_X1 U16335 ( .A(n18969), .ZN(n15130) );
  NAND2_X1 U16336 ( .A1(n13135), .A2(n15130), .ZN(n13099) );
  NAND2_X1 U16337 ( .A1(n13088), .A2(n13099), .ZN(P2_U2979) );
  AOI22_X1 U16338 ( .A1(n13788), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n13094), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n13089) );
  AOI22_X1 U16339 ( .A1(n13852), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13129), .ZN(n18981) );
  INV_X1 U16340 ( .A(n18981), .ZN(n15165) );
  NAND2_X1 U16341 ( .A1(n13135), .A2(n15165), .ZN(n13111) );
  NAND2_X1 U16342 ( .A1(n13089), .A2(n13111), .ZN(P2_U2974) );
  AOI22_X1 U16343 ( .A1(n13788), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n13094), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13090) );
  AOI22_X1 U16344 ( .A1(n13852), .A2(BUF1_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n13850), .ZN(n18974) );
  INV_X1 U16345 ( .A(n18974), .ZN(n15149) );
  NAND2_X1 U16346 ( .A1(n13135), .A2(n15149), .ZN(n13095) );
  NAND2_X1 U16347 ( .A1(n13090), .A2(n13095), .ZN(P2_U2977) );
  AOI22_X1 U16348 ( .A1(n13788), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n13094), .B2(
        P2_LWORD_REG_9__SCAN_IN), .ZN(n13092) );
  AOI22_X1 U16349 ( .A1(n13852), .A2(BUF1_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n13850), .ZN(n18976) );
  INV_X1 U16350 ( .A(n18976), .ZN(n13091) );
  NAND2_X1 U16351 ( .A1(n13135), .A2(n13091), .ZN(n13108) );
  NAND2_X1 U16352 ( .A1(n13092), .A2(n13108), .ZN(P2_U2976) );
  AOI22_X1 U16353 ( .A1(P2_EAX_REG_16__SCAN_IN), .A2(n13788), .B1(n13094), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13093) );
  AOI22_X1 U16354 ( .A1(n13852), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13129), .ZN(n19086) );
  INV_X1 U16355 ( .A(n19086), .ZN(n14053) );
  NAND2_X1 U16356 ( .A1(n13135), .A2(n14053), .ZN(n13114) );
  NAND2_X1 U16357 ( .A1(n13093), .A2(n13114), .ZN(P2_U2952) );
  AOI22_X1 U16358 ( .A1(P2_EAX_REG_26__SCAN_IN), .A2(n13788), .B1(n13137), 
        .B2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13096) );
  NAND2_X1 U16359 ( .A1(n13096), .A2(n13095), .ZN(P2_U2962) );
  AOI22_X1 U16360 ( .A1(P2_EAX_REG_22__SCAN_IN), .A2(n13788), .B1(n13137), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13098) );
  NAND2_X1 U16361 ( .A1(n13098), .A2(n13097), .ZN(P2_U2958) );
  AOI22_X1 U16362 ( .A1(P2_EAX_REG_28__SCAN_IN), .A2(n13788), .B1(n13137), 
        .B2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13100) );
  NAND2_X1 U16363 ( .A1(n13100), .A2(n13099), .ZN(P2_U2964) );
  AOI22_X1 U16364 ( .A1(P2_EAX_REG_29__SCAN_IN), .A2(n13788), .B1(n13137), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13101) );
  AOI22_X1 U16365 ( .A1(n13852), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n13129), .ZN(n18966) );
  INV_X1 U16366 ( .A(n18966), .ZN(n15123) );
  NAND2_X1 U16367 ( .A1(n13135), .A2(n15123), .ZN(n13105) );
  NAND2_X1 U16368 ( .A1(n13101), .A2(n13105), .ZN(P2_U2965) );
  AOI22_X1 U16369 ( .A1(P2_EAX_REG_27__SCAN_IN), .A2(n13788), .B1(n13137), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13103) );
  AOI22_X1 U16370 ( .A1(n13852), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n13129), .ZN(n18971) );
  INV_X1 U16371 ( .A(n18971), .ZN(n13102) );
  NAND2_X1 U16372 ( .A1(n13135), .A2(n13102), .ZN(n13118) );
  NAND2_X1 U16373 ( .A1(n13103), .A2(n13118), .ZN(P2_U2963) );
  AOI22_X1 U16374 ( .A1(P2_EAX_REG_18__SCAN_IN), .A2(n13788), .B1(n13137), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13104) );
  AOI22_X1 U16375 ( .A1(n13852), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13850), .ZN(n19104) );
  INV_X1 U16376 ( .A(n19104), .ZN(n15198) );
  NAND2_X1 U16377 ( .A1(n13135), .A2(n15198), .ZN(n13120) );
  NAND2_X1 U16378 ( .A1(n13104), .A2(n13120), .ZN(P2_U2954) );
  AOI22_X1 U16379 ( .A1(P2_EAX_REG_13__SCAN_IN), .A2(n13788), .B1(n13137), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13106) );
  NAND2_X1 U16380 ( .A1(n13106), .A2(n13105), .ZN(P2_U2980) );
  AOI22_X1 U16381 ( .A1(P2_EAX_REG_20__SCAN_IN), .A2(n13788), .B1(n13137), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13107) );
  AOI22_X1 U16382 ( .A1(n13852), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n13850), .ZN(n19115) );
  INV_X1 U16383 ( .A(n19115), .ZN(n15188) );
  NAND2_X1 U16384 ( .A1(n13135), .A2(n15188), .ZN(n13124) );
  NAND2_X1 U16385 ( .A1(n13107), .A2(n13124), .ZN(P2_U2956) );
  AOI22_X1 U16386 ( .A1(n13788), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n13137), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13109) );
  NAND2_X1 U16387 ( .A1(n13109), .A2(n13108), .ZN(P2_U2961) );
  AOI22_X1 U16388 ( .A1(n13788), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n13137), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13110) );
  OAI22_X1 U16389 ( .A1(n13850), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13852), .ZN(n19110) );
  INV_X1 U16390 ( .A(n19110), .ZN(n16234) );
  NAND2_X1 U16391 ( .A1(n13135), .A2(n16234), .ZN(n13122) );
  NAND2_X1 U16392 ( .A1(n13110), .A2(n13122), .ZN(P2_U2955) );
  AOI22_X1 U16393 ( .A1(n13788), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13137), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13112) );
  NAND2_X1 U16394 ( .A1(n13112), .A2(n13111), .ZN(P2_U2959) );
  AOI22_X1 U16395 ( .A1(n13788), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13137), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13113) );
  AOI22_X1 U16396 ( .A1(n13852), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13850), .ZN(n19098) );
  INV_X1 U16397 ( .A(n19098), .ZN(n19011) );
  NAND2_X1 U16398 ( .A1(n13135), .A2(n19011), .ZN(n13116) );
  NAND2_X1 U16399 ( .A1(n13113), .A2(n13116), .ZN(P2_U2953) );
  AOI22_X1 U16400 ( .A1(n13788), .A2(P2_EAX_REG_0__SCAN_IN), .B1(n13137), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n13115) );
  NAND2_X1 U16401 ( .A1(n13115), .A2(n13114), .ZN(P2_U2967) );
  AOI22_X1 U16402 ( .A1(n13788), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n13137), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n13117) );
  NAND2_X1 U16403 ( .A1(n13117), .A2(n13116), .ZN(P2_U2968) );
  AOI22_X1 U16404 ( .A1(n13788), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n13137), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13119) );
  NAND2_X1 U16405 ( .A1(n13119), .A2(n13118), .ZN(P2_U2978) );
  AOI22_X1 U16406 ( .A1(n13788), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13137), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n13121) );
  NAND2_X1 U16407 ( .A1(n13121), .A2(n13120), .ZN(P2_U2969) );
  AOI22_X1 U16408 ( .A1(n13788), .A2(P2_EAX_REG_3__SCAN_IN), .B1(n13137), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n13123) );
  NAND2_X1 U16409 ( .A1(n13123), .A2(n13122), .ZN(P2_U2970) );
  AOI22_X1 U16410 ( .A1(n13788), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13137), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n13125) );
  NAND2_X1 U16411 ( .A1(n13125), .A2(n13124), .ZN(P2_U2971) );
  AOI22_X1 U16412 ( .A1(n13788), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13137), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13126) );
  INV_X1 U16413 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16431) );
  OAI22_X1 U16414 ( .A1(n13129), .A2(n16431), .B1(n18190), .B2(n13852), .ZN(
        n18984) );
  NAND2_X1 U16415 ( .A1(n13135), .A2(n18984), .ZN(n13127) );
  NAND2_X1 U16416 ( .A1(n13126), .A2(n13127), .ZN(P2_U2957) );
  AOI22_X1 U16417 ( .A1(n13788), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n13137), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n13128) );
  NAND2_X1 U16418 ( .A1(n13128), .A2(n13127), .ZN(P2_U2972) );
  AOI22_X1 U16419 ( .A1(n13852), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13129), .ZN(n18960) );
  AOI22_X1 U16420 ( .A1(P2_EAX_REG_15__SCAN_IN), .A2(n13788), .B1(n13137), 
        .B2(P2_LWORD_REG_15__SCAN_IN), .ZN(n13130) );
  OAI21_X1 U16421 ( .B1(n18960), .B2(n13131), .A(n13130), .ZN(P2_U2982) );
  INV_X1 U16422 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19039) );
  INV_X1 U16423 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16425) );
  INV_X1 U16424 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17440) );
  AOI22_X1 U16425 ( .A1(n13852), .A2(n16425), .B1(n17440), .B2(n13850), .ZN(
        n18978) );
  NAND2_X1 U16426 ( .A1(n13135), .A2(n18978), .ZN(n13134) );
  NAND2_X1 U16427 ( .A1(n13137), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13132) );
  OAI211_X1 U16428 ( .C1(n13140), .C2(n19039), .A(n13134), .B(n13132), .ZN(
        P2_U2975) );
  INV_X1 U16429 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13186) );
  NAND2_X1 U16430 ( .A1(n13137), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13133) );
  OAI211_X1 U16431 ( .C1(n13140), .C2(n13186), .A(n13134), .B(n13133), .ZN(
        P2_U2960) );
  INV_X1 U16432 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19027) );
  NAND2_X1 U16433 ( .A1(n13135), .A2(n18963), .ZN(n13139) );
  NAND2_X1 U16434 ( .A1(n13137), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13136) );
  OAI211_X1 U16435 ( .C1(n13140), .C2(n19027), .A(n13139), .B(n13136), .ZN(
        P2_U2981) );
  INV_X1 U16436 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13183) );
  NAND2_X1 U16437 ( .A1(n13137), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13138) );
  OAI211_X1 U16438 ( .C1(n13140), .C2(n13183), .A(n13139), .B(n13138), .ZN(
        P2_U2966) );
  XNOR2_X1 U16439 ( .A(n13384), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13141) );
  XNOR2_X1 U16440 ( .A(n14121), .B(n13141), .ZN(n13350) );
  OAI21_X1 U16441 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13143), .A(
        n13142), .ZN(n13144) );
  INV_X1 U16442 ( .A(n13144), .ZN(n13351) );
  NAND2_X1 U16443 ( .A1(n18939), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13329) );
  OAI21_X1 U16444 ( .B1(n19067), .B2(n13145), .A(n13329), .ZN(n13146) );
  AOI21_X1 U16445 ( .B1(n13351), .B2(n16251), .A(n13146), .ZN(n13147) );
  OAI21_X1 U16446 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16262), .A(
        n13147), .ZN(n13148) );
  AOI21_X1 U16447 ( .B1(n16250), .B2(n13350), .A(n13148), .ZN(n13149) );
  OAI21_X1 U16448 ( .B1(n13728), .B2(n16272), .A(n13149), .ZN(P2_U3013) );
  OAI21_X1 U16449 ( .B1(n13152), .B2(n13151), .A(n13150), .ZN(n13452) );
  AOI21_X1 U16450 ( .B1(n13976), .B2(n13145), .A(n13153), .ZN(n13974) );
  OAI22_X1 U16451 ( .A1(n13976), .A2(n19067), .B1(n19652), .B2(n18925), .ZN(
        n13154) );
  AOI21_X1 U16452 ( .B1(n19059), .B2(n13974), .A(n13154), .ZN(n13159) );
  NOR2_X1 U16453 ( .A1(n13156), .A2(n13155), .ZN(n13444) );
  INV_X1 U16454 ( .A(n13444), .ZN(n13157) );
  NAND3_X1 U16455 ( .A1(n13157), .A2(n16250), .A3(n13443), .ZN(n13158) );
  OAI211_X1 U16456 ( .C1(n13452), .C2(n19075), .A(n13159), .B(n13158), .ZN(
        n13160) );
  AOI21_X1 U16457 ( .B1(n12146), .B2(n19078), .A(n13160), .ZN(n13161) );
  INV_X1 U16458 ( .A(n13161), .ZN(P2_U3012) );
  AND2_X1 U16459 ( .A1(n12899), .A2(n13167), .ZN(n13176) );
  INV_X1 U16460 ( .A(n13599), .ZN(n13557) );
  OAI22_X1 U16461 ( .A1(n13176), .A2(n13029), .B1(n13627), .B2(n13557), .ZN(
        n19781) );
  NAND3_X1 U16462 ( .A1(n13285), .A2(n13163), .A3(n15859), .ZN(n13162) );
  AND2_X1 U16463 ( .A1(n13162), .A2(n20669), .ZN(n20670) );
  OR2_X1 U16464 ( .A1(n19781), .A2(n20670), .ZN(n15829) );
  NAND2_X1 U16465 ( .A1(n15829), .A2(n14301), .ZN(n19787) );
  INV_X1 U16466 ( .A(n19787), .ZN(n13175) );
  INV_X1 U16467 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13174) );
  NAND2_X1 U16468 ( .A1(n13563), .A2(n13557), .ZN(n13171) );
  AND2_X1 U16469 ( .A1(n13163), .A2(n11368), .ZN(n13165) );
  OAI22_X1 U16470 ( .A1(n13166), .A2(n13165), .B1(n20024), .B2(n13164), .ZN(
        n13169) );
  INV_X1 U16471 ( .A(n13167), .ZN(n13168) );
  AOI22_X1 U16472 ( .A1(n13169), .A2(n13599), .B1(n12899), .B2(n13168), .ZN(
        n13170) );
  NAND2_X1 U16473 ( .A1(n13171), .A2(n13170), .ZN(n13172) );
  NAND2_X1 U16474 ( .A1(n13172), .A2(n13290), .ZN(n15826) );
  OR2_X1 U16475 ( .A1(n19787), .A2(n15826), .ZN(n13173) );
  OAI21_X1 U16476 ( .B1(n13175), .B2(n13174), .A(n13173), .ZN(P1_U3484) );
  INV_X1 U16477 ( .A(n20646), .ZN(n20503) );
  NAND2_X1 U16478 ( .A1(n20503), .A2(n20555), .ZN(n19783) );
  INV_X1 U16479 ( .A(n19783), .ZN(n14134) );
  NOR2_X1 U16480 ( .A1(n14134), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n13178)
         );
  NAND2_X1 U16481 ( .A1(n13176), .A2(n14301), .ZN(n14324) );
  OAI21_X1 U16482 ( .B1(n12921), .B2(n13627), .A(n20667), .ZN(n13177) );
  OAI21_X1 U16483 ( .B1(n13178), .B2(n20667), .A(n13177), .ZN(P1_U3487) );
  INV_X1 U16484 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13180) );
  AOI22_X1 U16485 ( .A1(n19757), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13179) );
  OAI21_X1 U16486 ( .B1(n13180), .B2(n13368), .A(n13179), .ZN(P2_U2923) );
  INV_X1 U16487 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n15155) );
  AOI22_X1 U16488 ( .A1(n19757), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13181) );
  OAI21_X1 U16489 ( .B1(n15155), .B2(n13368), .A(n13181), .ZN(P2_U2926) );
  AOI22_X1 U16490 ( .A1(n19757), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13182) );
  OAI21_X1 U16491 ( .B1(n13183), .B2(n13368), .A(n13182), .ZN(P2_U2921) );
  INV_X1 U16492 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n15141) );
  AOI22_X1 U16493 ( .A1(n19757), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13184) );
  OAI21_X1 U16494 ( .B1(n15141), .B2(n13368), .A(n13184), .ZN(P2_U2924) );
  AOI22_X1 U16495 ( .A1(n19757), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13185) );
  OAI21_X1 U16496 ( .B1(n13186), .B2(n13368), .A(n13185), .ZN(P2_U2927) );
  INV_X1 U16497 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13188) );
  AOI22_X1 U16498 ( .A1(n19757), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13187) );
  OAI21_X1 U16499 ( .B1(n13188), .B2(n13368), .A(n13187), .ZN(P2_U2922) );
  INV_X1 U16500 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13190) );
  AOI22_X1 U16501 ( .A1(n19757), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13189) );
  OAI21_X1 U16502 ( .B1(n13190), .B2(n13368), .A(n13189), .ZN(P2_U2925) );
  NAND2_X1 U16503 ( .A1(n12655), .A2(n13195), .ZN(n13706) );
  NAND2_X1 U16504 ( .A1(n12659), .A2(n13196), .ZN(n13700) );
  INV_X1 U16505 ( .A(n13700), .ZN(n13197) );
  OAI21_X2 U16506 ( .B1(n13218), .B2(n13197), .A(n13318), .ZN(n13198) );
  MUX2_X1 U16507 ( .A(n14115), .B(n13728), .S(n15110), .Z(n13199) );
  OAI21_X1 U16508 ( .B1(n19732), .B2(n15114), .A(n13199), .ZN(P2_U2886) );
  NAND2_X1 U16509 ( .A1(n19737), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n18830) );
  NOR2_X1 U16510 ( .A1(n10550), .A2(n18830), .ZN(n13200) );
  OAI21_X1 U16511 ( .B1(n12687), .B2(n19097), .A(n13200), .ZN(n13201) );
  INV_X1 U16512 ( .A(n13201), .ZN(n13202) );
  MUX2_X1 U16513 ( .A(n9815), .B(n10574), .S(n13198), .Z(n13203) );
  OAI21_X1 U16514 ( .B1(n19739), .B2(n15114), .A(n13203), .ZN(P2_U2887) );
  INV_X1 U16515 ( .A(n9616), .ZN(n13224) );
  NAND2_X1 U16516 ( .A1(n13224), .A2(n13779), .ZN(n13221) );
  OAI21_X1 U16517 ( .B1(n13204), .B2(n10529), .A(n19103), .ZN(n13207) );
  NOR2_X1 U16518 ( .A1(n13205), .A2(n10548), .ZN(n13206) );
  AOI21_X1 U16519 ( .B1(n9616), .B2(n13207), .A(n13206), .ZN(n13216) );
  INV_X1 U16520 ( .A(n13779), .ZN(n13747) );
  NOR2_X1 U16521 ( .A1(n13208), .A2(n13747), .ZN(n13213) );
  NOR2_X1 U16522 ( .A1(n12685), .A2(n19109), .ZN(n13211) );
  NAND2_X1 U16523 ( .A1(n12687), .A2(n10548), .ZN(n13209) );
  NAND2_X1 U16524 ( .A1(n13209), .A2(n19765), .ZN(n13210) );
  INV_X1 U16525 ( .A(n19103), .ZN(n13307) );
  AOI21_X1 U16526 ( .B1(n13211), .B2(n13210), .A(n13307), .ZN(n13212) );
  AOI21_X1 U16527 ( .B1(n13213), .B2(n13687), .A(n13212), .ZN(n13215) );
  NAND2_X1 U16528 ( .A1(n13205), .A2(n9622), .ZN(n13214) );
  NAND2_X1 U16529 ( .A1(n13214), .A2(n10559), .ZN(n13332) );
  INV_X1 U16530 ( .A(n13312), .ZN(n13217) );
  NOR2_X1 U16531 ( .A1(n13218), .A2(n13217), .ZN(n13219) );
  OAI211_X1 U16532 ( .C1(n13221), .C2(n13317), .A(n13220), .B(n13219), .ZN(
        n13722) );
  INV_X1 U16533 ( .A(n13722), .ZN(n13746) );
  NAND2_X1 U16534 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19742), .ZN(n15874) );
  OAI22_X1 U16535 ( .A1(n13746), .A2(n18832), .B1(n18835), .B2(n15874), .ZN(
        n13222) );
  INV_X1 U16536 ( .A(n15768), .ZN(n14027) );
  NAND2_X1 U16537 ( .A1(n13224), .A2(n13223), .ZN(n13690) );
  OR4_X1 U16538 ( .A1(n15768), .A2(n19708), .A3(n10753), .A4(n13690), .ZN(
        n13225) );
  OAI21_X1 U16539 ( .B1(n14027), .B2(n13226), .A(n13225), .ZN(P2_U3595) );
  INV_X1 U16540 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13231) );
  INV_X1 U16541 ( .A(n15859), .ZN(n13552) );
  NAND2_X1 U16542 ( .A1(n14877), .A2(n13552), .ZN(n13228) );
  NAND2_X1 U16543 ( .A1(n13228), .A2(n15840), .ZN(n13229) );
  NAND2_X1 U16544 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16170) );
  NAND2_X1 U16545 ( .A1(n20556), .A2(n16168), .ZN(n19901) );
  NOR2_X4 U16546 ( .A1(n19903), .A2(n19930), .ZN(n19929) );
  AOI22_X1 U16547 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13230) );
  OAI21_X1 U16548 ( .B1(n13231), .B2(n13436), .A(n13230), .ZN(P1_U2907) );
  AOI22_X1 U16549 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13232) );
  OAI21_X1 U16550 ( .B1(n11904), .B2(n13436), .A(n13232), .ZN(P1_U2912) );
  INV_X1 U16551 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13234) );
  AOI22_X1 U16552 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13233) );
  OAI21_X1 U16553 ( .B1(n13234), .B2(n13436), .A(n13233), .ZN(P1_U2908) );
  INV_X1 U16554 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13236) );
  AOI22_X1 U16555 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13235) );
  OAI21_X1 U16556 ( .B1(n13236), .B2(n13436), .A(n13235), .ZN(P1_U2910) );
  INV_X1 U16557 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13396) );
  AOI22_X1 U16558 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13237) );
  OAI21_X1 U16559 ( .B1(n13396), .B2(n13436), .A(n13237), .ZN(P1_U2911) );
  INV_X1 U16560 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13239) );
  AOI22_X1 U16561 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13238) );
  OAI21_X1 U16562 ( .B1(n13239), .B2(n13436), .A(n13238), .ZN(P1_U2906) );
  INV_X1 U16563 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n20808) );
  AOI22_X1 U16564 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13240) );
  OAI21_X1 U16565 ( .B1(n20808), .B2(n13436), .A(n13240), .ZN(P1_U2909) );
  OR2_X1 U16566 ( .A1(n13243), .A2(n13242), .ZN(n13244) );
  NAND2_X1 U16567 ( .A1(n13241), .A2(n13244), .ZN(n18997) );
  NOR2_X1 U16568 ( .A1(n13246), .A2(n13245), .ZN(n13247) );
  OR2_X1 U16569 ( .A1(n13251), .A2(n13247), .ZN(n13887) );
  NOR2_X1 U16570 ( .A1(n13887), .A2(n13198), .ZN(n13248) );
  AOI21_X1 U16571 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n15122), .A(n13248), .ZN(
        n13249) );
  OAI21_X1 U16572 ( .B1(n18997), .B2(n15114), .A(n13249), .ZN(P2_U2883) );
  XOR2_X1 U16573 ( .A(n13241), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13256)
         );
  OR2_X1 U16574 ( .A1(n13251), .A2(n13250), .ZN(n13253) );
  NAND2_X1 U16575 ( .A1(n13253), .A2(n13252), .ZN(n18945) );
  NOR2_X1 U16576 ( .A1(n18945), .A2(n13198), .ZN(n13254) );
  AOI21_X1 U16577 ( .B1(P2_EBX_REG_5__SCAN_IN), .B2(n13198), .A(n13254), .ZN(
        n13255) );
  OAI21_X1 U16578 ( .B1(n13256), .B2(n15114), .A(n13255), .ZN(P2_U2882) );
  MUX2_X1 U16579 ( .A(P2_EBX_REG_2__SCAN_IN), .B(n10647), .S(n15110), .Z(
        n13259) );
  INV_X1 U16580 ( .A(n13259), .ZN(n13260) );
  OAI21_X1 U16581 ( .B1(n19721), .B2(n15114), .A(n13260), .ZN(P2_U2885) );
  NAND3_X1 U16582 ( .A1(n20556), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16162) );
  INV_X1 U16583 ( .A(n16162), .ZN(n13263) );
  NAND2_X1 U16584 ( .A1(n20646), .A2(n13266), .ZN(n20668) );
  AND2_X1 U16585 ( .A1(n20668), .A2(n20556), .ZN(n13267) );
  NAND2_X1 U16586 ( .A1(n20556), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15837) );
  NAND2_X1 U16587 ( .A1(n20640), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13268) );
  NAND2_X1 U16588 ( .A1(n15837), .A2(n13268), .ZN(n13300) );
  INV_X1 U16589 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13652) );
  INV_X1 U16590 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n13655) );
  OAI22_X1 U16591 ( .A1(n14723), .A2(n13652), .B1(n16122), .B2(n13655), .ZN(
        n13269) );
  AOI21_X1 U16592 ( .B1(n16032), .B2(n13652), .A(n13269), .ZN(n13272) );
  OR2_X1 U16593 ( .A1(n13270), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20006) );
  NAND3_X1 U16594 ( .A1(n20006), .A2(n20005), .A3(n19968), .ZN(n13271) );
  OAI211_X1 U16595 ( .C1(n13654), .C2(n20022), .A(n13272), .B(n13271), .ZN(
        P1_U2998) );
  OR2_X1 U16596 ( .A1(n12943), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13274) );
  AND2_X1 U16597 ( .A1(n13274), .A2(n13273), .ZN(n13634) );
  INV_X1 U16598 ( .A(n13634), .ZN(n13283) );
  NAND2_X1 U16599 ( .A1(n13563), .A2(n13599), .ZN(n13548) );
  INV_X1 U16600 ( .A(n13275), .ZN(n13276) );
  NAND2_X1 U16601 ( .A1(n13276), .A2(n13630), .ZN(n13277) );
  NAND2_X1 U16602 ( .A1(n13548), .A2(n13277), .ZN(n13278) );
  INV_X1 U16603 ( .A(n13279), .ZN(n13282) );
  OAI21_X1 U16604 ( .B1(n13282), .B2(n13281), .A(n13280), .ZN(n13645) );
  NAND2_X2 U16605 ( .A1(n19899), .A2(n13290), .ZN(n14515) );
  OAI222_X1 U16606 ( .A1(n13283), .A2(n14532), .B1(n12926), .B2(n19899), .C1(
        n13645), .C2(n14515), .ZN(P1_U2872) );
  INV_X1 U16607 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13289) );
  INV_X1 U16608 ( .A(n13284), .ZN(n13286) );
  NAND2_X1 U16609 ( .A1(n13286), .A2(n13285), .ZN(n13287) );
  AND2_X1 U16610 ( .A1(n13288), .A2(n13287), .ZN(n20018) );
  OAI222_X1 U16611 ( .A1(n14515), .A2(n13654), .B1(n19899), .B2(n13289), .C1(
        n14532), .C2(n20018), .ZN(P1_U2871) );
  NAND2_X1 U16612 ( .A1(n11380), .A2(n13290), .ZN(n13291) );
  INV_X1 U16613 ( .A(n13291), .ZN(n13292) );
  NAND2_X1 U16614 ( .A1(n20021), .A2(DATAI_1_), .ZN(n13294) );
  NAND2_X1 U16615 ( .A1(n20020), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13293) );
  AND2_X1 U16616 ( .A1(n13294), .A2(n13293), .ZN(n20034) );
  INV_X1 U16617 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n19928) );
  OAI222_X1 U16618 ( .A1(n13654), .A2(n15997), .B1(n14573), .B2(n20034), .C1(
        n14571), .C2(n19928), .ZN(P1_U2903) );
  OR2_X1 U16619 ( .A1(n19934), .A2(n11367), .ZN(n13466) );
  INV_X1 U16620 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14570) );
  OR2_X1 U16621 ( .A1(n19934), .A2(n11366), .ZN(n13394) );
  INV_X1 U16622 ( .A(DATAI_15_), .ZN(n13297) );
  INV_X1 U16623 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13296) );
  MUX2_X1 U16624 ( .A(n13297), .B(n13296), .S(n20020), .Z(n14572) );
  INV_X1 U16625 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n19902) );
  OAI222_X1 U16626 ( .A1(n13466), .A2(n14570), .B1(n13394), .B2(n14572), .C1(
        n13481), .C2(n19902), .ZN(P1_U2967) );
  OAI21_X1 U16627 ( .B1(n13299), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13298), .ZN(n13409) );
  NAND2_X1 U16628 ( .A1(n20014), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13398) );
  OAI21_X1 U16629 ( .B1(n19962), .B2(n13300), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13301) );
  OAI211_X1 U16630 ( .C1(n13409), .C2(n16035), .A(n13398), .B(n13301), .ZN(
        n13302) );
  INV_X1 U16631 ( .A(n13302), .ZN(n13303) );
  OAI21_X1 U16632 ( .B1(n20022), .B2(n13645), .A(n13303), .ZN(P1_U2999) );
  NAND2_X1 U16633 ( .A1(n13307), .A2(n13779), .ZN(n13316) );
  AOI21_X1 U16634 ( .B1(n13304), .B2(n19765), .A(n10529), .ZN(n13314) );
  NAND2_X1 U16635 ( .A1(n13305), .A2(n10753), .ZN(n13310) );
  MUX2_X1 U16636 ( .A(n13307), .B(n13306), .S(n10753), .Z(n13308) );
  NAND3_X1 U16637 ( .A1(n13308), .A2(n13687), .A3(n19756), .ZN(n13309) );
  NAND4_X1 U16638 ( .A1(n13312), .A2(n13311), .A3(n13310), .A4(n13309), .ZN(
        n13313) );
  AOI21_X1 U16639 ( .B1(n13317), .B2(n13314), .A(n13313), .ZN(n13315) );
  OAI21_X1 U16640 ( .B1(n13317), .B2(n13316), .A(n13315), .ZN(n13319) );
  NAND2_X1 U16641 ( .A1(n13319), .A2(n13318), .ZN(n13348) );
  NAND2_X1 U16642 ( .A1(n13320), .A2(n12687), .ZN(n13322) );
  NAND2_X1 U16643 ( .A1(n13322), .A2(n9617), .ZN(n13323) );
  XNOR2_X1 U16644 ( .A(n13324), .B(n13325), .ZN(n19727) );
  NAND2_X1 U16645 ( .A1(n13685), .A2(n10753), .ZN(n13326) );
  NAND2_X1 U16646 ( .A1(n13326), .A2(n13706), .ZN(n13327) );
  INV_X1 U16647 ( .A(n13328), .ZN(n16290) );
  NAND2_X1 U16648 ( .A1(n13348), .A2(n16290), .ZN(n13826) );
  OAI21_X1 U16649 ( .B1(n13826), .B2(n14067), .A(n13329), .ZN(n13347) );
  NAND2_X1 U16650 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13822) );
  INV_X1 U16651 ( .A(n13822), .ZN(n13821) );
  NAND2_X1 U16652 ( .A1(n13344), .A2(n13705), .ZN(n13831) );
  AND2_X1 U16653 ( .A1(n10572), .A2(n13330), .ZN(n13342) );
  NAND2_X1 U16654 ( .A1(n13331), .A2(n10753), .ZN(n13723) );
  NAND2_X1 U16655 ( .A1(n13723), .A2(n13332), .ZN(n13333) );
  NAND2_X1 U16656 ( .A1(n13333), .A2(n10553), .ZN(n13340) );
  OAI22_X1 U16657 ( .A1(n13334), .A2(n12658), .B1(n19103), .B2(n19765), .ZN(
        n13335) );
  INV_X1 U16658 ( .A(n13335), .ZN(n13337) );
  AND3_X1 U16659 ( .A1(n13338), .A2(n13337), .A3(n13336), .ZN(n13339) );
  NAND2_X1 U16660 ( .A1(n13340), .A2(n13339), .ZN(n13341) );
  AOI21_X1 U16661 ( .B1(n13342), .B2(n10571), .A(n13341), .ZN(n13727) );
  NAND2_X1 U16662 ( .A1(n13727), .A2(n13700), .ZN(n13343) );
  NAND2_X1 U16663 ( .A1(n13344), .A2(n13343), .ZN(n15659) );
  INV_X1 U16664 ( .A(n15611), .ZN(n15660) );
  AOI211_X1 U16665 ( .C1(n14067), .C2(n13345), .A(n13821), .B(n15660), .ZN(
        n13346) );
  AOI211_X1 U16666 ( .C1(n19727), .C2(n15739), .A(n13347), .B(n13346), .ZN(
        n13353) );
  AOI22_X1 U16667 ( .A1(n16282), .A2(n13351), .B1(n16281), .B2(n13350), .ZN(
        n13352) );
  OAI211_X1 U16668 ( .C1(n13728), .C2(n16315), .A(n13353), .B(n13352), .ZN(
        P2_U3045) );
  INV_X1 U16669 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13355) );
  AOI22_X1 U16670 ( .A1(n19757), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13354) );
  OAI21_X1 U16671 ( .B1(n13355), .B2(n13368), .A(n13354), .ZN(P2_U2931) );
  INV_X1 U16672 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15181) );
  AOI22_X1 U16673 ( .A1(n19757), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13356) );
  OAI21_X1 U16674 ( .B1(n15181), .B2(n13368), .A(n13356), .ZN(P2_U2930) );
  INV_X1 U16675 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13358) );
  AOI22_X1 U16676 ( .A1(n19757), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13357) );
  OAI21_X1 U16677 ( .B1(n13358), .B2(n13368), .A(n13357), .ZN(P2_U2929) );
  INV_X1 U16678 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13360) );
  AOI22_X1 U16679 ( .A1(n19757), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13359) );
  OAI21_X1 U16680 ( .B1(n13360), .B2(n13368), .A(n13359), .ZN(P2_U2928) );
  INV_X1 U16681 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13362) );
  AOI22_X1 U16682 ( .A1(n19757), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13361) );
  OAI21_X1 U16683 ( .B1(n13362), .B2(n13368), .A(n13361), .ZN(P2_U2934) );
  INV_X1 U16684 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13364) );
  AOI22_X1 U16685 ( .A1(n19757), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13363) );
  OAI21_X1 U16686 ( .B1(n13364), .B2(n13368), .A(n13363), .ZN(P2_U2933) );
  INV_X1 U16687 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13366) );
  AOI22_X1 U16688 ( .A1(n19757), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13365) );
  OAI21_X1 U16689 ( .B1(n13366), .B2(n13368), .A(n13365), .ZN(P2_U2935) );
  INV_X1 U16690 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13369) );
  AOI22_X1 U16691 ( .A1(n19757), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13367) );
  OAI21_X1 U16692 ( .B1(n13369), .B2(n13368), .A(n13367), .ZN(P2_U2932) );
  NOR2_X1 U16693 ( .A1(n13241), .A2(n13370), .ZN(n13372) );
  OAI211_X1 U16694 ( .C1(n13372), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15119), .B(n13371), .ZN(n13376) );
  AOI21_X1 U16695 ( .B1(n13374), .B2(n13252), .A(n13373), .ZN(n14099) );
  NAND2_X1 U16696 ( .A1(n15110), .A2(n14099), .ZN(n13375) );
  OAI211_X1 U16697 ( .C1(n15110), .C2(n13967), .A(n13376), .B(n13375), .ZN(
        P2_U2881) );
  NOR2_X1 U16698 ( .A1(n13378), .A2(n13377), .ZN(n13379) );
  NOR2_X1 U16699 ( .A1(n13380), .A2(n13379), .ZN(n19019) );
  INV_X1 U16700 ( .A(n19019), .ZN(n14078) );
  NAND2_X1 U16701 ( .A1(n13328), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n19073) );
  OAI21_X1 U16702 ( .B1(n16305), .B2(n14078), .A(n19073), .ZN(n13386) );
  INV_X1 U16703 ( .A(n13381), .ZN(n13382) );
  OAI21_X1 U16704 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13383), .A(
        n13382), .ZN(n19074) );
  OAI21_X1 U16705 ( .B1(n14076), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13384), .ZN(n19071) );
  OAI22_X1 U16706 ( .A1(n16308), .A2(n19074), .B1(n16306), .B2(n19071), .ZN(
        n13385) );
  AOI211_X1 U16707 ( .C1(n19079), .C2(n15757), .A(n13386), .B(n13385), .ZN(
        n13388) );
  MUX2_X1 U16708 ( .A(n15660), .B(n13826), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13387) );
  NAND2_X1 U16709 ( .A1(n13388), .A2(n13387), .ZN(P2_U3046) );
  XOR2_X1 U16710 ( .A(n13371), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13393)
         );
  OR2_X1 U16711 ( .A1(n13389), .A2(n13373), .ZN(n13390) );
  NAND2_X1 U16712 ( .A1(n13418), .A2(n13390), .ZN(n14172) );
  MUX2_X1 U16713 ( .A(n14172), .B(n13391), .S(n15122), .Z(n13392) );
  OAI21_X1 U16714 ( .B1(n13393), .B2(n15114), .A(n13392), .ZN(P2_U2880) );
  MUX2_X1 U16715 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n20020), .Z(
        n14549) );
  NAND2_X1 U16716 ( .A1(n19944), .A2(n14549), .ZN(n19948) );
  NAND2_X1 U16717 ( .A1(n19934), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n13395) );
  OAI211_X1 U16718 ( .C1(n13466), .C2(n13396), .A(n19948), .B(n13395), .ZN(
        P1_U2946) );
  MUX2_X1 U16719 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n20020), .Z(
        n14579) );
  NAND2_X1 U16720 ( .A1(n19944), .A2(n14579), .ZN(n19952) );
  NAND2_X1 U16721 ( .A1(n19934), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13397) );
  OAI211_X1 U16722 ( .C1(n13466), .C2(n20808), .A(n19952), .B(n13397), .ZN(
        P1_U2948) );
  INV_X1 U16723 ( .A(n13398), .ZN(n13407) );
  INV_X1 U16724 ( .A(n13399), .ZN(n13400) );
  NAND2_X1 U16725 ( .A1(n13400), .A2(n16095), .ZN(n13402) );
  INV_X1 U16726 ( .A(n13402), .ZN(n13405) );
  AOI21_X1 U16727 ( .B1(n14882), .B2(n13402), .A(n13401), .ZN(n20012) );
  INV_X1 U16728 ( .A(n13403), .ZN(n13404) );
  AOI22_X1 U16729 ( .A1(n13405), .A2(n14882), .B1(n20012), .B2(n13404), .ZN(
        n13406) );
  AOI211_X1 U16730 ( .C1(n13634), .C2(n19981), .A(n13407), .B(n13406), .ZN(
        n13408) );
  OAI21_X1 U16731 ( .B1(n13409), .B2(n16126), .A(n13408), .ZN(P1_U3031) );
  INV_X1 U16732 ( .A(n19145), .ZN(n19711) );
  MUX2_X1 U16733 ( .A(P2_EBX_REG_3__SCAN_IN), .B(n13412), .S(n15110), .Z(
        n13413) );
  AOI21_X1 U16734 ( .B1(n19711), .B2(n15119), .A(n13413), .ZN(n13414) );
  INV_X1 U16735 ( .A(n13414), .ZN(P2_U2884) );
  XNOR2_X1 U16736 ( .A(n13415), .B(n13416), .ZN(n13421) );
  NAND2_X1 U16737 ( .A1(n13418), .A2(n13417), .ZN(n13419) );
  NAND2_X1 U16738 ( .A1(n13519), .A2(n13419), .ZN(n15748) );
  MUX2_X1 U16739 ( .A(n15748), .B(n11134), .S(n15122), .Z(n13420) );
  OAI21_X1 U16740 ( .B1(n13421), .B2(n15114), .A(n13420), .ZN(P2_U2879) );
  AOI22_X1 U16741 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13422) );
  OAI21_X1 U16742 ( .B1(n11818), .B2(n13436), .A(n13422), .ZN(P1_U2916) );
  INV_X1 U16743 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13424) );
  AOI22_X1 U16744 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13423) );
  OAI21_X1 U16745 ( .B1(n13424), .B2(n13436), .A(n13423), .ZN(P1_U2918) );
  INV_X1 U16746 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13426) );
  AOI22_X1 U16747 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13425) );
  OAI21_X1 U16748 ( .B1(n13426), .B2(n13436), .A(n13425), .ZN(P1_U2919) );
  INV_X1 U16749 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13428) );
  AOI22_X1 U16750 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13427) );
  OAI21_X1 U16751 ( .B1(n13428), .B2(n13436), .A(n13427), .ZN(P1_U2915) );
  INV_X1 U16752 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13430) );
  AOI22_X1 U16753 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13429) );
  OAI21_X1 U16754 ( .B1(n13430), .B2(n13436), .A(n13429), .ZN(P1_U2913) );
  INV_X1 U16755 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13432) );
  AOI22_X1 U16756 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13431) );
  OAI21_X1 U16757 ( .B1(n13432), .B2(n13436), .A(n13431), .ZN(P1_U2920) );
  INV_X1 U16758 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13434) );
  AOI22_X1 U16759 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13433) );
  OAI21_X1 U16760 ( .B1(n13434), .B2(n13436), .A(n13433), .ZN(P1_U2914) );
  INV_X1 U16761 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13437) );
  AOI22_X1 U16762 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13435) );
  OAI21_X1 U16763 ( .B1(n13437), .B2(n13436), .A(n13435), .ZN(P1_U2917) );
  NAND2_X1 U16764 ( .A1(n13439), .A2(n13438), .ZN(n13442) );
  INV_X1 U16765 ( .A(n13440), .ZN(n13441) );
  NAND2_X1 U16766 ( .A1(n13442), .A2(n13441), .ZN(n19723) );
  INV_X1 U16767 ( .A(n13443), .ZN(n13445) );
  NOR3_X1 U16768 ( .A1(n16306), .A2(n13445), .A3(n13444), .ZN(n13447) );
  OAI22_X1 U16769 ( .A1(n13826), .A2(n13823), .B1(n19652), .B2(n18925), .ZN(
        n13446) );
  AOI211_X1 U16770 ( .C1(n19723), .C2(n15739), .A(n13447), .B(n13446), .ZN(
        n13451) );
  INV_X1 U16771 ( .A(n13831), .ZN(n15655) );
  MUX2_X1 U16772 ( .A(n13821), .B(n13822), .S(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n13448) );
  INV_X1 U16773 ( .A(n13448), .ZN(n13449) );
  INV_X1 U16774 ( .A(n15659), .ZN(n13829) );
  AOI22_X1 U16775 ( .A1(n15655), .A2(n13449), .B1(n13829), .B2(n13448), .ZN(
        n13450) );
  OAI211_X1 U16776 ( .C1(n13452), .C2(n16308), .A(n13451), .B(n13450), .ZN(
        n13453) );
  AOI21_X1 U16777 ( .B1(n10647), .B2(n15757), .A(n13453), .ZN(n13454) );
  INV_X1 U16778 ( .A(n13454), .ZN(P2_U3044) );
  NAND2_X1 U16779 ( .A1(n20021), .A2(DATAI_0_), .ZN(n13456) );
  NAND2_X1 U16780 ( .A1(n20020), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13455) );
  INV_X1 U16781 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n19933) );
  OAI222_X1 U16782 ( .A1(n13645), .A2(n15997), .B1(n14573), .B2(n20027), .C1(
        n14571), .C2(n19933), .ZN(P1_U2904) );
  NAND2_X1 U16783 ( .A1(n13457), .A2(n13459), .ZN(n13664) );
  INV_X1 U16784 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13463) );
  NAND2_X1 U16785 ( .A1(n13461), .A2(n13460), .ZN(n13462) );
  NAND2_X1 U16786 ( .A1(n13535), .A2(n13462), .ZN(n19997) );
  OAI222_X1 U16787 ( .A1(n13664), .A2(n14515), .B1(n19899), .B2(n13463), .C1(
        n19997), .C2(n14532), .ZN(P1_U2870) );
  NAND2_X1 U16788 ( .A1(n20021), .A2(DATAI_2_), .ZN(n13465) );
  NAND2_X1 U16789 ( .A1(n20020), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13464) );
  AND2_X1 U16790 ( .A1(n13465), .A2(n13464), .ZN(n20037) );
  INV_X1 U16791 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n19926) );
  OAI222_X1 U16792 ( .A1(n13664), .A2(n15997), .B1(n14573), .B2(n20037), .C1(
        n14571), .C2(n19926), .ZN(P1_U2902) );
  AOI22_X1 U16793 ( .A1(n19959), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n19934), .ZN(n13467) );
  INV_X1 U16794 ( .A(n20037), .ZN(n16004) );
  NAND2_X1 U16795 ( .A1(n19944), .A2(n16004), .ZN(n13496) );
  NAND2_X1 U16796 ( .A1(n13467), .A2(n13496), .ZN(P1_U2939) );
  AOI22_X1 U16797 ( .A1(n19959), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n19934), .ZN(n13470) );
  NAND2_X1 U16798 ( .A1(n20021), .A2(DATAI_5_), .ZN(n13469) );
  NAND2_X1 U16799 ( .A1(n20020), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13468) );
  AND2_X1 U16800 ( .A1(n13469), .A2(n13468), .ZN(n20049) );
  INV_X1 U16801 ( .A(n20049), .ZN(n15996) );
  NAND2_X1 U16802 ( .A1(n19944), .A2(n15996), .ZN(n13500) );
  NAND2_X1 U16803 ( .A1(n13470), .A2(n13500), .ZN(P1_U2942) );
  AOI22_X1 U16804 ( .A1(n19959), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n19934), .ZN(n13471) );
  INV_X1 U16805 ( .A(n20027), .ZN(n14567) );
  NAND2_X1 U16806 ( .A1(n19944), .A2(n14567), .ZN(n13488) );
  NAND2_X1 U16807 ( .A1(n13471), .A2(n13488), .ZN(P1_U2937) );
  AOI22_X1 U16808 ( .A1(n19959), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n19954), .ZN(n13474) );
  NAND2_X1 U16809 ( .A1(n20021), .A2(DATAI_3_), .ZN(n13473) );
  NAND2_X1 U16810 ( .A1(n20020), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13472) );
  AND2_X1 U16811 ( .A1(n13473), .A2(n13472), .ZN(n20041) );
  INV_X1 U16812 ( .A(n20041), .ZN(n16001) );
  NAND2_X1 U16813 ( .A1(n19944), .A2(n16001), .ZN(n13476) );
  NAND2_X1 U16814 ( .A1(n13474), .A2(n13476), .ZN(P1_U2940) );
  AOI22_X1 U16815 ( .A1(n19959), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n19954), .ZN(n13475) );
  INV_X1 U16816 ( .A(n20034), .ZN(n16009) );
  NAND2_X1 U16817 ( .A1(n19944), .A2(n16009), .ZN(n13492) );
  NAND2_X1 U16818 ( .A1(n13475), .A2(n13492), .ZN(P1_U2938) );
  AOI22_X1 U16819 ( .A1(n19959), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n19954), .ZN(n13477) );
  NAND2_X1 U16820 ( .A1(n13477), .A2(n13476), .ZN(P1_U2955) );
  AOI22_X1 U16821 ( .A1(n19959), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n19954), .ZN(n13480) );
  NAND2_X1 U16822 ( .A1(n20021), .A2(DATAI_4_), .ZN(n13479) );
  NAND2_X1 U16823 ( .A1(n20020), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13478) );
  AND2_X1 U16824 ( .A1(n13479), .A2(n13478), .ZN(n20045) );
  INV_X1 U16825 ( .A(n20045), .ZN(n14563) );
  NAND2_X1 U16826 ( .A1(n19944), .A2(n14563), .ZN(n13498) );
  NAND2_X1 U16827 ( .A1(n13480), .A2(n13498), .ZN(P1_U2941) );
  AOI22_X1 U16828 ( .A1(n19959), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n19954), .ZN(n13484) );
  NAND2_X1 U16829 ( .A1(n20021), .A2(DATAI_6_), .ZN(n13483) );
  NAND2_X1 U16830 ( .A1(n20020), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13482) );
  AND2_X1 U16831 ( .A1(n13483), .A2(n13482), .ZN(n20052) );
  INV_X1 U16832 ( .A(n20052), .ZN(n14559) );
  NAND2_X1 U16833 ( .A1(n19944), .A2(n14559), .ZN(n13490) );
  NAND2_X1 U16834 ( .A1(n13484), .A2(n13490), .ZN(P1_U2943) );
  AOI22_X1 U16835 ( .A1(n19959), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n19954), .ZN(n13487) );
  NAND2_X1 U16836 ( .A1(n20021), .A2(DATAI_7_), .ZN(n13486) );
  NAND2_X1 U16837 ( .A1(n20020), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13485) );
  INV_X1 U16838 ( .A(n20059), .ZN(n14555) );
  NAND2_X1 U16839 ( .A1(n19944), .A2(n14555), .ZN(n13494) );
  NAND2_X1 U16840 ( .A1(n13487), .A2(n13494), .ZN(P1_U2944) );
  AOI22_X1 U16841 ( .A1(n19959), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n19954), .ZN(n13489) );
  NAND2_X1 U16842 ( .A1(n13489), .A2(n13488), .ZN(P1_U2952) );
  AOI22_X1 U16843 ( .A1(n19959), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n19954), .ZN(n13491) );
  NAND2_X1 U16844 ( .A1(n13491), .A2(n13490), .ZN(P1_U2958) );
  AOI22_X1 U16845 ( .A1(n19959), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n19954), .ZN(n13493) );
  NAND2_X1 U16846 ( .A1(n13493), .A2(n13492), .ZN(P1_U2953) );
  AOI22_X1 U16847 ( .A1(n19959), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n19954), .ZN(n13495) );
  NAND2_X1 U16848 ( .A1(n13495), .A2(n13494), .ZN(P1_U2959) );
  AOI22_X1 U16849 ( .A1(n19959), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n19954), .ZN(n13497) );
  NAND2_X1 U16850 ( .A1(n13497), .A2(n13496), .ZN(P1_U2954) );
  AOI22_X1 U16851 ( .A1(n19959), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n19954), .ZN(n13499) );
  NAND2_X1 U16852 ( .A1(n13499), .A2(n13498), .ZN(P1_U2956) );
  AOI22_X1 U16853 ( .A1(n19959), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n19954), .ZN(n13501) );
  NAND2_X1 U16854 ( .A1(n13501), .A2(n13500), .ZN(P1_U2957) );
  AOI21_X1 U16855 ( .B1(n13504), .B2(n13503), .A(n13502), .ZN(n20000) );
  INV_X1 U16856 ( .A(n20000), .ZN(n13509) );
  INV_X1 U16857 ( .A(n13664), .ZN(n13507) );
  AOI22_X1 U16858 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20014), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13505) );
  OAI21_X1 U16859 ( .B1(n19972), .B2(n13660), .A(n13505), .ZN(n13506) );
  AOI21_X1 U16860 ( .B1(n13507), .B2(n14671), .A(n13506), .ZN(n13508) );
  OAI21_X1 U16861 ( .B1(n13509), .B2(n16035), .A(n13508), .ZN(P1_U2997) );
  INV_X1 U16862 ( .A(n19723), .ZN(n18986) );
  XNOR2_X1 U16863 ( .A(n19721), .B(n19723), .ZN(n13513) );
  INV_X1 U16864 ( .A(n19727), .ZN(n13510) );
  NAND2_X1 U16865 ( .A1(n19732), .A2(n13510), .ZN(n13511) );
  XNOR2_X1 U16866 ( .A(n19732), .B(n19727), .ZN(n19009) );
  NAND2_X1 U16867 ( .A1(n19144), .A2(n19019), .ZN(n19018) );
  NAND2_X1 U16868 ( .A1(n19009), .A2(n19018), .ZN(n19008) );
  NAND2_X1 U16869 ( .A1(n13511), .A2(n19008), .ZN(n13512) );
  NAND2_X1 U16870 ( .A1(n13513), .A2(n13512), .ZN(n18987) );
  OAI21_X1 U16871 ( .B1(n13513), .B2(n13512), .A(n18987), .ZN(n13514) );
  NAND2_X1 U16872 ( .A1(n13514), .A2(n19017), .ZN(n13518) );
  INV_X1 U16873 ( .A(n16235), .ZN(n15156) );
  INV_X1 U16874 ( .A(n13515), .ZN(n13516) );
  AOI22_X1 U16875 ( .A1(n19012), .A2(n15198), .B1(n19015), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n13517) );
  OAI211_X1 U16876 ( .C1(n18986), .C2(n15206), .A(n13518), .B(n13517), .ZN(
        P2_U2917) );
  INV_X1 U16877 ( .A(n13520), .ZN(n13521) );
  OAI21_X1 U16878 ( .B1(n11136), .B2(n13521), .A(n13526), .ZN(n18928) );
  OAI211_X1 U16879 ( .C1(n9728), .C2(n9655), .A(n15119), .B(n9654), .ZN(n13523) );
  NAND2_X1 U16880 ( .A1(n15122), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n13522) );
  OAI211_X1 U16881 ( .C1(n15122), .C2(n18928), .A(n13523), .B(n13522), .ZN(
        P2_U2878) );
  XNOR2_X1 U16882 ( .A(n9654), .B(n13524), .ZN(n13531) );
  AND2_X1 U16883 ( .A1(n13526), .A2(n13525), .ZN(n13527) );
  NOR2_X1 U16884 ( .A1(n13672), .A2(n13527), .ZN(n16258) );
  NOR2_X1 U16885 ( .A1(n15110), .A2(n13528), .ZN(n13529) );
  AOI21_X1 U16886 ( .B1(n16258), .B2(n15110), .A(n13529), .ZN(n13530) );
  OAI21_X1 U16887 ( .B1(n13531), .B2(n15114), .A(n13530), .ZN(P2_U2877) );
  INV_X1 U16888 ( .A(n13533), .ZN(n13534) );
  XNOR2_X1 U16889 ( .A(n13532), .B(n13534), .ZN(n13755) );
  INV_X1 U16890 ( .A(n13755), .ZN(n13606) );
  AOI21_X1 U16891 ( .B1(n13536), .B2(n13535), .A(n13615), .ZN(n19980) );
  AOI22_X1 U16892 ( .A1(n19980), .A2(n19894), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14510), .ZN(n13537) );
  OAI21_X1 U16893 ( .B1(n13606), .B2(n14515), .A(n13537), .ZN(P1_U2869) );
  OAI21_X1 U16894 ( .B1(n13540), .B2(n13539), .A(n13538), .ZN(n19982) );
  AOI22_X1 U16895 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20014), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n13541) );
  OAI21_X1 U16896 ( .B1(n19972), .B2(n13767), .A(n13541), .ZN(n13542) );
  AOI21_X1 U16897 ( .B1(n13755), .B2(n14671), .A(n13542), .ZN(n13543) );
  OAI21_X1 U16898 ( .B1(n19982), .B2(n16035), .A(n13543), .ZN(P1_U2996) );
  NOR2_X1 U16899 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20555), .ZN(n13595) );
  NAND2_X1 U16900 ( .A1(n20024), .A2(n11367), .ZN(n13635) );
  OR2_X1 U16901 ( .A1(n13635), .A2(n13544), .ZN(n13545) );
  AND4_X1 U16902 ( .A1(n13548), .A2(n13547), .A3(n13546), .A4(n13545), .ZN(
        n13560) );
  NAND2_X1 U16903 ( .A1(n14877), .A2(n20669), .ZN(n13551) );
  INV_X1 U16904 ( .A(n13549), .ZN(n13550) );
  NAND2_X1 U16905 ( .A1(n13551), .A2(n13550), .ZN(n13553) );
  NAND2_X1 U16906 ( .A1(n13553), .A2(n13552), .ZN(n13556) );
  INV_X1 U16907 ( .A(n13554), .ZN(n13555) );
  NAND2_X1 U16908 ( .A1(n13556), .A2(n13555), .ZN(n13558) );
  NAND2_X1 U16909 ( .A1(n13558), .A2(n13557), .ZN(n13559) );
  INV_X1 U16910 ( .A(n13561), .ZN(n13562) );
  OR2_X1 U16911 ( .A1(n13563), .A2(n13562), .ZN(n13578) );
  XNOR2_X1 U16912 ( .A(n13564), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14887) );
  INV_X1 U16913 ( .A(n14877), .ZN(n15813) );
  XNOR2_X1 U16914 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13567) );
  INV_X1 U16915 ( .A(n13565), .ZN(n13566) );
  NAND2_X1 U16916 ( .A1(n13566), .A2(n14875), .ZN(n13581) );
  OAI22_X1 U16917 ( .A1(n15813), .A2(n13567), .B1(n13581), .B2(n14887), .ZN(
        n13573) );
  INV_X1 U16918 ( .A(n13569), .ZN(n13571) );
  NAND4_X1 U16919 ( .A1(n13571), .A2(n12070), .A3(n12048), .A4(n13570), .ZN(
        n13587) );
  INV_X1 U16920 ( .A(n13587), .ZN(n14879) );
  NOR2_X1 U16921 ( .A1(n13568), .A2(n14879), .ZN(n13572) );
  AOI211_X1 U16922 ( .C1(n13578), .C2(n14887), .A(n13573), .B(n13572), .ZN(
        n14893) );
  NAND2_X1 U16923 ( .A1(n13592), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13574) );
  OAI21_X1 U16924 ( .B1(n13592), .B2(n14893), .A(n13574), .ZN(n15820) );
  AOI22_X1 U16925 ( .A1(n13595), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15820), .B2(n20555), .ZN(n13589) );
  MUX2_X1 U16926 ( .A(n13575), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n13564), .Z(n13576) );
  NOR2_X1 U16927 ( .A1(n13576), .A2(n11234), .ZN(n13577) );
  NAND2_X1 U16928 ( .A1(n13578), .A2(n13577), .ZN(n13585) );
  NAND2_X1 U16929 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13579) );
  AOI22_X1 U16930 ( .A1(n11234), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n11227), .B2(n13579), .ZN(n13583) );
  AOI21_X1 U16931 ( .B1(n13564), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11227), .ZN(n13580) );
  NOR2_X1 U16932 ( .A1(n11278), .A2(n13580), .ZN(n20634) );
  NOR2_X1 U16933 ( .A1(n13581), .A2(n20634), .ZN(n13582) );
  AOI21_X1 U16934 ( .B1(n14877), .B2(n13583), .A(n13582), .ZN(n13584) );
  NAND2_X1 U16935 ( .A1(n13585), .A2(n13584), .ZN(n13586) );
  AOI21_X1 U16936 ( .B1(n20272), .B2(n13587), .A(n13586), .ZN(n20636) );
  MUX2_X1 U16937 ( .A(n11227), .B(n20636), .S(n15814), .Z(n15821) );
  INV_X1 U16938 ( .A(n15821), .ZN(n15825) );
  AOI22_X1 U16939 ( .A1(n15825), .A2(n20555), .B1(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13595), .ZN(n13588) );
  INV_X1 U16940 ( .A(n20157), .ZN(n20387) );
  OR2_X1 U16941 ( .A1(n11483), .A2(n20387), .ZN(n13591) );
  XNOR2_X1 U16942 ( .A(n13591), .B(n16158), .ZN(n19887) );
  OAI21_X1 U16943 ( .B1(n19887), .B2(n12048), .A(n15814), .ZN(n13594) );
  AOI21_X1 U16944 ( .B1(n13592), .B2(n16158), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n13593) );
  NAND2_X1 U16945 ( .A1(n13594), .A2(n13593), .ZN(n13597) );
  NAND2_X1 U16946 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n13595), .ZN(
        n13596) );
  NAND2_X1 U16947 ( .A1(n13597), .A2(n13596), .ZN(n15831) );
  INV_X1 U16948 ( .A(n15831), .ZN(n13598) );
  OAI21_X1 U16949 ( .B1(n15832), .B2(n13590), .A(n13598), .ZN(n13607) );
  NOR2_X1 U16950 ( .A1(n20556), .A2(n16170), .ZN(n14300) );
  OAI21_X1 U16951 ( .B1(n13607), .B2(P1_FLUSH_REG_SCAN_IN), .A(n14300), .ZN(
        n13600) );
  NAND2_X1 U16952 ( .A1(n20417), .A2(n20555), .ZN(n16165) );
  INV_X1 U16953 ( .A(n16165), .ZN(n20671) );
  AND2_X1 U16954 ( .A1(n20389), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20644) );
  NOR2_X1 U16955 ( .A1(n13568), .A2(n20644), .ZN(n13604) );
  NAND2_X1 U16956 ( .A1(n13601), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13602) );
  NOR2_X1 U16957 ( .A1(n13602), .A2(n20646), .ZN(n20651) );
  NAND2_X1 U16958 ( .A1(n13602), .A2(n20641), .ZN(n14873) );
  MUX2_X1 U16959 ( .A(n20651), .B(n20499), .S(n20268), .Z(n13603) );
  OAI21_X1 U16960 ( .B1(n13604), .B2(n13603), .A(n20653), .ZN(n13605) );
  OAI21_X1 U16961 ( .B1(n20653), .B2(n20274), .A(n13605), .ZN(P1_U3476) );
  INV_X1 U16962 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n19924) );
  OAI222_X1 U16963 ( .A1(n13606), .A2(n15997), .B1(n14573), .B2(n20041), .C1(
        n14571), .C2(n19924), .ZN(P1_U2901) );
  NOR2_X1 U16964 ( .A1(n13607), .A2(n16170), .ZN(n15841) );
  INV_X1 U16965 ( .A(n11568), .ZN(n20125) );
  OAI22_X1 U16966 ( .A1(n12818), .A2(n20646), .B1(n20125), .B2(n20644), .ZN(
        n13608) );
  OAI21_X1 U16967 ( .B1(n15841), .B2(n13608), .A(n20653), .ZN(n13609) );
  OAI21_X1 U16968 ( .B1(n20653), .B2(n20415), .A(n13609), .ZN(P1_U3478) );
  NAND2_X1 U16969 ( .A1(n13612), .A2(n13611), .ZN(n13613) );
  INV_X1 U16970 ( .A(n19967), .ZN(n13618) );
  OAI21_X1 U16971 ( .B1(n13615), .B2(n13614), .A(n13682), .ZN(n13616) );
  INV_X1 U16972 ( .A(n13616), .ZN(n19973) );
  AOI22_X1 U16973 ( .A1(n19973), .A2(n19894), .B1(P1_EBX_REG_4__SCAN_IN), .B2(
        n14510), .ZN(n13617) );
  OAI21_X1 U16974 ( .B1(n13618), .B2(n14515), .A(n13617), .ZN(P1_U2868) );
  INV_X1 U16975 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19922) );
  OAI222_X1 U16976 ( .A1(n13618), .A2(n15997), .B1(n14573), .B2(n20045), .C1(
        n14571), .C2(n19922), .ZN(P1_U2900) );
  AND2_X1 U16977 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20556), .ZN(n13620) );
  NAND2_X1 U16978 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20671), .ZN(n16164) );
  INV_X1 U16979 ( .A(n16164), .ZN(n13619) );
  AOI22_X1 U16980 ( .A1(n13621), .A2(n13620), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n13619), .ZN(n13622) );
  NAND2_X1 U16981 ( .A1(n16122), .A2(n13622), .ZN(n13623) );
  INV_X1 U16982 ( .A(n14317), .ZN(n13626) );
  AOI21_X1 U16983 ( .B1(n13627), .B2(n13639), .A(n19857), .ZN(n13754) );
  OAI21_X1 U16984 ( .B1(n19852), .B2(n19876), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13643) );
  NAND2_X1 U16985 ( .A1(n13629), .A2(n15835), .ZN(n13637) );
  NAND2_X1 U16986 ( .A1(n13630), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13632) );
  AND3_X1 U16987 ( .A1(n13637), .A2(n11372), .A3(n13632), .ZN(n13631) );
  NOR2_X1 U16988 ( .A1(n13632), .A2(n15835), .ZN(n13633) );
  AOI22_X1 U16989 ( .A1(P1_EBX_REG_0__SCAN_IN), .A2(n19875), .B1(n19884), .B2(
        n13634), .ZN(n13642) );
  INV_X1 U16990 ( .A(n13635), .ZN(n13636) );
  AND2_X1 U16991 ( .A1(n13639), .A2(n13636), .ZN(n13764) );
  NAND2_X1 U16992 ( .A1(n11568), .A2(n13764), .ZN(n13641) );
  NOR2_X1 U16993 ( .A1(n13637), .A2(n20024), .ZN(n13638) );
  NAND2_X1 U16994 ( .A1(n19835), .A2(n19831), .ZN(n19833) );
  NAND2_X1 U16995 ( .A1(n19833), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13640) );
  AND4_X1 U16996 ( .A1(n13643), .A2(n13642), .A3(n13641), .A4(n13640), .ZN(
        n13644) );
  OAI21_X1 U16997 ( .B1(n13754), .B2(n13645), .A(n13644), .ZN(P1_U2840) );
  INV_X1 U16998 ( .A(n13764), .ZN(n19886) );
  NAND2_X1 U16999 ( .A1(n19812), .A2(n13655), .ZN(n13648) );
  INV_X1 U17000 ( .A(n19831), .ZN(n19805) );
  AOI22_X1 U17001 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(n19875), .B1(n19805), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n13647) );
  OAI211_X1 U17002 ( .C1(n19867), .C2(n13652), .A(n13648), .B(n13647), .ZN(
        n13649) );
  AOI21_X1 U17003 ( .B1(n19884), .B2(n13284), .A(n13649), .ZN(n13650) );
  OAI21_X1 U17004 ( .B1(n13646), .B2(n19886), .A(n13650), .ZN(n13651) );
  AOI21_X1 U17005 ( .B1(n19852), .B2(n13652), .A(n13651), .ZN(n13653) );
  OAI21_X1 U17006 ( .B1(n13754), .B2(n13654), .A(n13653), .ZN(P1_U2839) );
  INV_X1 U17007 ( .A(n13568), .ZN(n20273) );
  NOR2_X1 U17008 ( .A1(n19835), .A2(n13655), .ZN(n13758) );
  INV_X1 U17009 ( .A(n13758), .ZN(n19882) );
  OAI21_X1 U17010 ( .B1(n19805), .B2(n13655), .A(n19833), .ZN(n13656) );
  INV_X1 U17011 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20578) );
  OAI22_X1 U17012 ( .A1(n13656), .A2(n20578), .B1(n19862), .B2(n19997), .ZN(
        n13657) );
  AOI21_X1 U17013 ( .B1(n19876), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n13657), .ZN(n13659) );
  NAND2_X1 U17014 ( .A1(n19875), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n13658) );
  OAI211_X1 U17015 ( .C1(n19882), .C2(P1_REIP_REG_2__SCAN_IN), .A(n13659), .B(
        n13658), .ZN(n13662) );
  NOR2_X1 U17016 ( .A1(n19892), .A2(n13660), .ZN(n13661) );
  AOI211_X1 U17017 ( .C1(n13764), .C2(n20273), .A(n13662), .B(n13661), .ZN(
        n13663) );
  OAI21_X1 U17018 ( .B1(n13754), .B2(n13664), .A(n13663), .ZN(P1_U2838) );
  XNOR2_X1 U17019 ( .A(n13665), .B(n13666), .ZN(n13670) );
  NAND2_X1 U17020 ( .A1(n13674), .A2(n13667), .ZN(n13668) );
  NAND2_X1 U17021 ( .A1(n13896), .A2(n13668), .ZN(n15724) );
  MUX2_X1 U17022 ( .A(n15724), .B(n13931), .S(n13198), .Z(n13669) );
  OAI21_X1 U17023 ( .B1(n13670), .B2(n15114), .A(n13669), .ZN(P2_U2875) );
  OR2_X1 U17024 ( .A1(n13672), .A2(n13671), .ZN(n13673) );
  NAND2_X1 U17025 ( .A1(n13674), .A2(n13673), .ZN(n16286) );
  INV_X1 U17026 ( .A(n13665), .ZN(n13675) );
  OAI211_X1 U17027 ( .C1(n9727), .C2(n9661), .A(n13675), .B(n15119), .ZN(
        n13677) );
  NAND2_X1 U17028 ( .A1(n13198), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n13676) );
  OAI211_X1 U17029 ( .C1(n15122), .C2(n16286), .A(n13677), .B(n13676), .ZN(
        P2_U2876) );
  NAND2_X1 U17030 ( .A1(n13610), .A2(n13679), .ZN(n13680) );
  AND2_X1 U17031 ( .A1(n13678), .A2(n13680), .ZN(n19871) );
  INV_X1 U17032 ( .A(n19871), .ZN(n13753) );
  INV_X1 U17033 ( .A(n14003), .ZN(n13681) );
  AOI21_X1 U17034 ( .B1(n13683), .B2(n13682), .A(n13681), .ZN(n19863) );
  AOI22_X1 U17035 ( .A1(n19863), .A2(n19894), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n14510), .ZN(n13684) );
  OAI21_X1 U17036 ( .B1(n13753), .B2(n14515), .A(n13684), .ZN(P1_U2867) );
  INV_X1 U17037 ( .A(n13842), .ZN(n13689) );
  INV_X1 U17038 ( .A(n13685), .ZN(n13686) );
  OAI22_X1 U17039 ( .A1(n13689), .A2(n13706), .B1(n13687), .B2(n13686), .ZN(
        n13688) );
  AOI21_X1 U17040 ( .B1(n13689), .B2(n13705), .A(n13688), .ZN(n19751) );
  INV_X1 U17041 ( .A(n13690), .ZN(n13693) );
  INV_X1 U17042 ( .A(n10929), .ZN(n13692) );
  AOI22_X1 U17043 ( .A1(n13693), .A2(n12687), .B1(n13692), .B2(n9618), .ZN(
        n13698) );
  INV_X1 U17044 ( .A(n13694), .ZN(n13696) );
  NOR3_X1 U17045 ( .A1(n13696), .A2(n13695), .A3(n13779), .ZN(n18833) );
  OAI21_X1 U17046 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n18833), .ZN(n13697) );
  NAND3_X1 U17047 ( .A1(n19751), .A2(n13698), .A3(n13697), .ZN(n13745) );
  INV_X1 U17048 ( .A(n13727), .ZN(n13731) );
  NAND2_X1 U17049 ( .A1(n9620), .A2(n13320), .ZN(n13726) );
  NOR2_X1 U17050 ( .A1(n10674), .A2(n10596), .ZN(n13714) );
  INV_X1 U17051 ( .A(n13714), .ZN(n13704) );
  NAND2_X1 U17052 ( .A1(n13320), .A2(n13699), .ZN(n13703) );
  NAND2_X1 U17053 ( .A1(n9617), .A2(n13700), .ZN(n13713) );
  NAND2_X1 U17054 ( .A1(n13713), .A2(n13701), .ZN(n13702) );
  NAND4_X1 U17055 ( .A1(n13726), .A2(n13704), .A3(n13703), .A4(n13702), .ZN(
        n13710) );
  INV_X1 U17056 ( .A(n13705), .ZN(n13707) );
  AND2_X1 U17057 ( .A1(n13707), .A2(n13706), .ZN(n13717) );
  NAND3_X1 U17058 ( .A1(n13320), .A2(n10596), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13708) );
  OAI21_X1 U17059 ( .B1(n13717), .B2(n13714), .A(n13708), .ZN(n13709) );
  MUX2_X1 U17060 ( .A(n13710), .B(n13709), .S(n10430), .Z(n13711) );
  MUX2_X1 U17061 ( .A(n10430), .B(n15767), .S(n13722), .Z(n13743) );
  INV_X1 U17062 ( .A(n13713), .ZN(n13716) );
  NOR2_X1 U17063 ( .A1(n13714), .A2(n9638), .ZN(n13715) );
  MUX2_X1 U17064 ( .A(n13717), .B(n13716), .S(n13715), .Z(n13720) );
  NAND2_X1 U17065 ( .A1(n13320), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13718) );
  MUX2_X1 U17066 ( .A(n13718), .B(n13726), .S(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n13719) );
  NAND2_X1 U17067 ( .A1(n13720), .A2(n13719), .ZN(n13721) );
  AOI21_X1 U17068 ( .B1(n10647), .B2(n13731), .A(n13721), .ZN(n15763) );
  MUX2_X1 U17069 ( .A(n13699), .B(n15763), .S(n13722), .Z(n13742) );
  INV_X1 U17070 ( .A(n13742), .ZN(n13740) );
  NAND2_X1 U17071 ( .A1(n19718), .A2(n19725), .ZN(n19197) );
  INV_X1 U17072 ( .A(n19197), .ZN(n19167) );
  INV_X1 U17073 ( .A(n13743), .ZN(n13737) );
  INV_X1 U17074 ( .A(n12655), .ZN(n13724) );
  NAND2_X1 U17075 ( .A1(n13724), .A2(n13723), .ZN(n13729) );
  OAI21_X1 U17076 ( .B1(n10672), .B2(n10670), .A(n13729), .ZN(n13725) );
  OAI211_X1 U17077 ( .C1(n13728), .C2(n13727), .A(n13726), .B(n13725), .ZN(
        n14071) );
  INV_X1 U17078 ( .A(n14071), .ZN(n13734) );
  MUX2_X1 U17079 ( .A(n13729), .B(n13320), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n13730) );
  AOI21_X1 U17080 ( .B1(n19079), .B2(n13731), .A(n13730), .ZN(n14023) );
  INV_X1 U17081 ( .A(n14023), .ZN(n13732) );
  AOI211_X1 U17082 ( .C1(n14071), .C2(n19735), .A(n20827), .B(n13732), .ZN(
        n13733) );
  AOI21_X1 U17083 ( .B1(n13734), .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n13733), .ZN(n13736) );
  NAND2_X1 U17084 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n13742), .ZN(
        n13735) );
  OAI211_X1 U17085 ( .C1(n13737), .C2(n19718), .A(n13736), .B(n13735), .ZN(
        n13738) );
  OAI22_X1 U17086 ( .A1(n13746), .A2(n13738), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n13743), .ZN(n13739) );
  AOI21_X1 U17087 ( .B1(n13740), .B2(n19167), .A(n13739), .ZN(n13741) );
  OAI22_X1 U17088 ( .A1(n13743), .A2(n13742), .B1(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n13741), .ZN(n13744) );
  AOI211_X1 U17089 ( .C1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n13746), .A(
        n13745), .B(n13744), .ZN(n16324) );
  AOI21_X1 U17090 ( .B1(n16324), .B2(n19726), .A(n19762), .ZN(n13751) );
  NOR3_X1 U17091 ( .A1(n13748), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n13747), 
        .ZN(n13750) );
  OR2_X1 U17092 ( .A1(n13749), .A2(n19350), .ZN(n19755) );
  INV_X1 U17093 ( .A(n19625), .ZN(n19627) );
  OAI21_X1 U17094 ( .B1(n19627), .B2(n19762), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n13752) );
  NAND2_X1 U17095 ( .A1(n13752), .A2(n15874), .ZN(P2_U3593) );
  OAI222_X1 U17096 ( .A1(n13753), .A2(n15997), .B1(n14573), .B2(n20049), .C1(
        n14571), .C2(n11600), .ZN(P1_U2899) );
  INV_X1 U17097 ( .A(n13754), .ZN(n19889) );
  NAND2_X1 U17098 ( .A1(n19889), .A2(n13755), .ZN(n13766) );
  AOI21_X1 U17099 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_2__SCAN_IN), 
        .A(n19835), .ZN(n13756) );
  OAI21_X1 U17100 ( .B1(n13756), .B2(n19805), .A(P1_REIP_REG_3__SCAN_IN), .ZN(
        n13762) );
  AOI22_X1 U17101 ( .A1(n19875), .A2(P1_EBX_REG_3__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n19876), .ZN(n13761) );
  NAND2_X1 U17102 ( .A1(n19980), .A2(n19884), .ZN(n13760) );
  INV_X1 U17103 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13757) );
  NAND3_X1 U17104 ( .A1(n13758), .A2(n13757), .A3(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n13759) );
  NAND4_X1 U17105 ( .A1(n13762), .A2(n13761), .A3(n13760), .A4(n13759), .ZN(
        n13763) );
  AOI21_X1 U17106 ( .B1(n20272), .B2(n13764), .A(n13763), .ZN(n13765) );
  OAI211_X1 U17107 ( .C1(n19892), .C2(n13767), .A(n13766), .B(n13765), .ZN(
        P1_U2837) );
  XNOR2_X1 U17108 ( .A(n13768), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15225) );
  NAND2_X1 U17109 ( .A1(n15225), .A2(n19762), .ZN(n13770) );
  INV_X1 U17110 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15470) );
  AOI21_X1 U17111 ( .B1(n14106), .B2(n13771), .A(n13775), .ZN(n14108) );
  AOI21_X1 U17112 ( .B1(n19068), .B2(n13772), .A(n13773), .ZN(n19058) );
  AOI22_X1 U17113 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n19762), .ZN(n14066) );
  AOI22_X1 U17114 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n13145), .B2(n19762), .ZN(
        n14065) );
  NAND2_X1 U17115 ( .A1(n14066), .A2(n14065), .ZN(n14064) );
  NOR2_X1 U17116 ( .A1(n13974), .A2(n14064), .ZN(n13801) );
  OAI21_X1 U17117 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n13153), .A(
        n13772), .ZN(n13870) );
  NAND2_X1 U17118 ( .A1(n13801), .A2(n13870), .ZN(n13884) );
  NOR2_X1 U17119 ( .A1(n19058), .A2(n13884), .ZN(n18941) );
  OAI21_X1 U17120 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n13773), .A(
        n13771), .ZN(n18944) );
  NAND2_X1 U17121 ( .A1(n18941), .A2(n18944), .ZN(n13962) );
  NOR2_X1 U17122 ( .A1(n14108), .A2(n13962), .ZN(n13912) );
  NOR2_X1 U17123 ( .A1(n18942), .A2(n13912), .ZN(n13776) );
  OAI21_X1 U17124 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n13775), .A(
        n13774), .ZN(n14162) );
  XNOR2_X1 U17125 ( .A(n13776), .B(n14162), .ZN(n13799) );
  NOR3_X1 U17126 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15873) );
  NAND2_X1 U17127 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15873), .ZN(n19628) );
  XNOR2_X1 U17128 ( .A(n13777), .B(n13778), .ZN(n18982) );
  NAND2_X1 U17129 ( .A1(n11212), .A2(n13779), .ZN(n13787) );
  NOR2_X1 U17130 ( .A1(n19761), .A2(n13787), .ZN(n13780) );
  NOR2_X1 U17131 ( .A1(n18982), .A2(n18947), .ZN(n13798) );
  NOR2_X1 U17132 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19768), .ZN(n13789) );
  AND2_X1 U17133 ( .A1(n9628), .A2(n13789), .ZN(n13781) );
  NOR2_X1 U17134 ( .A1(n19737), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19321) );
  INV_X1 U17135 ( .A(n19321), .ZN(n19624) );
  NOR2_X1 U17136 ( .A1(n19631), .A2(n19624), .ZN(n16316) );
  INV_X1 U17137 ( .A(n16316), .ZN(n13782) );
  NAND2_X1 U17138 ( .A1(n19628), .A2(n13782), .ZN(n13783) );
  OR2_X1 U17139 ( .A1(n18939), .A2(n13783), .ZN(n13784) );
  INV_X1 U17140 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n15052) );
  NOR2_X1 U17141 ( .A1(n13789), .A2(n15052), .ZN(n13785) );
  AND2_X1 U17142 ( .A1(n9628), .A2(n13785), .ZN(n13786) );
  AND2_X1 U17143 ( .A1(n13788), .A2(n13787), .ZN(n16172) );
  INV_X1 U17144 ( .A(n13789), .ZN(n13790) );
  AND3_X1 U17145 ( .A1(n13791), .A2(n15052), .A3(n13790), .ZN(n13792) );
  AOI22_X1 U17146 ( .A1(n13793), .A2(n18923), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n18922), .ZN(n13794) );
  OAI211_X1 U17147 ( .C1(n19659), .C2(n18927), .A(n13794), .B(n18925), .ZN(
        n13795) );
  AOI21_X1 U17148 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18931), .A(
        n13795), .ZN(n13796) );
  OAI21_X1 U17149 ( .B1(n18946), .B2(n14172), .A(n13796), .ZN(n13797) );
  AOI211_X1 U17150 ( .C1(n13799), .C2(n18949), .A(n13798), .B(n13797), .ZN(
        n13800) );
  INV_X1 U17151 ( .A(n13800), .ZN(P2_U2848) );
  NOR2_X1 U17152 ( .A1(n18942), .A2(n13801), .ZN(n13802) );
  XNOR2_X1 U17153 ( .A(n13802), .B(n13870), .ZN(n13815) );
  NOR2_X1 U17154 ( .A1(n19145), .A2(n14122), .ZN(n13814) );
  OR2_X1 U17155 ( .A1(n13804), .A2(n13803), .ZN(n13806) );
  NAND2_X1 U17156 ( .A1(n13806), .A2(n13805), .ZN(n18985) );
  INV_X1 U17157 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13871) );
  OAI22_X1 U17158 ( .A1(n13871), .A2(n18935), .B1(n12713), .B2(n18927), .ZN(
        n13810) );
  NAND2_X1 U17159 ( .A1(n18922), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n13807) );
  OAI21_X1 U17160 ( .B1(n13808), .B2(n18936), .A(n13807), .ZN(n13809) );
  NOR2_X1 U17161 ( .A1(n13810), .A2(n13809), .ZN(n13812) );
  NAND2_X1 U17162 ( .A1(n13412), .A2(n18902), .ZN(n13811) );
  OAI211_X1 U17163 ( .C1(n18985), .C2(n18947), .A(n13812), .B(n13811), .ZN(
        n13813) );
  AOI211_X1 U17164 ( .C1(n13815), .C2(n18949), .A(n13814), .B(n13813), .ZN(
        n13816) );
  INV_X1 U17165 ( .A(n13816), .ZN(P2_U2852) );
  XNOR2_X1 U17166 ( .A(n13818), .B(n13817), .ZN(n19061) );
  OAI21_X1 U17167 ( .B1(n13819), .B2(n16300), .A(n13820), .ZN(n19060) );
  NAND2_X1 U17168 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13821), .ZN(
        n13828) );
  NAND2_X1 U17169 ( .A1(n13823), .A2(n13822), .ZN(n13830) );
  INV_X1 U17170 ( .A(n13830), .ZN(n13824) );
  AOI21_X1 U17171 ( .B1(n13831), .B2(n13828), .A(n13824), .ZN(n13825) );
  NAND2_X1 U17172 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14167), .ZN(
        n16299) );
  INV_X1 U17173 ( .A(n13826), .ZN(n13827) );
  AOI21_X1 U17174 ( .B1(n13829), .B2(n13828), .A(n13827), .ZN(n15457) );
  OAI21_X1 U17175 ( .B1(n13831), .B2(n13830), .A(n15457), .ZN(n14168) );
  AOI21_X1 U17176 ( .B1(n15611), .B2(n13877), .A(n14168), .ZN(n16304) );
  NAND2_X1 U17177 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n13328), .ZN(n13832) );
  OAI221_X1 U17178 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n16299), .C1(
        n16300), .C2(n16304), .A(n13832), .ZN(n13838) );
  NAND2_X1 U17179 ( .A1(n13833), .A2(n13805), .ZN(n13836) );
  INV_X1 U17180 ( .A(n13834), .ZN(n13835) );
  NAND2_X1 U17181 ( .A1(n13836), .A2(n13835), .ZN(n18995) );
  OAI22_X1 U17182 ( .A1(n13887), .A2(n16315), .B1(n16305), .B2(n18995), .ZN(
        n13837) );
  AOI211_X1 U17183 ( .C1(n19060), .C2(n16282), .A(n13838), .B(n13837), .ZN(
        n13839) );
  OAI21_X1 U17184 ( .B1(n19061), .B2(n16306), .A(n13839), .ZN(P2_U3042) );
  NOR2_X2 U17185 ( .A1(n19494), .A2(n19707), .ZN(n19481) );
  OAI21_X1 U17186 ( .B1(n19481), .B2(n19515), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13849) );
  NOR2_X1 U17187 ( .A1(n13840), .A2(n19289), .ZN(n19226) );
  NAND2_X1 U17188 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19226), .ZN(
        n13848) );
  INV_X1 U17189 ( .A(n10807), .ZN(n13841) );
  AOI21_X1 U17190 ( .B1(n13841), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13846) );
  NAND3_X1 U17191 ( .A1(n19735), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19489) );
  NOR2_X1 U17192 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19489), .ZN(
        n19479) );
  INV_X1 U17193 ( .A(n19742), .ZN(n13844) );
  NAND2_X1 U17194 ( .A1(n19762), .A2(n18829), .ZN(n19767) );
  INV_X1 U17195 ( .A(n19767), .ZN(n13843) );
  OAI21_X1 U17196 ( .B1(n13846), .B2(n19479), .A(n19573), .ZN(n13847) );
  AOI22_X1 U17197 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19127), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19126), .ZN(n19549) );
  INV_X1 U17198 ( .A(n19606), .ZN(n19546) );
  AOI22_X1 U17199 ( .A1(n19515), .A2(n19603), .B1(n19481), .B2(n19546), .ZN(
        n13859) );
  INV_X1 U17200 ( .A(n13853), .ZN(n13856) );
  INV_X1 U17201 ( .A(n19226), .ZN(n13855) );
  OAI21_X1 U17202 ( .B1(n10807), .B2(n19479), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13854) );
  INV_X1 U17203 ( .A(n18984), .ZN(n13857) );
  NOR2_X2 U17204 ( .A1(n13857), .A2(n19523), .ZN(n19602) );
  AOI22_X1 U17205 ( .A1(n19480), .A2(n19602), .B1(n19601), .B2(n19479), .ZN(
        n13858) );
  OAI211_X1 U17206 ( .C1(n19484), .C2(n13860), .A(n13859), .B(n13858), .ZN(
        P2_U3149) );
  INV_X1 U17207 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13863) );
  AOI22_X1 U17208 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19127), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19126), .ZN(n19561) );
  AOI22_X1 U17209 ( .A1(n19515), .A2(n19617), .B1(n19481), .B2(n19556), .ZN(
        n13862) );
  NOR2_X2 U17210 ( .A1(n18981), .A2(n19523), .ZN(n19615) );
  AOI22_X1 U17211 ( .A1(n19480), .A2(n19615), .B1(n19479), .B2(n19613), .ZN(
        n13861) );
  OAI211_X1 U17212 ( .C1(n19484), .C2(n13863), .A(n13862), .B(n13861), .ZN(
        P2_U3151) );
  XNOR2_X1 U17213 ( .A(n13864), .B(n13865), .ZN(n13883) );
  NAND2_X1 U17214 ( .A1(n13867), .A2(n13866), .ZN(n13868) );
  XOR2_X1 U17215 ( .A(n13869), .B(n13868), .Z(n13876) );
  NAND2_X1 U17216 ( .A1(n13876), .A2(n16250), .ZN(n13875) );
  NOR2_X1 U17217 ( .A1(n16262), .A2(n13870), .ZN(n13873) );
  NAND2_X1 U17218 ( .A1(n18939), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n13878) );
  OAI21_X1 U17219 ( .B1(n19067), .B2(n13871), .A(n13878), .ZN(n13872) );
  OAI211_X1 U17220 ( .C1(n13883), .C2(n19075), .A(n13875), .B(n13874), .ZN(
        P2_U3011) );
  NAND2_X1 U17221 ( .A1(n13876), .A2(n16281), .ZN(n13882) );
  INV_X1 U17222 ( .A(n14168), .ZN(n15461) );
  INV_X1 U17223 ( .A(n14167), .ZN(n14098) );
  MUX2_X1 U17224 ( .A(n15461), .B(n14098), .S(n13877), .Z(n13879) );
  OAI211_X1 U17225 ( .C1(n18985), .C2(n16305), .A(n13879), .B(n13878), .ZN(
        n13880) );
  AOI21_X1 U17226 ( .B1(n12157), .B2(n15757), .A(n13880), .ZN(n13881) );
  OAI211_X1 U17227 ( .C1(n13883), .C2(n16308), .A(n13882), .B(n13881), .ZN(
        P2_U3043) );
  AND2_X1 U17228 ( .A1(n18893), .A2(n13884), .ZN(n13886) );
  AOI21_X1 U17229 ( .B1(n19058), .B2(n13886), .A(n19628), .ZN(n13885) );
  OAI21_X1 U17230 ( .B1(n19058), .B2(n13886), .A(n13885), .ZN(n13894) );
  INV_X1 U17231 ( .A(n13887), .ZN(n19064) );
  OAI21_X1 U17232 ( .B1(n18935), .B2(n19068), .A(n18925), .ZN(n13889) );
  OAI22_X1 U17233 ( .A1(n18927), .A2(n12720), .B1(n18947), .B2(n18995), .ZN(
        n13888) );
  AOI211_X1 U17234 ( .C1(P2_EBX_REG_4__SCAN_IN), .C2(n18922), .A(n13889), .B(
        n13888), .ZN(n13890) );
  OAI21_X1 U17235 ( .B1(n13891), .B2(n18936), .A(n13890), .ZN(n13892) );
  AOI21_X1 U17236 ( .B1(n19064), .B2(n18902), .A(n13892), .ZN(n13893) );
  OAI211_X1 U17237 ( .C1(n18997), .C2(n14122), .A(n13894), .B(n13893), .ZN(
        P2_U2851) );
  AOI21_X1 U17238 ( .B1(n13897), .B2(n13896), .A(n13895), .ZN(n15707) );
  INV_X1 U17239 ( .A(n15707), .ZN(n18913) );
  INV_X1 U17240 ( .A(n13898), .ZN(n13902) );
  INV_X1 U17241 ( .A(n13900), .ZN(n13906) );
  OAI211_X1 U17242 ( .C1(n13902), .C2(n13901), .A(n15119), .B(n13906), .ZN(
        n13904) );
  NAND2_X1 U17243 ( .A1(n13198), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13903) );
  OAI211_X1 U17244 ( .C1(n18913), .C2(n15122), .A(n13904), .B(n13903), .ZN(
        P2_U2874) );
  XNOR2_X1 U17245 ( .A(n13906), .B(n13905), .ZN(n13910) );
  NOR2_X1 U17246 ( .A1(n13895), .A2(n13907), .ZN(n13908) );
  OR2_X1 U17247 ( .A1(n14040), .A2(n13908), .ZN(n18900) );
  MUX2_X1 U17248 ( .A(n18900), .B(n18896), .S(n13198), .Z(n13909) );
  OAI21_X1 U17249 ( .B1(n13910), .B2(n15114), .A(n13909), .ZN(P2_U2873) );
  AOI21_X1 U17250 ( .B1(n15442), .B2(n13774), .A(n13911), .ZN(n15445) );
  NAND2_X1 U17251 ( .A1(n13912), .A2(n14162), .ZN(n13927) );
  NAND2_X1 U17252 ( .A1(n18893), .A2(n13927), .ZN(n13913) );
  XNOR2_X1 U17253 ( .A(n15445), .B(n13913), .ZN(n13922) );
  AOI22_X1 U17254 ( .A1(n13914), .A2(n18923), .B1(P2_EBX_REG_8__SCAN_IN), .B2(
        n18922), .ZN(n13915) );
  OAI211_X1 U17255 ( .C1(n12736), .C2(n18927), .A(n13915), .B(n18925), .ZN(
        n13916) );
  AOI21_X1 U17256 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18931), .A(
        n13916), .ZN(n13920) );
  AOI21_X1 U17257 ( .B1(n13918), .B2(n13917), .A(n16287), .ZN(n15749) );
  NAND2_X1 U17258 ( .A1(n18901), .A2(n15749), .ZN(n13919) );
  OAI211_X1 U17259 ( .C1(n15748), .C2(n18946), .A(n13920), .B(n13919), .ZN(
        n13921) );
  AOI21_X1 U17260 ( .B1(n13922), .B2(n18949), .A(n13921), .ZN(n13923) );
  INV_X1 U17261 ( .A(n13923), .ZN(P2_U2847) );
  AOI21_X1 U17262 ( .B1(n15425), .B2(n13929), .A(n13924), .ZN(n15426) );
  AOI21_X1 U17263 ( .B1(n16261), .B2(n13928), .A(n13926), .ZN(n16254) );
  NOR2_X1 U17264 ( .A1(n15445), .A2(n13927), .ZN(n18919) );
  OAI21_X1 U17265 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n13911), .A(
        n13928), .ZN(n18921) );
  NAND2_X1 U17266 ( .A1(n18919), .A2(n18921), .ZN(n13985) );
  NOR2_X1 U17267 ( .A1(n16254), .A2(n13985), .ZN(n13944) );
  OAI21_X1 U17268 ( .B1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n13926), .A(
        n13929), .ZN(n13945) );
  NAND2_X1 U17269 ( .A1(n13944), .A2(n13945), .ZN(n14898) );
  NAND2_X1 U17270 ( .A1(n18893), .A2(n14898), .ZN(n13930) );
  XNOR2_X1 U17271 ( .A(n15426), .B(n13930), .ZN(n13941) );
  OAI22_X1 U17272 ( .A1(n13932), .A2(n18936), .B1(n18954), .B2(n13931), .ZN(
        n13933) );
  INV_X1 U17273 ( .A(n13933), .ZN(n13934) );
  OAI211_X1 U17274 ( .C1(n12749), .C2(n18927), .A(n13934), .B(n18925), .ZN(
        n13935) );
  AOI21_X1 U17275 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18931), .A(
        n13935), .ZN(n13939) );
  AOI21_X1 U17276 ( .B1(n13937), .B2(n13947), .A(n13936), .ZN(n18968) );
  NAND2_X1 U17277 ( .A1(n18901), .A2(n18968), .ZN(n13938) );
  OAI211_X1 U17278 ( .C1(n15724), .C2(n18946), .A(n13939), .B(n13938), .ZN(
        n13940) );
  AOI21_X1 U17279 ( .B1(n13941), .B2(n18949), .A(n13940), .ZN(n13942) );
  INV_X1 U17280 ( .A(n13942), .ZN(P2_U2843) );
  INV_X1 U17281 ( .A(n13943), .ZN(n13956) );
  NOR2_X1 U17282 ( .A1(n18942), .A2(n19628), .ZN(n14079) );
  OAI211_X1 U17283 ( .C1(n13944), .C2(n13945), .A(n14079), .B(n14898), .ZN(
        n13955) );
  NOR2_X1 U17284 ( .A1(n19628), .A2(n18893), .ZN(n14118) );
  INV_X1 U17285 ( .A(n13945), .ZN(n16241) );
  OR2_X1 U17286 ( .A1(n13946), .A2(n13991), .ZN(n13948) );
  NAND2_X1 U17287 ( .A1(n13948), .A2(n13947), .ZN(n18972) );
  OR2_X1 U17288 ( .A1(n18947), .A2(n18972), .ZN(n13951) );
  NAND2_X1 U17289 ( .A1(n18922), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n13950) );
  AOI22_X1 U17290 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18931), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n18940), .ZN(n13949) );
  NAND4_X1 U17291 ( .A1(n13951), .A2(n13950), .A3(n13949), .A4(n18925), .ZN(
        n13953) );
  NOR2_X1 U17292 ( .A1(n16286), .A2(n18946), .ZN(n13952) );
  AOI211_X1 U17293 ( .C1(n14118), .C2(n16241), .A(n13953), .B(n13952), .ZN(
        n13954) );
  OAI211_X1 U17294 ( .C1(n13956), .C2(n18936), .A(n13955), .B(n13954), .ZN(
        P2_U2844) );
  INV_X1 U17295 ( .A(n13957), .ZN(n13959) );
  NAND3_X1 U17296 ( .A1(n16301), .A2(n13959), .A3(n13958), .ZN(n13960) );
  NAND2_X1 U17297 ( .A1(n13961), .A2(n13960), .ZN(n18983) );
  NAND2_X1 U17298 ( .A1(n18893), .A2(n13962), .ZN(n13963) );
  XNOR2_X1 U17299 ( .A(n14108), .B(n13963), .ZN(n13964) );
  NAND2_X1 U17300 ( .A1(n13964), .A2(n18949), .ZN(n13972) );
  OAI21_X1 U17301 ( .B1(n19657), .B2(n18927), .A(n18925), .ZN(n13965) );
  AOI21_X1 U17302 ( .B1(n18931), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n13965), .ZN(n13966) );
  OAI21_X1 U17303 ( .B1(n18954), .B2(n13967), .A(n13966), .ZN(n13970) );
  NOR2_X1 U17304 ( .A1(n13968), .A2(n18936), .ZN(n13969) );
  AOI211_X1 U17305 ( .C1(n14099), .C2(n18902), .A(n13970), .B(n13969), .ZN(
        n13971) );
  OAI211_X1 U17306 ( .C1(n18983), .C2(n18947), .A(n13972), .B(n13971), .ZN(
        P2_U2849) );
  NAND2_X1 U17307 ( .A1(n18893), .A2(n14064), .ZN(n13973) );
  XNOR2_X1 U17308 ( .A(n13974), .B(n13973), .ZN(n13975) );
  NAND2_X1 U17309 ( .A1(n13975), .A2(n18949), .ZN(n13984) );
  OAI22_X1 U17310 ( .A1(n18954), .A2(n13977), .B1(n18935), .B2(n13976), .ZN(
        n13979) );
  NOR2_X1 U17311 ( .A1(n18927), .A2(n19652), .ZN(n13978) );
  AOI211_X1 U17312 ( .C1(n18923), .C2(n13980), .A(n13979), .B(n13978), .ZN(
        n13981) );
  OAI21_X1 U17313 ( .B1(n18986), .B2(n18947), .A(n13981), .ZN(n13982) );
  AOI21_X1 U17314 ( .B1(n10647), .B2(n18902), .A(n13982), .ZN(n13983) );
  OAI211_X1 U17315 ( .C1(n19721), .C2(n14122), .A(n13984), .B(n13983), .ZN(
        P2_U2853) );
  NAND2_X1 U17316 ( .A1(n18893), .A2(n13985), .ZN(n13986) );
  XNOR2_X1 U17317 ( .A(n16254), .B(n13986), .ZN(n13998) );
  OAI22_X1 U17318 ( .A1(n13987), .A2(n18936), .B1(n18954), .B2(n13528), .ZN(
        n13988) );
  INV_X1 U17319 ( .A(n13988), .ZN(n13989) );
  OAI21_X1 U17320 ( .B1(n16261), .B2(n18935), .A(n13989), .ZN(n13997) );
  NAND2_X1 U17321 ( .A1(n16258), .A2(n18902), .ZN(n13994) );
  AOI21_X1 U17322 ( .B1(n13992), .B2(n13990), .A(n13991), .ZN(n18973) );
  AOI21_X1 U17323 ( .B1(n18901), .B2(n18973), .A(n13328), .ZN(n13993) );
  OAI211_X1 U17324 ( .C1(n18927), .C2(n13995), .A(n13994), .B(n13993), .ZN(
        n13996) );
  AOI211_X1 U17325 ( .C1(n13998), .C2(n18949), .A(n13997), .B(n13996), .ZN(
        n13999) );
  INV_X1 U17326 ( .A(n13999), .ZN(P2_U2845) );
  AND2_X1 U17327 ( .A1(n13678), .A2(n14001), .ZN(n14002) );
  NOR2_X1 U17328 ( .A1(n14000), .A2(n14002), .ZN(n19858) );
  INV_X1 U17329 ( .A(n19858), .ZN(n14006) );
  OAI222_X1 U17330 ( .A1(n14006), .A2(n15997), .B1(n14573), .B2(n20052), .C1(
        n14571), .C2(n11610), .ZN(P1_U2898) );
  INV_X1 U17331 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n14005) );
  AOI21_X1 U17332 ( .B1(n14004), .B2(n14003), .A(n16139), .ZN(n16147) );
  INV_X1 U17333 ( .A(n16147), .ZN(n19861) );
  OAI222_X1 U17334 ( .A1(n14006), .A2(n14515), .B1(n14005), .B2(n19899), .C1(
        n14532), .C2(n19861), .ZN(P1_U2866) );
  OR2_X1 U17335 ( .A1(n14000), .A2(n14009), .ZN(n14010) );
  AND2_X1 U17336 ( .A1(n14008), .A2(n14010), .ZN(n19896) );
  INV_X1 U17337 ( .A(n19896), .ZN(n14012) );
  OAI222_X1 U17338 ( .A1(n14012), .A2(n15997), .B1(n14573), .B2(n20059), .C1(
        n14011), .C2(n14571), .ZN(P1_U2897) );
  NAND2_X1 U17339 ( .A1(n14008), .A2(n14014), .ZN(n14015) );
  AND2_X1 U17340 ( .A1(n14013), .A2(n14015), .ZN(n19826) );
  INV_X1 U17341 ( .A(n19826), .ZN(n14021) );
  OAI21_X1 U17342 ( .B1(n14016), .B2(n14017), .A(n14145), .ZN(n14018) );
  INV_X1 U17343 ( .A(n14018), .ZN(n19819) );
  AOI22_X1 U17344 ( .A1(n19819), .A2(n19894), .B1(P1_EBX_REG_8__SCAN_IN), .B2(
        n14510), .ZN(n14019) );
  OAI21_X1 U17345 ( .B1(n14021), .B2(n14515), .A(n14019), .ZN(P1_U2864) );
  MUX2_X1 U17346 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n20020), .Z(
        n19935) );
  AOI22_X1 U17347 ( .A1(n14580), .A2(n19935), .B1(n16008), .B2(
        P1_EAX_REG_8__SCAN_IN), .ZN(n14020) );
  OAI21_X1 U17348 ( .B1(n14021), .B2(n15997), .A(n14020), .ZN(P1_U2896) );
  NOR2_X1 U17349 ( .A1(n12142), .A2(n16320), .ZN(n14025) );
  INV_X1 U17350 ( .A(n14066), .ZN(n14080) );
  AOI22_X1 U17351 ( .A1(n18942), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n14080), .B2(n18893), .ZN(n14069) );
  INV_X1 U17352 ( .A(n14069), .ZN(n14022) );
  OAI22_X1 U17353 ( .A1(n14023), .A2(n19708), .B1(n19726), .B2(n14022), .ZN(
        n14024) );
  OAI21_X1 U17354 ( .B1(n14025), .B2(n14024), .A(n14027), .ZN(n14026) );
  OAI21_X1 U17355 ( .B1(n14027), .B2(n10070), .A(n14026), .ZN(P2_U3601) );
  XNOR2_X1 U17356 ( .A(n14028), .B(n14029), .ZN(n16307) );
  OAI21_X1 U17357 ( .B1(n14033), .B2(n14031), .A(n14030), .ZN(n14032) );
  OAI21_X1 U17358 ( .B1(n10882), .B2(n14033), .A(n14032), .ZN(n16309) );
  NOR2_X1 U17359 ( .A1(n16309), .A2(n19075), .ZN(n14036) );
  NOR2_X1 U17360 ( .A1(n18945), .A2(n16272), .ZN(n14035) );
  INV_X1 U17361 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18934) );
  OAI22_X1 U17362 ( .A1(n18934), .A2(n19067), .B1(n16262), .B2(n18944), .ZN(
        n14034) );
  INV_X1 U17363 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n19655) );
  NOR2_X1 U17364 ( .A1(n19655), .A2(n18925), .ZN(n16313) );
  NOR4_X1 U17365 ( .A1(n14036), .A2(n14035), .A3(n14034), .A4(n16313), .ZN(
        n14037) );
  OAI21_X1 U17366 ( .B1(n19072), .B2(n16307), .A(n14037), .ZN(P2_U3009) );
  OR2_X1 U17367 ( .A1(n14040), .A2(n14039), .ZN(n14041) );
  AND2_X1 U17368 ( .A1(n14038), .A2(n14041), .ZN(n15677) );
  INV_X1 U17369 ( .A(n14043), .ZN(n14044) );
  OAI211_X1 U17370 ( .C1(n14042), .C2(n14045), .A(n14044), .B(n15119), .ZN(
        n14047) );
  NAND2_X1 U17371 ( .A1(n15122), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n14046) );
  OAI211_X1 U17372 ( .C1(n15042), .C2(n15122), .A(n14047), .B(n14046), .ZN(
        P2_U2872) );
  OAI21_X1 U17373 ( .B1(n14043), .B2(n14050), .A(n14049), .ZN(n14063) );
  OR2_X1 U17374 ( .A1(n15034), .A2(n14051), .ZN(n14052) );
  NAND2_X1 U17375 ( .A1(n15020), .A2(n14052), .ZN(n18883) );
  AOI22_X1 U17376 ( .A1(n18957), .A2(BUF1_REG_16__SCAN_IN), .B1(n18955), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n14055) );
  AOI22_X1 U17377 ( .A1(n16235), .A2(n14053), .B1(n19015), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n14054) );
  OAI211_X1 U17378 ( .C1(n15206), .C2(n18883), .A(n14055), .B(n14054), .ZN(
        n14056) );
  INV_X1 U17379 ( .A(n14056), .ZN(n14057) );
  OAI21_X1 U17380 ( .B1(n14063), .B2(n15185), .A(n14057), .ZN(P2_U2903) );
  NAND2_X1 U17381 ( .A1(n14038), .A2(n14058), .ZN(n14059) );
  NOR2_X1 U17382 ( .A1(n15110), .A2(n14060), .ZN(n14061) );
  AOI21_X1 U17383 ( .B1(n18885), .B2(n15110), .A(n14061), .ZN(n14062) );
  OAI21_X1 U17384 ( .B1(n14063), .B2(n15114), .A(n14062), .ZN(P2_U2871) );
  INV_X1 U17385 ( .A(n16320), .ZN(n14072) );
  OAI211_X1 U17386 ( .C1(n14066), .C2(n14065), .A(n18893), .B(n14064), .ZN(
        n14126) );
  OAI21_X1 U17387 ( .B1(n18893), .B2(n14067), .A(n14126), .ZN(n14068) );
  INV_X1 U17388 ( .A(n14068), .ZN(n15764) );
  NOR2_X1 U17389 ( .A1(n14069), .A2(n19726), .ZN(n15762) );
  AOI222_X1 U17390 ( .A1(n14073), .A2(n14072), .B1(n15764), .B2(n15762), .C1(
        n14071), .C2(n14070), .ZN(n14075) );
  NAND2_X1 U17391 ( .A1(n15768), .A2(n9619), .ZN(n14074) );
  OAI21_X1 U17392 ( .B1(n15768), .B2(n14075), .A(n14074), .ZN(P2_U3600) );
  INV_X1 U17393 ( .A(n14076), .ZN(n14077) );
  OAI22_X1 U17394 ( .A1(n18947), .A2(n14078), .B1(n18936), .B2(n14077), .ZN(
        n14084) );
  OAI21_X1 U17395 ( .B1(n18931), .B2(n14118), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14082) );
  NAND2_X1 U17396 ( .A1(n14080), .A2(n14079), .ZN(n14081) );
  OAI211_X1 U17397 ( .C1(n18954), .C2(n10574), .A(n14082), .B(n14081), .ZN(
        n14083) );
  AOI211_X1 U17398 ( .C1(P2_REIP_REG_0__SCAN_IN), .C2(n18940), .A(n14084), .B(
        n14083), .ZN(n14086) );
  NAND2_X1 U17399 ( .A1(n19079), .A2(n18902), .ZN(n14085) );
  OAI211_X1 U17400 ( .C1(n19739), .C2(n14122), .A(n14086), .B(n14085), .ZN(
        P2_U2855) );
  XNOR2_X1 U17401 ( .A(n14088), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14089) );
  XNOR2_X1 U17402 ( .A(n9604), .B(n14089), .ZN(n16135) );
  INV_X1 U17403 ( .A(n16135), .ZN(n14093) );
  AOI22_X1 U17404 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n20014), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n14090) );
  OAI21_X1 U17405 ( .B1(n19972), .B2(n19824), .A(n14090), .ZN(n14091) );
  AOI21_X1 U17406 ( .B1(n19826), .B2(n14671), .A(n14091), .ZN(n14092) );
  OAI21_X1 U17407 ( .B1(n14093), .B2(n16035), .A(n14092), .ZN(P1_U2991) );
  OAI21_X1 U17408 ( .B1(n14094), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n14095), .ZN(n14114) );
  XOR2_X1 U17409 ( .A(n14097), .B(n9597), .Z(n14112) );
  NOR2_X1 U17410 ( .A1(n18983), .A2(n16305), .ZN(n14104) );
  NAND3_X1 U17411 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14170) );
  AOI21_X1 U17412 ( .B1(n15611), .B2(n14170), .A(n14168), .ZN(n14102) );
  NOR3_X1 U17413 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14170), .A3(
        n14098), .ZN(n14169) );
  INV_X1 U17414 ( .A(n14099), .ZN(n14110) );
  NOR2_X1 U17415 ( .A1(n16315), .A2(n14110), .ZN(n14100) );
  AOI211_X1 U17416 ( .C1(P2_REIP_REG_6__SCAN_IN), .C2(n13328), .A(n14169), .B(
        n14100), .ZN(n14101) );
  OAI21_X1 U17417 ( .B1(n14102), .B2(n14166), .A(n14101), .ZN(n14103) );
  AOI211_X1 U17418 ( .C1(n14112), .C2(n16281), .A(n14104), .B(n14103), .ZN(
        n14105) );
  OAI21_X1 U17419 ( .B1(n16308), .B2(n14114), .A(n14105), .ZN(P2_U3040) );
  OAI22_X1 U17420 ( .A1(n14106), .A2(n19067), .B1(n19657), .B2(n18925), .ZN(
        n14107) );
  AOI21_X1 U17421 ( .B1(n19059), .B2(n14108), .A(n14107), .ZN(n14109) );
  OAI21_X1 U17422 ( .B1(n14110), .B2(n16272), .A(n14109), .ZN(n14111) );
  AOI21_X1 U17423 ( .B1(n14112), .B2(n16250), .A(n14111), .ZN(n14113) );
  OAI21_X1 U17424 ( .B1(n14114), .B2(n19075), .A(n14113), .ZN(P2_U3008) );
  OAI22_X1 U17425 ( .A1(n13145), .A2(n18935), .B1(n20772), .B2(n18927), .ZN(
        n14117) );
  NOR2_X1 U17426 ( .A1(n18954), .A2(n14115), .ZN(n14116) );
  AOI211_X1 U17427 ( .C1(n14118), .C2(n13145), .A(n14117), .B(n14116), .ZN(
        n14120) );
  NAND2_X1 U17428 ( .A1(n19727), .A2(n18901), .ZN(n14119) );
  OAI211_X1 U17429 ( .C1(n18936), .C2(n14121), .A(n14120), .B(n14119), .ZN(
        n14124) );
  NOR2_X1 U17430 ( .A1(n19732), .A2(n14122), .ZN(n14123) );
  AOI211_X1 U17431 ( .C1(n18902), .C2(n12141), .A(n14124), .B(n14123), .ZN(
        n14125) );
  OAI21_X1 U17432 ( .B1(n14126), .B2(n19628), .A(n14125), .ZN(P2_U2854) );
  NOR2_X1 U17433 ( .A1(n14128), .A2(n14129), .ZN(n14130) );
  OR2_X1 U17434 ( .A1(n14127), .A2(n14130), .ZN(n14735) );
  MUX2_X1 U17435 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n20020), .Z(
        n19937) );
  AOI22_X1 U17436 ( .A1(n14580), .A2(n19937), .B1(n16008), .B2(
        P1_EAX_REG_10__SCAN_IN), .ZN(n14131) );
  OAI21_X1 U17437 ( .B1(n14735), .B2(n15997), .A(n14131), .ZN(P1_U2894) );
  AND2_X1 U17438 ( .A1(n14143), .A2(n14132), .ZN(n14133) );
  OR2_X1 U17439 ( .A1(n14133), .A2(n14527), .ZN(n16121) );
  AOI22_X1 U17440 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19876), .B1(
        P1_EBX_REG_10__SCAN_IN), .B2(n19875), .ZN(n14135) );
  NAND2_X1 U17441 ( .A1(n19831), .A2(n14134), .ZN(n19864) );
  OAI211_X1 U17442 ( .C1(n16121), .C2(n19862), .A(n14135), .B(n19864), .ZN(
        n14138) );
  INV_X1 U17443 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n19846) );
  NAND4_X1 U17444 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_4__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n19834)
         );
  NAND2_X1 U17445 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19836) );
  NOR3_X1 U17446 ( .A1(n19846), .A2(n19834), .A3(n19836), .ZN(n19818) );
  NAND2_X1 U17447 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n19818), .ZN(n19806) );
  NOR2_X1 U17448 ( .A1(n20586), .A2(n19806), .ZN(n14449) );
  AOI21_X1 U17449 ( .B1(n19812), .B2(n14449), .A(P1_REIP_REG_10__SCAN_IN), 
        .ZN(n14136) );
  NAND2_X1 U17450 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n14449), .ZN(n14332) );
  NOR2_X1 U17451 ( .A1(n19805), .A2(n14332), .ZN(n14447) );
  INV_X1 U17452 ( .A(n19833), .ZN(n14446) );
  OR2_X1 U17453 ( .A1(n14447), .A2(n14446), .ZN(n15977) );
  OAI22_X1 U17454 ( .A1(n19892), .A2(n14731), .B1(n14136), .B2(n15977), .ZN(
        n14137) );
  NOR2_X1 U17455 ( .A1(n14138), .A2(n14137), .ZN(n14139) );
  OAI21_X1 U17456 ( .B1(n14735), .B2(n15982), .A(n14139), .ZN(P1_U2830) );
  AND2_X1 U17457 ( .A1(n14013), .A2(n14140), .ZN(n14141) );
  NOR2_X1 U17458 ( .A1(n14128), .A2(n14141), .ZN(n19814) );
  INV_X1 U17459 ( .A(n19814), .ZN(n14148) );
  AOI22_X1 U17460 ( .A1(n14580), .A2(n14549), .B1(n16008), .B2(
        P1_EAX_REG_9__SCAN_IN), .ZN(n14142) );
  OAI21_X1 U17461 ( .B1(n14148), .B2(n15997), .A(n14142), .ZN(P1_U2895) );
  INV_X1 U17462 ( .A(n14143), .ZN(n14144) );
  AOI21_X1 U17463 ( .B1(n14146), .B2(n14145), .A(n14144), .ZN(n19807) );
  AOI22_X1 U17464 ( .A1(n19807), .A2(n19894), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n14510), .ZN(n14147) );
  OAI21_X1 U17465 ( .B1(n14148), .B2(n14515), .A(n14147), .ZN(P1_U2863) );
  MUX2_X1 U17466 ( .A(n14150), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .S(
        n14844), .Z(n14151) );
  XNOR2_X1 U17467 ( .A(n14149), .B(n14151), .ZN(n16127) );
  INV_X1 U17468 ( .A(n19813), .ZN(n14153) );
  AOI22_X1 U17469 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n20014), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n14152) );
  OAI21_X1 U17470 ( .B1(n19972), .B2(n14153), .A(n14152), .ZN(n14154) );
  AOI21_X1 U17471 ( .B1(n19814), .B2(n14671), .A(n14154), .ZN(n14155) );
  OAI21_X1 U17472 ( .B1(n16127), .B2(n16035), .A(n14155), .ZN(P1_U2990) );
  INV_X1 U17473 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14156) );
  OAI222_X1 U17474 ( .A1(n16121), .A2(n14532), .B1(n19899), .B2(n14156), .C1(
        n14735), .C2(n14515), .ZN(P1_U2862) );
  XNOR2_X1 U17475 ( .A(n14158), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14159) );
  XNOR2_X1 U17476 ( .A(n14157), .B(n14159), .ZN(n14177) );
  NAND2_X1 U17477 ( .A1(n15433), .A2(n15432), .ZN(n14161) );
  XNOR2_X1 U17478 ( .A(n14160), .B(n14161), .ZN(n14175) );
  OAI22_X1 U17479 ( .A1(n19659), .A2(n18925), .B1(n16262), .B2(n14162), .ZN(
        n14164) );
  OAI22_X1 U17480 ( .A1(n16272), .A2(n14172), .B1(n9908), .B2(n19067), .ZN(
        n14163) );
  AOI211_X1 U17481 ( .C1(n14175), .C2(n16250), .A(n14164), .B(n14163), .ZN(
        n14165) );
  OAI21_X1 U17482 ( .B1(n14177), .B2(n19075), .A(n14165), .ZN(P2_U3007) );
  NOR2_X1 U17483 ( .A1(n14166), .A2(n14170), .ZN(n15459) );
  NAND2_X1 U17484 ( .A1(n15459), .A2(n14167), .ZN(n15752) );
  AOI211_X1 U17485 ( .C1(n15611), .C2(n14170), .A(n14169), .B(n14168), .ZN(
        n15754) );
  NAND2_X1 U17486 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n13328), .ZN(n14171) );
  OAI221_X1 U17487 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15752), .C1(
        n9951), .C2(n15754), .A(n14171), .ZN(n14174) );
  OAI22_X1 U17488 ( .A1(n18982), .A2(n16305), .B1(n16315), .B2(n14172), .ZN(
        n14173) );
  AOI211_X1 U17489 ( .C1(n14175), .C2(n16281), .A(n14174), .B(n14173), .ZN(
        n14176) );
  OAI21_X1 U17490 ( .B1(n14177), .B2(n16308), .A(n14176), .ZN(P2_U3039) );
  AND2_X1 U17491 ( .A1(n14179), .A2(n14178), .ZN(n14180) );
  NOR2_X1 U17492 ( .A1(n14189), .A2(n14180), .ZN(n15647) );
  INV_X1 U17493 ( .A(n15647), .ZN(n15028) );
  INV_X1 U17494 ( .A(n14182), .ZN(n14183) );
  AOI21_X1 U17495 ( .B1(n14184), .B2(n14049), .A(n14183), .ZN(n15208) );
  NAND2_X1 U17496 ( .A1(n15208), .A2(n15119), .ZN(n14186) );
  NAND2_X1 U17497 ( .A1(n15122), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n14185) );
  OAI211_X1 U17498 ( .C1(n15028), .C2(n15122), .A(n14186), .B(n14185), .ZN(
        P2_U2870) );
  OR2_X1 U17499 ( .A1(n14189), .A2(n14188), .ZN(n14190) );
  NAND2_X1 U17500 ( .A1(n14187), .A2(n14190), .ZN(n18872) );
  AOI21_X1 U17501 ( .B1(n14192), .B2(n14182), .A(n14191), .ZN(n15202) );
  NAND2_X1 U17502 ( .A1(n15202), .A2(n15119), .ZN(n14194) );
  NAND2_X1 U17503 ( .A1(n15122), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n14193) );
  OAI211_X1 U17504 ( .C1(n18872), .C2(n15122), .A(n14194), .B(n14193), .ZN(
        P2_U2869) );
  NAND2_X1 U17505 ( .A1(n14187), .A2(n14196), .ZN(n14197) );
  OR2_X1 U17506 ( .A1(n14191), .A2(n14199), .ZN(n14200) );
  AND2_X1 U17507 ( .A1(n14198), .A2(n14200), .ZN(n16237) );
  NAND2_X1 U17508 ( .A1(n16237), .A2(n15119), .ZN(n14202) );
  NAND2_X1 U17509 ( .A1(n15122), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n14201) );
  OAI211_X1 U17510 ( .C1(n15015), .C2(n15122), .A(n14202), .B(n14201), .ZN(
        P2_U2868) );
  INV_X1 U17511 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16794) );
  INV_X1 U17512 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n14209) );
  INV_X1 U17513 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16812) );
  NOR3_X1 U17514 ( .A1(n16794), .A2(n14209), .A3(n16812), .ZN(n14219) );
  NOR2_X1 U17515 ( .A1(n18204), .A2(n14203), .ZN(n14206) );
  INV_X1 U17516 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n16854) );
  INV_X1 U17517 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n20773) );
  INV_X1 U17518 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17189) );
  NOR2_X1 U17519 ( .A1(n20773), .A2(n17189), .ZN(n17184) );
  INV_X1 U17520 ( .A(n17184), .ZN(n16867) );
  NOR2_X1 U17521 ( .A1(n16854), .A2(n16867), .ZN(n17182) );
  NAND3_X1 U17522 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17195), .A3(n17182), .ZN(
        n14217) );
  INV_X1 U17523 ( .A(n14217), .ZN(n17180) );
  NAND2_X1 U17524 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17180), .ZN(n17179) );
  INV_X1 U17525 ( .A(n17179), .ZN(n17177) );
  NOR2_X1 U17526 ( .A1(n14209), .A2(n16812), .ZN(n14210) );
  NOR2_X1 U17527 ( .A1(n18204), .A2(n17179), .ZN(n17174) );
  AOI21_X1 U17528 ( .B1(n14210), .B2(n17174), .A(P3_EBX_REG_7__SCAN_IN), .ZN(
        n14211) );
  NOR2_X1 U17529 ( .A1(n17171), .A2(n14211), .ZN(n14212) );
  MUX2_X1 U17530 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B(n14212), .S(n17188), 
        .Z(P3_U2696) );
  OAI211_X1 U17531 ( .C1(n18612), .C2(n20789), .A(n9674), .B(n16821), .ZN(
        n18148) );
  NOR2_X1 U17532 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18148), .ZN(n14213) );
  NOR3_X1 U17533 ( .A1(n18763), .A2(n18808), .A3(n18820), .ZN(n18664) );
  INV_X1 U17534 ( .A(n18664), .ZN(n18751) );
  NAND2_X1 U17535 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18147) );
  NAND2_X1 U17536 ( .A1(n16821), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18765) );
  OAI21_X1 U17537 ( .B1(n14213), .B2(n18751), .A(n18509), .ZN(n18151) );
  INV_X1 U17538 ( .A(n18151), .ZN(n18155) );
  NOR2_X1 U17539 ( .A1(n18763), .A2(n16515), .ZN(n17762) );
  NAND2_X1 U17540 ( .A1(n18752), .A2(n18147), .ZN(n18811) );
  NOR2_X1 U17541 ( .A1(n17762), .A2(n18811), .ZN(n15771) );
  AOI21_X1 U17542 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15771), .ZN(n15772) );
  NOR2_X1 U17543 ( .A1(n18155), .A2(n15772), .ZN(n14215) );
  NAND3_X1 U17544 ( .A1(n18820), .A2(n18752), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18411) );
  INV_X1 U17545 ( .A(n18411), .ZN(n15774) );
  NOR2_X1 U17546 ( .A1(n18752), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18209) );
  OR2_X1 U17547 ( .A1(n18209), .A2(n18155), .ZN(n15770) );
  OR2_X1 U17548 ( .A1(n15774), .A2(n15770), .ZN(n14214) );
  MUX2_X1 U17549 ( .A(n14215), .B(n14214), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  AND2_X1 U17550 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16924) );
  NAND2_X1 U17551 ( .A1(n17120), .A2(n17195), .ZN(n17190) );
  INV_X1 U17552 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n16884) );
  NAND3_X1 U17553 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_12__SCAN_IN), .ZN(n17071) );
  NAND4_X1 U17554 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(P3_EBX_REG_8__SCAN_IN), .A4(P3_EBX_REG_4__SCAN_IN), .ZN(n14216) );
  NOR3_X1 U17555 ( .A1(n14217), .A2(n17071), .A3(n14216), .ZN(n14218) );
  NAND4_X1 U17556 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(n14219), .A4(n14218), .ZN(n17057) );
  INV_X1 U17557 ( .A(n17057), .ZN(n17031) );
  NAND2_X1 U17558 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17017), .ZN(n17003) );
  NOR2_X1 U17559 ( .A1(n18204), .A2(n17003), .ZN(n16991) );
  NAND3_X1 U17560 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n16977), .ZN(n16950) );
  NAND2_X1 U17561 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n16945), .ZN(n16930) );
  INV_X1 U17562 ( .A(n16930), .ZN(n16940) );
  NAND2_X1 U17563 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16940), .ZN(n16935) );
  NAND2_X1 U17564 ( .A1(n17188), .A2(n16935), .ZN(n14220) );
  OAI21_X1 U17565 ( .B1(n16924), .B2(n17190), .A(n14220), .ZN(n16925) );
  AOI22_X1 U17566 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14224) );
  AOI22_X1 U17567 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14223) );
  AOI22_X1 U17568 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14222) );
  AOI22_X1 U17569 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17079), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14221) );
  NAND4_X1 U17570 ( .A1(n14224), .A2(n14223), .A3(n14222), .A4(n14221), .ZN(
        n14230) );
  AOI22_X1 U17571 ( .A1(n14241), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14228) );
  AOI22_X1 U17572 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14227) );
  AOI22_X1 U17573 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14226) );
  AOI22_X1 U17574 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14225) );
  NAND4_X1 U17575 ( .A1(n14228), .A2(n14227), .A3(n14226), .A4(n14225), .ZN(
        n14229) );
  NOR2_X1 U17576 ( .A1(n14230), .A2(n14229), .ZN(n14295) );
  AOI22_X1 U17577 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14234) );
  AOI22_X1 U17578 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14233) );
  AOI22_X1 U17579 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14232) );
  AOI22_X1 U17580 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14231) );
  NAND4_X1 U17581 ( .A1(n14234), .A2(n14233), .A3(n14232), .A4(n14231), .ZN(
        n14240) );
  AOI22_X1 U17582 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14238) );
  AOI22_X1 U17583 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14237) );
  AOI22_X1 U17584 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14236) );
  AOI22_X1 U17585 ( .A1(n14241), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17079), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14235) );
  NAND4_X1 U17586 ( .A1(n14238), .A2(n14237), .A3(n14236), .A4(n14235), .ZN(
        n14239) );
  NOR2_X1 U17587 ( .A1(n14240), .A2(n14239), .ZN(n16933) );
  AOI22_X1 U17588 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n14241), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17079), .ZN(n14245) );
  AOI22_X1 U17589 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10280), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14244) );
  AOI22_X1 U17590 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n9591), .ZN(n14243) );
  AOI22_X1 U17591 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10141), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n9595), .ZN(n14242) );
  NAND4_X1 U17592 ( .A1(n14245), .A2(n14244), .A3(n14243), .A4(n14242), .ZN(
        n14251) );
  AOI22_X1 U17593 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17159), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14249) );
  AOI22_X1 U17594 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14248) );
  AOI22_X1 U17595 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14247) );
  AOI22_X1 U17596 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17156), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14246) );
  NAND4_X1 U17597 ( .A1(n14249), .A2(n14248), .A3(n14247), .A4(n14246), .ZN(
        n14250) );
  NOR2_X1 U17598 ( .A1(n14251), .A2(n14250), .ZN(n16942) );
  AOI22_X1 U17599 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17018), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14261) );
  AOI22_X1 U17600 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14260) );
  AOI22_X1 U17601 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14252) );
  OAI21_X1 U17602 ( .B1(n14284), .B2(n18164), .A(n14252), .ZN(n14258) );
  AOI22_X1 U17603 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14256) );
  AOI22_X1 U17604 ( .A1(n17079), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14255) );
  AOI22_X1 U17605 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14254) );
  AOI22_X1 U17606 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14253) );
  NAND4_X1 U17607 ( .A1(n14256), .A2(n14255), .A3(n14254), .A4(n14253), .ZN(
        n14257) );
  AOI211_X1 U17608 ( .C1(n14285), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n14258), .B(n14257), .ZN(n14259) );
  NAND3_X1 U17609 ( .A1(n14261), .A2(n14260), .A3(n14259), .ZN(n16947) );
  AOI22_X1 U17610 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14271) );
  AOI22_X1 U17611 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14270) );
  AOI22_X1 U17612 ( .A1(n17079), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14262) );
  OAI21_X1 U17613 ( .B1(n9674), .B2(n20823), .A(n14262), .ZN(n14268) );
  AOI22_X1 U17614 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14266) );
  AOI22_X1 U17615 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14265) );
  AOI22_X1 U17616 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14264) );
  AOI22_X1 U17617 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14263) );
  NAND4_X1 U17618 ( .A1(n14266), .A2(n14265), .A3(n14264), .A4(n14263), .ZN(
        n14267) );
  AOI211_X1 U17619 ( .C1(n17157), .C2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A(
        n14268), .B(n14267), .ZN(n14269) );
  NAND3_X1 U17620 ( .A1(n14271), .A2(n14270), .A3(n14269), .ZN(n16948) );
  NAND2_X1 U17621 ( .A1(n16947), .A2(n16948), .ZN(n16946) );
  NOR2_X1 U17622 ( .A1(n16942), .A2(n16946), .ZN(n16941) );
  AOI22_X1 U17623 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14281) );
  AOI22_X1 U17624 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14280) );
  AOI22_X1 U17625 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14272) );
  OAI21_X1 U17626 ( .B1(n14284), .B2(n18176), .A(n14272), .ZN(n14278) );
  AOI22_X1 U17627 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14276) );
  AOI22_X1 U17628 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14275) );
  AOI22_X1 U17629 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14274) );
  AOI22_X1 U17630 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17079), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14273) );
  NAND4_X1 U17631 ( .A1(n14276), .A2(n14275), .A3(n14274), .A4(n14273), .ZN(
        n14277) );
  AOI211_X1 U17632 ( .C1(n17158), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n14278), .B(n14277), .ZN(n14279) );
  NAND3_X1 U17633 ( .A1(n14281), .A2(n14280), .A3(n14279), .ZN(n16938) );
  NAND2_X1 U17634 ( .A1(n16941), .A2(n16938), .ZN(n16937) );
  NOR2_X1 U17635 ( .A1(n16933), .A2(n16937), .ZN(n16932) );
  AOI22_X1 U17636 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14294) );
  AOI22_X1 U17637 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14293) );
  AOI22_X1 U17638 ( .A1(n17079), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14283) );
  OAI21_X1 U17639 ( .B1(n14284), .B2(n18188), .A(n14283), .ZN(n14291) );
  AOI22_X1 U17640 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14289) );
  AOI22_X1 U17641 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14288) );
  AOI22_X1 U17642 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14287) );
  AOI22_X1 U17643 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14286) );
  NAND4_X1 U17644 ( .A1(n14289), .A2(n14288), .A3(n14287), .A4(n14286), .ZN(
        n14290) );
  AOI211_X1 U17645 ( .C1(n17081), .C2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n14291), .B(n14290), .ZN(n14292) );
  NAND3_X1 U17646 ( .A1(n14294), .A2(n14293), .A3(n14292), .ZN(n16928) );
  NAND2_X1 U17647 ( .A1(n16932), .A2(n16928), .ZN(n16927) );
  NOR2_X1 U17648 ( .A1(n14295), .A2(n16927), .ZN(n16922) );
  AOI21_X1 U17649 ( .B1(n14295), .B2(n16927), .A(n16922), .ZN(n17213) );
  AOI22_X1 U17650 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16925), .B1(n17213), 
        .B2(n17193), .ZN(n14299) );
  INV_X1 U17651 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n14297) );
  INV_X1 U17652 ( .A(n16935), .ZN(n14296) );
  NAND3_X1 U17653 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n14297), .A3(n14296), 
        .ZN(n14298) );
  NAND2_X1 U17654 ( .A1(n14299), .A2(n14298), .ZN(P3_U2675) );
  AOI22_X1 U17655 ( .A1(n14301), .A2(n15814), .B1(P1_FLUSH_REG_SCAN_IN), .B2(
        n14300), .ZN(n16160) );
  OAI21_X1 U17656 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n20389), .A(n16160), 
        .ZN(n16157) );
  INV_X1 U17657 ( .A(n16157), .ZN(n20637) );
  AOI21_X1 U17658 ( .B1(n14880), .B2(n14877), .A(n20637), .ZN(n14305) );
  OAI22_X1 U17659 ( .A1(n20125), .A2(n14879), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14302), .ZN(n15811) );
  OAI22_X1 U17660 ( .A1(n20555), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20633), .ZN(n14303) );
  AOI21_X1 U17661 ( .B1(n15811), .B2(n14880), .A(n14303), .ZN(n14304) );
  OAI22_X1 U17662 ( .A1(n14305), .A2(n11226), .B1(n14304), .B2(n20637), .ZN(
        P1_U3474) );
  AOI22_X1 U17663 ( .A1(n11148), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n14307) );
  NAND2_X1 U17664 ( .A1(n15046), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14306) );
  OAI211_X1 U17665 ( .C1(n11121), .C2(n15480), .A(n14307), .B(n14306), .ZN(
        n15043) );
  NOR2_X1 U17666 ( .A1(n15235), .A2(n13198), .ZN(n14308) );
  AOI21_X1 U17667 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n13198), .A(n14308), .ZN(
        n14309) );
  OAI21_X1 U17668 ( .B1(n14310), .B2(n15114), .A(n14309), .ZN(P2_U2857) );
  NAND2_X1 U17669 ( .A1(n14312), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14313) );
  NAND2_X1 U17670 ( .A1(n14314), .A2(n14313), .ZN(n14315) );
  XNOR2_X1 U17671 ( .A(n14315), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14744) );
  INV_X1 U17672 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20624) );
  NOR2_X1 U17673 ( .A1(n16122), .A2(n20624), .ZN(n14740) );
  AOI21_X1 U17674 ( .B1(n19962), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14740), .ZN(n14316) );
  OAI21_X1 U17675 ( .B1(n14317), .B2(n19972), .A(n14316), .ZN(n14318) );
  OAI21_X1 U17676 ( .B1(n14744), .B2(n16035), .A(n14319), .ZN(P1_U2968) );
  INV_X1 U17677 ( .A(n14586), .ZN(n14537) );
  INV_X1 U17678 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14345) );
  INV_X1 U17679 ( .A(n14321), .ZN(n14322) );
  AOI22_X1 U17680 ( .A1(n14327), .A2(n12921), .B1(n14322), .B2(n14362), .ZN(
        n14323) );
  AOI22_X1 U17681 ( .A1(n12943), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n13285), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14328) );
  OAI222_X1 U17682 ( .A1(n14515), .A2(n14537), .B1(n14345), .B2(n19899), .C1(
        n14745), .C2(n14532), .ZN(P1_U2842) );
  NAND2_X1 U17683 ( .A1(n14324), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n14326)
         );
  NAND3_X1 U17684 ( .A1(n14326), .A2(n14325), .A3(n19783), .ZN(P1_U2801) );
  MUX2_X1 U17685 ( .A(n14328), .B(n12939), .S(n14327), .Z(n14330) );
  AOI22_X1 U17686 ( .A1(n12943), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n13285), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14329) );
  XNOR2_X2 U17687 ( .A(n14330), .B(n14329), .ZN(n14738) );
  NAND2_X1 U17688 ( .A1(n14331), .A2(n19857), .ZN(n14340) );
  INV_X1 U17689 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14344) );
  NOR2_X1 U17690 ( .A1(n20620), .A2(n14344), .ZN(n14335) );
  INV_X1 U17691 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20615) );
  INV_X1 U17692 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20604) );
  NAND4_X1 U17693 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(P1_REIP_REG_12__SCAN_IN), .A4(P1_REIP_REG_11__SCAN_IN), .ZN(n15904) );
  NOR2_X1 U17694 ( .A1(n14332), .A2(n15904), .ZN(n15917) );
  INV_X1 U17695 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20602) );
  INV_X1 U17696 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20599) );
  NAND3_X1 U17697 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n15918) );
  NOR3_X1 U17698 ( .A1(n20602), .A2(n20599), .A3(n15918), .ZN(n15905) );
  NAND3_X1 U17699 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n15917), .A3(n15905), 
        .ZN(n15890) );
  NOR2_X1 U17700 ( .A1(n20604), .A2(n15890), .ZN(n15883) );
  NAND2_X1 U17701 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n15883), .ZN(n14434) );
  INV_X1 U17702 ( .A(n14434), .ZN(n14333) );
  AND2_X1 U17703 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n14333), .ZN(n14423) );
  NAND2_X1 U17704 ( .A1(n14423), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14381) );
  NAND2_X1 U17705 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14383) );
  NOR2_X1 U17706 ( .A1(n14381), .A2(n14383), .ZN(n14379) );
  NAND2_X1 U17707 ( .A1(n14379), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14364) );
  NOR2_X1 U17708 ( .A1(n20615), .A2(n14364), .ZN(n14365) );
  NAND2_X1 U17709 ( .A1(n19831), .A2(n14365), .ZN(n14334) );
  NAND2_X1 U17710 ( .A1(n19833), .A2(n14334), .ZN(n14370) );
  OAI21_X1 U17711 ( .B1(n14335), .B2(n19835), .A(n14370), .ZN(n14341) );
  INV_X1 U17712 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14459) );
  OAI22_X1 U17713 ( .A1(n19821), .A2(n14459), .B1(n14336), .B2(n19867), .ZN(
        n14338) );
  NAND3_X1 U17714 ( .A1(n19812), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n14365), 
        .ZN(n14343) );
  NOR3_X1 U17715 ( .A1(n14343), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14344), 
        .ZN(n14337) );
  AOI211_X1 U17716 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14341), .A(n14338), 
        .B(n14337), .ZN(n14339) );
  OAI211_X1 U17717 ( .C1(n14738), .C2(n19862), .A(n14340), .B(n14339), .ZN(
        P1_U2809) );
  NAND2_X1 U17718 ( .A1(n14586), .A2(n19857), .ZN(n14349) );
  INV_X1 U17719 ( .A(n14341), .ZN(n14342) );
  AOI21_X1 U17720 ( .B1(n14344), .B2(n14343), .A(n14342), .ZN(n14347) );
  OAI22_X1 U17721 ( .A1(n19821), .A2(n14345), .B1(n14584), .B2(n19867), .ZN(
        n14346) );
  AOI211_X1 U17722 ( .C1(n19852), .C2(n14582), .A(n14347), .B(n14346), .ZN(
        n14348) );
  OAI211_X1 U17723 ( .C1(n19862), .C2(n14745), .A(n14349), .B(n14348), .ZN(
        P1_U2810) );
  AOI21_X1 U17724 ( .B1(n14351), .B2(n14361), .A(n9646), .ZN(n14591) );
  NAND2_X1 U17725 ( .A1(n14591), .A2(n19857), .ZN(n14359) );
  INV_X1 U17726 ( .A(n14589), .ZN(n14357) );
  INV_X1 U17727 ( .A(n14365), .ZN(n14352) );
  NOR2_X1 U17728 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(n14352), .ZN(n14353) );
  AOI22_X1 U17729 ( .A1(n19812), .A2(n14353), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19876), .ZN(n14355) );
  NAND2_X1 U17730 ( .A1(n19875), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14354) );
  OAI211_X1 U17731 ( .C1(n14370), .C2(n20620), .A(n14355), .B(n14354), .ZN(
        n14356) );
  AOI21_X1 U17732 ( .B1(n19852), .B2(n14357), .A(n14356), .ZN(n14358) );
  OAI211_X1 U17733 ( .C1(n19862), .C2(n14460), .A(n14359), .B(n14358), .ZN(
        P1_U2811) );
  AOI21_X1 U17734 ( .B1(n14363), .B2(n14378), .A(n14362), .ZN(n14762) );
  NAND2_X1 U17735 ( .A1(n19852), .A2(n14605), .ZN(n14369) );
  NOR2_X1 U17736 ( .A1(n19867), .A2(n14602), .ZN(n14367) );
  NOR3_X1 U17737 ( .A1(n19835), .A2(n14365), .A3(n14364), .ZN(n14366) );
  AOI211_X1 U17738 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n19875), .A(n14367), .B(
        n14366), .ZN(n14368) );
  OAI211_X1 U17739 ( .C1(n14370), .C2(n20615), .A(n14369), .B(n14368), .ZN(
        n14371) );
  AOI21_X1 U17740 ( .B1(n14762), .B2(n19884), .A(n14371), .ZN(n14372) );
  OAI21_X1 U17741 ( .B1(n14603), .B2(n15982), .A(n14372), .ZN(P1_U2812) );
  AOI21_X1 U17742 ( .B1(n14375), .B2(n14373), .A(n14374), .ZN(n14614) );
  INV_X1 U17743 ( .A(n14614), .ZN(n14545) );
  NAND2_X1 U17744 ( .A1(n14392), .A2(n14376), .ZN(n14377) );
  NAND2_X1 U17745 ( .A1(n14378), .A2(n14377), .ZN(n14463) );
  INV_X1 U17746 ( .A(n14463), .ZN(n14772) );
  OAI21_X1 U17747 ( .B1(n19835), .B2(n14379), .A(n19831), .ZN(n14394) );
  INV_X1 U17748 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14464) );
  OAI22_X1 U17749 ( .A1(n19821), .A2(n14464), .B1(n14380), .B2(n19867), .ZN(
        n14385) );
  INV_X1 U17750 ( .A(n14381), .ZN(n14382) );
  NAND2_X1 U17751 ( .A1(n19812), .A2(n14382), .ZN(n14411) );
  NOR3_X1 U17752 ( .A1(n14411), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14383), 
        .ZN(n14384) );
  AOI211_X1 U17753 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n14394), .A(n14385), 
        .B(n14384), .ZN(n14386) );
  OAI21_X1 U17754 ( .B1(n19892), .B2(n14612), .A(n14386), .ZN(n14387) );
  AOI21_X1 U17755 ( .B1(n14772), .B2(n19884), .A(n14387), .ZN(n14388) );
  OAI21_X1 U17756 ( .B1(n14545), .B2(n15982), .A(n14388), .ZN(P1_U2813) );
  INV_X1 U17757 ( .A(n14373), .ZN(n14390) );
  AOI21_X1 U17758 ( .B1(n14391), .B2(n14406), .A(n14390), .ZN(n14623) );
  INV_X1 U17759 ( .A(n14623), .ZN(n14548) );
  AOI21_X1 U17760 ( .B1(n14393), .B2(n14403), .A(n9912), .ZN(n14783) );
  INV_X1 U17761 ( .A(n14619), .ZN(n14398) );
  AOI22_X1 U17762 ( .A1(n19875), .A2(P1_EBX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n19876), .ZN(n14397) );
  INV_X1 U17763 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20610) );
  NOR2_X1 U17764 ( .A1(n14411), .A2(n20610), .ZN(n14395) );
  OAI21_X1 U17765 ( .B1(n14395), .B2(P1_REIP_REG_26__SCAN_IN), .A(n14394), 
        .ZN(n14396) );
  OAI211_X1 U17766 ( .C1(n19892), .C2(n14398), .A(n14397), .B(n14396), .ZN(
        n14399) );
  AOI21_X1 U17767 ( .B1(n14783), .B2(n19884), .A(n14399), .ZN(n14400) );
  OAI21_X1 U17768 ( .B1(n14548), .B2(n15982), .A(n14400), .ZN(P1_U2814) );
  OR2_X1 U17769 ( .A1(n14419), .A2(n14401), .ZN(n14402) );
  NAND2_X1 U17770 ( .A1(n14403), .A2(n14402), .ZN(n14791) );
  AOI21_X1 U17772 ( .B1(n14407), .B2(n14405), .A(n14389), .ZN(n14632) );
  NAND2_X1 U17773 ( .A1(n14632), .A2(n19857), .ZN(n14415) );
  INV_X1 U17774 ( .A(n14630), .ZN(n14413) );
  OAI21_X1 U17775 ( .B1(n19835), .B2(n14423), .A(n19831), .ZN(n14435) );
  NOR2_X1 U17776 ( .A1(n19835), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14408) );
  OAI21_X1 U17777 ( .B1(n14435), .B2(n14408), .A(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14410) );
  AOI22_X1 U17778 ( .A1(n19875), .A2(P1_EBX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n19876), .ZN(n14409) );
  OAI211_X1 U17779 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14411), .A(n14410), 
        .B(n14409), .ZN(n14412) );
  AOI21_X1 U17780 ( .B1(n19852), .B2(n14413), .A(n14412), .ZN(n14414) );
  OAI211_X1 U17781 ( .C1(n19862), .C2(n14791), .A(n14415), .B(n14414), .ZN(
        P1_U2815) );
  OAI21_X1 U17782 ( .B1(n14416), .B2(n14417), .A(n14405), .ZN(n14638) );
  INV_X1 U17783 ( .A(n14418), .ZN(n14421) );
  INV_X1 U17784 ( .A(n14432), .ZN(n14420) );
  AOI21_X1 U17785 ( .B1(n14421), .B2(n14420), .A(n14419), .ZN(n14804) );
  INV_X1 U17786 ( .A(n14641), .ZN(n14428) );
  INV_X1 U17787 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14637) );
  INV_X1 U17788 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n14422) );
  NAND3_X1 U17789 ( .A1(n19812), .A2(n14423), .A3(n14422), .ZN(n14425) );
  NAND2_X1 U17790 ( .A1(n19875), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n14424) );
  OAI211_X1 U17791 ( .C1(n19867), .C2(n14637), .A(n14425), .B(n14424), .ZN(
        n14426) );
  AOI21_X1 U17792 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n14435), .A(n14426), 
        .ZN(n14427) );
  OAI21_X1 U17793 ( .B1(n19892), .B2(n14428), .A(n14427), .ZN(n14429) );
  AOI21_X1 U17794 ( .B1(n14804), .B2(n19884), .A(n14429), .ZN(n14430) );
  OAI21_X1 U17795 ( .B1(n14638), .B2(n15982), .A(n14430), .ZN(P1_U2816) );
  AOI21_X1 U17796 ( .B1(n14431), .B2(n9677), .A(n14416), .ZN(n14647) );
  INV_X1 U17797 ( .A(n14647), .ZN(n14558) );
  AOI21_X1 U17798 ( .B1(n14433), .B2(n14474), .A(n14432), .ZN(n14812) );
  AOI22_X1 U17799 ( .A1(n19875), .A2(P1_EBX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19876), .ZN(n14438) );
  NOR2_X1 U17800 ( .A1(n19835), .A2(n14434), .ZN(n14436) );
  OAI21_X1 U17801 ( .B1(n14436), .B2(P1_REIP_REG_23__SCAN_IN), .A(n14435), 
        .ZN(n14437) );
  OAI211_X1 U17802 ( .C1(n19892), .C2(n14645), .A(n14438), .B(n14437), .ZN(
        n14439) );
  AOI21_X1 U17803 ( .B1(n14812), .B2(n19884), .A(n14439), .ZN(n14440) );
  OAI21_X1 U17804 ( .B1(n14558), .B2(n15982), .A(n14440), .ZN(P1_U2817) );
  OR2_X1 U17805 ( .A1(n14127), .A2(n14442), .ZN(n14443) );
  NAND2_X1 U17806 ( .A1(n14441), .A2(n14443), .ZN(n14525) );
  OAI21_X1 U17807 ( .B1(n14525), .B2(n9978), .A(n14441), .ZN(n14517) );
  AND2_X1 U17808 ( .A1(n14517), .A2(n14516), .ZN(n14519) );
  OAI21_X1 U17809 ( .B1(n14519), .B2(n14445), .A(n14444), .ZN(n14728) );
  NAND2_X1 U17810 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14450) );
  INV_X1 U17811 ( .A(n14450), .ZN(n14448) );
  AOI21_X1 U17812 ( .B1(n14448), .B2(n14447), .A(n14446), .ZN(n15973) );
  NAND3_X1 U17813 ( .A1(n19812), .A2(P1_REIP_REG_10__SCAN_IN), .A3(n14449), 
        .ZN(n15986) );
  NOR2_X1 U17814 ( .A1(n14450), .A2(n15986), .ZN(n15958) );
  INV_X1 U17815 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20592) );
  NAND2_X1 U17816 ( .A1(n14451), .A2(n14452), .ZN(n14453) );
  AND2_X1 U17817 ( .A1(n14509), .A2(n14453), .ZN(n16086) );
  AOI22_X1 U17818 ( .A1(P1_EBX_REG_13__SCAN_IN), .A2(n19875), .B1(n19884), 
        .B2(n16086), .ZN(n14454) );
  OAI211_X1 U17819 ( .C1(n19867), .C2(n14455), .A(n14454), .B(n19864), .ZN(
        n14456) );
  AOI221_X1 U17820 ( .B1(n15973), .B2(P1_REIP_REG_13__SCAN_IN), .C1(n15958), 
        .C2(n20592), .A(n14456), .ZN(n14458) );
  NAND2_X1 U17821 ( .A1(n19852), .A2(n14725), .ZN(n14457) );
  OAI211_X1 U17822 ( .C1(n14728), .C2(n15982), .A(n14458), .B(n14457), .ZN(
        P1_U2827) );
  OAI22_X1 U17823 ( .A1(n14738), .A2(n14532), .B1(n19899), .B2(n14459), .ZN(
        P1_U2841) );
  INV_X1 U17824 ( .A(n14591), .ZN(n14540) );
  OAI222_X1 U17825 ( .A1(n14515), .A2(n14540), .B1(n14461), .B2(n19899), .C1(
        n14460), .C2(n14532), .ZN(P1_U2843) );
  AOI22_X1 U17826 ( .A1(n14762), .A2(n19894), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n14510), .ZN(n14462) );
  OAI21_X1 U17827 ( .B1(n14603), .B2(n14515), .A(n14462), .ZN(P1_U2844) );
  OAI222_X1 U17828 ( .A1(n14515), .A2(n14545), .B1(n14464), .B2(n19899), .C1(
        n14463), .C2(n14532), .ZN(P1_U2845) );
  AOI22_X1 U17829 ( .A1(n14783), .A2(n19894), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n14510), .ZN(n14465) );
  OAI21_X1 U17830 ( .B1(n14548), .B2(n14515), .A(n14465), .ZN(P1_U2846) );
  INV_X1 U17831 ( .A(n14632), .ZN(n14552) );
  INV_X1 U17832 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n20754) );
  OAI222_X1 U17833 ( .A1(n14515), .A2(n14552), .B1(n20754), .B2(n19899), .C1(
        n14791), .C2(n14532), .ZN(P1_U2847) );
  INV_X1 U17834 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14467) );
  INV_X1 U17835 ( .A(n14804), .ZN(n14466) );
  OAI222_X1 U17836 ( .A1(n14515), .A2(n14638), .B1(n19899), .B2(n14467), .C1(
        n14466), .C2(n14532), .ZN(P1_U2848) );
  AOI22_X1 U17837 ( .A1(n14812), .A2(n19894), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n14510), .ZN(n14468) );
  OAI21_X1 U17838 ( .B1(n14558), .B2(n14515), .A(n14468), .ZN(P1_U2849) );
  NAND2_X1 U17839 ( .A1(n14469), .A2(n14470), .ZN(n14471) );
  NAND2_X1 U17840 ( .A1(n14823), .A2(n14472), .ZN(n14473) );
  NAND2_X1 U17841 ( .A1(n14474), .A2(n14473), .ZN(n15893) );
  OAI22_X1 U17842 ( .A1(n15893), .A2(n14532), .B1(n15887), .B2(n19899), .ZN(
        n14475) );
  INV_X1 U17843 ( .A(n14475), .ZN(n14476) );
  OAI21_X1 U17844 ( .B1(n14562), .B2(n14515), .A(n14476), .ZN(P1_U2850) );
  INV_X1 U17845 ( .A(n14478), .ZN(n14667) );
  OAI21_X1 U17846 ( .B1(n14479), .B2(n14477), .A(n14667), .ZN(n15909) );
  NOR2_X1 U17847 ( .A1(n14833), .A2(n14480), .ZN(n14481) );
  OR2_X1 U17848 ( .A1(n14825), .A2(n14481), .ZN(n15914) );
  OAI22_X1 U17849 ( .A1(n15914), .A2(n14532), .B1(n15902), .B2(n19899), .ZN(
        n14482) );
  INV_X1 U17850 ( .A(n14482), .ZN(n14483) );
  OAI21_X1 U17851 ( .B1(n15909), .B2(n14515), .A(n14483), .ZN(P1_U2852) );
  XNOR2_X1 U17852 ( .A(n14485), .B(n14486), .ZN(n15930) );
  INV_X1 U17853 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14489) );
  NAND2_X1 U17854 ( .A1(n14857), .A2(n14487), .ZN(n14488) );
  NAND2_X1 U17855 ( .A1(n14834), .A2(n14488), .ZN(n16060) );
  OAI222_X1 U17856 ( .A1(n15930), .A2(n14515), .B1(n14489), .B2(n19899), .C1(
        n14532), .C2(n16060), .ZN(P1_U2854) );
  AOI21_X1 U17857 ( .B1(n14492), .B2(n14490), .A(n14491), .ZN(n14702) );
  OR2_X1 U17858 ( .A1(n14503), .A2(n14493), .ZN(n14494) );
  NAND2_X1 U17859 ( .A1(n14859), .A2(n14494), .ZN(n16072) );
  OAI22_X1 U17860 ( .A1(n16072), .A2(n14532), .B1(n15946), .B2(n19899), .ZN(
        n14495) );
  AOI21_X1 U17861 ( .B1(n14702), .B2(n19895), .A(n14495), .ZN(n14496) );
  INV_X1 U17862 ( .A(n14496), .ZN(P1_U2856) );
  INV_X1 U17863 ( .A(n14490), .ZN(n14499) );
  AOI21_X1 U17864 ( .B1(n14500), .B2(n14498), .A(n14499), .ZN(n16022) );
  INV_X1 U17865 ( .A(n16022), .ZN(n14574) );
  INV_X1 U17866 ( .A(n14509), .ZN(n14502) );
  AOI21_X1 U17867 ( .B1(n14502), .B2(n14508), .A(n14501), .ZN(n14504) );
  NOR2_X1 U17868 ( .A1(n14504), .A2(n14503), .ZN(n15952) );
  AOI22_X1 U17869 ( .A1(n15952), .A2(n19894), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n14510), .ZN(n14505) );
  OAI21_X1 U17870 ( .B1(n14574), .B2(n14515), .A(n14505), .ZN(P1_U2857) );
  NAND2_X1 U17871 ( .A1(n14444), .A2(n14506), .ZN(n14507) );
  XNOR2_X1 U17872 ( .A(n14509), .B(n14508), .ZN(n16078) );
  AOI22_X1 U17873 ( .A1(n16078), .A2(n19894), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n14510), .ZN(n14511) );
  OAI21_X1 U17874 ( .B1(n14576), .B2(n14515), .A(n14511), .ZN(P1_U2858) );
  NOR2_X1 U17875 ( .A1(n19899), .A2(n14512), .ZN(n14513) );
  AOI21_X1 U17876 ( .B1(n16086), .B2(n19894), .A(n14513), .ZN(n14514) );
  OAI21_X1 U17877 ( .B1(n14728), .B2(n14515), .A(n14514), .ZN(P1_U2859) );
  NOR2_X1 U17878 ( .A1(n14517), .A2(n14516), .ZN(n14518) );
  INV_X1 U17879 ( .A(n15976), .ZN(n16030) );
  OR2_X1 U17880 ( .A1(n14528), .A2(n14520), .ZN(n14521) );
  NAND2_X1 U17881 ( .A1(n14451), .A2(n14521), .ZN(n16104) );
  OAI22_X1 U17882 ( .A1(n16104), .A2(n14532), .B1(n15969), .B2(n19899), .ZN(
        n14522) );
  AOI21_X1 U17883 ( .B1(n16030), .B2(n19895), .A(n14522), .ZN(n14523) );
  INV_X1 U17884 ( .A(n14523), .ZN(P1_U2860) );
  XNOR2_X1 U17885 ( .A(n14525), .B(n14524), .ZN(n16039) );
  INV_X1 U17886 ( .A(n16039), .ZN(n15981) );
  INV_X1 U17887 ( .A(n14526), .ZN(n14530) );
  INV_X1 U17888 ( .A(n14527), .ZN(n14529) );
  AOI21_X1 U17889 ( .B1(n14530), .B2(n14529), .A(n14528), .ZN(n16105) );
  INV_X1 U17890 ( .A(n16105), .ZN(n14531) );
  OAI222_X1 U17891 ( .A1(n15981), .A2(n14515), .B1(n14533), .B2(n19899), .C1(
        n14532), .C2(n14531), .ZN(P1_U2861) );
  AOI22_X1 U17892 ( .A1(n16011), .A2(DATAI_30_), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n16008), .ZN(n14536) );
  NOR3_X1 U17893 ( .A1(n16008), .A2(n9769), .A3(n12070), .ZN(n14534) );
  MUX2_X1 U17894 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n20020), .Z(
        n19943) );
  AOI22_X1 U17895 ( .A1(n16010), .A2(n19943), .B1(BUF1_REG_30__SCAN_IN), .B2(
        n14566), .ZN(n14535) );
  OAI211_X1 U17896 ( .C1(n14537), .C2(n15997), .A(n14536), .B(n14535), .ZN(
        P1_U2874) );
  AOI22_X1 U17897 ( .A1(n16011), .A2(DATAI_29_), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n16008), .ZN(n14539) );
  MUX2_X1 U17898 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n20020), .Z(
        n19941) );
  AOI22_X1 U17899 ( .A1(n16010), .A2(n19941), .B1(BUF1_REG_29__SCAN_IN), .B2(
        n14566), .ZN(n14538) );
  OAI211_X1 U17900 ( .C1(n14540), .C2(n15997), .A(n14539), .B(n14538), .ZN(
        P1_U2875) );
  AOI22_X1 U17901 ( .A1(n16011), .A2(DATAI_28_), .B1(P1_EAX_REG_28__SCAN_IN), 
        .B2(n16008), .ZN(n14542) );
  MUX2_X1 U17902 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n20020), .Z(
        n19939) );
  AOI22_X1 U17903 ( .A1(n16010), .A2(n19939), .B1(BUF1_REG_28__SCAN_IN), .B2(
        n14566), .ZN(n14541) );
  OAI211_X1 U17904 ( .C1(n14603), .C2(n15997), .A(n14542), .B(n14541), .ZN(
        P1_U2876) );
  AOI22_X1 U17905 ( .A1(n16011), .A2(DATAI_27_), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n16008), .ZN(n14544) );
  AOI22_X1 U17906 ( .A1(n16010), .A2(n14579), .B1(BUF1_REG_27__SCAN_IN), .B2(
        n14566), .ZN(n14543) );
  OAI211_X1 U17907 ( .C1(n14545), .C2(n15997), .A(n14544), .B(n14543), .ZN(
        P1_U2877) );
  AOI22_X1 U17908 ( .A1(n16011), .A2(DATAI_26_), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n16008), .ZN(n14547) );
  AOI22_X1 U17909 ( .A1(n16010), .A2(n19937), .B1(BUF1_REG_26__SCAN_IN), .B2(
        n14566), .ZN(n14546) );
  OAI211_X1 U17910 ( .C1(n14548), .C2(n15997), .A(n14547), .B(n14546), .ZN(
        P1_U2878) );
  AOI22_X1 U17911 ( .A1(n16011), .A2(DATAI_25_), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(n16008), .ZN(n14551) );
  AOI22_X1 U17912 ( .A1(n16010), .A2(n14549), .B1(BUF1_REG_25__SCAN_IN), .B2(
        n14566), .ZN(n14550) );
  OAI211_X1 U17913 ( .C1(n14552), .C2(n15997), .A(n14551), .B(n14550), .ZN(
        P1_U2879) );
  AOI22_X1 U17914 ( .A1(n16011), .A2(DATAI_24_), .B1(P1_EAX_REG_24__SCAN_IN), 
        .B2(n16008), .ZN(n14554) );
  AOI22_X1 U17915 ( .A1(n16010), .A2(n19935), .B1(n14566), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n14553) );
  OAI211_X1 U17916 ( .C1(n14638), .C2(n15997), .A(n14554), .B(n14553), .ZN(
        P1_U2880) );
  AOI22_X1 U17917 ( .A1(n16011), .A2(DATAI_23_), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n16008), .ZN(n14557) );
  AOI22_X1 U17918 ( .A1(n16010), .A2(n14555), .B1(n14566), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n14556) );
  OAI211_X1 U17919 ( .C1(n14558), .C2(n15997), .A(n14557), .B(n14556), .ZN(
        P1_U2881) );
  AOI22_X1 U17920 ( .A1(n16011), .A2(DATAI_22_), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n16008), .ZN(n14561) );
  AOI22_X1 U17921 ( .A1(n16010), .A2(n14559), .B1(n14566), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n14560) );
  OAI211_X1 U17922 ( .C1(n14562), .C2(n15997), .A(n14561), .B(n14560), .ZN(
        P1_U2882) );
  AOI22_X1 U17923 ( .A1(n16011), .A2(DATAI_20_), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n16008), .ZN(n14565) );
  AOI22_X1 U17924 ( .A1(n16010), .A2(n14563), .B1(n14566), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n14564) );
  OAI211_X1 U17925 ( .C1(n15909), .C2(n15997), .A(n14565), .B(n14564), .ZN(
        P1_U2884) );
  INV_X1 U17926 ( .A(n14702), .ZN(n15947) );
  AOI22_X1 U17927 ( .A1(n16011), .A2(DATAI_16_), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n16008), .ZN(n14569) );
  AOI22_X1 U17928 ( .A1(n16010), .A2(n14567), .B1(n14566), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n14568) );
  OAI211_X1 U17929 ( .C1(n15947), .C2(n15997), .A(n14569), .B(n14568), .ZN(
        P1_U2888) );
  OAI222_X1 U17930 ( .A1(n14574), .A2(n15997), .B1(n14573), .B2(n14572), .C1(
        n14571), .C2(n14570), .ZN(P1_U2889) );
  AOI22_X1 U17931 ( .A1(n14580), .A2(n19943), .B1(n16008), .B2(
        P1_EAX_REG_14__SCAN_IN), .ZN(n14575) );
  OAI21_X1 U17932 ( .B1(n14576), .B2(n15997), .A(n14575), .ZN(P1_U2890) );
  AOI22_X1 U17933 ( .A1(n14580), .A2(n19941), .B1(n16008), .B2(
        P1_EAX_REG_13__SCAN_IN), .ZN(n14577) );
  OAI21_X1 U17934 ( .B1(n14728), .B2(n15997), .A(n14577), .ZN(P1_U2891) );
  AOI22_X1 U17935 ( .A1(n14580), .A2(n19939), .B1(n16008), .B2(
        P1_EAX_REG_12__SCAN_IN), .ZN(n14578) );
  OAI21_X1 U17936 ( .B1(n15976), .B2(n15997), .A(n14578), .ZN(P1_U2892) );
  AOI22_X1 U17937 ( .A1(n14580), .A2(n14579), .B1(n16008), .B2(
        P1_EAX_REG_11__SCAN_IN), .ZN(n14581) );
  OAI21_X1 U17938 ( .B1(n15981), .B2(n15997), .A(n14581), .ZN(P1_U2893) );
  NAND2_X1 U17939 ( .A1(n14582), .A2(n16032), .ZN(n14583) );
  NAND2_X1 U17940 ( .A1(n20014), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14749) );
  OAI211_X1 U17941 ( .C1(n14723), .C2(n14584), .A(n14583), .B(n14749), .ZN(
        n14585) );
  AOI21_X1 U17942 ( .B1(n19962), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14587), .ZN(n14588) );
  OAI21_X1 U17943 ( .B1(n14589), .B2(n19972), .A(n14588), .ZN(n14590) );
  AOI21_X1 U17944 ( .B1(n14591), .B2(n14671), .A(n14590), .ZN(n14592) );
  OAI21_X1 U17945 ( .B1(n14593), .B2(n16035), .A(n14592), .ZN(P1_U2970) );
  NAND2_X1 U17946 ( .A1(n14844), .A2(n14595), .ZN(n14616) );
  NAND2_X1 U17947 ( .A1(n14594), .A2(n14616), .ZN(n14599) );
  OAI21_X1 U17948 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n14596), .A(
        n14599), .ZN(n14598) );
  MUX2_X1 U17949 ( .A(n14609), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n14844), .Z(n14597) );
  OAI211_X1 U17950 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14599), .A(
        n14598), .B(n14597), .ZN(n14601) );
  XNOR2_X1 U17951 ( .A(n14601), .B(n14600), .ZN(n14764) );
  NAND2_X1 U17952 ( .A1(n20014), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14759) );
  OAI21_X1 U17953 ( .B1(n14723), .B2(n14602), .A(n14759), .ZN(n14604) );
  OAI21_X1 U17954 ( .B1(n16035), .B2(n14764), .A(n14606), .ZN(P1_U2971) );
  MUX2_X1 U17955 ( .A(n14608), .B(n14607), .S(n14841), .Z(n14610) );
  XNOR2_X1 U17956 ( .A(n14610), .B(n14609), .ZN(n14774) );
  NAND2_X1 U17957 ( .A1(n20014), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14768) );
  NAND2_X1 U17958 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14611) );
  OAI211_X1 U17959 ( .C1(n14612), .C2(n19972), .A(n14768), .B(n14611), .ZN(
        n14613) );
  AOI21_X1 U17960 ( .B1(n14614), .B2(n14671), .A(n14613), .ZN(n14615) );
  OAI21_X1 U17961 ( .B1(n16035), .B2(n14774), .A(n14615), .ZN(P1_U2972) );
  OAI211_X1 U17962 ( .C1(n14841), .C2(n14594), .A(n14617), .B(n14616), .ZN(
        n14618) );
  XOR2_X1 U17963 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n14618), .Z(
        n14785) );
  NAND2_X1 U17964 ( .A1(n14619), .A2(n16032), .ZN(n14620) );
  NAND2_X1 U17965 ( .A1(n20014), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14779) );
  OAI211_X1 U17966 ( .C1(n14723), .C2(n14621), .A(n14620), .B(n14779), .ZN(
        n14622) );
  AOI21_X1 U17967 ( .B1(n14623), .B2(n14671), .A(n14622), .ZN(n14624) );
  OAI21_X1 U17968 ( .B1(n16035), .B2(n14785), .A(n14624), .ZN(P1_U2973) );
  NOR3_X1 U17969 ( .A1(n14594), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14627) );
  NAND2_X1 U17970 ( .A1(n14625), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14634) );
  NOR2_X1 U17971 ( .A1(n14634), .A2(n14801), .ZN(n14626) );
  MUX2_X1 U17972 ( .A(n14627), .B(n14626), .S(n14844), .Z(n14628) );
  XNOR2_X1 U17973 ( .A(n14628), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14794) );
  NOR2_X1 U17974 ( .A1(n16122), .A2(n20610), .ZN(n14787) );
  AOI21_X1 U17975 ( .B1(n19962), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14787), .ZN(n14629) );
  OAI21_X1 U17976 ( .B1(n14630), .B2(n19972), .A(n14629), .ZN(n14631) );
  AOI21_X1 U17977 ( .B1(n14632), .B2(n14671), .A(n14631), .ZN(n14633) );
  OAI21_X1 U17978 ( .B1(n16035), .B2(n14794), .A(n14633), .ZN(P1_U2974) );
  NOR2_X1 U17979 ( .A1(n14594), .A2(n14844), .ZN(n14635) );
  MUX2_X1 U17980 ( .A(n12874), .B(n14635), .S(n14634), .Z(n14636) );
  XNOR2_X1 U17981 ( .A(n14636), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14806) );
  NAND2_X1 U17982 ( .A1(n20014), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14800) );
  OAI21_X1 U17983 ( .B1(n14723), .B2(n14637), .A(n14800), .ZN(n14640) );
  NOR2_X1 U17984 ( .A1(n14638), .A2(n20022), .ZN(n14639) );
  AOI211_X1 U17985 ( .C1(n16032), .C2(n14641), .A(n14640), .B(n14639), .ZN(
        n14642) );
  OAI21_X1 U17986 ( .B1(n14806), .B2(n16035), .A(n14642), .ZN(P1_U2975) );
  XNOR2_X1 U17987 ( .A(n14844), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14643) );
  XNOR2_X1 U17988 ( .A(n14594), .B(n14643), .ZN(n14814) );
  INV_X1 U17989 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20608) );
  NOR2_X1 U17990 ( .A1(n16122), .A2(n20608), .ZN(n14807) );
  AOI21_X1 U17991 ( .B1(n19962), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n14807), .ZN(n14644) );
  OAI21_X1 U17992 ( .B1(n14645), .B2(n19972), .A(n14644), .ZN(n14646) );
  AOI21_X1 U17993 ( .B1(n14647), .B2(n14671), .A(n14646), .ZN(n14648) );
  OAI21_X1 U17994 ( .B1(n14814), .B2(n16035), .A(n14648), .ZN(P1_U2976) );
  INV_X1 U17995 ( .A(n14652), .ZN(n14650) );
  OR2_X1 U17996 ( .A1(n14650), .A2(n14649), .ZN(n14656) );
  NAND2_X1 U17997 ( .A1(n14652), .A2(n14651), .ZN(n14654) );
  NAND2_X1 U17998 ( .A1(n14654), .A2(n14653), .ZN(n14655) );
  NAND2_X1 U17999 ( .A1(n14656), .A2(n14655), .ZN(n14822) );
  INV_X1 U18000 ( .A(n15882), .ZN(n14658) );
  NOR2_X1 U18001 ( .A1(n16122), .A2(n15884), .ZN(n14815) );
  AOI21_X1 U18002 ( .B1(n19962), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n14815), .ZN(n14657) );
  OAI21_X1 U18003 ( .B1(n14658), .B2(n19972), .A(n14657), .ZN(n14659) );
  AOI21_X1 U18004 ( .B1(n15889), .B2(n14671), .A(n14659), .ZN(n14660) );
  OAI21_X1 U18005 ( .B1(n16035), .B2(n14822), .A(n14660), .ZN(P1_U2977) );
  NOR2_X1 U18006 ( .A1(n14674), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14664) );
  NOR2_X1 U18007 ( .A1(n14661), .A2(n14662), .ZN(n14663) );
  MUX2_X1 U18008 ( .A(n14664), .B(n14663), .S(n12874), .Z(n14665) );
  XNOR2_X1 U18009 ( .A(n14665), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14832) );
  INV_X1 U18010 ( .A(n14469), .ZN(n14666) );
  AOI21_X1 U18011 ( .B1(n14668), .B2(n14667), .A(n14666), .ZN(n15998) );
  NAND2_X1 U18012 ( .A1(n20014), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14827) );
  NAND2_X1 U18013 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14669) );
  OAI211_X1 U18014 ( .C1(n15901), .C2(n19972), .A(n14827), .B(n14669), .ZN(
        n14670) );
  AOI21_X1 U18015 ( .B1(n15998), .B2(n14671), .A(n14670), .ZN(n14672) );
  OAI21_X1 U18016 ( .B1(n16035), .B2(n14832), .A(n14672), .ZN(P1_U2978) );
  NAND2_X1 U18017 ( .A1(n9601), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14673) );
  MUX2_X1 U18018 ( .A(n14674), .B(n14673), .S(n14844), .Z(n14675) );
  XNOR2_X1 U18019 ( .A(n14675), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15869) );
  NAND2_X1 U18020 ( .A1(n15869), .A2(n19968), .ZN(n14679) );
  INV_X1 U18021 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n14676) );
  OAI22_X1 U18022 ( .A1(n14723), .A2(n15903), .B1(n16122), .B2(n14676), .ZN(
        n14677) );
  AOI21_X1 U18023 ( .B1(n15912), .B2(n16032), .A(n14677), .ZN(n14678) );
  OAI211_X1 U18024 ( .C1(n20022), .C2(n15909), .A(n14679), .B(n14678), .ZN(
        P1_U2979) );
  NOR2_X1 U18025 ( .A1(n14844), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14680) );
  MUX2_X1 U18026 ( .A(n12874), .B(n14680), .S(n14661), .Z(n14681) );
  XNOR2_X1 U18027 ( .A(n14681), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14840) );
  AND2_X1 U18028 ( .A1(n14683), .A2(n14682), .ZN(n14684) );
  NOR2_X1 U18029 ( .A1(n16122), .A2(n20602), .ZN(n14836) );
  AOI21_X1 U18030 ( .B1(n19962), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n14836), .ZN(n14685) );
  OAI21_X1 U18031 ( .B1(n15915), .B2(n19972), .A(n14685), .ZN(n14686) );
  AOI21_X1 U18032 ( .B1(n10076), .B2(n14671), .A(n14686), .ZN(n14687) );
  OAI21_X1 U18033 ( .B1(n14840), .B2(n16035), .A(n14687), .ZN(P1_U2980) );
  OAI21_X1 U18034 ( .B1(n14689), .B2(n14688), .A(n14661), .ZN(n16061) );
  OAI22_X1 U18035 ( .A1(n14723), .A2(n15926), .B1(n16122), .B2(n20599), .ZN(
        n14691) );
  NOR2_X1 U18036 ( .A1(n15930), .A2(n20022), .ZN(n14690) );
  AOI211_X1 U18037 ( .C1(n16032), .C2(n15929), .A(n14691), .B(n14690), .ZN(
        n14692) );
  OAI21_X1 U18038 ( .B1(n16035), .B2(n16061), .A(n14692), .ZN(P1_U2981) );
  INV_X1 U18039 ( .A(n14863), .ZN(n14695) );
  AOI21_X1 U18040 ( .B1(n14694), .B2(n14696), .A(n14695), .ZN(n14698) );
  XNOR2_X1 U18041 ( .A(n14698), .B(n14697), .ZN(n16069) );
  INV_X1 U18042 ( .A(n15950), .ZN(n14700) );
  AOI22_X1 U18043 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20014), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n14699) );
  OAI21_X1 U18044 ( .B1(n14700), .B2(n19972), .A(n14699), .ZN(n14701) );
  AOI21_X1 U18045 ( .B1(n14702), .B2(n14671), .A(n14701), .ZN(n14703) );
  OAI21_X1 U18046 ( .B1(n16035), .B2(n16069), .A(n14703), .ZN(P1_U2983) );
  NOR2_X1 U18047 ( .A1(n14844), .A2(n16098), .ZN(n14719) );
  NOR2_X1 U18048 ( .A1(n14844), .A2(n14705), .ZN(n14715) );
  NOR3_X1 U18049 ( .A1(n14717), .A2(n14719), .A3(n14715), .ZN(n14843) );
  INV_X1 U18050 ( .A(n14706), .ZN(n14708) );
  OAI21_X1 U18051 ( .B1(n14843), .B2(n14708), .A(n14707), .ZN(n14710) );
  XNOR2_X1 U18052 ( .A(n14844), .B(n16081), .ZN(n14709) );
  XNOR2_X1 U18053 ( .A(n14710), .B(n14709), .ZN(n16079) );
  INV_X1 U18054 ( .A(n16079), .ZN(n14714) );
  AOI22_X1 U18055 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20014), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n14711) );
  OAI21_X1 U18056 ( .B1(n19972), .B2(n15962), .A(n14711), .ZN(n14712) );
  AOI21_X1 U18057 ( .B1(n15964), .B2(n14671), .A(n14712), .ZN(n14713) );
  OAI21_X1 U18058 ( .B1(n14714), .B2(n16035), .A(n14713), .ZN(P1_U2985) );
  AOI21_X1 U18059 ( .B1(n14717), .B2(n14716), .A(n14715), .ZN(n16028) );
  INV_X1 U18060 ( .A(n14720), .ZN(n14718) );
  NOR2_X1 U18061 ( .A1(n14719), .A2(n14718), .ZN(n16027) );
  NAND2_X1 U18062 ( .A1(n16028), .A2(n16027), .ZN(n16026) );
  NAND2_X1 U18063 ( .A1(n16026), .A2(n14720), .ZN(n14721) );
  XOR2_X1 U18064 ( .A(n14722), .B(n14721), .Z(n16088) );
  NAND2_X1 U18065 ( .A1(n16088), .A2(n19968), .ZN(n14727) );
  OAI22_X1 U18066 ( .A1(n14723), .A2(n14455), .B1(n16122), .B2(n20592), .ZN(
        n14724) );
  AOI21_X1 U18067 ( .B1(n16032), .B2(n14725), .A(n14724), .ZN(n14726) );
  OAI211_X1 U18068 ( .C1(n20022), .C2(n14728), .A(n14727), .B(n14726), .ZN(
        P1_U2986) );
  MUX2_X1 U18069 ( .A(n14729), .B(n14704), .S(n14844), .Z(n14730) );
  XOR2_X1 U18070 ( .A(n16114), .B(n14730), .Z(n16118) );
  AOI22_X1 U18071 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20014), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14734) );
  INV_X1 U18072 ( .A(n14731), .ZN(n14732) );
  NAND2_X1 U18073 ( .A1(n16032), .A2(n14732), .ZN(n14733) );
  OAI211_X1 U18074 ( .C1(n14735), .C2(n20022), .A(n14734), .B(n14733), .ZN(
        n14736) );
  AOI21_X1 U18075 ( .B1(n16118), .B2(n19968), .A(n14736), .ZN(n14737) );
  INV_X1 U18076 ( .A(n14737), .ZN(P1_U2989) );
  NOR2_X1 U18077 ( .A1(n14738), .A2(n20017), .ZN(n14742) );
  INV_X1 U18078 ( .A(n14766), .ZN(n14747) );
  INV_X1 U18079 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14881) );
  AOI211_X1 U18080 ( .C1(n14748), .C2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n14747), .B(n14881), .ZN(n14741) );
  INV_X1 U18081 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14746) );
  NOR4_X1 U18082 ( .A1(n14751), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14750), .A4(n14746), .ZN(n14739) );
  OAI21_X1 U18083 ( .B1(n14744), .B2(n16126), .A(n14743), .ZN(P1_U3000) );
  NOR3_X1 U18084 ( .A1(n14748), .A2(n14747), .A3(n14746), .ZN(n14754) );
  INV_X1 U18085 ( .A(n14749), .ZN(n14753) );
  NOR3_X1 U18086 ( .A1(n14751), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14750), .ZN(n14752) );
  NAND3_X1 U18087 ( .A1(n14765), .A2(n14757), .A3(n14756), .ZN(n14760) );
  NAND3_X1 U18088 ( .A1(n14767), .A2(n14766), .A3(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14758) );
  NAND3_X1 U18089 ( .A1(n14760), .A2(n14759), .A3(n14758), .ZN(n14761) );
  AOI21_X1 U18090 ( .B1(n14762), .B2(n19981), .A(n14761), .ZN(n14763) );
  OAI21_X1 U18091 ( .B1(n14764), .B2(n16126), .A(n14763), .ZN(P1_U3003) );
  INV_X1 U18092 ( .A(n14765), .ZN(n14770) );
  NAND3_X1 U18093 ( .A1(n14767), .A2(n14766), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14769) );
  OAI211_X1 U18094 ( .C1(n14770), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14769), .B(n14768), .ZN(n14771) );
  AOI21_X1 U18095 ( .B1(n14772), .B2(n19981), .A(n14771), .ZN(n14773) );
  OAI21_X1 U18096 ( .B1(n14774), .B2(n16126), .A(n14773), .ZN(P1_U3004) );
  NAND3_X1 U18097 ( .A1(n14775), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14776) );
  OR2_X1 U18098 ( .A1(n14810), .A2(n14776), .ZN(n14789) );
  INV_X1 U18099 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14777) );
  AOI21_X1 U18100 ( .B1(n14789), .B2(n14786), .A(n14777), .ZN(n14782) );
  INV_X1 U18101 ( .A(n14810), .ZN(n14798) );
  NAND3_X1 U18102 ( .A1(n14798), .A2(n14778), .A3(n14777), .ZN(n14780) );
  NAND2_X1 U18103 ( .A1(n14780), .A2(n14779), .ZN(n14781) );
  AOI211_X1 U18104 ( .C1(n14783), .C2(n19981), .A(n14782), .B(n14781), .ZN(
        n14784) );
  OAI21_X1 U18105 ( .B1(n14785), .B2(n16126), .A(n14784), .ZN(P1_U3005) );
  INV_X1 U18106 ( .A(n14786), .ZN(n14788) );
  AOI21_X1 U18107 ( .B1(n14788), .B2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n14787), .ZN(n14790) );
  OAI211_X1 U18108 ( .C1(n14791), .C2(n20017), .A(n14790), .B(n14789), .ZN(
        n14792) );
  INV_X1 U18109 ( .A(n14792), .ZN(n14793) );
  OAI21_X1 U18110 ( .B1(n14794), .B2(n16126), .A(n14793), .ZN(P1_U3006) );
  INV_X1 U18111 ( .A(n14795), .ZN(n14796) );
  AOI21_X1 U18112 ( .B1(n19988), .B2(n14797), .A(n14796), .ZN(n14802) );
  NAND3_X1 U18113 ( .A1(n14798), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n14801), .ZN(n14799) );
  OAI211_X1 U18114 ( .C1(n14802), .C2(n14801), .A(n14800), .B(n14799), .ZN(
        n14803) );
  AOI21_X1 U18115 ( .B1(n14804), .B2(n19981), .A(n14803), .ZN(n14805) );
  OAI21_X1 U18116 ( .B1(n14806), .B2(n16126), .A(n14805), .ZN(P1_U3007) );
  AOI21_X1 U18117 ( .B1(n14808), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n14807), .ZN(n14809) );
  OAI21_X1 U18118 ( .B1(n14810), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n14809), .ZN(n14811) );
  AOI21_X1 U18119 ( .B1(n14812), .B2(n19981), .A(n14811), .ZN(n14813) );
  OAI21_X1 U18120 ( .B1(n14814), .B2(n16126), .A(n14813), .ZN(P1_U3008) );
  INV_X1 U18121 ( .A(n15893), .ZN(n14820) );
  XNOR2_X1 U18122 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14818) );
  INV_X1 U18123 ( .A(n14828), .ZN(n14816) );
  AOI21_X1 U18124 ( .B1(n14816), .B2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n14815), .ZN(n14817) );
  OAI21_X1 U18125 ( .B1(n14829), .B2(n14818), .A(n14817), .ZN(n14819) );
  AOI21_X1 U18126 ( .B1(n14820), .B2(n19981), .A(n14819), .ZN(n14821) );
  OAI21_X1 U18127 ( .B1(n14822), .B2(n16126), .A(n14821), .ZN(P1_U3009) );
  OAI21_X1 U18128 ( .B1(n14825), .B2(n14824), .A(n14823), .ZN(n14826) );
  INV_X1 U18129 ( .A(n14826), .ZN(n15987) );
  OAI221_X1 U18130 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n14829), 
        .C1(n12896), .C2(n14828), .A(n14827), .ZN(n14830) );
  AOI21_X1 U18131 ( .B1(n15987), .B2(n19981), .A(n14830), .ZN(n14831) );
  OAI21_X1 U18132 ( .B1(n14832), .B2(n16126), .A(n14831), .ZN(P1_U3010) );
  AOI21_X1 U18133 ( .B1(n14835), .B2(n14834), .A(n14833), .ZN(n15990) );
  AOI21_X1 U18134 ( .B1(n15862), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n14836), .ZN(n14837) );
  OAI21_X1 U18135 ( .B1(n15861), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n14837), .ZN(n14838) );
  AOI21_X1 U18136 ( .B1(n15990), .B2(n19981), .A(n14838), .ZN(n14839) );
  OAI21_X1 U18137 ( .B1(n14840), .B2(n16126), .A(n14839), .ZN(P1_U3012) );
  NAND2_X1 U18138 ( .A1(n14841), .A2(n16076), .ZN(n14849) );
  NOR2_X1 U18139 ( .A1(n14843), .A2(n14842), .ZN(n14847) );
  OAI21_X1 U18140 ( .B1(n14845), .B2(n14844), .A(n14864), .ZN(n14846) );
  OAI21_X1 U18141 ( .B1(n14847), .B2(n14846), .A(n9703), .ZN(n14848) );
  MUX2_X1 U18142 ( .A(n14841), .B(n14849), .S(n14848), .Z(n14850) );
  XNOR2_X1 U18143 ( .A(n14850), .B(n12890), .ZN(n16020) );
  NOR2_X1 U18144 ( .A1(n16091), .A2(n14851), .ZN(n16068) );
  INV_X1 U18145 ( .A(n14852), .ZN(n16065) );
  INV_X1 U18146 ( .A(n20008), .ZN(n16134) );
  NOR2_X1 U18147 ( .A1(n14855), .A2(n14853), .ZN(n16082) );
  OAI21_X1 U18148 ( .B1(n14855), .B2(n14854), .A(n16093), .ZN(n14856) );
  OAI211_X1 U18149 ( .C1(n16082), .C2(n16095), .A(n19989), .B(n14856), .ZN(
        n16087) );
  AOI21_X1 U18150 ( .B1(n16081), .B2(n16134), .A(n16087), .ZN(n16077) );
  OAI21_X1 U18151 ( .B1(n20008), .B2(n16065), .A(n16077), .ZN(n16063) );
  OAI221_X1 U18152 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n16070), 
        .C1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n16068), .A(n16063), .ZN(
        n14862) );
  INV_X1 U18153 ( .A(n14857), .ZN(n14858) );
  AOI21_X1 U18154 ( .B1(n14860), .B2(n14859), .A(n14858), .ZN(n15993) );
  AOI22_X1 U18155 ( .A1(n15993), .A2(n19981), .B1(n20014), .B2(
        P1_REIP_REG_17__SCAN_IN), .ZN(n14861) );
  OAI211_X1 U18156 ( .C1(n16020), .C2(n16126), .A(n14862), .B(n14861), .ZN(
        P1_U3014) );
  NAND2_X1 U18157 ( .A1(n14864), .A2(n14863), .ZN(n14867) );
  NAND2_X1 U18158 ( .A1(n14694), .A2(n14865), .ZN(n14866) );
  XOR2_X1 U18159 ( .A(n14867), .B(n14866), .Z(n16025) );
  INV_X1 U18160 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20594) );
  OAI22_X1 U18161 ( .A1(n16122), .A2(n20594), .B1(n16077), .B2(n14869), .ZN(
        n14868) );
  AOI21_X1 U18162 ( .B1(n15952), .B2(n19981), .A(n14868), .ZN(n14871) );
  NAND2_X1 U18163 ( .A1(n16068), .A2(n14869), .ZN(n14870) );
  OAI211_X1 U18164 ( .C1(n16025), .C2(n16126), .A(n14871), .B(n14870), .ZN(
        P1_U3016) );
  NOR2_X1 U18165 ( .A1(n13601), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14872) );
  OAI22_X1 U18166 ( .A1(n14873), .A2(n14872), .B1(n13646), .B2(n20644), .ZN(
        n14874) );
  MUX2_X1 U18167 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14874), .S(
        n20653), .Z(P1_U3477) );
  NOR2_X1 U18168 ( .A1(n13590), .A2(n13564), .ZN(n14876) );
  AOI22_X1 U18169 ( .A1(n14877), .A2(n11225), .B1(n14876), .B2(n14875), .ZN(
        n14878) );
  OAI21_X1 U18170 ( .B1(n13646), .B2(n14879), .A(n14878), .ZN(n15815) );
  INV_X1 U18171 ( .A(n15815), .ZN(n14885) );
  INV_X1 U18172 ( .A(n14880), .ZN(n20635) );
  OAI22_X1 U18173 ( .A1(n14881), .A2(n20011), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14888) );
  NOR2_X1 U18174 ( .A1(n20555), .A2(n14882), .ZN(n14890) );
  NOR3_X1 U18175 ( .A1(n13590), .A2(n13564), .A3(n20633), .ZN(n14883) );
  AOI21_X1 U18176 ( .B1(n14888), .B2(n14890), .A(n14883), .ZN(n14884) );
  OAI21_X1 U18177 ( .B1(n14885), .B2(n20635), .A(n14884), .ZN(n14886) );
  MUX2_X1 U18178 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14886), .S(
        n16157), .Z(P1_U3473) );
  INV_X1 U18179 ( .A(n14887), .ZN(n14891) );
  INV_X1 U18180 ( .A(n14888), .ZN(n14889) );
  AOI22_X1 U18181 ( .A1(n14891), .A2(n15846), .B1(n14890), .B2(n14889), .ZN(
        n14892) );
  OAI21_X1 U18182 ( .B1(n14893), .B2(n20635), .A(n14892), .ZN(n14894) );
  MUX2_X1 U18183 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14894), .S(
        n16157), .Z(P1_U3472) );
  OAI21_X1 U18184 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n14895), .A(
        n14913), .ZN(n18863) );
  AND2_X1 U18185 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n14906), .ZN(
        n14904) );
  OAI21_X1 U18186 ( .B1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n14904), .A(
        n14897), .ZN(n15382) );
  NOR2_X1 U18187 ( .A1(n15426), .A2(n14898), .ZN(n18910) );
  OAI21_X1 U18188 ( .B1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n13924), .A(
        n14900), .ZN(n18912) );
  NAND2_X1 U18189 ( .A1(n18910), .A2(n18912), .ZN(n18892) );
  AOI21_X1 U18190 ( .B1(n15409), .B2(n14900), .A(n14901), .ZN(n18895) );
  OR2_X1 U18191 ( .A1(n14901), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14903) );
  INV_X1 U18192 ( .A(n14906), .ZN(n14902) );
  NAND2_X1 U18193 ( .A1(n14903), .A2(n14902), .ZN(n15400) );
  INV_X1 U18194 ( .A(n14904), .ZN(n14905) );
  OAI21_X1 U18195 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n14906), .A(
        n14905), .ZN(n18887) );
  NAND2_X1 U18196 ( .A1(n18888), .A2(n18887), .ZN(n18886) );
  NAND2_X1 U18197 ( .A1(n15382), .A2(n15017), .ZN(n15016) );
  NAND2_X1 U18198 ( .A1(n15016), .A2(n18893), .ZN(n18875) );
  OAI21_X1 U18199 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n14907), .A(
        n14908), .ZN(n18876) );
  NAND2_X1 U18200 ( .A1(n18875), .A2(n18876), .ZN(n18874) );
  NAND2_X1 U18201 ( .A1(n18874), .A2(n18893), .ZN(n15003) );
  INV_X1 U18202 ( .A(n14908), .ZN(n14910) );
  INV_X1 U18203 ( .A(n14895), .ZN(n14909) );
  OAI21_X1 U18204 ( .B1(n14910), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n14909), .ZN(n15363) );
  NAND2_X1 U18205 ( .A1(n15003), .A2(n15363), .ZN(n15002) );
  NAND2_X1 U18206 ( .A1(n18863), .A2(n18862), .ZN(n18861) );
  INV_X1 U18207 ( .A(n14912), .ZN(n14915) );
  NAND2_X1 U18208 ( .A1(n11216), .A2(n14913), .ZN(n14914) );
  NAND2_X1 U18209 ( .A1(n14915), .A2(n14914), .ZN(n15340) );
  NAND2_X1 U18210 ( .A1(n14991), .A2(n15340), .ZN(n14990) );
  NAND2_X1 U18211 ( .A1(n14990), .A2(n18893), .ZN(n15805) );
  OAI21_X1 U18212 ( .B1(n14912), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n14916), .ZN(n15806) );
  NAND2_X1 U18213 ( .A1(n15805), .A2(n15806), .ZN(n15804) );
  AOI21_X1 U18214 ( .B1(n15303), .B2(n14916), .A(n14919), .ZN(n15306) );
  INV_X1 U18215 ( .A(n15306), .ZN(n16223) );
  NAND2_X1 U18216 ( .A1(n16222), .A2(n16223), .ZN(n16221) );
  NAND2_X1 U18217 ( .A1(n16221), .A2(n18893), .ZN(n14977) );
  OR2_X1 U18218 ( .A1(n14919), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14920) );
  NAND2_X1 U18219 ( .A1(n14918), .A2(n14920), .ZN(n15295) );
  NAND2_X1 U18220 ( .A1(n14977), .A2(n15295), .ZN(n14976) );
  NAND2_X1 U18221 ( .A1(n14976), .A2(n18893), .ZN(n14964) );
  NAND2_X1 U18222 ( .A1(n14918), .A2(n15282), .ZN(n14921) );
  NAND2_X1 U18223 ( .A1(n14923), .A2(n14921), .ZN(n15279) );
  NAND2_X1 U18224 ( .A1(n14964), .A2(n15279), .ZN(n14963) );
  NAND2_X1 U18225 ( .A1(n14963), .A2(n18893), .ZN(n16211) );
  NAND2_X1 U18226 ( .A1(n14923), .A2(n14922), .ZN(n14924) );
  NAND2_X1 U18227 ( .A1(n14925), .A2(n14924), .ZN(n16212) );
  NAND2_X1 U18228 ( .A1(n16211), .A2(n16212), .ZN(n16210) );
  NAND2_X1 U18229 ( .A1(n16210), .A2(n18893), .ZN(n14945) );
  INV_X1 U18230 ( .A(n14928), .ZN(n14927) );
  NAND2_X1 U18231 ( .A1(n14925), .A2(n14952), .ZN(n14926) );
  NAND2_X1 U18232 ( .A1(n14927), .A2(n14926), .ZN(n15261) );
  NAND2_X1 U18233 ( .A1(n14945), .A2(n15261), .ZN(n14944) );
  NAND2_X1 U18234 ( .A1(n14944), .A2(n18893), .ZN(n16198) );
  OR2_X1 U18235 ( .A1(n14928), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14929) );
  NAND2_X1 U18236 ( .A1(n11217), .A2(n14929), .ZN(n16199) );
  NAND2_X1 U18237 ( .A1(n16198), .A2(n16199), .ZN(n16197) );
  NAND2_X1 U18238 ( .A1(n16197), .A2(n18893), .ZN(n14931) );
  NAND2_X1 U18239 ( .A1(n14931), .A2(n14930), .ZN(n16176) );
  OAI211_X1 U18240 ( .C1(n14931), .C2(n14930), .A(n18949), .B(n16176), .ZN(
        n14942) );
  NOR2_X1 U18241 ( .A1(n15136), .A2(n14932), .ZN(n14933) );
  NOR2_X1 U18242 ( .A1(n15499), .A2(n18947), .ZN(n14940) );
  NOR2_X1 U18243 ( .A1(n14935), .A2(n18936), .ZN(n14939) );
  OAI22_X1 U18244 ( .A1(n14936), .A2(n18935), .B1(n19693), .B2(n18927), .ZN(
        n14938) );
  NOR2_X1 U18245 ( .A1(n18954), .A2(n11205), .ZN(n14937) );
  NOR4_X1 U18246 ( .A1(n14940), .A2(n14939), .A3(n14938), .A4(n14937), .ZN(
        n14941) );
  OAI211_X1 U18247 ( .C1(n15503), .C2(n18946), .A(n14942), .B(n14941), .ZN(
        P2_U2826) );
  XNOR2_X1 U18248 ( .A(n15074), .B(n14943), .ZN(n15529) );
  OAI211_X1 U18249 ( .C1(n14945), .C2(n15261), .A(n18949), .B(n14944), .ZN(
        n14958) );
  OR2_X1 U18250 ( .A1(n14947), .A2(n14946), .ZN(n14948) );
  NAND2_X1 U18251 ( .A1(n14949), .A2(n14948), .ZN(n15241) );
  AND2_X1 U18252 ( .A1(n15148), .A2(n14950), .ZN(n14951) );
  NOR2_X1 U18253 ( .A1(n15134), .A2(n14951), .ZN(n15526) );
  INV_X1 U18254 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19690) );
  OAI22_X1 U18255 ( .A1(n14952), .A2(n18935), .B1(n19690), .B2(n18927), .ZN(
        n14954) );
  NOR2_X1 U18256 ( .A1(n18954), .A2(n11196), .ZN(n14953) );
  AOI211_X1 U18257 ( .C1(n15526), .C2(n18901), .A(n14954), .B(n14953), .ZN(
        n14955) );
  OAI21_X1 U18258 ( .B1(n15241), .B2(n18936), .A(n14955), .ZN(n14956) );
  INV_X1 U18259 ( .A(n14956), .ZN(n14957) );
  OAI211_X1 U18260 ( .C1(n15529), .C2(n18946), .A(n14958), .B(n14957), .ZN(
        P2_U2828) );
  NOR2_X1 U18261 ( .A1(n14974), .A2(n14959), .ZN(n14960) );
  OR2_X1 U18262 ( .A1(n15076), .A2(n14960), .ZN(n15278) );
  INV_X1 U18263 ( .A(n14961), .ZN(n14971) );
  XNOR2_X1 U18264 ( .A(n14979), .B(n14962), .ZN(n15550) );
  OAI211_X1 U18265 ( .C1(n15279), .C2(n14964), .A(n18949), .B(n14963), .ZN(
        n14967) );
  OAI22_X1 U18266 ( .A1(n15282), .A2(n18935), .B1(n19686), .B2(n18927), .ZN(
        n14965) );
  INV_X1 U18267 ( .A(n14965), .ZN(n14966) );
  NAND2_X1 U18268 ( .A1(n14967), .A2(n14966), .ZN(n14968) );
  AOI21_X1 U18269 ( .B1(n18922), .B2(P2_EBX_REG_25__SCAN_IN), .A(n14968), .ZN(
        n14969) );
  OAI21_X1 U18270 ( .B1(n15550), .B2(n18947), .A(n14969), .ZN(n14970) );
  AOI21_X1 U18271 ( .B1(n14971), .B2(n18923), .A(n14970), .ZN(n14972) );
  OAI21_X1 U18272 ( .B1(n15278), .B2(n18946), .A(n14972), .ZN(P2_U2830) );
  AND2_X1 U18273 ( .A1(n9668), .A2(n14973), .ZN(n14975) );
  OR2_X1 U18274 ( .A1(n14975), .A2(n14974), .ZN(n15564) );
  OAI211_X1 U18275 ( .C1(n14977), .C2(n15295), .A(n18949), .B(n14976), .ZN(
        n14987) );
  OAI21_X1 U18276 ( .B1(n14978), .B2(n14980), .A(n14979), .ZN(n14981) );
  INV_X1 U18277 ( .A(n14981), .ZN(n16229) );
  AOI22_X1 U18278 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18931), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n18940), .ZN(n14982) );
  OAI21_X1 U18279 ( .B1(n18954), .B2(n15090), .A(n14982), .ZN(n14985) );
  NOR2_X1 U18280 ( .A1(n14983), .A2(n18936), .ZN(n14984) );
  AOI211_X1 U18281 ( .C1(n18901), .C2(n16229), .A(n14985), .B(n14984), .ZN(
        n14986) );
  OAI211_X1 U18282 ( .C1(n18946), .C2(n15564), .A(n14987), .B(n14986), .ZN(
        P2_U2831) );
  AND2_X1 U18283 ( .A1(n15117), .A2(n14988), .ZN(n14989) );
  NOR2_X1 U18284 ( .A1(n9696), .A2(n14989), .ZN(n15595) );
  INV_X1 U18285 ( .A(n15595), .ZN(n15111) );
  OAI211_X1 U18286 ( .C1(n14991), .C2(n15340), .A(n18949), .B(n14990), .ZN(
        n15001) );
  INV_X1 U18287 ( .A(n14992), .ZN(n14999) );
  OAI22_X1 U18288 ( .A1(n18954), .A2(n15112), .B1(n20763), .B2(n18927), .ZN(
        n14998) );
  NAND2_X1 U18289 ( .A1(n14993), .A2(n14994), .ZN(n14995) );
  AND2_X1 U18290 ( .A1(n15174), .A2(n14995), .ZN(n15597) );
  INV_X1 U18291 ( .A(n15597), .ZN(n14996) );
  OAI22_X1 U18292 ( .A1(n14996), .A2(n18947), .B1(n18935), .B2(n11216), .ZN(
        n14997) );
  AOI211_X1 U18293 ( .C1(n14999), .C2(n18923), .A(n14998), .B(n14997), .ZN(
        n15000) );
  OAI211_X1 U18294 ( .C1(n18946), .C2(n15111), .A(n15001), .B(n15000), .ZN(
        P2_U2834) );
  OAI211_X1 U18295 ( .C1(n15003), .C2(n15363), .A(n18949), .B(n15002), .ZN(
        n15014) );
  INV_X1 U18296 ( .A(n15004), .ZN(n15005) );
  XNOR2_X1 U18297 ( .A(n15006), .B(n15005), .ZN(n16236) );
  INV_X1 U18298 ( .A(n16236), .ZN(n15010) );
  AOI21_X1 U18299 ( .B1(P2_REIP_REG_19__SCAN_IN), .B2(n18940), .A(n18939), 
        .ZN(n15007) );
  OAI21_X1 U18300 ( .B1(n15364), .B2(n18935), .A(n15007), .ZN(n15008) );
  AOI21_X1 U18301 ( .B1(n18922), .B2(P2_EBX_REG_19__SCAN_IN), .A(n15008), .ZN(
        n15009) );
  OAI21_X1 U18302 ( .B1(n15010), .B2(n18947), .A(n15009), .ZN(n15011) );
  AOI21_X1 U18303 ( .B1(n15012), .B2(n18923), .A(n15011), .ZN(n15013) );
  OAI211_X1 U18304 ( .C1(n18946), .C2(n15015), .A(n15014), .B(n15013), .ZN(
        P2_U2836) );
  OAI211_X1 U18305 ( .C1(n15382), .C2(n15017), .A(n18949), .B(n15016), .ZN(
        n15027) );
  INV_X1 U18306 ( .A(n15018), .ZN(n15025) );
  NAND2_X1 U18307 ( .A1(n15020), .A2(n15019), .ZN(n15021) );
  NAND2_X1 U18308 ( .A1(n15197), .A2(n15021), .ZN(n15650) );
  NOR2_X1 U18309 ( .A1(n15650), .A2(n18947), .ZN(n15024) );
  AOI22_X1 U18310 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n18931), .B1(
        P2_EBX_REG_17__SCAN_IN), .B2(n18922), .ZN(n15022) );
  OAI211_X1 U18311 ( .C1(n18927), .C2(n19671), .A(n15022), .B(n16290), .ZN(
        n15023) );
  AOI211_X1 U18312 ( .C1(n15025), .C2(n18923), .A(n15024), .B(n15023), .ZN(
        n15026) );
  OAI211_X1 U18313 ( .C1(n15028), .C2(n18946), .A(n15027), .B(n15026), .ZN(
        P2_U2838) );
  OAI211_X1 U18314 ( .C1(n15030), .C2(n15400), .A(n18949), .B(n15029), .ZN(
        n15041) );
  INV_X1 U18315 ( .A(n15031), .ZN(n15039) );
  AND2_X1 U18316 ( .A1(n15032), .A2(n15033), .ZN(n15035) );
  OR2_X1 U18317 ( .A1(n15035), .A2(n15034), .ZN(n18961) );
  NOR2_X1 U18318 ( .A1(n18961), .A2(n18947), .ZN(n15038) );
  AOI22_X1 U18319 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18931), .B1(
        P2_EBX_REG_15__SCAN_IN), .B2(n18922), .ZN(n15036) );
  OAI211_X1 U18320 ( .C1(n18927), .C2(n19667), .A(n15036), .B(n18925), .ZN(
        n15037) );
  AOI211_X1 U18321 ( .C1(n15039), .C2(n18923), .A(n15038), .B(n15037), .ZN(
        n15040) );
  OAI211_X1 U18322 ( .C1(n18946), .C2(n15042), .A(n15041), .B(n15040), .ZN(
        P2_U2840) );
  NAND2_X1 U18323 ( .A1(n15044), .A2(n15043), .ZN(n15050) );
  AOI22_X1 U18324 ( .A1(n11148), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n15048) );
  NAND2_X1 U18325 ( .A1(n15046), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n15047) );
  OAI211_X1 U18326 ( .C1(n11121), .C2(n15470), .A(n15048), .B(n15047), .ZN(
        n15049) );
  NAND2_X1 U18327 ( .A1(n16175), .A2(n15110), .ZN(n15051) );
  OAI21_X1 U18328 ( .B1(n15110), .B2(n15052), .A(n15051), .ZN(P2_U2856) );
  XNOR2_X1 U18329 ( .A(n15053), .B(n15054), .ZN(n15129) );
  NOR2_X1 U18330 ( .A1(n15503), .A2(n13198), .ZN(n15055) );
  AOI21_X1 U18331 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n13198), .A(n15055), .ZN(
        n15056) );
  OAI21_X1 U18332 ( .B1(n15129), .B2(n15114), .A(n15056), .ZN(P2_U2858) );
  INV_X1 U18333 ( .A(n15057), .ZN(n15058) );
  NOR2_X1 U18334 ( .A1(n15059), .A2(n15058), .ZN(n15061) );
  XNOR2_X1 U18335 ( .A(n15061), .B(n15060), .ZN(n15140) );
  NAND2_X1 U18336 ( .A1(n15063), .A2(n15062), .ZN(n15064) );
  NAND2_X1 U18337 ( .A1(n15065), .A2(n15064), .ZN(n16195) );
  NOR2_X1 U18338 ( .A1(n16195), .A2(n13198), .ZN(n15066) );
  AOI21_X1 U18339 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n13198), .A(n15066), .ZN(
        n15067) );
  OAI21_X1 U18340 ( .B1(n15140), .B2(n15114), .A(n15067), .ZN(P2_U2859) );
  INV_X1 U18341 ( .A(n15071), .ZN(n15145) );
  NOR2_X1 U18342 ( .A1(n15529), .A2(n13198), .ZN(n15072) );
  AOI21_X1 U18343 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n13198), .A(n15072), .ZN(
        n15073) );
  OAI21_X1 U18344 ( .B1(n15145), .B2(n15114), .A(n15073), .ZN(P2_U2860) );
  OAI21_X1 U18345 ( .B1(n15076), .B2(n15075), .A(n15074), .ZN(n15538) );
  AOI21_X1 U18346 ( .B1(n15077), .B2(n15079), .A(n15078), .ZN(n15153) );
  NAND2_X1 U18347 ( .A1(n15153), .A2(n15119), .ZN(n15081) );
  NAND2_X1 U18348 ( .A1(n15122), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15080) );
  OAI211_X1 U18349 ( .C1(n15122), .C2(n15538), .A(n15081), .B(n15080), .ZN(
        P2_U2861) );
  XNOR2_X1 U18350 ( .A(n15082), .B(n15083), .ZN(n15161) );
  MUX2_X1 U18351 ( .A(n15278), .B(n9879), .S(n15122), .Z(n15084) );
  OAI21_X1 U18352 ( .B1(n15161), .B2(n15114), .A(n15084), .ZN(P2_U2862) );
  NAND2_X1 U18353 ( .A1(n12687), .A2(n15086), .ZN(n15087) );
  XNOR2_X1 U18354 ( .A(n15088), .B(n15087), .ZN(n15089) );
  XNOR2_X1 U18355 ( .A(n15085), .B(n15089), .ZN(n16228) );
  MUX2_X1 U18356 ( .A(n15564), .B(n15090), .S(n15122), .Z(n15091) );
  OAI21_X1 U18357 ( .B1(n16228), .B2(n15114), .A(n15091), .ZN(P2_U2863) );
  OAI21_X1 U18358 ( .B1(n15092), .B2(n15095), .A(n15094), .ZN(n15170) );
  NAND2_X1 U18359 ( .A1(n15096), .A2(n15097), .ZN(n15098) );
  NAND2_X1 U18360 ( .A1(n9668), .A2(n15098), .ZN(n15572) );
  NOR2_X1 U18361 ( .A1(n15572), .A2(n13198), .ZN(n15099) );
  AOI21_X1 U18362 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n15122), .A(n15099), .ZN(
        n15100) );
  OAI21_X1 U18363 ( .B1(n15170), .B2(n15114), .A(n15100), .ZN(P2_U2864) );
  OR2_X1 U18364 ( .A1(n9696), .A2(n15101), .ZN(n15102) );
  NAND2_X1 U18365 ( .A1(n15096), .A2(n15102), .ZN(n15584) );
  AOI21_X1 U18366 ( .B1(n15105), .B2(n15103), .A(n15104), .ZN(n15171) );
  NAND2_X1 U18367 ( .A1(n15171), .A2(n15119), .ZN(n15107) );
  NAND2_X1 U18368 ( .A1(n15122), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15106) );
  OAI211_X1 U18369 ( .C1(n15584), .C2(n15122), .A(n15107), .B(n15106), .ZN(
        P2_U2865) );
  OAI21_X1 U18370 ( .B1(n15108), .B2(n15109), .A(n15103), .ZN(n15186) );
  MUX2_X1 U18371 ( .A(n15112), .B(n15111), .S(n15110), .Z(n15113) );
  OAI21_X1 U18372 ( .B1(n15186), .B2(n15114), .A(n15113), .ZN(P2_U2866) );
  NAND2_X1 U18373 ( .A1(n14195), .A2(n15115), .ZN(n15116) );
  NAND2_X1 U18374 ( .A1(n15117), .A2(n15116), .ZN(n18859) );
  AOI21_X1 U18375 ( .B1(n15118), .B2(n14198), .A(n15108), .ZN(n15187) );
  NAND2_X1 U18376 ( .A1(n15187), .A2(n15119), .ZN(n15121) );
  NAND2_X1 U18377 ( .A1(n15122), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n15120) );
  OAI211_X1 U18378 ( .C1(n18859), .C2(n15122), .A(n15121), .B(n15120), .ZN(
        P2_U2867) );
  INV_X1 U18379 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n15125) );
  AOI22_X1 U18380 ( .A1(n16235), .A2(n15123), .B1(n19015), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n15124) );
  OAI21_X1 U18381 ( .B1(n15132), .B2(n15125), .A(n15124), .ZN(n15127) );
  NOR2_X1 U18382 ( .A1(n15499), .A2(n15206), .ZN(n15126) );
  AOI211_X1 U18383 ( .C1(n18957), .C2(BUF1_REG_29__SCAN_IN), .A(n15127), .B(
        n15126), .ZN(n15128) );
  OAI21_X1 U18384 ( .B1(n15129), .B2(n15185), .A(n15128), .ZN(P2_U2890) );
  AOI22_X1 U18385 ( .A1(n16235), .A2(n15130), .B1(n19015), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n15131) );
  OAI21_X1 U18386 ( .B1(n15132), .B2(n18183), .A(n15131), .ZN(n15138) );
  NOR2_X1 U18387 ( .A1(n15134), .A2(n15133), .ZN(n15135) );
  OR2_X1 U18388 ( .A1(n15136), .A2(n15135), .ZN(n16194) );
  NOR2_X1 U18389 ( .A1(n16194), .A2(n15206), .ZN(n15137) );
  AOI211_X1 U18390 ( .C1(n18957), .C2(BUF1_REG_28__SCAN_IN), .A(n15138), .B(
        n15137), .ZN(n15139) );
  OAI21_X1 U18391 ( .B1(n15140), .B2(n15185), .A(n15139), .ZN(P2_U2891) );
  OAI22_X1 U18392 ( .A1(n15156), .A2(n18971), .B1(n19014), .B2(n15141), .ZN(
        n15142) );
  AOI21_X1 U18393 ( .B1(n18955), .B2(BUF2_REG_27__SCAN_IN), .A(n15142), .ZN(
        n15144) );
  AOI22_X1 U18394 ( .A1(n15526), .A2(n19016), .B1(n18957), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15143) );
  OAI211_X1 U18395 ( .C1(n15145), .C2(n15185), .A(n15144), .B(n15143), .ZN(
        P2_U2892) );
  NAND2_X1 U18396 ( .A1(n9712), .A2(n15146), .ZN(n15147) );
  NAND2_X1 U18397 ( .A1(n15148), .A2(n15147), .ZN(n16207) );
  AOI22_X1 U18398 ( .A1(n16235), .A2(n15149), .B1(n19015), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15151) );
  AOI22_X1 U18399 ( .A1(n18957), .A2(BUF1_REG_26__SCAN_IN), .B1(n18955), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n15150) );
  OAI211_X1 U18400 ( .C1(n16207), .C2(n15206), .A(n15151), .B(n15150), .ZN(
        n15152) );
  AOI21_X1 U18401 ( .B1(n15153), .B2(n19017), .A(n15152), .ZN(n15154) );
  INV_X1 U18402 ( .A(n15154), .ZN(P2_U2893) );
  OAI22_X1 U18403 ( .A1(n15156), .A2(n18976), .B1(n19014), .B2(n15155), .ZN(
        n15159) );
  INV_X1 U18404 ( .A(n18957), .ZN(n15157) );
  INV_X1 U18405 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16395) );
  OAI22_X1 U18406 ( .A1(n15550), .A2(n15206), .B1(n15157), .B2(n16395), .ZN(
        n15158) );
  AOI211_X1 U18407 ( .C1(n18955), .C2(BUF2_REG_25__SCAN_IN), .A(n15159), .B(
        n15158), .ZN(n15160) );
  OAI21_X1 U18408 ( .B1(n15161), .B2(n15185), .A(n15160), .ZN(P2_U2894) );
  NOR2_X1 U18409 ( .A1(n15162), .A2(n15163), .ZN(n15164) );
  OR2_X1 U18410 ( .A1(n14978), .A2(n15164), .ZN(n16218) );
  AOI22_X1 U18411 ( .A1(n16235), .A2(n15165), .B1(n19015), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n15167) );
  AOI22_X1 U18412 ( .A1(n18957), .A2(BUF1_REG_23__SCAN_IN), .B1(n18955), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n15166) );
  OAI211_X1 U18413 ( .C1(n16218), .C2(n15206), .A(n15167), .B(n15166), .ZN(
        n15168) );
  INV_X1 U18414 ( .A(n15168), .ZN(n15169) );
  OAI21_X1 U18415 ( .B1(n15170), .B2(n15185), .A(n15169), .ZN(P2_U2896) );
  NAND2_X1 U18416 ( .A1(n15171), .A2(n19017), .ZN(n15179) );
  AOI22_X1 U18417 ( .A1(n16235), .A2(n15172), .B1(n19015), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n15178) );
  AOI22_X1 U18418 ( .A1(n18957), .A2(BUF1_REG_22__SCAN_IN), .B1(n18955), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n15177) );
  AND2_X1 U18419 ( .A1(n15174), .A2(n15173), .ZN(n15175) );
  NOR2_X1 U18420 ( .A1(n15162), .A2(n15175), .ZN(n15802) );
  NAND2_X1 U18421 ( .A1(n15802), .A2(n19016), .ZN(n15176) );
  NAND4_X1 U18422 ( .A1(n15179), .A2(n15178), .A3(n15177), .A4(n15176), .ZN(
        P2_U2897) );
  NAND2_X1 U18423 ( .A1(n16235), .A2(n18984), .ZN(n15180) );
  OAI21_X1 U18424 ( .B1(n19014), .B2(n15181), .A(n15180), .ZN(n15182) );
  AOI21_X1 U18425 ( .B1(n15597), .B2(n19016), .A(n15182), .ZN(n15184) );
  AOI22_X1 U18426 ( .A1(n18957), .A2(BUF1_REG_21__SCAN_IN), .B1(n18955), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n15183) );
  OAI211_X1 U18427 ( .C1(n15186), .C2(n15185), .A(n15184), .B(n15183), .ZN(
        P2_U2898) );
  NAND2_X1 U18428 ( .A1(n15187), .A2(n19017), .ZN(n15195) );
  AOI22_X1 U18429 ( .A1(n16235), .A2(n15188), .B1(n19015), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n15194) );
  AOI22_X1 U18430 ( .A1(n18957), .A2(BUF1_REG_20__SCAN_IN), .B1(n18955), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n15193) );
  OR2_X1 U18431 ( .A1(n15190), .A2(n15189), .ZN(n15191) );
  AND2_X1 U18432 ( .A1(n14993), .A2(n15191), .ZN(n18857) );
  NAND2_X1 U18433 ( .A1(n18857), .A2(n19016), .ZN(n15192) );
  NAND4_X1 U18434 ( .A1(n15195), .A2(n15194), .A3(n15193), .A4(n15192), .ZN(
        P2_U2899) );
  XNOR2_X1 U18435 ( .A(n15197), .B(n15196), .ZN(n18871) );
  AOI22_X1 U18436 ( .A1(n18957), .A2(BUF1_REG_18__SCAN_IN), .B1(n18955), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n15200) );
  AOI22_X1 U18437 ( .A1(n16235), .A2(n15198), .B1(n19015), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n15199) );
  OAI211_X1 U18438 ( .C1(n18871), .C2(n15206), .A(n15200), .B(n15199), .ZN(
        n15201) );
  AOI21_X1 U18439 ( .B1(n15202), .B2(n19017), .A(n15201), .ZN(n15203) );
  INV_X1 U18440 ( .A(n15203), .ZN(P2_U2901) );
  AOI22_X1 U18441 ( .A1(n18957), .A2(BUF1_REG_17__SCAN_IN), .B1(n18955), .B2(
        BUF2_REG_17__SCAN_IN), .ZN(n15205) );
  AOI22_X1 U18442 ( .A1(n16235), .A2(n19011), .B1(n19015), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n15204) );
  OAI211_X1 U18443 ( .C1(n15206), .C2(n15650), .A(n15205), .B(n15204), .ZN(
        n15207) );
  AOI21_X1 U18444 ( .B1(n15208), .B2(n19017), .A(n15207), .ZN(n15209) );
  INV_X1 U18445 ( .A(n15209), .ZN(P2_U2902) );
  NOR2_X2 U18446 ( .A1(n15230), .A2(n15480), .ZN(n15210) );
  XNOR2_X1 U18447 ( .A(n15210), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15478) );
  NAND2_X1 U18448 ( .A1(n15217), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n15214) );
  XNOR2_X1 U18449 ( .A(n15216), .B(n15214), .ZN(n16181) );
  NAND2_X1 U18450 ( .A1(n16181), .A2(n15220), .ZN(n15215) );
  NAND2_X1 U18451 ( .A1(n15215), .A2(n15480), .ZN(n15232) );
  OR2_X1 U18452 ( .A1(n15215), .A2(n15480), .ZN(n15233) );
  NOR2_X1 U18453 ( .A1(n15216), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n15218) );
  MUX2_X1 U18454 ( .A(n15219), .B(n15218), .S(n15217), .Z(n16173) );
  NAND2_X1 U18455 ( .A1(n16173), .A2(n15220), .ZN(n15221) );
  XNOR2_X1 U18456 ( .A(n15221), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15222) );
  XNOR2_X1 U18457 ( .A(n15223), .B(n15222), .ZN(n15474) );
  NAND2_X1 U18458 ( .A1(n13328), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n15452) );
  NAND2_X1 U18459 ( .A1(n19069), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15224) );
  OAI211_X1 U18460 ( .C1(n16262), .C2(n15225), .A(n15452), .B(n15224), .ZN(
        n15226) );
  AOI21_X1 U18461 ( .B1(n16175), .B2(n19078), .A(n15226), .ZN(n15227) );
  OAI21_X1 U18462 ( .B1(n15474), .B2(n19072), .A(n15227), .ZN(n15228) );
  INV_X1 U18463 ( .A(n15228), .ZN(n15229) );
  OAI21_X1 U18464 ( .B1(n15478), .B2(n19075), .A(n15229), .ZN(P2_U2983) );
  NAND2_X1 U18465 ( .A1(n15233), .A2(n15232), .ZN(n15234) );
  XNOR2_X1 U18466 ( .A(n15237), .B(n15236), .ZN(n16184) );
  NAND2_X1 U18467 ( .A1(n13328), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15481) );
  NAND2_X1 U18468 ( .A1(n19069), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15238) );
  OAI211_X1 U18469 ( .C1(n16262), .C2(n16184), .A(n15481), .B(n15238), .ZN(
        n15239) );
  NOR2_X1 U18470 ( .A1(n15241), .A2(n15240), .ZN(n15245) );
  NAND2_X1 U18471 ( .A1(n15243), .A2(n15242), .ZN(n15244) );
  XOR2_X1 U18472 ( .A(n15245), .B(n15244), .Z(n15257) );
  AOI22_X1 U18473 ( .A1(n15257), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n15245), .B2(n15244), .ZN(n15248) );
  XOR2_X1 U18474 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n15246), .Z(
        n15247) );
  XNOR2_X1 U18475 ( .A(n15248), .B(n15247), .ZN(n15522) );
  AOI21_X1 U18476 ( .B1(n15517), .B2(n15249), .A(n15250), .ZN(n15520) );
  INV_X1 U18477 ( .A(n16199), .ZN(n15253) );
  INV_X1 U18478 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15251) );
  NAND2_X1 U18479 ( .A1(n13328), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15511) );
  OAI21_X1 U18480 ( .B1(n19067), .B2(n15251), .A(n15511), .ZN(n15252) );
  AOI21_X1 U18481 ( .B1(n19059), .B2(n15253), .A(n15252), .ZN(n15254) );
  OAI21_X1 U18482 ( .B1(n16195), .B2(n16272), .A(n15254), .ZN(n15255) );
  AOI21_X1 U18483 ( .B1(n15520), .B2(n16251), .A(n15255), .ZN(n15256) );
  OAI21_X1 U18484 ( .B1(n15522), .B2(n19072), .A(n15256), .ZN(P2_U2986) );
  XNOR2_X1 U18485 ( .A(n15257), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15534) );
  INV_X1 U18486 ( .A(n15249), .ZN(n15259) );
  AOI21_X1 U18487 ( .B1(n15523), .B2(n15258), .A(n15259), .ZN(n15532) );
  NOR2_X1 U18488 ( .A1(n15529), .A2(n16272), .ZN(n15263) );
  NAND2_X1 U18489 ( .A1(n13328), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15524) );
  NAND2_X1 U18490 ( .A1(n19069), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15260) );
  OAI211_X1 U18491 ( .C1(n16262), .C2(n15261), .A(n15524), .B(n15260), .ZN(
        n15262) );
  AOI211_X1 U18492 ( .C1(n15532), .C2(n16251), .A(n15263), .B(n15262), .ZN(
        n15264) );
  OAI21_X1 U18493 ( .B1(n15534), .B2(n19072), .A(n15264), .ZN(P2_U2987) );
  BUF_X1 U18494 ( .A(n15265), .Z(n15266) );
  OAI21_X1 U18495 ( .B1(n15266), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15258), .ZN(n15546) );
  INV_X1 U18496 ( .A(n15276), .ZN(n15268) );
  OAI21_X1 U18497 ( .B1(n15267), .B2(n15268), .A(n15275), .ZN(n15269) );
  XOR2_X1 U18498 ( .A(n15270), .B(n15269), .Z(n15535) );
  NAND2_X1 U18499 ( .A1(n15535), .A2(n16250), .ZN(n15274) );
  INV_X1 U18500 ( .A(n15538), .ZN(n16209) );
  NAND2_X1 U18501 ( .A1(n18939), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15539) );
  NAND2_X1 U18502 ( .A1(n19069), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15271) );
  OAI211_X1 U18503 ( .C1(n16262), .C2(n16212), .A(n15539), .B(n15271), .ZN(
        n15272) );
  AOI21_X1 U18504 ( .B1(n16209), .B2(n19078), .A(n15272), .ZN(n15273) );
  OAI211_X1 U18505 ( .C1(n15546), .C2(n19075), .A(n15274), .B(n15273), .ZN(
        P2_U2988) );
  NAND2_X1 U18506 ( .A1(n15276), .A2(n15275), .ZN(n15277) );
  XNOR2_X1 U18507 ( .A(n15267), .B(n15277), .ZN(n15558) );
  INV_X1 U18508 ( .A(n15278), .ZN(n15552) );
  INV_X1 U18509 ( .A(n15279), .ZN(n15280) );
  NAND2_X1 U18510 ( .A1(n19059), .A2(n15280), .ZN(n15281) );
  NAND2_X1 U18511 ( .A1(n13328), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15548) );
  OAI211_X1 U18512 ( .C1(n19067), .C2(n15282), .A(n15281), .B(n15548), .ZN(
        n15286) );
  INV_X1 U18513 ( .A(n15283), .ZN(n15284) );
  NOR3_X1 U18514 ( .A1(n15547), .A2(n15266), .A3(n19075), .ZN(n15285) );
  AOI211_X1 U18515 ( .C1(n19078), .C2(n15552), .A(n15286), .B(n15285), .ZN(
        n15287) );
  OAI21_X1 U18516 ( .B1(n19072), .B2(n15558), .A(n15287), .ZN(P2_U2989) );
  NAND2_X1 U18518 ( .A1(n15342), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15312) );
  NOR2_X1 U18519 ( .A1(n15312), .A2(n15574), .ZN(n15300) );
  OAI21_X1 U18520 ( .B1(n15300), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15283), .ZN(n15569) );
  INV_X1 U18521 ( .A(n15291), .ZN(n15293) );
  NAND2_X1 U18522 ( .A1(n15293), .A2(n15292), .ZN(n15294) );
  XNOR2_X1 U18523 ( .A(n15290), .B(n15294), .ZN(n15567) );
  NOR2_X1 U18524 ( .A1(n18925), .A2(n19684), .ZN(n15562) );
  NOR2_X1 U18525 ( .A1(n16262), .A2(n15295), .ZN(n15296) );
  AOI211_X1 U18526 ( .C1(n19069), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15562), .B(n15296), .ZN(n15297) );
  OAI21_X1 U18527 ( .B1(n15564), .B2(n16272), .A(n15297), .ZN(n15298) );
  AOI21_X1 U18528 ( .B1(n15567), .B2(n16250), .A(n15298), .ZN(n15299) );
  OAI21_X1 U18529 ( .B1(n15569), .B2(n19075), .A(n15299), .ZN(P2_U2990) );
  INV_X1 U18530 ( .A(n15312), .ZN(n15302) );
  INV_X1 U18531 ( .A(n15300), .ZN(n15301) );
  OAI21_X1 U18532 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15302), .A(
        n15301), .ZN(n15583) );
  NAND2_X1 U18533 ( .A1(n13328), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15575) );
  OAI21_X1 U18534 ( .B1(n19067), .B2(n15303), .A(n15575), .ZN(n15305) );
  NOR2_X1 U18535 ( .A1(n15572), .A2(n16272), .ZN(n15304) );
  AOI211_X1 U18536 ( .C1(n19059), .C2(n15306), .A(n15305), .B(n15304), .ZN(
        n15311) );
  OR2_X1 U18537 ( .A1(n15308), .A2(n15307), .ZN(n15571) );
  NAND3_X1 U18538 ( .A1(n15571), .A2(n15309), .A3(n16250), .ZN(n15310) );
  OAI211_X1 U18539 ( .C1(n15583), .C2(n19075), .A(n15311), .B(n15310), .ZN(
        P2_U2991) );
  OAI21_X1 U18540 ( .B1(n15342), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15312), .ZN(n15594) );
  NAND2_X1 U18541 ( .A1(n15315), .A2(n15314), .ZN(n15316) );
  XNOR2_X1 U18542 ( .A(n15313), .B(n15316), .ZN(n15592) );
  NOR2_X1 U18543 ( .A1(n15584), .A2(n16272), .ZN(n15319) );
  NAND2_X1 U18544 ( .A1(n13328), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n15585) );
  NAND2_X1 U18545 ( .A1(n19069), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15317) );
  OAI211_X1 U18546 ( .C1(n16262), .C2(n15806), .A(n15585), .B(n15317), .ZN(
        n15318) );
  AOI211_X1 U18547 ( .C1(n15592), .C2(n16250), .A(n15319), .B(n15318), .ZN(
        n15320) );
  OAI21_X1 U18548 ( .B1(n15594), .B2(n19075), .A(n15320), .ZN(P2_U2992) );
  INV_X1 U18549 ( .A(n15423), .ZN(n15321) );
  NAND3_X1 U18550 ( .A1(n15323), .A2(n9699), .A3(n15416), .ZN(n15324) );
  OAI21_X1 U18551 ( .B1(n15325), .B2(n15324), .A(n15417), .ZN(n15407) );
  INV_X1 U18552 ( .A(n15404), .ZN(n15326) );
  INV_X1 U18553 ( .A(n15394), .ZN(n15327) );
  INV_X1 U18554 ( .A(n15328), .ZN(n15388) );
  NAND2_X1 U18555 ( .A1(n15331), .A2(n15330), .ZN(n15380) );
  NAND2_X1 U18556 ( .A1(n9598), .A2(n15332), .ZN(n15347) );
  INV_X1 U18557 ( .A(n15348), .ZN(n15333) );
  NAND2_X1 U18558 ( .A1(n15336), .A2(n15335), .ZN(n15337) );
  XNOR2_X1 U18559 ( .A(n15338), .B(n15337), .ZN(n15607) );
  NOR2_X1 U18560 ( .A1(n18925), .A2(n20763), .ZN(n15596) );
  AOI21_X1 U18561 ( .B1(n19069), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15596), .ZN(n15339) );
  OAI21_X1 U18562 ( .B1(n16262), .B2(n15340), .A(n15339), .ZN(n15344) );
  NOR2_X1 U18563 ( .A1(n15289), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15341) );
  OR2_X1 U18564 ( .A1(n15342), .A2(n15341), .ZN(n15601) );
  NOR2_X1 U18565 ( .A1(n15601), .A2(n19075), .ZN(n15343) );
  OAI21_X1 U18566 ( .B1(n15607), .B2(n19072), .A(n15345), .ZN(P2_U2993) );
  NAND2_X1 U18567 ( .A1(n15347), .A2(n15346), .ZN(n15351) );
  NAND2_X1 U18568 ( .A1(n15349), .A2(n15348), .ZN(n15350) );
  XNOR2_X1 U18569 ( .A(n15351), .B(n15350), .ZN(n15620) );
  INV_X1 U18570 ( .A(n15352), .ZN(n15353) );
  NAND2_X1 U18571 ( .A1(n15353), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15622) );
  AOI21_X1 U18572 ( .B1(n15612), .B2(n15622), .A(n15289), .ZN(n15618) );
  NOR2_X1 U18573 ( .A1(n18925), .A2(n19677), .ZN(n15614) );
  NOR2_X1 U18574 ( .A1(n16262), .A2(n18863), .ZN(n15354) );
  AOI211_X1 U18575 ( .C1(n19069), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15614), .B(n15354), .ZN(n15355) );
  OAI21_X1 U18576 ( .B1(n18859), .B2(n16272), .A(n15355), .ZN(n15356) );
  AOI21_X1 U18577 ( .B1(n15618), .B2(n16251), .A(n15356), .ZN(n15357) );
  OAI21_X1 U18578 ( .B1(n15620), .B2(n19072), .A(n15357), .ZN(P2_U2994) );
  NAND2_X1 U18579 ( .A1(n15359), .A2(n15358), .ZN(n15362) );
  INV_X1 U18580 ( .A(n15372), .ZN(n15360) );
  XOR2_X1 U18581 ( .A(n15362), .B(n15361), .Z(n15634) );
  NOR2_X1 U18582 ( .A1(n15363), .A2(n16262), .ZN(n15366) );
  NAND2_X1 U18583 ( .A1(n18939), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15623) );
  OAI21_X1 U18584 ( .B1(n19067), .B2(n15364), .A(n15623), .ZN(n15365) );
  AOI211_X1 U18585 ( .C1(n15628), .C2(n19078), .A(n15366), .B(n15365), .ZN(
        n15368) );
  NAND2_X1 U18586 ( .A1(n15352), .A2(n20778), .ZN(n15621) );
  NAND3_X1 U18587 ( .A1(n15622), .A2(n16251), .A3(n15621), .ZN(n15367) );
  OAI211_X1 U18588 ( .C1(n15634), .C2(n19072), .A(n15368), .B(n15367), .ZN(
        P2_U2995) );
  NAND2_X1 U18589 ( .A1(n15369), .A2(n15610), .ZN(n15370) );
  NAND2_X1 U18590 ( .A1(n15352), .A2(n15370), .ZN(n15645) );
  NAND2_X1 U18591 ( .A1(n15372), .A2(n15371), .ZN(n15374) );
  XOR2_X1 U18592 ( .A(n15374), .B(n9599), .Z(n15635) );
  NAND2_X1 U18593 ( .A1(n15635), .A2(n16250), .ZN(n15378) );
  INV_X1 U18594 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19673) );
  OAI22_X1 U18595 ( .A1(n19673), .A2(n16290), .B1(n16262), .B2(n18876), .ZN(
        n15376) );
  NOR2_X1 U18596 ( .A1(n18872), .A2(n16272), .ZN(n15375) );
  AOI211_X1 U18597 ( .C1(n19069), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15376), .B(n15375), .ZN(n15377) );
  OAI211_X1 U18598 ( .C1(n19075), .C2(n15645), .A(n15378), .B(n15377), .ZN(
        P2_U2996) );
  XOR2_X1 U18599 ( .A(n15380), .B(n15379), .Z(n15664) );
  NAND2_X1 U18600 ( .A1(n18939), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15648) );
  NAND2_X1 U18601 ( .A1(n19069), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15381) );
  OAI211_X1 U18602 ( .C1(n15382), .C2(n16262), .A(n15648), .B(n15381), .ZN(
        n15383) );
  AOI21_X1 U18603 ( .B1(n15647), .B2(n19078), .A(n15383), .ZN(n15387) );
  INV_X1 U18604 ( .A(n15384), .ZN(n16244) );
  NAND2_X1 U18605 ( .A1(n16244), .A2(n15656), .ZN(n15408) );
  NOR2_X2 U18606 ( .A1(n15408), .A2(n15682), .ZN(n15398) );
  NAND2_X1 U18607 ( .A1(n15398), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15654) );
  INV_X1 U18608 ( .A(n15654), .ZN(n15385) );
  OAI211_X1 U18609 ( .C1(n15385), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16251), .B(n15369), .ZN(n15386) );
  OAI211_X1 U18610 ( .C1(n15664), .C2(n19072), .A(n15387), .B(n15386), .ZN(
        P2_U2997) );
  XNOR2_X1 U18611 ( .A(n15389), .B(n15388), .ZN(n15673) );
  OAI211_X1 U18612 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15398), .A(
        n9596), .B(n16251), .ZN(n15393) );
  NAND2_X1 U18613 ( .A1(n18939), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n15665) );
  NAND2_X1 U18614 ( .A1(n19069), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15390) );
  OAI211_X1 U18615 ( .C1(n16262), .C2(n18887), .A(n15665), .B(n15390), .ZN(
        n15391) );
  AOI21_X1 U18616 ( .B1(n18885), .B2(n19078), .A(n15391), .ZN(n15392) );
  OAI211_X1 U18617 ( .C1(n15673), .C2(n19072), .A(n15393), .B(n15392), .ZN(
        P2_U2998) );
  NAND2_X1 U18618 ( .A1(n15395), .A2(n15394), .ZN(n15397) );
  XOR2_X1 U18619 ( .A(n15397), .B(n15396), .Z(n15686) );
  AOI21_X1 U18620 ( .B1(n15682), .B2(n15408), .A(n15398), .ZN(n15674) );
  NAND2_X1 U18621 ( .A1(n15674), .A2(n16251), .ZN(n15403) );
  NAND2_X1 U18622 ( .A1(n18939), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n15678) );
  NAND2_X1 U18623 ( .A1(n19069), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15399) );
  OAI211_X1 U18624 ( .C1(n15400), .C2(n16262), .A(n15678), .B(n15399), .ZN(
        n15401) );
  AOI21_X1 U18625 ( .B1(n15677), .B2(n19078), .A(n15401), .ZN(n15402) );
  OAI211_X1 U18626 ( .C1(n15686), .C2(n19072), .A(n15403), .B(n15402), .ZN(
        P2_U2999) );
  NAND2_X1 U18627 ( .A1(n15405), .A2(n15404), .ZN(n15406) );
  XNOR2_X1 U18628 ( .A(n15407), .B(n15406), .ZN(n15701) );
  NAND2_X1 U18629 ( .A1(n16244), .A2(n15692), .ZN(n15414) );
  INV_X1 U18630 ( .A(n15408), .ZN(n15666) );
  AOI21_X1 U18631 ( .B1(n15691), .B2(n15414), .A(n15666), .ZN(n15687) );
  NAND2_X1 U18632 ( .A1(n15687), .A2(n16251), .ZN(n15413) );
  INV_X1 U18633 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19666) );
  OAI22_X1 U18634 ( .A1(n15409), .A2(n19067), .B1(n19666), .B2(n16290), .ZN(
        n15411) );
  NOR2_X1 U18635 ( .A1(n18900), .A2(n16272), .ZN(n15410) );
  AOI211_X1 U18636 ( .C1(n19059), .C2(n18895), .A(n15411), .B(n15410), .ZN(
        n15412) );
  OAI211_X1 U18637 ( .C1(n19072), .C2(n15701), .A(n15413), .B(n15412), .ZN(
        P2_U3000) );
  NOR2_X1 U18638 ( .A1(n15384), .A2(n15726), .ZN(n15716) );
  OAI21_X1 U18639 ( .B1(n15716), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15414), .ZN(n15714) );
  AND2_X1 U18640 ( .A1(n18939), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n15706) );
  INV_X1 U18641 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18918) );
  OAI22_X1 U18642 ( .A1(n18918), .A2(n19067), .B1(n16262), .B2(n18912), .ZN(
        n15415) );
  AOI211_X1 U18643 ( .C1(n19078), .C2(n15707), .A(n15706), .B(n15415), .ZN(
        n15421) );
  NAND2_X1 U18644 ( .A1(n15417), .A2(n15416), .ZN(n15419) );
  XOR2_X1 U18645 ( .A(n15419), .B(n15418), .Z(n15712) );
  NAND2_X1 U18646 ( .A1(n15712), .A2(n16250), .ZN(n15420) );
  OAI211_X1 U18647 ( .C1(n15714), .C2(n19075), .A(n15421), .B(n15420), .ZN(
        P2_U3001) );
  NAND2_X1 U18648 ( .A1(n15384), .A2(n15726), .ZN(n15717) );
  NAND2_X1 U18649 ( .A1(n15717), .A2(n16251), .ZN(n15431) );
  NAND2_X1 U18650 ( .A1(n9699), .A2(n15423), .ZN(n15424) );
  XNOR2_X1 U18651 ( .A(n15422), .B(n15424), .ZN(n15715) );
  OAI22_X1 U18652 ( .A1(n15425), .A2(n19067), .B1(n12749), .B2(n18925), .ZN(
        n15429) );
  INV_X1 U18653 ( .A(n15426), .ZN(n15427) );
  OAI22_X1 U18654 ( .A1(n15724), .A2(n16272), .B1(n16262), .B2(n15427), .ZN(
        n15428) );
  AOI211_X1 U18655 ( .C1(n15715), .C2(n16250), .A(n15429), .B(n15428), .ZN(
        n15430) );
  OAI21_X1 U18656 ( .B1(n15716), .B2(n15431), .A(n15430), .ZN(P2_U3002) );
  NAND2_X1 U18657 ( .A1(n14160), .A2(n15432), .ZN(n15434) );
  NAND2_X1 U18658 ( .A1(n15434), .A2(n15433), .ZN(n15438) );
  AND2_X1 U18659 ( .A1(n15436), .A2(n15435), .ZN(n15437) );
  XNOR2_X1 U18660 ( .A(n15438), .B(n15437), .ZN(n15761) );
  NAND2_X1 U18661 ( .A1(n15441), .A2(n15440), .ZN(n15747) );
  NAND3_X1 U18662 ( .A1(n15439), .A2(n15747), .A3(n16251), .ZN(n15447) );
  NOR2_X1 U18663 ( .A1(n15748), .A2(n16272), .ZN(n15444) );
  OAI22_X1 U18664 ( .A1(n15442), .A2(n19067), .B1(n12736), .B2(n16290), .ZN(
        n15443) );
  AOI211_X1 U18665 ( .C1(n19059), .C2(n15445), .A(n15444), .B(n15443), .ZN(
        n15446) );
  OAI211_X1 U18666 ( .C1(n15761), .C2(n19072), .A(n15447), .B(n15446), .ZN(
        P2_U3006) );
  AOI222_X1 U18667 ( .A1(n12712), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12770), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C1(n12795), .C2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n15448) );
  NAND2_X1 U18668 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15750) );
  NOR2_X1 U18669 ( .A1(n15750), .A2(n15752), .ZN(n16292) );
  NAND2_X1 U18670 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16292), .ZN(
        n16273) );
  INV_X1 U18671 ( .A(n16273), .ZN(n15450) );
  NAND2_X1 U18672 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15464) );
  INV_X1 U18673 ( .A(n15464), .ZN(n16274) );
  NAND2_X1 U18674 ( .A1(n15450), .A2(n16274), .ZN(n15690) );
  NAND2_X1 U18675 ( .A1(n10913), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15451) );
  NOR2_X1 U18676 ( .A1(n15631), .A2(n15458), .ZN(n15605) );
  NAND2_X1 U18677 ( .A1(n15605), .A2(n15465), .ZN(n15554) );
  NAND2_X1 U18678 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15455) );
  OR2_X1 U18679 ( .A1(n15554), .A2(n15455), .ZN(n15494) );
  NOR2_X1 U18680 ( .A1(n15494), .A2(n15468), .ZN(n15497) );
  INV_X1 U18681 ( .A(n15452), .ZN(n15453) );
  INV_X1 U18682 ( .A(n15455), .ZN(n15456) );
  OR2_X1 U18683 ( .A1(n15554), .A2(n15456), .ZN(n15467) );
  NAND2_X1 U18684 ( .A1(n15457), .A2(n15660), .ZN(n15740) );
  INV_X1 U18685 ( .A(n15458), .ZN(n15608) );
  NAND3_X1 U18686 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(n15459), .ZN(n15460) );
  NAND2_X1 U18687 ( .A1(n15611), .A2(n15460), .ZN(n15463) );
  AND2_X1 U18688 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15461), .ZN(
        n15462) );
  NAND2_X1 U18689 ( .A1(n15463), .A2(n15462), .ZN(n16293) );
  NOR2_X1 U18690 ( .A1(n15636), .A2(n15719), .ZN(n15609) );
  NAND4_X1 U18691 ( .A1(n15465), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15608), .A4(n15609), .ZN(n15466) );
  NAND2_X1 U18692 ( .A1(n15740), .A2(n15466), .ZN(n15560) );
  OAI21_X1 U18693 ( .B1(n15468), .B2(n15496), .A(n15611), .ZN(n15469) );
  NAND2_X1 U18694 ( .A1(n15536), .A2(n15469), .ZN(n15483) );
  AOI21_X1 U18695 ( .B1(n15480), .B2(n15611), .A(n15483), .ZN(n15471) );
  NOR2_X1 U18696 ( .A1(n15471), .A2(n15470), .ZN(n15472) );
  AOI211_X1 U18697 ( .C1(n15757), .C2(n16175), .A(n15473), .B(n15472), .ZN(
        n15477) );
  INV_X1 U18698 ( .A(n15474), .ZN(n15475) );
  NAND2_X1 U18699 ( .A1(n15475), .A2(n16281), .ZN(n15476) );
  OAI211_X1 U18700 ( .C1(n15478), .C2(n16308), .A(n15477), .B(n15476), .ZN(
        P2_U3015) );
  NAND3_X1 U18701 ( .A1(n15497), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15480), .ZN(n15485) );
  INV_X1 U18702 ( .A(n15481), .ZN(n15482) );
  OAI21_X1 U18703 ( .B1(n15235), .B2(n16315), .A(n15488), .ZN(n15489) );
  OAI21_X1 U18704 ( .B1(n15492), .B2(n16308), .A(n15491), .ZN(P2_U3016) );
  INV_X1 U18705 ( .A(n15494), .ZN(n15493) );
  NAND2_X1 U18706 ( .A1(n15493), .A2(n15523), .ZN(n15528) );
  AND2_X1 U18707 ( .A1(n15528), .A2(n15536), .ZN(n15518) );
  OR2_X1 U18708 ( .A1(n15494), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15512) );
  AOI21_X1 U18709 ( .B1(n15518), .B2(n15512), .A(n15496), .ZN(n15495) );
  INV_X1 U18710 ( .A(n15495), .ZN(n15506) );
  NAND2_X1 U18711 ( .A1(n15497), .A2(n15496), .ZN(n15502) );
  OAI21_X1 U18712 ( .B1(n15499), .B2(n16305), .A(n15498), .ZN(n15500) );
  INV_X1 U18713 ( .A(n15500), .ZN(n15501) );
  OAI211_X1 U18714 ( .C1(n16315), .C2(n15503), .A(n15502), .B(n15501), .ZN(
        n15504) );
  INV_X1 U18715 ( .A(n15504), .ZN(n15505) );
  OAI211_X1 U18716 ( .C1(n15507), .C2(n16308), .A(n15506), .B(n15505), .ZN(
        n15508) );
  INV_X1 U18717 ( .A(n15508), .ZN(n15509) );
  OAI21_X1 U18718 ( .B1(n15510), .B2(n16306), .A(n15509), .ZN(P2_U3017) );
  INV_X1 U18719 ( .A(n16195), .ZN(n15515) );
  NOR2_X1 U18720 ( .A1(n16194), .A2(n16305), .ZN(n15514) );
  OAI21_X1 U18721 ( .B1(n15512), .B2(n15523), .A(n15511), .ZN(n15513) );
  AOI211_X1 U18722 ( .C1(n15515), .C2(n15757), .A(n15514), .B(n15513), .ZN(
        n15516) );
  OAI21_X1 U18723 ( .B1(n15518), .B2(n15517), .A(n15516), .ZN(n15519) );
  AOI21_X1 U18724 ( .B1(n15520), .B2(n16282), .A(n15519), .ZN(n15521) );
  OAI21_X1 U18725 ( .B1(n15522), .B2(n16306), .A(n15521), .ZN(P2_U3018) );
  NOR2_X1 U18726 ( .A1(n15536), .A2(n15523), .ZN(n15531) );
  INV_X1 U18727 ( .A(n15524), .ZN(n15525) );
  AOI21_X1 U18728 ( .B1(n15526), .B2(n15739), .A(n15525), .ZN(n15527) );
  OAI211_X1 U18729 ( .C1(n15529), .C2(n16315), .A(n15528), .B(n15527), .ZN(
        n15530) );
  AOI211_X1 U18730 ( .C1(n15532), .C2(n16282), .A(n15531), .B(n15530), .ZN(
        n15533) );
  OAI21_X1 U18731 ( .B1(n15534), .B2(n16306), .A(n15533), .ZN(P2_U3019) );
  NAND2_X1 U18732 ( .A1(n15535), .A2(n16281), .ZN(n15545) );
  INV_X1 U18733 ( .A(n15536), .ZN(n15543) );
  OAI21_X1 U18734 ( .B1(n15554), .B2(n10914), .A(n15537), .ZN(n15542) );
  NOR2_X1 U18735 ( .A1(n15538), .A2(n16315), .ZN(n15541) );
  OAI21_X1 U18736 ( .B1(n16207), .B2(n16305), .A(n15539), .ZN(n15540) );
  AOI211_X1 U18737 ( .C1(n15543), .C2(n15542), .A(n15541), .B(n15540), .ZN(
        n15544) );
  OAI211_X1 U18738 ( .C1(n16308), .C2(n15546), .A(n15545), .B(n15544), .ZN(
        P2_U3020) );
  NOR3_X1 U18739 ( .A1(n15547), .A2(n15266), .A3(n16308), .ZN(n15556) );
  OR2_X1 U18740 ( .A1(n15560), .A2(n10914), .ZN(n15549) );
  OAI211_X1 U18741 ( .C1(n15550), .C2(n16305), .A(n15549), .B(n15548), .ZN(
        n15551) );
  AOI21_X1 U18742 ( .B1(n15552), .B2(n15757), .A(n15551), .ZN(n15553) );
  OAI21_X1 U18743 ( .B1(n15554), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15553), .ZN(n15555) );
  NOR2_X1 U18744 ( .A1(n15556), .A2(n15555), .ZN(n15557) );
  OAI21_X1 U18745 ( .B1(n16306), .B2(n15558), .A(n15557), .ZN(P2_U3021) );
  NAND2_X1 U18746 ( .A1(n15605), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15590) );
  NAND2_X1 U18747 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15570) );
  NOR3_X1 U18748 ( .A1(n15590), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15570), .ZN(n15566) );
  NOR2_X1 U18749 ( .A1(n15560), .A2(n15559), .ZN(n15561) );
  AOI211_X1 U18750 ( .C1(n16229), .C2(n15739), .A(n15562), .B(n15561), .ZN(
        n15563) );
  OAI21_X1 U18751 ( .B1(n15564), .B2(n16315), .A(n15563), .ZN(n15565) );
  AOI211_X1 U18752 ( .C1(n15567), .C2(n16281), .A(n15566), .B(n15565), .ZN(
        n15568) );
  OAI21_X1 U18753 ( .B1(n15569), .B2(n16308), .A(n15568), .ZN(P2_U3022) );
  OAI21_X1 U18754 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n15570), .ZN(n15580) );
  NAND3_X1 U18755 ( .A1(n15571), .A2(n15309), .A3(n16281), .ZN(n15579) );
  INV_X1 U18756 ( .A(n15572), .ZN(n16220) );
  NAND4_X1 U18757 ( .A1(n15608), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A4(n15609), .ZN(n15573) );
  NAND2_X1 U18758 ( .A1(n15740), .A2(n15573), .ZN(n15600) );
  OR2_X1 U18759 ( .A1(n15600), .A2(n15574), .ZN(n15576) );
  OAI211_X1 U18760 ( .C1(n16218), .C2(n16305), .A(n15576), .B(n15575), .ZN(
        n15577) );
  AOI21_X1 U18761 ( .B1(n16220), .B2(n15757), .A(n15577), .ZN(n15578) );
  OAI211_X1 U18762 ( .C1(n15580), .C2(n15590), .A(n15579), .B(n15578), .ZN(
        n15581) );
  INV_X1 U18763 ( .A(n15581), .ZN(n15582) );
  OAI21_X1 U18764 ( .B1(n15583), .B2(n16308), .A(n15582), .ZN(P2_U3023) );
  INV_X1 U18765 ( .A(n15584), .ZN(n15803) );
  NAND2_X1 U18766 ( .A1(n15802), .A2(n15739), .ZN(n15586) );
  OAI211_X1 U18767 ( .C1(n15600), .C2(n15587), .A(n15586), .B(n15585), .ZN(
        n15588) );
  AOI21_X1 U18768 ( .B1(n15803), .B2(n15757), .A(n15588), .ZN(n15589) );
  OAI21_X1 U18769 ( .B1(n15590), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15589), .ZN(n15591) );
  AOI21_X1 U18770 ( .B1(n15592), .B2(n16281), .A(n15591), .ZN(n15593) );
  OAI21_X1 U18771 ( .B1(n15594), .B2(n16308), .A(n15593), .ZN(P2_U3024) );
  NAND2_X1 U18772 ( .A1(n15595), .A2(n15757), .ZN(n15599) );
  AOI21_X1 U18773 ( .B1(n15597), .B2(n15739), .A(n15596), .ZN(n15598) );
  OAI211_X1 U18774 ( .C1(n15604), .C2(n15600), .A(n15599), .B(n15598), .ZN(
        n15603) );
  NOR2_X1 U18775 ( .A1(n15601), .A2(n16308), .ZN(n15602) );
  OAI21_X1 U18776 ( .B1(n15607), .B2(n16306), .A(n15606), .ZN(P2_U3025) );
  AOI211_X1 U18777 ( .C1(n15612), .C2(n20778), .A(n15608), .B(n15631), .ZN(
        n15617) );
  INV_X1 U18778 ( .A(n15740), .ZN(n15689) );
  NOR2_X1 U18779 ( .A1(n15689), .A2(n15609), .ZN(n15637) );
  AOI21_X1 U18780 ( .B1(n15611), .B2(n15610), .A(n15637), .ZN(n15626) );
  NOR2_X1 U18781 ( .A1(n15626), .A2(n15612), .ZN(n15613) );
  AOI211_X1 U18782 ( .C1(n15739), .C2(n18857), .A(n15614), .B(n15613), .ZN(
        n15615) );
  OAI21_X1 U18783 ( .B1(n18859), .B2(n16315), .A(n15615), .ZN(n15616) );
  AOI211_X1 U18784 ( .C1(n15618), .C2(n16282), .A(n15617), .B(n15616), .ZN(
        n15619) );
  OAI21_X1 U18785 ( .B1(n15620), .B2(n16306), .A(n15619), .ZN(P2_U3026) );
  NAND3_X1 U18786 ( .A1(n15622), .A2(n16282), .A3(n15621), .ZN(n15630) );
  INV_X1 U18787 ( .A(n15623), .ZN(n15624) );
  AOI21_X1 U18788 ( .B1(n15739), .B2(n16236), .A(n15624), .ZN(n15625) );
  OAI21_X1 U18789 ( .B1(n15626), .B2(n20778), .A(n15625), .ZN(n15627) );
  AOI21_X1 U18790 ( .B1(n15628), .B2(n15757), .A(n15627), .ZN(n15629) );
  OAI211_X1 U18791 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15631), .A(
        n15630), .B(n15629), .ZN(n15632) );
  INV_X1 U18792 ( .A(n15632), .ZN(n15633) );
  OAI21_X1 U18793 ( .B1(n15634), .B2(n16306), .A(n15633), .ZN(P2_U3027) );
  NAND2_X1 U18794 ( .A1(n15635), .A2(n16281), .ZN(n15644) );
  INV_X1 U18795 ( .A(n18872), .ZN(n15642) );
  NOR2_X1 U18796 ( .A1(n15636), .A2(n15690), .ZN(n15638) );
  MUX2_X1 U18797 ( .A(n15638), .B(n15637), .S(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .Z(n15639) );
  AOI21_X1 U18798 ( .B1(n18939), .B2(P2_REIP_REG_18__SCAN_IN), .A(n15639), 
        .ZN(n15640) );
  OAI21_X1 U18799 ( .B1(n16305), .B2(n18871), .A(n15640), .ZN(n15641) );
  AOI21_X1 U18800 ( .B1(n15642), .B2(n15757), .A(n15641), .ZN(n15643) );
  OAI211_X1 U18801 ( .C1(n15645), .C2(n16308), .A(n15644), .B(n15643), .ZN(
        P2_U3028) );
  INV_X1 U18802 ( .A(n15690), .ZN(n15727) );
  NAND2_X1 U18803 ( .A1(n15727), .A2(n15656), .ZN(n15675) );
  OAI22_X1 U18804 ( .A1(n9596), .A2(n16308), .B1(n15646), .B2(n15675), .ZN(
        n15653) );
  NAND2_X1 U18805 ( .A1(n15647), .A2(n15757), .ZN(n15649) );
  OAI211_X1 U18806 ( .C1(n16305), .C2(n15650), .A(n15649), .B(n15648), .ZN(
        n15651) );
  OAI21_X1 U18807 ( .B1(n16282), .B2(n15655), .A(n15654), .ZN(n15658) );
  INV_X1 U18808 ( .A(n15656), .ZN(n15657) );
  OAI21_X1 U18809 ( .B1(n15719), .B2(n15657), .A(n15740), .ZN(n15676) );
  OAI211_X1 U18810 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15659), .A(
        n15658), .B(n15676), .ZN(n15670) );
  NOR2_X1 U18811 ( .A1(n15660), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15661) );
  OAI21_X1 U18812 ( .B1(n15670), .B2(n15661), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15662) );
  OAI211_X1 U18813 ( .C1(n15664), .C2(n16306), .A(n15663), .B(n15662), .ZN(
        P2_U3029) );
  OAI21_X1 U18814 ( .B1(n16305), .B2(n18883), .A(n15665), .ZN(n15669) );
  NAND2_X1 U18815 ( .A1(n15666), .A2(n16282), .ZN(n15667) );
  AOI211_X1 U18816 ( .C1(n15667), .C2(n15675), .A(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n15682), .ZN(n15668) );
  AOI211_X1 U18817 ( .C1(n15757), .C2(n18885), .A(n15669), .B(n15668), .ZN(
        n15672) );
  NAND2_X1 U18818 ( .A1(n15670), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15671) );
  OAI211_X1 U18819 ( .C1(n16306), .C2(n15673), .A(n15672), .B(n15671), .ZN(
        P2_U3030) );
  NAND2_X1 U18820 ( .A1(n15674), .A2(n16282), .ZN(n15685) );
  INV_X1 U18821 ( .A(n15675), .ZN(n15683) );
  NOR2_X1 U18822 ( .A1(n15676), .A2(n15682), .ZN(n15681) );
  NAND2_X1 U18823 ( .A1(n15677), .A2(n15757), .ZN(n15679) );
  OAI211_X1 U18824 ( .C1(n16305), .C2(n18961), .A(n15679), .B(n15678), .ZN(
        n15680) );
  AOI211_X1 U18825 ( .C1(n15683), .C2(n15682), .A(n15681), .B(n15680), .ZN(
        n15684) );
  OAI211_X1 U18826 ( .C1(n15686), .C2(n16306), .A(n15685), .B(n15684), .ZN(
        P2_U3031) );
  NAND2_X1 U18827 ( .A1(n15687), .A2(n16282), .ZN(n15700) );
  INV_X1 U18828 ( .A(n15719), .ZN(n15688) );
  OAI22_X1 U18829 ( .A1(n15690), .A2(n15692), .B1(n15689), .B2(n15688), .ZN(
        n15702) );
  NAND3_X1 U18830 ( .A1(n15727), .A2(n15692), .A3(n15691), .ZN(n15697) );
  INV_X1 U18831 ( .A(n15032), .ZN(n15694) );
  AOI21_X1 U18832 ( .B1(n15695), .B2(n15693), .A(n15694), .ZN(n18962) );
  AOI22_X1 U18833 ( .A1(n15739), .A2(n18962), .B1(n18939), .B2(
        P2_REIP_REG_14__SCAN_IN), .ZN(n15696) );
  OAI211_X1 U18834 ( .C1(n18900), .C2(n16315), .A(n15697), .B(n15696), .ZN(
        n15698) );
  AOI21_X1 U18835 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15702), .A(
        n15698), .ZN(n15699) );
  OAI211_X1 U18836 ( .C1(n15701), .C2(n16306), .A(n15700), .B(n15699), .ZN(
        P2_U3032) );
  INV_X1 U18837 ( .A(n15702), .ZN(n15710) );
  AOI21_X1 U18838 ( .B1(n15727), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15709) );
  OR2_X1 U18839 ( .A1(n15703), .A2(n13936), .ZN(n15704) );
  NAND2_X1 U18840 ( .A1(n15693), .A2(n15704), .ZN(n18967) );
  NOR2_X1 U18841 ( .A1(n16305), .A2(n18967), .ZN(n15705) );
  AOI211_X1 U18842 ( .C1(n15707), .C2(n15757), .A(n15706), .B(n15705), .ZN(
        n15708) );
  OAI21_X1 U18843 ( .B1(n15710), .B2(n15709), .A(n15708), .ZN(n15711) );
  AOI21_X1 U18844 ( .B1(n15712), .B2(n16281), .A(n15711), .ZN(n15713) );
  OAI21_X1 U18845 ( .B1(n15714), .B2(n16308), .A(n15713), .ZN(P2_U3033) );
  INV_X1 U18846 ( .A(n15715), .ZN(n15730) );
  INV_X1 U18847 ( .A(n15716), .ZN(n15718) );
  NAND3_X1 U18848 ( .A1(n15718), .A2(n16282), .A3(n15717), .ZN(n15729) );
  NAND2_X1 U18849 ( .A1(n15740), .A2(n15719), .ZN(n15721) );
  NAND2_X1 U18850 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n13328), .ZN(n15720) );
  OAI21_X1 U18851 ( .B1(n15726), .B2(n15721), .A(n15720), .ZN(n15722) );
  AOI21_X1 U18852 ( .B1(n15739), .B2(n18968), .A(n15722), .ZN(n15723) );
  OAI21_X1 U18853 ( .B1(n15724), .B2(n16315), .A(n15723), .ZN(n15725) );
  AOI21_X1 U18854 ( .B1(n15727), .B2(n15726), .A(n15725), .ZN(n15728) );
  OAI211_X1 U18855 ( .C1(n15730), .C2(n16306), .A(n15729), .B(n15728), .ZN(
        P2_U3034) );
  INV_X1 U18856 ( .A(n15731), .ZN(n15732) );
  OAI21_X1 U18857 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n15732), .A(
        n9673), .ZN(n16256) );
  INV_X1 U18858 ( .A(n16266), .ZN(n15733) );
  NAND2_X1 U18859 ( .A1(n15734), .A2(n15733), .ZN(n15738) );
  NOR2_X1 U18860 ( .A1(n15736), .A2(n15735), .ZN(n15737) );
  XNOR2_X1 U18861 ( .A(n15738), .B(n15737), .ZN(n16255) );
  AOI22_X1 U18862 ( .A1(n16258), .A2(n15757), .B1(n15739), .B2(n18973), .ZN(
        n15744) );
  NAND2_X1 U18863 ( .A1(n15740), .A2(n16293), .ZN(n16277) );
  NAND2_X1 U18864 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n13328), .ZN(n15741) );
  OAI221_X1 U18865 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16273), 
        .C1(n16275), .C2(n16277), .A(n15741), .ZN(n15742) );
  INV_X1 U18866 ( .A(n15742), .ZN(n15743) );
  OAI211_X1 U18867 ( .C1(n16255), .C2(n16306), .A(n15744), .B(n15743), .ZN(
        n15745) );
  INV_X1 U18868 ( .A(n15745), .ZN(n15746) );
  OAI21_X1 U18869 ( .B1(n16256), .B2(n16308), .A(n15746), .ZN(P2_U3036) );
  NAND3_X1 U18870 ( .A1(n15439), .A2(n15747), .A3(n16282), .ZN(n15760) );
  INV_X1 U18871 ( .A(n15748), .ZN(n15758) );
  INV_X1 U18872 ( .A(n15749), .ZN(n18980) );
  OAI22_X1 U18873 ( .A1(n16305), .A2(n18980), .B1(n12736), .B2(n16290), .ZN(
        n15756) );
  OAI21_X1 U18874 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n15750), .ZN(n15751) );
  OAI22_X1 U18875 ( .A1(n15754), .A2(n15753), .B1(n15752), .B2(n15751), .ZN(
        n15755) );
  AOI211_X1 U18876 ( .C1(n15758), .C2(n15757), .A(n15756), .B(n15755), .ZN(
        n15759) );
  OAI211_X1 U18877 ( .C1(n15761), .C2(n16306), .A(n15760), .B(n15759), .ZN(
        P2_U3038) );
  INV_X1 U18878 ( .A(n15762), .ZN(n15765) );
  OAI222_X1 U18879 ( .A1(n15765), .A2(n15764), .B1(n19708), .B2(n15763), .C1(
        n16320), .C2(n19721), .ZN(n15766) );
  MUX2_X1 U18880 ( .A(n15766), .B(n10596), .S(n15768), .Z(P2_U3599) );
  OAI22_X1 U18881 ( .A1(n19145), .A2(n16320), .B1(n15767), .B2(n19708), .ZN(
        n15769) );
  MUX2_X1 U18882 ( .A(n15769), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15768), .Z(P2_U3596) );
  NAND2_X1 U18883 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18319) );
  AOI221_X1 U18884 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18319), .C1(n15771), 
        .C2(n18319), .A(n15770), .ZN(n18154) );
  INV_X1 U18885 ( .A(n15772), .ZN(n15773) );
  NAND2_X1 U18886 ( .A1(n18623), .A2(n18411), .ZN(n18344) );
  OAI211_X1 U18887 ( .C1(n15774), .C2(n15773), .A(n18151), .B(n18344), .ZN(
        n18152) );
  AOI22_X1 U18888 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18154), .B1(
        n18152), .B2(n18156), .ZN(P3_U2865) );
  NAND2_X1 U18889 ( .A1(n18601), .A2(n18814), .ZN(n15778) );
  NAND3_X1 U18890 ( .A1(n18601), .A2(n15776), .A3(n18814), .ZN(n15878) );
  OAI211_X1 U18891 ( .C1(n15778), .C2(n17348), .A(n15777), .B(n15878), .ZN(
        n15779) );
  NAND2_X1 U18892 ( .A1(n18808), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18160) );
  NAND2_X1 U18893 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18664), .ZN(n15781) );
  INV_X1 U18894 ( .A(n18766), .ZN(n18821) );
  AOI21_X1 U18895 ( .B1(n15782), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15784) );
  NOR2_X1 U18896 ( .A1(n15784), .A2(n15783), .ZN(n18599) );
  NAND3_X1 U18897 ( .A1(n18782), .A2(n18821), .A3(n18599), .ZN(n15785) );
  OAI21_X1 U18898 ( .B1(n18782), .B2(n16821), .A(n15785), .ZN(P3_U3284) );
  INV_X1 U18899 ( .A(n15786), .ZN(n17824) );
  INV_X1 U18900 ( .A(n17826), .ZN(n17462) );
  NAND2_X1 U18901 ( .A1(n15787), .A2(n17462), .ZN(n16374) );
  OAI21_X1 U18902 ( .B1(n17996), .B2(n16374), .A(n15788), .ZN(n15789) );
  AOI21_X1 U18903 ( .B1(n18142), .B2(n16377), .A(n15789), .ZN(n15852) );
  AOI21_X1 U18904 ( .B1(n18028), .B2(n17818), .A(n15790), .ZN(n16376) );
  OAI22_X1 U18905 ( .A1(n17996), .A2(n16358), .B1(n18125), .B2(n16362), .ZN(
        n15791) );
  INV_X1 U18906 ( .A(n15791), .ZN(n15855) );
  OAI21_X1 U18907 ( .B1(n9846), .B2(n16376), .A(n15855), .ZN(n15792) );
  AOI21_X1 U18908 ( .B1(n15793), .B2(n17463), .A(n15792), .ZN(n15798) );
  NAND2_X1 U18909 ( .A1(n15795), .A2(n15794), .ZN(n15796) );
  XOR2_X1 U18910 ( .A(n15796), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(
        n16361) );
  AOI22_X1 U18911 ( .A1(n9846), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n18057), 
        .B2(n16361), .ZN(n15797) );
  OAI221_X1 U18912 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15852), 
        .C1(n16359), .C2(n15798), .A(n15797), .ZN(P3_U2833) );
  AOI22_X1 U18913 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18931), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18940), .ZN(n15810) );
  OAI22_X1 U18914 ( .A1(n15800), .A2(n18936), .B1(n18954), .B2(n15799), .ZN(
        n15801) );
  INV_X1 U18915 ( .A(n15801), .ZN(n15809) );
  AOI22_X1 U18916 ( .A1(n15803), .A2(n18902), .B1(n15802), .B2(n18901), .ZN(
        n15808) );
  OAI211_X1 U18917 ( .C1(n15806), .C2(n15805), .A(n18949), .B(n15804), .ZN(
        n15807) );
  NAND4_X1 U18918 ( .A1(n15810), .A2(n15809), .A3(n15808), .A4(n15807), .ZN(
        P2_U2833) );
  INV_X1 U18919 ( .A(n15811), .ZN(n15812) );
  OAI211_X1 U18920 ( .C1(n11226), .C2(n15813), .A(n15812), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n15816) );
  OAI211_X1 U18921 ( .C1(n15816), .C2(n20493), .A(n15815), .B(n15814), .ZN(
        n15818) );
  NAND2_X1 U18922 ( .A1(n15816), .A2(n20493), .ZN(n15817) );
  NAND2_X1 U18923 ( .A1(n15818), .A2(n15817), .ZN(n15819) );
  AOI222_X1 U18924 ( .A1(n15820), .A2(n15819), .B1(n15820), .B2(n20274), .C1(
        n15819), .C2(n20274), .ZN(n15822) );
  INV_X1 U18925 ( .A(n15822), .ZN(n15824) );
  AOI21_X1 U18926 ( .B1(n15822), .B2(n15821), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n15823) );
  AOI21_X1 U18927 ( .B1(n15825), .B2(n15824), .A(n15823), .ZN(n15834) );
  NOR2_X1 U18928 ( .A1(P1_MORE_REG_SCAN_IN), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(
        n15828) );
  OAI211_X1 U18929 ( .C1(n15829), .C2(n15828), .A(n15827), .B(n15826), .ZN(
        n15830) );
  NOR2_X1 U18930 ( .A1(n15831), .A2(n15830), .ZN(n15833) );
  OAI211_X1 U18931 ( .C1(n15834), .C2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n15833), .B(n15832), .ZN(n15842) );
  INV_X1 U18932 ( .A(n15835), .ZN(n15839) );
  OAI21_X1 U18933 ( .B1(n20669), .B2(n15837), .A(n15836), .ZN(n15838) );
  OAI21_X1 U18934 ( .B1(n15840), .B2(n15839), .A(n15838), .ZN(n16167) );
  AOI221_X1 U18935 ( .B1(n20556), .B2(n20555), .C1(n15842), .C2(n20555), .A(
        n16167), .ZN(n16169) );
  AOI21_X1 U18936 ( .B1(n15843), .B2(n15842), .A(n15841), .ZN(n15844) );
  OAI211_X1 U18937 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20669), .A(n15844), 
        .B(n16164), .ZN(n15845) );
  NOR2_X1 U18938 ( .A1(n16169), .A2(n15845), .ZN(n15849) );
  NAND2_X1 U18939 ( .A1(n20671), .A2(n15846), .ZN(n15847) );
  NAND2_X1 U18940 ( .A1(n20556), .A2(n15847), .ZN(n15848) );
  OAI22_X1 U18941 ( .A1(n15849), .A2(n20556), .B1(n16169), .B2(n15848), .ZN(
        P1_U3161) );
  INV_X1 U18942 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16343) );
  INV_X1 U18943 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18742) );
  NOR2_X1 U18944 ( .A1(n18094), .A2(n18742), .ZN(n16348) );
  NOR3_X1 U18945 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15852), .A3(
        n16359), .ZN(n15853) );
  OAI221_X1 U18946 ( .B1(n16343), .B2(n15856), .C1(n16343), .C2(n15855), .A(
        n15854), .ZN(P3_U2832) );
  INV_X1 U18947 ( .A(HOLD), .ZN(n20561) );
  INV_X1 U18948 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20575) );
  NAND2_X1 U18949 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n15857) );
  OAI21_X1 U18950 ( .B1(n20561), .B2(n11362), .A(n15857), .ZN(n15858) );
  OAI21_X1 U18951 ( .B1(n20561), .B2(n20575), .A(n15858), .ZN(n15860) );
  OAI211_X1 U18952 ( .C1(n20669), .C2(n11362), .A(n15860), .B(n15859), .ZN(
        P1_U3195) );
  AND2_X1 U18953 ( .A1(n19929), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  INV_X1 U18954 ( .A(n15861), .ZN(n15863) );
  AOI21_X1 U18955 ( .B1(n15864), .B2(n15863), .A(n15862), .ZN(n15865) );
  INV_X1 U18956 ( .A(n15865), .ZN(n15866) );
  AOI22_X1 U18957 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15866), .B1(
        n20014), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n15871) );
  AOI22_X1 U18958 ( .A1(n15869), .A2(n20004), .B1(n15868), .B2(n15867), .ZN(
        n15870) );
  OAI211_X1 U18959 ( .C1(n20017), .C2(n15914), .A(n15871), .B(n15870), .ZN(
        P1_U3011) );
  NOR3_X1 U18960 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19762), .A3(n19756), 
        .ZN(n16317) );
  INV_X1 U18961 ( .A(n15874), .ZN(n16318) );
  NOR4_X1 U18962 ( .A1(n15873), .A2(n15872), .A3(n16317), .A4(n16318), .ZN(
        P2_U3178) );
  OAI221_X1 U18963 ( .B1(n18835), .B2(n15874), .C1(n16319), .C2(n15874), .A(
        n19523), .ZN(n19743) );
  NOR2_X1 U18964 ( .A1(n15875), .A2(n19743), .ZN(P2_U3047) );
  AOI21_X2 U18965 ( .B1(n15878), .B2(n10071), .A(n18658), .ZN(n17196) );
  NAND2_X1 U18966 ( .A1(n17120), .A2(n17196), .ZN(n17342) );
  INV_X1 U18967 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17432) );
  AOI22_X1 U18968 ( .A1(n17341), .A2(BUF2_REG_0__SCAN_IN), .B1(n17340), .B2(
        n15880), .ZN(n15881) );
  OAI221_X1 U18969 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17342), .C1(n17432), 
        .C2(n17196), .A(n15881), .ZN(P3_U2735) );
  AOI22_X1 U18970 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19876), .B1(
        n15882), .B2(n19852), .ZN(n15886) );
  INV_X1 U18971 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n15884) );
  NAND3_X1 U18972 ( .A1(n19812), .A2(n15884), .A3(n15883), .ZN(n15885) );
  OAI211_X1 U18973 ( .C1(n19821), .C2(n15887), .A(n15886), .B(n15885), .ZN(
        n15888) );
  AOI21_X1 U18974 ( .B1(n15889), .B2(n19857), .A(n15888), .ZN(n15892) );
  NOR2_X1 U18975 ( .A1(n19835), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15894) );
  INV_X1 U18976 ( .A(n15890), .ZN(n15895) );
  OAI21_X1 U18977 ( .B1(n19835), .B2(n15895), .A(n19831), .ZN(n15906) );
  OAI21_X1 U18978 ( .B1(n15894), .B2(n15906), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n15891) );
  OAI211_X1 U18979 ( .C1(n15893), .C2(n19862), .A(n15892), .B(n15891), .ZN(
        P1_U2818) );
  INV_X1 U18980 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15897) );
  AOI22_X1 U18981 ( .A1(P1_EBX_REG_21__SCAN_IN), .A2(n19875), .B1(n15895), 
        .B2(n15894), .ZN(n15896) );
  OAI21_X1 U18982 ( .B1(n15897), .B2(n19867), .A(n15896), .ZN(n15898) );
  AOI21_X1 U18983 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n15906), .A(n15898), 
        .ZN(n15900) );
  AOI22_X1 U18984 ( .A1(n15998), .A2(n19857), .B1(n15987), .B2(n19884), .ZN(
        n15899) );
  OAI211_X1 U18985 ( .C1(n15901), .C2(n19892), .A(n15900), .B(n15899), .ZN(
        P1_U2819) );
  OAI22_X1 U18986 ( .A1(n15903), .A2(n19867), .B1(n15902), .B2(n19821), .ZN(
        n15911) );
  AOI21_X1 U18987 ( .B1(n15905), .B2(n15943), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n15908) );
  INV_X1 U18988 ( .A(n15906), .ZN(n15907) );
  OAI22_X1 U18989 ( .A1(n15909), .A2(n15982), .B1(n15908), .B2(n15907), .ZN(
        n15910) );
  AOI211_X1 U18990 ( .C1(n15912), .C2(n19852), .A(n15911), .B(n15910), .ZN(
        n15913) );
  OAI21_X1 U18991 ( .B1(n19862), .B2(n15914), .A(n15913), .ZN(P1_U2820) );
  OAI22_X1 U18992 ( .A1(n15915), .A2(n19892), .B1(n15992), .B2(n19821), .ZN(
        n15916) );
  AOI211_X1 U18993 ( .C1(n19876), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n19879), .B(n15916), .ZN(n15924) );
  AOI22_X1 U18994 ( .A1(n10076), .A2(n19857), .B1(n15990), .B2(n19884), .ZN(
        n15923) );
  NAND4_X1 U18995 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .A4(n15943), .ZN(n15920) );
  NOR2_X1 U18996 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15920), .ZN(n15928) );
  OAI21_X1 U18997 ( .B1(n19835), .B2(n15917), .A(n19831), .ZN(n15942) );
  AOI21_X1 U18998 ( .B1(n15918), .B2(n19833), .A(n15942), .ZN(n15919) );
  INV_X1 U18999 ( .A(n15919), .ZN(n15937) );
  OAI21_X1 U19000 ( .B1(n15928), .B2(n15937), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15922) );
  OR3_X1 U19001 ( .A1(n20599), .A2(n15920), .A3(P1_REIP_REG_19__SCAN_IN), .ZN(
        n15921) );
  NAND4_X1 U19002 ( .A1(n15924), .A2(n15923), .A3(n15922), .A4(n15921), .ZN(
        P1_U2821) );
  AOI22_X1 U19003 ( .A1(P1_EBX_REG_18__SCAN_IN), .A2(n19875), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n15937), .ZN(n15925) );
  OAI211_X1 U19004 ( .C1(n19867), .C2(n15926), .A(n15925), .B(n19864), .ZN(
        n15927) );
  AOI211_X1 U19005 ( .C1(n19852), .C2(n15929), .A(n15928), .B(n15927), .ZN(
        n15932) );
  INV_X1 U19006 ( .A(n15930), .ZN(n16005) );
  NAND2_X1 U19007 ( .A1(n16005), .A2(n19857), .ZN(n15931) );
  OAI211_X1 U19008 ( .C1(n16060), .C2(n19862), .A(n15932), .B(n15931), .ZN(
        P1_U2822) );
  OAI22_X1 U19009 ( .A1(n15933), .A2(n19867), .B1(n15995), .B2(n19821), .ZN(
        n15934) );
  AOI211_X1 U19010 ( .C1(n19852), .C2(n16016), .A(n19879), .B(n15934), .ZN(
        n15941) );
  OAI21_X1 U19011 ( .B1(n14491), .B2(n15935), .A(n14485), .ZN(n15936) );
  INV_X1 U19012 ( .A(n15936), .ZN(n16017) );
  AOI22_X1 U19013 ( .A1(n16017), .A2(n19857), .B1(n19884), .B2(n15993), .ZN(
        n15940) );
  AND3_X1 U19014 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .A3(n15943), .ZN(n15938) );
  OAI21_X1 U19015 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n15938), .A(n15937), 
        .ZN(n15939) );
  NAND3_X1 U19016 ( .A1(n15941), .A2(n15940), .A3(n15939), .ZN(P1_U2823) );
  INV_X1 U19017 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20597) );
  INV_X1 U19018 ( .A(n15942), .ZN(n15967) );
  NAND2_X1 U19019 ( .A1(n15943), .A2(n20594), .ZN(n15955) );
  AOI21_X1 U19020 ( .B1(n19876), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n19879), .ZN(n15945) );
  NAND3_X1 U19021 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n15943), .A3(n20597), 
        .ZN(n15944) );
  OAI211_X1 U19022 ( .C1(n19821), .C2(n15946), .A(n15945), .B(n15944), .ZN(
        n15949) );
  OAI22_X1 U19023 ( .A1(n15947), .A2(n15982), .B1(n19862), .B2(n16072), .ZN(
        n15948) );
  AOI211_X1 U19024 ( .C1(n15950), .C2(n19852), .A(n15949), .B(n15948), .ZN(
        n15951) );
  OAI221_X1 U19025 ( .B1(n20597), .B2(n15967), .C1(n20597), .C2(n15955), .A(
        n15951), .ZN(P1_U2824) );
  AOI22_X1 U19026 ( .A1(n16021), .A2(n19852), .B1(n19884), .B2(n15952), .ZN(
        n15957) );
  AOI22_X1 U19027 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n19876), .B1(
        P1_EBX_REG_15__SCAN_IN), .B2(n19875), .ZN(n15953) );
  OAI211_X1 U19028 ( .C1(n15967), .C2(n20594), .A(n19864), .B(n15953), .ZN(
        n15954) );
  AOI21_X1 U19029 ( .B1(n16022), .B2(n19857), .A(n15954), .ZN(n15956) );
  NAND3_X1 U19030 ( .A1(n15957), .A2(n15956), .A3(n15955), .ZN(P1_U2825) );
  AOI21_X1 U19031 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n15958), .A(
        P1_REIP_REG_14__SCAN_IN), .ZN(n15968) );
  INV_X1 U19032 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15960) );
  OAI22_X1 U19033 ( .A1(n15960), .A2(n19867), .B1(n15959), .B2(n19821), .ZN(
        n15961) );
  AOI211_X1 U19034 ( .C1(n16078), .C2(n19884), .A(n19879), .B(n15961), .ZN(
        n15966) );
  INV_X1 U19035 ( .A(n15962), .ZN(n15963) );
  AOI22_X1 U19036 ( .A1(n15964), .A2(n19857), .B1(n15963), .B2(n19852), .ZN(
        n15965) );
  OAI211_X1 U19037 ( .C1(n15968), .C2(n15967), .A(n15966), .B(n15965), .ZN(
        P1_U2826) );
  OAI22_X1 U19038 ( .A1(n15969), .A2(n19821), .B1(n19862), .B2(n16104), .ZN(
        n15970) );
  AOI211_X1 U19039 ( .C1(n19876), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n19879), .B(n15970), .ZN(n15975) );
  INV_X1 U19040 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20588) );
  INV_X1 U19041 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15971) );
  OAI21_X1 U19042 ( .B1(n20588), .B2(n15986), .A(n15971), .ZN(n15972) );
  AOI22_X1 U19043 ( .A1(n16031), .A2(n19852), .B1(n15973), .B2(n15972), .ZN(
        n15974) );
  OAI211_X1 U19044 ( .C1(n15982), .C2(n15976), .A(n15975), .B(n15974), .ZN(
        P1_U2828) );
  INV_X1 U19045 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15980) );
  INV_X1 U19046 ( .A(n15977), .ZN(n15978) );
  AOI22_X1 U19047 ( .A1(n19884), .A2(n16105), .B1(P1_REIP_REG_11__SCAN_IN), 
        .B2(n15978), .ZN(n15979) );
  OAI211_X1 U19048 ( .C1(n19867), .C2(n15980), .A(n15979), .B(n19864), .ZN(
        n15984) );
  OAI22_X1 U19049 ( .A1(n16042), .A2(n19892), .B1(n15982), .B2(n15981), .ZN(
        n15983) );
  AOI211_X1 U19050 ( .C1(P1_EBX_REG_11__SCAN_IN), .C2(n19875), .A(n15984), .B(
        n15983), .ZN(n15985) );
  OAI21_X1 U19051 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15986), .A(n15985), 
        .ZN(P1_U2829) );
  AOI22_X1 U19052 ( .A1(n15998), .A2(n19895), .B1(n15987), .B2(n19894), .ZN(
        n15988) );
  OAI21_X1 U19053 ( .B1(n19899), .B2(n15989), .A(n15988), .ZN(P1_U2851) );
  AOI22_X1 U19054 ( .A1(n10076), .A2(n19895), .B1(n15990), .B2(n19894), .ZN(
        n15991) );
  OAI21_X1 U19055 ( .B1(n19899), .B2(n15992), .A(n15991), .ZN(P1_U2853) );
  AOI22_X1 U19056 ( .A1(n16017), .A2(n19895), .B1(n19894), .B2(n15993), .ZN(
        n15994) );
  OAI21_X1 U19057 ( .B1(n19899), .B2(n15995), .A(n15994), .ZN(P1_U2855) );
  INV_X1 U19058 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16403) );
  AOI22_X1 U19059 ( .A1(n16010), .A2(n15996), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n16008), .ZN(n16000) );
  INV_X1 U19060 ( .A(n15997), .ZN(n16012) );
  AOI22_X1 U19061 ( .A1(n15998), .A2(n16012), .B1(n16011), .B2(DATAI_21_), 
        .ZN(n15999) );
  OAI211_X1 U19062 ( .C1(n16015), .C2(n16403), .A(n16000), .B(n15999), .ZN(
        P1_U2883) );
  INV_X1 U19063 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16406) );
  AOI22_X1 U19064 ( .A1(n16010), .A2(n16001), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n16008), .ZN(n16003) );
  AOI22_X1 U19065 ( .A1(n10076), .A2(n16012), .B1(n16011), .B2(DATAI_19_), 
        .ZN(n16002) );
  OAI211_X1 U19066 ( .C1(n16015), .C2(n16406), .A(n16003), .B(n16002), .ZN(
        P1_U2885) );
  INV_X1 U19067 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16408) );
  AOI22_X1 U19068 ( .A1(n16010), .A2(n16004), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n16008), .ZN(n16007) );
  AOI22_X1 U19069 ( .A1(n16005), .A2(n16012), .B1(n16011), .B2(DATAI_18_), 
        .ZN(n16006) );
  OAI211_X1 U19070 ( .C1(n16015), .C2(n16408), .A(n16007), .B(n16006), .ZN(
        P1_U2886) );
  INV_X1 U19071 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16410) );
  AOI22_X1 U19072 ( .A1(n16010), .A2(n16009), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n16008), .ZN(n16014) );
  AOI22_X1 U19073 ( .A1(n16017), .A2(n16012), .B1(n16011), .B2(DATAI_17_), 
        .ZN(n16013) );
  OAI211_X1 U19074 ( .C1(n16015), .C2(n16410), .A(n16014), .B(n16013), .ZN(
        P1_U2887) );
  AOI22_X1 U19075 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n20014), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16019) );
  AOI22_X1 U19076 ( .A1(n16017), .A2(n14671), .B1(n16016), .B2(n16032), .ZN(
        n16018) );
  OAI211_X1 U19077 ( .C1(n16035), .C2(n16020), .A(n16019), .B(n16018), .ZN(
        P1_U2982) );
  AOI22_X1 U19078 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20014), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16024) );
  AOI22_X1 U19079 ( .A1(n16022), .A2(n14671), .B1(n16021), .B2(n16032), .ZN(
        n16023) );
  OAI211_X1 U19080 ( .C1(n16025), .C2(n16035), .A(n16024), .B(n16023), .ZN(
        P1_U2984) );
  OAI21_X1 U19081 ( .B1(n16028), .B2(n16027), .A(n16026), .ZN(n16029) );
  INV_X1 U19082 ( .A(n16029), .ZN(n16099) );
  AOI22_X1 U19083 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20014), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16034) );
  AOI22_X1 U19084 ( .A1(n16032), .A2(n16031), .B1(n14671), .B2(n16030), .ZN(
        n16033) );
  OAI211_X1 U19085 ( .C1(n16099), .C2(n16035), .A(n16034), .B(n16033), .ZN(
        P1_U2987) );
  AOI22_X1 U19086 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20014), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16041) );
  NOR2_X1 U19087 ( .A1(n14729), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16037) );
  NOR2_X1 U19088 ( .A1(n14704), .A2(n16114), .ZN(n16036) );
  MUX2_X1 U19089 ( .A(n16037), .B(n16036), .S(n14844), .Z(n16038) );
  XOR2_X1 U19090 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n16038), .Z(
        n16107) );
  AOI22_X1 U19091 ( .A1(n19968), .A2(n16107), .B1(n14671), .B2(n16039), .ZN(
        n16040) );
  OAI211_X1 U19092 ( .C1(n19972), .C2(n16042), .A(n16041), .B(n16040), .ZN(
        P1_U2988) );
  AOI22_X1 U19093 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20014), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16048) );
  NAND2_X1 U19094 ( .A1(n16045), .A2(n16044), .ZN(n16046) );
  XNOR2_X1 U19095 ( .A(n16043), .B(n16046), .ZN(n16141) );
  AOI22_X1 U19096 ( .A1(n16141), .A2(n19968), .B1(n14671), .B2(n19896), .ZN(
        n16047) );
  OAI211_X1 U19097 ( .C1(n19972), .C2(n19839), .A(n16048), .B(n16047), .ZN(
        P1_U2992) );
  AOI22_X1 U19098 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20014), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16053) );
  XNOR2_X1 U19099 ( .A(n16050), .B(n16149), .ZN(n16051) );
  XNOR2_X1 U19100 ( .A(n16049), .B(n16051), .ZN(n16146) );
  AOI22_X1 U19101 ( .A1(n16146), .A2(n19968), .B1(n14671), .B2(n19858), .ZN(
        n16052) );
  OAI211_X1 U19102 ( .C1(n19972), .C2(n19850), .A(n16053), .B(n16052), .ZN(
        P1_U2993) );
  AOI22_X1 U19103 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20014), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16059) );
  OAI21_X1 U19104 ( .B1(n16056), .B2(n16055), .A(n16054), .ZN(n16057) );
  INV_X1 U19105 ( .A(n16057), .ZN(n16152) );
  AOI22_X1 U19106 ( .A1(n16152), .A2(n19968), .B1(n14671), .B2(n19871), .ZN(
        n16058) );
  OAI211_X1 U19107 ( .C1(n19972), .C2(n19874), .A(n16059), .B(n16058), .ZN(
        P1_U2994) );
  OAI22_X1 U19108 ( .A1(n16061), .A2(n16126), .B1(n20017), .B2(n16060), .ZN(
        n16062) );
  AOI21_X1 U19109 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n16063), .A(
        n16062), .ZN(n16067) );
  NAND3_X1 U19110 ( .A1(n16065), .A2(n16068), .A3(n16064), .ZN(n16066) );
  OAI211_X1 U19111 ( .C1(n20599), .C2(n16122), .A(n16067), .B(n16066), .ZN(
        P1_U3013) );
  OAI21_X1 U19112 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n16068), .ZN(n16071) );
  OAI222_X1 U19113 ( .A1(n16072), .A2(n20017), .B1(n16071), .B2(n16070), .C1(
        n16126), .C2(n16069), .ZN(n16073) );
  INV_X1 U19114 ( .A(n16073), .ZN(n16075) );
  NAND2_X1 U19115 ( .A1(n20014), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n16074) );
  OAI211_X1 U19116 ( .C1(n16077), .C2(n16076), .A(n16075), .B(n16074), .ZN(
        P1_U3015) );
  AOI22_X1 U19117 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16087), .B1(
        n20014), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16085) );
  AOI22_X1 U19118 ( .A1(n16079), .A2(n20004), .B1(n19981), .B2(n16078), .ZN(
        n16084) );
  AOI21_X1 U19119 ( .B1(n19993), .B2(n19988), .A(n19994), .ZN(n16080) );
  INV_X1 U19120 ( .A(n16080), .ZN(n16123) );
  NAND3_X1 U19121 ( .A1(n16082), .A2(n16081), .A3(n16123), .ZN(n16083) );
  NAND3_X1 U19122 ( .A1(n16085), .A2(n16084), .A3(n16083), .ZN(P1_U3017) );
  AOI22_X1 U19123 ( .A1(n20014), .A2(P1_REIP_REG_13__SCAN_IN), .B1(n19981), 
        .B2(n16086), .ZN(n16090) );
  AOI22_X1 U19124 ( .A1(n16088), .A2(n20004), .B1(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16087), .ZN(n16089) );
  OAI211_X1 U19125 ( .C1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n16091), .A(
        n16090), .B(n16089), .ZN(P1_U3018) );
  INV_X1 U19126 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16110) );
  NOR2_X1 U19127 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16110), .ZN(
        n16101) );
  NAND2_X1 U19128 ( .A1(n16094), .A2(n16123), .ZN(n19987) );
  NOR2_X1 U19129 ( .A1(n16092), .A2(n19987), .ZN(n16106) );
  INV_X1 U19130 ( .A(n16093), .ZN(n19990) );
  OR2_X1 U19131 ( .A1(n16095), .A2(n16094), .ZN(n19992) );
  OAI211_X1 U19132 ( .C1(n19990), .C2(n19993), .A(n19992), .B(n19989), .ZN(
        n19983) );
  AOI21_X1 U19133 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16096), .A(
        n20008), .ZN(n16097) );
  NOR2_X1 U19134 ( .A1(n19983), .A2(n16097), .ZN(n16111) );
  OAI22_X1 U19135 ( .A1(n16099), .A2(n16126), .B1(n16111), .B2(n16098), .ZN(
        n16100) );
  AOI21_X1 U19136 ( .B1(n16101), .B2(n16106), .A(n16100), .ZN(n16103) );
  NAND2_X1 U19137 ( .A1(n20014), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n16102) );
  OAI211_X1 U19138 ( .C1(n20017), .C2(n16104), .A(n16103), .B(n16102), .ZN(
        P1_U3019) );
  AOI22_X1 U19139 ( .A1(n20014), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n19981), 
        .B2(n16105), .ZN(n16109) );
  AOI22_X1 U19140 ( .A1(n16107), .A2(n20004), .B1(n16110), .B2(n16106), .ZN(
        n16108) );
  OAI211_X1 U19141 ( .C1(n16111), .C2(n16110), .A(n16109), .B(n16108), .ZN(
        P1_U3020) );
  OAI211_X1 U19142 ( .C1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n16124), .B(n16123), .ZN(n16115) );
  OAI21_X1 U19143 ( .B1(n16113), .B2(n19983), .A(n16112), .ZN(n16131) );
  OAI22_X1 U19144 ( .A1(n16116), .A2(n16115), .B1(n16114), .B2(n16131), .ZN(
        n16117) );
  AOI21_X1 U19145 ( .B1(n16118), .B2(n20004), .A(n16117), .ZN(n16120) );
  NAND2_X1 U19146 ( .A1(n20014), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n16119) );
  OAI211_X1 U19147 ( .C1(n20017), .C2(n16121), .A(n16120), .B(n16119), .ZN(
        P1_U3021) );
  NOR2_X1 U19148 ( .A1(n16122), .A2(n20586), .ZN(n16129) );
  NAND2_X1 U19149 ( .A1(n16124), .A2(n16123), .ZN(n16125) );
  OAI22_X1 U19150 ( .A1(n16127), .A2(n16126), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16125), .ZN(n16128) );
  AOI211_X1 U19151 ( .C1(n19981), .C2(n19807), .A(n16129), .B(n16128), .ZN(
        n16130) );
  OAI21_X1 U19152 ( .B1(n14150), .B2(n16131), .A(n16130), .ZN(P1_U3022) );
  INV_X1 U19153 ( .A(n19987), .ZN(n19976) );
  NAND3_X1 U19154 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16145), .A3(
        n19976), .ZN(n16144) );
  AOI22_X1 U19155 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n16132), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n12954), .ZN(n16138) );
  AOI22_X1 U19156 ( .A1(n20014), .A2(P1_REIP_REG_8__SCAN_IN), .B1(n19981), 
        .B2(n19819), .ZN(n16137) );
  AOI21_X1 U19157 ( .B1(n16134), .B2(n16133), .A(n19983), .ZN(n16156) );
  OAI21_X1 U19158 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n20008), .A(
        n16156), .ZN(n16140) );
  AOI22_X1 U19159 ( .A1(n16135), .A2(n20004), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n16140), .ZN(n16136) );
  OAI211_X1 U19160 ( .C1(n16144), .C2(n16138), .A(n16137), .B(n16136), .ZN(
        P1_U3023) );
  AOI21_X1 U19161 ( .B1(n9734), .B2(n9920), .A(n14016), .ZN(n19893) );
  AOI22_X1 U19162 ( .A1(n20014), .A2(P1_REIP_REG_7__SCAN_IN), .B1(n19981), 
        .B2(n19893), .ZN(n16143) );
  AOI22_X1 U19163 ( .A1(n16141), .A2(n20004), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16140), .ZN(n16142) );
  OAI211_X1 U19164 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n16144), .A(
        n16143), .B(n16142), .ZN(P1_U3024) );
  NAND2_X1 U19165 ( .A1(n16145), .A2(n19976), .ZN(n16150) );
  AOI222_X1 U19166 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20014), .B1(n19981), 
        .B2(n16147), .C1(n20004), .C2(n16146), .ZN(n16148) );
  OAI221_X1 U19167 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16150), .C1(
        n16149), .C2(n16156), .A(n16148), .ZN(P1_U3025) );
  AOI22_X1 U19168 ( .A1(n20014), .A2(P1_REIP_REG_5__SCAN_IN), .B1(n19981), 
        .B2(n19863), .ZN(n16154) );
  NOR3_X1 U19169 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n19975), .A3(
        n19987), .ZN(n16151) );
  AOI21_X1 U19170 ( .B1(n16152), .B2(n20004), .A(n16151), .ZN(n16153) );
  OAI211_X1 U19171 ( .C1(n16156), .C2(n16155), .A(n16154), .B(n16153), .ZN(
        P1_U3026) );
  OR3_X1 U19172 ( .A1(n19887), .A2(n20635), .A3(n12048), .ZN(n16159) );
  OAI22_X1 U19173 ( .A1(n16160), .A2(n16159), .B1(n16158), .B2(n16157), .ZN(
        P1_U3468) );
  NAND4_X1 U19174 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n12008), .A4(n20669), .ZN(n16161) );
  NAND2_X1 U19175 ( .A1(n16162), .A2(n16161), .ZN(n20557) );
  OAI21_X1 U19176 ( .B1(n16169), .B2(n20556), .A(n20555), .ZN(n16163) );
  OAI211_X1 U19177 ( .C1(n16165), .C2(n20669), .A(n16164), .B(n16163), .ZN(
        n16166) );
  AOI221_X1 U19178 ( .B1(n16168), .B2(n16167), .C1(n20557), .C2(n16167), .A(
        n16166), .ZN(P1_U3162) );
  NOR2_X1 U19179 ( .A1(n16169), .A2(n20556), .ZN(n16171) );
  OAI22_X1 U19180 ( .A1(n20389), .A2(n16171), .B1(n16170), .B2(n20556), .ZN(
        P1_U3466) );
  AOI22_X1 U19181 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n16172), .B1(
        P2_REIP_REG_31__SCAN_IN), .B2(n18940), .ZN(n16180) );
  AOI22_X1 U19182 ( .A1(n16173), .A2(n18923), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n18931), .ZN(n16179) );
  INV_X1 U19183 ( .A(n16174), .ZN(n18956) );
  AOI22_X1 U19184 ( .A1(n16175), .A2(n18902), .B1(n18901), .B2(n18956), .ZN(
        n16178) );
  NAND2_X1 U19185 ( .A1(n18893), .A2(n16176), .ZN(n16183) );
  NAND4_X1 U19186 ( .A1(n18949), .A2(n16184), .A3(n18893), .A4(n16183), .ZN(
        n16177) );
  NAND4_X1 U19187 ( .A1(n16180), .A2(n16179), .A3(n16178), .A4(n16177), .ZN(
        P2_U2824) );
  AOI22_X1 U19188 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n18931), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n18940), .ZN(n16192) );
  AOI22_X1 U19189 ( .A1(n16181), .A2(n18923), .B1(P2_EBX_REG_30__SCAN_IN), 
        .B2(n18922), .ZN(n16191) );
  INV_X1 U19190 ( .A(n15235), .ZN(n16182) );
  AOI22_X1 U19191 ( .A1(n16182), .A2(n18902), .B1(n18901), .B2(n15487), .ZN(
        n16190) );
  AOI21_X1 U19192 ( .B1(n16184), .B2(n16183), .A(n19628), .ZN(n16188) );
  INV_X1 U19193 ( .A(n16183), .ZN(n16186) );
  NAND2_X1 U19194 ( .A1(n16188), .A2(n16187), .ZN(n16189) );
  NAND4_X1 U19195 ( .A1(n16192), .A2(n16191), .A3(n16190), .A4(n16189), .ZN(
        P2_U2825) );
  AOI22_X1 U19196 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18931), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n18940), .ZN(n16203) );
  AOI22_X1 U19197 ( .A1(n16193), .A2(n18923), .B1(P2_EBX_REG_28__SCAN_IN), 
        .B2(n18922), .ZN(n16202) );
  OAI22_X1 U19198 ( .A1(n16195), .A2(n18946), .B1(n16194), .B2(n18947), .ZN(
        n16196) );
  INV_X1 U19199 ( .A(n16196), .ZN(n16201) );
  OAI211_X1 U19200 ( .C1(n16199), .C2(n16198), .A(n18949), .B(n16197), .ZN(
        n16200) );
  NAND4_X1 U19201 ( .A1(n16203), .A2(n16202), .A3(n16201), .A4(n16200), .ZN(
        P2_U2827) );
  AOI22_X1 U19202 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18931), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n18940), .ZN(n16216) );
  OAI22_X1 U19203 ( .A1(n16205), .A2(n18936), .B1(n18954), .B2(n16204), .ZN(
        n16206) );
  INV_X1 U19204 ( .A(n16206), .ZN(n16215) );
  INV_X1 U19205 ( .A(n16207), .ZN(n16208) );
  AOI22_X1 U19206 ( .A1(n16209), .A2(n18902), .B1(n16208), .B2(n18901), .ZN(
        n16214) );
  OAI211_X1 U19207 ( .C1(n16212), .C2(n16211), .A(n18949), .B(n16210), .ZN(
        n16213) );
  NAND4_X1 U19208 ( .A1(n16216), .A2(n16215), .A3(n16214), .A4(n16213), .ZN(
        P2_U2829) );
  AOI22_X1 U19209 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18931), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n18940), .ZN(n16227) );
  AOI22_X1 U19210 ( .A1(n16217), .A2(n18923), .B1(P2_EBX_REG_23__SCAN_IN), 
        .B2(n18922), .ZN(n16226) );
  INV_X1 U19211 ( .A(n16218), .ZN(n16219) );
  AOI22_X1 U19212 ( .A1(n16220), .A2(n18902), .B1(n16219), .B2(n18901), .ZN(
        n16225) );
  OAI211_X1 U19213 ( .C1(n16223), .C2(n16222), .A(n18949), .B(n16221), .ZN(
        n16224) );
  NAND4_X1 U19214 ( .A1(n16227), .A2(n16226), .A3(n16225), .A4(n16224), .ZN(
        P2_U2832) );
  AOI22_X1 U19215 ( .A1(n16235), .A2(n18978), .B1(n19015), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n16233) );
  AOI22_X1 U19216 ( .A1(n18955), .A2(BUF2_REG_24__SCAN_IN), .B1(n18957), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n16232) );
  INV_X1 U19217 ( .A(n16228), .ZN(n16230) );
  AOI22_X1 U19218 ( .A1(n16230), .A2(n19017), .B1(n19016), .B2(n16229), .ZN(
        n16231) );
  NAND3_X1 U19219 ( .A1(n16233), .A2(n16232), .A3(n16231), .ZN(P2_U2895) );
  AOI22_X1 U19220 ( .A1(n16235), .A2(n16234), .B1(n19015), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n16240) );
  AOI22_X1 U19221 ( .A1(n18955), .A2(BUF2_REG_19__SCAN_IN), .B1(n18957), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n16239) );
  AOI22_X1 U19222 ( .A1(n16237), .A2(n19017), .B1(n19016), .B2(n16236), .ZN(
        n16238) );
  NAND3_X1 U19223 ( .A1(n16240), .A2(n16239), .A3(n16238), .ZN(P2_U2900) );
  AOI22_X1 U19224 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19069), .B1(
        n19059), .B2(n16241), .ZN(n16242) );
  OAI21_X1 U19225 ( .B1(n12748), .B2(n16290), .A(n16242), .ZN(n16243) );
  INV_X1 U19226 ( .A(n16243), .ZN(n16253) );
  AOI21_X1 U19227 ( .B1(n16276), .B2(n9673), .A(n16244), .ZN(n16283) );
  NAND2_X1 U19228 ( .A1(n9686), .A2(n16245), .ZN(n16249) );
  NAND2_X1 U19229 ( .A1(n16247), .A2(n16246), .ZN(n16248) );
  XNOR2_X1 U19230 ( .A(n16249), .B(n16248), .ZN(n16280) );
  AOI22_X1 U19231 ( .A1(n16283), .A2(n16251), .B1(n16250), .B2(n16280), .ZN(
        n16252) );
  OAI211_X1 U19232 ( .C1(n16272), .C2(n16286), .A(n16253), .B(n16252), .ZN(
        P2_U3003) );
  AOI22_X1 U19233 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n13328), .B1(n19059), 
        .B2(n16254), .ZN(n16260) );
  OAI22_X1 U19234 ( .A1(n16256), .A2(n19075), .B1(n16255), .B2(n19072), .ZN(
        n16257) );
  AOI21_X1 U19235 ( .B1(n19078), .B2(n16258), .A(n16257), .ZN(n16259) );
  OAI211_X1 U19236 ( .C1(n16261), .C2(n19067), .A(n16260), .B(n16259), .ZN(
        P2_U3004) );
  OAI22_X1 U19237 ( .A1(n9906), .A2(n19067), .B1(n16262), .B2(n18921), .ZN(
        n16263) );
  AOI21_X1 U19238 ( .B1(P2_REIP_REG_9__SCAN_IN), .B2(n18939), .A(n16263), .ZN(
        n16271) );
  OAI21_X1 U19239 ( .B1(n16264), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15731), .ZN(n16295) );
  OR2_X1 U19240 ( .A1(n16267), .A2(n16266), .ZN(n16268) );
  XNOR2_X1 U19241 ( .A(n16265), .B(n16268), .ZN(n16294) );
  OAI22_X1 U19242 ( .A1(n16295), .A2(n19075), .B1(n19072), .B2(n16294), .ZN(
        n16269) );
  INV_X1 U19243 ( .A(n16269), .ZN(n16270) );
  OAI211_X1 U19244 ( .C1(n16272), .C2(n18928), .A(n16271), .B(n16270), .ZN(
        P2_U3005) );
  AOI211_X1 U19245 ( .C1(n16275), .C2(n16276), .A(n16274), .B(n16273), .ZN(
        n16279) );
  OAI22_X1 U19246 ( .A1(n16277), .A2(n16276), .B1(n16305), .B2(n18972), .ZN(
        n16278) );
  AOI211_X1 U19247 ( .C1(n18939), .C2(P2_REIP_REG_11__SCAN_IN), .A(n16279), 
        .B(n16278), .ZN(n16285) );
  AOI22_X1 U19248 ( .A1(n16283), .A2(n16282), .B1(n16281), .B2(n16280), .ZN(
        n16284) );
  OAI211_X1 U19249 ( .C1(n16315), .C2(n16286), .A(n16285), .B(n16284), .ZN(
        P2_U3035) );
  OR2_X1 U19250 ( .A1(n16288), .A2(n16287), .ZN(n16289) );
  NAND2_X1 U19251 ( .A1(n16289), .A2(n13990), .ZN(n18977) );
  OAI22_X1 U19252 ( .A1(n16305), .A2(n18977), .B1(n12742), .B2(n16290), .ZN(
        n16291) );
  AOI221_X1 U19253 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16293), .C1(
        n16292), .C2(n16293), .A(n16291), .ZN(n16298) );
  OAI22_X1 U19254 ( .A1(n16295), .A2(n16308), .B1(n16306), .B2(n16294), .ZN(
        n16296) );
  INV_X1 U19255 ( .A(n16296), .ZN(n16297) );
  OAI211_X1 U19256 ( .C1(n16315), .C2(n18928), .A(n16298), .B(n16297), .ZN(
        P2_U3037) );
  AOI221_X1 U19257 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n16300), .C2(n16303), .A(
        n16299), .ZN(n16312) );
  OAI21_X1 U19258 ( .B1(n13834), .B2(n16302), .A(n16301), .ZN(n18993) );
  OAI22_X1 U19259 ( .A1(n18993), .A2(n16305), .B1(n16304), .B2(n16303), .ZN(
        n16311) );
  OAI22_X1 U19260 ( .A1(n16309), .A2(n16308), .B1(n16307), .B2(n16306), .ZN(
        n16310) );
  NOR4_X1 U19261 ( .A1(n16313), .A2(n16312), .A3(n16311), .A4(n16310), .ZN(
        n16314) );
  OAI21_X1 U19262 ( .B1(n16315), .B2(n18945), .A(n16314), .ZN(P2_U3041) );
  AOI211_X1 U19263 ( .C1(n16319), .C2(n16318), .A(n16317), .B(n16316), .ZN(
        n16323) );
  OAI22_X1 U19264 ( .A1(n19625), .A2(n19756), .B1(n18829), .B2(n16320), .ZN(
        n16321) );
  MUX2_X1 U19265 ( .A(n16321), .B(n19625), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n16322) );
  OAI211_X1 U19266 ( .C1(n16324), .C2(n18832), .A(n16323), .B(n16322), .ZN(
        P2_U3176) );
  AOI22_X1 U19267 ( .A1(n18795), .A2(n17875), .B1(n18797), .B2(n18600), .ZN(
        n16325) );
  OAI21_X4 U19268 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18811), .A(n16494), 
        .ZN(n17811) );
  NAND2_X1 U19269 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17761) );
  INV_X1 U19270 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17730) );
  INV_X1 U19271 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17716) );
  NOR2_X1 U19272 ( .A1(n17730), .A2(n17716), .ZN(n17712) );
  NAND2_X1 U19273 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17637) );
  NOR2_X1 U19274 ( .A1(n17637), .A2(n17636), .ZN(n16694) );
  NAND2_X1 U19275 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17612) );
  NAND2_X1 U19276 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17575) );
  NOR2_X1 U19277 ( .A1(n20720), .A2(n17544), .ZN(n17538) );
  NAND2_X1 U19278 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17505) );
  NOR2_X2 U19279 ( .A1(n9670), .A2(n17505), .ZN(n17487) );
  NAND2_X1 U19280 ( .A1(n16364), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16326) );
  INV_X1 U19281 ( .A(n17471), .ZN(n17458) );
  NAND3_X1 U19282 ( .A1(n17458), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16355) );
  NOR2_X1 U19283 ( .A1(n20747), .A2(n16355), .ZN(n16327) );
  AOI21_X1 U19284 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17596), .A(
        n18545), .ZN(n17611) );
  INV_X1 U19285 ( .A(n17611), .ZN(n17661) );
  NAND2_X1 U19286 ( .A1(n16327), .A2(n17661), .ZN(n16345) );
  XNOR2_X1 U19287 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16329) );
  INV_X1 U19288 ( .A(n17596), .ZN(n17564) );
  NOR2_X1 U19289 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17564), .ZN(
        n16366) );
  INV_X1 U19290 ( .A(n16365), .ZN(n16516) );
  OAI22_X1 U19291 ( .A1(n17812), .A2(n16516), .B1(n18507), .B2(n16327), .ZN(
        n16328) );
  OR2_X1 U19292 ( .A1(n16328), .A2(n17798), .ZN(n16357) );
  NOR2_X1 U19293 ( .A1(n16366), .A2(n16357), .ZN(n16346) );
  OAI22_X1 U19294 ( .A1(n16345), .A2(n16329), .B1(n16346), .B2(n16541), .ZN(
        n16330) );
  AOI211_X1 U19295 ( .C1(n17609), .C2(n16531), .A(n16331), .B(n16330), .ZN(
        n16339) );
  INV_X1 U19296 ( .A(n16333), .ZN(n16335) );
  NOR2_X2 U19297 ( .A1(n16375), .A2(n17815), .ZN(n17724) );
  OAI211_X1 U19298 ( .C1(n17816), .C2(n16340), .A(n16339), .B(n16338), .ZN(
        P3_U2799) );
  NOR2_X2 U19299 ( .A1(n16342), .A2(n17618), .ZN(n17517) );
  NAND3_X1 U19300 ( .A1(n16344), .A2(n17517), .A3(n16343), .ZN(n16353) );
  INV_X1 U19301 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16545) );
  XNOR2_X1 U19302 ( .A(n16545), .B(n16364), .ZN(n16544) );
  AOI22_X1 U19303 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16346), .B1(
        n16345), .B2(n16545), .ZN(n16347) );
  AOI211_X1 U19304 ( .C1(n17609), .C2(n16544), .A(n16348), .B(n16347), .ZN(
        n16352) );
  OAI22_X1 U19305 ( .A1(n16362), .A2(n17816), .B1(n16358), .B2(n16334), .ZN(
        n16350) );
  AOI22_X1 U19306 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16350), .B1(
        n17723), .B2(n16349), .ZN(n16351) );
  OAI211_X1 U19307 ( .C1(n16354), .C2(n16353), .A(n16352), .B(n16351), .ZN(
        P3_U2800) );
  OAI21_X1 U19308 ( .B1(n18507), .B2(n16355), .A(n20747), .ZN(n16356) );
  AOI22_X1 U19309 ( .A1(n9846), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n16357), 
        .B2(n16356), .ZN(n16370) );
  AOI211_X1 U19310 ( .C1(n16359), .C2(n16374), .A(n16358), .B(n16334), .ZN(
        n16360) );
  AOI21_X1 U19311 ( .B1(n17723), .B2(n16361), .A(n16360), .ZN(n16369) );
  INV_X1 U19312 ( .A(n16362), .ZN(n16363) );
  OAI211_X1 U19313 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16377), .A(
        n17803), .B(n16363), .ZN(n16368) );
  AOI21_X1 U19314 ( .B1(n20747), .B2(n16365), .A(n16364), .ZN(n16553) );
  OAI21_X1 U19315 ( .B1(n16366), .B2(n17609), .A(n16553), .ZN(n16367) );
  NAND4_X1 U19316 ( .A1(n16370), .A2(n16369), .A3(n16368), .A4(n16367), .ZN(
        P3_U2801) );
  NAND2_X1 U19317 ( .A1(n18600), .A2(n17312), .ZN(n18014) );
  AOI22_X1 U19318 ( .A1(n17875), .A2(n17883), .B1(n17962), .B2(n17990), .ZN(
        n17927) );
  NAND2_X1 U19319 ( .A1(n16371), .A2(n17927), .ZN(n17896) );
  NAND2_X1 U19320 ( .A1(n17896), .A2(n17880), .ZN(n17885) );
  NOR2_X1 U19321 ( .A1(n18143), .A2(n17868), .ZN(n17856) );
  NOR2_X1 U19322 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n16372), .ZN(
        n17470) );
  AOI22_X1 U19323 ( .A1(n9846), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n17856), 
        .B2(n17470), .ZN(n16381) );
  INV_X1 U19324 ( .A(n17477), .ZN(n16373) );
  AOI21_X1 U19325 ( .B1(n17722), .B2(n16373), .A(n9676), .ZN(n17467) );
  AOI22_X1 U19326 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n10223), .B1(
        n17722), .B2(n17463), .ZN(n17466) );
  NOR2_X1 U19327 ( .A1(n17467), .A2(n17466), .ZN(n17465) );
  NAND4_X1 U19328 ( .A1(n17722), .A2(n17477), .A3(n18140), .A4(n17463), .ZN(
        n16379) );
  NAND3_X1 U19329 ( .A1(n18057), .A2(n9676), .A3(n17466), .ZN(n16378) );
  NAND4_X1 U19330 ( .A1(n16381), .A2(n16380), .A3(n16379), .A4(n16378), .ZN(
        P3_U2834) );
  NOR3_X1 U19331 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), 
        .A3(P3_BE_N_REG_0__SCAN_IN), .ZN(n16383) );
  NOR4_X1 U19332 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16382) );
  INV_X2 U19333 ( .A(n16477), .ZN(U215) );
  NAND4_X1 U19334 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16383), .A3(n16382), .A4(
        U215), .ZN(U213) );
  INV_X1 U19335 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16479) );
  INV_X2 U19336 ( .A(U214), .ZN(n16441) );
  OAI222_X1 U19337 ( .A1(U212), .A2(n16479), .B1(n16443), .B2(n16385), .C1(
        U214), .C2(n16480), .ZN(U216) );
  INV_X1 U19338 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16387) );
  AOI22_X1 U19339 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16440), .ZN(n16386) );
  OAI21_X1 U19340 ( .B1(n16387), .B2(n16443), .A(n16386), .ZN(U217) );
  INV_X1 U19341 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16389) );
  AOI22_X1 U19342 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16440), .ZN(n16388) );
  OAI21_X1 U19343 ( .B1(n16389), .B2(n16443), .A(n16388), .ZN(U218) );
  INV_X1 U19344 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16391) );
  AOI22_X1 U19345 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16440), .ZN(n16390) );
  OAI21_X1 U19346 ( .B1(n16391), .B2(n16443), .A(n16390), .ZN(U219) );
  INV_X1 U19347 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n19107) );
  AOI22_X1 U19348 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16440), .ZN(n16392) );
  OAI21_X1 U19349 ( .B1(n19107), .B2(n16443), .A(n16392), .ZN(U220) );
  INV_X1 U19350 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n20709) );
  INV_X1 U19351 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20707) );
  INV_X1 U19352 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n16393) );
  OAI222_X1 U19353 ( .A1(U212), .A2(n20709), .B1(n16443), .B2(n20707), .C1(
        U214), .C2(n16393), .ZN(U221) );
  AOI22_X1 U19354 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16440), .ZN(n16394) );
  OAI21_X1 U19355 ( .B1(n16395), .B2(n16443), .A(n16394), .ZN(U222) );
  INV_X1 U19356 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16397) );
  AOI22_X1 U19357 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16440), .ZN(n16396) );
  OAI21_X1 U19358 ( .B1(n16397), .B2(n16443), .A(n16396), .ZN(U223) );
  INV_X1 U19359 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16399) );
  AOI22_X1 U19360 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16440), .ZN(n16398) );
  OAI21_X1 U19361 ( .B1(n16399), .B2(n16443), .A(n16398), .ZN(U224) );
  INV_X1 U19362 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16401) );
  AOI22_X1 U19363 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16440), .ZN(n16400) );
  OAI21_X1 U19364 ( .B1(n16401), .B2(n16443), .A(n16400), .ZN(U225) );
  AOI22_X1 U19365 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16440), .ZN(n16402) );
  OAI21_X1 U19366 ( .B1(n16403), .B2(n16443), .A(n16402), .ZN(U226) );
  INV_X1 U19367 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n19118) );
  AOI22_X1 U19368 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16440), .ZN(n16404) );
  OAI21_X1 U19369 ( .B1(n19118), .B2(n16443), .A(n16404), .ZN(U227) );
  AOI22_X1 U19370 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16440), .ZN(n16405) );
  OAI21_X1 U19371 ( .B1(n16406), .B2(n16443), .A(n16405), .ZN(U228) );
  AOI22_X1 U19372 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16440), .ZN(n16407) );
  OAI21_X1 U19373 ( .B1(n16408), .B2(n16443), .A(n16407), .ZN(U229) );
  AOI22_X1 U19374 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16440), .ZN(n16409) );
  OAI21_X1 U19375 ( .B1(n16410), .B2(n16443), .A(n16409), .ZN(U230) );
  INV_X1 U19376 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n19094) );
  AOI22_X1 U19377 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16440), .ZN(n16411) );
  OAI21_X1 U19378 ( .B1(n19094), .B2(n16443), .A(n16411), .ZN(U231) );
  AOI22_X1 U19379 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16440), .ZN(n16412) );
  OAI21_X1 U19380 ( .B1(n13296), .B2(n16443), .A(n16412), .ZN(U232) );
  AOI22_X1 U19381 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16440), .ZN(n16413) );
  OAI21_X1 U19382 ( .B1(n12672), .B2(n16443), .A(n16413), .ZN(U233) );
  INV_X1 U19383 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16415) );
  AOI22_X1 U19384 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16440), .ZN(n16414) );
  OAI21_X1 U19385 ( .B1(n16415), .B2(n16443), .A(n16414), .ZN(U234) );
  INV_X1 U19386 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16417) );
  AOI22_X1 U19387 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16440), .ZN(n16416) );
  OAI21_X1 U19388 ( .B1(n16417), .B2(n16443), .A(n16416), .ZN(U235) );
  INV_X1 U19389 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16419) );
  AOI22_X1 U19390 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16440), .ZN(n16418) );
  OAI21_X1 U19391 ( .B1(n16419), .B2(n16443), .A(n16418), .ZN(U236) );
  INV_X1 U19392 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16421) );
  AOI22_X1 U19393 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16440), .ZN(n16420) );
  OAI21_X1 U19394 ( .B1(n16421), .B2(n16443), .A(n16420), .ZN(U237) );
  INV_X1 U19395 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16423) );
  AOI22_X1 U19396 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16440), .ZN(n16422) );
  OAI21_X1 U19397 ( .B1(n16423), .B2(n16443), .A(n16422), .ZN(U238) );
  AOI22_X1 U19398 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16440), .ZN(n16424) );
  OAI21_X1 U19399 ( .B1(n16425), .B2(n16443), .A(n16424), .ZN(U239) );
  INV_X1 U19400 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16427) );
  AOI22_X1 U19401 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16440), .ZN(n16426) );
  OAI21_X1 U19402 ( .B1(n16427), .B2(n16443), .A(n16426), .ZN(U240) );
  INV_X1 U19403 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16429) );
  AOI22_X1 U19404 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16440), .ZN(n16428) );
  OAI21_X1 U19405 ( .B1(n16429), .B2(n16443), .A(n16428), .ZN(U241) );
  AOI22_X1 U19406 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16440), .ZN(n16430) );
  OAI21_X1 U19407 ( .B1(n16431), .B2(n16443), .A(n16430), .ZN(U242) );
  INV_X1 U19408 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16433) );
  AOI22_X1 U19409 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16440), .ZN(n16432) );
  OAI21_X1 U19410 ( .B1(n16433), .B2(n16443), .A(n16432), .ZN(U243) );
  INV_X1 U19411 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16435) );
  AOI22_X1 U19412 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16440), .ZN(n16434) );
  OAI21_X1 U19413 ( .B1(n16435), .B2(n16443), .A(n16434), .ZN(U244) );
  INV_X1 U19414 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16437) );
  AOI22_X1 U19415 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16440), .ZN(n16436) );
  OAI21_X1 U19416 ( .B1(n16437), .B2(n16443), .A(n16436), .ZN(U245) );
  INV_X1 U19417 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16439) );
  AOI22_X1 U19418 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16440), .ZN(n16438) );
  OAI21_X1 U19419 ( .B1(n16439), .B2(n16443), .A(n16438), .ZN(U246) );
  INV_X1 U19420 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16444) );
  AOI22_X1 U19421 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16441), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16440), .ZN(n16442) );
  OAI21_X1 U19422 ( .B1(n16444), .B2(n16443), .A(n16442), .ZN(U247) );
  OAI22_X1 U19423 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16477), .ZN(n16445) );
  INV_X1 U19424 ( .A(n16445), .ZN(U251) );
  OAI22_X1 U19425 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16477), .ZN(n16446) );
  INV_X1 U19426 ( .A(n16446), .ZN(U252) );
  OAI22_X1 U19427 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16477), .ZN(n16447) );
  INV_X1 U19428 ( .A(n16447), .ZN(U253) );
  OAI22_X1 U19429 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16477), .ZN(n16448) );
  INV_X1 U19430 ( .A(n16448), .ZN(U254) );
  OAI22_X1 U19431 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16477), .ZN(n16449) );
  INV_X1 U19432 ( .A(n16449), .ZN(U255) );
  OAI22_X1 U19433 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16477), .ZN(n16450) );
  INV_X1 U19434 ( .A(n16450), .ZN(U256) );
  OAI22_X1 U19435 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16477), .ZN(n16451) );
  INV_X1 U19436 ( .A(n16451), .ZN(U257) );
  OAI22_X1 U19437 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16477), .ZN(n16452) );
  INV_X1 U19438 ( .A(n16452), .ZN(U258) );
  OAI22_X1 U19439 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16477), .ZN(n16453) );
  INV_X1 U19440 ( .A(n16453), .ZN(U259) );
  OAI22_X1 U19441 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16468), .ZN(n16454) );
  INV_X1 U19442 ( .A(n16454), .ZN(U260) );
  OAI22_X1 U19443 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16468), .ZN(n16455) );
  INV_X1 U19444 ( .A(n16455), .ZN(U261) );
  OAI22_X1 U19445 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16477), .ZN(n16456) );
  INV_X1 U19446 ( .A(n16456), .ZN(U262) );
  OAI22_X1 U19447 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16468), .ZN(n16457) );
  INV_X1 U19448 ( .A(n16457), .ZN(U263) );
  OAI22_X1 U19449 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16477), .ZN(n16458) );
  INV_X1 U19450 ( .A(n16458), .ZN(U264) );
  OAI22_X1 U19451 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16477), .ZN(n16459) );
  INV_X1 U19452 ( .A(n16459), .ZN(U265) );
  OAI22_X1 U19453 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16468), .ZN(n16460) );
  INV_X1 U19454 ( .A(n16460), .ZN(U266) );
  OAI22_X1 U19455 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16468), .ZN(n16461) );
  INV_X1 U19456 ( .A(n16461), .ZN(U267) );
  OAI22_X1 U19457 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16468), .ZN(n16462) );
  INV_X1 U19458 ( .A(n16462), .ZN(U268) );
  OAI22_X1 U19459 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16468), .ZN(n16463) );
  INV_X1 U19460 ( .A(n16463), .ZN(U269) );
  OAI22_X1 U19461 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16468), .ZN(n16464) );
  INV_X1 U19462 ( .A(n16464), .ZN(U270) );
  OAI22_X1 U19463 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16468), .ZN(n16465) );
  INV_X1 U19464 ( .A(n16465), .ZN(U271) );
  OAI22_X1 U19465 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16477), .ZN(n16466) );
  INV_X1 U19466 ( .A(n16466), .ZN(U272) );
  OAI22_X1 U19467 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16477), .ZN(n16467) );
  INV_X1 U19468 ( .A(n16467), .ZN(U273) );
  OAI22_X1 U19469 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16468), .ZN(n16469) );
  INV_X1 U19470 ( .A(n16469), .ZN(U274) );
  OAI22_X1 U19471 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16477), .ZN(n16470) );
  INV_X1 U19472 ( .A(n16470), .ZN(U275) );
  OAI22_X1 U19473 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16477), .ZN(n16471) );
  INV_X1 U19474 ( .A(n16471), .ZN(U276) );
  INV_X1 U19475 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n19102) );
  AOI22_X1 U19476 ( .A1(n16477), .A2(n20709), .B1(n19102), .B2(U215), .ZN(U277) );
  OAI22_X1 U19477 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16477), .ZN(n16472) );
  INV_X1 U19478 ( .A(n16472), .ZN(U278) );
  OAI22_X1 U19479 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16477), .ZN(n16473) );
  INV_X1 U19480 ( .A(n16473), .ZN(U279) );
  OAI22_X1 U19481 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16477), .ZN(n16474) );
  INV_X1 U19482 ( .A(n16474), .ZN(U280) );
  OAI22_X1 U19483 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16477), .ZN(n16475) );
  INV_X1 U19484 ( .A(n16475), .ZN(U281) );
  AOI22_X1 U19485 ( .A1(n16477), .A2(n16479), .B1(n18200), .B2(U215), .ZN(U282) );
  INV_X1 U19486 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16478) );
  AOI222_X1 U19487 ( .A1(n16480), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16479), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16478), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16481) );
  INV_X2 U19488 ( .A(n16483), .ZN(n16482) );
  INV_X1 U19489 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18702) );
  INV_X1 U19490 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19663) );
  AOI22_X1 U19491 ( .A1(n16482), .A2(n18702), .B1(n19663), .B2(n16483), .ZN(
        U347) );
  INV_X1 U19492 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18700) );
  INV_X1 U19493 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19662) );
  AOI22_X1 U19494 ( .A1(n16481), .A2(n18700), .B1(n19662), .B2(n16483), .ZN(
        U348) );
  INV_X1 U19495 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18697) );
  INV_X1 U19496 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19661) );
  AOI22_X1 U19497 ( .A1(n16482), .A2(n18697), .B1(n19661), .B2(n16483), .ZN(
        U349) );
  INV_X1 U19498 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18696) );
  INV_X1 U19499 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19660) );
  AOI22_X1 U19500 ( .A1(n16482), .A2(n18696), .B1(n19660), .B2(n16483), .ZN(
        U350) );
  INV_X1 U19501 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18695) );
  INV_X1 U19502 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19658) );
  AOI22_X1 U19503 ( .A1(n16482), .A2(n18695), .B1(n19658), .B2(n16483), .ZN(
        U351) );
  INV_X1 U19504 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18693) );
  INV_X1 U19505 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19656) );
  AOI22_X1 U19506 ( .A1(n16482), .A2(n18693), .B1(n19656), .B2(n16483), .ZN(
        U352) );
  INV_X1 U19507 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18691) );
  INV_X1 U19508 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19654) );
  AOI22_X1 U19509 ( .A1(n16482), .A2(n18691), .B1(n19654), .B2(n16483), .ZN(
        U353) );
  INV_X1 U19510 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18689) );
  AOI22_X1 U19511 ( .A1(n16482), .A2(n18689), .B1(n19653), .B2(n16483), .ZN(
        U354) );
  INV_X1 U19512 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18741) );
  INV_X1 U19513 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20825) );
  AOI22_X1 U19514 ( .A1(n16482), .A2(n18741), .B1(n20825), .B2(n16483), .ZN(
        U355) );
  INV_X1 U19515 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18738) );
  INV_X1 U19516 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19694) );
  AOI22_X1 U19517 ( .A1(n16482), .A2(n18738), .B1(n19694), .B2(n16483), .ZN(
        U356) );
  INV_X1 U19518 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18735) );
  INV_X1 U19519 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19692) );
  AOI22_X1 U19520 ( .A1(n16482), .A2(n18735), .B1(n19692), .B2(n16483), .ZN(
        U357) );
  INV_X1 U19521 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18734) );
  INV_X1 U19522 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19689) );
  AOI22_X1 U19523 ( .A1(n16482), .A2(n18734), .B1(n19689), .B2(n16483), .ZN(
        U358) );
  INV_X1 U19524 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18732) );
  INV_X1 U19525 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20769) );
  AOI22_X1 U19526 ( .A1(n16482), .A2(n18732), .B1(n20769), .B2(n16483), .ZN(
        U359) );
  INV_X1 U19527 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18730) );
  INV_X1 U19528 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19687) );
  AOI22_X1 U19529 ( .A1(n16482), .A2(n18730), .B1(n19687), .B2(n16483), .ZN(
        U360) );
  INV_X1 U19530 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18728) );
  INV_X1 U19531 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19685) );
  AOI22_X1 U19532 ( .A1(n16482), .A2(n18728), .B1(n19685), .B2(n16483), .ZN(
        U361) );
  INV_X1 U19533 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18726) );
  INV_X1 U19534 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19683) );
  AOI22_X1 U19535 ( .A1(n16482), .A2(n18726), .B1(n19683), .B2(n16483), .ZN(
        U362) );
  INV_X1 U19536 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18724) );
  INV_X1 U19537 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19681) );
  AOI22_X1 U19538 ( .A1(n16482), .A2(n18724), .B1(n19681), .B2(n16483), .ZN(
        U363) );
  INV_X1 U19539 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18722) );
  INV_X1 U19540 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19679) );
  AOI22_X1 U19541 ( .A1(n16482), .A2(n18722), .B1(n19679), .B2(n16483), .ZN(
        U364) );
  INV_X1 U19542 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18687) );
  INV_X1 U19543 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19651) );
  AOI22_X1 U19544 ( .A1(n16482), .A2(n18687), .B1(n19651), .B2(n16483), .ZN(
        U365) );
  INV_X1 U19545 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18720) );
  INV_X1 U19546 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19678) );
  AOI22_X1 U19547 ( .A1(n16482), .A2(n18720), .B1(n19678), .B2(n16483), .ZN(
        U366) );
  INV_X1 U19548 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n20760) );
  INV_X1 U19549 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19676) );
  AOI22_X1 U19550 ( .A1(n16482), .A2(n20760), .B1(n19676), .B2(n16483), .ZN(
        U367) );
  INV_X1 U19551 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18718) );
  INV_X1 U19552 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19674) );
  AOI22_X1 U19553 ( .A1(n16482), .A2(n18718), .B1(n19674), .B2(n16483), .ZN(
        U368) );
  INV_X1 U19554 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18715) );
  INV_X1 U19555 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19672) );
  AOI22_X1 U19556 ( .A1(n16482), .A2(n18715), .B1(n19672), .B2(n16483), .ZN(
        U369) );
  INV_X1 U19557 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18714) );
  INV_X1 U19558 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19670) );
  AOI22_X1 U19559 ( .A1(n16482), .A2(n18714), .B1(n19670), .B2(n16483), .ZN(
        U370) );
  INV_X1 U19560 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18712) );
  INV_X1 U19561 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19668) );
  AOI22_X1 U19562 ( .A1(n16481), .A2(n18712), .B1(n19668), .B2(n16483), .ZN(
        U371) );
  INV_X1 U19563 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18709) );
  INV_X1 U19564 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20755) );
  AOI22_X1 U19565 ( .A1(n16482), .A2(n18709), .B1(n20755), .B2(n16483), .ZN(
        U372) );
  INV_X1 U19566 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18708) );
  INV_X1 U19567 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19665) );
  AOI22_X1 U19568 ( .A1(n16482), .A2(n18708), .B1(n19665), .B2(n16483), .ZN(
        U373) );
  INV_X1 U19569 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18706) );
  INV_X1 U19570 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19664) );
  AOI22_X1 U19571 ( .A1(n16482), .A2(n18706), .B1(n19664), .B2(n16483), .ZN(
        U374) );
  INV_X1 U19572 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18704) );
  INV_X1 U19573 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20824) );
  AOI22_X1 U19574 ( .A1(n16481), .A2(n18704), .B1(n20824), .B2(n16483), .ZN(
        U375) );
  INV_X1 U19575 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18684) );
  INV_X1 U19576 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19650) );
  AOI22_X1 U19577 ( .A1(n16481), .A2(n18684), .B1(n19650), .B2(n16483), .ZN(
        U376) );
  INV_X1 U19578 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18683) );
  NAND2_X1 U19579 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18683), .ZN(n18673) );
  AOI22_X1 U19580 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18673), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18677), .ZN(n18750) );
  AOI21_X1 U19581 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18750), .ZN(n16484) );
  INV_X1 U19582 ( .A(n16484), .ZN(P3_U2633) );
  NAND2_X1 U19583 ( .A1(n18821), .A2(n18820), .ZN(n16488) );
  AND2_X1 U19584 ( .A1(n16486), .A2(n16485), .ZN(n16492) );
  OAI21_X1 U19585 ( .B1(n16492), .B2(n17398), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16487) );
  OAI21_X1 U19586 ( .B1(n16488), .B2(n18808), .A(n16487), .ZN(P3_U2634) );
  AOI21_X1 U19587 ( .B1(n18677), .B2(n18683), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16489) );
  AOI22_X1 U19588 ( .A1(n18817), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16489), 
        .B2(n18818), .ZN(P3_U2635) );
  NOR2_X1 U19589 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18669) );
  OAI21_X1 U19590 ( .B1(n18669), .B2(BS16), .A(n18750), .ZN(n18748) );
  OAI21_X1 U19591 ( .B1(n18750), .B2(n16515), .A(n18748), .ZN(P3_U2636) );
  INV_X1 U19592 ( .A(n16490), .ZN(n16493) );
  NOR3_X1 U19593 ( .A1(n16493), .A2(n16492), .A3(n16491), .ZN(n18603) );
  NOR2_X1 U19594 ( .A1(n18603), .A2(n18658), .ZN(n18801) );
  INV_X1 U19595 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18149) );
  OAI21_X1 U19596 ( .B1(n18801), .B2(n18149), .A(n16494), .ZN(P3_U2637) );
  NOR4_X1 U19597 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n16498) );
  NOR4_X1 U19598 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16497) );
  NOR4_X1 U19599 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n16496) );
  NOR4_X1 U19600 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16495) );
  NAND4_X1 U19601 ( .A1(n16498), .A2(n16497), .A3(n16496), .A4(n16495), .ZN(
        n16504) );
  NOR4_X1 U19602 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16502) );
  AOI211_X1 U19603 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16501) );
  NOR4_X1 U19604 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16500) );
  NOR4_X1 U19605 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16499) );
  NAND4_X1 U19606 ( .A1(n16502), .A2(n16501), .A3(n16500), .A4(n16499), .ZN(
        n16503) );
  NOR2_X1 U19607 ( .A1(n16504), .A2(n16503), .ZN(n18792) );
  INV_X1 U19608 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16506) );
  NOR3_X1 U19609 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16507) );
  OAI21_X1 U19610 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16507), .A(n18792), .ZN(
        n16505) );
  OAI21_X1 U19611 ( .B1(n18792), .B2(n16506), .A(n16505), .ZN(P3_U2638) );
  INV_X1 U19612 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18685) );
  INV_X1 U19613 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18749) );
  AOI21_X1 U19614 ( .B1(n18685), .B2(n18749), .A(n16507), .ZN(n16509) );
  INV_X1 U19615 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16508) );
  INV_X1 U19616 ( .A(n18792), .ZN(n18789) );
  AOI22_X1 U19617 ( .A1(n18792), .A2(n16509), .B1(n16508), .B2(n18789), .ZN(
        P3_U2639) );
  NAND2_X1 U19618 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18763), .ZN(n16510) );
  NOR2_X1 U19619 ( .A1(n18752), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18539) );
  INV_X1 U19620 ( .A(n18539), .ZN(n18435) );
  NOR3_X1 U19621 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n18666) );
  NOR2_X1 U19622 ( .A1(n9846), .A2(n18661), .ZN(n16776) );
  INV_X1 U19623 ( .A(n18823), .ZN(n18810) );
  OAI211_X1 U19624 ( .C1(n18804), .C2(n18803), .A(n18814), .B(n16515), .ZN(
        n16511) );
  INV_X1 U19625 ( .A(n16511), .ZN(n18653) );
  AOI211_X4 U19626 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18804), .A(n18653), .B(
        n16514), .ZN(n16843) );
  INV_X1 U19627 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18729) );
  INV_X1 U19628 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18725) );
  INV_X1 U19629 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18710) );
  INV_X1 U19630 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18707) );
  INV_X1 U19631 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18694) );
  INV_X1 U19632 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18690) );
  NAND3_X1 U19633 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16832) );
  NOR2_X1 U19634 ( .A1(n18690), .A2(n16832), .ZN(n16808) );
  NAND2_X1 U19635 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16808), .ZN(n16797) );
  NOR2_X1 U19636 ( .A1(n18694), .A2(n16797), .ZN(n16782) );
  NAND3_X1 U19637 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_8__SCAN_IN), 
        .A3(n16782), .ZN(n16750) );
  NAND2_X1 U19638 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16751) );
  NOR3_X1 U19639 ( .A1(n18703), .A2(n16750), .A3(n16751), .ZN(n16725) );
  NAND2_X1 U19640 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16725), .ZN(n16703) );
  NOR3_X1 U19641 ( .A1(n18710), .A2(n18707), .A3(n16703), .ZN(n16651) );
  NAND3_X1 U19642 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16659) );
  NAND2_X1 U19643 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16660) );
  NOR2_X1 U19644 ( .A1(n16659), .A2(n16660), .ZN(n16648) );
  NAND3_X1 U19645 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16651), .A3(n16648), 
        .ZN(n16625) );
  NAND2_X1 U19646 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n16613) );
  NOR3_X1 U19647 ( .A1(n18725), .A2(n16625), .A3(n16613), .ZN(n16605) );
  NAND2_X1 U19648 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16605), .ZN(n16594) );
  NOR2_X1 U19649 ( .A1(n18729), .A2(n16594), .ZN(n16583) );
  NAND2_X1 U19650 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16583), .ZN(n16533) );
  NOR2_X1 U19651 ( .A1(n16868), .A2(n16533), .ZN(n16576) );
  NAND4_X1 U19652 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16576), .ZN(n16535) );
  NOR3_X1 U19653 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18742), .A3(n16535), 
        .ZN(n16512) );
  AOI21_X1 U19654 ( .B1(n16843), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16512), .ZN(
        n16540) );
  NAND2_X1 U19655 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18804), .ZN(n16513) );
  AOI211_X4 U19656 ( .C1(n16515), .C2(n18814), .A(n16514), .B(n16513), .ZN(
        n16845) );
  NOR3_X1 U19657 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16852) );
  INV_X1 U19658 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16846) );
  NAND2_X1 U19659 ( .A1(n16852), .A2(n16846), .ZN(n16844) );
  NOR2_X1 U19660 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16844), .ZN(n16820) );
  NAND2_X1 U19661 ( .A1(n16820), .A2(n16812), .ZN(n16811) );
  NOR2_X1 U19662 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16811), .ZN(n16795) );
  NAND2_X1 U19663 ( .A1(n16795), .A2(n16794), .ZN(n16791) );
  NOR2_X1 U19664 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16791), .ZN(n16771) );
  NAND2_X1 U19665 ( .A1(n16771), .A2(n17056), .ZN(n16760) );
  INV_X1 U19666 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17118) );
  NAND2_X1 U19667 ( .A1(n16748), .A2(n17118), .ZN(n16743) );
  NAND2_X1 U19668 ( .A1(n16730), .A2(n17070), .ZN(n16721) );
  NAND2_X1 U19669 ( .A1(n16704), .A2(n20697), .ZN(n16700) );
  INV_X1 U19670 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16679) );
  NAND2_X1 U19671 ( .A1(n16686), .A2(n16679), .ZN(n16678) );
  INV_X1 U19672 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16656) );
  NAND2_X1 U19673 ( .A1(n16663), .A2(n16656), .ZN(n16654) );
  INV_X1 U19674 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16976) );
  NAND2_X1 U19675 ( .A1(n16643), .A2(n16976), .ZN(n16635) );
  NAND2_X1 U19676 ( .A1(n16623), .A2(n16883), .ZN(n16619) );
  INV_X1 U19677 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16887) );
  NAND2_X1 U19678 ( .A1(n16612), .A2(n16887), .ZN(n16599) );
  NOR2_X1 U19679 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16599), .ZN(n16584) );
  INV_X1 U19680 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16578) );
  NAND2_X1 U19681 ( .A1(n16584), .A2(n16578), .ZN(n16577) );
  NOR2_X1 U19682 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16577), .ZN(n16562) );
  INV_X1 U19683 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16888) );
  NAND2_X1 U19684 ( .A1(n16562), .A2(n16888), .ZN(n16542) );
  NOR2_X1 U19685 ( .A1(n16874), .A2(n16542), .ZN(n16548) );
  INV_X1 U19686 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16894) );
  INV_X1 U19687 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16517) );
  NAND2_X1 U19688 ( .A1(n9732), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16518) );
  AOI21_X1 U19689 ( .B1(n16517), .B2(n16518), .A(n16516), .ZN(n17461) );
  OAI21_X1 U19690 ( .B1(n9732), .B2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16518), .ZN(n17479) );
  INV_X1 U19691 ( .A(n17479), .ZN(n16573) );
  NAND2_X1 U19692 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17487), .ZN(
        n17460) );
  AOI21_X1 U19693 ( .B1(n9944), .B2(n17460), .A(n9732), .ZN(n17491) );
  INV_X1 U19694 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16595) );
  INV_X1 U19695 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17513) );
  NOR2_X1 U19696 ( .A1(n17804), .A2(n9702), .ZN(n16525) );
  AND2_X1 U19697 ( .A1(n17538), .A2(n16525), .ZN(n17497) );
  NAND2_X1 U19698 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17497), .ZN(
        n16521) );
  OR2_X1 U19699 ( .A1(n17513), .A2(n16521), .ZN(n16520) );
  INV_X1 U19700 ( .A(n17460), .ZN(n16519) );
  AOI21_X1 U19701 ( .B1(n16595), .B2(n16520), .A(n16519), .ZN(n17499) );
  XOR2_X1 U19702 ( .A(n17513), .B(n16521), .Z(n17509) );
  OAI21_X1 U19703 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17497), .A(
        n16521), .ZN(n16522) );
  INV_X1 U19704 ( .A(n16522), .ZN(n17525) );
  NAND2_X1 U19705 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16525), .ZN(
        n16523) );
  AOI21_X1 U19706 ( .B1(n17544), .B2(n16523), .A(n17497), .ZN(n17542) );
  XNOR2_X1 U19707 ( .A(n20720), .B(n16525), .ZN(n17555) );
  INV_X1 U19708 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17541) );
  NAND2_X1 U19709 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16524), .ZN(
        n17539) );
  AOI21_X1 U19710 ( .B1(n17541), .B2(n17539), .A(n16525), .ZN(n17565) );
  INV_X1 U19711 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17578) );
  INV_X1 U19712 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16682) );
  NAND2_X1 U19713 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16526), .ZN(
        n16529) );
  NOR2_X1 U19714 ( .A1(n16682), .A2(n16529), .ZN(n16528) );
  NAND2_X1 U19715 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16528), .ZN(
        n16527) );
  AOI22_X1 U19716 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16524), .B1(
        n17578), .B2(n16527), .ZN(n17573) );
  INV_X1 U19717 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17585) );
  INV_X1 U19718 ( .A(n16528), .ZN(n17572) );
  XOR2_X1 U19719 ( .A(n17585), .B(n17572), .Z(n17588) );
  AOI21_X1 U19720 ( .B1(n16682), .B2(n16529), .A(n16528), .ZN(n17600) );
  INV_X1 U19721 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16530) );
  NOR2_X1 U19722 ( .A1(n17804), .A2(n16738), .ZN(n16747) );
  NAND2_X1 U19723 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n16747), .ZN(
        n17647) );
  INV_X1 U19724 ( .A(n17647), .ZN(n16727) );
  AND2_X1 U19725 ( .A1(n16694), .A2(n16727), .ZN(n17607) );
  NAND2_X1 U19726 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17607), .ZN(
        n16693) );
  AOI22_X1 U19727 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16526), .B1(
        n16530), .B2(n16693), .ZN(n17608) );
  OAI21_X1 U19728 ( .B1(n16693), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n16531), .ZN(n16532) );
  INV_X1 U19729 ( .A(n16532), .ZN(n16685) );
  NOR2_X1 U19730 ( .A1(n17608), .A2(n16685), .ZN(n16684) );
  NOR2_X1 U19731 ( .A1(n17600), .A2(n16673), .ZN(n16672) );
  NOR2_X1 U19732 ( .A1(n16672), .A2(n16837), .ZN(n16667) );
  NOR2_X1 U19733 ( .A1(n17588), .A2(n16667), .ZN(n16666) );
  NOR2_X1 U19734 ( .A1(n16666), .A2(n16837), .ZN(n16653) );
  NOR2_X1 U19735 ( .A1(n17573), .A2(n16653), .ZN(n16652) );
  NOR2_X1 U19736 ( .A1(n16652), .A2(n16837), .ZN(n16642) );
  NOR2_X1 U19737 ( .A1(n17565), .A2(n16642), .ZN(n16641) );
  NOR2_X1 U19738 ( .A1(n17542), .A2(n16627), .ZN(n16626) );
  NOR2_X1 U19739 ( .A1(n16626), .A2(n16837), .ZN(n16615) );
  NOR2_X1 U19740 ( .A1(n17525), .A2(n16615), .ZN(n16614) );
  NOR2_X1 U19741 ( .A1(n16614), .A2(n16837), .ZN(n16607) );
  NOR2_X1 U19742 ( .A1(n17509), .A2(n16607), .ZN(n16606) );
  NOR2_X1 U19743 ( .A1(n16606), .A2(n16837), .ZN(n16593) );
  NOR2_X1 U19744 ( .A1(n17499), .A2(n16593), .ZN(n16592) );
  NOR2_X1 U19745 ( .A1(n16592), .A2(n16837), .ZN(n16586) );
  NOR2_X1 U19746 ( .A1(n17491), .A2(n16586), .ZN(n16585) );
  NOR2_X1 U19747 ( .A1(n16563), .A2(n16837), .ZN(n16552) );
  NAND2_X1 U19748 ( .A1(n16531), .A2(n18661), .ZN(n16866) );
  NOR3_X1 U19749 ( .A1(n16544), .A2(n16543), .A3(n16866), .ZN(n16538) );
  NAND3_X1 U19750 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16534) );
  AND2_X1 U19751 ( .A1(n16833), .A2(n16533), .ZN(n16582) );
  NOR2_X1 U19752 ( .A1(n16877), .A2(n16582), .ZN(n16581) );
  INV_X1 U19753 ( .A(n16581), .ZN(n16589) );
  AOI21_X1 U19754 ( .B1(n16833), .B2(n16534), .A(n16589), .ZN(n16561) );
  NOR2_X1 U19755 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16535), .ZN(n16547) );
  INV_X1 U19756 ( .A(n16547), .ZN(n16536) );
  AOI21_X1 U19757 ( .B1(n16561), .B2(n16536), .A(n18740), .ZN(n16537) );
  OAI211_X1 U19758 ( .C1(n16541), .C2(n16865), .A(n16540), .B(n16539), .ZN(
        P3_U2640) );
  NAND2_X1 U19759 ( .A1(n16845), .A2(n16542), .ZN(n16557) );
  OAI22_X1 U19760 ( .A1(n16561), .A2(n18742), .B1(n16545), .B2(n16865), .ZN(
        n16546) );
  OAI21_X1 U19761 ( .B1(n16843), .B2(n16548), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16549) );
  OAI211_X1 U19762 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16557), .A(n16550), .B(
        n16549), .ZN(P3_U2641) );
  INV_X1 U19763 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18737) );
  AOI211_X1 U19764 ( .C1(n16553), .C2(n16552), .A(n16551), .B(n16839), .ZN(
        n16556) );
  NAND3_X1 U19765 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16576), .ZN(n16554) );
  OAI22_X1 U19766 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16554), .B1(n20747), 
        .B2(n16865), .ZN(n16555) );
  AOI211_X1 U19767 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16843), .A(n16556), .B(
        n16555), .ZN(n16560) );
  INV_X1 U19768 ( .A(n16557), .ZN(n16558) );
  OAI21_X1 U19769 ( .B1(n16562), .B2(n16888), .A(n16558), .ZN(n16559) );
  OAI211_X1 U19770 ( .C1(n16561), .C2(n18737), .A(n16560), .B(n16559), .ZN(
        P3_U2642) );
  AOI22_X1 U19771 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16824), .B1(
        n16843), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16570) );
  AOI211_X1 U19772 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16577), .A(n16562), .B(
        n16874), .ZN(n16566) );
  AOI211_X1 U19773 ( .C1(n17461), .C2(n16564), .A(n16563), .B(n16839), .ZN(
        n16565) );
  AOI211_X1 U19774 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16589), .A(n16566), 
        .B(n16565), .ZN(n16569) );
  NAND2_X1 U19775 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16567) );
  OAI211_X1 U19776 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16576), .B(n16567), .ZN(n16568) );
  NAND3_X1 U19777 ( .A1(n16570), .A2(n16569), .A3(n16568), .ZN(P3_U2643) );
  INV_X1 U19778 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18733) );
  AOI211_X1 U19779 ( .C1(n16573), .C2(n16572), .A(n16571), .B(n16839), .ZN(
        n16575) );
  INV_X1 U19780 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17482) );
  OAI22_X1 U19781 ( .A1(n17482), .A2(n16865), .B1(n16875), .B2(n16578), .ZN(
        n16574) );
  AOI211_X1 U19782 ( .C1(n16576), .C2(n18733), .A(n16575), .B(n16574), .ZN(
        n16580) );
  OAI211_X1 U19783 ( .C1(n16584), .C2(n16578), .A(n16845), .B(n16577), .ZN(
        n16579) );
  OAI211_X1 U19784 ( .C1(n16581), .C2(n18733), .A(n16580), .B(n16579), .ZN(
        P3_U2644) );
  AOI22_X1 U19785 ( .A1(n16843), .A2(P3_EBX_REG_26__SCAN_IN), .B1(n16583), 
        .B2(n16582), .ZN(n16591) );
  AOI211_X1 U19786 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16599), .A(n16584), .B(
        n16874), .ZN(n16588) );
  AOI211_X1 U19787 ( .C1(n17491), .C2(n16586), .A(n16585), .B(n16839), .ZN(
        n16587) );
  AOI211_X1 U19788 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16589), .A(n16588), 
        .B(n16587), .ZN(n16590) );
  OAI211_X1 U19789 ( .C1(n9944), .C2(n16865), .A(n16591), .B(n16590), .ZN(
        P3_U2645) );
  INV_X1 U19790 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18727) );
  OAI21_X1 U19791 ( .B1(n16605), .B2(n16868), .A(n16855), .ZN(n16618) );
  AOI21_X1 U19792 ( .B1(n16833), .B2(n18727), .A(n16618), .ZN(n16602) );
  AOI211_X1 U19793 ( .C1(n17499), .C2(n16593), .A(n16592), .B(n16839), .ZN(
        n16598) );
  NOR3_X1 U19794 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16868), .A3(n16594), 
        .ZN(n16597) );
  OAI22_X1 U19795 ( .A1(n16595), .A2(n16865), .B1(n16875), .B2(n16887), .ZN(
        n16596) );
  NOR3_X1 U19796 ( .A1(n16598), .A2(n16597), .A3(n16596), .ZN(n16601) );
  OAI211_X1 U19797 ( .C1(n16612), .C2(n16887), .A(n16845), .B(n16599), .ZN(
        n16600) );
  OAI211_X1 U19798 ( .C1(n16602), .C2(n18729), .A(n16601), .B(n16600), .ZN(
        P3_U2646) );
  AOI21_X1 U19799 ( .B1(n16619), .B2(P3_EBX_REG_24__SCAN_IN), .A(n16874), .ZN(
        n16603) );
  AOI21_X1 U19800 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16843), .A(n16603), .ZN(
        n16611) );
  NOR2_X1 U19801 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16868), .ZN(n16604) );
  AOI22_X1 U19802 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16824), .B1(
        n16605), .B2(n16604), .ZN(n16610) );
  AOI211_X1 U19803 ( .C1(n17509), .C2(n16607), .A(n16606), .B(n16839), .ZN(
        n16608) );
  AOI21_X1 U19804 ( .B1(n16618), .B2(P3_REIP_REG_24__SCAN_IN), .A(n16608), 
        .ZN(n16609) );
  OAI211_X1 U19805 ( .C1(n16612), .C2(n16611), .A(n16610), .B(n16609), .ZN(
        P3_U2647) );
  AOI22_X1 U19806 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n16824), .B1(
        n16843), .B2(P3_EBX_REG_23__SCAN_IN), .ZN(n16622) );
  NAND2_X1 U19807 ( .A1(n16833), .A2(n16651), .ZN(n16687) );
  NAND3_X1 U19808 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16648), .A3(n16696), 
        .ZN(n16640) );
  NOR2_X1 U19809 ( .A1(n16613), .A2(n16640), .ZN(n16617) );
  AOI211_X1 U19810 ( .C1(n17525), .C2(n16615), .A(n16614), .B(n16839), .ZN(
        n16616) );
  AOI221_X1 U19811 ( .B1(n16618), .B2(P3_REIP_REG_23__SCAN_IN), .C1(n16617), 
        .C2(n18725), .A(n16616), .ZN(n16621) );
  OAI211_X1 U19812 ( .C1(n16623), .C2(n16883), .A(n16845), .B(n16619), .ZN(
        n16620) );
  NAND3_X1 U19813 ( .A1(n16622), .A2(n16621), .A3(n16620), .ZN(P3_U2648) );
  AOI211_X1 U19814 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16635), .A(n16623), .B(
        n16874), .ZN(n16624) );
  AOI21_X1 U19815 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n16843), .A(n16624), .ZN(
        n16632) );
  AOI21_X1 U19816 ( .B1(n16833), .B2(n16625), .A(n16877), .ZN(n16646) );
  OAI21_X1 U19817 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n16640), .A(n16646), 
        .ZN(n16630) );
  INV_X1 U19818 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18721) );
  NOR3_X1 U19819 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n18721), .A3(n16640), 
        .ZN(n16629) );
  AOI211_X1 U19820 ( .C1(n17542), .C2(n16627), .A(n16626), .B(n16839), .ZN(
        n16628) );
  AOI211_X1 U19821 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16630), .A(n16629), 
        .B(n16628), .ZN(n16631) );
  OAI211_X1 U19822 ( .C1(n17544), .C2(n16865), .A(n16632), .B(n16631), .ZN(
        P3_U2649) );
  AOI211_X1 U19823 ( .C1(n17555), .C2(n16634), .A(n16633), .B(n16839), .ZN(
        n16638) );
  OAI211_X1 U19824 ( .C1(n16643), .C2(n16976), .A(n16845), .B(n16635), .ZN(
        n16636) );
  OAI21_X1 U19825 ( .B1(n16976), .B2(n16875), .A(n16636), .ZN(n16637) );
  AOI211_X1 U19826 ( .C1(n16824), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16638), .B(n16637), .ZN(n16639) );
  OAI221_X1 U19827 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n16640), .C1(n18721), 
        .C2(n16646), .A(n16639), .ZN(P3_U2650) );
  INV_X1 U19828 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16885) );
  AOI211_X1 U19829 ( .C1(n17565), .C2(n16642), .A(n16641), .B(n16839), .ZN(
        n16645) );
  AOI211_X1 U19830 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16654), .A(n16643), .B(
        n16874), .ZN(n16644) );
  AOI211_X1 U19831 ( .C1(n16824), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16645), .B(n16644), .ZN(n16650) );
  INV_X1 U19832 ( .A(n16646), .ZN(n16647) );
  OAI221_X1 U19833 ( .B1(P3_REIP_REG_20__SCAN_IN), .B2(n16648), .C1(
        P3_REIP_REG_20__SCAN_IN), .C2(n16696), .A(n16647), .ZN(n16649) );
  OAI211_X1 U19834 ( .C1(n16885), .C2(n16875), .A(n16650), .B(n16649), .ZN(
        P3_U2651) );
  NAND2_X1 U19835 ( .A1(n16868), .A2(n16855), .ZN(n16880) );
  OAI21_X1 U19836 ( .B1(n16651), .B2(n16868), .A(n16855), .ZN(n16683) );
  AOI21_X1 U19837 ( .B1(n16659), .B2(n16880), .A(n16683), .ZN(n16665) );
  INV_X1 U19838 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18719) );
  AOI211_X1 U19839 ( .C1(n17573), .C2(n16653), .A(n16652), .B(n16839), .ZN(
        n16658) );
  OAI211_X1 U19840 ( .C1(n16663), .C2(n16656), .A(n16845), .B(n16654), .ZN(
        n16655) );
  OAI211_X1 U19841 ( .C1(n16875), .C2(n16656), .A(n18094), .B(n16655), .ZN(
        n16657) );
  AOI211_X1 U19842 ( .C1(n16824), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16658), .B(n16657), .ZN(n16662) );
  NOR2_X1 U19843 ( .A1(n16659), .A2(n16687), .ZN(n16669) );
  OAI211_X1 U19844 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n16669), .B(n16660), .ZN(n16661) );
  OAI211_X1 U19845 ( .C1(n16665), .C2(n18719), .A(n16662), .B(n16661), .ZN(
        P3_U2652) );
  AOI211_X1 U19846 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16678), .A(n16663), .B(
        n16874), .ZN(n16664) );
  AOI211_X1 U19847 ( .C1(n16843), .C2(P3_EBX_REG_18__SCAN_IN), .A(n9846), .B(
        n16664), .ZN(n16671) );
  INV_X1 U19848 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18717) );
  INV_X1 U19849 ( .A(n16665), .ZN(n16677) );
  AOI211_X1 U19850 ( .C1(n17588), .C2(n16667), .A(n16666), .B(n16839), .ZN(
        n16668) );
  AOI221_X1 U19851 ( .B1(n16669), .B2(n18717), .C1(n16677), .C2(
        P3_REIP_REG_18__SCAN_IN), .A(n16668), .ZN(n16670) );
  OAI211_X1 U19852 ( .C1(n17585), .C2(n16865), .A(n16671), .B(n16670), .ZN(
        P3_U2653) );
  AOI211_X1 U19853 ( .C1(n17600), .C2(n16673), .A(n16672), .B(n16839), .ZN(
        n16676) );
  INV_X1 U19854 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18716) );
  NAND4_X1 U19855 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .A3(n16696), .A4(n18716), .ZN(n16674) );
  OAI211_X1 U19856 ( .C1(n16875), .C2(n16679), .A(n18094), .B(n16674), .ZN(
        n16675) );
  AOI211_X1 U19857 ( .C1(P3_REIP_REG_17__SCAN_IN), .C2(n16677), .A(n16676), 
        .B(n16675), .ZN(n16681) );
  OAI211_X1 U19858 ( .C1(n16686), .C2(n16679), .A(n16845), .B(n16678), .ZN(
        n16680) );
  OAI211_X1 U19859 ( .C1(n16865), .C2(n16682), .A(n16681), .B(n16680), .ZN(
        P3_U2654) );
  INV_X1 U19860 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18713) );
  INV_X1 U19861 ( .A(n16683), .ZN(n16709) );
  AOI22_X1 U19862 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16824), .B1(
        n16843), .B2(P3_EBX_REG_16__SCAN_IN), .ZN(n16692) );
  AOI211_X1 U19863 ( .C1(n17608), .C2(n16685), .A(n16684), .B(n16839), .ZN(
        n16690) );
  AOI211_X1 U19864 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16700), .A(n16686), .B(
        n16874), .ZN(n16689) );
  INV_X1 U19865 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18711) );
  AOI221_X1 U19866 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(P3_REIP_REG_15__SCAN_IN), .C1(n18713), .C2(n18711), .A(n16687), .ZN(n16688) );
  NOR4_X1 U19867 ( .A1(n9846), .A2(n16690), .A3(n16689), .A4(n16688), .ZN(
        n16691) );
  OAI211_X1 U19868 ( .C1(n18713), .C2(n16709), .A(n16692), .B(n16691), .ZN(
        P3_U2655) );
  INV_X1 U19869 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17626) );
  OAI21_X1 U19870 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17607), .A(
        n16693), .ZN(n17623) );
  NOR2_X1 U19871 ( .A1(n17804), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16861) );
  INV_X1 U19872 ( .A(n16861), .ZN(n16737) );
  NOR3_X1 U19873 ( .A1(n16738), .A2(n17674), .A3(n16737), .ZN(n16726) );
  AOI21_X1 U19874 ( .B1(n16694), .B2(n16726), .A(n16837), .ZN(n16695) );
  XNOR2_X1 U19875 ( .A(n17623), .B(n16695), .ZN(n16699) );
  AOI22_X1 U19876 ( .A1(n16843), .A2(P3_EBX_REG_15__SCAN_IN), .B1(n16696), 
        .B2(n18711), .ZN(n16697) );
  OAI211_X1 U19877 ( .C1(n18711), .C2(n16709), .A(n16697), .B(n18094), .ZN(
        n16698) );
  AOI21_X1 U19878 ( .B1(n16699), .B2(n18661), .A(n16698), .ZN(n16702) );
  OAI211_X1 U19879 ( .C1(n16704), .C2(n20697), .A(n16845), .B(n16700), .ZN(
        n16701) );
  OAI211_X1 U19880 ( .C1(n16865), .C2(n17626), .A(n16702), .B(n16701), .ZN(
        P3_U2656) );
  NOR2_X1 U19881 ( .A1(n16868), .A2(n16703), .ZN(n16714) );
  AOI21_X1 U19882 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(n16714), .A(
        P3_REIP_REG_14__SCAN_IN), .ZN(n16710) );
  AOI22_X1 U19883 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16824), .B1(
        n16843), .B2(P3_EBX_REG_14__SCAN_IN), .ZN(n16708) );
  INV_X1 U19884 ( .A(n17637), .ZN(n17652) );
  NAND2_X1 U19885 ( .A1(n17652), .A2(n16727), .ZN(n16711) );
  AOI21_X1 U19886 ( .B1(n17636), .B2(n16711), .A(n17607), .ZN(n17639) );
  AOI21_X1 U19887 ( .B1(n17652), .B2(n16726), .A(n16837), .ZN(n16715) );
  XOR2_X1 U19888 ( .A(n17639), .B(n16715), .Z(n16706) );
  AOI211_X1 U19889 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16721), .A(n16704), .B(
        n16874), .ZN(n16705) );
  AOI211_X1 U19890 ( .C1(n18661), .C2(n16706), .A(n9846), .B(n16705), .ZN(
        n16707) );
  OAI211_X1 U19891 ( .C1(n16710), .C2(n16709), .A(n16708), .B(n16707), .ZN(
        P3_U2657) );
  INV_X1 U19892 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20680) );
  NOR2_X1 U19893 ( .A1(n20680), .A2(n17647), .ZN(n16712) );
  OAI21_X1 U19894 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16712), .A(
        n16711), .ZN(n17650) );
  AOI21_X1 U19895 ( .B1(n16531), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n16839), .ZN(n16870) );
  INV_X1 U19896 ( .A(n16870), .ZN(n16713) );
  AOI211_X1 U19897 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n16531), .A(
        n17650), .B(n16713), .ZN(n16720) );
  INV_X1 U19898 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18705) );
  OAI21_X1 U19899 ( .B1(n16725), .B2(n16868), .A(n16855), .ZN(n16741) );
  AOI21_X1 U19900 ( .B1(n16833), .B2(n18705), .A(n16741), .ZN(n16718) );
  AOI21_X1 U19901 ( .B1(n16714), .B2(n18707), .A(n9846), .ZN(n16717) );
  NAND3_X1 U19902 ( .A1(n18661), .A2(n16715), .A3(n17650), .ZN(n16716) );
  OAI211_X1 U19903 ( .C1(n16718), .C2(n18707), .A(n16717), .B(n16716), .ZN(
        n16719) );
  AOI211_X1 U19904 ( .C1(n16824), .C2(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16720), .B(n16719), .ZN(n16723) );
  OAI211_X1 U19905 ( .C1(n16730), .C2(n17070), .A(n16845), .B(n16721), .ZN(
        n16722) );
  OAI211_X1 U19906 ( .C1(n17070), .C2(n16875), .A(n16723), .B(n16722), .ZN(
        P3_U2658) );
  INV_X1 U19907 ( .A(n16741), .ZN(n16735) );
  NOR2_X1 U19908 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16868), .ZN(n16724) );
  AOI22_X1 U19909 ( .A1(n16843), .A2(P3_EBX_REG_12__SCAN_IN), .B1(n16725), 
        .B2(n16724), .ZN(n16734) );
  NOR2_X1 U19910 ( .A1(n16726), .A2(n16837), .ZN(n16728) );
  AOI22_X1 U19911 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17647), .B1(
        n16727), .B2(n20680), .ZN(n17662) );
  XOR2_X1 U19912 ( .A(n16728), .B(n17662), .Z(n16729) );
  OAI21_X1 U19913 ( .B1(n16839), .B2(n16729), .A(n18094), .ZN(n16732) );
  AOI211_X1 U19914 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16743), .A(n16730), .B(
        n16874), .ZN(n16731) );
  AOI211_X1 U19915 ( .C1(n16824), .C2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16732), .B(n16731), .ZN(n16733) );
  OAI211_X1 U19916 ( .C1(n18705), .C2(n16735), .A(n16734), .B(n16733), .ZN(
        P3_U2659) );
  AOI22_X1 U19917 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n16824), .B1(
        n16843), .B2(P3_EBX_REG_11__SCAN_IN), .ZN(n16746) );
  OAI21_X1 U19918 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16747), .A(
        n17647), .ZN(n16736) );
  INV_X1 U19919 ( .A(n16736), .ZN(n17677) );
  OAI21_X1 U19920 ( .B1(n16738), .B2(n16737), .A(n16531), .ZN(n16739) );
  XNOR2_X1 U19921 ( .A(n17677), .B(n16739), .ZN(n16742) );
  NOR2_X1 U19922 ( .A1(n16868), .A2(n16750), .ZN(n16749) );
  INV_X1 U19923 ( .A(n16749), .ZN(n16766) );
  OAI21_X1 U19924 ( .B1(n16751), .B2(n16766), .A(n18703), .ZN(n16740) );
  AOI22_X1 U19925 ( .A1(n18661), .A2(n16742), .B1(n16741), .B2(n16740), .ZN(
        n16745) );
  OAI211_X1 U19926 ( .C1(n16748), .C2(n17118), .A(n16845), .B(n16743), .ZN(
        n16744) );
  NAND4_X1 U19927 ( .A1(n16746), .A2(n16745), .A3(n18094), .A4(n16744), .ZN(
        P3_U2660) );
  INV_X1 U19928 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17685) );
  AND3_X1 U19929 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17714), .A3(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16783) );
  NAND2_X1 U19930 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16783), .ZN(
        n16772) );
  INV_X1 U19931 ( .A(n16772), .ZN(n16763) );
  NAND2_X1 U19932 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16763), .ZN(
        n16759) );
  AOI21_X1 U19933 ( .B1(n17685), .B2(n16759), .A(n16747), .ZN(n17688) );
  OAI21_X1 U19934 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16759), .A(
        n16531), .ZN(n16764) );
  XOR2_X1 U19935 ( .A(n17688), .B(n16764), .Z(n16757) );
  AOI211_X1 U19936 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16760), .A(n16748), .B(
        n16874), .ZN(n16755) );
  AOI21_X1 U19937 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n16749), .A(
        P3_REIP_REG_10__SCAN_IN), .ZN(n16753) );
  OR2_X1 U19938 ( .A1(n16750), .A2(n16877), .ZN(n16758) );
  OAI21_X1 U19939 ( .B1(n16751), .B2(n16758), .A(n16880), .ZN(n16752) );
  OAI22_X1 U19940 ( .A1(n16753), .A2(n16752), .B1(n17685), .B2(n16865), .ZN(
        n16754) );
  AOI211_X1 U19941 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16843), .A(n16755), .B(
        n16754), .ZN(n16756) );
  OAI211_X1 U19942 ( .C1(n16757), .C2(n16839), .A(n16756), .B(n18094), .ZN(
        P3_U2661) );
  INV_X1 U19943 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18699) );
  NAND2_X1 U19944 ( .A1(n16880), .A2(n16758), .ZN(n16774) );
  OAI21_X1 U19945 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16763), .A(
        n16759), .ZN(n17703) );
  NOR2_X1 U19946 ( .A1(n16839), .A2(n16531), .ZN(n16785) );
  INV_X1 U19947 ( .A(n16785), .ZN(n16864) );
  OAI22_X1 U19948 ( .A1(n16875), .A2(n17056), .B1(n17703), .B2(n16864), .ZN(
        n16769) );
  INV_X1 U19949 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16762) );
  OAI211_X1 U19950 ( .C1(n16771), .C2(n17056), .A(n16845), .B(n16760), .ZN(
        n16761) );
  OAI21_X1 U19951 ( .B1(n16865), .B2(n16762), .A(n16761), .ZN(n16768) );
  INV_X1 U19952 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16876) );
  OAI221_X1 U19953 ( .B1(n17703), .B2(n16763), .C1(n17703), .C2(n16876), .A(
        n18661), .ZN(n16765) );
  OAI22_X1 U19954 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16766), .B1(n16765), 
        .B2(n16764), .ZN(n16767) );
  NOR4_X1 U19955 ( .A1(n9846), .A2(n16769), .A3(n16768), .A4(n16767), .ZN(
        n16770) );
  OAI21_X1 U19956 ( .B1(n18699), .B2(n16774), .A(n16770), .ZN(P3_U2662) );
  INV_X1 U19957 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n16781) );
  AOI211_X1 U19958 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16791), .A(n16771), .B(
        n16874), .ZN(n16778) );
  AOI21_X1 U19959 ( .B1(n16783), .B2(n16876), .A(n16837), .ZN(n16786) );
  OAI21_X1 U19960 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16783), .A(
        n16772), .ZN(n17718) );
  OAI21_X1 U19961 ( .B1(n16786), .B2(n17718), .A(n18094), .ZN(n16773) );
  AOI21_X1 U19962 ( .B1(n16786), .B2(n17718), .A(n16773), .ZN(n16775) );
  INV_X1 U19963 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18698) );
  OAI22_X1 U19964 ( .A1(n16776), .A2(n16775), .B1(n18698), .B2(n16774), .ZN(
        n16777) );
  AOI211_X1 U19965 ( .C1(n16824), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16778), .B(n16777), .ZN(n16780) );
  NAND4_X1 U19966 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n16833), .A3(n16782), 
        .A4(n18698), .ZN(n16779) );
  OAI211_X1 U19967 ( .C1(n16781), .C2(n16875), .A(n16780), .B(n16779), .ZN(
        P3_U2663) );
  NAND2_X1 U19968 ( .A1(n16833), .A2(n16782), .ZN(n16789) );
  INV_X1 U19969 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n20777) );
  AOI221_X1 U19970 ( .B1(n18694), .B2(n16833), .C1(n16797), .C2(n16833), .A(
        n16877), .ZN(n16788) );
  NAND2_X1 U19971 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17714), .ZN(
        n16799) );
  AOI21_X1 U19972 ( .B1(n17730), .B2(n16799), .A(n16783), .ZN(n17735) );
  NAND2_X1 U19973 ( .A1(n17714), .A2(n16861), .ZN(n16800) );
  AOI21_X1 U19974 ( .B1(n17735), .B2(n16800), .A(n16839), .ZN(n16784) );
  OAI22_X1 U19975 ( .A1(n17735), .A2(n16786), .B1(n16785), .B2(n16784), .ZN(
        n16787) );
  OAI221_X1 U19976 ( .B1(P3_REIP_REG_7__SCAN_IN), .B2(n16789), .C1(n20777), 
        .C2(n16788), .A(n16787), .ZN(n16790) );
  AOI211_X1 U19977 ( .C1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n16824), .A(
        n9846), .B(n16790), .ZN(n16793) );
  OAI211_X1 U19978 ( .C1(n16795), .C2(n16794), .A(n16845), .B(n16791), .ZN(
        n16792) );
  OAI211_X1 U19979 ( .C1(n16794), .C2(n16875), .A(n16793), .B(n16792), .ZN(
        P3_U2664) );
  AOI21_X1 U19980 ( .B1(n16833), .B2(n16797), .A(n16877), .ZN(n16818) );
  AOI211_X1 U19981 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16811), .A(n16795), .B(
        n16874), .ZN(n16796) );
  AOI21_X1 U19982 ( .B1(n16824), .B2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16796), .ZN(n16807) );
  NOR3_X1 U19983 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16868), .A3(n16797), .ZN(
        n16805) );
  INV_X1 U19984 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16810) );
  NAND2_X1 U19985 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16798), .ZN(
        n16825) );
  NOR2_X1 U19986 ( .A1(n16810), .A2(n16825), .ZN(n16809) );
  OAI21_X1 U19987 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16809), .A(
        n16799), .ZN(n17744) );
  NAND2_X1 U19988 ( .A1(n17744), .A2(n16800), .ZN(n16803) );
  INV_X1 U19989 ( .A(n17744), .ZN(n16801) );
  OAI211_X1 U19990 ( .C1(n16809), .C2(n16837), .A(n16801), .B(n16870), .ZN(
        n16802) );
  OAI211_X1 U19991 ( .C1(n16866), .C2(n16803), .A(n18094), .B(n16802), .ZN(
        n16804) );
  AOI211_X1 U19992 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16843), .A(n16805), .B(
        n16804), .ZN(n16806) );
  OAI211_X1 U19993 ( .C1(n18694), .C2(n16818), .A(n16807), .B(n16806), .ZN(
        P3_U2665) );
  AOI21_X1 U19994 ( .B1(n16833), .B2(n16808), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n16819) );
  AOI22_X1 U19995 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n16824), .B1(
        n16843), .B2(P3_EBX_REG_5__SCAN_IN), .ZN(n16817) );
  AOI21_X1 U19996 ( .B1(n16810), .B2(n16825), .A(n16809), .ZN(n17759) );
  AOI21_X1 U19997 ( .B1(n16798), .B2(n16861), .A(n16837), .ZN(n16826) );
  XOR2_X1 U19998 ( .A(n17759), .B(n16826), .Z(n16815) );
  OAI211_X1 U19999 ( .C1(n16812), .C2(n16820), .A(n16811), .B(n16845), .ZN(
        n16813) );
  INV_X1 U20000 ( .A(n16813), .ZN(n16814) );
  AOI211_X1 U20001 ( .C1(n18661), .C2(n16815), .A(n9846), .B(n16814), .ZN(
        n16816) );
  OAI211_X1 U20002 ( .C1(n16819), .C2(n16818), .A(n16817), .B(n16816), .ZN(
        P3_U2666) );
  AOI21_X1 U20003 ( .B1(n16833), .B2(n16832), .A(n16877), .ZN(n16840) );
  AOI211_X1 U20004 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16844), .A(n16820), .B(
        n16874), .ZN(n16823) );
  NOR2_X1 U20005 ( .A1(n18161), .A2(n18810), .ZN(n18825) );
  INV_X1 U20006 ( .A(n18825), .ZN(n16882) );
  OAI221_X1 U20007 ( .B1(n16882), .B2(n9593), .C1(n16882), .C2(n16821), .A(
        n18094), .ZN(n16822) );
  AOI211_X1 U20008 ( .C1(n16824), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n16823), .B(n16822), .ZN(n16831) );
  NOR2_X1 U20009 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17761), .ZN(
        n17773) );
  NOR2_X1 U20010 ( .A1(n17804), .A2(n17761), .ZN(n16836) );
  OAI21_X1 U20011 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16836), .A(
        n16825), .ZN(n17770) );
  AOI22_X1 U20012 ( .A1(n16861), .A2(n17773), .B1(n16826), .B2(n17770), .ZN(
        n16827) );
  AOI221_X1 U20013 ( .B1(n16531), .B2(n16827), .C1(n17770), .C2(n16827), .A(
        n16839), .ZN(n16829) );
  NOR3_X1 U20014 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16868), .A3(n16832), .ZN(
        n16828) );
  AOI211_X1 U20015 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16843), .A(n16829), .B(
        n16828), .ZN(n16830) );
  OAI211_X1 U20016 ( .C1(n16840), .C2(n18690), .A(n16831), .B(n16830), .ZN(
        P3_U2667) );
  INV_X1 U20017 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16849) );
  INV_X1 U20018 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18686) );
  NOR2_X1 U20019 ( .A1(n18685), .A2(n18686), .ZN(n16851) );
  INV_X1 U20020 ( .A(n16851), .ZN(n16835) );
  NAND2_X1 U20021 ( .A1(n16833), .A2(n16832), .ZN(n16834) );
  NOR2_X1 U20022 ( .A1(n18784), .A2(n18612), .ZN(n18610) );
  OAI21_X1 U20023 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18610), .A(
        n9593), .ZN(n18754) );
  OAI22_X1 U20024 ( .A1(n16835), .A2(n16834), .B1(n16882), .B2(n18754), .ZN(
        n16842) );
  INV_X1 U20025 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18688) );
  NAND2_X1 U20026 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16850) );
  AOI21_X1 U20027 ( .B1(n16849), .B2(n16850), .A(n16836), .ZN(n17786) );
  AOI21_X1 U20028 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n16861), .A(
        n16837), .ZN(n16860) );
  XNOR2_X1 U20029 ( .A(n17786), .B(n16860), .ZN(n16838) );
  OAI22_X1 U20030 ( .A1(n16840), .A2(n18688), .B1(n16839), .B2(n16838), .ZN(
        n16841) );
  AOI211_X1 U20031 ( .C1(n16843), .C2(P3_EBX_REG_3__SCAN_IN), .A(n16842), .B(
        n16841), .ZN(n16848) );
  OAI211_X1 U20032 ( .C1(n16852), .C2(n16846), .A(n16845), .B(n16844), .ZN(
        n16847) );
  OAI211_X1 U20033 ( .C1(n16865), .C2(n16849), .A(n16848), .B(n16847), .ZN(
        P3_U2668) );
  OAI21_X1 U20034 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16850), .ZN(n17794) );
  AOI211_X1 U20035 ( .C1(n18685), .C2(n18686), .A(n16851), .B(n16868), .ZN(
        n16859) );
  NAND2_X1 U20036 ( .A1(n20773), .A2(n17189), .ZN(n16853) );
  AOI211_X1 U20037 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16853), .A(n16852), .B(
        n16874), .ZN(n16858) );
  INV_X1 U20038 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17797) );
  OAI22_X1 U20039 ( .A1(n17797), .A2(n16865), .B1(n16875), .B2(n16854), .ZN(
        n16857) );
  NOR2_X1 U20040 ( .A1(n18784), .A2(n18778), .ZN(n18630) );
  NOR2_X1 U20041 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18630), .ZN(
        n18614) );
  INV_X1 U20042 ( .A(n18614), .ZN(n18608) );
  OAI21_X1 U20043 ( .B1(n18612), .B2(n18784), .A(n18608), .ZN(n18764) );
  OAI22_X1 U20044 ( .A1(n18686), .A2(n16855), .B1(n18764), .B2(n16882), .ZN(
        n16856) );
  NOR4_X1 U20045 ( .A1(n16859), .A2(n16858), .A3(n16857), .A4(n16856), .ZN(
        n16863) );
  OAI211_X1 U20046 ( .C1(n16861), .C2(n17794), .A(n18661), .B(n16860), .ZN(
        n16862) );
  OAI211_X1 U20047 ( .C1(n16864), .C2(n17794), .A(n16863), .B(n16862), .ZN(
        P3_U2669) );
  AOI22_X1 U20048 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(n18778), .B2(n18784), .ZN(
        n18775) );
  AOI22_X1 U20049 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16877), .B1(n18775), 
        .B2(n18825), .ZN(n16873) );
  OAI211_X1 U20050 ( .C1(n16876), .C2(n16866), .A(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B(n16865), .ZN(n16871) );
  OAI21_X1 U20051 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n16867), .ZN(n17191) );
  OAI22_X1 U20052 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16868), .B1(n16874), 
        .B2(n17191), .ZN(n16869) );
  AOI221_X1 U20053 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16871), .C1(
        n16870), .C2(n16871), .A(n16869), .ZN(n16872) );
  OAI211_X1 U20054 ( .C1(n16875), .C2(n17189), .A(n16873), .B(n16872), .ZN(
        P3_U2670) );
  AOI21_X1 U20055 ( .B1(n16875), .B2(n16874), .A(n20773), .ZN(n16879) );
  NOR3_X1 U20056 ( .A1(n18821), .A2(n16877), .A3(n16876), .ZN(n16878) );
  AOI211_X1 U20057 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(n16880), .A(n16879), .B(
        n16878), .ZN(n16881) );
  OAI21_X1 U20058 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n16882), .A(
        n16881), .ZN(P3_U2671) );
  NOR2_X1 U20059 ( .A1(n16884), .A2(n16883), .ZN(n16890) );
  NOR2_X1 U20060 ( .A1(n16885), .A2(n17003), .ZN(n16975) );
  INV_X1 U20061 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n16931) );
  NAND2_X1 U20062 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .ZN(n16886) );
  NOR4_X1 U20063 ( .A1(n16888), .A2(n16931), .A3(n16887), .A4(n16886), .ZN(
        n16889) );
  NAND4_X1 U20064 ( .A1(n16890), .A2(n16924), .A3(n16975), .A4(n16889), .ZN(
        n16893) );
  NOR2_X1 U20065 ( .A1(n16894), .A2(n16893), .ZN(n16919) );
  NAND2_X1 U20066 ( .A1(n17188), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16892) );
  NAND2_X1 U20067 ( .A1(n16919), .A2(n17120), .ZN(n16891) );
  OAI22_X1 U20068 ( .A1(n16919), .A2(n16892), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16891), .ZN(P3_U2672) );
  NAND2_X1 U20069 ( .A1(n16894), .A2(n16893), .ZN(n16895) );
  NAND2_X1 U20070 ( .A1(n16895), .A2(n17188), .ZN(n16918) );
  AOI22_X1 U20071 ( .A1(n17018), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17079), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16899) );
  AOI22_X1 U20072 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16898) );
  AOI22_X1 U20073 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16897) );
  AOI22_X1 U20074 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16896) );
  NAND4_X1 U20075 ( .A1(n16899), .A2(n16898), .A3(n16897), .A4(n16896), .ZN(
        n16906) );
  AOI22_X1 U20076 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10140), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16904) );
  AOI22_X1 U20077 ( .A1(n10280), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16903) );
  INV_X1 U20078 ( .A(n16900), .ZN(n17166) );
  AOI22_X1 U20079 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16902) );
  AOI22_X1 U20080 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16901) );
  NAND4_X1 U20081 ( .A1(n16904), .A2(n16903), .A3(n16902), .A4(n16901), .ZN(
        n16905) );
  NOR2_X1 U20082 ( .A1(n16906), .A2(n16905), .ZN(n16917) );
  AOI22_X1 U20083 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16916) );
  AOI22_X1 U20084 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10140), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16915) );
  AOI22_X1 U20085 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16907) );
  OAI21_X1 U20086 ( .B1(n16983), .B2(n20713), .A(n16907), .ZN(n16913) );
  AOI22_X1 U20087 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16911) );
  AOI22_X1 U20088 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17018), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16910) );
  AOI22_X1 U20089 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16909) );
  AOI22_X1 U20090 ( .A1(n14241), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16908) );
  NAND4_X1 U20091 ( .A1(n16911), .A2(n16910), .A3(n16909), .A4(n16908), .ZN(
        n16912) );
  AOI211_X1 U20092 ( .C1(n17079), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n16913), .B(n16912), .ZN(n16914) );
  NAND3_X1 U20093 ( .A1(n16916), .A2(n16915), .A3(n16914), .ZN(n16921) );
  NAND2_X1 U20094 ( .A1(n16922), .A2(n16921), .ZN(n16920) );
  XNOR2_X1 U20095 ( .A(n16917), .B(n16920), .ZN(n17208) );
  OAI22_X1 U20096 ( .A1(n16919), .A2(n16918), .B1(n17208), .B2(n17188), .ZN(
        P3_U2673) );
  OAI21_X1 U20097 ( .B1(n16922), .B2(n16921), .A(n16920), .ZN(n17212) );
  NOR2_X1 U20098 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16935), .ZN(n16923) );
  AOI22_X1 U20099 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16925), .B1(n16924), 
        .B2(n16923), .ZN(n16926) );
  OAI21_X1 U20100 ( .B1(n17212), .B2(n17188), .A(n16926), .ZN(P3_U2674) );
  OAI21_X1 U20101 ( .B1(n16932), .B2(n16928), .A(n16927), .ZN(n17221) );
  NAND3_X1 U20102 ( .A1(n16935), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17188), 
        .ZN(n16929) );
  OAI221_X1 U20103 ( .B1(n16935), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17188), 
        .C2(n17221), .A(n16929), .ZN(P3_U2676) );
  OAI21_X1 U20104 ( .B1(n16931), .B2(n17193), .A(n16930), .ZN(n16934) );
  AOI21_X1 U20105 ( .B1(n16933), .B2(n16937), .A(n16932), .ZN(n17222) );
  AOI22_X1 U20106 ( .A1(n16935), .A2(n16934), .B1(n17222), .B2(n17193), .ZN(
        n16936) );
  INV_X1 U20107 ( .A(n16936), .ZN(P3_U2677) );
  AOI21_X1 U20108 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17188), .A(n16945), .ZN(
        n16939) );
  OAI21_X1 U20109 ( .B1(n16941), .B2(n16938), .A(n16937), .ZN(n17231) );
  OAI22_X1 U20110 ( .A1(n16940), .A2(n16939), .B1(n17188), .B2(n17231), .ZN(
        P3_U2678) );
  INV_X1 U20111 ( .A(n16950), .ZN(n16964) );
  AOI22_X1 U20112 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17188), .B1(
        P3_EBX_REG_23__SCAN_IN), .B2(n16964), .ZN(n16944) );
  AOI21_X1 U20113 ( .B1(n16942), .B2(n16946), .A(n16941), .ZN(n17232) );
  INV_X1 U20114 ( .A(n17232), .ZN(n16943) );
  OAI22_X1 U20115 ( .A1(n16945), .A2(n16944), .B1(n17188), .B2(n16943), .ZN(
        P3_U2679) );
  OAI21_X1 U20116 ( .B1(n16948), .B2(n16947), .A(n16946), .ZN(n17242) );
  NAND3_X1 U20117 ( .A1(n16950), .A2(P3_EBX_REG_23__SCAN_IN), .A3(n17188), 
        .ZN(n16949) );
  OAI221_X1 U20118 ( .B1(n16950), .B2(P3_EBX_REG_23__SCAN_IN), .C1(n17188), 
        .C2(n17242), .A(n16949), .ZN(P3_U2680) );
  AOI22_X1 U20119 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17188), .B1(
        P3_EBX_REG_21__SCAN_IN), .B2(n16977), .ZN(n16963) );
  AOI22_X1 U20120 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16961) );
  AOI22_X1 U20121 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17018), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16960) );
  AOI22_X1 U20122 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16951) );
  OAI21_X1 U20123 ( .B1(n16952), .B2(n20713), .A(n16951), .ZN(n16958) );
  AOI22_X1 U20124 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(n9591), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16956) );
  AOI22_X1 U20125 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16955) );
  AOI22_X1 U20126 ( .A1(n14241), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17079), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16954) );
  AOI22_X1 U20127 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16953) );
  NAND4_X1 U20128 ( .A1(n16956), .A2(n16955), .A3(n16954), .A4(n16953), .ZN(
        n16957) );
  AOI211_X1 U20129 ( .C1(n17166), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n16958), .B(n16957), .ZN(n16959) );
  NAND3_X1 U20130 ( .A1(n16961), .A2(n16960), .A3(n16959), .ZN(n17244) );
  INV_X1 U20131 ( .A(n17244), .ZN(n16962) );
  OAI22_X1 U20132 ( .A1(n16964), .A2(n16963), .B1(n16962), .B2(n17188), .ZN(
        P3_U2681) );
  AOI22_X1 U20133 ( .A1(n17080), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16968) );
  AOI22_X1 U20134 ( .A1(n14241), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10140), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16967) );
  AOI22_X1 U20135 ( .A1(n17018), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17079), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16966) );
  AOI22_X1 U20136 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16965) );
  NAND4_X1 U20137 ( .A1(n16968), .A2(n16967), .A3(n16966), .A4(n16965), .ZN(
        n16974) );
  AOI22_X1 U20138 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16972) );
  AOI22_X1 U20139 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16971) );
  AOI22_X1 U20140 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16970) );
  AOI22_X1 U20141 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16969) );
  NAND4_X1 U20142 ( .A1(n16972), .A2(n16971), .A3(n16970), .A4(n16969), .ZN(
        n16973) );
  NOR2_X1 U20143 ( .A1(n16974), .A2(n16973), .ZN(n17250) );
  NOR2_X1 U20144 ( .A1(n17193), .A2(n16975), .ZN(n16990) );
  AOI22_X1 U20145 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16990), .B1(n16977), 
        .B2(n16976), .ZN(n16978) );
  OAI21_X1 U20146 ( .B1(n17250), .B2(n17188), .A(n16978), .ZN(P3_U2682) );
  AOI22_X1 U20147 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16982) );
  AOI22_X1 U20148 ( .A1(n10153), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10152), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16981) );
  AOI22_X1 U20149 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16980) );
  AOI22_X1 U20150 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16979) );
  NAND4_X1 U20151 ( .A1(n16982), .A2(n16981), .A3(n16980), .A4(n16979), .ZN(
        n16989) );
  AOI22_X1 U20152 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16987) );
  AOI22_X1 U20153 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16986) );
  AOI22_X1 U20154 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10099), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16985) );
  AOI22_X1 U20155 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10140), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16984) );
  NAND4_X1 U20156 ( .A1(n16987), .A2(n16986), .A3(n16985), .A4(n16984), .ZN(
        n16988) );
  NOR2_X1 U20157 ( .A1(n16989), .A2(n16988), .ZN(n17258) );
  OAI21_X1 U20158 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16991), .A(n16990), .ZN(
        n16992) );
  OAI21_X1 U20159 ( .B1(n17258), .B2(n17188), .A(n16992), .ZN(P3_U2683) );
  AOI22_X1 U20160 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10152), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16996) );
  AOI22_X1 U20161 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16995) );
  AOI22_X1 U20162 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16994) );
  AOI22_X1 U20163 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16993) );
  NAND4_X1 U20164 ( .A1(n16996), .A2(n16995), .A3(n16994), .A4(n16993), .ZN(
        n17002) );
  AOI22_X1 U20165 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17079), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17000) );
  AOI22_X1 U20166 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16999) );
  AOI22_X1 U20167 ( .A1(n17018), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16998) );
  AOI22_X1 U20168 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10140), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16997) );
  NAND4_X1 U20169 ( .A1(n17000), .A2(n16999), .A3(n16998), .A4(n16997), .ZN(
        n17001) );
  NOR2_X1 U20170 ( .A1(n17002), .A2(n17001), .ZN(n17262) );
  OAI21_X1 U20171 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17017), .A(n17003), .ZN(
        n17004) );
  AOI22_X1 U20172 ( .A1(n17193), .A2(n17262), .B1(n17004), .B2(n17188), .ZN(
        P3_U2684) );
  AOI21_X1 U20173 ( .B1(n20688), .B2(n17029), .A(n17193), .ZN(n17005) );
  INV_X1 U20174 ( .A(n17005), .ZN(n17016) );
  AOI22_X1 U20175 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17009) );
  AOI22_X1 U20176 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10099), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17008) );
  AOI22_X1 U20177 ( .A1(n17080), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10152), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17007) );
  AOI22_X1 U20178 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17006) );
  NAND4_X1 U20179 ( .A1(n17009), .A2(n17008), .A3(n17007), .A4(n17006), .ZN(
        n17015) );
  AOI22_X1 U20180 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10140), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17013) );
  AOI22_X1 U20181 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17012) );
  AOI22_X1 U20182 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17018), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17011) );
  AOI22_X1 U20183 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17010) );
  NAND4_X1 U20184 ( .A1(n17013), .A2(n17012), .A3(n17011), .A4(n17010), .ZN(
        n17014) );
  NOR2_X1 U20185 ( .A1(n17015), .A2(n17014), .ZN(n17267) );
  OAI22_X1 U20186 ( .A1(n17017), .A2(n17016), .B1(n17267), .B2(n17188), .ZN(
        P3_U2685) );
  AOI22_X1 U20187 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17018), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17022) );
  AOI22_X1 U20188 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n9591), .ZN(n17021) );
  AOI22_X1 U20189 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n10141), .ZN(n17020) );
  AOI22_X1 U20190 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n9595), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17019) );
  NAND4_X1 U20191 ( .A1(n17022), .A2(n17021), .A3(n17020), .A4(n17019), .ZN(
        n17028) );
  AOI22_X1 U20192 ( .A1(n14241), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17026) );
  AOI22_X1 U20193 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17079), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17025) );
  AOI22_X1 U20194 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17153), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n17156), .ZN(n17024) );
  AOI22_X1 U20195 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n10280), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17151), .ZN(n17023) );
  NAND4_X1 U20196 ( .A1(n17026), .A2(n17025), .A3(n17024), .A4(n17023), .ZN(
        n17027) );
  NOR2_X1 U20197 ( .A1(n17028), .A2(n17027), .ZN(n17272) );
  OAI21_X1 U20198 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17045), .A(n17029), .ZN(
        n17030) );
  AOI22_X1 U20199 ( .A1(n17193), .A2(n17272), .B1(n17030), .B2(n17188), .ZN(
        P3_U2686) );
  OAI21_X1 U20200 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17031), .A(n17188), .ZN(
        n17044) );
  AOI22_X1 U20201 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17035) );
  AOI22_X1 U20202 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17034) );
  AOI22_X1 U20203 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17033) );
  AOI22_X1 U20204 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17032) );
  NAND4_X1 U20205 ( .A1(n17035), .A2(n17034), .A3(n17033), .A4(n17032), .ZN(
        n17043) );
  AOI22_X1 U20206 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17041) );
  AOI22_X1 U20207 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17040) );
  AOI22_X1 U20208 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10152), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17039) );
  AOI22_X1 U20209 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17140), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17038) );
  NAND4_X1 U20210 ( .A1(n17041), .A2(n17040), .A3(n17039), .A4(n17038), .ZN(
        n17042) );
  NOR2_X1 U20211 ( .A1(n17043), .A2(n17042), .ZN(n17279) );
  OAI22_X1 U20212 ( .A1(n17045), .A2(n17044), .B1(n17279), .B2(n17188), .ZN(
        P3_U2687) );
  AOI22_X1 U20213 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17049) );
  AOI22_X1 U20214 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17048) );
  AOI22_X1 U20215 ( .A1(n10153), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17047) );
  AOI22_X1 U20216 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17046) );
  NAND4_X1 U20217 ( .A1(n17049), .A2(n17048), .A3(n17047), .A4(n17046), .ZN(
        n17055) );
  AOI22_X1 U20218 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17053) );
  AOI22_X1 U20219 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17052) );
  AOI22_X1 U20220 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17051) );
  AOI22_X1 U20221 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10099), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17050) );
  NAND4_X1 U20222 ( .A1(n17053), .A2(n17052), .A3(n17051), .A4(n17050), .ZN(
        n17054) );
  NOR2_X1 U20223 ( .A1(n17055), .A2(n17054), .ZN(n17285) );
  INV_X1 U20224 ( .A(n17071), .ZN(n17058) );
  NAND2_X1 U20225 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17171), .ZN(n17170) );
  NAND2_X1 U20226 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17121), .ZN(n17117) );
  NOR2_X1 U20227 ( .A1(n17118), .A2(n17117), .ZN(n17101) );
  OAI221_X1 U20228 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17058), .C1(
        P3_EBX_REG_15__SCAN_IN), .C2(n17101), .A(n17057), .ZN(n17059) );
  AOI22_X1 U20229 ( .A1(n17193), .A2(n17285), .B1(n17059), .B2(n17188), .ZN(
        P3_U2688) );
  AOI22_X1 U20230 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n9591), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17069) );
  AOI22_X1 U20231 ( .A1(n14241), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17068) );
  AOI22_X1 U20232 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17060) );
  OAI21_X1 U20233 ( .B1(n10089), .B2(n20713), .A(n17060), .ZN(n17066) );
  AOI22_X1 U20234 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10280), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17064) );
  AOI22_X1 U20235 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17063) );
  AOI22_X1 U20236 ( .A1(n17018), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17079), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17062) );
  AOI22_X1 U20237 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17061) );
  NAND4_X1 U20238 ( .A1(n17064), .A2(n17063), .A3(n17062), .A4(n17061), .ZN(
        n17065) );
  AOI211_X1 U20239 ( .C1(n17157), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n17066), .B(n17065), .ZN(n17067) );
  NAND3_X1 U20240 ( .A1(n17069), .A2(n17068), .A3(n17067), .ZN(n17287) );
  INV_X1 U20241 ( .A(n17287), .ZN(n17074) );
  INV_X1 U20242 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17102) );
  NAND2_X1 U20243 ( .A1(n17120), .A2(n17101), .ZN(n17088) );
  NOR3_X1 U20244 ( .A1(n17070), .A2(n17102), .A3(n17088), .ZN(n17090) );
  AOI21_X1 U20245 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17188), .A(n17090), .ZN(
        n17073) );
  NOR2_X1 U20246 ( .A1(n17071), .A2(n17088), .ZN(n17072) );
  OAI22_X1 U20247 ( .A1(n17074), .A2(n17188), .B1(n17073), .B2(n17072), .ZN(
        P3_U2689) );
  AOI22_X1 U20248 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17078) );
  AOI22_X1 U20249 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17077) );
  AOI22_X1 U20250 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10280), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17076) );
  AOI22_X1 U20251 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17075) );
  NAND4_X1 U20252 ( .A1(n17078), .A2(n17077), .A3(n17076), .A4(n17075), .ZN(
        n17087) );
  AOI22_X1 U20253 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17079), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17085) );
  AOI22_X1 U20254 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17084) );
  AOI22_X1 U20255 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17083) );
  AOI22_X1 U20256 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17082) );
  NAND4_X1 U20257 ( .A1(n17085), .A2(n17084), .A3(n17083), .A4(n17082), .ZN(
        n17086) );
  NOR2_X1 U20258 ( .A1(n17087), .A2(n17086), .ZN(n17291) );
  INV_X1 U20259 ( .A(n17088), .ZN(n17103) );
  AOI22_X1 U20260 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17188), .B1(
        P3_EBX_REG_12__SCAN_IN), .B2(n17103), .ZN(n17089) );
  OAI22_X1 U20261 ( .A1(n17291), .A2(n17188), .B1(n17090), .B2(n17089), .ZN(
        P3_U2690) );
  AOI22_X1 U20262 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17079), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17094) );
  AOI22_X1 U20263 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17093) );
  AOI22_X1 U20264 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17153), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17092) );
  AOI22_X1 U20265 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10141), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17091) );
  NAND4_X1 U20266 ( .A1(n17094), .A2(n17093), .A3(n17092), .A4(n17091), .ZN(
        n17100) );
  AOI22_X1 U20267 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17098) );
  AOI22_X1 U20268 ( .A1(n17018), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17097) );
  AOI22_X1 U20269 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n9591), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17096) );
  AOI22_X1 U20270 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10280), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17095) );
  NAND4_X1 U20271 ( .A1(n17098), .A2(n17097), .A3(n17096), .A4(n17095), .ZN(
        n17099) );
  NOR2_X1 U20272 ( .A1(n17100), .A2(n17099), .ZN(n17295) );
  NOR2_X1 U20273 ( .A1(n17193), .A2(n17101), .ZN(n17105) );
  AOI22_X1 U20274 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17105), .B1(n17103), 
        .B2(n17102), .ZN(n17104) );
  OAI21_X1 U20275 ( .B1(n17295), .B2(n17188), .A(n17104), .ZN(P3_U2691) );
  INV_X1 U20276 ( .A(n17105), .ZN(n17119) );
  AOI22_X1 U20277 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17115) );
  AOI22_X1 U20278 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17114) );
  AOI22_X1 U20279 ( .A1(n14241), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17106) );
  OAI21_X1 U20280 ( .B1(n17155), .B2(n18182), .A(n17106), .ZN(n17112) );
  AOI22_X1 U20281 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17153), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17110) );
  AOI22_X1 U20282 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17109) );
  AOI22_X1 U20283 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17108) );
  AOI22_X1 U20284 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17107) );
  NAND4_X1 U20285 ( .A1(n17110), .A2(n17109), .A3(n17108), .A4(n17107), .ZN(
        n17111) );
  AOI211_X1 U20286 ( .C1(n17140), .C2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n17112), .B(n17111), .ZN(n17113) );
  NAND3_X1 U20287 ( .A1(n17115), .A2(n17114), .A3(n17113), .ZN(n17298) );
  NAND2_X1 U20288 ( .A1(n17193), .A2(n17298), .ZN(n17116) );
  OAI221_X1 U20289 ( .B1(n17119), .B2(n17118), .C1(n17119), .C2(n17117), .A(
        n17116), .ZN(P3_U2692) );
  NAND2_X1 U20290 ( .A1(n17120), .A2(n17121), .ZN(n17135) );
  NOR2_X1 U20291 ( .A1(n17193), .A2(n17121), .ZN(n17147) );
  AOI22_X1 U20292 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17133) );
  AOI22_X1 U20293 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17132) );
  AOI22_X1 U20294 ( .A1(n17018), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17122) );
  OAI21_X1 U20295 ( .B1(n17155), .B2(n18176), .A(n17122), .ZN(n17130) );
  AOI22_X1 U20296 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17128) );
  AOI22_X1 U20297 ( .A1(n14241), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17153), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17127) );
  AOI22_X1 U20298 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17126) );
  AOI22_X1 U20299 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17125) );
  NAND4_X1 U20300 ( .A1(n17128), .A2(n17127), .A3(n17126), .A4(n17125), .ZN(
        n17129) );
  AOI211_X1 U20301 ( .C1(n17157), .C2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n17130), .B(n17129), .ZN(n17131) );
  NAND3_X1 U20302 ( .A1(n17133), .A2(n17132), .A3(n17131), .ZN(n17301) );
  AOI22_X1 U20303 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17147), .B1(n17193), 
        .B2(n17301), .ZN(n17134) );
  OAI21_X1 U20304 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17135), .A(n17134), .ZN(
        P3_U2693) );
  AOI22_X1 U20305 ( .A1(n14241), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n17159), .ZN(n17139) );
  AOI22_X1 U20306 ( .A1(n14285), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17138) );
  AOI22_X1 U20307 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17166), .B1(
        n10280), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17137) );
  AOI22_X1 U20308 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10141), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17156), .ZN(n17136) );
  NAND4_X1 U20309 ( .A1(n17139), .A2(n17138), .A3(n17137), .A4(n17136), .ZN(
        n17146) );
  AOI22_X1 U20310 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17123), .B1(
        n17140), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17144) );
  AOI22_X1 U20311 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17153), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17143) );
  AOI22_X1 U20312 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17079), .B1(
        n17081), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17142) );
  AOI22_X1 U20313 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17151), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n9591), .ZN(n17141) );
  NAND4_X1 U20314 ( .A1(n17144), .A2(n17143), .A3(n17142), .A4(n17141), .ZN(
        n17145) );
  NOR2_X1 U20315 ( .A1(n17146), .A2(n17145), .ZN(n17305) );
  INV_X1 U20316 ( .A(n17170), .ZN(n17148) );
  OAI21_X1 U20317 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17148), .A(n17147), .ZN(
        n17149) );
  OAI21_X1 U20318 ( .B1(n17305), .B2(n17188), .A(n17149), .ZN(P3_U2694) );
  AOI22_X1 U20319 ( .A1(n10153), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17169) );
  AOI22_X1 U20320 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17168) );
  AOI22_X1 U20321 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10140), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17154) );
  OAI21_X1 U20322 ( .B1(n17155), .B2(n18164), .A(n17154), .ZN(n17165) );
  AOI22_X1 U20323 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17163) );
  AOI22_X1 U20324 ( .A1(n17081), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17162) );
  AOI22_X1 U20325 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17161) );
  AOI22_X1 U20326 ( .A1(n17079), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17160) );
  NAND4_X1 U20327 ( .A1(n17163), .A2(n17162), .A3(n17161), .A4(n17160), .ZN(
        n17164) );
  AOI211_X1 U20328 ( .C1(n17166), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n17165), .B(n17164), .ZN(n17167) );
  NAND3_X1 U20329 ( .A1(n17169), .A2(n17168), .A3(n17167), .ZN(n17308) );
  INV_X1 U20330 ( .A(n17308), .ZN(n17173) );
  OAI21_X1 U20331 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17171), .A(n17170), .ZN(
        n17172) );
  AOI22_X1 U20332 ( .A1(n17193), .A2(n17173), .B1(n17172), .B2(n17188), .ZN(
        P3_U2695) );
  NAND2_X1 U20333 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17174), .ZN(n17176) );
  INV_X1 U20334 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18199) );
  NAND3_X1 U20335 ( .A1(n17176), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n17188), .ZN(
        n17175) );
  OAI221_X1 U20336 ( .B1(n17176), .B2(P3_EBX_REG_6__SCAN_IN), .C1(n17188), 
        .C2(n18199), .A(n17175), .ZN(P3_U2697) );
  INV_X1 U20337 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18194) );
  OAI211_X1 U20338 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n17177), .A(n17176), .B(
        n17188), .ZN(n17178) );
  OAI21_X1 U20339 ( .B1(n17188), .B2(n18194), .A(n17178), .ZN(P3_U2698) );
  OAI21_X1 U20340 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17180), .A(n17179), .ZN(
        n17181) );
  AOI22_X1 U20341 ( .A1(n17193), .A2(n18188), .B1(n17181), .B2(n17188), .ZN(
        P3_U2699) );
  INV_X1 U20342 ( .A(n17190), .ZN(n17192) );
  NAND2_X1 U20343 ( .A1(n17182), .A2(n17192), .ZN(n17185) );
  NAND3_X1 U20344 ( .A1(n17185), .A2(P3_EBX_REG_3__SCAN_IN), .A3(n17188), .ZN(
        n17183) );
  OAI221_X1 U20345 ( .B1(n17185), .B2(P3_EBX_REG_3__SCAN_IN), .C1(n17188), 
        .C2(n18182), .A(n17183), .ZN(P3_U2700) );
  AOI21_X1 U20346 ( .B1(n17195), .B2(n17184), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n17187) );
  NAND2_X1 U20347 ( .A1(n17188), .A2(n17185), .ZN(n17186) );
  OAI22_X1 U20348 ( .A1(n17187), .A2(n17186), .B1(n18176), .B2(n17188), .ZN(
        P3_U2701) );
  INV_X1 U20349 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18170) );
  OAI222_X1 U20350 ( .A1(n17191), .A2(n17190), .B1(n17189), .B2(n17195), .C1(
        n18170), .C2(n17188), .ZN(P3_U2702) );
  AOI22_X1 U20351 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17193), .B1(
        n17192), .B2(n20773), .ZN(n17194) );
  OAI21_X1 U20352 ( .B1(n17195), .B2(n20773), .A(n17194), .ZN(P3_U2703) );
  INV_X1 U20353 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17426) );
  NAND4_X1 U20354 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .A3(P3_EAX_REG_4__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17197) );
  NOR2_X1 U20355 ( .A1(n17343), .A2(n17197), .ZN(n17198) );
  NAND4_X1 U20356 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .A3(P3_EAX_REG_0__SCAN_IN), .A4(n17198), .ZN(n17309) );
  NAND2_X1 U20357 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .ZN(n17286) );
  NAND4_X1 U20358 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(P3_EAX_REG_8__SCAN_IN), .A4(n17199), .ZN(n17280) );
  NAND2_X1 U20359 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(P3_EAX_REG_17__SCAN_IN), 
        .ZN(n17243) );
  NAND4_X1 U20360 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_22__SCAN_IN), .A4(P3_EAX_REG_19__SCAN_IN), .ZN(n17200)
         );
  NOR3_X2 U20361 ( .A1(n17275), .A2(n17243), .A3(n17200), .ZN(n17239) );
  NAND2_X1 U20362 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17239), .ZN(n17238) );
  NOR2_X2 U20363 ( .A1(n17238), .A2(n18204), .ZN(n17234) );
  NAND2_X1 U20364 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17214), .ZN(n17209) );
  INV_X1 U20365 ( .A(n17209), .ZN(n17205) );
  NAND2_X1 U20366 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17205), .ZN(n17204) );
  NAND3_X1 U20367 ( .A1(n17327), .A2(P3_EAX_REG_31__SCAN_IN), .A3(n17204), 
        .ZN(n17203) );
  NAND2_X1 U20368 ( .A1(n17201), .A2(n17332), .ZN(n17249) );
  NAND2_X1 U20369 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17273), .ZN(n17202) );
  OAI211_X1 U20370 ( .C1(P3_EAX_REG_31__SCAN_IN), .C2(n17204), .A(n17203), .B(
        n17202), .ZN(P3_U2704) );
  NAND2_X1 U20371 ( .A1(n18191), .A2(n17332), .ZN(n17237) );
  AOI22_X1 U20372 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17274), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17273), .ZN(n17207) );
  OAI211_X1 U20373 ( .C1(n17205), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17327), .B(
        n17204), .ZN(n17206) );
  OAI211_X1 U20374 ( .C1(n17208), .C2(n17335), .A(n17207), .B(n17206), .ZN(
        P3_U2705) );
  AOI22_X1 U20375 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17274), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17273), .ZN(n17211) );
  OAI211_X1 U20376 ( .C1(n17214), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17327), .B(
        n17209), .ZN(n17210) );
  OAI211_X1 U20377 ( .C1(n17212), .C2(n17335), .A(n17211), .B(n17210), .ZN(
        P3_U2706) );
  INV_X1 U20378 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n18183) );
  AOI22_X1 U20379 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17274), .B1(n17340), .B2(
        n17213), .ZN(n17217) );
  AOI211_X1 U20380 ( .C1(n17426), .C2(n17218), .A(n17214), .B(n17332), .ZN(
        n17215) );
  INV_X1 U20381 ( .A(n17215), .ZN(n17216) );
  OAI211_X1 U20382 ( .C1(n17249), .C2(n18183), .A(n17217), .B(n17216), .ZN(
        P3_U2707) );
  AOI22_X1 U20383 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17274), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17273), .ZN(n17220) );
  OAI211_X1 U20384 ( .C1(n17223), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17327), .B(
        n17218), .ZN(n17219) );
  OAI211_X1 U20385 ( .C1(n17221), .C2(n17335), .A(n17220), .B(n17219), .ZN(
        P3_U2708) );
  AOI22_X1 U20386 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17274), .B1(n17340), .B2(
        n17222), .ZN(n17226) );
  AOI211_X1 U20387 ( .C1(n17422), .C2(n17227), .A(n17223), .B(n17332), .ZN(
        n17224) );
  INV_X1 U20388 ( .A(n17224), .ZN(n17225) );
  OAI211_X1 U20389 ( .C1(n17249), .C2(n19102), .A(n17226), .B(n17225), .ZN(
        P3_U2709) );
  AOI22_X1 U20390 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17274), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17273), .ZN(n17230) );
  OAI211_X1 U20391 ( .C1(n17228), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17327), .B(
        n17227), .ZN(n17229) );
  OAI211_X1 U20392 ( .C1(n17231), .C2(n17335), .A(n17230), .B(n17229), .ZN(
        P3_U2710) );
  AOI22_X1 U20393 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n17273), .B1(n17340), .B2(
        n17232), .ZN(n17236) );
  OAI211_X1 U20394 ( .C1(n17234), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17327), .B(
        n17233), .ZN(n17235) );
  OAI211_X1 U20395 ( .C1(n17237), .C2(n17440), .A(n17236), .B(n17235), .ZN(
        P3_U2711) );
  AOI22_X1 U20396 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17274), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17273), .ZN(n17241) );
  OAI211_X1 U20397 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17239), .A(n17327), .B(
        n17238), .ZN(n17240) );
  OAI211_X1 U20398 ( .C1(n17242), .C2(n17335), .A(n17241), .B(n17240), .ZN(
        P3_U2712) );
  NAND2_X1 U20399 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17263), .ZN(n17259) );
  NAND3_X1 U20400 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(n17255), .ZN(n17248) );
  AOI22_X1 U20401 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17273), .B1(n17340), .B2(
        n17244), .ZN(n17247) );
  NAND2_X1 U20402 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17255), .ZN(n17254) );
  NAND2_X1 U20403 ( .A1(n17327), .A2(n17254), .ZN(n17253) );
  OAI21_X1 U20404 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17342), .A(n17253), .ZN(
        n17245) );
  AOI22_X1 U20405 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17274), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17245), .ZN(n17246) );
  OAI211_X1 U20406 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17248), .A(n17247), .B(
        n17246), .ZN(P3_U2713) );
  INV_X1 U20407 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17412) );
  INV_X1 U20408 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n18189) );
  OAI22_X1 U20409 ( .A1(n17250), .A2(n17335), .B1(n18189), .B2(n17249), .ZN(
        n17251) );
  AOI21_X1 U20410 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17274), .A(n17251), .ZN(
        n17252) );
  OAI221_X1 U20411 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17254), .C1(n17412), 
        .C2(n17253), .A(n17252), .ZN(P3_U2714) );
  AOI22_X1 U20412 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17274), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17273), .ZN(n17257) );
  OAI211_X1 U20413 ( .C1(n17255), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17327), .B(
        n17254), .ZN(n17256) );
  OAI211_X1 U20414 ( .C1(n17258), .C2(n17335), .A(n17257), .B(n17256), .ZN(
        P3_U2715) );
  AOI22_X1 U20415 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17274), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17273), .ZN(n17261) );
  OAI211_X1 U20416 ( .C1(n17263), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17327), .B(
        n17259), .ZN(n17260) );
  OAI211_X1 U20417 ( .C1(n17262), .C2(n17335), .A(n17261), .B(n17260), .ZN(
        P3_U2716) );
  AOI22_X1 U20418 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17274), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17273), .ZN(n17266) );
  INV_X1 U20419 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17406) );
  INV_X1 U20420 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17404) );
  OR2_X1 U20421 ( .A1(n17404), .A2(n17275), .ZN(n17268) );
  AOI211_X1 U20422 ( .C1(n17406), .C2(n17268), .A(n17263), .B(n17332), .ZN(
        n17264) );
  INV_X1 U20423 ( .A(n17264), .ZN(n17265) );
  OAI211_X1 U20424 ( .C1(n17267), .C2(n17335), .A(n17266), .B(n17265), .ZN(
        P3_U2717) );
  AOI22_X1 U20425 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17274), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17273), .ZN(n17271) );
  INV_X1 U20426 ( .A(n17275), .ZN(n17269) );
  OAI211_X1 U20427 ( .C1(n17269), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17327), .B(
        n17268), .ZN(n17270) );
  OAI211_X1 U20428 ( .C1(n17272), .C2(n17335), .A(n17271), .B(n17270), .ZN(
        P3_U2718) );
  AOI22_X1 U20429 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17274), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17273), .ZN(n17278) );
  OAI211_X1 U20430 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17276), .A(n17327), .B(
        n17275), .ZN(n17277) );
  OAI211_X1 U20431 ( .C1(n17279), .C2(n17335), .A(n17278), .B(n17277), .ZN(
        P3_U2719) );
  NOR2_X1 U20432 ( .A1(n18204), .A2(n17280), .ZN(n17282) );
  NAND2_X1 U20433 ( .A1(n17327), .A2(n17280), .ZN(n17289) );
  INV_X1 U20434 ( .A(n17289), .ZN(n17281) );
  MUX2_X1 U20435 ( .A(n17282), .B(n17281), .S(P3_EAX_REG_15__SCAN_IN), .Z(
        n17283) );
  AOI21_X1 U20436 ( .B1(BUF2_REG_15__SCAN_IN), .B2(n17341), .A(n17283), .ZN(
        n17284) );
  OAI21_X1 U20437 ( .B1(n17285), .B2(n17335), .A(n17284), .ZN(P3_U2720) );
  NOR2_X1 U20438 ( .A1(n18204), .A2(n17309), .ZN(n17314) );
  NOR2_X1 U20439 ( .A1(n17286), .A2(n17302), .ZN(n17297) );
  NAND2_X1 U20440 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17297), .ZN(n17290) );
  AOI22_X1 U20441 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17341), .B1(n17340), .B2(
        n17287), .ZN(n17288) );
  OAI221_X1 U20442 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17290), .C1(n17453), 
        .C2(n17289), .A(n17288), .ZN(P3_U2721) );
  INV_X1 U20443 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17451) );
  INV_X1 U20444 ( .A(n17290), .ZN(n17293) );
  AOI21_X1 U20445 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17327), .A(n17297), .ZN(
        n17292) );
  OAI222_X1 U20446 ( .A1(n17338), .A2(n17451), .B1(n17293), .B2(n17292), .C1(
        n17335), .C2(n17291), .ZN(P3_U2722) );
  INV_X1 U20447 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17448) );
  INV_X1 U20448 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17375) );
  INV_X1 U20449 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17373) );
  OAI22_X1 U20450 ( .A1(n17302), .A2(n17375), .B1(n17373), .B2(n17332), .ZN(
        n17294) );
  INV_X1 U20451 ( .A(n17294), .ZN(n17296) );
  OAI222_X1 U20452 ( .A1(n17338), .A2(n17448), .B1(n17297), .B2(n17296), .C1(
        n17335), .C2(n17295), .ZN(P3_U2723) );
  NAND2_X1 U20453 ( .A1(n17302), .A2(P3_EAX_REG_11__SCAN_IN), .ZN(n17300) );
  AOI22_X1 U20454 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17341), .B1(n17340), .B2(
        n17298), .ZN(n17299) );
  OAI221_X1 U20455 ( .B1(n17302), .B2(P3_EAX_REG_11__SCAN_IN), .C1(n17300), 
        .C2(n17332), .A(n17299), .ZN(P3_U2724) );
  AOI22_X1 U20456 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17341), .B1(n17340), .B2(
        n17301), .ZN(n17304) );
  OAI211_X1 U20457 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n17307), .A(n17327), .B(
        n17302), .ZN(n17303) );
  NAND2_X1 U20458 ( .A1(n17304), .A2(n17303), .ZN(P3_U2725) );
  INV_X1 U20459 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17442) );
  AOI22_X1 U20460 ( .A1(n17314), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17327), .ZN(n17306) );
  OAI222_X1 U20461 ( .A1(n17338), .A2(n17442), .B1(n17307), .B2(n17306), .C1(
        n17335), .C2(n17305), .ZN(P3_U2726) );
  INV_X1 U20462 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17381) );
  AOI22_X1 U20463 ( .A1(n17340), .A2(n17308), .B1(n17314), .B2(n17381), .ZN(
        n17311) );
  NAND3_X1 U20464 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17327), .A3(n17309), .ZN(
        n17310) );
  OAI211_X1 U20465 ( .C1(n17338), .C2(n17440), .A(n17311), .B(n17310), .ZN(
        P3_U2727) );
  INV_X1 U20466 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18201) );
  INV_X1 U20467 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n20804) );
  INV_X1 U20468 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17388) );
  INV_X1 U20469 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17391) );
  NOR2_X1 U20470 ( .A1(n17432), .A2(n17342), .ZN(n17345) );
  NAND2_X1 U20471 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17345), .ZN(n17331) );
  NAND2_X1 U20472 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17337), .ZN(n17323) );
  NOR2_X1 U20473 ( .A1(n17388), .A2(n17323), .ZN(n17326) );
  NAND2_X1 U20474 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17326), .ZN(n17315) );
  NOR2_X1 U20475 ( .A1(n20804), .A2(n17315), .ZN(n17319) );
  AOI21_X1 U20476 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17327), .A(n17319), .ZN(
        n17313) );
  OAI222_X1 U20477 ( .A1(n17338), .A2(n18201), .B1(n17314), .B2(n17313), .C1(
        n17335), .C2(n17312), .ZN(P3_U2728) );
  INV_X1 U20478 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n20806) );
  INV_X1 U20479 ( .A(n17315), .ZN(n17322) );
  AOI21_X1 U20480 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17327), .A(n17322), .ZN(
        n17318) );
  INV_X1 U20481 ( .A(n17316), .ZN(n17317) );
  OAI222_X1 U20482 ( .A1(n20806), .A2(n17338), .B1(n17319), .B2(n17318), .C1(
        n17335), .C2(n17317), .ZN(P3_U2729) );
  AOI21_X1 U20483 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17327), .A(n17326), .ZN(
        n17321) );
  OAI222_X1 U20484 ( .A1(n18190), .A2(n17338), .B1(n17322), .B2(n17321), .C1(
        n17335), .C2(n17320), .ZN(P3_U2730) );
  INV_X1 U20485 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18184) );
  INV_X1 U20486 ( .A(n17323), .ZN(n17330) );
  AOI21_X1 U20487 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17327), .A(n17330), .ZN(
        n17325) );
  OAI222_X1 U20488 ( .A1(n18184), .A2(n17338), .B1(n17326), .B2(n17325), .C1(
        n17335), .C2(n9841), .ZN(P3_U2731) );
  INV_X1 U20489 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18177) );
  AOI21_X1 U20490 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17327), .A(n17337), .ZN(
        n17329) );
  OAI222_X1 U20491 ( .A1(n18177), .A2(n17338), .B1(n17330), .B2(n17329), .C1(
        n17335), .C2(n17328), .ZN(P3_U2732) );
  INV_X1 U20492 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18171) );
  OAI21_X1 U20493 ( .B1(n17391), .B2(n17332), .A(n17331), .ZN(n17333) );
  INV_X1 U20494 ( .A(n17333), .ZN(n17336) );
  OAI222_X1 U20495 ( .A1(n18171), .A2(n17338), .B1(n17337), .B2(n17336), .C1(
        n17335), .C2(n17334), .ZN(P3_U2733) );
  AOI22_X1 U20496 ( .A1(n17341), .A2(BUF2_REG_1__SCAN_IN), .B1(n17340), .B2(
        n17339), .ZN(n17347) );
  NOR2_X1 U20497 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17342), .ZN(n17344) );
  OAI22_X1 U20498 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17345), .B1(n17344), .B2(
        n17343), .ZN(n17346) );
  NAND2_X1 U20499 ( .A1(n17347), .A2(n17346), .ZN(P3_U2734) );
  INV_X1 U20500 ( .A(n17812), .ZN(n17648) );
  NAND2_X1 U20501 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17648), .ZN(n17352) );
  NOR2_X4 U20502 ( .A1(n17394), .A2(n17368), .ZN(n17365) );
  AND2_X1 U20503 ( .A1(n17365), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20504 ( .A(P3_UWORD_REG_14__SCAN_IN), .ZN(n20719) );
  INV_X1 U20505 ( .A(n17367), .ZN(n17350) );
  AOI22_X1 U20506 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17350), .B1(n17365), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17349) );
  OAI21_X1 U20507 ( .B1(n17352), .B2(n20719), .A(n17349), .ZN(P3_U2737) );
  INV_X1 U20508 ( .A(P3_UWORD_REG_13__SCAN_IN), .ZN(n20710) );
  AOI22_X1 U20509 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17350), .B1(n17365), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17351) );
  OAI21_X1 U20510 ( .B1(n17352), .B2(n20710), .A(n17351), .ZN(P3_U2738) );
  AOI22_X1 U20511 ( .A1(n17394), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17353) );
  OAI21_X1 U20512 ( .B1(n17426), .B2(n17367), .A(n17353), .ZN(P3_U2739) );
  INV_X1 U20513 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17424) );
  AOI22_X1 U20514 ( .A1(n17394), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17354) );
  OAI21_X1 U20515 ( .B1(n17424), .B2(n17367), .A(n17354), .ZN(P3_U2740) );
  AOI22_X1 U20516 ( .A1(n17394), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17355) );
  OAI21_X1 U20517 ( .B1(n17422), .B2(n17367), .A(n17355), .ZN(P3_U2741) );
  INV_X1 U20518 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17420) );
  AOI22_X1 U20519 ( .A1(n17394), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17356) );
  OAI21_X1 U20520 ( .B1(n17420), .B2(n17367), .A(n17356), .ZN(P3_U2742) );
  INV_X1 U20521 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17418) );
  AOI22_X1 U20522 ( .A1(n17394), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17357) );
  OAI21_X1 U20523 ( .B1(n17418), .B2(n17367), .A(n17357), .ZN(P3_U2743) );
  INV_X1 U20524 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17416) );
  AOI22_X1 U20525 ( .A1(n17394), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17358) );
  OAI21_X1 U20526 ( .B1(n17416), .B2(n17367), .A(n17358), .ZN(P3_U2744) );
  INV_X1 U20527 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17414) );
  AOI22_X1 U20528 ( .A1(n17394), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17359) );
  OAI21_X1 U20529 ( .B1(n17414), .B2(n17367), .A(n17359), .ZN(P3_U2745) );
  AOI22_X1 U20530 ( .A1(n17394), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17360) );
  OAI21_X1 U20531 ( .B1(n17412), .B2(n17367), .A(n17360), .ZN(P3_U2746) );
  INV_X1 U20532 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17410) );
  AOI22_X1 U20533 ( .A1(n17394), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17361) );
  OAI21_X1 U20534 ( .B1(n17410), .B2(n17367), .A(n17361), .ZN(P3_U2747) );
  INV_X1 U20535 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17408) );
  AOI22_X1 U20536 ( .A1(n17394), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(
        P3_DATAO_REG_19__SCAN_IN), .B2(n17365), .ZN(n17362) );
  OAI21_X1 U20537 ( .B1(n17408), .B2(n17367), .A(n17362), .ZN(P3_U2748) );
  AOI22_X1 U20538 ( .A1(n17394), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17363) );
  OAI21_X1 U20539 ( .B1(n17406), .B2(n17367), .A(n17363), .ZN(P3_U2749) );
  AOI22_X1 U20540 ( .A1(n17394), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17364) );
  OAI21_X1 U20541 ( .B1(n17404), .B2(n17367), .A(n17364), .ZN(P3_U2750) );
  INV_X1 U20542 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17402) );
  AOI22_X1 U20543 ( .A1(n17394), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17366) );
  OAI21_X1 U20544 ( .B1(n17402), .B2(n17367), .A(n17366), .ZN(P3_U2751) );
  AOI22_X1 U20545 ( .A1(n17394), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(
        P3_DATAO_REG_15__SCAN_IN), .B2(n17365), .ZN(n17369) );
  OAI21_X1 U20546 ( .B1(n17457), .B2(n17396), .A(n17369), .ZN(P3_U2752) );
  AOI22_X1 U20547 ( .A1(n17394), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17370) );
  OAI21_X1 U20548 ( .B1(n17453), .B2(n17396), .A(n17370), .ZN(P3_U2753) );
  AOI22_X1 U20549 ( .A1(n17394), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17371) );
  OAI21_X1 U20550 ( .B1(n20748), .B2(n17396), .A(n17371), .ZN(P3_U2754) );
  AOI22_X1 U20551 ( .A1(n17394), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17372) );
  OAI21_X1 U20552 ( .B1(n17373), .B2(n17396), .A(n17372), .ZN(P3_U2755) );
  AOI22_X1 U20553 ( .A1(n17394), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17374) );
  OAI21_X1 U20554 ( .B1(n17375), .B2(n17396), .A(n17374), .ZN(P3_U2756) );
  INV_X1 U20555 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17377) );
  AOI22_X1 U20556 ( .A1(n17394), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17376) );
  OAI21_X1 U20557 ( .B1(n17377), .B2(n17396), .A(n17376), .ZN(P3_U2757) );
  INV_X1 U20558 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17379) );
  AOI22_X1 U20559 ( .A1(n17394), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17378) );
  OAI21_X1 U20560 ( .B1(n17379), .B2(n17396), .A(n17378), .ZN(P3_U2758) );
  AOI22_X1 U20561 ( .A1(n17394), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17380) );
  OAI21_X1 U20562 ( .B1(n17381), .B2(n17396), .A(n17380), .ZN(P3_U2759) );
  INV_X1 U20563 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17383) );
  AOI22_X1 U20564 ( .A1(n17394), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17382) );
  OAI21_X1 U20565 ( .B1(n17383), .B2(n17396), .A(n17382), .ZN(P3_U2760) );
  AOI22_X1 U20566 ( .A1(n17394), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17384) );
  OAI21_X1 U20567 ( .B1(n20804), .B2(n17396), .A(n17384), .ZN(P3_U2761) );
  INV_X1 U20568 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17386) );
  AOI22_X1 U20569 ( .A1(n17394), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17385) );
  OAI21_X1 U20570 ( .B1(n17386), .B2(n17396), .A(n17385), .ZN(P3_U2762) );
  AOI22_X1 U20571 ( .A1(n17394), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17387) );
  OAI21_X1 U20572 ( .B1(n17388), .B2(n17396), .A(n17387), .ZN(P3_U2763) );
  INV_X1 U20573 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n20712) );
  AOI22_X1 U20574 ( .A1(n17394), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17389) );
  OAI21_X1 U20575 ( .B1(n20712), .B2(n17396), .A(n17389), .ZN(P3_U2764) );
  AOI22_X1 U20576 ( .A1(n17394), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17390) );
  OAI21_X1 U20577 ( .B1(n17391), .B2(n17396), .A(n17390), .ZN(P3_U2765) );
  INV_X1 U20578 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17393) );
  AOI22_X1 U20579 ( .A1(n17394), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17392) );
  OAI21_X1 U20580 ( .B1(n17393), .B2(n17396), .A(n17392), .ZN(P3_U2766) );
  AOI22_X1 U20581 ( .A1(n17394), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17365), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17395) );
  OAI21_X1 U20582 ( .B1(n17432), .B2(n17396), .A(n17395), .ZN(P3_U2767) );
  AOI22_X1 U20583 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17454), .ZN(n17401) );
  OAI21_X1 U20584 ( .B1(n17402), .B2(n20803), .A(n17401), .ZN(P3_U2768) );
  AOI22_X1 U20585 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17454), .ZN(n17403) );
  OAI21_X1 U20586 ( .B1(n17404), .B2(n20803), .A(n17403), .ZN(P3_U2769) );
  AOI22_X1 U20587 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17454), .ZN(n17405) );
  OAI21_X1 U20588 ( .B1(n17406), .B2(n20803), .A(n17405), .ZN(P3_U2770) );
  AOI22_X1 U20589 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17454), .ZN(n17407) );
  OAI21_X1 U20590 ( .B1(n17408), .B2(n20803), .A(n17407), .ZN(P3_U2771) );
  AOI22_X1 U20591 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17454), .ZN(n17409) );
  OAI21_X1 U20592 ( .B1(n17410), .B2(n20803), .A(n17409), .ZN(P3_U2772) );
  AOI22_X1 U20593 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17454), .ZN(n17411) );
  OAI21_X1 U20594 ( .B1(n17412), .B2(n20803), .A(n17411), .ZN(P3_U2773) );
  AOI22_X1 U20595 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17454), .ZN(n17413) );
  OAI21_X1 U20596 ( .B1(n17414), .B2(n20803), .A(n17413), .ZN(P3_U2774) );
  AOI22_X1 U20597 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17454), .ZN(n17415) );
  OAI21_X1 U20598 ( .B1(n17416), .B2(n20803), .A(n17415), .ZN(P3_U2775) );
  AOI22_X1 U20599 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17454), .ZN(n17417) );
  OAI21_X1 U20600 ( .B1(n17418), .B2(n20803), .A(n17417), .ZN(P3_U2776) );
  AOI22_X1 U20601 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17454), .ZN(n17419) );
  OAI21_X1 U20602 ( .B1(n17420), .B2(n20803), .A(n17419), .ZN(P3_U2777) );
  AOI22_X1 U20603 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17454), .ZN(n17421) );
  OAI21_X1 U20604 ( .B1(n17422), .B2(n20803), .A(n17421), .ZN(P3_U2778) );
  AOI22_X1 U20605 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17454), .ZN(n17423) );
  OAI21_X1 U20606 ( .B1(n17424), .B2(n20803), .A(n17423), .ZN(P3_U2779) );
  AOI22_X1 U20607 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17454), .ZN(n17425) );
  OAI21_X1 U20608 ( .B1(n17426), .B2(n20803), .A(n17425), .ZN(P3_U2780) );
  INV_X1 U20609 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17428) );
  AOI22_X1 U20610 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17454), .ZN(n17427) );
  OAI21_X1 U20611 ( .B1(n17428), .B2(n20803), .A(n17427), .ZN(P3_U2781) );
  AOI22_X1 U20612 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17455), .B1(
        P3_EAX_REG_30__SCAN_IN), .B2(n17449), .ZN(n17429) );
  OAI21_X1 U20613 ( .B1(n17430), .B2(n20719), .A(n17429), .ZN(P3_U2782) );
  AOI22_X1 U20614 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17454), .ZN(n17431) );
  OAI21_X1 U20615 ( .B1(n17432), .B2(n20803), .A(n17431), .ZN(P3_U2783) );
  INV_X1 U20616 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18165) );
  AOI22_X1 U20617 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17449), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17454), .ZN(n17433) );
  OAI21_X1 U20618 ( .B1(n18165), .B2(n20805), .A(n17433), .ZN(P3_U2784) );
  AOI22_X1 U20619 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17449), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17454), .ZN(n17434) );
  OAI21_X1 U20620 ( .B1(n18171), .B2(n20805), .A(n17434), .ZN(P3_U2785) );
  AOI22_X1 U20621 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17449), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17454), .ZN(n17435) );
  OAI21_X1 U20622 ( .B1(n18177), .B2(n20805), .A(n17435), .ZN(P3_U2786) );
  AOI22_X1 U20623 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17449), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17454), .ZN(n17436) );
  OAI21_X1 U20624 ( .B1(n18184), .B2(n20805), .A(n17436), .ZN(P3_U2787) );
  AOI22_X1 U20625 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17449), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17454), .ZN(n17437) );
  OAI21_X1 U20626 ( .B1(n18190), .B2(n20805), .A(n17437), .ZN(P3_U2788) );
  AOI22_X1 U20627 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17449), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17454), .ZN(n17438) );
  OAI21_X1 U20628 ( .B1(n18201), .B2(n20805), .A(n17438), .ZN(P3_U2790) );
  AOI22_X1 U20629 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17449), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17454), .ZN(n17439) );
  OAI21_X1 U20630 ( .B1(n17440), .B2(n20805), .A(n17439), .ZN(P3_U2791) );
  AOI22_X1 U20631 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17449), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17454), .ZN(n17441) );
  OAI21_X1 U20632 ( .B1(n17442), .B2(n20805), .A(n17441), .ZN(P3_U2792) );
  INV_X1 U20633 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17444) );
  AOI22_X1 U20634 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17449), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17454), .ZN(n17443) );
  OAI21_X1 U20635 ( .B1(n17444), .B2(n20805), .A(n17443), .ZN(P3_U2793) );
  INV_X1 U20636 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17446) );
  AOI22_X1 U20637 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17449), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17454), .ZN(n17445) );
  OAI21_X1 U20638 ( .B1(n17446), .B2(n20805), .A(n17445), .ZN(P3_U2794) );
  AOI22_X1 U20639 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17449), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17454), .ZN(n17447) );
  OAI21_X1 U20640 ( .B1(n17448), .B2(n20805), .A(n17447), .ZN(P3_U2795) );
  AOI22_X1 U20641 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17449), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17454), .ZN(n17450) );
  OAI21_X1 U20642 ( .B1(n17451), .B2(n20805), .A(n17450), .ZN(P3_U2796) );
  AOI22_X1 U20643 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17454), .ZN(n17452) );
  OAI21_X1 U20644 ( .B1(n17453), .B2(n20803), .A(n17452), .ZN(P3_U2797) );
  AOI22_X1 U20645 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17454), .ZN(n17456) );
  OAI21_X1 U20646 ( .B1(n17457), .B2(n20803), .A(n17456), .ZN(P3_U2798) );
  INV_X1 U20647 ( .A(n17762), .ZN(n17715) );
  OAI21_X1 U20648 ( .B1(n17458), .B2(n17715), .A(n17811), .ZN(n17459) );
  AOI21_X1 U20649 ( .B1(n17648), .B2(n17460), .A(n17459), .ZN(n17489) );
  OAI21_X1 U20650 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17564), .A(
        n17489), .ZN(n17481) );
  AOI22_X1 U20651 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17481), .B1(
        n17609), .B2(n17461), .ZN(n17476) );
  NOR2_X1 U20652 ( .A1(n17803), .A2(n17724), .ZN(n17559) );
  OAI22_X1 U20653 ( .A1(n17824), .A2(n17816), .B1(n17462), .B2(n16334), .ZN(
        n17494) );
  NOR2_X1 U20654 ( .A1(n17818), .A2(n17494), .ZN(n17464) );
  NOR3_X1 U20655 ( .A1(n17559), .A2(n17464), .A3(n17463), .ZN(n17469) );
  AOI211_X1 U20656 ( .C1(n17467), .C2(n17466), .A(n17465), .B(n17632), .ZN(
        n17468) );
  AOI211_X1 U20657 ( .C1(n17517), .C2(n17470), .A(n17469), .B(n17468), .ZN(
        n17475) );
  NAND2_X1 U20658 ( .A1(n9846), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17474) );
  NOR2_X1 U20659 ( .A1(n17611), .A2(n17471), .ZN(n17483) );
  OAI211_X1 U20660 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17483), .B(n17472), .ZN(n17473) );
  NAND4_X1 U20661 ( .A1(n17476), .A2(n17475), .A3(n17474), .A4(n17473), .ZN(
        P3_U2802) );
  NOR2_X1 U20662 ( .A1(n9676), .A2(n17477), .ZN(n17478) );
  XOR2_X1 U20663 ( .A(n17478), .B(n17722), .Z(n17831) );
  OAI22_X1 U20664 ( .A1(n18094), .A2(n18733), .B1(n17663), .B2(n17479), .ZN(
        n17480) );
  AOI221_X1 U20665 ( .B1(n17483), .B2(n17482), .C1(n17481), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17480), .ZN(n17486) );
  INV_X1 U20666 ( .A(n17517), .ZN(n17532) );
  NOR2_X1 U20667 ( .A1(n17817), .A2(n17532), .ZN(n17484) );
  AOI22_X1 U20668 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17494), .B1(
        n17484), .B2(n17818), .ZN(n17485) );
  OAI211_X1 U20669 ( .C1(n17831), .C2(n17632), .A(n17486), .B(n17485), .ZN(
        P3_U2803) );
  INV_X1 U20670 ( .A(n17841), .ZN(n17843) );
  NAND3_X1 U20671 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17843), .A3(
        n17833), .ZN(n17838) );
  AOI21_X1 U20672 ( .B1(n17487), .B2(n18545), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17488) );
  INV_X1 U20673 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18731) );
  OAI22_X1 U20674 ( .A1(n17489), .A2(n17488), .B1(n18094), .B2(n18731), .ZN(
        n17490) );
  AOI221_X1 U20675 ( .B1(n17609), .B2(n17491), .C1(n17596), .C2(n17491), .A(
        n17490), .ZN(n17496) );
  OAI21_X1 U20676 ( .B1(n17493), .B2(n17833), .A(n17492), .ZN(n17836) );
  AOI22_X1 U20677 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17494), .B1(
        n17723), .B2(n17836), .ZN(n17495) );
  OAI211_X1 U20678 ( .C1(n17532), .C2(n17838), .A(n17496), .B(n17495), .ZN(
        P3_U2804) );
  OAI21_X1 U20679 ( .B1(n17497), .B2(n17812), .A(n17811), .ZN(n17498) );
  AOI21_X1 U20680 ( .B1(n18545), .B2(n9670), .A(n17498), .ZN(n17528) );
  OAI21_X1 U20681 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17564), .A(
        n17528), .ZN(n17512) );
  AOI22_X1 U20682 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17512), .B1(
        n17609), .B2(n17499), .ZN(n17508) );
  XOR2_X1 U20683 ( .A(n17500), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17852) );
  XOR2_X1 U20684 ( .A(n17501), .B(n17845), .Z(n17854) );
  OAI21_X1 U20685 ( .B1(n17722), .B2(n10038), .A(n17502), .ZN(n17503) );
  XOR2_X1 U20686 ( .A(n17503), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17850) );
  OAI22_X1 U20687 ( .A1(n17816), .A2(n17854), .B1(n17632), .B2(n17850), .ZN(
        n17504) );
  AOI21_X1 U20688 ( .B1(n17724), .B2(n17852), .A(n17504), .ZN(n17507) );
  NAND2_X1 U20689 ( .A1(n9846), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17848) );
  NOR2_X1 U20690 ( .A1(n17611), .A2(n9670), .ZN(n17514) );
  OAI211_X1 U20691 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17514), .B(n17505), .ZN(n17506) );
  NAND4_X1 U20692 ( .A1(n17508), .A2(n17507), .A3(n17848), .A4(n17506), .ZN(
        P3_U2805) );
  AOI22_X1 U20693 ( .A1(n17803), .A2(n17859), .B1(n17724), .B2(n17858), .ZN(
        n17531) );
  AOI22_X1 U20694 ( .A1(n9846), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n17609), 
        .B2(n17509), .ZN(n17510) );
  INV_X1 U20695 ( .A(n17510), .ZN(n17511) );
  AOI221_X1 U20696 ( .B1(n17514), .B2(n17513), .C1(n17512), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17511), .ZN(n17519) );
  OAI21_X1 U20697 ( .B1(n17516), .B2(n17520), .A(n17515), .ZN(n17857) );
  NOR2_X1 U20698 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17867), .ZN(
        n17855) );
  AOI22_X1 U20699 ( .A1(n17723), .A2(n17857), .B1(n17517), .B2(n17855), .ZN(
        n17518) );
  OAI211_X1 U20700 ( .C1(n17531), .C2(n17520), .A(n17519), .B(n17518), .ZN(
        P3_U2806) );
  OAI22_X1 U20701 ( .A1(n17722), .A2(n17886), .B1(n17521), .B2(n17536), .ZN(
        n17522) );
  NOR2_X1 U20702 ( .A1(n17522), .A2(n17560), .ZN(n17523) );
  XOR2_X1 U20703 ( .A(n17523), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(
        n17871) );
  AOI21_X1 U20704 ( .B1(n17524), .B2(n18545), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17527) );
  OAI21_X1 U20705 ( .B1(n17609), .B2(n17596), .A(n17525), .ZN(n17526) );
  NAND2_X1 U20706 ( .A1(n9846), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17872) );
  OAI211_X1 U20707 ( .C1(n17528), .C2(n17527), .A(n17526), .B(n17872), .ZN(
        n17529) );
  AOI21_X1 U20708 ( .B1(n17723), .B2(n17871), .A(n17529), .ZN(n17530) );
  OAI221_X1 U20709 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17532), 
        .C1(n17867), .C2(n17531), .A(n17530), .ZN(P3_U2807) );
  INV_X1 U20710 ( .A(n17533), .ZN(n17535) );
  INV_X1 U20711 ( .A(n17560), .ZN(n17534) );
  OAI221_X1 U20712 ( .B1(n17536), .B2(n17535), .C1(n17536), .C2(n17549), .A(
        n17534), .ZN(n17537) );
  XOR2_X1 U20713 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17537), .Z(
        n17891) );
  NOR2_X1 U20714 ( .A1(n17962), .A2(n16334), .ZN(n17629) );
  NOR2_X1 U20715 ( .A1(n17883), .A2(n17816), .ZN(n17628) );
  NOR2_X1 U20716 ( .A1(n17629), .A2(n17628), .ZN(n17617) );
  OAI21_X1 U20717 ( .B1(n17880), .B2(n17559), .A(n17617), .ZN(n17556) );
  OR2_X1 U20718 ( .A1(n9702), .A2(n17611), .ZN(n17553) );
  AOI211_X1 U20719 ( .C1(n20720), .C2(n17544), .A(n17538), .B(n17553), .ZN(
        n17546) );
  AOI22_X1 U20720 ( .A1(n17648), .A2(n17539), .B1(n17762), .B2(n9702), .ZN(
        n17540) );
  NAND2_X1 U20721 ( .A1(n17540), .A2(n17811), .ZN(n17563) );
  AOI21_X1 U20722 ( .B1(n17596), .B2(n17541), .A(n17563), .ZN(n17552) );
  AOI22_X1 U20723 ( .A1(n9846), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n17609), 
        .B2(n17542), .ZN(n17543) );
  OAI21_X1 U20724 ( .B1(n17552), .B2(n17544), .A(n17543), .ZN(n17545) );
  AOI211_X1 U20725 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17556), .A(
        n17546), .B(n17545), .ZN(n17548) );
  NAND3_X1 U20726 ( .A1(n17880), .A2(n17601), .A3(n17886), .ZN(n17547) );
  OAI211_X1 U20727 ( .C1(n17632), .C2(n17891), .A(n17548), .B(n17547), .ZN(
        P3_U2808) );
  NAND3_X1 U20728 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17722), .A3(
        n17549), .ZN(n17569) );
  OAI22_X1 U20729 ( .A1(n17893), .A2(n17569), .B1(n17590), .B2(n17550), .ZN(
        n17551) );
  XNOR2_X1 U20730 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17551), .ZN(
        n17903) );
  NAND2_X1 U20731 ( .A1(n9846), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n17901) );
  OAI221_X1 U20732 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17553), .C1(
        n20720), .C2(n17552), .A(n17901), .ZN(n17554) );
  AOI21_X1 U20733 ( .B1(n17609), .B2(n17555), .A(n17554), .ZN(n17558) );
  NOR2_X1 U20734 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17893), .ZN(
        n17899) );
  NAND2_X1 U20735 ( .A1(n17932), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17894) );
  NOR2_X1 U20736 ( .A1(n17618), .A2(n17894), .ZN(n17581) );
  AOI22_X1 U20737 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17556), .B1(
        n17899), .B2(n17581), .ZN(n17557) );
  OAI211_X1 U20738 ( .C1(n17903), .C2(n17632), .A(n17558), .B(n17557), .ZN(
        P3_U2809) );
  INV_X1 U20739 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n20679) );
  NOR2_X1 U20740 ( .A1(n20679), .A2(n17894), .ZN(n17906) );
  OAI21_X1 U20741 ( .B1(n17559), .B2(n17906), .A(n17617), .ZN(n17580) );
  AOI221_X1 U20742 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17569), 
        .C1(n20679), .C2(n17589), .A(n17560), .ZN(n17561) );
  XOR2_X1 U20743 ( .A(n17878), .B(n17561), .Z(n17920) );
  NAND2_X1 U20744 ( .A1(n17906), .A2(n17878), .ZN(n17913) );
  OAI22_X1 U20745 ( .A1(n17632), .A2(n17920), .B1(n17618), .B2(n17913), .ZN(
        n17562) );
  AOI21_X1 U20746 ( .B1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n17580), .A(
        n17562), .ZN(n17568) );
  NAND2_X1 U20747 ( .A1(n9846), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17918) );
  OAI221_X1 U20748 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n16524), .C1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n18545), .A(n17563), .ZN(
        n17567) );
  OAI21_X1 U20749 ( .B1(n17609), .B2(n17596), .A(n17565), .ZN(n17566) );
  NAND4_X1 U20750 ( .A1(n17568), .A2(n17918), .A3(n17567), .A4(n17566), .ZN(
        P3_U2810) );
  OAI21_X1 U20751 ( .B1(n17589), .B2(n17590), .A(n17569), .ZN(n17570) );
  XOR2_X1 U20752 ( .A(n17570), .B(n20679), .Z(n17926) );
  AOI21_X1 U20753 ( .B1(n17574), .B2(n17762), .A(n17798), .ZN(n17571) );
  INV_X1 U20754 ( .A(n17571), .ZN(n17597) );
  AOI21_X1 U20755 ( .B1(n17648), .B2(n17572), .A(n17597), .ZN(n17584) );
  AOI22_X1 U20756 ( .A1(n9846), .A2(P3_REIP_REG_19__SCAN_IN), .B1(n17609), 
        .B2(n17573), .ZN(n17577) );
  NOR2_X1 U20757 ( .A1(n17611), .A2(n17574), .ZN(n17583) );
  OAI211_X1 U20758 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17583), .B(n17575), .ZN(n17576) );
  OAI211_X1 U20759 ( .C1(n17584), .C2(n17578), .A(n17577), .B(n17576), .ZN(
        n17579) );
  AOI221_X1 U20760 ( .B1(n17581), .B2(n20679), .C1(n17580), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n17579), .ZN(n17582) );
  OAI21_X1 U20761 ( .B1(n17926), .B2(n17632), .A(n17582), .ZN(P3_U2811) );
  NAND2_X1 U20762 ( .A1(n17932), .A2(n17898), .ZN(n17939) );
  INV_X1 U20763 ( .A(n17583), .ZN(n17586) );
  NAND2_X1 U20764 ( .A1(n9846), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17937) );
  OAI221_X1 U20765 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17586), .C1(
        n17585), .C2(n17584), .A(n17937), .ZN(n17587) );
  AOI21_X1 U20766 ( .B1(n17609), .B2(n17588), .A(n17587), .ZN(n17593) );
  OAI21_X1 U20767 ( .B1(n17932), .B2(n17618), .A(n17617), .ZN(n17602) );
  OAI21_X1 U20768 ( .B1(n17898), .B2(n10223), .A(n17589), .ZN(n17591) );
  XOR2_X1 U20769 ( .A(n17591), .B(n17590), .Z(n17935) );
  AOI22_X1 U20770 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17602), .B1(
        n17723), .B2(n17935), .ZN(n17592) );
  OAI211_X1 U20771 ( .C1(n17618), .C2(n17939), .A(n17593), .B(n17592), .ZN(
        P3_U2812) );
  AOI21_X1 U20772 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17595), .A(
        n17594), .ZN(n17948) );
  NAND2_X1 U20773 ( .A1(n9846), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n17945) );
  OAI221_X1 U20774 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16526), .C1(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n18545), .A(n17597), .ZN(
        n17598) );
  NAND2_X1 U20775 ( .A1(n17945), .A2(n17598), .ZN(n17599) );
  AOI21_X1 U20776 ( .B1(n17600), .B2(n17805), .A(n17599), .ZN(n17604) );
  NOR2_X1 U20777 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17957), .ZN(
        n17944) );
  AOI22_X1 U20778 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17602), .B1(
        n17601), .B2(n17944), .ZN(n17603) );
  OAI211_X1 U20779 ( .C1(n17948), .C2(n17632), .A(n17604), .B(n17603), .ZN(
        P3_U2813) );
  NAND2_X1 U20780 ( .A1(n17722), .A2(n18015), .ZN(n17690) );
  INV_X1 U20781 ( .A(n17690), .ZN(n17699) );
  AOI22_X1 U20782 ( .A1(n17699), .A2(n17929), .B1(n17605), .B2(n10223), .ZN(
        n17606) );
  XOR2_X1 U20783 ( .A(n17957), .B(n17606), .Z(n17954) );
  AOI21_X1 U20784 ( .B1(n17762), .B2(n17610), .A(n17798), .ZN(n17635) );
  OAI21_X1 U20785 ( .B1(n17607), .B2(n17812), .A(n17635), .ZN(n17625) );
  AOI22_X1 U20786 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17625), .B1(
        n17609), .B2(n17608), .ZN(n17614) );
  NOR2_X1 U20787 ( .A1(n17611), .A2(n17610), .ZN(n17627) );
  OAI211_X1 U20788 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17627), .B(n17612), .ZN(n17613) );
  OAI211_X1 U20789 ( .C1(n18713), .C2(n18094), .A(n17614), .B(n17613), .ZN(
        n17615) );
  AOI21_X1 U20790 ( .B1(n17723), .B2(n17954), .A(n17615), .ZN(n17616) );
  OAI221_X1 U20791 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17618), 
        .C1(n17957), .C2(n17617), .A(n17616), .ZN(P3_U2814) );
  INV_X1 U20792 ( .A(n17619), .ZN(n17655) );
  NAND3_X1 U20793 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17722), .A3(
        n17655), .ZN(n17621) );
  NOR2_X1 U20794 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n10209), .ZN(
        n18001) );
  AOI21_X1 U20795 ( .B1(n17621), .B2(n17620), .A(n18001), .ZN(n17622) );
  XNOR2_X1 U20796 ( .A(n17622), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17969) );
  NAND2_X1 U20797 ( .A1(n9846), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n17971) );
  OAI21_X1 U20798 ( .B1(n17663), .B2(n17623), .A(n17971), .ZN(n17624) );
  AOI221_X1 U20799 ( .B1(n17627), .B2(n17626), .C1(n17625), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17624), .ZN(n17631) );
  OAI21_X1 U20800 ( .B1(n17640), .B2(n17995), .A(n10208), .ZN(n17966) );
  NAND2_X1 U20801 ( .A1(n17633), .A2(n10208), .ZN(n17964) );
  AOI22_X1 U20802 ( .A1(n17629), .A2(n17966), .B1(n17628), .B2(n17964), .ZN(
        n17630) );
  OAI211_X1 U20803 ( .C1(n17632), .C2(n17969), .A(n17631), .B(n17630), .ZN(
        P3_U2815) );
  NAND2_X1 U20804 ( .A1(n18013), .A2(n17975), .ZN(n17646) );
  INV_X1 U20805 ( .A(n17646), .ZN(n17993) );
  OAI221_X1 U20806 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17993), .A(n17633), .ZN(
        n17988) );
  NAND2_X1 U20807 ( .A1(n17634), .A2(n18545), .ZN(n17676) );
  AOI221_X1 U20808 ( .B1(n17637), .B2(n17636), .C1(n17676), .C2(n17636), .A(
        n17635), .ZN(n17638) );
  NOR2_X1 U20809 ( .A1(n18094), .A2(n18710), .ZN(n17982) );
  AOI211_X1 U20810 ( .C1(n17639), .C2(n17805), .A(n17638), .B(n17982), .ZN(
        n17645) );
  NAND2_X1 U20811 ( .A1(n17975), .A2(n18015), .ZN(n17989) );
  NOR2_X1 U20812 ( .A1(n17640), .A2(n17995), .ZN(n17641) );
  AOI221_X1 U20813 ( .B1(n17660), .B2(n17979), .C1(n17989), .C2(n17979), .A(
        n17641), .ZN(n17985) );
  AOI22_X1 U20814 ( .A1(n17699), .A2(n17974), .B1(n17642), .B2(n10209), .ZN(
        n17643) );
  XOR2_X1 U20815 ( .A(n17979), .B(n17643), .Z(n17984) );
  AOI22_X1 U20816 ( .A1(n17724), .A2(n17985), .B1(n17723), .B2(n17984), .ZN(
        n17644) );
  OAI211_X1 U20817 ( .C1(n17816), .C2(n17988), .A(n17645), .B(n17644), .ZN(
        P3_U2816) );
  AOI22_X1 U20818 ( .A1(n17803), .A2(n17646), .B1(n17724), .B2(n17989), .ZN(
        n17672) );
  AOI21_X1 U20819 ( .B1(n17648), .B2(n17647), .A(n17798), .ZN(n17649) );
  OAI21_X1 U20820 ( .B1(n17634), .B2(n17715), .A(n17649), .ZN(n17665) );
  NOR2_X1 U20821 ( .A1(n18094), .A2(n18707), .ZN(n17654) );
  OAI211_X1 U20822 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17634), .B(n17661), .ZN(n17651) );
  OAI22_X1 U20823 ( .A1(n17652), .A2(n17651), .B1(n17650), .B2(n17663), .ZN(
        n17653) );
  AOI211_X1 U20824 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17665), .A(
        n17654), .B(n17653), .ZN(n17659) );
  AOI21_X1 U20825 ( .B1(n10209), .B2(n10223), .A(n17655), .ZN(n17656) );
  AOI21_X1 U20826 ( .B1(n10223), .B2(n17667), .A(n17656), .ZN(n17657) );
  XOR2_X1 U20827 ( .A(n17657), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n18002) );
  INV_X1 U20828 ( .A(n18021), .ZN(n18000) );
  NOR2_X1 U20829 ( .A1(n17709), .A2(n18000), .ZN(n17669) );
  AOI22_X1 U20830 ( .A1(n17723), .A2(n18002), .B1(n18001), .B2(n17669), .ZN(
        n17658) );
  OAI211_X1 U20831 ( .C1(n17672), .C2(n17660), .A(n17659), .B(n17658), .ZN(
        P3_U2817) );
  AND2_X1 U20832 ( .A1(n17661), .A2(n17634), .ZN(n17666) );
  OAI22_X1 U20833 ( .A1(n18094), .A2(n18705), .B1(n17663), .B2(n17662), .ZN(
        n17664) );
  AOI221_X1 U20834 ( .B1(n17666), .B2(n20680), .C1(n17665), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17664), .ZN(n17671) );
  OAI21_X1 U20835 ( .B1(n18000), .B2(n17690), .A(n17667), .ZN(n17668) );
  XOR2_X1 U20836 ( .A(n17668), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18005) );
  AOI22_X1 U20837 ( .A1(n17723), .A2(n18005), .B1(n17669), .B2(n10209), .ZN(
        n17670) );
  OAI211_X1 U20838 ( .C1(n17672), .C2(n10209), .A(n17671), .B(n17670), .ZN(
        P3_U2818) );
  NOR3_X1 U20839 ( .A1(n17743), .A2(n17747), .A3(n18507), .ZN(n17731) );
  NAND2_X1 U20840 ( .A1(n17673), .A2(n17731), .ZN(n17687) );
  OAI21_X1 U20841 ( .B1(n17702), .B2(n17674), .A(n17687), .ZN(n17675) );
  AOI22_X1 U20842 ( .A1(n17677), .A2(n17805), .B1(n17676), .B2(n17675), .ZN(
        n17684) );
  INV_X1 U20843 ( .A(n17680), .ZN(n18020) );
  AOI21_X1 U20844 ( .B1(n18020), .B2(n17699), .A(n9709), .ZN(n17678) );
  XOR2_X1 U20845 ( .A(n17679), .B(n17678), .Z(n18012) );
  NOR2_X1 U20846 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17680), .ZN(
        n18011) );
  INV_X1 U20847 ( .A(n17709), .ZN(n17681) );
  AOI22_X1 U20848 ( .A1(n17723), .A2(n18012), .B1(n18011), .B2(n17681), .ZN(
        n17683) );
  NOR2_X1 U20849 ( .A1(n18020), .A2(n17709), .ZN(n17693) );
  INV_X1 U20850 ( .A(n18013), .ZN(n17997) );
  AOI22_X1 U20851 ( .A1(n17995), .A2(n17724), .B1(n17803), .B2(n17997), .ZN(
        n17708) );
  INV_X1 U20852 ( .A(n17708), .ZN(n17692) );
  OAI21_X1 U20853 ( .B1(n17693), .B2(n17692), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17682) );
  NAND2_X1 U20854 ( .A1(n9846), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n18025) );
  NAND4_X1 U20855 ( .A1(n17684), .A2(n17683), .A3(n17682), .A4(n18025), .ZN(
        P3_U2819) );
  NAND3_X1 U20856 ( .A1(n17712), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        n17731), .ZN(n17701) );
  OAI21_X1 U20857 ( .B1(n17702), .B2(n17685), .A(n17701), .ZN(n17686) );
  AOI22_X1 U20858 ( .A1(n17688), .A2(n17805), .B1(n17687), .B2(n17686), .ZN(
        n17697) );
  OAI21_X1 U20859 ( .B1(n18045), .B2(n17690), .A(n17689), .ZN(n17691) );
  XOR2_X1 U20860 ( .A(n17691), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .Z(
        n18030) );
  AOI22_X1 U20861 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17692), .B1(
        n17723), .B2(n18030), .ZN(n17696) );
  NAND2_X1 U20862 ( .A1(n9846), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n17695) );
  OAI21_X1 U20863 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n17693), .ZN(n17694) );
  NAND4_X1 U20864 ( .A1(n17697), .A2(n17696), .A3(n17695), .A4(n17694), .ZN(
        P3_U2820) );
  NOR2_X1 U20865 ( .A1(n17699), .A2(n17698), .ZN(n17700) );
  XOR2_X1 U20866 ( .A(n17700), .B(n18045), .Z(n18042) );
  NOR2_X1 U20867 ( .A1(n18094), .A2(n18699), .ZN(n18041) );
  INV_X1 U20868 ( .A(n17701), .ZN(n17705) );
  INV_X1 U20869 ( .A(n17702), .ZN(n17806) );
  AOI22_X1 U20870 ( .A1(n17712), .A2(n17731), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17806), .ZN(n17704) );
  OAI22_X1 U20871 ( .A1(n17705), .A2(n17704), .B1(n17795), .B2(n17703), .ZN(
        n17706) );
  AOI211_X1 U20872 ( .C1(n17723), .C2(n18042), .A(n18041), .B(n17706), .ZN(
        n17707) );
  OAI221_X1 U20873 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17709), .C1(
        n18045), .C2(n17708), .A(n17707), .ZN(P3_U2821) );
  OAI21_X1 U20874 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17711), .A(
        n17710), .ZN(n18062) );
  NAND2_X1 U20875 ( .A1(n17714), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17713) );
  AOI211_X1 U20876 ( .C1(n17716), .C2(n17713), .A(n17712), .B(n18507), .ZN(
        n17720) );
  OAI21_X1 U20877 ( .B1(n17715), .B2(n17714), .A(n17811), .ZN(n17729) );
  INV_X1 U20878 ( .A(n17729), .ZN(n17717) );
  OAI22_X1 U20879 ( .A1(n17795), .A2(n17718), .B1(n17717), .B2(n17716), .ZN(
        n17719) );
  AOI211_X1 U20880 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n9846), .A(n17720), .B(
        n17719), .ZN(n17726) );
  OAI21_X1 U20881 ( .B1(n17722), .B2(n18059), .A(n17721), .ZN(n18056) );
  AOI22_X1 U20882 ( .A1(n17724), .A2(n18059), .B1(n17723), .B2(n18056), .ZN(
        n17725) );
  OAI211_X1 U20883 ( .C1(n17816), .C2(n18062), .A(n17726), .B(n17725), .ZN(
        P3_U2822) );
  OAI21_X1 U20884 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17728), .A(
        n17727), .ZN(n18071) );
  NOR2_X1 U20885 ( .A1(n18094), .A2(n20777), .ZN(n18067) );
  AOI221_X1 U20886 ( .B1(n17731), .B2(n17730), .C1(n17729), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18067), .ZN(n17737) );
  NOR2_X1 U20887 ( .A1(n17733), .A2(n17732), .ZN(n17734) );
  XOR2_X1 U20888 ( .A(n17734), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18068) );
  AOI22_X1 U20889 ( .A1(n17803), .A2(n18068), .B1(n17735), .B2(n17805), .ZN(
        n17736) );
  OAI211_X1 U20890 ( .C1(n17815), .C2(n18071), .A(n17737), .B(n17736), .ZN(
        P3_U2823) );
  OAI21_X1 U20891 ( .B1(n17740), .B2(n17739), .A(n17738), .ZN(n18075) );
  NOR2_X1 U20892 ( .A1(n17743), .A2(n18507), .ZN(n17748) );
  OAI21_X1 U20893 ( .B1(n17742), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n17741), .ZN(n18080) );
  OAI22_X1 U20894 ( .A1(n17816), .A2(n18080), .B1(n18094), .B2(n18694), .ZN(
        n17746) );
  OAI21_X1 U20895 ( .B1(n18507), .B2(n17743), .A(n17806), .ZN(n17756) );
  OAI22_X1 U20896 ( .A1(n17795), .A2(n17744), .B1(n17747), .B2(n17756), .ZN(
        n17745) );
  AOI211_X1 U20897 ( .C1(n17748), .C2(n17747), .A(n17746), .B(n17745), .ZN(
        n17749) );
  OAI21_X1 U20898 ( .B1(n17815), .B2(n18075), .A(n17749), .ZN(P3_U2824) );
  OAI21_X1 U20899 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17751), .A(
        n17750), .ZN(n18082) );
  AOI21_X1 U20900 ( .B1(n16798), .B2(n17811), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17757) );
  OAI21_X1 U20901 ( .B1(n17754), .B2(n17753), .A(n17752), .ZN(n17755) );
  XOR2_X1 U20902 ( .A(n17755), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(
        n18088) );
  OAI22_X1 U20903 ( .A1(n17757), .A2(n17756), .B1(n17816), .B2(n18088), .ZN(
        n17758) );
  AOI21_X1 U20904 ( .B1(n17759), .B2(n17805), .A(n17758), .ZN(n17760) );
  NAND2_X1 U20905 ( .A1(n9846), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18081) );
  OAI211_X1 U20906 ( .C1(n17815), .C2(n18082), .A(n17760), .B(n18081), .ZN(
        P3_U2825) );
  AOI21_X1 U20907 ( .B1(n17762), .B2(n17761), .A(n17798), .ZN(n17784) );
  OAI21_X1 U20908 ( .B1(n17765), .B2(n17764), .A(n17763), .ZN(n17766) );
  XOR2_X1 U20909 ( .A(n17766), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(
        n18100) );
  OAI22_X1 U20910 ( .A1(n17816), .A2(n18100), .B1(n18094), .B2(n18690), .ZN(
        n17772) );
  OAI21_X1 U20911 ( .B1(n17769), .B2(n17768), .A(n17767), .ZN(n18093) );
  OAI22_X1 U20912 ( .A1(n17795), .A2(n17770), .B1(n17815), .B2(n18093), .ZN(
        n17771) );
  AOI211_X1 U20913 ( .C1(n18545), .C2(n17773), .A(n17772), .B(n17771), .ZN(
        n17774) );
  OAI21_X1 U20914 ( .B1(n17784), .B2(n17775), .A(n17774), .ZN(P3_U2826) );
  OAI21_X1 U20915 ( .B1(n17778), .B2(n17777), .A(n17776), .ZN(n18104) );
  AOI21_X1 U20916 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17811), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17783) );
  OAI21_X1 U20917 ( .B1(n17781), .B2(n17780), .A(n17779), .ZN(n17782) );
  XOR2_X1 U20918 ( .A(n17782), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(
        n18105) );
  OAI22_X1 U20919 ( .A1(n17784), .A2(n17783), .B1(n17815), .B2(n18105), .ZN(
        n17785) );
  AOI21_X1 U20920 ( .B1(n17786), .B2(n17805), .A(n17785), .ZN(n17787) );
  NAND2_X1 U20921 ( .A1(n9846), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18108) );
  OAI211_X1 U20922 ( .C1(n17816), .C2(n18104), .A(n17787), .B(n18108), .ZN(
        P3_U2827) );
  OAI21_X1 U20923 ( .B1(n17790), .B2(n17789), .A(n17788), .ZN(n18124) );
  OAI21_X1 U20924 ( .B1(n17793), .B2(n17792), .A(n17791), .ZN(n18119) );
  OAI22_X1 U20925 ( .A1(n17795), .A2(n17794), .B1(n17815), .B2(n18119), .ZN(
        n17796) );
  AOI221_X1 U20926 ( .B1(n17798), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18545), .C2(n17797), .A(n17796), .ZN(n17799) );
  NAND2_X1 U20927 ( .A1(n9846), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18122) );
  OAI211_X1 U20928 ( .C1(n17816), .C2(n18124), .A(n17799), .B(n18122), .ZN(
        P3_U2828) );
  OAI21_X1 U20929 ( .B1(n17801), .B2(n17809), .A(n17800), .ZN(n18137) );
  NAND2_X1 U20930 ( .A1(n18781), .A2(n17810), .ZN(n17802) );
  XNOR2_X1 U20931 ( .A(n17802), .B(n17801), .ZN(n18133) );
  AOI22_X1 U20932 ( .A1(n17803), .A2(n18133), .B1(n9846), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17808) );
  AOI22_X1 U20933 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17806), .B1(
        n17805), .B2(n17804), .ZN(n17807) );
  OAI211_X1 U20934 ( .C1(n17815), .C2(n18137), .A(n17808), .B(n17807), .ZN(
        P3_U2829) );
  AOI21_X1 U20935 ( .B1(n17810), .B2(n18781), .A(n17809), .ZN(n18139) );
  INV_X1 U20936 ( .A(n18139), .ZN(n18141) );
  NAND3_X1 U20937 ( .A1(n18763), .A2(n17812), .A3(n17811), .ZN(n17813) );
  AOI22_X1 U20938 ( .A1(n9846), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17813), .ZN(n17814) );
  OAI221_X1 U20939 ( .B1(n18139), .B2(n17816), .C1(n18141), .C2(n17815), .A(
        n17814), .ZN(P3_U2830) );
  INV_X1 U20940 ( .A(n17856), .ZN(n17839) );
  OAI22_X1 U20941 ( .A1(n17818), .A2(n18143), .B1(n17817), .B2(n17839), .ZN(
        n17828) );
  NAND2_X1 U20942 ( .A1(n18130), .A2(n18618), .ZN(n18092) );
  INV_X1 U20943 ( .A(n18092), .ZN(n18113) );
  AOI21_X1 U20944 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18618), .A(
        n17819), .ZN(n17881) );
  OAI21_X1 U20945 ( .B1(n17881), .B2(n17820), .A(n18092), .ZN(n17860) );
  OAI21_X1 U20946 ( .B1(n18113), .B2(n17843), .A(n17860), .ZN(n17840) );
  AOI22_X1 U20947 ( .A1(n18621), .A2(n17845), .B1(n18611), .B2(n17821), .ZN(
        n17823) );
  OAI211_X1 U20948 ( .C1(n17824), .C2(n18794), .A(n17823), .B(n17822), .ZN(
        n17825) );
  AOI211_X1 U20949 ( .C1(n17990), .C2(n17826), .A(n17840), .B(n17825), .ZN(
        n17832) );
  OAI211_X1 U20950 ( .C1(n18130), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n17832), .ZN(n17827) );
  AOI22_X1 U20951 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18121), .B1(
        n17828), .B2(n17827), .ZN(n17830) );
  NAND2_X1 U20952 ( .A1(n9846), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17829) );
  OAI211_X1 U20953 ( .C1(n17831), .C2(n17947), .A(n17830), .B(n17829), .ZN(
        P3_U2835) );
  NOR3_X1 U20954 ( .A1(n17832), .A2(n18143), .A3(n17833), .ZN(n17835) );
  OAI22_X1 U20955 ( .A1(n17833), .A2(n18128), .B1(n18094), .B2(n18731), .ZN(
        n17834) );
  AOI211_X1 U20956 ( .C1(n18057), .C2(n17836), .A(n17835), .B(n17834), .ZN(
        n17837) );
  OAI21_X1 U20957 ( .B1(n17839), .B2(n17838), .A(n17837), .ZN(P3_U2836) );
  AOI221_X1 U20958 ( .B1(n17841), .B2(n18639), .C1(n17862), .C2(n18639), .A(
        n17840), .ZN(n17846) );
  NAND3_X1 U20959 ( .A1(n17843), .A2(n17842), .A3(n17845), .ZN(n17844) );
  OAI21_X1 U20960 ( .B1(n17846), .B2(n17845), .A(n17844), .ZN(n17847) );
  AOI22_X1 U20961 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18121), .B1(
        n18127), .B2(n17847), .ZN(n17849) );
  OAI211_X1 U20962 ( .C1(n17850), .C2(n17947), .A(n17849), .B(n17848), .ZN(
        n17851) );
  AOI21_X1 U20963 ( .B1(n18058), .B2(n17852), .A(n17851), .ZN(n17853) );
  OAI21_X1 U20964 ( .B1(n18125), .B2(n17854), .A(n17853), .ZN(P3_U2837) );
  AOI22_X1 U20965 ( .A1(n18057), .A2(n17857), .B1(n17856), .B2(n17855), .ZN(
        n17866) );
  AOI22_X1 U20966 ( .A1(n17875), .A2(n17859), .B1(n17990), .B2(n17858), .ZN(
        n17861) );
  NAND3_X1 U20967 ( .A1(n17861), .A2(n18128), .A3(n17860), .ZN(n17864) );
  AOI211_X1 U20968 ( .C1(n18639), .C2(n17862), .A(n17867), .B(n17864), .ZN(
        n17863) );
  NOR2_X1 U20969 ( .A1(n9846), .A2(n17863), .ZN(n17870) );
  OAI211_X1 U20970 ( .C1(n18051), .C2(n17864), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17870), .ZN(n17865) );
  OAI211_X1 U20971 ( .C1(n18727), .C2(n18094), .A(n17866), .B(n17865), .ZN(
        P3_U2838) );
  OAI21_X1 U20972 ( .B1(n18121), .B2(n17868), .A(n17867), .ZN(n17869) );
  AOI22_X1 U20973 ( .A1(n18057), .A2(n17871), .B1(n17870), .B2(n17869), .ZN(
        n17873) );
  NAND2_X1 U20974 ( .A1(n17873), .A2(n17872), .ZN(P3_U2839) );
  NAND2_X1 U20975 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17874), .ZN(
        n17882) );
  NOR2_X1 U20976 ( .A1(n17875), .A2(n17990), .ZN(n18019) );
  OAI21_X1 U20977 ( .B1(n17876), .B2(n17894), .A(n18639), .ZN(n17877) );
  OAI221_X1 U20978 ( .B1(n18130), .B2(n17930), .C1(n18130), .C2(n17906), .A(
        n17877), .ZN(n17904) );
  AOI21_X1 U20979 ( .B1(n18621), .B2(n17878), .A(n17904), .ZN(n17879) );
  OAI21_X1 U20980 ( .B1(n17880), .B2(n18019), .A(n17879), .ZN(n17892) );
  AOI211_X1 U20981 ( .C1(n18028), .C2(n17882), .A(n17881), .B(n17892), .ZN(
        n17887) );
  NOR2_X1 U20982 ( .A1(n17883), .A2(n18794), .ZN(n17963) );
  AOI21_X1 U20983 ( .B1(n17990), .B2(n17884), .A(n17963), .ZN(n17909) );
  AOI22_X1 U20984 ( .A1(n17887), .A2(n17909), .B1(n17886), .B2(n17885), .ZN(
        n17888) );
  AOI22_X1 U20985 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18121), .B1(
        n18127), .B2(n17888), .ZN(n17890) );
  NAND2_X1 U20986 ( .A1(n9846), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17889) );
  OAI211_X1 U20987 ( .C1(n17891), .C2(n17947), .A(n17890), .B(n17889), .ZN(
        P3_U2840) );
  NAND2_X1 U20988 ( .A1(n18618), .A2(n18613), .ZN(n18126) );
  NAND2_X1 U20989 ( .A1(n18127), .A2(n17909), .ZN(n17953) );
  AOI211_X1 U20990 ( .C1(n17893), .C2(n18126), .A(n17953), .B(n17892), .ZN(
        n17895) );
  NOR2_X1 U20991 ( .A1(n18781), .A2(n17950), .ZN(n18035) );
  NAND2_X1 U20992 ( .A1(n17929), .A2(n18035), .ZN(n17951) );
  OAI21_X1 U20993 ( .B1(n17894), .B2(n17951), .A(n18611), .ZN(n17905) );
  AOI21_X1 U20994 ( .B1(n17895), .B2(n17905), .A(n9846), .ZN(n17900) );
  INV_X1 U20995 ( .A(n17896), .ZN(n17914) );
  NOR4_X1 U20996 ( .A1(n17914), .A2(n17898), .A3(n17897), .A4(n18143), .ZN(
        n17922) );
  AOI22_X1 U20997 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17900), .B1(
        n17899), .B2(n17922), .ZN(n17902) );
  OAI211_X1 U20998 ( .C1(n17903), .C2(n17947), .A(n17902), .B(n17901), .ZN(
        P3_U2841) );
  NAND3_X1 U20999 ( .A1(n20679), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(n18126), 
        .ZN(n17912) );
  INV_X1 U21000 ( .A(n17904), .ZN(n17910) );
  OAI211_X1 U21001 ( .C1(n17906), .C2(n18019), .A(n18128), .B(n17905), .ZN(
        n17907) );
  INV_X1 U21002 ( .A(n17907), .ZN(n17908) );
  NAND3_X1 U21003 ( .A1(n17910), .A2(n17909), .A3(n17908), .ZN(n17911) );
  NAND2_X1 U21004 ( .A1(n18094), .A2(n17911), .ZN(n17921) );
  NAND2_X1 U21005 ( .A1(n17912), .A2(n17921), .ZN(n17917) );
  INV_X1 U21006 ( .A(n17913), .ZN(n17916) );
  NOR2_X1 U21007 ( .A1(n17914), .A2(n18143), .ZN(n17915) );
  AOI22_X1 U21008 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17917), .B1(
        n17916), .B2(n17915), .ZN(n17919) );
  OAI211_X1 U21009 ( .C1(n17920), .C2(n17947), .A(n17919), .B(n17918), .ZN(
        P3_U2842) );
  NAND2_X1 U21010 ( .A1(n9846), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17925) );
  INV_X1 U21011 ( .A(n17921), .ZN(n17923) );
  AOI22_X1 U21012 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17923), .B1(
        n17922), .B2(n20679), .ZN(n17924) );
  OAI211_X1 U21013 ( .C1(n17926), .C2(n17947), .A(n17925), .B(n17924), .ZN(
        P3_U2843) );
  OAI22_X1 U21014 ( .A1(n18048), .A2(n18613), .B1(n18114), .B2(n18091), .ZN(
        n18101) );
  NAND2_X1 U21015 ( .A1(n18127), .A2(n18101), .ZN(n18089) );
  NOR2_X1 U21016 ( .A1(n17961), .A2(n18089), .ZN(n17999) );
  INV_X1 U21017 ( .A(n17927), .ZN(n17928) );
  AOI22_X1 U21018 ( .A1(n17929), .A2(n17999), .B1(n18127), .B2(n17928), .ZN(
        n17958) );
  NAND2_X1 U21019 ( .A1(n18611), .A2(n18781), .ZN(n18112) );
  NAND3_X1 U21020 ( .A1(n17930), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18112), .ZN(n17934) );
  OAI22_X1 U21021 ( .A1(n17932), .A2(n18019), .B1(n17931), .B2(n18613), .ZN(
        n17933) );
  AOI211_X1 U21022 ( .C1(n18092), .C2(n17934), .A(n17953), .B(n17933), .ZN(
        n17941) );
  AOI221_X1 U21023 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17941), 
        .C1(n18113), .C2(n17941), .A(n9846), .ZN(n17936) );
  AOI22_X1 U21024 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17936), .B1(
        n18057), .B2(n17935), .ZN(n17938) );
  OAI211_X1 U21025 ( .C1(n17958), .C2(n17939), .A(n17938), .B(n17937), .ZN(
        P3_U2844) );
  INV_X1 U21026 ( .A(n17958), .ZN(n17943) );
  INV_X1 U21027 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17940) );
  NOR3_X1 U21028 ( .A1(n9846), .A2(n17941), .A3(n17940), .ZN(n17942) );
  AOI21_X1 U21029 ( .B1(n17944), .B2(n17943), .A(n17942), .ZN(n17946) );
  OAI211_X1 U21030 ( .C1(n17948), .C2(n17947), .A(n17946), .B(n17945), .ZN(
        P3_U2845) );
  NOR2_X1 U21031 ( .A1(n17949), .A2(n18613), .ZN(n18038) );
  AOI21_X1 U21032 ( .B1(n18621), .B2(n17950), .A(n18038), .ZN(n18018) );
  OAI21_X1 U21033 ( .B1(n10208), .B2(n18611), .A(n17951), .ZN(n17952) );
  OAI211_X1 U21034 ( .C1(n18022), .C2(n17959), .A(n18018), .B(n17952), .ZN(
        n17967) );
  OAI221_X1 U21035 ( .B1(n17953), .B2(n18051), .C1(n17953), .C2(n17967), .A(
        n18094), .ZN(n17956) );
  AOI22_X1 U21036 ( .A1(n9846), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18057), 
        .B2(n17954), .ZN(n17955) );
  OAI221_X1 U21037 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17958), 
        .C1(n17957), .C2(n17956), .A(n17955), .ZN(P3_U2846) );
  NAND2_X1 U21038 ( .A1(n17959), .A2(n18101), .ZN(n17960) );
  OAI21_X1 U21039 ( .B1(n17961), .B2(n17960), .A(n10208), .ZN(n17968) );
  NOR2_X1 U21040 ( .A1(n17962), .A2(n18014), .ZN(n17965) );
  AOI222_X1 U21041 ( .A1(n17968), .A2(n17967), .B1(n17966), .B2(n17965), .C1(
        n17964), .C2(n17963), .ZN(n17973) );
  INV_X1 U21042 ( .A(n17969), .ZN(n17970) );
  AOI22_X1 U21043 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18121), .B1(
        n18057), .B2(n17970), .ZN(n17972) );
  OAI211_X1 U21044 ( .C1(n17973), .C2(n18143), .A(n17972), .B(n17971), .ZN(
        P3_U2847) );
  INV_X1 U21045 ( .A(n17974), .ZN(n17978) );
  NOR2_X1 U21046 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17978), .ZN(
        n17983) );
  INV_X1 U21047 ( .A(n18018), .ZN(n17977) );
  AOI21_X1 U21048 ( .B1(n17975), .B2(n18035), .A(n18618), .ZN(n17976) );
  NOR2_X1 U21049 ( .A1(n17977), .A2(n17976), .ZN(n17992) );
  AOI21_X1 U21050 ( .B1(n18051), .B2(n17978), .A(n18143), .ZN(n17980) );
  AOI211_X1 U21051 ( .C1(n17992), .C2(n17980), .A(n9846), .B(n17979), .ZN(
        n17981) );
  AOI211_X1 U21052 ( .C1(n17999), .C2(n17983), .A(n17982), .B(n17981), .ZN(
        n17987) );
  AOI22_X1 U21053 ( .A1(n18058), .A2(n17985), .B1(n18057), .B2(n17984), .ZN(
        n17986) );
  OAI211_X1 U21054 ( .C1(n18125), .C2(n17988), .A(n17987), .B(n17986), .ZN(
        P3_U2848) );
  AOI22_X1 U21055 ( .A1(n17990), .A2(n17989), .B1(n18028), .B2(n18000), .ZN(
        n17991) );
  OAI211_X1 U21056 ( .C1(n17993), .C2(n18794), .A(n17992), .B(n17991), .ZN(
        n18006) );
  OAI21_X1 U21057 ( .B1(n18022), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18127), .ZN(n17994) );
  OAI21_X1 U21058 ( .B1(n18006), .B2(n17994), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18004) );
  OAI22_X1 U21059 ( .A1(n17997), .A2(n18125), .B1(n17996), .B2(n17995), .ZN(
        n17998) );
  NOR2_X1 U21060 ( .A1(n17999), .A2(n17998), .ZN(n18046) );
  NOR2_X1 U21061 ( .A1(n18046), .A2(n18000), .ZN(n18008) );
  AOI22_X1 U21062 ( .A1(n18057), .A2(n18002), .B1(n18001), .B2(n18008), .ZN(
        n18003) );
  OAI221_X1 U21063 ( .B1(n9846), .B2(n18004), .C1(n18094), .C2(n18707), .A(
        n18003), .ZN(P3_U2849) );
  AOI22_X1 U21064 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18121), .B1(
        n18057), .B2(n18005), .ZN(n18010) );
  NOR2_X1 U21065 ( .A1(n18143), .A2(n10209), .ZN(n18007) );
  OAI22_X1 U21066 ( .A1(n18008), .A2(n18007), .B1(n18006), .B2(n10209), .ZN(
        n18009) );
  OAI211_X1 U21067 ( .C1(n18705), .C2(n18094), .A(n18010), .B(n18009), .ZN(
        P3_U2850) );
  INV_X1 U21068 ( .A(n18046), .ZN(n18027) );
  AOI22_X1 U21069 ( .A1(n18057), .A2(n18012), .B1(n18011), .B2(n18027), .ZN(
        n18026) );
  AOI21_X1 U21070 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18035), .A(
        n18618), .ZN(n18016) );
  OAI22_X1 U21071 ( .A1(n18015), .A2(n18014), .B1(n18794), .B2(n18013), .ZN(
        n18036) );
  NOR3_X1 U21072 ( .A1(n18016), .A2(n18036), .A3(n18143), .ZN(n18017) );
  OAI211_X1 U21073 ( .C1(n18020), .C2(n18019), .A(n18018), .B(n18017), .ZN(
        n18029) );
  OAI22_X1 U21074 ( .A1(n18022), .A2(n18021), .B1(n18618), .B2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18023) );
  OAI211_X1 U21075 ( .C1(n18029), .C2(n18023), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18094), .ZN(n18024) );
  NAND3_X1 U21076 ( .A1(n18026), .A2(n18025), .A3(n18024), .ZN(P3_U2851) );
  NAND2_X1 U21077 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18027), .ZN(
        n18034) );
  INV_X1 U21078 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18033) );
  OAI221_X1 U21079 ( .B1(n18029), .B2(n18028), .C1(n18029), .C2(n18045), .A(
        n18094), .ZN(n18032) );
  AOI22_X1 U21080 ( .A1(n9846), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18057), 
        .B2(n18030), .ZN(n18031) );
  OAI221_X1 U21081 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n18034), 
        .C1(n18033), .C2(n18032), .A(n18031), .ZN(P3_U2852) );
  AOI211_X1 U21082 ( .C1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n18618), .A(
        n18113), .B(n18035), .ZN(n18037) );
  OR4_X1 U21083 ( .A1(n18121), .A2(n18038), .A3(n18037), .A4(n18036), .ZN(
        n18040) );
  OAI221_X1 U21084 ( .B1(n18040), .B2(n18621), .C1(n18040), .C2(n18039), .A(
        n18094), .ZN(n18044) );
  AOI21_X1 U21085 ( .B1(n18057), .B2(n18042), .A(n18041), .ZN(n18043) );
  OAI221_X1 U21086 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18046), .C1(
        n18045), .C2(n18044), .A(n18043), .ZN(P3_U2853) );
  NAND2_X1 U21087 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18047) );
  NOR3_X1 U21088 ( .A1(n18072), .A2(n18047), .A3(n18089), .ZN(n18055) );
  INV_X1 U21089 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18077) );
  NAND2_X1 U21090 ( .A1(n18639), .A2(n18048), .ZN(n18117) );
  NAND2_X1 U21091 ( .A1(n18112), .A2(n18117), .ZN(n18090) );
  AOI21_X1 U21092 ( .B1(n18639), .B2(n18072), .A(n18090), .ZN(n18049) );
  OAI21_X1 U21093 ( .B1(n18113), .B2(n18050), .A(n18049), .ZN(n18073) );
  AOI211_X1 U21094 ( .C1(n18051), .C2(n18077), .A(n20725), .B(n18073), .ZN(
        n18064) );
  OAI21_X1 U21095 ( .B1(n18064), .B2(n18129), .A(n18128), .ZN(n18053) );
  NOR2_X1 U21096 ( .A1(n18094), .A2(n18698), .ZN(n18052) );
  AOI221_X1 U21097 ( .B1(n18055), .B2(n18054), .C1(n18053), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18052), .ZN(n18061) );
  AOI22_X1 U21098 ( .A1(n18059), .A2(n18058), .B1(n18057), .B2(n18056), .ZN(
        n18060) );
  OAI211_X1 U21099 ( .C1(n18125), .C2(n18062), .A(n18061), .B(n18060), .ZN(
        P3_U2854) );
  INV_X1 U21100 ( .A(n18140), .ZN(n18136) );
  NAND3_X1 U21101 ( .A1(n18063), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n18101), .ZN(n18065) );
  AOI211_X1 U21102 ( .C1(n20725), .C2(n18065), .A(n18064), .B(n18143), .ZN(
        n18066) );
  AOI211_X1 U21103 ( .C1(n18121), .C2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18067), .B(n18066), .ZN(n18070) );
  NAND2_X1 U21104 ( .A1(n18142), .A2(n18068), .ZN(n18069) );
  OAI211_X1 U21105 ( .C1(n18071), .C2(n18136), .A(n18070), .B(n18069), .ZN(
        P3_U2855) );
  NOR2_X1 U21106 ( .A1(n18072), .A2(n18089), .ZN(n18078) );
  AOI21_X1 U21107 ( .B1(n18073), .B2(n18127), .A(n18121), .ZN(n18074) );
  INV_X1 U21108 ( .A(n18074), .ZN(n18084) );
  OAI22_X1 U21109 ( .A1(n18094), .A2(n18694), .B1(n18136), .B2(n18075), .ZN(
        n18076) );
  AOI221_X1 U21110 ( .B1(n18078), .B2(n18077), .C1(n18084), .C2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n18076), .ZN(n18079) );
  OAI21_X1 U21111 ( .B1(n18125), .B2(n18080), .A(n18079), .ZN(P3_U2856) );
  NOR3_X1 U21112 ( .A1(n18110), .A2(n18097), .A3(n18089), .ZN(n18086) );
  OAI21_X1 U21113 ( .B1(n18136), .B2(n18082), .A(n18081), .ZN(n18083) );
  AOI221_X1 U21114 ( .B1(n18086), .B2(n18085), .C1(n18084), .C2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n18083), .ZN(n18087) );
  OAI21_X1 U21115 ( .B1(n18125), .B2(n18088), .A(n18087), .ZN(P3_U2857) );
  NOR2_X1 U21116 ( .A1(n18110), .A2(n18089), .ZN(n18098) );
  AOI211_X1 U21117 ( .C1(n18092), .C2(n18091), .A(n18110), .B(n18090), .ZN(
        n18102) );
  OAI21_X1 U21118 ( .B1(n18102), .B2(n18129), .A(n18128), .ZN(n18096) );
  OAI22_X1 U21119 ( .A1(n18094), .A2(n18690), .B1(n18136), .B2(n18093), .ZN(
        n18095) );
  AOI221_X1 U21120 ( .B1(n18098), .B2(n18097), .C1(n18096), .C2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n18095), .ZN(n18099) );
  OAI21_X1 U21121 ( .B1(n18125), .B2(n18100), .A(n18099), .ZN(P3_U2858) );
  INV_X1 U21122 ( .A(n18101), .ZN(n18103) );
  AOI211_X1 U21123 ( .C1(n18103), .C2(n18110), .A(n18102), .B(n18143), .ZN(
        n18107) );
  OAI22_X1 U21124 ( .A1(n18136), .A2(n18105), .B1(n18125), .B2(n18104), .ZN(
        n18106) );
  NOR2_X1 U21125 ( .A1(n18107), .A2(n18106), .ZN(n18109) );
  OAI211_X1 U21126 ( .C1(n18128), .C2(n18110), .A(n18109), .B(n18108), .ZN(
        P3_U2859) );
  NAND3_X1 U21127 ( .A1(n18639), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18111) );
  OAI211_X1 U21128 ( .C1(n18113), .C2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n18112), .B(n18111), .ZN(n18116) );
  NOR2_X1 U21129 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18114), .ZN(
        n18115) );
  AOI22_X1 U21130 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18116), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18115), .ZN(n18118) );
  OAI211_X1 U21131 ( .C1(n18796), .C2(n18119), .A(n18118), .B(n18117), .ZN(
        n18120) );
  AOI22_X1 U21132 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18121), .B1(
        n18127), .B2(n18120), .ZN(n18123) );
  OAI211_X1 U21133 ( .C1(n18125), .C2(n18124), .A(n18123), .B(n18122), .ZN(
        P3_U2860) );
  NAND3_X1 U21134 ( .A1(n18127), .A2(n18781), .A3(n18126), .ZN(n18145) );
  INV_X1 U21135 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18761) );
  AOI21_X1 U21136 ( .B1(n18128), .B2(n18145), .A(n18761), .ZN(n18132) );
  AOI211_X1 U21137 ( .C1(n18130), .C2(n18781), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18129), .ZN(n18131) );
  AOI211_X1 U21138 ( .C1(n18142), .C2(n18133), .A(n18132), .B(n18131), .ZN(
        n18135) );
  NAND2_X1 U21139 ( .A1(n9846), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18134) );
  OAI211_X1 U21140 ( .C1(n18137), .C2(n18136), .A(n18135), .B(n18134), .ZN(
        P3_U2861) );
  AND2_X1 U21141 ( .A1(n9846), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18138) );
  AOI221_X1 U21142 ( .B1(n18142), .B2(n18141), .C1(n18140), .C2(n18139), .A(
        n18138), .ZN(n18146) );
  OAI211_X1 U21143 ( .C1(n18621), .C2(n18143), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n18094), .ZN(n18144) );
  NAND3_X1 U21144 ( .A1(n18146), .A2(n18145), .A3(n18144), .ZN(P3_U2862) );
  AOI21_X1 U21145 ( .B1(n18149), .B2(n18148), .A(n18147), .ZN(n18655) );
  OAI21_X1 U21146 ( .B1(n18655), .B2(n18209), .A(n18151), .ZN(n18150) );
  OAI221_X1 U21147 ( .B1(n18622), .B2(n18811), .C1(n18622), .C2(n18151), .A(
        n18150), .ZN(P3_U2863) );
  NAND2_X1 U21148 ( .A1(n18644), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18298) );
  INV_X1 U21149 ( .A(n18298), .ZN(n18345) );
  NAND2_X1 U21150 ( .A1(n18156), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18410) );
  INV_X1 U21151 ( .A(n18410), .ZN(n18390) );
  NOR2_X1 U21152 ( .A1(n18345), .A2(n18390), .ZN(n18153) );
  OAI22_X1 U21153 ( .A1(n18154), .A2(n18644), .B1(n18153), .B2(n18152), .ZN(
        P3_U2866) );
  AND2_X1 U21154 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18155), .ZN(
        P3_U2867) );
  NOR2_X1 U21155 ( .A1(n18644), .A2(n18319), .ZN(n18543) );
  NAND2_X1 U21156 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18543), .ZN(
        n18597) );
  INV_X1 U21157 ( .A(n18597), .ZN(n18570) );
  NOR2_X1 U21158 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18210) );
  NOR2_X1 U21159 ( .A1(n18570), .A2(n18261), .ZN(n18233) );
  AOI21_X1 U21160 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18509), .ZN(n18321) );
  INV_X1 U21161 ( .A(n18321), .ZN(n18158) );
  NAND2_X1 U21162 ( .A1(n18623), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18389) );
  INV_X1 U21163 ( .A(n18389), .ZN(n18157) );
  NOR2_X1 U21164 ( .A1(n18156), .A2(n18644), .ZN(n18482) );
  NAND2_X1 U21165 ( .A1(n18157), .A2(n18482), .ZN(n18499) );
  INV_X1 U21166 ( .A(n18499), .ZN(n18592) );
  NAND2_X1 U21167 ( .A1(n18622), .A2(n18543), .ZN(n18537) );
  INV_X1 U21168 ( .A(n18537), .ZN(n18512) );
  NOR2_X1 U21169 ( .A1(n18592), .A2(n18512), .ZN(n18510) );
  OAI22_X1 U21170 ( .A1(n18233), .A2(n18158), .B1(n18510), .B2(n18507), .ZN(
        n18208) );
  NAND2_X1 U21171 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18545), .ZN(n18549) );
  INV_X1 U21172 ( .A(n18549), .ZN(n18506) );
  AND2_X1 U21173 ( .A1(n18414), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18540) );
  NOR2_X1 U21174 ( .A1(n18539), .A2(n18233), .ZN(n18202) );
  AOI22_X1 U21175 ( .A1(n18506), .A2(n18592), .B1(n18540), .B2(n18202), .ZN(
        n18163) );
  NOR2_X1 U21176 ( .A1(n18160), .A2(n18159), .ZN(n18203) );
  NAND2_X1 U21177 ( .A1(n18161), .A2(n18203), .ZN(n18515) );
  INV_X1 U21178 ( .A(n18515), .ZN(n18546) );
  INV_X1 U21179 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n19093) );
  NOR2_X2 U21180 ( .A1(n18507), .A2(n19093), .ZN(n18541) );
  AOI22_X1 U21181 ( .A1(n18546), .A2(n18261), .B1(n18541), .B2(n18512), .ZN(
        n18162) );
  OAI211_X1 U21182 ( .C1(n18164), .C2(n18208), .A(n18163), .B(n18162), .ZN(
        P3_U2868) );
  NOR2_X2 U21183 ( .A1(n18509), .A2(n18165), .ZN(n18550) );
  AND2_X1 U21184 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18545), .ZN(n18552) );
  AOI22_X1 U21185 ( .A1(n18550), .A2(n18202), .B1(n18552), .B2(n18592), .ZN(
        n18169) );
  INV_X1 U21186 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n18166) );
  NOR2_X2 U21187 ( .A1(n18507), .A2(n18166), .ZN(n18551) );
  INV_X1 U21188 ( .A(n18203), .ZN(n18196) );
  NOR2_X1 U21189 ( .A1(n18196), .A2(n18167), .ZN(n18213) );
  AOI22_X1 U21190 ( .A1(n18551), .A2(n18512), .B1(n18213), .B2(n18261), .ZN(
        n18168) );
  OAI211_X1 U21191 ( .C1(n18170), .C2(n18208), .A(n18169), .B(n18168), .ZN(
        P3_U2869) );
  NOR2_X1 U21192 ( .A1(n19102), .A2(n18507), .ZN(n18518) );
  NOR2_X2 U21193 ( .A1(n18509), .A2(n18171), .ZN(n18556) );
  AOI22_X1 U21194 ( .A1(n18518), .A2(n18592), .B1(n18556), .B2(n18202), .ZN(
        n18175) );
  NAND2_X1 U21195 ( .A1(n18172), .A2(n18203), .ZN(n18521) );
  INV_X1 U21196 ( .A(n18521), .ZN(n18558) );
  INV_X1 U21197 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n18173) );
  NOR2_X2 U21198 ( .A1(n18507), .A2(n18173), .ZN(n18557) );
  AOI22_X1 U21199 ( .A1(n18558), .A2(n18261), .B1(n18557), .B2(n18512), .ZN(
        n18174) );
  OAI211_X1 U21200 ( .C1(n18176), .C2(n18208), .A(n18175), .B(n18174), .ZN(
        P3_U2870) );
  NOR2_X2 U21201 ( .A1(n20785), .A2(n18507), .ZN(n18563) );
  NOR2_X2 U21202 ( .A1(n18509), .A2(n18177), .ZN(n18562) );
  AOI22_X1 U21203 ( .A1(n18563), .A2(n18592), .B1(n18562), .B2(n18202), .ZN(
        n18181) );
  INV_X1 U21204 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n18178) );
  NOR2_X2 U21205 ( .A1(n18507), .A2(n18178), .ZN(n18564) );
  NOR2_X1 U21206 ( .A1(n18196), .A2(n18179), .ZN(n18218) );
  AOI22_X1 U21207 ( .A1(n18564), .A2(n18512), .B1(n18218), .B2(n18261), .ZN(
        n18180) );
  OAI211_X1 U21208 ( .C1(n18182), .C2(n18208), .A(n18181), .B(n18180), .ZN(
        P3_U2871) );
  NOR2_X2 U21209 ( .A1(n18183), .A2(n18507), .ZN(n18524) );
  NOR2_X2 U21210 ( .A1(n18509), .A2(n18184), .ZN(n18569) );
  AOI22_X1 U21211 ( .A1(n18524), .A2(n18592), .B1(n18569), .B2(n18202), .ZN(
        n18187) );
  NAND2_X1 U21212 ( .A1(n18185), .A2(n18203), .ZN(n18527) );
  INV_X1 U21213 ( .A(n18527), .ZN(n18571) );
  INV_X1 U21214 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n20687) );
  NOR2_X2 U21215 ( .A1(n18507), .A2(n20687), .ZN(n18568) );
  AOI22_X1 U21216 ( .A1(n18571), .A2(n18261), .B1(n18568), .B2(n18512), .ZN(
        n18186) );
  OAI211_X1 U21217 ( .C1(n18188), .C2(n18208), .A(n18187), .B(n18186), .ZN(
        P3_U2872) );
  NOR2_X2 U21218 ( .A1(n18507), .A2(n18189), .ZN(n18578) );
  NOR2_X2 U21219 ( .A1(n18509), .A2(n18190), .ZN(n18576) );
  AOI22_X1 U21220 ( .A1(n18578), .A2(n18512), .B1(n18576), .B2(n18202), .ZN(
        n18193) );
  NOR2_X1 U21221 ( .A1(n18196), .A2(n18191), .ZN(n18223) );
  AND2_X1 U21222 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18545), .ZN(n18577) );
  AOI22_X1 U21223 ( .A1(n18223), .A2(n18261), .B1(n18577), .B2(n18592), .ZN(
        n18192) );
  OAI211_X1 U21224 ( .C1(n18194), .C2(n18208), .A(n18193), .B(n18192), .ZN(
        P3_U2873) );
  NOR2_X2 U21225 ( .A1(n12676), .A2(n18507), .ZN(n18584) );
  NOR2_X2 U21226 ( .A1(n18509), .A2(n20806), .ZN(n18582) );
  AOI22_X1 U21227 ( .A1(n18584), .A2(n18592), .B1(n18582), .B2(n18202), .ZN(
        n18198) );
  AND2_X1 U21228 ( .A1(n18545), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18583) );
  NOR2_X1 U21229 ( .A1(n18196), .A2(n18195), .ZN(n18226) );
  AOI22_X1 U21230 ( .A1(n18583), .A2(n18512), .B1(n18226), .B2(n18261), .ZN(
        n18197) );
  OAI211_X1 U21231 ( .C1(n18199), .C2(n18208), .A(n18198), .B(n18197), .ZN(
        P3_U2874) );
  NOR2_X2 U21232 ( .A1(n18507), .A2(n18200), .ZN(n18591) );
  NOR2_X2 U21233 ( .A1(n18201), .A2(n18509), .ZN(n18589) );
  AOI22_X1 U21234 ( .A1(n18591), .A2(n18592), .B1(n18589), .B2(n18202), .ZN(
        n18207) );
  NAND2_X1 U21235 ( .A1(n18204), .A2(n18203), .ZN(n18598) );
  INV_X1 U21236 ( .A(n18598), .ZN(n18500) );
  INV_X1 U21237 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n18205) );
  NOR2_X2 U21238 ( .A1(n18205), .A2(n18507), .ZN(n18593) );
  AOI22_X1 U21239 ( .A1(n18500), .A2(n18261), .B1(n18593), .B2(n18512), .ZN(
        n18206) );
  OAI211_X1 U21240 ( .C1(n20823), .C2(n18208), .A(n18207), .B(n18206), .ZN(
        P3_U2875) );
  NOR2_X2 U21241 ( .A1(n18389), .A2(n18253), .ZN(n18292) );
  NAND2_X1 U21242 ( .A1(n18623), .A2(n18435), .ZN(n18479) );
  NOR2_X1 U21243 ( .A1(n18253), .A2(n18479), .ZN(n18229) );
  AOI22_X1 U21244 ( .A1(n18506), .A2(n18512), .B1(n18540), .B2(n18229), .ZN(
        n18212) );
  NOR2_X1 U21245 ( .A1(n18509), .A2(n18209), .ZN(n18542) );
  AND2_X1 U21246 ( .A1(n18623), .A2(n18542), .ZN(n18481) );
  AOI22_X1 U21247 ( .A1(n18545), .A2(n18543), .B1(n18210), .B2(n18481), .ZN(
        n18230) );
  AOI22_X1 U21248 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18230), .B1(
        n18541), .B2(n18570), .ZN(n18211) );
  OAI211_X1 U21249 ( .C1(n18515), .C2(n18282), .A(n18212), .B(n18211), .ZN(
        P3_U2876) );
  AOI22_X1 U21250 ( .A1(n18551), .A2(n18570), .B1(n18550), .B2(n18229), .ZN(
        n18215) );
  AOI22_X1 U21251 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18230), .B1(
        n18552), .B2(n18512), .ZN(n18214) );
  OAI211_X1 U21252 ( .C1(n18555), .C2(n18282), .A(n18215), .B(n18214), .ZN(
        P3_U2877) );
  AOI22_X1 U21253 ( .A1(n18557), .A2(n18570), .B1(n18556), .B2(n18229), .ZN(
        n18217) );
  AOI22_X1 U21254 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18230), .B1(
        n18518), .B2(n18512), .ZN(n18216) );
  OAI211_X1 U21255 ( .C1(n18521), .C2(n18282), .A(n18217), .B(n18216), .ZN(
        P3_U2878) );
  INV_X1 U21256 ( .A(n18218), .ZN(n18567) );
  AOI22_X1 U21257 ( .A1(n18563), .A2(n18512), .B1(n18562), .B2(n18229), .ZN(
        n18220) );
  AOI22_X1 U21258 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18230), .B1(
        n18564), .B2(n18570), .ZN(n18219) );
  OAI211_X1 U21259 ( .C1(n18567), .C2(n18282), .A(n18220), .B(n18219), .ZN(
        P3_U2879) );
  AOI22_X1 U21260 ( .A1(n18524), .A2(n18512), .B1(n18569), .B2(n18229), .ZN(
        n18222) );
  AOI22_X1 U21261 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18230), .B1(
        n18568), .B2(n18570), .ZN(n18221) );
  OAI211_X1 U21262 ( .C1(n18527), .C2(n18282), .A(n18222), .B(n18221), .ZN(
        P3_U2880) );
  AOI22_X1 U21263 ( .A1(n18578), .A2(n18570), .B1(n18576), .B2(n18229), .ZN(
        n18225) );
  AOI22_X1 U21264 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18230), .B1(
        n18577), .B2(n18512), .ZN(n18224) );
  OAI211_X1 U21265 ( .C1(n18581), .C2(n18282), .A(n18225), .B(n18224), .ZN(
        P3_U2881) );
  INV_X1 U21266 ( .A(n18226), .ZN(n18587) );
  AOI22_X1 U21267 ( .A1(n18584), .A2(n18512), .B1(n18582), .B2(n18229), .ZN(
        n18228) );
  AOI22_X1 U21268 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18230), .B1(
        n18583), .B2(n18570), .ZN(n18227) );
  OAI211_X1 U21269 ( .C1(n18587), .C2(n18282), .A(n18228), .B(n18227), .ZN(
        P3_U2882) );
  AOI22_X1 U21270 ( .A1(n18593), .A2(n18570), .B1(n18589), .B2(n18229), .ZN(
        n18232) );
  AOI22_X1 U21271 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18230), .B1(
        n18591), .B2(n18512), .ZN(n18231) );
  OAI211_X1 U21272 ( .C1(n18598), .C2(n18282), .A(n18232), .B(n18231), .ZN(
        P3_U2883) );
  NOR2_X1 U21273 ( .A1(n18623), .A2(n18253), .ZN(n18297) );
  NAND2_X1 U21274 ( .A1(n18297), .A2(n18622), .ZN(n18305) );
  INV_X1 U21275 ( .A(n18305), .ZN(n18315) );
  NOR2_X1 U21276 ( .A1(n18292), .A2(n18315), .ZN(n18274) );
  NOR2_X1 U21277 ( .A1(n18539), .A2(n18274), .ZN(n18249) );
  AOI22_X1 U21278 ( .A1(n18541), .A2(n18261), .B1(n18540), .B2(n18249), .ZN(
        n18236) );
  OAI21_X1 U21279 ( .B1(n18233), .B2(n18411), .A(n18274), .ZN(n18234) );
  OAI211_X1 U21280 ( .C1(n18315), .C2(n18752), .A(n18414), .B(n18234), .ZN(
        n18250) );
  AOI22_X1 U21281 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18250), .B1(
        n18506), .B2(n18570), .ZN(n18235) );
  OAI211_X1 U21282 ( .C1(n18515), .C2(n18305), .A(n18236), .B(n18235), .ZN(
        P3_U2884) );
  AOI22_X1 U21283 ( .A1(n18550), .A2(n18249), .B1(n18552), .B2(n18570), .ZN(
        n18238) );
  AOI22_X1 U21284 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18250), .B1(
        n18551), .B2(n18261), .ZN(n18237) );
  OAI211_X1 U21285 ( .C1(n18555), .C2(n18305), .A(n18238), .B(n18237), .ZN(
        P3_U2885) );
  AOI22_X1 U21286 ( .A1(n18518), .A2(n18570), .B1(n18556), .B2(n18249), .ZN(
        n18240) );
  AOI22_X1 U21287 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18250), .B1(
        n18557), .B2(n18261), .ZN(n18239) );
  OAI211_X1 U21288 ( .C1(n18521), .C2(n18305), .A(n18240), .B(n18239), .ZN(
        P3_U2886) );
  AOI22_X1 U21289 ( .A1(n18563), .A2(n18570), .B1(n18562), .B2(n18249), .ZN(
        n18242) );
  AOI22_X1 U21290 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18250), .B1(
        n18564), .B2(n18261), .ZN(n18241) );
  OAI211_X1 U21291 ( .C1(n18567), .C2(n18305), .A(n18242), .B(n18241), .ZN(
        P3_U2887) );
  AOI22_X1 U21292 ( .A1(n18524), .A2(n18570), .B1(n18569), .B2(n18249), .ZN(
        n18244) );
  AOI22_X1 U21293 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18250), .B1(
        n18568), .B2(n18261), .ZN(n18243) );
  OAI211_X1 U21294 ( .C1(n18527), .C2(n18305), .A(n18244), .B(n18243), .ZN(
        P3_U2888) );
  AOI22_X1 U21295 ( .A1(n18577), .A2(n18570), .B1(n18576), .B2(n18249), .ZN(
        n18246) );
  AOI22_X1 U21296 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18250), .B1(
        n18578), .B2(n18261), .ZN(n18245) );
  OAI211_X1 U21297 ( .C1(n18581), .C2(n18305), .A(n18246), .B(n18245), .ZN(
        P3_U2889) );
  AOI22_X1 U21298 ( .A1(n18583), .A2(n18261), .B1(n18582), .B2(n18249), .ZN(
        n18248) );
  AOI22_X1 U21299 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18250), .B1(
        n18584), .B2(n18570), .ZN(n18247) );
  OAI211_X1 U21300 ( .C1(n18587), .C2(n18305), .A(n18248), .B(n18247), .ZN(
        P3_U2890) );
  AOI22_X1 U21301 ( .A1(n18593), .A2(n18261), .B1(n18589), .B2(n18249), .ZN(
        n18252) );
  AOI22_X1 U21302 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18250), .B1(
        n18591), .B2(n18570), .ZN(n18251) );
  OAI211_X1 U21303 ( .C1(n18598), .C2(n18305), .A(n18252), .B(n18251), .ZN(
        P3_U2891) );
  AND2_X1 U21304 ( .A1(n18435), .A2(n18297), .ZN(n18270) );
  AOI22_X1 U21305 ( .A1(n18541), .A2(n18292), .B1(n18540), .B2(n18270), .ZN(
        n18256) );
  OAI21_X1 U21306 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18253), .A(n18343), 
        .ZN(n18254) );
  NAND3_X1 U21307 ( .A1(n18414), .A2(n18344), .A3(n18254), .ZN(n18271) );
  AOI22_X1 U21308 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18271), .B1(
        n18506), .B2(n18261), .ZN(n18255) );
  OAI211_X1 U21309 ( .C1(n18515), .C2(n18343), .A(n18256), .B(n18255), .ZN(
        P3_U2892) );
  AOI22_X1 U21310 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18271), .B1(
        n18550), .B2(n18270), .ZN(n18258) );
  AOI22_X1 U21311 ( .A1(n18551), .A2(n18292), .B1(n18552), .B2(n18261), .ZN(
        n18257) );
  OAI211_X1 U21312 ( .C1(n18555), .C2(n18343), .A(n18258), .B(n18257), .ZN(
        P3_U2893) );
  AOI22_X1 U21313 ( .A1(n18557), .A2(n18292), .B1(n18556), .B2(n18270), .ZN(
        n18260) );
  AOI22_X1 U21314 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18271), .B1(
        n18518), .B2(n18261), .ZN(n18259) );
  OAI211_X1 U21315 ( .C1(n18521), .C2(n18343), .A(n18260), .B(n18259), .ZN(
        P3_U2894) );
  AOI22_X1 U21316 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18271), .B1(
        n18562), .B2(n18270), .ZN(n18263) );
  AOI22_X1 U21317 ( .A1(n18564), .A2(n18292), .B1(n18563), .B2(n18261), .ZN(
        n18262) );
  OAI211_X1 U21318 ( .C1(n18567), .C2(n18343), .A(n18263), .B(n18262), .ZN(
        P3_U2895) );
  AOI22_X1 U21319 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18271), .B1(
        n18569), .B2(n18270), .ZN(n18265) );
  AOI22_X1 U21320 ( .A1(n18524), .A2(n18261), .B1(n18568), .B2(n18292), .ZN(
        n18264) );
  OAI211_X1 U21321 ( .C1(n18527), .C2(n18343), .A(n18265), .B(n18264), .ZN(
        P3_U2896) );
  AOI22_X1 U21322 ( .A1(n18577), .A2(n18261), .B1(n18576), .B2(n18270), .ZN(
        n18267) );
  AOI22_X1 U21323 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18271), .B1(
        n18578), .B2(n18292), .ZN(n18266) );
  OAI211_X1 U21324 ( .C1(n18581), .C2(n18343), .A(n18267), .B(n18266), .ZN(
        P3_U2897) );
  AOI22_X1 U21325 ( .A1(n18583), .A2(n18292), .B1(n18582), .B2(n18270), .ZN(
        n18269) );
  AOI22_X1 U21326 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18271), .B1(
        n18584), .B2(n18261), .ZN(n18268) );
  OAI211_X1 U21327 ( .C1(n18587), .C2(n18343), .A(n18269), .B(n18268), .ZN(
        P3_U2898) );
  AOI22_X1 U21328 ( .A1(n18591), .A2(n18261), .B1(n18589), .B2(n18270), .ZN(
        n18273) );
  AOI22_X1 U21329 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18271), .B1(
        n18593), .B2(n18292), .ZN(n18272) );
  OAI211_X1 U21330 ( .C1(n18598), .C2(n18343), .A(n18273), .B(n18272), .ZN(
        P3_U2899) );
  NAND2_X1 U21331 ( .A1(n18627), .A2(n18345), .ZN(n18296) );
  NOR2_X1 U21332 ( .A1(n18335), .A2(n18363), .ZN(n18320) );
  NOR2_X1 U21333 ( .A1(n18539), .A2(n18320), .ZN(n18291) );
  AOI22_X1 U21334 ( .A1(n18506), .A2(n18292), .B1(n18540), .B2(n18291), .ZN(
        n18277) );
  OAI21_X1 U21335 ( .B1(n18274), .B2(n18411), .A(n18320), .ZN(n18275) );
  OAI211_X1 U21336 ( .C1(n18363), .C2(n18752), .A(n18414), .B(n18275), .ZN(
        n18293) );
  AOI22_X1 U21337 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18293), .B1(
        n18541), .B2(n18315), .ZN(n18276) );
  OAI211_X1 U21338 ( .C1(n18515), .C2(n18296), .A(n18277), .B(n18276), .ZN(
        P3_U2900) );
  AOI22_X1 U21339 ( .A1(n18550), .A2(n18291), .B1(n18552), .B2(n18292), .ZN(
        n18279) );
  AOI22_X1 U21340 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18293), .B1(
        n18551), .B2(n18315), .ZN(n18278) );
  OAI211_X1 U21341 ( .C1(n18555), .C2(n18296), .A(n18279), .B(n18278), .ZN(
        P3_U2901) );
  INV_X1 U21342 ( .A(n18518), .ZN(n18561) );
  AOI22_X1 U21343 ( .A1(n18557), .A2(n18315), .B1(n18556), .B2(n18291), .ZN(
        n18281) );
  AOI22_X1 U21344 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18293), .B1(
        n18558), .B2(n18363), .ZN(n18280) );
  OAI211_X1 U21345 ( .C1(n18561), .C2(n18282), .A(n18281), .B(n18280), .ZN(
        P3_U2902) );
  AOI22_X1 U21346 ( .A1(n18564), .A2(n18315), .B1(n18562), .B2(n18291), .ZN(
        n18284) );
  AOI22_X1 U21347 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18293), .B1(
        n18563), .B2(n18292), .ZN(n18283) );
  OAI211_X1 U21348 ( .C1(n18567), .C2(n18296), .A(n18284), .B(n18283), .ZN(
        P3_U2903) );
  AOI22_X1 U21349 ( .A1(n18524), .A2(n18292), .B1(n18569), .B2(n18291), .ZN(
        n18286) );
  AOI22_X1 U21350 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18293), .B1(
        n18568), .B2(n18315), .ZN(n18285) );
  OAI211_X1 U21351 ( .C1(n18527), .C2(n18296), .A(n18286), .B(n18285), .ZN(
        P3_U2904) );
  AOI22_X1 U21352 ( .A1(n18578), .A2(n18315), .B1(n18576), .B2(n18291), .ZN(
        n18288) );
  AOI22_X1 U21353 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18293), .B1(
        n18577), .B2(n18292), .ZN(n18287) );
  OAI211_X1 U21354 ( .C1(n18581), .C2(n18296), .A(n18288), .B(n18287), .ZN(
        P3_U2905) );
  AOI22_X1 U21355 ( .A1(n18584), .A2(n18292), .B1(n18582), .B2(n18291), .ZN(
        n18290) );
  AOI22_X1 U21356 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18293), .B1(
        n18583), .B2(n18315), .ZN(n18289) );
  OAI211_X1 U21357 ( .C1(n18587), .C2(n18296), .A(n18290), .B(n18289), .ZN(
        P3_U2906) );
  AOI22_X1 U21358 ( .A1(n18591), .A2(n18292), .B1(n18589), .B2(n18291), .ZN(
        n18295) );
  AOI22_X1 U21359 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18293), .B1(
        n18593), .B2(n18315), .ZN(n18294) );
  OAI211_X1 U21360 ( .C1(n18598), .C2(n18296), .A(n18295), .B(n18294), .ZN(
        P3_U2907) );
  NOR2_X1 U21361 ( .A1(n18298), .A2(n18479), .ZN(n18314) );
  AOI22_X1 U21362 ( .A1(n18541), .A2(n18335), .B1(n18540), .B2(n18314), .ZN(
        n18300) );
  AOI22_X1 U21363 ( .A1(n18545), .A2(n18297), .B1(n18345), .B2(n18481), .ZN(
        n18316) );
  NOR2_X2 U21364 ( .A1(n18389), .A2(n18298), .ZN(n18380) );
  AOI22_X1 U21365 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18316), .B1(
        n18380), .B2(n18546), .ZN(n18299) );
  OAI211_X1 U21366 ( .C1(n18549), .C2(n18305), .A(n18300), .B(n18299), .ZN(
        P3_U2908) );
  AOI22_X1 U21367 ( .A1(n18551), .A2(n18335), .B1(n18550), .B2(n18314), .ZN(
        n18302) );
  AOI22_X1 U21368 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18316), .B1(
        n18552), .B2(n18315), .ZN(n18301) );
  OAI211_X1 U21369 ( .C1(n18388), .C2(n18555), .A(n18302), .B(n18301), .ZN(
        P3_U2909) );
  AOI22_X1 U21370 ( .A1(n18557), .A2(n18335), .B1(n18556), .B2(n18314), .ZN(
        n18304) );
  AOI22_X1 U21371 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18316), .B1(
        n18380), .B2(n18558), .ZN(n18303) );
  OAI211_X1 U21372 ( .C1(n18561), .C2(n18305), .A(n18304), .B(n18303), .ZN(
        P3_U2910) );
  AOI22_X1 U21373 ( .A1(n18563), .A2(n18315), .B1(n18562), .B2(n18314), .ZN(
        n18307) );
  AOI22_X1 U21374 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18316), .B1(
        n18564), .B2(n18335), .ZN(n18306) );
  OAI211_X1 U21375 ( .C1(n18388), .C2(n18567), .A(n18307), .B(n18306), .ZN(
        P3_U2911) );
  AOI22_X1 U21376 ( .A1(n18524), .A2(n18315), .B1(n18569), .B2(n18314), .ZN(
        n18309) );
  AOI22_X1 U21377 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18316), .B1(
        n18568), .B2(n18335), .ZN(n18308) );
  OAI211_X1 U21378 ( .C1(n18388), .C2(n18527), .A(n18309), .B(n18308), .ZN(
        P3_U2912) );
  AOI22_X1 U21379 ( .A1(n18578), .A2(n18335), .B1(n18576), .B2(n18314), .ZN(
        n18311) );
  AOI22_X1 U21380 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18316), .B1(
        n18577), .B2(n18315), .ZN(n18310) );
  OAI211_X1 U21381 ( .C1(n18388), .C2(n18581), .A(n18311), .B(n18310), .ZN(
        P3_U2913) );
  AOI22_X1 U21382 ( .A1(n18584), .A2(n18315), .B1(n18582), .B2(n18314), .ZN(
        n18313) );
  AOI22_X1 U21383 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18316), .B1(
        n18583), .B2(n18335), .ZN(n18312) );
  OAI211_X1 U21384 ( .C1(n18388), .C2(n18587), .A(n18313), .B(n18312), .ZN(
        P3_U2914) );
  AOI22_X1 U21385 ( .A1(n18591), .A2(n18315), .B1(n18589), .B2(n18314), .ZN(
        n18318) );
  AOI22_X1 U21386 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18316), .B1(
        n18593), .B2(n18335), .ZN(n18317) );
  OAI211_X1 U21387 ( .C1(n18388), .C2(n18598), .A(n18318), .B(n18317), .ZN(
        P3_U2915) );
  NOR2_X1 U21388 ( .A1(n18319), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18391) );
  NAND2_X1 U21389 ( .A1(n18622), .A2(n18391), .ZN(n18338) );
  INV_X1 U21390 ( .A(n18338), .ZN(n18406) );
  NOR2_X1 U21391 ( .A1(n18380), .A2(n18406), .ZN(n18366) );
  NOR2_X1 U21392 ( .A1(n18539), .A2(n18366), .ZN(n18339) );
  AOI22_X1 U21393 ( .A1(n18541), .A2(n18363), .B1(n18540), .B2(n18339), .ZN(
        n18324) );
  OAI21_X1 U21394 ( .B1(n18411), .B2(n18320), .A(n18366), .ZN(n18322) );
  NAND2_X1 U21395 ( .A1(n18322), .A2(n18321), .ZN(n18340) );
  AOI22_X1 U21396 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18340), .B1(
        n18406), .B2(n18546), .ZN(n18323) );
  OAI211_X1 U21397 ( .C1(n18549), .C2(n18343), .A(n18324), .B(n18323), .ZN(
        P3_U2916) );
  AOI22_X1 U21398 ( .A1(n18551), .A2(n18363), .B1(n18550), .B2(n18339), .ZN(
        n18326) );
  AOI22_X1 U21399 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18340), .B1(
        n18552), .B2(n18335), .ZN(n18325) );
  OAI211_X1 U21400 ( .C1(n18338), .C2(n18555), .A(n18326), .B(n18325), .ZN(
        P3_U2917) );
  AOI22_X1 U21401 ( .A1(n18557), .A2(n18363), .B1(n18556), .B2(n18339), .ZN(
        n18328) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18340), .B1(
        n18406), .B2(n18558), .ZN(n18327) );
  OAI211_X1 U21403 ( .C1(n18561), .C2(n18343), .A(n18328), .B(n18327), .ZN(
        P3_U2918) );
  AOI22_X1 U21404 ( .A1(n18563), .A2(n18335), .B1(n18562), .B2(n18339), .ZN(
        n18330) );
  AOI22_X1 U21405 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18340), .B1(
        n18564), .B2(n18363), .ZN(n18329) );
  OAI211_X1 U21406 ( .C1(n18338), .C2(n18567), .A(n18330), .B(n18329), .ZN(
        P3_U2919) );
  AOI22_X1 U21407 ( .A1(n18524), .A2(n18335), .B1(n18569), .B2(n18339), .ZN(
        n18332) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18340), .B1(
        n18568), .B2(n18363), .ZN(n18331) );
  OAI211_X1 U21409 ( .C1(n18338), .C2(n18527), .A(n18332), .B(n18331), .ZN(
        P3_U2920) );
  AOI22_X1 U21410 ( .A1(n18578), .A2(n18363), .B1(n18576), .B2(n18339), .ZN(
        n18334) );
  AOI22_X1 U21411 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18340), .B1(
        n18577), .B2(n18335), .ZN(n18333) );
  OAI211_X1 U21412 ( .C1(n18338), .C2(n18581), .A(n18334), .B(n18333), .ZN(
        P3_U2921) );
  AOI22_X1 U21413 ( .A1(n18584), .A2(n18335), .B1(n18582), .B2(n18339), .ZN(
        n18337) );
  AOI22_X1 U21414 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18340), .B1(
        n18583), .B2(n18363), .ZN(n18336) );
  OAI211_X1 U21415 ( .C1(n18338), .C2(n18587), .A(n18337), .B(n18336), .ZN(
        P3_U2922) );
  INV_X1 U21416 ( .A(n18591), .ZN(n18505) );
  AOI22_X1 U21417 ( .A1(n18593), .A2(n18363), .B1(n18589), .B2(n18339), .ZN(
        n18342) );
  AOI22_X1 U21418 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18340), .B1(
        n18406), .B2(n18500), .ZN(n18341) );
  OAI211_X1 U21419 ( .C1(n18505), .C2(n18343), .A(n18342), .B(n18341), .ZN(
        P3_U2923) );
  INV_X1 U21420 ( .A(n18391), .ZN(n18346) );
  NOR2_X2 U21421 ( .A1(n18622), .A2(n18346), .ZN(n18431) );
  NAND3_X1 U21422 ( .A1(n18542), .A2(n18345), .A3(n18344), .ZN(n18362) );
  NOR2_X1 U21423 ( .A1(n18539), .A2(n18346), .ZN(n18361) );
  AOI22_X1 U21424 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18362), .B1(
        n18540), .B2(n18361), .ZN(n18348) );
  AOI22_X1 U21425 ( .A1(n18506), .A2(n18363), .B1(n18380), .B2(n18541), .ZN(
        n18347) );
  OAI211_X1 U21426 ( .C1(n18425), .C2(n18515), .A(n18348), .B(n18347), .ZN(
        P3_U2924) );
  AOI22_X1 U21427 ( .A1(n18550), .A2(n18361), .B1(n18552), .B2(n18363), .ZN(
        n18350) );
  AOI22_X1 U21428 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18362), .B1(
        n18380), .B2(n18551), .ZN(n18349) );
  OAI211_X1 U21429 ( .C1(n18425), .C2(n18555), .A(n18350), .B(n18349), .ZN(
        P3_U2925) );
  AOI22_X1 U21430 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18362), .B1(
        n18556), .B2(n18361), .ZN(n18352) );
  AOI22_X1 U21431 ( .A1(n18380), .A2(n18557), .B1(n18518), .B2(n18363), .ZN(
        n18351) );
  OAI211_X1 U21432 ( .C1(n18425), .C2(n18521), .A(n18352), .B(n18351), .ZN(
        P3_U2926) );
  AOI22_X1 U21433 ( .A1(n18563), .A2(n18363), .B1(n18562), .B2(n18361), .ZN(
        n18354) );
  AOI22_X1 U21434 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18362), .B1(
        n18380), .B2(n18564), .ZN(n18353) );
  OAI211_X1 U21435 ( .C1(n18425), .C2(n18567), .A(n18354), .B(n18353), .ZN(
        P3_U2927) );
  AOI22_X1 U21436 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18362), .B1(
        n18569), .B2(n18361), .ZN(n18356) );
  AOI22_X1 U21437 ( .A1(n18380), .A2(n18568), .B1(n18524), .B2(n18363), .ZN(
        n18355) );
  OAI211_X1 U21438 ( .C1(n18425), .C2(n18527), .A(n18356), .B(n18355), .ZN(
        P3_U2928) );
  AOI22_X1 U21439 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18362), .B1(
        n18576), .B2(n18361), .ZN(n18358) );
  AOI22_X1 U21440 ( .A1(n18380), .A2(n18578), .B1(n18577), .B2(n18363), .ZN(
        n18357) );
  OAI211_X1 U21441 ( .C1(n18425), .C2(n18581), .A(n18358), .B(n18357), .ZN(
        P3_U2929) );
  AOI22_X1 U21442 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18362), .B1(
        n18582), .B2(n18361), .ZN(n18360) );
  AOI22_X1 U21443 ( .A1(n18380), .A2(n18583), .B1(n18584), .B2(n18363), .ZN(
        n18359) );
  OAI211_X1 U21444 ( .C1(n18425), .C2(n18587), .A(n18360), .B(n18359), .ZN(
        P3_U2930) );
  AOI22_X1 U21445 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18362), .B1(
        n18589), .B2(n18361), .ZN(n18365) );
  AOI22_X1 U21446 ( .A1(n18380), .A2(n18593), .B1(n18591), .B2(n18363), .ZN(
        n18364) );
  OAI211_X1 U21447 ( .C1(n18425), .C2(n18598), .A(n18365), .B(n18364), .ZN(
        P3_U2931) );
  NAND2_X1 U21448 ( .A1(n18627), .A2(n18390), .ZN(n18383) );
  AOI21_X1 U21449 ( .B1(n18383), .B2(n18425), .A(n18539), .ZN(n18384) );
  AOI22_X1 U21450 ( .A1(n18406), .A2(n18541), .B1(n18540), .B2(n18384), .ZN(
        n18369) );
  AOI221_X1 U21451 ( .B1(n18366), .B2(n18425), .C1(n18411), .C2(n18425), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18367) );
  OAI21_X1 U21452 ( .B1(n18452), .B2(n18367), .A(n18414), .ZN(n18385) );
  AOI22_X1 U21453 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18385), .B1(
        n18452), .B2(n18546), .ZN(n18368) );
  OAI211_X1 U21454 ( .C1(n18549), .C2(n18388), .A(n18369), .B(n18368), .ZN(
        P3_U2932) );
  AOI22_X1 U21455 ( .A1(n18380), .A2(n18552), .B1(n18384), .B2(n18550), .ZN(
        n18371) );
  AOI22_X1 U21456 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18385), .B1(
        n18406), .B2(n18551), .ZN(n18370) );
  OAI211_X1 U21457 ( .C1(n18383), .C2(n18555), .A(n18371), .B(n18370), .ZN(
        P3_U2933) );
  AOI22_X1 U21458 ( .A1(n18406), .A2(n18557), .B1(n18384), .B2(n18556), .ZN(
        n18373) );
  AOI22_X1 U21459 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18385), .B1(
        n18452), .B2(n18558), .ZN(n18372) );
  OAI211_X1 U21460 ( .C1(n18388), .C2(n18561), .A(n18373), .B(n18372), .ZN(
        P3_U2934) );
  AOI22_X1 U21461 ( .A1(n18380), .A2(n18563), .B1(n18384), .B2(n18562), .ZN(
        n18375) );
  AOI22_X1 U21462 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18385), .B1(
        n18406), .B2(n18564), .ZN(n18374) );
  OAI211_X1 U21463 ( .C1(n18383), .C2(n18567), .A(n18375), .B(n18374), .ZN(
        P3_U2935) );
  INV_X1 U21464 ( .A(n18524), .ZN(n18575) );
  AOI22_X1 U21465 ( .A1(n18406), .A2(n18568), .B1(n18384), .B2(n18569), .ZN(
        n18377) );
  AOI22_X1 U21466 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18385), .B1(
        n18452), .B2(n18571), .ZN(n18376) );
  OAI211_X1 U21467 ( .C1(n18388), .C2(n18575), .A(n18377), .B(n18376), .ZN(
        P3_U2936) );
  AOI22_X1 U21468 ( .A1(n18380), .A2(n18577), .B1(n18384), .B2(n18576), .ZN(
        n18379) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18385), .B1(
        n18406), .B2(n18578), .ZN(n18378) );
  OAI211_X1 U21470 ( .C1(n18383), .C2(n18581), .A(n18379), .B(n18378), .ZN(
        P3_U2937) );
  AOI22_X1 U21471 ( .A1(n18380), .A2(n18584), .B1(n18384), .B2(n18582), .ZN(
        n18382) );
  AOI22_X1 U21472 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18385), .B1(
        n18406), .B2(n18583), .ZN(n18381) );
  OAI211_X1 U21473 ( .C1(n18383), .C2(n18587), .A(n18382), .B(n18381), .ZN(
        P3_U2938) );
  AOI22_X1 U21474 ( .A1(n18406), .A2(n18593), .B1(n18384), .B2(n18589), .ZN(
        n18387) );
  AOI22_X1 U21475 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18385), .B1(
        n18452), .B2(n18500), .ZN(n18386) );
  OAI211_X1 U21476 ( .C1(n18388), .C2(n18505), .A(n18387), .B(n18386), .ZN(
        P3_U2939) );
  NOR2_X2 U21477 ( .A1(n18389), .A2(n18410), .ZN(n18475) );
  NOR2_X1 U21478 ( .A1(n18410), .A2(n18479), .ZN(n18436) );
  AOI22_X1 U21479 ( .A1(n18431), .A2(n18541), .B1(n18540), .B2(n18436), .ZN(
        n18393) );
  AOI22_X1 U21480 ( .A1(n18545), .A2(n18391), .B1(n18390), .B2(n18481), .ZN(
        n18407) );
  AOI22_X1 U21481 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18407), .B1(
        n18506), .B2(n18406), .ZN(n18392) );
  OAI211_X1 U21482 ( .C1(n18515), .C2(n18469), .A(n18393), .B(n18392), .ZN(
        P3_U2940) );
  AOI22_X1 U21483 ( .A1(n18406), .A2(n18552), .B1(n18550), .B2(n18436), .ZN(
        n18395) );
  AOI22_X1 U21484 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18407), .B1(
        n18431), .B2(n18551), .ZN(n18394) );
  OAI211_X1 U21485 ( .C1(n18555), .C2(n18469), .A(n18395), .B(n18394), .ZN(
        P3_U2941) );
  AOI22_X1 U21486 ( .A1(n18406), .A2(n18518), .B1(n18556), .B2(n18436), .ZN(
        n18397) );
  AOI22_X1 U21487 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18407), .B1(
        n18431), .B2(n18557), .ZN(n18396) );
  OAI211_X1 U21488 ( .C1(n18521), .C2(n18469), .A(n18397), .B(n18396), .ZN(
        P3_U2942) );
  AOI22_X1 U21489 ( .A1(n18406), .A2(n18563), .B1(n18562), .B2(n18436), .ZN(
        n18399) );
  AOI22_X1 U21490 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18407), .B1(
        n18431), .B2(n18564), .ZN(n18398) );
  OAI211_X1 U21491 ( .C1(n18567), .C2(n18469), .A(n18399), .B(n18398), .ZN(
        P3_U2943) );
  AOI22_X1 U21492 ( .A1(n18406), .A2(n18524), .B1(n18569), .B2(n18436), .ZN(
        n18401) );
  AOI22_X1 U21493 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18407), .B1(
        n18431), .B2(n18568), .ZN(n18400) );
  OAI211_X1 U21494 ( .C1(n18527), .C2(n18469), .A(n18401), .B(n18400), .ZN(
        P3_U2944) );
  AOI22_X1 U21495 ( .A1(n18431), .A2(n18578), .B1(n18576), .B2(n18436), .ZN(
        n18403) );
  AOI22_X1 U21496 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18407), .B1(
        n18406), .B2(n18577), .ZN(n18402) );
  OAI211_X1 U21497 ( .C1(n18581), .C2(n18469), .A(n18403), .B(n18402), .ZN(
        P3_U2945) );
  AOI22_X1 U21498 ( .A1(n18406), .A2(n18584), .B1(n18582), .B2(n18436), .ZN(
        n18405) );
  AOI22_X1 U21499 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18407), .B1(
        n18431), .B2(n18583), .ZN(n18404) );
  OAI211_X1 U21500 ( .C1(n18587), .C2(n18469), .A(n18405), .B(n18404), .ZN(
        P3_U2946) );
  AOI22_X1 U21501 ( .A1(n18431), .A2(n18593), .B1(n18589), .B2(n18436), .ZN(
        n18409) );
  AOI22_X1 U21502 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18407), .B1(
        n18406), .B2(n18591), .ZN(n18408) );
  OAI211_X1 U21503 ( .C1(n18598), .C2(n18469), .A(n18409), .B(n18408), .ZN(
        P3_U2947) );
  NAND2_X1 U21504 ( .A1(n18483), .A2(n18622), .ZN(n18504) );
  INV_X1 U21505 ( .A(n18504), .ZN(n18496) );
  NOR2_X1 U21506 ( .A1(n18475), .A2(n18496), .ZN(n18457) );
  NOR2_X1 U21507 ( .A1(n18539), .A2(n18457), .ZN(n18430) );
  AOI22_X1 U21508 ( .A1(n18506), .A2(n18431), .B1(n18540), .B2(n18430), .ZN(
        n18416) );
  NOR2_X1 U21509 ( .A1(n18452), .A2(n18431), .ZN(n18412) );
  OAI21_X1 U21510 ( .B1(n18412), .B2(n18411), .A(n18457), .ZN(n18413) );
  OAI211_X1 U21511 ( .C1(n18496), .C2(n18752), .A(n18414), .B(n18413), .ZN(
        n18432) );
  AOI22_X1 U21512 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18432), .B1(
        n18452), .B2(n18541), .ZN(n18415) );
  OAI211_X1 U21513 ( .C1(n18515), .C2(n18504), .A(n18416), .B(n18415), .ZN(
        P3_U2948) );
  AOI22_X1 U21514 ( .A1(n18452), .A2(n18551), .B1(n18550), .B2(n18430), .ZN(
        n18418) );
  AOI22_X1 U21515 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18432), .B1(
        n18431), .B2(n18552), .ZN(n18417) );
  OAI211_X1 U21516 ( .C1(n18555), .C2(n18504), .A(n18418), .B(n18417), .ZN(
        P3_U2949) );
  AOI22_X1 U21517 ( .A1(n18452), .A2(n18557), .B1(n18556), .B2(n18430), .ZN(
        n18420) );
  AOI22_X1 U21518 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18432), .B1(
        n18558), .B2(n18496), .ZN(n18419) );
  OAI211_X1 U21519 ( .C1(n18425), .C2(n18561), .A(n18420), .B(n18419), .ZN(
        P3_U2950) );
  AOI22_X1 U21520 ( .A1(n18431), .A2(n18563), .B1(n18562), .B2(n18430), .ZN(
        n18422) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18432), .B1(
        n18452), .B2(n18564), .ZN(n18421) );
  OAI211_X1 U21522 ( .C1(n18567), .C2(n18504), .A(n18422), .B(n18421), .ZN(
        P3_U2951) );
  AOI22_X1 U21523 ( .A1(n18452), .A2(n18568), .B1(n18569), .B2(n18430), .ZN(
        n18424) );
  AOI22_X1 U21524 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18432), .B1(
        n18571), .B2(n18496), .ZN(n18423) );
  OAI211_X1 U21525 ( .C1(n18425), .C2(n18575), .A(n18424), .B(n18423), .ZN(
        P3_U2952) );
  AOI22_X1 U21526 ( .A1(n18431), .A2(n18577), .B1(n18576), .B2(n18430), .ZN(
        n18427) );
  AOI22_X1 U21527 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18432), .B1(
        n18452), .B2(n18578), .ZN(n18426) );
  OAI211_X1 U21528 ( .C1(n18581), .C2(n18504), .A(n18427), .B(n18426), .ZN(
        P3_U2953) );
  AOI22_X1 U21529 ( .A1(n18431), .A2(n18584), .B1(n18582), .B2(n18430), .ZN(
        n18429) );
  AOI22_X1 U21530 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18432), .B1(
        n18452), .B2(n18583), .ZN(n18428) );
  OAI211_X1 U21531 ( .C1(n18587), .C2(n18504), .A(n18429), .B(n18428), .ZN(
        P3_U2954) );
  AOI22_X1 U21532 ( .A1(n18431), .A2(n18591), .B1(n18589), .B2(n18430), .ZN(
        n18434) );
  AOI22_X1 U21533 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18432), .B1(
        n18452), .B2(n18593), .ZN(n18433) );
  OAI211_X1 U21534 ( .C1(n18598), .C2(n18504), .A(n18434), .B(n18433), .ZN(
        P3_U2955) );
  NAND2_X1 U21535 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18483), .ZN(
        n18456) );
  AND2_X1 U21536 ( .A1(n18435), .A2(n18483), .ZN(n18451) );
  AOI22_X1 U21537 ( .A1(n18506), .A2(n18452), .B1(n18540), .B2(n18451), .ZN(
        n18438) );
  AOI22_X1 U21538 ( .A1(n18545), .A2(n18436), .B1(n18542), .B2(n18483), .ZN(
        n18453) );
  AOI22_X1 U21539 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18453), .B1(
        n18541), .B2(n18475), .ZN(n18437) );
  OAI211_X1 U21540 ( .C1(n18515), .C2(n18456), .A(n18438), .B(n18437), .ZN(
        P3_U2956) );
  AOI22_X1 U21541 ( .A1(n18551), .A2(n18475), .B1(n18550), .B2(n18451), .ZN(
        n18440) );
  AOI22_X1 U21542 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18453), .B1(
        n18452), .B2(n18552), .ZN(n18439) );
  OAI211_X1 U21543 ( .C1(n18555), .C2(n18456), .A(n18440), .B(n18439), .ZN(
        P3_U2957) );
  AOI22_X1 U21544 ( .A1(n18452), .A2(n18518), .B1(n18556), .B2(n18451), .ZN(
        n18442) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18453), .B1(
        n18557), .B2(n18475), .ZN(n18441) );
  OAI211_X1 U21546 ( .C1(n18521), .C2(n18456), .A(n18442), .B(n18441), .ZN(
        P3_U2958) );
  AOI22_X1 U21547 ( .A1(n18564), .A2(n18475), .B1(n18562), .B2(n18451), .ZN(
        n18444) );
  AOI22_X1 U21548 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18453), .B1(
        n18452), .B2(n18563), .ZN(n18443) );
  OAI211_X1 U21549 ( .C1(n18567), .C2(n18456), .A(n18444), .B(n18443), .ZN(
        P3_U2959) );
  AOI22_X1 U21550 ( .A1(n18569), .A2(n18451), .B1(n18568), .B2(n18475), .ZN(
        n18446) );
  AOI22_X1 U21551 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18453), .B1(
        n18452), .B2(n18524), .ZN(n18445) );
  OAI211_X1 U21552 ( .C1(n18527), .C2(n18456), .A(n18446), .B(n18445), .ZN(
        P3_U2960) );
  AOI22_X1 U21553 ( .A1(n18578), .A2(n18475), .B1(n18576), .B2(n18451), .ZN(
        n18448) );
  AOI22_X1 U21554 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18453), .B1(
        n18452), .B2(n18577), .ZN(n18447) );
  OAI211_X1 U21555 ( .C1(n18581), .C2(n18456), .A(n18448), .B(n18447), .ZN(
        P3_U2961) );
  AOI22_X1 U21556 ( .A1(n18452), .A2(n18584), .B1(n18582), .B2(n18451), .ZN(
        n18450) );
  AOI22_X1 U21557 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18453), .B1(
        n18583), .B2(n18475), .ZN(n18449) );
  OAI211_X1 U21558 ( .C1(n18587), .C2(n18456), .A(n18450), .B(n18449), .ZN(
        P3_U2962) );
  AOI22_X1 U21559 ( .A1(n18452), .A2(n18591), .B1(n18589), .B2(n18451), .ZN(
        n18455) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18453), .B1(
        n18593), .B2(n18475), .ZN(n18454) );
  OAI211_X1 U21561 ( .C1(n18598), .C2(n18456), .A(n18455), .B(n18454), .ZN(
        P3_U2963) );
  NAND2_X1 U21562 ( .A1(n18627), .A2(n18482), .ZN(n18574) );
  INV_X1 U21563 ( .A(n18574), .ZN(n18590) );
  NOR2_X1 U21564 ( .A1(n18533), .A2(n18590), .ZN(n18508) );
  NOR2_X1 U21565 ( .A1(n18539), .A2(n18508), .ZN(n18474) );
  AOI22_X1 U21566 ( .A1(n18506), .A2(n18475), .B1(n18540), .B2(n18474), .ZN(
        n18460) );
  OAI22_X1 U21567 ( .A1(n18457), .A2(n18507), .B1(n18508), .B2(n18509), .ZN(
        n18458) );
  OAI21_X1 U21568 ( .B1(n18590), .B2(n18752), .A(n18458), .ZN(n18476) );
  AOI22_X1 U21569 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18476), .B1(
        n18541), .B2(n18496), .ZN(n18459) );
  OAI211_X1 U21570 ( .C1(n18515), .C2(n18574), .A(n18460), .B(n18459), .ZN(
        P3_U2964) );
  AOI22_X1 U21571 ( .A1(n18550), .A2(n18474), .B1(n18552), .B2(n18475), .ZN(
        n18462) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18476), .B1(
        n18551), .B2(n18496), .ZN(n18461) );
  OAI211_X1 U21573 ( .C1(n18555), .C2(n18574), .A(n18462), .B(n18461), .ZN(
        P3_U2965) );
  AOI22_X1 U21574 ( .A1(n18518), .A2(n18475), .B1(n18556), .B2(n18474), .ZN(
        n18464) );
  AOI22_X1 U21575 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18476), .B1(
        n18557), .B2(n18496), .ZN(n18463) );
  OAI211_X1 U21576 ( .C1(n18521), .C2(n18574), .A(n18464), .B(n18463), .ZN(
        P3_U2966) );
  AOI22_X1 U21577 ( .A1(n18564), .A2(n18496), .B1(n18562), .B2(n18474), .ZN(
        n18466) );
  AOI22_X1 U21578 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18476), .B1(
        n18563), .B2(n18475), .ZN(n18465) );
  OAI211_X1 U21579 ( .C1(n18567), .C2(n18574), .A(n18466), .B(n18465), .ZN(
        P3_U2967) );
  AOI22_X1 U21580 ( .A1(n18569), .A2(n18474), .B1(n18568), .B2(n18496), .ZN(
        n18468) );
  AOI22_X1 U21581 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18476), .B1(
        n18571), .B2(n18590), .ZN(n18467) );
  OAI211_X1 U21582 ( .C1(n18575), .C2(n18469), .A(n18468), .B(n18467), .ZN(
        P3_U2968) );
  AOI22_X1 U21583 ( .A1(n18578), .A2(n18496), .B1(n18576), .B2(n18474), .ZN(
        n18471) );
  AOI22_X1 U21584 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18476), .B1(
        n18577), .B2(n18475), .ZN(n18470) );
  OAI211_X1 U21585 ( .C1(n18581), .C2(n18574), .A(n18471), .B(n18470), .ZN(
        P3_U2969) );
  AOI22_X1 U21586 ( .A1(n18584), .A2(n18475), .B1(n18582), .B2(n18474), .ZN(
        n18473) );
  AOI22_X1 U21587 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18476), .B1(
        n18583), .B2(n18496), .ZN(n18472) );
  OAI211_X1 U21588 ( .C1(n18587), .C2(n18574), .A(n18473), .B(n18472), .ZN(
        P3_U2970) );
  AOI22_X1 U21589 ( .A1(n18591), .A2(n18475), .B1(n18589), .B2(n18474), .ZN(
        n18478) );
  AOI22_X1 U21590 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18476), .B1(
        n18593), .B2(n18496), .ZN(n18477) );
  OAI211_X1 U21591 ( .C1(n18598), .C2(n18574), .A(n18478), .B(n18477), .ZN(
        P3_U2971) );
  INV_X1 U21592 ( .A(n18482), .ZN(n18480) );
  NOR2_X1 U21593 ( .A1(n18480), .A2(n18479), .ZN(n18544) );
  AOI22_X1 U21594 ( .A1(n18506), .A2(n18496), .B1(n18540), .B2(n18544), .ZN(
        n18485) );
  AOI22_X1 U21595 ( .A1(n18545), .A2(n18483), .B1(n18482), .B2(n18481), .ZN(
        n18501) );
  AOI22_X1 U21596 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18501), .B1(
        n18541), .B2(n18533), .ZN(n18484) );
  OAI211_X1 U21597 ( .C1(n18515), .C2(n18499), .A(n18485), .B(n18484), .ZN(
        P3_U2972) );
  AOI22_X1 U21598 ( .A1(n18551), .A2(n18533), .B1(n18550), .B2(n18544), .ZN(
        n18487) );
  AOI22_X1 U21599 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18501), .B1(
        n18552), .B2(n18496), .ZN(n18486) );
  OAI211_X1 U21600 ( .C1(n18555), .C2(n18499), .A(n18487), .B(n18486), .ZN(
        P3_U2973) );
  AOI22_X1 U21601 ( .A1(n18557), .A2(n18533), .B1(n18556), .B2(n18544), .ZN(
        n18489) );
  AOI22_X1 U21602 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18501), .B1(
        n18558), .B2(n18592), .ZN(n18488) );
  OAI211_X1 U21603 ( .C1(n18561), .C2(n18504), .A(n18489), .B(n18488), .ZN(
        P3_U2974) );
  AOI22_X1 U21604 ( .A1(n18563), .A2(n18496), .B1(n18562), .B2(n18544), .ZN(
        n18491) );
  AOI22_X1 U21605 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18501), .B1(
        n18564), .B2(n18533), .ZN(n18490) );
  OAI211_X1 U21606 ( .C1(n18567), .C2(n18499), .A(n18491), .B(n18490), .ZN(
        P3_U2975) );
  AOI22_X1 U21607 ( .A1(n18524), .A2(n18496), .B1(n18569), .B2(n18544), .ZN(
        n18493) );
  AOI22_X1 U21608 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18501), .B1(
        n18568), .B2(n18533), .ZN(n18492) );
  OAI211_X1 U21609 ( .C1(n18527), .C2(n18499), .A(n18493), .B(n18492), .ZN(
        P3_U2976) );
  AOI22_X1 U21610 ( .A1(n18577), .A2(n18496), .B1(n18576), .B2(n18544), .ZN(
        n18495) );
  AOI22_X1 U21611 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18501), .B1(
        n18578), .B2(n18533), .ZN(n18494) );
  OAI211_X1 U21612 ( .C1(n18581), .C2(n18499), .A(n18495), .B(n18494), .ZN(
        P3_U2977) );
  AOI22_X1 U21613 ( .A1(n18584), .A2(n18496), .B1(n18582), .B2(n18544), .ZN(
        n18498) );
  AOI22_X1 U21614 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18501), .B1(
        n18583), .B2(n18533), .ZN(n18497) );
  OAI211_X1 U21615 ( .C1(n18587), .C2(n18499), .A(n18498), .B(n18497), .ZN(
        P3_U2978) );
  AOI22_X1 U21616 ( .A1(n18593), .A2(n18533), .B1(n18589), .B2(n18544), .ZN(
        n18503) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18501), .B1(
        n18500), .B2(n18592), .ZN(n18502) );
  OAI211_X1 U21618 ( .C1(n18505), .C2(n18504), .A(n18503), .B(n18502), .ZN(
        P3_U2979) );
  NOR2_X1 U21619 ( .A1(n18539), .A2(n18510), .ZN(n18532) );
  AOI22_X1 U21620 ( .A1(n18506), .A2(n18533), .B1(n18540), .B2(n18532), .ZN(
        n18514) );
  OAI22_X1 U21621 ( .A1(n18510), .A2(n18509), .B1(n18508), .B2(n18507), .ZN(
        n18511) );
  OAI21_X1 U21622 ( .B1(n18512), .B2(n18752), .A(n18511), .ZN(n18534) );
  AOI22_X1 U21623 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18534), .B1(
        n18541), .B2(n18590), .ZN(n18513) );
  OAI211_X1 U21624 ( .C1(n18515), .C2(n18537), .A(n18514), .B(n18513), .ZN(
        P3_U2980) );
  AOI22_X1 U21625 ( .A1(n18551), .A2(n18590), .B1(n18550), .B2(n18532), .ZN(
        n18517) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18534), .B1(
        n18552), .B2(n18533), .ZN(n18516) );
  OAI211_X1 U21627 ( .C1(n18555), .C2(n18537), .A(n18517), .B(n18516), .ZN(
        P3_U2981) );
  AOI22_X1 U21628 ( .A1(n18518), .A2(n18533), .B1(n18556), .B2(n18532), .ZN(
        n18520) );
  AOI22_X1 U21629 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18534), .B1(
        n18557), .B2(n18590), .ZN(n18519) );
  OAI211_X1 U21630 ( .C1(n18521), .C2(n18537), .A(n18520), .B(n18519), .ZN(
        P3_U2982) );
  AOI22_X1 U21631 ( .A1(n18563), .A2(n18533), .B1(n18562), .B2(n18532), .ZN(
        n18523) );
  AOI22_X1 U21632 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18534), .B1(
        n18564), .B2(n18590), .ZN(n18522) );
  OAI211_X1 U21633 ( .C1(n18567), .C2(n18537), .A(n18523), .B(n18522), .ZN(
        P3_U2983) );
  AOI22_X1 U21634 ( .A1(n18524), .A2(n18533), .B1(n18569), .B2(n18532), .ZN(
        n18526) );
  AOI22_X1 U21635 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18534), .B1(
        n18568), .B2(n18590), .ZN(n18525) );
  OAI211_X1 U21636 ( .C1(n18527), .C2(n18537), .A(n18526), .B(n18525), .ZN(
        P3_U2984) );
  AOI22_X1 U21637 ( .A1(n18577), .A2(n18533), .B1(n18576), .B2(n18532), .ZN(
        n18529) );
  AOI22_X1 U21638 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18534), .B1(
        n18578), .B2(n18590), .ZN(n18528) );
  OAI211_X1 U21639 ( .C1(n18581), .C2(n18537), .A(n18529), .B(n18528), .ZN(
        P3_U2985) );
  AOI22_X1 U21640 ( .A1(n18584), .A2(n18533), .B1(n18582), .B2(n18532), .ZN(
        n18531) );
  AOI22_X1 U21641 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18534), .B1(
        n18583), .B2(n18590), .ZN(n18530) );
  OAI211_X1 U21642 ( .C1(n18587), .C2(n18537), .A(n18531), .B(n18530), .ZN(
        P3_U2986) );
  AOI22_X1 U21643 ( .A1(n18591), .A2(n18533), .B1(n18589), .B2(n18532), .ZN(
        n18536) );
  AOI22_X1 U21644 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18534), .B1(
        n18593), .B2(n18590), .ZN(n18535) );
  OAI211_X1 U21645 ( .C1(n18598), .C2(n18537), .A(n18536), .B(n18535), .ZN(
        P3_U2987) );
  INV_X1 U21646 ( .A(n18543), .ZN(n18538) );
  NOR2_X1 U21647 ( .A1(n18539), .A2(n18538), .ZN(n18588) );
  AOI22_X1 U21648 ( .A1(n18541), .A2(n18592), .B1(n18540), .B2(n18588), .ZN(
        n18548) );
  AOI22_X1 U21649 ( .A1(n18545), .A2(n18544), .B1(n18543), .B2(n18542), .ZN(
        n18594) );
  AOI22_X1 U21650 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18594), .B1(
        n18546), .B2(n18570), .ZN(n18547) );
  OAI211_X1 U21651 ( .C1(n18549), .C2(n18574), .A(n18548), .B(n18547), .ZN(
        P3_U2988) );
  AOI22_X1 U21652 ( .A1(n18551), .A2(n18592), .B1(n18550), .B2(n18588), .ZN(
        n18554) );
  AOI22_X1 U21653 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18594), .B1(
        n18552), .B2(n18590), .ZN(n18553) );
  OAI211_X1 U21654 ( .C1(n18555), .C2(n18597), .A(n18554), .B(n18553), .ZN(
        P3_U2989) );
  AOI22_X1 U21655 ( .A1(n18557), .A2(n18592), .B1(n18556), .B2(n18588), .ZN(
        n18560) );
  AOI22_X1 U21656 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18594), .B1(
        n18558), .B2(n18570), .ZN(n18559) );
  OAI211_X1 U21657 ( .C1(n18561), .C2(n18574), .A(n18560), .B(n18559), .ZN(
        P3_U2990) );
  AOI22_X1 U21658 ( .A1(n18563), .A2(n18590), .B1(n18562), .B2(n18588), .ZN(
        n18566) );
  AOI22_X1 U21659 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18594), .B1(
        n18564), .B2(n18592), .ZN(n18565) );
  OAI211_X1 U21660 ( .C1(n18567), .C2(n18597), .A(n18566), .B(n18565), .ZN(
        P3_U2991) );
  AOI22_X1 U21661 ( .A1(n18569), .A2(n18588), .B1(n18568), .B2(n18592), .ZN(
        n18573) );
  AOI22_X1 U21662 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18594), .B1(
        n18571), .B2(n18570), .ZN(n18572) );
  OAI211_X1 U21663 ( .C1(n18575), .C2(n18574), .A(n18573), .B(n18572), .ZN(
        P3_U2992) );
  AOI22_X1 U21664 ( .A1(n18577), .A2(n18590), .B1(n18576), .B2(n18588), .ZN(
        n18580) );
  AOI22_X1 U21665 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18594), .B1(
        n18578), .B2(n18592), .ZN(n18579) );
  OAI211_X1 U21666 ( .C1(n18581), .C2(n18597), .A(n18580), .B(n18579), .ZN(
        P3_U2993) );
  AOI22_X1 U21667 ( .A1(n18583), .A2(n18592), .B1(n18582), .B2(n18588), .ZN(
        n18586) );
  AOI22_X1 U21668 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18594), .B1(
        n18584), .B2(n18590), .ZN(n18585) );
  OAI211_X1 U21669 ( .C1(n18587), .C2(n18597), .A(n18586), .B(n18585), .ZN(
        P3_U2994) );
  AOI22_X1 U21670 ( .A1(n18591), .A2(n18590), .B1(n18589), .B2(n18588), .ZN(
        n18596) );
  AOI22_X1 U21671 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18594), .B1(
        n18593), .B2(n18592), .ZN(n18595) );
  OAI211_X1 U21672 ( .C1(n18598), .C2(n18597), .A(n18596), .B(n18595), .ZN(
        P3_U2995) );
  AOI211_X1 U21673 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18626), .A(
        n18600), .B(n18599), .ZN(n18650) );
  OAI22_X1 U21674 ( .A1(n18602), .A2(n18601), .B1(n18795), .B2(n18613), .ZN(
        n18798) );
  AOI221_X1 U21675 ( .B1(P3_MORE_REG_SCAN_IN), .B2(n18603), .C1(
        P3_FLUSH_REG_SCAN_IN), .C2(n18603), .A(n18798), .ZN(n18649) );
  AOI21_X1 U21676 ( .B1(n18606), .B2(n18605), .A(n18604), .ZN(n18629) );
  OAI21_X1 U21677 ( .B1(n18607), .B2(n18631), .A(n18612), .ZN(n18609) );
  OAI211_X1 U21678 ( .C1(n18610), .C2(n18629), .A(n18609), .B(n18608), .ZN(
        n18758) );
  NOR2_X1 U21679 ( .A1(n18626), .A2(n18758), .ZN(n18616) );
  AOI211_X1 U21680 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18611), .A(
        n18632), .B(n18631), .ZN(n18634) );
  OAI22_X1 U21681 ( .A1(n18614), .A2(n18613), .B1(n18634), .B2(n18612), .ZN(
        n18755) );
  NAND2_X1 U21682 ( .A1(n20789), .A2(n18755), .ZN(n18615) );
  OAI22_X1 U21683 ( .A1(n18616), .A2(n20789), .B1(n18626), .B2(n18615), .ZN(
        n18647) );
  NAND2_X1 U21684 ( .A1(n18618), .A2(n18617), .ZN(n18620) );
  INV_X1 U21685 ( .A(n18634), .ZN(n18619) );
  AOI22_X1 U21686 ( .A1(n18775), .A2(n18620), .B1(n18778), .B2(n18619), .ZN(
        n18772) );
  AOI22_X1 U21687 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18621), .B1(
        n18620), .B2(n18784), .ZN(n18624) );
  INV_X1 U21688 ( .A(n18624), .ZN(n18780) );
  NOR3_X1 U21689 ( .A1(n18623), .A2(n18622), .A3(n18780), .ZN(n18625) );
  OAI22_X1 U21690 ( .A1(n18772), .A2(n18625), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18624), .ZN(n18628) );
  INV_X1 U21691 ( .A(n18626), .ZN(n18640) );
  AOI21_X1 U21692 ( .B1(n18628), .B2(n18640), .A(n18627), .ZN(n18642) );
  NOR3_X1 U21693 ( .A1(n18630), .A2(n18629), .A3(n18771), .ZN(n18638) );
  NOR2_X1 U21694 ( .A1(n18632), .A2(n18631), .ZN(n18636) );
  OAI22_X1 U21695 ( .A1(n18636), .A2(n18635), .B1(n18634), .B2(n18633), .ZN(
        n18637) );
  AOI211_X1 U21696 ( .C1(n18639), .C2(n18764), .A(n18638), .B(n18637), .ZN(
        n18767) );
  MUX2_X1 U21697 ( .A(n18771), .B(n18767), .S(n18640), .Z(n18643) );
  OR2_X1 U21698 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18643), .ZN(
        n18641) );
  AOI221_X1 U21699 ( .B1(n18642), .B2(n18641), .C1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C2(n18643), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18646) );
  OAI21_X1 U21700 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n18643), .ZN(n18645) );
  AOI222_X1 U21701 ( .A1(n18647), .A2(n18646), .B1(n18647), .B2(n18645), .C1(
        n18646), .C2(n18644), .ZN(n18648) );
  NAND4_X1 U21702 ( .A1(n18650), .A2(n18649), .A3(n18648), .A4(n18794), .ZN(
        n18651) );
  INV_X1 U21703 ( .A(n18651), .ZN(n18659) );
  AOI22_X1 U21704 ( .A1(n18779), .A2(n18667), .B1(n18805), .B2(n17394), .ZN(
        n18656) );
  AOI211_X1 U21705 ( .C1(n18653), .C2(n18652), .A(n18658), .B(n18651), .ZN(
        n18654) );
  NOR2_X1 U21706 ( .A1(n18654), .A2(n18808), .ZN(n18753) );
  NAND2_X1 U21707 ( .A1(n18805), .A2(n18820), .ZN(n18660) );
  OAI211_X1 U21708 ( .C1(n18807), .C2(n18752), .A(n18753), .B(n18660), .ZN(
        n18663) );
  OAI22_X1 U21709 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18656), .B1(n18655), 
        .B2(n18663), .ZN(n18657) );
  OAI21_X1 U21710 ( .B1(n18659), .B2(n18658), .A(n18657), .ZN(P3_U2996) );
  NOR3_X1 U21711 ( .A1(n18763), .A2(n18808), .A3(n18660), .ZN(n18665) );
  AOI211_X1 U21712 ( .C1(n18805), .C2(n17394), .A(n18661), .B(n18665), .ZN(
        n18662) );
  OAI21_X1 U21713 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n18663), .A(n18662), 
        .ZN(P3_U2997) );
  NOR4_X1 U21714 ( .A1(n18667), .A2(n18666), .A3(n18665), .A4(n18664), .ZN(
        P3_U2998) );
  INV_X1 U21715 ( .A(P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20704) );
  NOR2_X1 U21716 ( .A1(n20704), .A2(n18750), .ZN(P3_U2999) );
  AND2_X1 U21717 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18668), .ZN(
        P3_U3000) );
  AND2_X1 U21718 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18668), .ZN(
        P3_U3001) );
  AND2_X1 U21719 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18668), .ZN(
        P3_U3002) );
  AND2_X1 U21720 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18668), .ZN(
        P3_U3003) );
  AND2_X1 U21721 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18668), .ZN(
        P3_U3004) );
  AND2_X1 U21722 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18668), .ZN(
        P3_U3005) );
  AND2_X1 U21723 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18668), .ZN(
        P3_U3006) );
  AND2_X1 U21724 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18668), .ZN(
        P3_U3007) );
  AND2_X1 U21725 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18668), .ZN(
        P3_U3008) );
  AND2_X1 U21726 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18668), .ZN(
        P3_U3009) );
  AND2_X1 U21727 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18668), .ZN(
        P3_U3010) );
  AND2_X1 U21728 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18668), .ZN(
        P3_U3011) );
  AND2_X1 U21729 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18668), .ZN(
        P3_U3012) );
  AND2_X1 U21730 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18668), .ZN(
        P3_U3013) );
  AND2_X1 U21731 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18668), .ZN(
        P3_U3014) );
  AND2_X1 U21732 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18668), .ZN(
        P3_U3015) );
  AND2_X1 U21733 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18668), .ZN(
        P3_U3016) );
  AND2_X1 U21734 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18668), .ZN(
        P3_U3017) );
  AND2_X1 U21735 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18668), .ZN(
        P3_U3018) );
  AND2_X1 U21736 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18668), .ZN(
        P3_U3019) );
  AND2_X1 U21737 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18668), .ZN(
        P3_U3020) );
  AND2_X1 U21738 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18668), .ZN(P3_U3021) );
  AND2_X1 U21739 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18668), .ZN(P3_U3022) );
  AND2_X1 U21740 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18668), .ZN(P3_U3023) );
  AND2_X1 U21741 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18668), .ZN(P3_U3024) );
  AND2_X1 U21742 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18668), .ZN(P3_U3025) );
  AND2_X1 U21743 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18668), .ZN(P3_U3026) );
  AND2_X1 U21744 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18668), .ZN(P3_U3027) );
  AND2_X1 U21745 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18668), .ZN(P3_U3028) );
  OAI21_X1 U21746 ( .B1(n18669), .B2(n20561), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18670) );
  AOI22_X1 U21747 ( .A1(n18677), .A2(n18683), .B1(n18818), .B2(n18670), .ZN(
        n18672) );
  INV_X1 U21748 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18671) );
  NAND3_X1 U21749 ( .A1(NA), .A2(n18677), .A3(n18671), .ZN(n18676) );
  OAI211_X1 U21750 ( .C1(n18814), .C2(n18673), .A(n18672), .B(n18676), .ZN(
        P3_U3029) );
  OAI22_X1 U21751 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(n20561), .B2(n18683), .ZN(n18678)
         );
  OAI21_X1 U21752 ( .B1(P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18680) );
  NAND2_X1 U21753 ( .A1(n18805), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18675) );
  OAI211_X1 U21754 ( .C1(n18678), .C2(n18680), .A(n18674), .B(n18675), .ZN(
        P3_U3030) );
  INV_X1 U21755 ( .A(n18675), .ZN(n18679) );
  AOI21_X1 U21756 ( .B1(n18677), .B2(n18676), .A(n18679), .ZN(n18682) );
  INV_X1 U21757 ( .A(NA), .ZN(n20566) );
  AOI21_X1 U21758 ( .B1(n18679), .B2(n20566), .A(n18678), .ZN(n18681) );
  OAI22_X1 U21759 ( .A1(n18682), .A2(n18683), .B1(n18681), .B2(n18680), .ZN(
        P3_U3031) );
  NAND2_X2 U21760 ( .A1(n18817), .A2(n18683), .ZN(n18739) );
  OAI222_X1 U21761 ( .A1(n18685), .A2(n18743), .B1(n18684), .B2(n18817), .C1(
        n18686), .C2(n18739), .ZN(P3_U3032) );
  OAI222_X1 U21762 ( .A1(n18739), .A2(n18688), .B1(n18687), .B2(n18817), .C1(
        n18686), .C2(n18743), .ZN(P3_U3033) );
  OAI222_X1 U21763 ( .A1(n18739), .A2(n18690), .B1(n18689), .B2(n18817), .C1(
        n18688), .C2(n18743), .ZN(P3_U3034) );
  INV_X1 U21764 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18692) );
  OAI222_X1 U21765 ( .A1(n18739), .A2(n18692), .B1(n18691), .B2(n18817), .C1(
        n18690), .C2(n18743), .ZN(P3_U3035) );
  OAI222_X1 U21766 ( .A1(n18739), .A2(n18694), .B1(n18693), .B2(n18817), .C1(
        n18692), .C2(n18743), .ZN(P3_U3036) );
  OAI222_X1 U21767 ( .A1(n18739), .A2(n20777), .B1(n18695), .B2(n18817), .C1(
        n18694), .C2(n18743), .ZN(P3_U3037) );
  OAI222_X1 U21768 ( .A1(n20777), .A2(n18743), .B1(n18696), .B2(n18817), .C1(
        n18698), .C2(n18739), .ZN(P3_U3038) );
  OAI222_X1 U21769 ( .A1(n18698), .A2(n18743), .B1(n18697), .B2(n18817), .C1(
        n18699), .C2(n18739), .ZN(P3_U3039) );
  INV_X1 U21770 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18701) );
  OAI222_X1 U21771 ( .A1(n18739), .A2(n18701), .B1(n18700), .B2(n18817), .C1(
        n18699), .C2(n18743), .ZN(P3_U3040) );
  OAI222_X1 U21772 ( .A1(n18739), .A2(n18703), .B1(n18702), .B2(n18817), .C1(
        n18701), .C2(n18743), .ZN(P3_U3041) );
  OAI222_X1 U21773 ( .A1(n18739), .A2(n18705), .B1(n18704), .B2(n18817), .C1(
        n18703), .C2(n18743), .ZN(P3_U3042) );
  OAI222_X1 U21774 ( .A1(n18739), .A2(n18707), .B1(n18706), .B2(n18817), .C1(
        n18705), .C2(n18743), .ZN(P3_U3043) );
  OAI222_X1 U21775 ( .A1(n18739), .A2(n18710), .B1(n18708), .B2(n18817), .C1(
        n18707), .C2(n18743), .ZN(P3_U3044) );
  OAI222_X1 U21776 ( .A1(n18710), .A2(n18743), .B1(n18709), .B2(n18817), .C1(
        n18711), .C2(n18739), .ZN(P3_U3045) );
  OAI222_X1 U21777 ( .A1(n18739), .A2(n18713), .B1(n18712), .B2(n18817), .C1(
        n18711), .C2(n18743), .ZN(P3_U3046) );
  OAI222_X1 U21778 ( .A1(n18739), .A2(n18716), .B1(n18714), .B2(n18817), .C1(
        n18713), .C2(n18743), .ZN(P3_U3047) );
  OAI222_X1 U21779 ( .A1(n18716), .A2(n18743), .B1(n18715), .B2(n18817), .C1(
        n18717), .C2(n18739), .ZN(P3_U3048) );
  OAI222_X1 U21780 ( .A1(n18739), .A2(n18719), .B1(n18718), .B2(n18817), .C1(
        n18717), .C2(n18743), .ZN(P3_U3049) );
  INV_X1 U21781 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n20738) );
  OAI222_X1 U21782 ( .A1(n18739), .A2(n20738), .B1(n20760), .B2(n18817), .C1(
        n18719), .C2(n18743), .ZN(P3_U3050) );
  OAI222_X1 U21783 ( .A1(n20738), .A2(n18743), .B1(n18720), .B2(n18817), .C1(
        n18721), .C2(n18739), .ZN(P3_U3051) );
  INV_X1 U21784 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18723) );
  OAI222_X1 U21785 ( .A1(n18739), .A2(n18723), .B1(n18722), .B2(n18817), .C1(
        n18721), .C2(n18743), .ZN(P3_U3052) );
  OAI222_X1 U21786 ( .A1(n18739), .A2(n18725), .B1(n18724), .B2(n18817), .C1(
        n18723), .C2(n18743), .ZN(P3_U3053) );
  OAI222_X1 U21787 ( .A1(n18739), .A2(n18727), .B1(n18726), .B2(n18817), .C1(
        n18725), .C2(n18743), .ZN(P3_U3054) );
  OAI222_X1 U21788 ( .A1(n18739), .A2(n18729), .B1(n18728), .B2(n18817), .C1(
        n18727), .C2(n18743), .ZN(P3_U3055) );
  OAI222_X1 U21789 ( .A1(n18739), .A2(n18731), .B1(n18730), .B2(n18817), .C1(
        n18729), .C2(n18743), .ZN(P3_U3056) );
  OAI222_X1 U21790 ( .A1(n18739), .A2(n18733), .B1(n18732), .B2(n18817), .C1(
        n18731), .C2(n18743), .ZN(P3_U3057) );
  INV_X1 U21791 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18736) );
  OAI222_X1 U21792 ( .A1(n18739), .A2(n18736), .B1(n18734), .B2(n18817), .C1(
        n18733), .C2(n18743), .ZN(P3_U3058) );
  OAI222_X1 U21793 ( .A1(n18736), .A2(n18743), .B1(n18735), .B2(n18817), .C1(
        n18737), .C2(n18739), .ZN(P3_U3059) );
  OAI222_X1 U21794 ( .A1(n18739), .A2(n18742), .B1(n18738), .B2(n18817), .C1(
        n18737), .C2(n18743), .ZN(P3_U3060) );
  OAI222_X1 U21795 ( .A1(n18743), .A2(n18742), .B1(n18741), .B2(n18817), .C1(
        n18740), .C2(n18739), .ZN(P3_U3061) );
  OAI22_X1 U21796 ( .A1(n18818), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18817), .ZN(n18744) );
  INV_X1 U21797 ( .A(n18744), .ZN(P3_U3274) );
  INV_X1 U21798 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18787) );
  INV_X1 U21799 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n20791) );
  AOI22_X1 U21800 ( .A1(n18817), .A2(n18787), .B1(n20791), .B2(n18818), .ZN(
        P3_U3275) );
  OAI22_X1 U21801 ( .A1(n18818), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18817), .ZN(n18745) );
  INV_X1 U21802 ( .A(n18745), .ZN(P3_U3276) );
  OAI22_X1 U21803 ( .A1(n18818), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18817), .ZN(n18746) );
  INV_X1 U21804 ( .A(n18746), .ZN(P3_U3277) );
  OAI21_X1 U21805 ( .B1(n18750), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18748), 
        .ZN(n18747) );
  INV_X1 U21806 ( .A(n18747), .ZN(P3_U3280) );
  OAI21_X1 U21807 ( .B1(n18750), .B2(n18749), .A(n18748), .ZN(P3_U3281) );
  OAI21_X1 U21808 ( .B1(n18753), .B2(n18752), .A(n18751), .ZN(P3_U3282) );
  INV_X1 U21809 ( .A(n18782), .ZN(n18785) );
  INV_X1 U21810 ( .A(n18754), .ZN(n18757) );
  NOR2_X1 U21811 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18766), .ZN(
        n18756) );
  AOI22_X1 U21812 ( .A1(n18779), .A2(n18757), .B1(n18756), .B2(n18755), .ZN(
        n18760) );
  AOI21_X1 U21813 ( .B1(n18821), .B2(n18758), .A(n18785), .ZN(n18759) );
  OAI22_X1 U21814 ( .A1(n18785), .A2(n18760), .B1(n18759), .B2(n20789), .ZN(
        P3_U3285) );
  OAI22_X1 U21815 ( .A1(n18762), .A2(n18761), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18774) );
  INV_X1 U21816 ( .A(n18774), .ZN(n18769) );
  NOR2_X1 U21817 ( .A1(n18763), .A2(n18781), .ZN(n18773) );
  OAI22_X1 U21818 ( .A1(n18767), .A2(n18766), .B1(n18765), .B2(n18764), .ZN(
        n18768) );
  AOI21_X1 U21819 ( .B1(n18769), .B2(n18773), .A(n18768), .ZN(n18770) );
  AOI22_X1 U21820 ( .A1(n18785), .A2(n18771), .B1(n18770), .B2(n18782), .ZN(
        P3_U3288) );
  INV_X1 U21821 ( .A(n18772), .ZN(n18776) );
  AOI222_X1 U21822 ( .A1(n18776), .A2(n18821), .B1(n18779), .B2(n18775), .C1(
        n18774), .C2(n18773), .ZN(n18777) );
  AOI22_X1 U21823 ( .A1(n18785), .A2(n18778), .B1(n18777), .B2(n18782), .ZN(
        P3_U3289) );
  AOI222_X1 U21824 ( .A1(n18781), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18821), 
        .B2(n18780), .C1(n18784), .C2(n18779), .ZN(n18783) );
  AOI22_X1 U21825 ( .A1(n18785), .A2(n18784), .B1(n18783), .B2(n18782), .ZN(
        P3_U3290) );
  AOI211_X1 U21826 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_REIP_REG_1__SCAN_IN), .B(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18786) );
  AOI21_X1 U21827 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18786), .ZN(n18788) );
  AOI22_X1 U21828 ( .A1(n18792), .A2(n18788), .B1(n18787), .B2(n18789), .ZN(
        P3_U3292) );
  NOR2_X1 U21829 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n18791) );
  INV_X1 U21830 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18790) );
  AOI22_X1 U21831 ( .A1(n18792), .A2(n18791), .B1(n18790), .B2(n18789), .ZN(
        P3_U3293) );
  INV_X1 U21832 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18824) );
  OAI22_X1 U21833 ( .A1(n18818), .A2(n18824), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n18817), .ZN(n18793) );
  INV_X1 U21834 ( .A(n18793), .ZN(P3_U3294) );
  INV_X1 U21835 ( .A(P3_MORE_REG_SCAN_IN), .ZN(n18802) );
  OAI22_X1 U21836 ( .A1(n18797), .A2(n18796), .B1(n18795), .B2(n18794), .ZN(
        n18799) );
  OAI21_X1 U21837 ( .B1(n18799), .B2(n18798), .A(n18801), .ZN(n18800) );
  OAI21_X1 U21838 ( .B1(n18802), .B2(n18801), .A(n18800), .ZN(P3_U3295) );
  OAI21_X1 U21839 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18804), .A(n18803), 
        .ZN(n18806) );
  AOI211_X1 U21840 ( .C1(n18822), .C2(n18806), .A(n18805), .B(n18820), .ZN(
        n18809) );
  OAI21_X1 U21841 ( .B1(n18809), .B2(n18808), .A(n18807), .ZN(n18816) );
  OAI21_X1 U21842 ( .B1(n18812), .B2(n18811), .A(n18810), .ZN(n18813) );
  AOI21_X1 U21843 ( .B1(n17394), .B2(n18814), .A(n18813), .ZN(n18815) );
  MUX2_X1 U21844 ( .A(n18816), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n18815), 
        .Z(P3_U3296) );
  OAI22_X1 U21845 ( .A1(n18818), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18817), .ZN(n18819) );
  INV_X1 U21846 ( .A(n18819), .ZN(P3_U3297) );
  AOI21_X1 U21847 ( .B1(n18821), .B2(n18820), .A(n18823), .ZN(n18827) );
  AOI22_X1 U21848 ( .A1(n18827), .A2(n18824), .B1(n18823), .B2(n18822), .ZN(
        P3_U3298) );
  INV_X1 U21849 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18826) );
  AOI21_X1 U21850 ( .B1(n18827), .B2(n18826), .A(n18825), .ZN(P3_U3299) );
  NAND2_X1 U21851 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19649), .ZN(n19639) );
  AOI22_X1 U21852 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19639), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n19633), .ZN(n19705) );
  AOI21_X1 U21853 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19705), .ZN(n18828) );
  INV_X1 U21854 ( .A(n18828), .ZN(P2_U2815) );
  INV_X1 U21855 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n20695) );
  OAI22_X1 U21856 ( .A1(n19758), .A2(n20695), .B1(n18830), .B2(n18829), .ZN(
        P2_U2816) );
  OR2_X1 U21857 ( .A1(n19641), .A2(n19776), .ZN(n19636) );
  AOI21_X1 U21858 ( .B1(n19633), .B2(n19636), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18831) );
  AOI21_X1 U21859 ( .B1(n19776), .B2(P2_CODEFETCH_REG_SCAN_IN), .A(n18831), 
        .ZN(P2_U2817) );
  OAI21_X1 U21860 ( .B1(n19641), .B2(BS16), .A(n19705), .ZN(n19703) );
  OAI21_X1 U21861 ( .B1(n19705), .B2(n11212), .A(n19703), .ZN(P2_U2818) );
  NOR2_X1 U21862 ( .A1(n18833), .A2(n18832), .ZN(n19753) );
  OAI21_X1 U21863 ( .B1(n19753), .B2(n18835), .A(n18834), .ZN(P2_U2819) );
  NOR2_X1 U21864 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20822) );
  AOI211_X1 U21865 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_12__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18836) );
  INV_X1 U21866 ( .A(P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20728) );
  INV_X1 U21867 ( .A(P2_DATAWIDTH_REG_13__SCAN_IN), .ZN(n20686) );
  AND4_X1 U21868 ( .A1(n20822), .A2(n18836), .A3(n20728), .A4(n20686), .ZN(
        n18844) );
  NOR4_X1 U21869 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n18843) );
  NOR4_X1 U21870 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n18842) );
  NOR4_X1 U21871 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18840) );
  NOR4_X1 U21872 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_15__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18839) );
  NOR4_X1 U21873 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18838) );
  NOR4_X1 U21874 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18837) );
  AND4_X1 U21875 ( .A1(n18840), .A2(n18839), .A3(n18838), .A4(n18837), .ZN(
        n18841) );
  NAND4_X1 U21876 ( .A1(n18844), .A2(n18843), .A3(n18842), .A4(n18841), .ZN(
        n18853) );
  NOR2_X1 U21877 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18853), .ZN(n18847) );
  INV_X1 U21878 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18845) );
  AOI22_X1 U21879 ( .A1(n18847), .A2(n18848), .B1(n18853), .B2(n18845), .ZN(
        P2_U2820) );
  OR3_X1 U21880 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18852) );
  INV_X1 U21881 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18846) );
  AOI22_X1 U21882 ( .A1(n18847), .A2(n18852), .B1(n18853), .B2(n18846), .ZN(
        P2_U2821) );
  INV_X1 U21883 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19704) );
  NAND2_X1 U21884 ( .A1(n18847), .A2(n19704), .ZN(n18851) );
  INV_X1 U21885 ( .A(n18853), .ZN(n18855) );
  OAI21_X1 U21886 ( .B1(n18848), .B2(n20772), .A(n18855), .ZN(n18849) );
  OAI21_X1 U21887 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18855), .A(n18849), 
        .ZN(n18850) );
  OAI221_X1 U21888 ( .B1(n18851), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18851), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18850), .ZN(P2_U2822) );
  INV_X1 U21889 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18854) );
  OAI221_X1 U21890 ( .B1(n18855), .B2(n18854), .C1(n18853), .C2(n18852), .A(
        n18851), .ZN(P2_U2823) );
  AOI22_X1 U21891 ( .A1(n18856), .A2(n18923), .B1(P2_REIP_REG_20__SCAN_IN), 
        .B2(n18940), .ZN(n18867) );
  AOI22_X1 U21892 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18931), .B1(
        P2_EBX_REG_20__SCAN_IN), .B2(n18922), .ZN(n18866) );
  INV_X1 U21893 ( .A(n18857), .ZN(n18858) );
  OAI22_X1 U21894 ( .A1(n18859), .A2(n18946), .B1(n18858), .B2(n18947), .ZN(
        n18860) );
  INV_X1 U21895 ( .A(n18860), .ZN(n18865) );
  OAI211_X1 U21896 ( .C1(n18863), .C2(n18862), .A(n18949), .B(n18861), .ZN(
        n18864) );
  NAND4_X1 U21897 ( .A1(n18867), .A2(n18866), .A3(n18865), .A4(n18864), .ZN(
        P2_U2835) );
  AOI22_X1 U21898 ( .A1(n18868), .A2(n18923), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n18922), .ZN(n18869) );
  OAI211_X1 U21899 ( .C1(n19673), .C2(n18927), .A(n18869), .B(n18925), .ZN(
        n18870) );
  AOI21_X1 U21900 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18931), .A(
        n18870), .ZN(n18879) );
  OAI22_X1 U21901 ( .A1(n18872), .A2(n18946), .B1(n18871), .B2(n18947), .ZN(
        n18873) );
  INV_X1 U21902 ( .A(n18873), .ZN(n18878) );
  OAI211_X1 U21903 ( .C1(n18876), .C2(n18875), .A(n18949), .B(n18874), .ZN(
        n18877) );
  NAND3_X1 U21904 ( .A1(n18879), .A2(n18878), .A3(n18877), .ZN(P2_U2837) );
  AOI22_X1 U21905 ( .A1(P2_EBX_REG_16__SCAN_IN), .A2(n18922), .B1(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18931), .ZN(n18880) );
  OAI21_X1 U21906 ( .B1(n18881), .B2(n18936), .A(n18880), .ZN(n18882) );
  AOI211_X1 U21907 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n18940), .A(n18939), 
        .B(n18882), .ZN(n18891) );
  NOR2_X1 U21908 ( .A1(n18883), .A2(n18947), .ZN(n18884) );
  AOI21_X1 U21909 ( .B1(n18885), .B2(n18902), .A(n18884), .ZN(n18890) );
  OAI211_X1 U21910 ( .C1(n18888), .C2(n18887), .A(n18949), .B(n18886), .ZN(
        n18889) );
  NAND3_X1 U21911 ( .A1(n18891), .A2(n18890), .A3(n18889), .ZN(P2_U2839) );
  NAND2_X1 U21912 ( .A1(n18893), .A2(n18892), .ZN(n18894) );
  XOR2_X1 U21913 ( .A(n18895), .B(n18894), .Z(n18906) );
  OAI21_X1 U21914 ( .B1(n19666), .B2(n18927), .A(n18925), .ZN(n18899) );
  OAI22_X1 U21915 ( .A1(n18897), .A2(n18936), .B1(n18896), .B2(n18954), .ZN(
        n18898) );
  AOI211_X1 U21916 ( .C1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n18931), .A(
        n18899), .B(n18898), .ZN(n18905) );
  INV_X1 U21917 ( .A(n18900), .ZN(n18903) );
  AOI22_X1 U21918 ( .A1(n18903), .A2(n18902), .B1(n18962), .B2(n18901), .ZN(
        n18904) );
  OAI211_X1 U21919 ( .C1(n19628), .C2(n18906), .A(n18905), .B(n18904), .ZN(
        P2_U2841) );
  INV_X1 U21920 ( .A(n18907), .ZN(n18908) );
  OAI22_X1 U21921 ( .A1(n18908), .A2(n18936), .B1(n11151), .B2(n18954), .ZN(
        n18909) );
  AOI211_X1 U21922 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n18940), .A(n18939), 
        .B(n18909), .ZN(n18917) );
  NOR2_X1 U21923 ( .A1(n18942), .A2(n18910), .ZN(n18911) );
  XNOR2_X1 U21924 ( .A(n18912), .B(n18911), .ZN(n18915) );
  OAI22_X1 U21925 ( .A1(n18913), .A2(n18946), .B1(n18967), .B2(n18947), .ZN(
        n18914) );
  AOI21_X1 U21926 ( .B1(n18915), .B2(n18949), .A(n18914), .ZN(n18916) );
  OAI211_X1 U21927 ( .C1(n18918), .C2(n18935), .A(n18917), .B(n18916), .ZN(
        P2_U2842) );
  NOR2_X1 U21928 ( .A1(n18942), .A2(n18919), .ZN(n18920) );
  XOR2_X1 U21929 ( .A(n18921), .B(n18920), .Z(n18933) );
  AOI22_X1 U21930 ( .A1(n18924), .A2(n18923), .B1(P2_EBX_REG_9__SCAN_IN), .B2(
        n18922), .ZN(n18926) );
  OAI211_X1 U21931 ( .C1(n12742), .C2(n18927), .A(n18926), .B(n18925), .ZN(
        n18930) );
  OAI22_X1 U21932 ( .A1(n18928), .A2(n18946), .B1(n18947), .B2(n18977), .ZN(
        n18929) );
  AOI211_X1 U21933 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n18931), .A(
        n18930), .B(n18929), .ZN(n18932) );
  OAI21_X1 U21934 ( .B1(n19628), .B2(n18933), .A(n18932), .ZN(P2_U2846) );
  OAI22_X1 U21935 ( .A1(n18937), .A2(n18936), .B1(n18935), .B2(n18934), .ZN(
        n18938) );
  AOI211_X1 U21936 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n18940), .A(n18939), .B(
        n18938), .ZN(n18952) );
  NOR2_X1 U21937 ( .A1(n18942), .A2(n18941), .ZN(n18943) );
  XNOR2_X1 U21938 ( .A(n18944), .B(n18943), .ZN(n18950) );
  OAI22_X1 U21939 ( .A1(n18993), .A2(n18947), .B1(n18946), .B2(n18945), .ZN(
        n18948) );
  AOI21_X1 U21940 ( .B1(n18950), .B2(n18949), .A(n18948), .ZN(n18951) );
  OAI211_X1 U21941 ( .C1(n18954), .C2(n18953), .A(n18952), .B(n18951), .ZN(
        P2_U2850) );
  AOI22_X1 U21942 ( .A1(n18956), .A2(n19016), .B1(n18955), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n18959) );
  AOI22_X1 U21943 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19015), .B1(n18957), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n18958) );
  NAND2_X1 U21944 ( .A1(n18959), .A2(n18958), .ZN(P2_U2888) );
  INV_X1 U21945 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19025) );
  OAI222_X1 U21946 ( .A1(n18961), .A2(n18994), .B1(n19025), .B2(n19014), .C1(
        n18960), .C2(n19022), .ZN(P2_U2904) );
  INV_X1 U21947 ( .A(n18962), .ZN(n18965) );
  AOI22_X1 U21948 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19015), .B1(n18963), 
        .B2(n19012), .ZN(n18964) );
  OAI21_X1 U21949 ( .B1(n18994), .B2(n18965), .A(n18964), .ZN(P2_U2905) );
  INV_X1 U21950 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19029) );
  OAI222_X1 U21951 ( .A1(n18967), .A2(n18994), .B1(n19029), .B2(n19014), .C1(
        n19022), .C2(n18966), .ZN(P2_U2906) );
  INV_X1 U21952 ( .A(n18968), .ZN(n18970) );
  INV_X1 U21953 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19031) );
  OAI222_X1 U21954 ( .A1(n18970), .A2(n18994), .B1(n19031), .B2(n19014), .C1(
        n19022), .C2(n18969), .ZN(P2_U2907) );
  INV_X1 U21955 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19033) );
  OAI222_X1 U21956 ( .A1(n18972), .A2(n18994), .B1(n19033), .B2(n19014), .C1(
        n19022), .C2(n18971), .ZN(P2_U2908) );
  INV_X1 U21957 ( .A(n18973), .ZN(n18975) );
  INV_X1 U21958 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19035) );
  OAI222_X1 U21959 ( .A1(n18975), .A2(n18994), .B1(n19035), .B2(n19014), .C1(
        n19022), .C2(n18974), .ZN(P2_U2909) );
  INV_X1 U21960 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19037) );
  OAI222_X1 U21961 ( .A1(n18977), .A2(n18994), .B1(n19037), .B2(n19014), .C1(
        n19022), .C2(n18976), .ZN(P2_U2910) );
  AOI22_X1 U21962 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19015), .B1(n18978), .B2(
        n19012), .ZN(n18979) );
  OAI21_X1 U21963 ( .B1(n18994), .B2(n18980), .A(n18979), .ZN(P2_U2911) );
  INV_X1 U21964 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19041) );
  OAI222_X1 U21965 ( .A1(n18982), .A2(n18994), .B1(n19041), .B2(n19014), .C1(
        n19022), .C2(n18981), .ZN(P2_U2912) );
  INV_X1 U21966 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19043) );
  OAI222_X1 U21967 ( .A1(n18983), .A2(n18994), .B1(n19043), .B2(n19014), .C1(
        n19022), .C2(n19125), .ZN(P2_U2913) );
  AOI22_X1 U21968 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19015), .B1(n18984), .B2(
        n19012), .ZN(n18992) );
  INV_X1 U21969 ( .A(n18985), .ZN(n19710) );
  XNOR2_X1 U21970 ( .A(n19711), .B(n18985), .ZN(n19004) );
  NAND2_X1 U21971 ( .A1(n19721), .A2(n18986), .ZN(n18988) );
  NAND2_X1 U21972 ( .A1(n18988), .A2(n18987), .ZN(n19003) );
  NAND2_X1 U21973 ( .A1(n19004), .A2(n19003), .ZN(n19002) );
  OAI21_X1 U21974 ( .B1(n19711), .B2(n19710), .A(n19002), .ZN(n18989) );
  NAND2_X1 U21975 ( .A1(n18989), .A2(n18995), .ZN(n18998) );
  INV_X1 U21976 ( .A(n18997), .ZN(n18990) );
  NAND3_X1 U21977 ( .A1(n18998), .A2(n18990), .A3(n19017), .ZN(n18991) );
  OAI211_X1 U21978 ( .C1(n18994), .C2(n18993), .A(n18992), .B(n18991), .ZN(
        P2_U2914) );
  INV_X1 U21979 ( .A(n18995), .ZN(n18996) );
  AOI22_X1 U21980 ( .A1(n19016), .A2(n18996), .B1(n19015), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n19001) );
  XNOR2_X1 U21981 ( .A(n18998), .B(n18997), .ZN(n18999) );
  NAND2_X1 U21982 ( .A1(n18999), .A2(n19017), .ZN(n19000) );
  OAI211_X1 U21983 ( .C1(n19115), .C2(n19022), .A(n19001), .B(n19000), .ZN(
        P2_U2915) );
  OAI21_X1 U21984 ( .B1(n19004), .B2(n19003), .A(n19002), .ZN(n19005) );
  NAND2_X1 U21985 ( .A1(n19005), .A2(n19017), .ZN(n19007) );
  AOI22_X1 U21986 ( .A1(n19710), .A2(n19016), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19015), .ZN(n19006) );
  OAI211_X1 U21987 ( .C1(n19110), .C2(n19022), .A(n19007), .B(n19006), .ZN(
        P2_U2916) );
  INV_X1 U21988 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19053) );
  OAI21_X1 U21989 ( .B1(n19009), .B2(n19018), .A(n19008), .ZN(n19010) );
  AOI222_X1 U21990 ( .A1(n19012), .A2(n19011), .B1(n19016), .B2(n19727), .C1(
        n19010), .C2(n19017), .ZN(n19013) );
  OAI21_X1 U21991 ( .B1(n19014), .B2(n19053), .A(n19013), .ZN(P2_U2918) );
  AOI22_X1 U21992 ( .A1(n19016), .A2(n19019), .B1(n19015), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n19021) );
  OAI211_X1 U21993 ( .C1(n19144), .C2(n19019), .A(n19018), .B(n19017), .ZN(
        n19020) );
  OAI211_X1 U21994 ( .C1(n19086), .C2(n19022), .A(n19021), .B(n19020), .ZN(
        P2_U2919) );
  AOI22_X1 U21995 ( .A1(n19757), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19024) );
  OAI21_X1 U21996 ( .B1(n19025), .B2(n19056), .A(n19024), .ZN(P2_U2936) );
  AOI22_X1 U21997 ( .A1(n19757), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19026) );
  OAI21_X1 U21998 ( .B1(n19027), .B2(n19056), .A(n19026), .ZN(P2_U2937) );
  AOI22_X1 U21999 ( .A1(n19757), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19028) );
  OAI21_X1 U22000 ( .B1(n19029), .B2(n19056), .A(n19028), .ZN(P2_U2938) );
  AOI22_X1 U22001 ( .A1(n19757), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19030) );
  OAI21_X1 U22002 ( .B1(n19031), .B2(n19056), .A(n19030), .ZN(P2_U2939) );
  AOI22_X1 U22003 ( .A1(n19757), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19032) );
  OAI21_X1 U22004 ( .B1(n19033), .B2(n19056), .A(n19032), .ZN(P2_U2940) );
  AOI22_X1 U22005 ( .A1(n19757), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19034) );
  OAI21_X1 U22006 ( .B1(n19035), .B2(n19056), .A(n19034), .ZN(P2_U2941) );
  AOI22_X1 U22007 ( .A1(n19757), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19036) );
  OAI21_X1 U22008 ( .B1(n19037), .B2(n19056), .A(n19036), .ZN(P2_U2942) );
  AOI22_X1 U22009 ( .A1(n19757), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19038) );
  OAI21_X1 U22010 ( .B1(n19039), .B2(n19056), .A(n19038), .ZN(P2_U2943) );
  AOI22_X1 U22011 ( .A1(n19757), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19040) );
  OAI21_X1 U22012 ( .B1(n19041), .B2(n19056), .A(n19040), .ZN(P2_U2944) );
  AOI22_X1 U22013 ( .A1(n19757), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19042) );
  OAI21_X1 U22014 ( .B1(n19043), .B2(n19056), .A(n19042), .ZN(P2_U2945) );
  INV_X1 U22015 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19045) );
  AOI22_X1 U22016 ( .A1(n19757), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19044) );
  OAI21_X1 U22017 ( .B1(n19045), .B2(n19056), .A(n19044), .ZN(P2_U2946) );
  INV_X1 U22018 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19047) );
  AOI22_X1 U22019 ( .A1(n19757), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19046) );
  OAI21_X1 U22020 ( .B1(n19047), .B2(n19056), .A(n19046), .ZN(P2_U2947) );
  INV_X1 U22021 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19049) );
  AOI22_X1 U22022 ( .A1(n19757), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19048) );
  OAI21_X1 U22023 ( .B1(n19049), .B2(n19056), .A(n19048), .ZN(P2_U2948) );
  INV_X1 U22024 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19051) );
  AOI22_X1 U22025 ( .A1(n19757), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19050) );
  OAI21_X1 U22026 ( .B1(n19051), .B2(n19056), .A(n19050), .ZN(P2_U2949) );
  AOI22_X1 U22027 ( .A1(n19757), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19052) );
  OAI21_X1 U22028 ( .B1(n19053), .B2(n19056), .A(n19052), .ZN(P2_U2950) );
  INV_X1 U22029 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19057) );
  AOI22_X1 U22030 ( .A1(n19757), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19054), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19055) );
  OAI21_X1 U22031 ( .B1(n19057), .B2(n19056), .A(n19055), .ZN(P2_U2951) );
  AOI22_X1 U22032 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n13328), .B1(n19059), 
        .B2(n19058), .ZN(n19066) );
  INV_X1 U22033 ( .A(n19060), .ZN(n19062) );
  OAI22_X1 U22034 ( .A1(n19062), .A2(n19075), .B1(n19061), .B2(n19072), .ZN(
        n19063) );
  AOI21_X1 U22035 ( .B1(n19078), .B2(n19064), .A(n19063), .ZN(n19065) );
  OAI211_X1 U22036 ( .C1(n19068), .C2(n19067), .A(n19066), .B(n19065), .ZN(
        P2_U3010) );
  OAI21_X1 U22037 ( .B1(n19070), .B2(n19069), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19081) );
  NOR2_X1 U22038 ( .A1(n19072), .A2(n19071), .ZN(n19077) );
  OAI21_X1 U22039 ( .B1(n19075), .B2(n19074), .A(n19073), .ZN(n19076) );
  AOI211_X1 U22040 ( .C1(n19079), .C2(n19078), .A(n19077), .B(n19076), .ZN(
        n19080) );
  NAND2_X1 U22041 ( .A1(n19081), .A2(n19080), .ZN(P2_U3014) );
  NAND2_X1 U22042 ( .A1(n19085), .A2(n19166), .ZN(n19082) );
  AOI21_X1 U22043 ( .B1(n19082), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19714), 
        .ZN(n19088) );
  NOR2_X1 U22044 ( .A1(n19348), .A2(n19197), .ZN(n19131) );
  INV_X1 U22045 ( .A(n19131), .ZN(n19083) );
  AND2_X1 U22046 ( .A1(n19570), .A2(n19083), .ZN(n19091) );
  AOI22_X2 U22047 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19126), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n19127), .ZN(n19578) );
  INV_X1 U22048 ( .A(n19578), .ZN(n19466) );
  NOR2_X2 U22049 ( .A1(n19765), .A2(n19108), .ZN(n19566) );
  AOI22_X1 U22050 ( .A1(n19466), .A2(n19618), .B1(n19566), .B2(n19131), .ZN(
        n19096) );
  INV_X1 U22051 ( .A(n19088), .ZN(n19092) );
  OAI21_X1 U22052 ( .B1(n19089), .B2(n19131), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19090) );
  OAI22_X2 U22053 ( .A1(n19094), .A2(n19117), .B1(n19093), .B2(n19116), .ZN(
        n19575) );
  AOI22_X1 U22054 ( .A1(n19087), .A2(n19132), .B1(n19156), .B2(n19575), .ZN(
        n19095) );
  OAI211_X1 U22055 ( .C1(n19135), .C2(n19097), .A(n19096), .B(n19095), .ZN(
        P2_U3048) );
  INV_X1 U22056 ( .A(n19583), .ZN(n19532) );
  NOR2_X2 U22057 ( .A1(n12687), .A2(n19108), .ZN(n19579) );
  AOI22_X1 U22058 ( .A1(n19532), .A2(n19618), .B1(n19579), .B2(n19131), .ZN(
        n19101) );
  AOI22_X1 U22059 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19127), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19126), .ZN(n19535) );
  AOI22_X1 U22060 ( .A1(n19099), .A2(n19132), .B1(n19156), .B2(n19580), .ZN(
        n19100) );
  OAI211_X1 U22061 ( .C1(n19135), .C2(n12486), .A(n19101), .B(n19100), .ZN(
        P2_U3049) );
  NOR2_X2 U22062 ( .A1(n19103), .A2(n19108), .ZN(n19584) );
  AOI22_X1 U22063 ( .A1(n19499), .A2(n19618), .B1(n19584), .B2(n19131), .ZN(
        n19106) );
  NOR2_X2 U22064 ( .A1(n19104), .A2(n19523), .ZN(n19585) );
  AOI22_X1 U22065 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19127), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19126), .ZN(n19502) );
  AOI22_X1 U22066 ( .A1(n19585), .A2(n19132), .B1(n19156), .B2(n19586), .ZN(
        n19105) );
  OAI211_X1 U22067 ( .C1(n19135), .C2(n10706), .A(n19106), .B(n19105), .ZN(
        P2_U3050) );
  NOR2_X2 U22068 ( .A1(n19109), .A2(n19108), .ZN(n19590) );
  AOI22_X1 U22069 ( .A1(n19538), .A2(n19618), .B1(n19590), .B2(n19131), .ZN(
        n19113) );
  AOI22_X1 U22070 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19127), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19126), .ZN(n19541) );
  AOI22_X1 U22071 ( .A1(n19111), .A2(n19132), .B1(n19156), .B2(n19591), .ZN(
        n19112) );
  OAI211_X1 U22072 ( .C1(n19135), .C2(n19114), .A(n19113), .B(n19112), .ZN(
        P2_U3051) );
  INV_X1 U22073 ( .A(n19600), .ZN(n19505) );
  AOI22_X1 U22074 ( .A1(n19505), .A2(n19618), .B1(n19595), .B2(n19131), .ZN(
        n19120) );
  NOR2_X2 U22075 ( .A1(n19115), .A2(n19523), .ZN(n19596) );
  OAI22_X2 U22076 ( .A1(n19118), .A2(n19117), .B1(n20687), .B2(n19116), .ZN(
        n19597) );
  AOI22_X1 U22077 ( .A1(n19596), .A2(n19132), .B1(n19156), .B2(n19597), .ZN(
        n19119) );
  OAI211_X1 U22078 ( .C1(n19135), .C2(n19121), .A(n19120), .B(n19119), .ZN(
        P2_U3052) );
  AOI22_X1 U22079 ( .A1(n19546), .A2(n19618), .B1(n19601), .B2(n19131), .ZN(
        n19123) );
  AOI22_X1 U22080 ( .A1(n19602), .A2(n19132), .B1(n19156), .B2(n19603), .ZN(
        n19122) );
  OAI211_X1 U22081 ( .C1(n19135), .C2(n13370), .A(n19123), .B(n19122), .ZN(
        P2_U3053) );
  AOI22_X1 U22082 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19126), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19127), .ZN(n19612) );
  AOI22_X1 U22083 ( .A1(n19618), .A2(n19550), .B1(n19607), .B2(n19131), .ZN(
        n19129) );
  NOR2_X2 U22084 ( .A1(n19125), .A2(n19523), .ZN(n19608) );
  AOI22_X1 U22085 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19127), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19126), .ZN(n19553) );
  INV_X1 U22086 ( .A(n19553), .ZN(n19609) );
  AOI22_X1 U22087 ( .A1(n19608), .A2(n19132), .B1(n19156), .B2(n19609), .ZN(
        n19128) );
  OAI211_X1 U22088 ( .C1(n19135), .C2(n19130), .A(n19129), .B(n19128), .ZN(
        P2_U3054) );
  AOI22_X1 U22089 ( .A1(n19556), .A2(n19618), .B1(n19613), .B2(n19131), .ZN(
        n19134) );
  AOI22_X1 U22090 ( .A1(n19615), .A2(n19132), .B1(n19156), .B2(n19617), .ZN(
        n19133) );
  OAI211_X1 U22091 ( .C1(n19135), .C2(n12617), .A(n19134), .B(n19133), .ZN(
        P2_U3055) );
  NAND2_X1 U22092 ( .A1(n19167), .A2(n19735), .ZN(n19140) );
  INV_X1 U22093 ( .A(n19136), .ZN(n19137) );
  NOR2_X1 U22094 ( .A1(n20827), .A2(n19140), .ZN(n19161) );
  INV_X1 U22095 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19350) );
  NOR3_X1 U22096 ( .A1(n19137), .A2(n19161), .A3(n19350), .ZN(n19139) );
  AOI211_X2 U22097 ( .C1(n19140), .C2(n19350), .A(n19321), .B(n19139), .ZN(
        n19162) );
  AOI22_X1 U22098 ( .A1(n19162), .A2(n19087), .B1(n19566), .B2(n19161), .ZN(
        n19147) );
  NAND2_X1 U22099 ( .A1(n19145), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19322) );
  INV_X1 U22100 ( .A(n19322), .ZN(n19138) );
  NAND2_X1 U22101 ( .A1(n19138), .A2(n19143), .ZN(n19141) );
  AOI21_X1 U22102 ( .B1(n19141), .B2(n19140), .A(n19139), .ZN(n19142) );
  OAI211_X1 U22103 ( .C1(n19161), .C2(n19737), .A(n19142), .B(n19573), .ZN(
        n19163) );
  AOI22_X1 U22104 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19163), .B1(
        n19188), .B2(n19575), .ZN(n19146) );
  OAI211_X1 U22105 ( .C1(n19578), .C2(n19166), .A(n19147), .B(n19146), .ZN(
        P2_U3056) );
  AOI22_X1 U22106 ( .A1(n19162), .A2(n19099), .B1(n19579), .B2(n19161), .ZN(
        n19149) );
  AOI22_X1 U22107 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19163), .B1(
        n19188), .B2(n19580), .ZN(n19148) );
  OAI211_X1 U22108 ( .C1(n19583), .C2(n19166), .A(n19149), .B(n19148), .ZN(
        P2_U3057) );
  AOI22_X1 U22109 ( .A1(n19162), .A2(n19585), .B1(n19584), .B2(n19161), .ZN(
        n19151) );
  AOI22_X1 U22110 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19163), .B1(
        n19156), .B2(n19499), .ZN(n19150) );
  OAI211_X1 U22111 ( .C1(n19502), .C2(n19196), .A(n19151), .B(n19150), .ZN(
        P2_U3058) );
  AOI22_X1 U22112 ( .A1(n19162), .A2(n19111), .B1(n19590), .B2(n19161), .ZN(
        n19153) );
  AOI22_X1 U22113 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19163), .B1(
        n19188), .B2(n19591), .ZN(n19152) );
  OAI211_X1 U22114 ( .C1(n19594), .C2(n19166), .A(n19153), .B(n19152), .ZN(
        P2_U3059) );
  AOI22_X1 U22115 ( .A1(n19162), .A2(n19596), .B1(n19595), .B2(n19161), .ZN(
        n19155) );
  AOI22_X1 U22116 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19163), .B1(
        n19188), .B2(n19597), .ZN(n19154) );
  OAI211_X1 U22117 ( .C1(n19600), .C2(n19166), .A(n19155), .B(n19154), .ZN(
        P2_U3060) );
  AOI22_X1 U22118 ( .A1(n19162), .A2(n19602), .B1(n19601), .B2(n19161), .ZN(
        n19158) );
  AOI22_X1 U22119 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19163), .B1(
        n19156), .B2(n19546), .ZN(n19157) );
  OAI211_X1 U22120 ( .C1(n19549), .C2(n19196), .A(n19158), .B(n19157), .ZN(
        P2_U3061) );
  AOI22_X1 U22121 ( .A1(n19162), .A2(n19608), .B1(n19607), .B2(n19161), .ZN(
        n19160) );
  AOI22_X1 U22122 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19163), .B1(
        n19188), .B2(n19609), .ZN(n19159) );
  OAI211_X1 U22123 ( .C1(n19612), .C2(n19166), .A(n19160), .B(n19159), .ZN(
        P2_U3062) );
  INV_X1 U22124 ( .A(n19556), .ZN(n19623) );
  AOI22_X1 U22125 ( .A1(n19162), .A2(n19615), .B1(n19613), .B2(n19161), .ZN(
        n19165) );
  AOI22_X1 U22126 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19163), .B1(
        n19188), .B2(n19617), .ZN(n19164) );
  OAI211_X1 U22127 ( .C1(n19623), .C2(n19166), .A(n19165), .B(n19164), .ZN(
        P2_U3063) );
  NAND2_X1 U22128 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19167), .ZN(
        n19203) );
  NOR2_X1 U22129 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19203), .ZN(
        n19191) );
  OAI21_X1 U22130 ( .B1(n19169), .B2(n19191), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19168) );
  OR2_X1 U22131 ( .A1(n19411), .A2(n19197), .ZN(n19172) );
  NAND2_X1 U22132 ( .A1(n19168), .A2(n19172), .ZN(n19192) );
  AOI22_X1 U22133 ( .A1(n19192), .A2(n19087), .B1(n19566), .B2(n19191), .ZN(
        n19177) );
  INV_X1 U22134 ( .A(n19169), .ZN(n19170) );
  AOI21_X1 U22135 ( .B1(n19170), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19175) );
  INV_X1 U22136 ( .A(n19707), .ZN(n19171) );
  OAI21_X1 U22137 ( .B1(n19221), .B2(n19188), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19173) );
  NAND3_X1 U22138 ( .A1(n19173), .A2(n19520), .A3(n19172), .ZN(n19174) );
  OAI211_X1 U22139 ( .C1(n19191), .C2(n19175), .A(n19174), .B(n19573), .ZN(
        n19193) );
  AOI22_X1 U22140 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19193), .B1(
        n19221), .B2(n19575), .ZN(n19176) );
  OAI211_X1 U22141 ( .C1(n19578), .C2(n19196), .A(n19177), .B(n19176), .ZN(
        P2_U3064) );
  AOI22_X1 U22142 ( .A1(n19192), .A2(n19099), .B1(n19579), .B2(n19191), .ZN(
        n19179) );
  AOI22_X1 U22143 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19193), .B1(
        n19221), .B2(n19580), .ZN(n19178) );
  OAI211_X1 U22144 ( .C1(n19583), .C2(n19196), .A(n19179), .B(n19178), .ZN(
        P2_U3065) );
  AOI22_X1 U22145 ( .A1(n19192), .A2(n19585), .B1(n19584), .B2(n19191), .ZN(
        n19181) );
  AOI22_X1 U22146 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19193), .B1(
        n19221), .B2(n19586), .ZN(n19180) );
  OAI211_X1 U22147 ( .C1(n19589), .C2(n19196), .A(n19181), .B(n19180), .ZN(
        P2_U3066) );
  AOI22_X1 U22148 ( .A1(n19192), .A2(n19111), .B1(n19590), .B2(n19191), .ZN(
        n19183) );
  AOI22_X1 U22149 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19193), .B1(
        n19221), .B2(n19591), .ZN(n19182) );
  OAI211_X1 U22150 ( .C1(n19594), .C2(n19196), .A(n19183), .B(n19182), .ZN(
        P2_U3067) );
  AOI22_X1 U22151 ( .A1(n19192), .A2(n19596), .B1(n19595), .B2(n19191), .ZN(
        n19185) );
  AOI22_X1 U22152 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19193), .B1(
        n19221), .B2(n19597), .ZN(n19184) );
  OAI211_X1 U22153 ( .C1(n19600), .C2(n19196), .A(n19185), .B(n19184), .ZN(
        P2_U3068) );
  AOI22_X1 U22154 ( .A1(n19192), .A2(n19602), .B1(n19601), .B2(n19191), .ZN(
        n19187) );
  AOI22_X1 U22155 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19193), .B1(
        n19221), .B2(n19603), .ZN(n19186) );
  OAI211_X1 U22156 ( .C1(n19606), .C2(n19196), .A(n19187), .B(n19186), .ZN(
        P2_U3069) );
  AOI22_X1 U22157 ( .A1(n19192), .A2(n19608), .B1(n19607), .B2(n19191), .ZN(
        n19190) );
  AOI22_X1 U22158 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19193), .B1(
        n19188), .B2(n19550), .ZN(n19189) );
  OAI211_X1 U22159 ( .C1(n19553), .C2(n19219), .A(n19190), .B(n19189), .ZN(
        P2_U3070) );
  AOI22_X1 U22160 ( .A1(n19192), .A2(n19615), .B1(n19613), .B2(n19191), .ZN(
        n19195) );
  AOI22_X1 U22161 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19193), .B1(
        n19221), .B2(n19617), .ZN(n19194) );
  OAI211_X1 U22162 ( .C1(n19623), .C2(n19196), .A(n19195), .B(n19194), .ZN(
        P2_U3071) );
  NOR2_X1 U22163 ( .A1(n19438), .A2(n19197), .ZN(n19220) );
  AOI22_X1 U22164 ( .A1(n19575), .A2(n19246), .B1(n19220), .B2(n19566), .ZN(
        n19206) );
  OAI21_X1 U22165 ( .B1(n19322), .B2(n19707), .A(n19520), .ZN(n19204) );
  INV_X1 U22166 ( .A(n19203), .ZN(n19200) );
  INV_X1 U22167 ( .A(n19220), .ZN(n19198) );
  OAI211_X1 U22168 ( .C1(n10792), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19198), 
        .B(n19714), .ZN(n19199) );
  OAI211_X1 U22169 ( .C1(n19204), .C2(n19200), .A(n19573), .B(n19199), .ZN(
        n19223) );
  INV_X1 U22170 ( .A(n10792), .ZN(n19201) );
  OAI21_X1 U22171 ( .B1(n19201), .B2(n19220), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19202) );
  OAI21_X1 U22172 ( .B1(n19204), .B2(n19203), .A(n19202), .ZN(n19222) );
  AOI22_X1 U22173 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19223), .B1(
        n19087), .B2(n19222), .ZN(n19205) );
  OAI211_X1 U22174 ( .C1(n19578), .C2(n19219), .A(n19206), .B(n19205), .ZN(
        P2_U3072) );
  AOI22_X1 U22175 ( .A1(n19532), .A2(n19221), .B1(n19220), .B2(n19579), .ZN(
        n19208) );
  AOI22_X1 U22176 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19223), .B1(
        n19099), .B2(n19222), .ZN(n19207) );
  OAI211_X1 U22177 ( .C1(n19535), .C2(n19254), .A(n19208), .B(n19207), .ZN(
        P2_U3073) );
  AOI22_X1 U22178 ( .A1(n19246), .A2(n19586), .B1(n19220), .B2(n19584), .ZN(
        n19210) );
  AOI22_X1 U22179 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19223), .B1(
        n19585), .B2(n19222), .ZN(n19209) );
  OAI211_X1 U22180 ( .C1(n19589), .C2(n19219), .A(n19210), .B(n19209), .ZN(
        P2_U3074) );
  AOI22_X1 U22181 ( .A1(n19538), .A2(n19221), .B1(n19220), .B2(n19590), .ZN(
        n19212) );
  AOI22_X1 U22182 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19223), .B1(
        n19111), .B2(n19222), .ZN(n19211) );
  OAI211_X1 U22183 ( .C1(n19541), .C2(n19254), .A(n19212), .B(n19211), .ZN(
        P2_U3075) );
  AOI22_X1 U22184 ( .A1(n19597), .A2(n19246), .B1(n19220), .B2(n19595), .ZN(
        n19214) );
  AOI22_X1 U22185 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19223), .B1(
        n19596), .B2(n19222), .ZN(n19213) );
  OAI211_X1 U22186 ( .C1(n19600), .C2(n19219), .A(n19214), .B(n19213), .ZN(
        P2_U3076) );
  AOI22_X1 U22187 ( .A1(n19246), .A2(n19603), .B1(n19601), .B2(n19220), .ZN(
        n19216) );
  AOI22_X1 U22188 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19223), .B1(
        n19602), .B2(n19222), .ZN(n19215) );
  OAI211_X1 U22189 ( .C1(n19606), .C2(n19219), .A(n19216), .B(n19215), .ZN(
        P2_U3077) );
  AOI22_X1 U22190 ( .A1(n19609), .A2(n19246), .B1(n19220), .B2(n19607), .ZN(
        n19218) );
  AOI22_X1 U22191 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19223), .B1(
        n19608), .B2(n19222), .ZN(n19217) );
  OAI211_X1 U22192 ( .C1(n19612), .C2(n19219), .A(n19218), .B(n19217), .ZN(
        P2_U3078) );
  AOI22_X1 U22193 ( .A1(n19556), .A2(n19221), .B1(n19613), .B2(n19220), .ZN(
        n19225) );
  AOI22_X1 U22194 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19223), .B1(
        n19615), .B2(n19222), .ZN(n19224) );
  OAI211_X1 U22195 ( .C1(n19561), .C2(n19254), .A(n19225), .B(n19224), .ZN(
        P2_U3079) );
  NAND2_X1 U22196 ( .A1(n19226), .A2(n19718), .ZN(n19232) );
  NAND2_X1 U22197 ( .A1(n19718), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19287) );
  NOR2_X1 U22198 ( .A1(n19348), .A2(n19287), .ZN(n19249) );
  OAI21_X1 U22199 ( .B1(n19229), .B2(n19249), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19227) );
  OAI21_X1 U22200 ( .B1(n19232), .B2(n19714), .A(n19227), .ZN(n19250) );
  AOI22_X1 U22201 ( .A1(n19250), .A2(n19087), .B1(n19566), .B2(n19249), .ZN(
        n19235) );
  OAI21_X1 U22202 ( .B1(n19246), .B2(n19281), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19231) );
  AOI211_X1 U22203 ( .C1(n19229), .C2(n19737), .A(n19249), .B(n19520), .ZN(
        n19230) );
  AOI211_X1 U22204 ( .C1(n19232), .C2(n19231), .A(n19523), .B(n19230), .ZN(
        n19233) );
  AOI22_X1 U22205 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19251), .B1(
        n19281), .B2(n19575), .ZN(n19234) );
  OAI211_X1 U22206 ( .C1(n19578), .C2(n19254), .A(n19235), .B(n19234), .ZN(
        P2_U3080) );
  AOI22_X1 U22207 ( .A1(n19250), .A2(n19099), .B1(n19579), .B2(n19249), .ZN(
        n19237) );
  AOI22_X1 U22208 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19251), .B1(
        n19281), .B2(n19580), .ZN(n19236) );
  OAI211_X1 U22209 ( .C1(n19583), .C2(n19254), .A(n19237), .B(n19236), .ZN(
        P2_U3081) );
  AOI22_X1 U22210 ( .A1(n19250), .A2(n19585), .B1(n19584), .B2(n19249), .ZN(
        n19239) );
  AOI22_X1 U22211 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19251), .B1(
        n19281), .B2(n19586), .ZN(n19238) );
  OAI211_X1 U22212 ( .C1(n19589), .C2(n19254), .A(n19239), .B(n19238), .ZN(
        P2_U3082) );
  AOI22_X1 U22213 ( .A1(n19250), .A2(n19111), .B1(n19590), .B2(n19249), .ZN(
        n19241) );
  AOI22_X1 U22214 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19251), .B1(
        n19281), .B2(n19591), .ZN(n19240) );
  OAI211_X1 U22215 ( .C1(n19594), .C2(n19254), .A(n19241), .B(n19240), .ZN(
        P2_U3083) );
  INV_X1 U22216 ( .A(n19597), .ZN(n19508) );
  AOI22_X1 U22217 ( .A1(n19250), .A2(n19596), .B1(n19595), .B2(n19249), .ZN(
        n19243) );
  AOI22_X1 U22218 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19251), .B1(
        n19246), .B2(n19505), .ZN(n19242) );
  OAI211_X1 U22219 ( .C1(n19508), .C2(n19275), .A(n19243), .B(n19242), .ZN(
        P2_U3084) );
  AOI22_X1 U22220 ( .A1(n19250), .A2(n19602), .B1(n19601), .B2(n19249), .ZN(
        n19245) );
  AOI22_X1 U22221 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19251), .B1(
        n19281), .B2(n19603), .ZN(n19244) );
  OAI211_X1 U22222 ( .C1(n19606), .C2(n19254), .A(n19245), .B(n19244), .ZN(
        P2_U3085) );
  AOI22_X1 U22223 ( .A1(n19250), .A2(n19608), .B1(n19607), .B2(n19249), .ZN(
        n19248) );
  AOI22_X1 U22224 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19251), .B1(
        n19246), .B2(n19550), .ZN(n19247) );
  OAI211_X1 U22225 ( .C1(n19553), .C2(n19275), .A(n19248), .B(n19247), .ZN(
        P2_U3086) );
  AOI22_X1 U22226 ( .A1(n19250), .A2(n19615), .B1(n19613), .B2(n19249), .ZN(
        n19253) );
  AOI22_X1 U22227 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19251), .B1(
        n19281), .B2(n19617), .ZN(n19252) );
  OAI211_X1 U22228 ( .C1(n19623), .C2(n19254), .A(n19253), .B(n19252), .ZN(
        P2_U3087) );
  OR2_X1 U22229 ( .A1(n19322), .A2(n19493), .ZN(n19255) );
  AND2_X1 U22230 ( .A1(n19255), .A2(n19520), .ZN(n19258) );
  INV_X1 U22231 ( .A(n19287), .ZN(n19316) );
  NAND2_X1 U22232 ( .A1(n19316), .A2(n19735), .ZN(n19261) );
  AOI21_X1 U22233 ( .B1(n10800), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19256) );
  NOR2_X1 U22234 ( .A1(n20827), .A2(n19261), .ZN(n19280) );
  OAI21_X1 U22235 ( .B1(n19256), .B2(n19280), .A(n19573), .ZN(n19257) );
  AOI21_X1 U22236 ( .B1(n19258), .B2(n19261), .A(n19257), .ZN(n19266) );
  AOI22_X1 U22237 ( .A1(n19575), .A2(n19307), .B1(n19566), .B2(n19280), .ZN(
        n19264) );
  INV_X1 U22238 ( .A(n19258), .ZN(n19262) );
  INV_X1 U22239 ( .A(n10800), .ZN(n19259) );
  OAI21_X1 U22240 ( .B1(n19259), .B2(n19280), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19260) );
  AOI22_X1 U22241 ( .A1(n19087), .A2(n19282), .B1(n19281), .B2(n19466), .ZN(
        n19263) );
  OAI211_X1 U22242 ( .C1(n19266), .C2(n19265), .A(n19264), .B(n19263), .ZN(
        P2_U3088) );
  AOI22_X1 U22243 ( .A1(n19307), .A2(n19580), .B1(n19280), .B2(n19579), .ZN(
        n19268) );
  AOI22_X1 U22244 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19283), .B1(
        n19099), .B2(n19282), .ZN(n19267) );
  OAI211_X1 U22245 ( .C1(n19583), .C2(n19275), .A(n19268), .B(n19267), .ZN(
        P2_U3089) );
  AOI22_X1 U22246 ( .A1(n19281), .A2(n19499), .B1(n19584), .B2(n19280), .ZN(
        n19270) );
  AOI22_X1 U22247 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19283), .B1(
        n19585), .B2(n19282), .ZN(n19269) );
  OAI211_X1 U22248 ( .C1(n19502), .C2(n19315), .A(n19270), .B(n19269), .ZN(
        P2_U3090) );
  AOI22_X1 U22249 ( .A1(n19281), .A2(n19538), .B1(n19280), .B2(n19590), .ZN(
        n19272) );
  AOI22_X1 U22250 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19283), .B1(
        n19111), .B2(n19282), .ZN(n19271) );
  OAI211_X1 U22251 ( .C1(n19541), .C2(n19315), .A(n19272), .B(n19271), .ZN(
        P2_U3091) );
  AOI22_X1 U22252 ( .A1(n19597), .A2(n19307), .B1(n19595), .B2(n19280), .ZN(
        n19274) );
  AOI22_X1 U22253 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19283), .B1(
        n19596), .B2(n19282), .ZN(n19273) );
  OAI211_X1 U22254 ( .C1(n19600), .C2(n19275), .A(n19274), .B(n19273), .ZN(
        P2_U3092) );
  AOI22_X1 U22255 ( .A1(n19281), .A2(n19546), .B1(n19601), .B2(n19280), .ZN(
        n19277) );
  AOI22_X1 U22256 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19283), .B1(
        n19602), .B2(n19282), .ZN(n19276) );
  OAI211_X1 U22257 ( .C1(n19549), .C2(n19315), .A(n19277), .B(n19276), .ZN(
        P2_U3093) );
  AOI22_X1 U22258 ( .A1(n19281), .A2(n19550), .B1(n19607), .B2(n19280), .ZN(
        n19279) );
  AOI22_X1 U22259 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19283), .B1(
        n19608), .B2(n19282), .ZN(n19278) );
  OAI211_X1 U22260 ( .C1(n19553), .C2(n19315), .A(n19279), .B(n19278), .ZN(
        P2_U3094) );
  AOI22_X1 U22261 ( .A1(n19281), .A2(n19556), .B1(n19613), .B2(n19280), .ZN(
        n19285) );
  AOI22_X1 U22262 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19283), .B1(
        n19615), .B2(n19282), .ZN(n19284) );
  OAI211_X1 U22263 ( .C1(n19561), .C2(n19315), .A(n19285), .B(n19284), .ZN(
        P2_U3095) );
  INV_X1 U22264 ( .A(n19562), .ZN(n19567) );
  NOR3_X2 U22265 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n19567), .ZN(n19310) );
  OAI21_X1 U22266 ( .B1(n19290), .B2(n19310), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19286) );
  OAI21_X1 U22267 ( .B1(n19287), .B2(n19411), .A(n19286), .ZN(n19311) );
  AOI22_X1 U22268 ( .A1(n19311), .A2(n19087), .B1(n19566), .B2(n19310), .ZN(
        n19296) );
  OAI21_X1 U22269 ( .B1(n19307), .B2(n19344), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19293) );
  NAND2_X1 U22270 ( .A1(n19289), .A2(n19316), .ZN(n19292) );
  AOI211_X1 U22271 ( .C1(n19290), .C2(n19737), .A(n19310), .B(n19520), .ZN(
        n19291) );
  AOI211_X1 U22272 ( .C1(n19293), .C2(n19292), .A(n19523), .B(n19291), .ZN(
        n19294) );
  AOI22_X1 U22273 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19312), .B1(
        n19344), .B2(n19575), .ZN(n19295) );
  OAI211_X1 U22274 ( .C1(n19578), .C2(n19315), .A(n19296), .B(n19295), .ZN(
        P2_U3096) );
  AOI22_X1 U22275 ( .A1(n19311), .A2(n19099), .B1(n19579), .B2(n19310), .ZN(
        n19298) );
  AOI22_X1 U22276 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19312), .B1(
        n19307), .B2(n19532), .ZN(n19297) );
  OAI211_X1 U22277 ( .C1(n19535), .C2(n19342), .A(n19298), .B(n19297), .ZN(
        P2_U3097) );
  AOI22_X1 U22278 ( .A1(n19311), .A2(n19585), .B1(n19584), .B2(n19310), .ZN(
        n19300) );
  AOI22_X1 U22279 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19312), .B1(
        n19307), .B2(n19499), .ZN(n19299) );
  OAI211_X1 U22280 ( .C1(n19502), .C2(n19342), .A(n19300), .B(n19299), .ZN(
        P2_U3098) );
  AOI22_X1 U22281 ( .A1(n19311), .A2(n19111), .B1(n19590), .B2(n19310), .ZN(
        n19302) );
  AOI22_X1 U22282 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19312), .B1(
        n19307), .B2(n19538), .ZN(n19301) );
  OAI211_X1 U22283 ( .C1(n19541), .C2(n19342), .A(n19302), .B(n19301), .ZN(
        P2_U3099) );
  AOI22_X1 U22284 ( .A1(n19311), .A2(n19596), .B1(n19595), .B2(n19310), .ZN(
        n19304) );
  AOI22_X1 U22285 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19312), .B1(
        n19344), .B2(n19597), .ZN(n19303) );
  OAI211_X1 U22286 ( .C1(n19600), .C2(n19315), .A(n19304), .B(n19303), .ZN(
        P2_U3100) );
  AOI22_X1 U22287 ( .A1(n19311), .A2(n19602), .B1(n19601), .B2(n19310), .ZN(
        n19306) );
  AOI22_X1 U22288 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19312), .B1(
        n19307), .B2(n19546), .ZN(n19305) );
  OAI211_X1 U22289 ( .C1(n19549), .C2(n19342), .A(n19306), .B(n19305), .ZN(
        P2_U3101) );
  AOI22_X1 U22290 ( .A1(n19311), .A2(n19608), .B1(n19607), .B2(n19310), .ZN(
        n19309) );
  AOI22_X1 U22291 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19312), .B1(
        n19307), .B2(n19550), .ZN(n19308) );
  OAI211_X1 U22292 ( .C1(n19553), .C2(n19342), .A(n19309), .B(n19308), .ZN(
        P2_U3102) );
  AOI22_X1 U22293 ( .A1(n19311), .A2(n19615), .B1(n19613), .B2(n19310), .ZN(
        n19314) );
  AOI22_X1 U22294 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19312), .B1(
        n19344), .B2(n19617), .ZN(n19313) );
  OAI211_X1 U22295 ( .C1(n19623), .C2(n19315), .A(n19314), .B(n19313), .ZN(
        P2_U3103) );
  OR2_X1 U22296 ( .A1(n19567), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19325) );
  INV_X1 U22297 ( .A(n19438), .ZN(n19317) );
  NAND2_X1 U22298 ( .A1(n19317), .A2(n19316), .ZN(n19352) );
  AND2_X1 U22299 ( .A1(n19352), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19318) );
  NAND2_X1 U22300 ( .A1(n19319), .A2(n19318), .ZN(n19323) );
  INV_X1 U22301 ( .A(n19323), .ZN(n19320) );
  AOI211_X2 U22302 ( .C1(n19325), .C2(n19350), .A(n19321), .B(n19320), .ZN(
        n19343) );
  AOI22_X1 U22303 ( .A1(n19343), .A2(n19087), .B1(n19355), .B2(n19566), .ZN(
        n19329) );
  OR2_X1 U22304 ( .A1(n19322), .A2(n19568), .ZN(n19715) );
  OAI211_X1 U22305 ( .C1(n19355), .C2(n19737), .A(n19323), .B(n19573), .ZN(
        n19324) );
  AOI21_X1 U22306 ( .B1(n19715), .B2(n19325), .A(n19324), .ZN(n19326) );
  AOI22_X1 U22307 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19345), .B1(
        n19371), .B2(n19575), .ZN(n19328) );
  OAI211_X1 U22308 ( .C1(n19578), .C2(n19342), .A(n19329), .B(n19328), .ZN(
        P2_U3104) );
  AOI22_X1 U22309 ( .A1(n19343), .A2(n19099), .B1(n19355), .B2(n19579), .ZN(
        n19331) );
  AOI22_X1 U22310 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19345), .B1(
        n19371), .B2(n19580), .ZN(n19330) );
  OAI211_X1 U22311 ( .C1(n19583), .C2(n19342), .A(n19331), .B(n19330), .ZN(
        P2_U3105) );
  AOI22_X1 U22312 ( .A1(n19343), .A2(n19585), .B1(n19355), .B2(n19584), .ZN(
        n19333) );
  AOI22_X1 U22313 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19345), .B1(
        n19371), .B2(n19586), .ZN(n19332) );
  OAI211_X1 U22314 ( .C1(n19589), .C2(n19342), .A(n19333), .B(n19332), .ZN(
        P2_U3106) );
  AOI22_X1 U22315 ( .A1(n19343), .A2(n19111), .B1(n19355), .B2(n19590), .ZN(
        n19335) );
  AOI22_X1 U22316 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19345), .B1(
        n19344), .B2(n19538), .ZN(n19334) );
  OAI211_X1 U22317 ( .C1(n19541), .C2(n19379), .A(n19335), .B(n19334), .ZN(
        P2_U3107) );
  AOI22_X1 U22318 ( .A1(n19343), .A2(n19596), .B1(n19355), .B2(n19595), .ZN(
        n19337) );
  AOI22_X1 U22319 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19345), .B1(
        n19371), .B2(n19597), .ZN(n19336) );
  OAI211_X1 U22320 ( .C1(n19600), .C2(n19342), .A(n19337), .B(n19336), .ZN(
        P2_U3108) );
  AOI22_X1 U22321 ( .A1(n19343), .A2(n19602), .B1(n19601), .B2(n19355), .ZN(
        n19339) );
  AOI22_X1 U22322 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19345), .B1(
        n19371), .B2(n19603), .ZN(n19338) );
  OAI211_X1 U22323 ( .C1(n19606), .C2(n19342), .A(n19339), .B(n19338), .ZN(
        P2_U3109) );
  AOI22_X1 U22324 ( .A1(n19343), .A2(n19608), .B1(n19355), .B2(n19607), .ZN(
        n19341) );
  AOI22_X1 U22325 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19345), .B1(
        n19371), .B2(n19609), .ZN(n19340) );
  OAI211_X1 U22326 ( .C1(n19612), .C2(n19342), .A(n19341), .B(n19340), .ZN(
        P2_U3110) );
  AOI22_X1 U22327 ( .A1(n19343), .A2(n19615), .B1(n19613), .B2(n19355), .ZN(
        n19347) );
  AOI22_X1 U22328 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19345), .B1(
        n19344), .B2(n19556), .ZN(n19346) );
  OAI211_X1 U22329 ( .C1(n19561), .C2(n19379), .A(n19347), .B(n19346), .ZN(
        P2_U3111) );
  NAND2_X1 U22330 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19725), .ZN(
        n19443) );
  NOR2_X1 U22331 ( .A1(n19348), .A2(n19443), .ZN(n19374) );
  AOI22_X1 U22332 ( .A1(n19575), .A2(n19404), .B1(n19566), .B2(n19374), .ZN(
        n19360) );
  NAND2_X1 U22333 ( .A1(n19401), .A2(n19379), .ZN(n19349) );
  AOI21_X1 U22334 ( .B1(n19349), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19714), 
        .ZN(n19354) );
  OAI21_X1 U22335 ( .B1(n9606), .B2(n19350), .A(n19737), .ZN(n19351) );
  AOI21_X1 U22336 ( .B1(n19354), .B2(n19352), .A(n19351), .ZN(n19353) );
  OAI21_X1 U22337 ( .B1(n19374), .B2(n19353), .A(n19573), .ZN(n19376) );
  OAI21_X1 U22338 ( .B1(n19355), .B2(n19374), .A(n19354), .ZN(n19358) );
  OAI21_X1 U22339 ( .B1(n9606), .B2(n19374), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19357) );
  NAND2_X1 U22340 ( .A1(n19358), .A2(n19357), .ZN(n19375) );
  AOI22_X1 U22341 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19376), .B1(
        n19087), .B2(n19375), .ZN(n19359) );
  OAI211_X1 U22342 ( .C1(n19578), .C2(n19379), .A(n19360), .B(n19359), .ZN(
        P2_U3112) );
  AOI22_X1 U22343 ( .A1(n19404), .A2(n19580), .B1(n19579), .B2(n19374), .ZN(
        n19362) );
  AOI22_X1 U22344 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19376), .B1(
        n19375), .B2(n19099), .ZN(n19361) );
  OAI211_X1 U22345 ( .C1(n19583), .C2(n19379), .A(n19362), .B(n19361), .ZN(
        P2_U3113) );
  AOI22_X1 U22346 ( .A1(n19404), .A2(n19586), .B1(n19584), .B2(n19374), .ZN(
        n19364) );
  AOI22_X1 U22347 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19376), .B1(
        n19375), .B2(n19585), .ZN(n19363) );
  OAI211_X1 U22348 ( .C1(n19589), .C2(n19379), .A(n19364), .B(n19363), .ZN(
        P2_U3114) );
  AOI22_X1 U22349 ( .A1(n19404), .A2(n19591), .B1(n19374), .B2(n19590), .ZN(
        n19366) );
  AOI22_X1 U22350 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19376), .B1(
        n19375), .B2(n19111), .ZN(n19365) );
  OAI211_X1 U22351 ( .C1(n19594), .C2(n19379), .A(n19366), .B(n19365), .ZN(
        P2_U3115) );
  AOI22_X1 U22352 ( .A1(n19505), .A2(n19371), .B1(n19595), .B2(n19374), .ZN(
        n19368) );
  AOI22_X1 U22353 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19376), .B1(
        n19375), .B2(n19596), .ZN(n19367) );
  OAI211_X1 U22354 ( .C1(n19508), .C2(n19401), .A(n19368), .B(n19367), .ZN(
        P2_U3116) );
  AOI22_X1 U22355 ( .A1(n19404), .A2(n19603), .B1(n19601), .B2(n19374), .ZN(
        n19370) );
  AOI22_X1 U22356 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19376), .B1(
        n19375), .B2(n19602), .ZN(n19369) );
  OAI211_X1 U22357 ( .C1(n19606), .C2(n19379), .A(n19370), .B(n19369), .ZN(
        P2_U3117) );
  AOI22_X1 U22358 ( .A1(n19550), .A2(n19371), .B1(n19607), .B2(n19374), .ZN(
        n19373) );
  AOI22_X1 U22359 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19376), .B1(
        n19375), .B2(n19608), .ZN(n19372) );
  OAI211_X1 U22360 ( .C1(n19553), .C2(n19401), .A(n19373), .B(n19372), .ZN(
        P2_U3118) );
  AOI22_X1 U22361 ( .A1(n19404), .A2(n19617), .B1(n19613), .B2(n19374), .ZN(
        n19378) );
  AOI22_X1 U22362 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19376), .B1(
        n19375), .B2(n19615), .ZN(n19377) );
  OAI211_X1 U22363 ( .C1(n19623), .C2(n19379), .A(n19378), .B(n19377), .ZN(
        P2_U3119) );
  NOR3_X2 U22364 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20827), .A3(
        n19443), .ZN(n19412) );
  AOI22_X1 U22365 ( .A1(n19575), .A2(n19428), .B1(n19566), .B2(n19412), .ZN(
        n19390) );
  NAND2_X1 U22366 ( .A1(n19711), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19569) );
  OAI21_X1 U22367 ( .B1(n19569), .B2(n19380), .A(n19520), .ZN(n19388) );
  NOR2_X1 U22368 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19443), .ZN(
        n19384) );
  INV_X1 U22369 ( .A(n10727), .ZN(n19385) );
  OAI21_X1 U22370 ( .B1(n19385), .B2(n19350), .A(n19737), .ZN(n19382) );
  INV_X1 U22371 ( .A(n19412), .ZN(n19381) );
  AOI21_X1 U22372 ( .B1(n19382), .B2(n19381), .A(n19523), .ZN(n19383) );
  OAI21_X1 U22373 ( .B1(n19388), .B2(n19384), .A(n19383), .ZN(n19406) );
  INV_X1 U22374 ( .A(n19384), .ZN(n19387) );
  OAI21_X1 U22375 ( .B1(n19385), .B2(n19412), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19386) );
  OAI21_X1 U22376 ( .B1(n19388), .B2(n19387), .A(n19386), .ZN(n19405) );
  AOI22_X1 U22377 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19406), .B1(
        n19087), .B2(n19405), .ZN(n19389) );
  OAI211_X1 U22378 ( .C1(n19578), .C2(n19401), .A(n19390), .B(n19389), .ZN(
        P2_U3120) );
  AOI22_X1 U22379 ( .A1(n19532), .A2(n19404), .B1(n19579), .B2(n19412), .ZN(
        n19392) );
  AOI22_X1 U22380 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19406), .B1(
        n19099), .B2(n19405), .ZN(n19391) );
  OAI211_X1 U22381 ( .C1(n19535), .C2(n19437), .A(n19392), .B(n19391), .ZN(
        P2_U3121) );
  AOI22_X1 U22382 ( .A1(n19499), .A2(n19404), .B1(n19584), .B2(n19412), .ZN(
        n19394) );
  AOI22_X1 U22383 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19406), .B1(
        n19585), .B2(n19405), .ZN(n19393) );
  OAI211_X1 U22384 ( .C1(n19502), .C2(n19437), .A(n19394), .B(n19393), .ZN(
        P2_U3122) );
  AOI22_X1 U22385 ( .A1(n19428), .A2(n19591), .B1(n19590), .B2(n19412), .ZN(
        n19396) );
  AOI22_X1 U22386 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19406), .B1(
        n19111), .B2(n19405), .ZN(n19395) );
  OAI211_X1 U22387 ( .C1(n19594), .C2(n19401), .A(n19396), .B(n19395), .ZN(
        P2_U3123) );
  AOI22_X1 U22388 ( .A1(n19597), .A2(n19428), .B1(n19595), .B2(n19412), .ZN(
        n19398) );
  AOI22_X1 U22389 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19406), .B1(
        n19596), .B2(n19405), .ZN(n19397) );
  OAI211_X1 U22390 ( .C1(n19600), .C2(n19401), .A(n19398), .B(n19397), .ZN(
        P2_U3124) );
  AOI22_X1 U22391 ( .A1(n19428), .A2(n19603), .B1(n19601), .B2(n19412), .ZN(
        n19400) );
  AOI22_X1 U22392 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19406), .B1(
        n19602), .B2(n19405), .ZN(n19399) );
  OAI211_X1 U22393 ( .C1(n19606), .C2(n19401), .A(n19400), .B(n19399), .ZN(
        P2_U3125) );
  AOI22_X1 U22394 ( .A1(n19404), .A2(n19550), .B1(n19607), .B2(n19412), .ZN(
        n19403) );
  AOI22_X1 U22395 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19406), .B1(
        n19608), .B2(n19405), .ZN(n19402) );
  OAI211_X1 U22396 ( .C1(n19553), .C2(n19437), .A(n19403), .B(n19402), .ZN(
        P2_U3126) );
  AOI22_X1 U22397 ( .A1(n19556), .A2(n19404), .B1(n19613), .B2(n19412), .ZN(
        n19408) );
  AOI22_X1 U22398 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19406), .B1(
        n19615), .B2(n19405), .ZN(n19407) );
  OAI211_X1 U22399 ( .C1(n19561), .C2(n19437), .A(n19408), .B(n19407), .ZN(
        P2_U3127) );
  NOR3_X2 U22400 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19735), .A3(
        n19443), .ZN(n19431) );
  OAI21_X1 U22401 ( .B1(n19409), .B2(n19431), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19410) );
  OAI21_X1 U22402 ( .B1(n19443), .B2(n19411), .A(n19410), .ZN(n19432) );
  AOI22_X1 U22403 ( .A1(n19432), .A2(n19087), .B1(n19566), .B2(n19431), .ZN(
        n19417) );
  AOI221_X1 U22404 ( .B1(n19433), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19428), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19412), .ZN(n19413) );
  AOI211_X1 U22405 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19414), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19413), .ZN(n19415) );
  OAI21_X1 U22406 ( .B1(n19415), .B2(n19431), .A(n19573), .ZN(n19434) );
  AOI22_X1 U22407 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19434), .B1(
        n19433), .B2(n19575), .ZN(n19416) );
  OAI211_X1 U22408 ( .C1(n19578), .C2(n19437), .A(n19417), .B(n19416), .ZN(
        P2_U3128) );
  AOI22_X1 U22409 ( .A1(n19432), .A2(n19099), .B1(n19579), .B2(n19431), .ZN(
        n19419) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19434), .B1(
        n19433), .B2(n19580), .ZN(n19418) );
  OAI211_X1 U22411 ( .C1(n19583), .C2(n19437), .A(n19419), .B(n19418), .ZN(
        P2_U3129) );
  AOI22_X1 U22412 ( .A1(n19432), .A2(n19585), .B1(n19584), .B2(n19431), .ZN(
        n19421) );
  AOI22_X1 U22413 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19434), .B1(
        n19433), .B2(n19586), .ZN(n19420) );
  OAI211_X1 U22414 ( .C1(n19589), .C2(n19437), .A(n19421), .B(n19420), .ZN(
        P2_U3130) );
  AOI22_X1 U22415 ( .A1(n19432), .A2(n19111), .B1(n19590), .B2(n19431), .ZN(
        n19423) );
  AOI22_X1 U22416 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19434), .B1(
        n19433), .B2(n19591), .ZN(n19422) );
  OAI211_X1 U22417 ( .C1(n19594), .C2(n19437), .A(n19423), .B(n19422), .ZN(
        P2_U3131) );
  AOI22_X1 U22418 ( .A1(n19432), .A2(n19596), .B1(n19595), .B2(n19431), .ZN(
        n19425) );
  AOI22_X1 U22419 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19434), .B1(
        n19428), .B2(n19505), .ZN(n19424) );
  OAI211_X1 U22420 ( .C1(n19508), .C2(n19465), .A(n19425), .B(n19424), .ZN(
        P2_U3132) );
  AOI22_X1 U22421 ( .A1(n19432), .A2(n19602), .B1(n19601), .B2(n19431), .ZN(
        n19427) );
  AOI22_X1 U22422 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19434), .B1(
        n19433), .B2(n19603), .ZN(n19426) );
  OAI211_X1 U22423 ( .C1(n19606), .C2(n19437), .A(n19427), .B(n19426), .ZN(
        P2_U3133) );
  AOI22_X1 U22424 ( .A1(n19432), .A2(n19608), .B1(n19607), .B2(n19431), .ZN(
        n19430) );
  AOI22_X1 U22425 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19434), .B1(
        n19428), .B2(n19550), .ZN(n19429) );
  OAI211_X1 U22426 ( .C1(n19553), .C2(n19465), .A(n19430), .B(n19429), .ZN(
        P2_U3134) );
  AOI22_X1 U22427 ( .A1(n19432), .A2(n19615), .B1(n19613), .B2(n19431), .ZN(
        n19436) );
  AOI22_X1 U22428 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19434), .B1(
        n19433), .B2(n19617), .ZN(n19435) );
  OAI211_X1 U22429 ( .C1(n19623), .C2(n19437), .A(n19436), .B(n19435), .ZN(
        P2_U3135) );
  OR2_X1 U22430 ( .A1(n19735), .A2(n19443), .ZN(n19441) );
  INV_X1 U22431 ( .A(n19442), .ZN(n19439) );
  NOR2_X1 U22432 ( .A1(n19438), .A2(n19443), .ZN(n19460) );
  OAI21_X1 U22433 ( .B1(n19439), .B2(n19460), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19440) );
  OAI21_X1 U22434 ( .B1(n19441), .B2(n19714), .A(n19440), .ZN(n19461) );
  AOI22_X1 U22435 ( .A1(n19461), .A2(n19087), .B1(n19566), .B2(n19460), .ZN(
        n19447) );
  AOI21_X1 U22436 ( .B1(n19442), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19445) );
  OAI22_X1 U22437 ( .A1(n19569), .A2(n19707), .B1(n19735), .B2(n19443), .ZN(
        n19444) );
  OAI211_X1 U22438 ( .C1(n19460), .C2(n19445), .A(n19444), .B(n19573), .ZN(
        n19462) );
  AOI22_X1 U22439 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19462), .B1(
        n19481), .B2(n19575), .ZN(n19446) );
  OAI211_X1 U22440 ( .C1(n19578), .C2(n19465), .A(n19447), .B(n19446), .ZN(
        P2_U3136) );
  AOI22_X1 U22441 ( .A1(n19461), .A2(n19099), .B1(n19579), .B2(n19460), .ZN(
        n19449) );
  AOI22_X1 U22442 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19462), .B1(
        n19481), .B2(n19580), .ZN(n19448) );
  OAI211_X1 U22443 ( .C1(n19583), .C2(n19465), .A(n19449), .B(n19448), .ZN(
        P2_U3137) );
  AOI22_X1 U22444 ( .A1(n19461), .A2(n19585), .B1(n19584), .B2(n19460), .ZN(
        n19451) );
  AOI22_X1 U22445 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19462), .B1(
        n19481), .B2(n19586), .ZN(n19450) );
  OAI211_X1 U22446 ( .C1(n19589), .C2(n19465), .A(n19451), .B(n19450), .ZN(
        P2_U3138) );
  AOI22_X1 U22447 ( .A1(n19461), .A2(n19111), .B1(n19590), .B2(n19460), .ZN(
        n19453) );
  AOI22_X1 U22448 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19462), .B1(
        n19481), .B2(n19591), .ZN(n19452) );
  OAI211_X1 U22449 ( .C1(n19594), .C2(n19465), .A(n19453), .B(n19452), .ZN(
        P2_U3139) );
  AOI22_X1 U22450 ( .A1(n19461), .A2(n19596), .B1(n19595), .B2(n19460), .ZN(
        n19455) );
  AOI22_X1 U22451 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19462), .B1(
        n19481), .B2(n19597), .ZN(n19454) );
  OAI211_X1 U22452 ( .C1(n19600), .C2(n19465), .A(n19455), .B(n19454), .ZN(
        P2_U3140) );
  AOI22_X1 U22453 ( .A1(n19461), .A2(n19602), .B1(n19601), .B2(n19460), .ZN(
        n19457) );
  AOI22_X1 U22454 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19462), .B1(
        n19481), .B2(n19603), .ZN(n19456) );
  OAI211_X1 U22455 ( .C1(n19606), .C2(n19465), .A(n19457), .B(n19456), .ZN(
        P2_U3141) );
  AOI22_X1 U22456 ( .A1(n19461), .A2(n19608), .B1(n19607), .B2(n19460), .ZN(
        n19459) );
  AOI22_X1 U22457 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19462), .B1(
        n19481), .B2(n19609), .ZN(n19458) );
  OAI211_X1 U22458 ( .C1(n19612), .C2(n19465), .A(n19459), .B(n19458), .ZN(
        P2_U3142) );
  AOI22_X1 U22459 ( .A1(n19461), .A2(n19615), .B1(n19613), .B2(n19460), .ZN(
        n19464) );
  AOI22_X1 U22460 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19462), .B1(
        n19481), .B2(n19617), .ZN(n19463) );
  OAI211_X1 U22461 ( .C1(n19623), .C2(n19465), .A(n19464), .B(n19463), .ZN(
        P2_U3143) );
  AOI22_X1 U22462 ( .A1(n19480), .A2(n19087), .B1(n19479), .B2(n19566), .ZN(
        n19468) );
  AOI22_X1 U22463 ( .A1(n19515), .A2(n19575), .B1(n19481), .B2(n19466), .ZN(
        n19467) );
  OAI211_X1 U22464 ( .C1(n19484), .C2(n12440), .A(n19468), .B(n19467), .ZN(
        P2_U3144) );
  AOI22_X1 U22465 ( .A1(n19480), .A2(n19099), .B1(n19479), .B2(n19579), .ZN(
        n19470) );
  AOI22_X1 U22466 ( .A1(n19515), .A2(n19580), .B1(n19481), .B2(n19532), .ZN(
        n19469) );
  OAI211_X1 U22467 ( .C1(n19484), .C2(n19471), .A(n19470), .B(n19469), .ZN(
        P2_U3145) );
  AOI22_X1 U22468 ( .A1(n19480), .A2(n19585), .B1(n19479), .B2(n19584), .ZN(
        n19473) );
  AOI22_X1 U22469 ( .A1(n19515), .A2(n19586), .B1(n19481), .B2(n19499), .ZN(
        n19472) );
  OAI211_X1 U22470 ( .C1(n19484), .C2(n12509), .A(n19473), .B(n19472), .ZN(
        P2_U3146) );
  INV_X1 U22471 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n19476) );
  AOI22_X1 U22472 ( .A1(n19480), .A2(n19111), .B1(n19479), .B2(n19590), .ZN(
        n19475) );
  AOI22_X1 U22473 ( .A1(n19515), .A2(n19591), .B1(n19481), .B2(n19538), .ZN(
        n19474) );
  OAI211_X1 U22474 ( .C1(n19484), .C2(n19476), .A(n19475), .B(n19474), .ZN(
        P2_U3147) );
  AOI22_X1 U22475 ( .A1(n19480), .A2(n19596), .B1(n19479), .B2(n19595), .ZN(
        n19478) );
  AOI22_X1 U22476 ( .A1(n19481), .A2(n19505), .B1(n19515), .B2(n19597), .ZN(
        n19477) );
  OAI211_X1 U22477 ( .C1(n19484), .C2(n12556), .A(n19478), .B(n19477), .ZN(
        P2_U3148) );
  AOI22_X1 U22478 ( .A1(n19480), .A2(n19608), .B1(n19479), .B2(n19607), .ZN(
        n19483) );
  AOI22_X1 U22479 ( .A1(n19481), .A2(n19550), .B1(n19515), .B2(n19609), .ZN(
        n19482) );
  OAI211_X1 U22480 ( .C1(n19484), .C2(n12419), .A(n19483), .B(n19482), .ZN(
        P2_U3150) );
  NOR2_X1 U22481 ( .A1(n20827), .A2(n19489), .ZN(n19525) );
  INV_X1 U22482 ( .A(n19525), .ZN(n19485) );
  AND2_X1 U22483 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19485), .ZN(n19486) );
  NAND2_X1 U22484 ( .A1(n19487), .A2(n19486), .ZN(n19490) );
  OAI21_X1 U22485 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19489), .A(n19350), 
        .ZN(n19488) );
  AND2_X1 U22486 ( .A1(n19490), .A2(n19488), .ZN(n19514) );
  AOI22_X1 U22487 ( .A1(n19514), .A2(n19087), .B1(n19566), .B2(n19525), .ZN(
        n19496) );
  OAI21_X1 U22488 ( .B1(n19569), .B2(n19493), .A(n19489), .ZN(n19491) );
  AND2_X1 U22489 ( .A1(n19491), .A2(n19490), .ZN(n19492) );
  OAI211_X1 U22490 ( .C1(n19525), .C2(n19737), .A(n19492), .B(n19573), .ZN(
        n19516) );
  AOI22_X1 U22491 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19516), .B1(
        n19555), .B2(n19575), .ZN(n19495) );
  OAI211_X1 U22492 ( .C1(n19578), .C2(n19513), .A(n19496), .B(n19495), .ZN(
        P2_U3152) );
  AOI22_X1 U22493 ( .A1(n19514), .A2(n19099), .B1(n19579), .B2(n19525), .ZN(
        n19498) );
  AOI22_X1 U22494 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19516), .B1(
        n19555), .B2(n19580), .ZN(n19497) );
  OAI211_X1 U22495 ( .C1(n19583), .C2(n19513), .A(n19498), .B(n19497), .ZN(
        P2_U3153) );
  AOI22_X1 U22496 ( .A1(n19514), .A2(n19585), .B1(n19584), .B2(n19525), .ZN(
        n19501) );
  AOI22_X1 U22497 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19516), .B1(
        n19515), .B2(n19499), .ZN(n19500) );
  OAI211_X1 U22498 ( .C1(n19502), .C2(n19545), .A(n19501), .B(n19500), .ZN(
        P2_U3154) );
  AOI22_X1 U22499 ( .A1(n19514), .A2(n19111), .B1(n19590), .B2(n19525), .ZN(
        n19504) );
  AOI22_X1 U22500 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19516), .B1(
        n19555), .B2(n19591), .ZN(n19503) );
  OAI211_X1 U22501 ( .C1(n19594), .C2(n19513), .A(n19504), .B(n19503), .ZN(
        P2_U3155) );
  AOI22_X1 U22502 ( .A1(n19514), .A2(n19596), .B1(n19595), .B2(n19525), .ZN(
        n19507) );
  AOI22_X1 U22503 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19516), .B1(
        n19515), .B2(n19505), .ZN(n19506) );
  OAI211_X1 U22504 ( .C1(n19508), .C2(n19545), .A(n19507), .B(n19506), .ZN(
        P2_U3156) );
  AOI22_X1 U22505 ( .A1(n19514), .A2(n19602), .B1(n19601), .B2(n19525), .ZN(
        n19510) );
  AOI22_X1 U22506 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19516), .B1(
        n19555), .B2(n19603), .ZN(n19509) );
  OAI211_X1 U22507 ( .C1(n19606), .C2(n19513), .A(n19510), .B(n19509), .ZN(
        P2_U3157) );
  AOI22_X1 U22508 ( .A1(n19514), .A2(n19608), .B1(n19607), .B2(n19525), .ZN(
        n19512) );
  AOI22_X1 U22509 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19516), .B1(
        n19555), .B2(n19609), .ZN(n19511) );
  OAI211_X1 U22510 ( .C1(n19612), .C2(n19513), .A(n19512), .B(n19511), .ZN(
        P2_U3158) );
  AOI22_X1 U22511 ( .A1(n19514), .A2(n19615), .B1(n19613), .B2(n19525), .ZN(
        n19518) );
  AOI22_X1 U22512 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19516), .B1(
        n19515), .B2(n19556), .ZN(n19517) );
  OAI211_X1 U22513 ( .C1(n19561), .C2(n19545), .A(n19518), .B(n19517), .ZN(
        P2_U3159) );
  INV_X1 U22514 ( .A(n19622), .ZN(n19542) );
  NOR3_X2 U22515 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19718), .A3(
        n19567), .ZN(n19554) );
  AOI22_X1 U22516 ( .A1(n19575), .A2(n19542), .B1(n19566), .B2(n19554), .ZN(
        n19531) );
  NOR3_X1 U22517 ( .A1(n19526), .A2(n19554), .A3(n19350), .ZN(n19524) );
  OAI21_X1 U22518 ( .B1(n19555), .B2(n19542), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19521) );
  NAND2_X1 U22519 ( .A1(n19521), .A2(n19520), .ZN(n19529) );
  AOI221_X1 U22520 ( .B1(n19737), .B2(n19529), .C1(n19737), .C2(n19525), .A(
        n19554), .ZN(n19522) );
  NOR2_X1 U22521 ( .A1(n19554), .A2(n19525), .ZN(n19528) );
  OAI21_X1 U22522 ( .B1(n19526), .B2(n19554), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19527) );
  AOI22_X1 U22523 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19558), .B1(
        n19087), .B2(n19557), .ZN(n19530) );
  OAI211_X1 U22524 ( .C1(n19578), .C2(n19545), .A(n19531), .B(n19530), .ZN(
        P2_U3160) );
  AOI22_X1 U22525 ( .A1(n19532), .A2(n19555), .B1(n19579), .B2(n19554), .ZN(
        n19534) );
  AOI22_X1 U22526 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19558), .B1(
        n19099), .B2(n19557), .ZN(n19533) );
  OAI211_X1 U22527 ( .C1(n19535), .C2(n19622), .A(n19534), .B(n19533), .ZN(
        P2_U3161) );
  AOI22_X1 U22528 ( .A1(n19542), .A2(n19586), .B1(n19584), .B2(n19554), .ZN(
        n19537) );
  AOI22_X1 U22529 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19558), .B1(
        n19585), .B2(n19557), .ZN(n19536) );
  OAI211_X1 U22530 ( .C1(n19589), .C2(n19545), .A(n19537), .B(n19536), .ZN(
        P2_U3162) );
  AOI22_X1 U22531 ( .A1(n19538), .A2(n19555), .B1(n19590), .B2(n19554), .ZN(
        n19540) );
  AOI22_X1 U22532 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19558), .B1(
        n19111), .B2(n19557), .ZN(n19539) );
  OAI211_X1 U22533 ( .C1(n19541), .C2(n19622), .A(n19540), .B(n19539), .ZN(
        P2_U3163) );
  AOI22_X1 U22534 ( .A1(n19597), .A2(n19542), .B1(n19595), .B2(n19554), .ZN(
        n19544) );
  AOI22_X1 U22535 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19558), .B1(
        n19596), .B2(n19557), .ZN(n19543) );
  OAI211_X1 U22536 ( .C1(n19600), .C2(n19545), .A(n19544), .B(n19543), .ZN(
        P2_U3164) );
  AOI22_X1 U22537 ( .A1(n19546), .A2(n19555), .B1(n19601), .B2(n19554), .ZN(
        n19548) );
  AOI22_X1 U22538 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19558), .B1(
        n19602), .B2(n19557), .ZN(n19547) );
  OAI211_X1 U22539 ( .C1(n19549), .C2(n19622), .A(n19548), .B(n19547), .ZN(
        P2_U3165) );
  AOI22_X1 U22540 ( .A1(n19555), .A2(n19550), .B1(n19607), .B2(n19554), .ZN(
        n19552) );
  AOI22_X1 U22541 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19558), .B1(
        n19608), .B2(n19557), .ZN(n19551) );
  OAI211_X1 U22542 ( .C1(n19553), .C2(n19622), .A(n19552), .B(n19551), .ZN(
        P2_U3166) );
  AOI22_X1 U22543 ( .A1(n19556), .A2(n19555), .B1(n19613), .B2(n19554), .ZN(
        n19560) );
  AOI22_X1 U22544 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19558), .B1(
        n19615), .B2(n19557), .ZN(n19559) );
  OAI211_X1 U22545 ( .C1(n19561), .C2(n19622), .A(n19560), .B(n19559), .ZN(
        P2_U3167) );
  NAND2_X1 U22546 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19562), .ZN(
        n19565) );
  INV_X1 U22547 ( .A(n19571), .ZN(n19563) );
  INV_X1 U22548 ( .A(n19570), .ZN(n19614) );
  OAI21_X1 U22549 ( .B1(n19563), .B2(n19614), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19564) );
  OAI21_X1 U22550 ( .B1(n19565), .B2(n19714), .A(n19564), .ZN(n19616) );
  AOI22_X1 U22551 ( .A1(n19616), .A2(n19087), .B1(n19614), .B2(n19566), .ZN(
        n19577) );
  OAI22_X1 U22552 ( .A1(n19569), .A2(n19568), .B1(n19567), .B2(n19718), .ZN(
        n19574) );
  OAI211_X1 U22553 ( .C1(n19571), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19570), 
        .B(n19714), .ZN(n19572) );
  NAND3_X1 U22554 ( .A1(n19574), .A2(n19573), .A3(n19572), .ZN(n19619) );
  AOI22_X1 U22555 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19619), .B1(
        n19618), .B2(n19575), .ZN(n19576) );
  OAI211_X1 U22556 ( .C1(n19578), .C2(n19622), .A(n19577), .B(n19576), .ZN(
        P2_U3168) );
  AOI22_X1 U22557 ( .A1(n19616), .A2(n19099), .B1(n19614), .B2(n19579), .ZN(
        n19582) );
  AOI22_X1 U22558 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19619), .B1(
        n19618), .B2(n19580), .ZN(n19581) );
  OAI211_X1 U22559 ( .C1(n19583), .C2(n19622), .A(n19582), .B(n19581), .ZN(
        P2_U3169) );
  AOI22_X1 U22560 ( .A1(n19616), .A2(n19585), .B1(n19614), .B2(n19584), .ZN(
        n19588) );
  AOI22_X1 U22561 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19619), .B1(
        n19618), .B2(n19586), .ZN(n19587) );
  OAI211_X1 U22562 ( .C1(n19589), .C2(n19622), .A(n19588), .B(n19587), .ZN(
        P2_U3170) );
  AOI22_X1 U22563 ( .A1(n19616), .A2(n19111), .B1(n19614), .B2(n19590), .ZN(
        n19593) );
  AOI22_X1 U22564 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19619), .B1(
        n19618), .B2(n19591), .ZN(n19592) );
  OAI211_X1 U22565 ( .C1(n19594), .C2(n19622), .A(n19593), .B(n19592), .ZN(
        P2_U3171) );
  AOI22_X1 U22566 ( .A1(n19616), .A2(n19596), .B1(n19614), .B2(n19595), .ZN(
        n19599) );
  AOI22_X1 U22567 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19619), .B1(
        n19618), .B2(n19597), .ZN(n19598) );
  OAI211_X1 U22568 ( .C1(n19600), .C2(n19622), .A(n19599), .B(n19598), .ZN(
        P2_U3172) );
  AOI22_X1 U22569 ( .A1(n19616), .A2(n19602), .B1(n19614), .B2(n19601), .ZN(
        n19605) );
  AOI22_X1 U22570 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19619), .B1(
        n19618), .B2(n19603), .ZN(n19604) );
  OAI211_X1 U22571 ( .C1(n19606), .C2(n19622), .A(n19605), .B(n19604), .ZN(
        P2_U3173) );
  AOI22_X1 U22572 ( .A1(n19616), .A2(n19608), .B1(n19614), .B2(n19607), .ZN(
        n19611) );
  AOI22_X1 U22573 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19619), .B1(
        n19618), .B2(n19609), .ZN(n19610) );
  OAI211_X1 U22574 ( .C1(n19612), .C2(n19622), .A(n19611), .B(n19610), .ZN(
        P2_U3174) );
  AOI22_X1 U22575 ( .A1(n19616), .A2(n19615), .B1(n19614), .B2(n19613), .ZN(
        n19621) );
  AOI22_X1 U22576 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19619), .B1(
        n19618), .B2(n19617), .ZN(n19620) );
  OAI211_X1 U22577 ( .C1(n19623), .C2(n19622), .A(n19621), .B(n19620), .ZN(
        P2_U3175) );
  OAI211_X1 U22578 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19756), .A(n19625), 
        .B(n19624), .ZN(n19630) );
  NOR2_X1 U22579 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19762), .ZN(n19626) );
  OAI211_X1 U22580 ( .C1(n19627), .C2(n19626), .A(n19768), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19629) );
  OAI211_X1 U22581 ( .C1(n19631), .C2(n19630), .A(n19629), .B(n19628), .ZN(
        P2_U3177) );
  AND2_X1 U22582 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19632), .ZN(
        P2_U3179) );
  AND2_X1 U22583 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19632), .ZN(
        P2_U3180) );
  AND2_X1 U22584 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19632), .ZN(
        P2_U3181) );
  AND2_X1 U22585 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19632), .ZN(
        P2_U3182) );
  INV_X1 U22586 ( .A(P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20744) );
  NOR2_X1 U22587 ( .A1(n20744), .A2(n19705), .ZN(P2_U3183) );
  AND2_X1 U22588 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19632), .ZN(
        P2_U3184) );
  AND2_X1 U22589 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19632), .ZN(
        P2_U3185) );
  AND2_X1 U22590 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19632), .ZN(
        P2_U3186) );
  AND2_X1 U22591 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19632), .ZN(
        P2_U3187) );
  AND2_X1 U22592 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19632), .ZN(
        P2_U3188) );
  AND2_X1 U22593 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19632), .ZN(
        P2_U3189) );
  AND2_X1 U22594 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19632), .ZN(
        P2_U3190) );
  AND2_X1 U22595 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19632), .ZN(
        P2_U3191) );
  AND2_X1 U22596 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19632), .ZN(
        P2_U3192) );
  AND2_X1 U22597 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19632), .ZN(
        P2_U3193) );
  INV_X1 U22598 ( .A(P2_DATAWIDTH_REG_16__SCAN_IN), .ZN(n20775) );
  NOR2_X1 U22599 ( .A1(n20775), .A2(n19705), .ZN(P2_U3194) );
  AND2_X1 U22600 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19632), .ZN(
        P2_U3195) );
  AND2_X1 U22601 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19632), .ZN(
        P2_U3196) );
  NOR2_X1 U22602 ( .A1(n20686), .A2(n19705), .ZN(P2_U3197) );
  INV_X1 U22603 ( .A(P2_DATAWIDTH_REG_12__SCAN_IN), .ZN(n20726) );
  NOR2_X1 U22604 ( .A1(n20726), .A2(n19705), .ZN(P2_U3198) );
  AND2_X1 U22605 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19632), .ZN(
        P2_U3199) );
  AND2_X1 U22606 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19632), .ZN(
        P2_U3200) );
  AND2_X1 U22607 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19632), .ZN(P2_U3201) );
  AND2_X1 U22608 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19632), .ZN(P2_U3202) );
  AND2_X1 U22609 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19632), .ZN(P2_U3203) );
  AND2_X1 U22610 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19632), .ZN(P2_U3204) );
  AND2_X1 U22611 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19632), .ZN(P2_U3205) );
  AND2_X1 U22612 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19632), .ZN(P2_U3206) );
  NOR2_X1 U22613 ( .A1(n20728), .A2(n19705), .ZN(P2_U3207) );
  AND2_X1 U22614 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19632), .ZN(P2_U3208) );
  INV_X1 U22615 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19774) );
  INV_X1 U22616 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19642) );
  NOR2_X1 U22617 ( .A1(n19642), .A2(n19756), .ZN(n19640) );
  OR3_X1 U22618 ( .A1(n19774), .A2(n19633), .A3(n19640), .ZN(n19634) );
  NOR3_X1 U22619 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n20566), .ZN(n19646) );
  AOI21_X1 U22620 ( .B1(n19649), .B2(n19634), .A(n19646), .ZN(n19635) );
  OAI221_X1 U22621 ( .B1(n19636), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .C1(
        n19636), .C2(n20561), .A(n19635), .ZN(P2_U3209) );
  AOI21_X1 U22622 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20561), .A(n19649), 
        .ZN(n19643) );
  NOR3_X1 U22623 ( .A1(n19643), .A2(n19774), .A3(n19633), .ZN(n19637) );
  NOR2_X1 U22624 ( .A1(n19637), .A2(n19640), .ZN(n19638) );
  OAI211_X1 U22625 ( .C1(n20561), .C2(n19639), .A(n19638), .B(n19766), .ZN(
        P2_U3210) );
  AOI22_X1 U22626 ( .A1(n19641), .A2(n19774), .B1(n19640), .B2(n20566), .ZN(
        n19648) );
  OAI21_X1 U22627 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n19647) );
  NOR2_X1 U22628 ( .A1(n19642), .A2(n19649), .ZN(n19644) );
  AOI21_X1 U22629 ( .B1(n19768), .B2(n19644), .A(n19643), .ZN(n19645) );
  OAI22_X1 U22630 ( .A1(n19648), .A2(n19647), .B1(n19646), .B2(n19645), .ZN(
        P2_U3211) );
  NAND2_X2 U22631 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19776), .ZN(n19695) );
  NAND2_X2 U22632 ( .A1(n19776), .A2(n19649), .ZN(n19698) );
  OAI222_X1 U22633 ( .A1(n19695), .A2(n20772), .B1(n19650), .B2(n19776), .C1(
        n19652), .C2(n19698), .ZN(P2_U3212) );
  OAI222_X1 U22634 ( .A1(n19695), .A2(n19652), .B1(n19651), .B2(n19776), .C1(
        n12713), .C2(n19698), .ZN(P2_U3213) );
  OAI222_X1 U22635 ( .A1(n19695), .A2(n12713), .B1(n19653), .B2(n19776), .C1(
        n12720), .C2(n19698), .ZN(P2_U3214) );
  OAI222_X1 U22636 ( .A1(n19698), .A2(n19655), .B1(n19654), .B2(n19776), .C1(
        n12720), .C2(n19695), .ZN(P2_U3215) );
  OAI222_X1 U22637 ( .A1(n19698), .A2(n19657), .B1(n19656), .B2(n19776), .C1(
        n19655), .C2(n19695), .ZN(P2_U3216) );
  OAI222_X1 U22638 ( .A1(n19698), .A2(n19659), .B1(n19658), .B2(n19776), .C1(
        n19657), .C2(n19695), .ZN(P2_U3217) );
  OAI222_X1 U22639 ( .A1(n19698), .A2(n12736), .B1(n19660), .B2(n19776), .C1(
        n19659), .C2(n19695), .ZN(P2_U3218) );
  OAI222_X1 U22640 ( .A1(n19698), .A2(n12742), .B1(n19661), .B2(n19776), .C1(
        n12736), .C2(n19695), .ZN(P2_U3219) );
  OAI222_X1 U22641 ( .A1(n19698), .A2(n13995), .B1(n19662), .B2(n19776), .C1(
        n12742), .C2(n19695), .ZN(P2_U3220) );
  OAI222_X1 U22642 ( .A1(n19698), .A2(n12748), .B1(n19663), .B2(n19776), .C1(
        n13995), .C2(n19695), .ZN(P2_U3221) );
  OAI222_X1 U22643 ( .A1(n19698), .A2(n12749), .B1(n20824), .B2(n19776), .C1(
        n12748), .C2(n19695), .ZN(P2_U3222) );
  OAI222_X1 U22644 ( .A1(n19698), .A2(n12756), .B1(n19664), .B2(n19776), .C1(
        n12749), .C2(n19695), .ZN(P2_U3223) );
  OAI222_X1 U22645 ( .A1(n19698), .A2(n19666), .B1(n19665), .B2(n19776), .C1(
        n12756), .C2(n19695), .ZN(P2_U3224) );
  OAI222_X1 U22646 ( .A1(n19698), .A2(n19667), .B1(n20755), .B2(n19776), .C1(
        n19666), .C2(n19695), .ZN(P2_U3225) );
  OAI222_X1 U22647 ( .A1(n19698), .A2(n19669), .B1(n19668), .B2(n19776), .C1(
        n19667), .C2(n19695), .ZN(P2_U3226) );
  OAI222_X1 U22648 ( .A1(n19698), .A2(n19671), .B1(n19670), .B2(n19776), .C1(
        n19669), .C2(n19695), .ZN(P2_U3227) );
  OAI222_X1 U22649 ( .A1(n19698), .A2(n19673), .B1(n19672), .B2(n19776), .C1(
        n19671), .C2(n19695), .ZN(P2_U3228) );
  OAI222_X1 U22650 ( .A1(n19698), .A2(n19675), .B1(n19674), .B2(n19776), .C1(
        n19673), .C2(n19695), .ZN(P2_U3229) );
  OAI222_X1 U22651 ( .A1(n19698), .A2(n19677), .B1(n19676), .B2(n19776), .C1(
        n19675), .C2(n19695), .ZN(P2_U3230) );
  OAI222_X1 U22652 ( .A1(n19698), .A2(n20763), .B1(n19678), .B2(n19776), .C1(
        n19677), .C2(n19695), .ZN(P2_U3231) );
  INV_X1 U22653 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19680) );
  OAI222_X1 U22654 ( .A1(n19698), .A2(n19680), .B1(n19679), .B2(n19776), .C1(
        n20763), .C2(n19695), .ZN(P2_U3232) );
  OAI222_X1 U22655 ( .A1(n19698), .A2(n19682), .B1(n19681), .B2(n19776), .C1(
        n19680), .C2(n19695), .ZN(P2_U3233) );
  OAI222_X1 U22656 ( .A1(n19698), .A2(n19684), .B1(n19683), .B2(n19776), .C1(
        n19682), .C2(n19695), .ZN(P2_U3234) );
  OAI222_X1 U22657 ( .A1(n19698), .A2(n19686), .B1(n19685), .B2(n19776), .C1(
        n19684), .C2(n19695), .ZN(P2_U3235) );
  INV_X1 U22658 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19688) );
  OAI222_X1 U22659 ( .A1(n19698), .A2(n19688), .B1(n19687), .B2(n19776), .C1(
        n19686), .C2(n19695), .ZN(P2_U3236) );
  OAI222_X1 U22660 ( .A1(n19698), .A2(n19690), .B1(n20769), .B2(n19776), .C1(
        n19688), .C2(n19695), .ZN(P2_U3237) );
  OAI222_X1 U22661 ( .A1(n19695), .A2(n19690), .B1(n19689), .B2(n19776), .C1(
        n19691), .C2(n19698), .ZN(P2_U3238) );
  OAI222_X1 U22662 ( .A1(n19698), .A2(n19693), .B1(n19692), .B2(n19776), .C1(
        n19691), .C2(n19695), .ZN(P2_U3239) );
  INV_X1 U22663 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19696) );
  OAI222_X1 U22664 ( .A1(n19698), .A2(n19696), .B1(n19694), .B2(n19776), .C1(
        n19693), .C2(n19695), .ZN(P2_U3240) );
  INV_X1 U22665 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19697) );
  OAI222_X1 U22666 ( .A1(n19698), .A2(n19697), .B1(n20825), .B2(n19776), .C1(
        n19696), .C2(n19695), .ZN(P2_U3241) );
  OAI22_X1 U22667 ( .A1(n19777), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19776), .ZN(n19699) );
  INV_X1 U22668 ( .A(n19699), .ZN(P2_U3585) );
  MUX2_X1 U22669 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n19777), .Z(P2_U3586) );
  OAI22_X1 U22670 ( .A1(n19777), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19776), .ZN(n19700) );
  INV_X1 U22671 ( .A(n19700), .ZN(P2_U3587) );
  OAI22_X1 U22672 ( .A1(n19777), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19776), .ZN(n19701) );
  INV_X1 U22673 ( .A(n19701), .ZN(P2_U3588) );
  OAI21_X1 U22674 ( .B1(n19705), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19703), 
        .ZN(n19702) );
  INV_X1 U22675 ( .A(n19702), .ZN(P2_U3591) );
  OAI21_X1 U22676 ( .B1(n19705), .B2(n19704), .A(n19703), .ZN(P2_U3592) );
  INV_X1 U22677 ( .A(n19743), .ZN(n19745) );
  INV_X1 U22678 ( .A(n19728), .ZN(n19706) );
  OR2_X1 U22679 ( .A1(n19707), .A2(n19706), .ZN(n19719) );
  NAND2_X1 U22680 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19708), .ZN(n19709) );
  OAI21_X1 U22681 ( .B1(n19732), .B2(n19709), .A(n19736), .ZN(n19720) );
  NAND2_X1 U22682 ( .A1(n19719), .A2(n19720), .ZN(n19712) );
  AOI22_X1 U22683 ( .A1(n19712), .A2(n19711), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19710), .ZN(n19713) );
  OAI21_X1 U22684 ( .B1(n19715), .B2(n19714), .A(n19713), .ZN(n19716) );
  INV_X1 U22685 ( .A(n19716), .ZN(n19717) );
  AOI22_X1 U22686 ( .A1(n19745), .A2(n19718), .B1(n19717), .B2(n19743), .ZN(
        P2_U3602) );
  OAI21_X1 U22687 ( .B1(n19721), .B2(n19720), .A(n19719), .ZN(n19722) );
  AOI21_X1 U22688 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19723), .A(n19722), 
        .ZN(n19724) );
  AOI22_X1 U22689 ( .A1(n19745), .A2(n19725), .B1(n19724), .B2(n19743), .ZN(
        P2_U3603) );
  OAI21_X1 U22690 ( .B1(n11212), .B2(n19726), .A(n19736), .ZN(n19731) );
  NAND2_X1 U22691 ( .A1(n19727), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19730) );
  NAND2_X1 U22692 ( .A1(n19732), .A2(n19728), .ZN(n19729) );
  OAI211_X1 U22693 ( .C1(n19732), .C2(n19731), .A(n19730), .B(n19729), .ZN(
        n19733) );
  INV_X1 U22694 ( .A(n19733), .ZN(n19734) );
  AOI22_X1 U22695 ( .A1(n19745), .A2(n19735), .B1(n19734), .B2(n19743), .ZN(
        P2_U3604) );
  INV_X1 U22696 ( .A(n19736), .ZN(n19738) );
  OAI22_X1 U22697 ( .A1(n19739), .A2(n19738), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19737), .ZN(n19740) );
  AOI21_X1 U22698 ( .B1(n19742), .B2(n19741), .A(n19740), .ZN(n19744) );
  AOI22_X1 U22699 ( .A1(n19745), .A2(n20827), .B1(n19744), .B2(n19743), .ZN(
        P2_U3605) );
  INV_X1 U22700 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19746) );
  AOI22_X1 U22701 ( .A1(n19776), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19746), 
        .B2(n19777), .ZN(P2_U3608) );
  AOI21_X1 U22702 ( .B1(n19748), .B2(n19747), .A(n19761), .ZN(n19749) );
  AOI21_X1 U22703 ( .B1(n10565), .B2(n19750), .A(n19749), .ZN(n19752) );
  OAI21_X1 U22704 ( .B1(n19752), .B2(n10929), .A(n19751), .ZN(n19754) );
  MUX2_X1 U22705 ( .A(P2_MORE_REG_SCAN_IN), .B(n19754), .S(n19753), .Z(
        P2_U3609) );
  AOI22_X1 U22706 ( .A1(n19757), .A2(n19756), .B1(n19737), .B2(n19755), .ZN(
        n19760) );
  INV_X1 U22707 ( .A(n19758), .ZN(n19759) );
  NAND2_X1 U22708 ( .A1(n19760), .A2(n19759), .ZN(n19775) );
  AOI211_X1 U22709 ( .C1(P2_STATEBS16_REG_SCAN_IN), .C2(n19763), .A(n19762), 
        .B(n19761), .ZN(n19772) );
  NAND3_X1 U22710 ( .A1(n19766), .A2(n19765), .A3(n19764), .ZN(n19770) );
  OAI21_X1 U22711 ( .B1(n19768), .B2(n19350), .A(n19767), .ZN(n19769) );
  NAND2_X1 U22712 ( .A1(n19770), .A2(n19769), .ZN(n19771) );
  OAI21_X1 U22713 ( .B1(n19772), .B2(n19771), .A(n19775), .ZN(n19773) );
  OAI21_X1 U22714 ( .B1(n19775), .B2(n19774), .A(n19773), .ZN(P2_U3610) );
  OAI22_X1 U22715 ( .A1(n19777), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19776), .ZN(n19778) );
  INV_X1 U22716 ( .A(n19778), .ZN(P2_U3611) );
  AOI21_X1 U22717 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20575), .A(n20564), 
        .ZN(n19785) );
  INV_X1 U22718 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19779) );
  AOI21_X1 U22719 ( .B1(n19785), .B2(n19779), .A(n20666), .ZN(P1_U2802) );
  OAI21_X1 U22720 ( .B1(n19781), .B2(n19780), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19782) );
  OAI21_X1 U22721 ( .B1(n19783), .B2(n20556), .A(n19782), .ZN(P1_U2803) );
  NOR2_X1 U22722 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19786) );
  OAI21_X1 U22723 ( .B1(n19786), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20676), .ZN(
        n19784) );
  OAI21_X1 U22724 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20664), .A(n19784), 
        .ZN(P1_U2804) );
  NOR2_X1 U22725 ( .A1(n20666), .A2(n19785), .ZN(n20632) );
  OAI21_X1 U22726 ( .B1(BS16), .B2(n19786), .A(n20632), .ZN(n20630) );
  OAI21_X1 U22727 ( .B1(n20632), .B2(n20640), .A(n20630), .ZN(P1_U2805) );
  AOI21_X1 U22728 ( .B1(n19787), .B2(P1_FLUSH_REG_SCAN_IN), .A(n19968), .ZN(
        n19788) );
  INV_X1 U22729 ( .A(n19788), .ZN(P1_U2806) );
  NOR4_X1 U22730 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19792) );
  NOR4_X1 U22731 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19791) );
  NOR4_X1 U22732 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19790) );
  NOR4_X1 U22733 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19789) );
  NAND4_X1 U22734 ( .A1(n19792), .A2(n19791), .A3(n19790), .A4(n19789), .ZN(
        n19798) );
  NOR4_X1 U22735 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19796) );
  AOI211_X1 U22736 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_5__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19795) );
  NOR4_X1 U22737 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19794) );
  NOR4_X1 U22738 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19793) );
  NAND4_X1 U22739 ( .A1(n19796), .A2(n19795), .A3(n19794), .A4(n19793), .ZN(
        n19797) );
  NOR2_X1 U22740 ( .A1(n19798), .A2(n19797), .ZN(n20663) );
  INV_X1 U22741 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19800) );
  NOR3_X1 U22742 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19801) );
  OAI21_X1 U22743 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19801), .A(n20663), .ZN(
        n19799) );
  OAI21_X1 U22744 ( .B1(n20663), .B2(n19800), .A(n19799), .ZN(P1_U2807) );
  INV_X1 U22745 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20631) );
  AOI21_X1 U22746 ( .B1(n13655), .B2(n20631), .A(n19801), .ZN(n19803) );
  INV_X1 U22747 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19802) );
  INV_X1 U22748 ( .A(n20663), .ZN(n20660) );
  AOI22_X1 U22749 ( .A1(n20663), .A2(n19803), .B1(n19802), .B2(n20660), .ZN(
        P1_U2808) );
  INV_X1 U22750 ( .A(n19806), .ZN(n19804) );
  NOR2_X1 U22751 ( .A1(n19835), .A2(n19804), .ZN(n19817) );
  NOR2_X1 U22752 ( .A1(n19817), .A2(n19805), .ZN(n19830) );
  NOR2_X1 U22753 ( .A1(n19806), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n19811) );
  AOI22_X1 U22754 ( .A1(P1_EBX_REG_9__SCAN_IN), .A2(n19875), .B1(n19884), .B2(
        n19807), .ZN(n19808) );
  OAI211_X1 U22755 ( .C1(n19867), .C2(n19809), .A(n19864), .B(n19808), .ZN(
        n19810) );
  AOI21_X1 U22756 ( .B1(n19812), .B2(n19811), .A(n19810), .ZN(n19816) );
  AOI22_X1 U22757 ( .A1(n19814), .A2(n19857), .B1(n19852), .B2(n19813), .ZN(
        n19815) );
  OAI211_X1 U22758 ( .C1(n19830), .C2(n20586), .A(n19816), .B(n19815), .ZN(
        P1_U2831) );
  INV_X1 U22759 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n19829) );
  AOI22_X1 U22760 ( .A1(n19884), .A2(n19819), .B1(n19818), .B2(n19817), .ZN(
        n19820) );
  OAI21_X1 U22761 ( .B1(n19822), .B2(n19821), .A(n19820), .ZN(n19823) );
  AOI211_X1 U22762 ( .C1(n19876), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n19879), .B(n19823), .ZN(n19828) );
  INV_X1 U22763 ( .A(n19824), .ZN(n19825) );
  AOI22_X1 U22764 ( .A1(n19826), .A2(n19857), .B1(n19825), .B2(n19852), .ZN(
        n19827) );
  OAI211_X1 U22765 ( .C1(n19830), .C2(n19829), .A(n19828), .B(n19827), .ZN(
        P1_U2832) );
  INV_X1 U22766 ( .A(n19834), .ZN(n19832) );
  OAI21_X1 U22767 ( .B1(n19835), .B2(n19832), .A(n19831), .ZN(n19880) );
  AOI21_X1 U22768 ( .B1(n19836), .B2(n19833), .A(n19880), .ZN(n19854) );
  NOR2_X1 U22769 ( .A1(n19835), .A2(n19834), .ZN(n19870) );
  INV_X1 U22770 ( .A(n19870), .ZN(n19837) );
  NOR3_X1 U22771 ( .A1(n19837), .A2(P1_REIP_REG_7__SCAN_IN), .A3(n19836), .ZN(
        n19838) );
  AOI211_X1 U22772 ( .C1(n19876), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n19879), .B(n19838), .ZN(n19844) );
  AOI22_X1 U22773 ( .A1(P1_EBX_REG_7__SCAN_IN), .A2(n19875), .B1(n19884), .B2(
        n19893), .ZN(n19843) );
  NAND2_X1 U22774 ( .A1(n19896), .A2(n19857), .ZN(n19842) );
  INV_X1 U22775 ( .A(n19839), .ZN(n19840) );
  NAND2_X1 U22776 ( .A1(n19852), .A2(n19840), .ZN(n19841) );
  AND4_X1 U22777 ( .A1(n19844), .A2(n19843), .A3(n19842), .A4(n19841), .ZN(
        n19845) );
  OAI21_X1 U22778 ( .B1(n19854), .B2(n19846), .A(n19845), .ZN(P1_U2833) );
  INV_X1 U22779 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n19855) );
  NAND3_X1 U22780 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19870), .A3(n19855), 
        .ZN(n19847) );
  OAI211_X1 U22781 ( .C1(n19867), .C2(n19848), .A(n19864), .B(n19847), .ZN(
        n19849) );
  AOI21_X1 U22782 ( .B1(P1_EBX_REG_6__SCAN_IN), .B2(n19875), .A(n19849), .ZN(
        n19860) );
  INV_X1 U22783 ( .A(n19850), .ZN(n19851) );
  NAND2_X1 U22784 ( .A1(n19852), .A2(n19851), .ZN(n19853) );
  OAI21_X1 U22785 ( .B1(n19855), .B2(n19854), .A(n19853), .ZN(n19856) );
  AOI21_X1 U22786 ( .B1(n19858), .B2(n19857), .A(n19856), .ZN(n19859) );
  OAI211_X1 U22787 ( .C1(n19862), .C2(n19861), .A(n19860), .B(n19859), .ZN(
        P1_U2834) );
  INV_X1 U22788 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n19869) );
  INV_X1 U22789 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19866) );
  AOI22_X1 U22790 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(n19875), .B1(n19884), .B2(
        n19863), .ZN(n19865) );
  OAI211_X1 U22791 ( .C1(n19867), .C2(n19866), .A(n19865), .B(n19864), .ZN(
        n19868) );
  AOI221_X1 U22792 ( .B1(n19880), .B2(P1_REIP_REG_5__SCAN_IN), .C1(n19870), 
        .C2(n19869), .A(n19868), .ZN(n19873) );
  NAND2_X1 U22793 ( .A1(n19889), .A2(n19871), .ZN(n19872) );
  OAI211_X1 U22794 ( .C1(n19892), .C2(n19874), .A(n19873), .B(n19872), .ZN(
        P1_U2835) );
  AOI22_X1 U22795 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19876), .B1(
        P1_EBX_REG_4__SCAN_IN), .B2(n19875), .ZN(n19877) );
  INV_X1 U22796 ( .A(n19877), .ZN(n19878) );
  AOI211_X1 U22797 ( .C1(P1_REIP_REG_4__SCAN_IN), .C2(n19880), .A(n19879), .B(
        n19878), .ZN(n19891) );
  NAND2_X1 U22798 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n19881) );
  NOR3_X1 U22799 ( .A1(n19882), .A2(P1_REIP_REG_4__SCAN_IN), .A3(n19881), .ZN(
        n19883) );
  AOI21_X1 U22800 ( .B1(n19973), .B2(n19884), .A(n19883), .ZN(n19885) );
  OAI21_X1 U22801 ( .B1(n19887), .B2(n19886), .A(n19885), .ZN(n19888) );
  AOI21_X1 U22802 ( .B1(n19889), .B2(n19967), .A(n19888), .ZN(n19890) );
  OAI211_X1 U22803 ( .C1(n19971), .C2(n19892), .A(n19891), .B(n19890), .ZN(
        P1_U2836) );
  AOI22_X1 U22804 ( .A1(n19896), .A2(n19895), .B1(n19894), .B2(n19893), .ZN(
        n19897) );
  OAI21_X1 U22805 ( .B1(n19899), .B2(n19898), .A(n19897), .ZN(P1_U2865) );
  AOI22_X1 U22806 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n19903), .B1(n19929), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19900) );
  OAI21_X1 U22807 ( .B1(n19902), .B2(n19901), .A(n19900), .ZN(P1_U2921) );
  INV_X1 U22808 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n19905) );
  AOI22_X1 U22809 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19904) );
  OAI21_X1 U22810 ( .B1(n19905), .B2(n19932), .A(n19904), .ZN(P1_U2922) );
  INV_X1 U22811 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n19907) );
  AOI22_X1 U22812 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19906) );
  OAI21_X1 U22813 ( .B1(n19907), .B2(n19932), .A(n19906), .ZN(P1_U2923) );
  INV_X1 U22814 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n19909) );
  AOI22_X1 U22815 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19908) );
  OAI21_X1 U22816 ( .B1(n19909), .B2(n19932), .A(n19908), .ZN(P1_U2924) );
  INV_X1 U22817 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n19911) );
  AOI22_X1 U22818 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19910) );
  OAI21_X1 U22819 ( .B1(n19911), .B2(n19932), .A(n19910), .ZN(P1_U2925) );
  INV_X1 U22820 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n19913) );
  AOI22_X1 U22821 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19912) );
  OAI21_X1 U22822 ( .B1(n19913), .B2(n19932), .A(n19912), .ZN(P1_U2926) );
  INV_X1 U22823 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n19915) );
  AOI22_X1 U22824 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19914) );
  OAI21_X1 U22825 ( .B1(n19915), .B2(n19932), .A(n19914), .ZN(P1_U2927) );
  INV_X1 U22826 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n19917) );
  AOI22_X1 U22827 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19916) );
  OAI21_X1 U22828 ( .B1(n19917), .B2(n19932), .A(n19916), .ZN(P1_U2928) );
  AOI22_X1 U22829 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19918) );
  OAI21_X1 U22830 ( .B1(n14011), .B2(n19932), .A(n19918), .ZN(P1_U2929) );
  AOI22_X1 U22831 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19919) );
  OAI21_X1 U22832 ( .B1(n11610), .B2(n19932), .A(n19919), .ZN(P1_U2930) );
  AOI22_X1 U22833 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19920) );
  OAI21_X1 U22834 ( .B1(n11600), .B2(n19932), .A(n19920), .ZN(P1_U2931) );
  AOI22_X1 U22835 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19921) );
  OAI21_X1 U22836 ( .B1(n19922), .B2(n19932), .A(n19921), .ZN(P1_U2932) );
  AOI22_X1 U22837 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19923) );
  OAI21_X1 U22838 ( .B1(n19924), .B2(n19932), .A(n19923), .ZN(P1_U2933) );
  AOI22_X1 U22839 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19925) );
  OAI21_X1 U22840 ( .B1(n19926), .B2(n19932), .A(n19925), .ZN(P1_U2934) );
  AOI22_X1 U22841 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19927) );
  OAI21_X1 U22842 ( .B1(n19928), .B2(n19932), .A(n19927), .ZN(P1_U2935) );
  AOI22_X1 U22843 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n19930), .B1(n19929), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19931) );
  OAI21_X1 U22844 ( .B1(n19933), .B2(n19932), .A(n19931), .ZN(P1_U2936) );
  AOI22_X1 U22845 ( .A1(n19959), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n19934), .ZN(n19936) );
  NAND2_X1 U22846 ( .A1(n19944), .A2(n19935), .ZN(n19946) );
  NAND2_X1 U22847 ( .A1(n19936), .A2(n19946), .ZN(P1_U2945) );
  AOI22_X1 U22848 ( .A1(n19959), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n19954), .ZN(n19938) );
  NAND2_X1 U22849 ( .A1(n19944), .A2(n19937), .ZN(n19950) );
  NAND2_X1 U22850 ( .A1(n19938), .A2(n19950), .ZN(P1_U2947) );
  AOI22_X1 U22851 ( .A1(n19959), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n19954), .ZN(n19940) );
  NAND2_X1 U22852 ( .A1(n19944), .A2(n19939), .ZN(n19955) );
  NAND2_X1 U22853 ( .A1(n19940), .A2(n19955), .ZN(P1_U2949) );
  AOI22_X1 U22854 ( .A1(n19959), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n19954), .ZN(n19942) );
  NAND2_X1 U22855 ( .A1(n19944), .A2(n19941), .ZN(n19957) );
  NAND2_X1 U22856 ( .A1(n19942), .A2(n19957), .ZN(P1_U2950) );
  AOI22_X1 U22857 ( .A1(n19959), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n19954), .ZN(n19945) );
  NAND2_X1 U22858 ( .A1(n19944), .A2(n19943), .ZN(n19960) );
  NAND2_X1 U22859 ( .A1(n19945), .A2(n19960), .ZN(P1_U2951) );
  AOI22_X1 U22860 ( .A1(n19959), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n19954), .ZN(n19947) );
  NAND2_X1 U22861 ( .A1(n19947), .A2(n19946), .ZN(P1_U2960) );
  AOI22_X1 U22862 ( .A1(n19959), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n19954), .ZN(n19949) );
  NAND2_X1 U22863 ( .A1(n19949), .A2(n19948), .ZN(P1_U2961) );
  AOI22_X1 U22864 ( .A1(n19959), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n19954), .ZN(n19951) );
  NAND2_X1 U22865 ( .A1(n19951), .A2(n19950), .ZN(P1_U2962) );
  AOI22_X1 U22866 ( .A1(n19959), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n19954), .ZN(n19953) );
  NAND2_X1 U22867 ( .A1(n19953), .A2(n19952), .ZN(P1_U2963) );
  AOI22_X1 U22868 ( .A1(n19959), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n19954), .ZN(n19956) );
  NAND2_X1 U22869 ( .A1(n19956), .A2(n19955), .ZN(P1_U2964) );
  AOI22_X1 U22870 ( .A1(n19959), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n19954), .ZN(n19958) );
  NAND2_X1 U22871 ( .A1(n19958), .A2(n19957), .ZN(P1_U2965) );
  AOI22_X1 U22872 ( .A1(n19959), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n19954), .ZN(n19961) );
  NAND2_X1 U22873 ( .A1(n19961), .A2(n19960), .ZN(P1_U2966) );
  AOI22_X1 U22874 ( .A1(n19962), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20014), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n19970) );
  OAI21_X1 U22875 ( .B1(n19965), .B2(n19964), .A(n19963), .ZN(n19966) );
  INV_X1 U22876 ( .A(n19966), .ZN(n19974) );
  AOI22_X1 U22877 ( .A1(n19974), .A2(n19968), .B1(n14671), .B2(n19967), .ZN(
        n19969) );
  OAI211_X1 U22878 ( .C1(n19972), .C2(n19971), .A(n19970), .B(n19969), .ZN(
        P1_U2995) );
  AOI22_X1 U22879 ( .A1(n20014), .A2(P1_REIP_REG_4__SCAN_IN), .B1(n19981), 
        .B2(n19973), .ZN(n19979) );
  AOI22_X1 U22880 ( .A1(n19974), .A2(n20004), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n19983), .ZN(n19978) );
  OAI211_X1 U22881 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n19976), .B(n19975), .ZN(n19977) );
  NAND3_X1 U22882 ( .A1(n19979), .A2(n19978), .A3(n19977), .ZN(P1_U3027) );
  AOI22_X1 U22883 ( .A1(n20014), .A2(P1_REIP_REG_3__SCAN_IN), .B1(n19981), 
        .B2(n19980), .ZN(n19986) );
  INV_X1 U22884 ( .A(n19982), .ZN(n19984) );
  AOI22_X1 U22885 ( .A1(n19984), .A2(n20004), .B1(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n19983), .ZN(n19985) );
  OAI211_X1 U22886 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n19987), .A(
        n19986), .B(n19985), .ZN(P1_U3028) );
  NAND2_X1 U22887 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n19988), .ZN(
        n20003) );
  OAI21_X1 U22888 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n19990), .A(
        n19989), .ZN(n19991) );
  INV_X1 U22889 ( .A(n19991), .ZN(n20002) );
  INV_X1 U22890 ( .A(n19992), .ZN(n19999) );
  NAND3_X1 U22891 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n19994), .A3(
        n19993), .ZN(n19996) );
  NAND2_X1 U22892 ( .A1(n20014), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n19995) );
  OAI211_X1 U22893 ( .C1(n20017), .C2(n19997), .A(n19996), .B(n19995), .ZN(
        n19998) );
  AOI211_X1 U22894 ( .C1(n20000), .C2(n20004), .A(n19999), .B(n19998), .ZN(
        n20001) );
  OAI221_X1 U22895 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20003), .C1(
        n20762), .C2(n20002), .A(n20001), .ZN(P1_U3029) );
  NAND3_X1 U22896 ( .A1(n20006), .A2(n20005), .A3(n20004), .ZN(n20010) );
  OR3_X1 U22897 ( .A1(n20008), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n20007), .ZN(n20009) );
  OAI211_X1 U22898 ( .C1(n20012), .C2(n20011), .A(n20010), .B(n20009), .ZN(
        n20013) );
  INV_X1 U22899 ( .A(n20013), .ZN(n20016) );
  NAND2_X1 U22900 ( .A1(n20014), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20015) );
  OAI211_X1 U22901 ( .C1(n20018), .C2(n20017), .A(n20016), .B(n20015), .ZN(
        P1_U3030) );
  NOR2_X1 U22902 ( .A1(n20019), .A2(n20653), .ZN(P1_U3032) );
  AOI22_X1 U22903 ( .A1(DATAI_16_), .A2(n20057), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20056), .ZN(n20507) );
  NOR2_X2 U22904 ( .A1(n20055), .A2(n20024), .ZN(n20495) );
  NAND2_X1 U22905 ( .A1(n20655), .A2(n20274), .ZN(n20123) );
  AOI22_X1 U22906 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20056), .B1(DATAI_24_), 
        .B2(n20057), .ZN(n20456) );
  INV_X1 U22907 ( .A(n20456), .ZN(n20504) );
  AOI22_X1 U22908 ( .A1(n20495), .A2(n10081), .B1(n20058), .B2(n20504), .ZN(
        n20033) );
  NAND2_X1 U22909 ( .A1(n20029), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20444) );
  NAND2_X1 U22910 ( .A1(n20084), .A2(n20553), .ZN(n20025) );
  AOI21_X1 U22911 ( .B1(n20025), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20646), 
        .ZN(n20028) );
  OR2_X1 U22912 ( .A1(n20272), .A2(n20273), .ZN(n20093) );
  INV_X1 U22913 ( .A(n13646), .ZN(n20447) );
  OR2_X1 U22914 ( .A1(n20093), .A2(n20447), .ZN(n20030) );
  INV_X1 U22915 ( .A(n20326), .ZN(n20097) );
  OR2_X1 U22916 ( .A1(n20097), .A2(n20275), .ZN(n20159) );
  AOI22_X1 U22917 ( .A1(n20028), .A2(n20030), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20159), .ZN(n20026) );
  OAI211_X1 U22918 ( .C1(n10081), .C2(n20389), .A(n20328), .B(n20026), .ZN(
        n20061) );
  NOR2_X2 U22919 ( .A1(n20027), .A2(n20066), .ZN(n20496) );
  INV_X1 U22920 ( .A(n20028), .ZN(n20031) );
  OR2_X1 U22921 ( .A1(n20029), .A2(n12008), .ZN(n20330) );
  AOI22_X1 U22922 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20061), .B1(
        n20496), .B2(n20060), .ZN(n20032) );
  OAI211_X1 U22923 ( .C1(n20507), .C2(n20084), .A(n20033), .B(n20032), .ZN(
        P1_U3033) );
  AOI22_X1 U22924 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20056), .B1(DATAI_17_), 
        .B2(n20057), .ZN(n20513) );
  NOR2_X2 U22925 ( .A1(n20055), .A2(n11366), .ZN(n20508) );
  AOI22_X1 U22926 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20056), .B1(DATAI_25_), 
        .B2(n20057), .ZN(n20460) );
  INV_X1 U22927 ( .A(n20460), .ZN(n20510) );
  AOI22_X1 U22928 ( .A1(n20508), .A2(n10081), .B1(n20058), .B2(n20510), .ZN(
        n20036) );
  NOR2_X2 U22929 ( .A1(n20034), .A2(n20066), .ZN(n20509) );
  AOI22_X1 U22930 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20061), .B1(
        n20509), .B2(n20060), .ZN(n20035) );
  OAI211_X1 U22931 ( .C1(n20513), .C2(n20084), .A(n20036), .B(n20035), .ZN(
        P1_U3034) );
  AOI22_X1 U22932 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20056), .B1(DATAI_18_), 
        .B2(n20057), .ZN(n20519) );
  NOR2_X2 U22933 ( .A1(n20055), .A2(n12911), .ZN(n20514) );
  AOI22_X1 U22934 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20056), .B1(DATAI_26_), 
        .B2(n20057), .ZN(n20464) );
  INV_X1 U22935 ( .A(n20464), .ZN(n20516) );
  AOI22_X1 U22936 ( .A1(n20514), .A2(n10081), .B1(n20058), .B2(n20516), .ZN(
        n20039) );
  NOR2_X2 U22937 ( .A1(n20037), .A2(n20066), .ZN(n20515) );
  AOI22_X1 U22938 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20061), .B1(
        n20515), .B2(n20060), .ZN(n20038) );
  OAI211_X1 U22939 ( .C1(n20519), .C2(n20084), .A(n20039), .B(n20038), .ZN(
        P1_U3035) );
  AOI22_X1 U22940 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20056), .B1(DATAI_19_), 
        .B2(n20057), .ZN(n20525) );
  NOR2_X2 U22941 ( .A1(n20055), .A2(n20040), .ZN(n20520) );
  AOI22_X1 U22942 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20056), .B1(DATAI_27_), 
        .B2(n20057), .ZN(n20468) );
  INV_X1 U22943 ( .A(n20468), .ZN(n20522) );
  AOI22_X1 U22944 ( .A1(n20520), .A2(n10081), .B1(n20058), .B2(n20522), .ZN(
        n20043) );
  NOR2_X2 U22945 ( .A1(n20041), .A2(n20066), .ZN(n20521) );
  AOI22_X1 U22946 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20061), .B1(
        n20521), .B2(n20060), .ZN(n20042) );
  OAI211_X1 U22947 ( .C1(n20525), .C2(n20084), .A(n20043), .B(n20042), .ZN(
        P1_U3036) );
  AOI22_X1 U22948 ( .A1(DATAI_20_), .A2(n20057), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n20056), .ZN(n20531) );
  NOR2_X2 U22949 ( .A1(n20055), .A2(n20044), .ZN(n20526) );
  AOI22_X1 U22950 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20056), .B1(DATAI_28_), 
        .B2(n20057), .ZN(n20472) );
  INV_X1 U22951 ( .A(n20472), .ZN(n20528) );
  AOI22_X1 U22952 ( .A1(n20526), .A2(n10081), .B1(n20058), .B2(n20528), .ZN(
        n20047) );
  NOR2_X2 U22953 ( .A1(n20045), .A2(n20066), .ZN(n20527) );
  AOI22_X1 U22954 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20061), .B1(
        n20527), .B2(n20060), .ZN(n20046) );
  OAI211_X1 U22955 ( .C1(n20531), .C2(n20084), .A(n20047), .B(n20046), .ZN(
        P1_U3037) );
  AOI22_X1 U22956 ( .A1(DATAI_21_), .A2(n20057), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20056), .ZN(n20537) );
  NOR2_X2 U22957 ( .A1(n20055), .A2(n20048), .ZN(n20532) );
  AOI22_X1 U22958 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20056), .B1(DATAI_29_), 
        .B2(n20057), .ZN(n20476) );
  INV_X1 U22959 ( .A(n20476), .ZN(n20534) );
  AOI22_X1 U22960 ( .A1(n20532), .A2(n10081), .B1(n20058), .B2(n20534), .ZN(
        n20051) );
  NOR2_X2 U22961 ( .A1(n20049), .A2(n20066), .ZN(n20533) );
  AOI22_X1 U22962 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20061), .B1(
        n20533), .B2(n20060), .ZN(n20050) );
  OAI211_X1 U22963 ( .C1(n20537), .C2(n20084), .A(n20051), .B(n20050), .ZN(
        P1_U3038) );
  AOI22_X1 U22964 ( .A1(DATAI_22_), .A2(n20057), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n20056), .ZN(n20543) );
  NOR2_X2 U22965 ( .A1(n20055), .A2(n11566), .ZN(n20538) );
  AOI22_X1 U22966 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20056), .B1(DATAI_30_), 
        .B2(n20057), .ZN(n20480) );
  INV_X1 U22967 ( .A(n20480), .ZN(n20540) );
  AOI22_X1 U22968 ( .A1(n20538), .A2(n10081), .B1(n20058), .B2(n20540), .ZN(
        n20054) );
  NOR2_X2 U22969 ( .A1(n20052), .A2(n20066), .ZN(n20539) );
  AOI22_X1 U22970 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20061), .B1(
        n20539), .B2(n20060), .ZN(n20053) );
  OAI211_X1 U22971 ( .C1(n20543), .C2(n20084), .A(n20054), .B(n20053), .ZN(
        P1_U3039) );
  AOI22_X1 U22972 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20056), .B1(DATAI_23_), 
        .B2(n20057), .ZN(n20554) );
  NOR2_X2 U22973 ( .A1(n20055), .A2(n9769), .ZN(n20545) );
  AOI22_X1 U22974 ( .A1(DATAI_31_), .A2(n20057), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20056), .ZN(n20488) );
  INV_X1 U22975 ( .A(n20488), .ZN(n20548) );
  AOI22_X1 U22976 ( .A1(n20545), .A2(n10081), .B1(n20058), .B2(n20548), .ZN(
        n20063) );
  NOR2_X2 U22977 ( .A1(n20059), .A2(n20066), .ZN(n20547) );
  AOI22_X1 U22978 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20061), .B1(
        n20547), .B2(n20060), .ZN(n20062) );
  OAI211_X1 U22979 ( .C1(n20554), .C2(n20084), .A(n20063), .B(n20062), .ZN(
        P1_U3040) );
  INV_X1 U22980 ( .A(n20093), .ZN(n20126) );
  INV_X1 U22981 ( .A(n20064), .ZN(n20416) );
  NOR2_X1 U22982 ( .A1(n20123), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20069) );
  INV_X1 U22983 ( .A(n20069), .ZN(n20065) );
  NOR2_X1 U22984 ( .A1(n20415), .A2(n20065), .ZN(n20085) );
  AOI21_X1 U22985 ( .B1(n20126), .B2(n20416), .A(n20085), .ZN(n20067) );
  OAI22_X1 U22986 ( .A1(n20067), .A2(n20646), .B1(n20065), .B2(n12008), .ZN(
        n20086) );
  AOI22_X1 U22987 ( .A1(n20496), .A2(n20086), .B1(n20495), .B2(n20085), .ZN(
        n20071) );
  OAI211_X1 U22988 ( .C1(n20127), .C2(n20640), .A(n20641), .B(n20067), .ZN(
        n20068) );
  OAI211_X1 U22989 ( .C1(n20641), .C2(n20069), .A(n20501), .B(n20068), .ZN(
        n20088) );
  INV_X1 U22990 ( .A(n20303), .ZN(n20413) );
  INV_X1 U22991 ( .A(n20507), .ZN(n20453) );
  AOI22_X1 U22992 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20088), .B1(
        n20116), .B2(n20453), .ZN(n20070) );
  OAI211_X1 U22993 ( .C1(n20456), .C2(n20084), .A(n20071), .B(n20070), .ZN(
        P1_U3041) );
  AOI22_X1 U22994 ( .A1(n20509), .A2(n20086), .B1(n20508), .B2(n20085), .ZN(
        n20073) );
  INV_X1 U22995 ( .A(n20513), .ZN(n20457) );
  AOI22_X1 U22996 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20088), .B1(
        n20116), .B2(n20457), .ZN(n20072) );
  OAI211_X1 U22997 ( .C1(n20460), .C2(n20084), .A(n20073), .B(n20072), .ZN(
        P1_U3042) );
  AOI22_X1 U22998 ( .A1(n20515), .A2(n20086), .B1(n20514), .B2(n20085), .ZN(
        n20075) );
  INV_X1 U22999 ( .A(n20084), .ZN(n20087) );
  AOI22_X1 U23000 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20088), .B1(
        n20087), .B2(n20516), .ZN(n20074) );
  OAI211_X1 U23001 ( .C1(n20519), .C2(n20114), .A(n20075), .B(n20074), .ZN(
        P1_U3043) );
  AOI22_X1 U23002 ( .A1(n20521), .A2(n20086), .B1(n20520), .B2(n20085), .ZN(
        n20077) );
  AOI22_X1 U23003 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20088), .B1(
        n20087), .B2(n20522), .ZN(n20076) );
  OAI211_X1 U23004 ( .C1(n20525), .C2(n20114), .A(n20077), .B(n20076), .ZN(
        P1_U3044) );
  AOI22_X1 U23005 ( .A1(n20527), .A2(n20086), .B1(n20526), .B2(n20085), .ZN(
        n20079) );
  INV_X1 U23006 ( .A(n20531), .ZN(n20469) );
  AOI22_X1 U23007 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20088), .B1(
        n20116), .B2(n20469), .ZN(n20078) );
  OAI211_X1 U23008 ( .C1(n20472), .C2(n20084), .A(n20079), .B(n20078), .ZN(
        P1_U3045) );
  AOI22_X1 U23009 ( .A1(n20533), .A2(n20086), .B1(n20532), .B2(n20085), .ZN(
        n20081) );
  INV_X1 U23010 ( .A(n20537), .ZN(n20473) );
  AOI22_X1 U23011 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20088), .B1(
        n20116), .B2(n20473), .ZN(n20080) );
  OAI211_X1 U23012 ( .C1(n20476), .C2(n20084), .A(n20081), .B(n20080), .ZN(
        P1_U3046) );
  AOI22_X1 U23013 ( .A1(n20539), .A2(n20086), .B1(n20538), .B2(n20085), .ZN(
        n20083) );
  INV_X1 U23014 ( .A(n20543), .ZN(n20477) );
  AOI22_X1 U23015 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20088), .B1(
        n20116), .B2(n20477), .ZN(n20082) );
  OAI211_X1 U23016 ( .C1(n20480), .C2(n20084), .A(n20083), .B(n20082), .ZN(
        P1_U3047) );
  AOI22_X1 U23017 ( .A1(n20547), .A2(n20086), .B1(n20545), .B2(n20085), .ZN(
        n20090) );
  AOI22_X1 U23018 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20088), .B1(
        n20087), .B2(n20548), .ZN(n20089) );
  OAI211_X1 U23019 ( .C1(n20554), .C2(n20114), .A(n20090), .B(n20089), .ZN(
        P1_U3048) );
  INV_X1 U23020 ( .A(n20123), .ZN(n20091) );
  NAND2_X1 U23021 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20091), .ZN(
        n20130) );
  NOR2_X1 U23022 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20130), .ZN(
        n20115) );
  AOI22_X1 U23023 ( .A1(n20116), .A2(n20504), .B1(n20495), .B2(n20115), .ZN(
        n20101) );
  NAND2_X1 U23024 ( .A1(n20153), .A2(n20114), .ZN(n20092) );
  AOI21_X1 U23025 ( .B1(n20092), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20646), 
        .ZN(n20096) );
  OR2_X1 U23026 ( .A1(n20093), .A2(n13646), .ZN(n20098) );
  NOR2_X1 U23027 ( .A1(n20115), .A2(n20389), .ZN(n20094) );
  AOI21_X1 U23028 ( .B1(n20096), .B2(n20098), .A(n20094), .ZN(n20095) );
  OAI21_X1 U23029 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20326), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20213) );
  NAND3_X1 U23030 ( .A1(n20328), .A2(n20095), .A3(n20213), .ZN(n20118) );
  INV_X1 U23031 ( .A(n20096), .ZN(n20099) );
  NAND2_X1 U23032 ( .A1(n20097), .A2(n20655), .ZN(n20216) );
  AOI22_X1 U23033 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20118), .B1(
        n20496), .B2(n20117), .ZN(n20100) );
  OAI211_X1 U23034 ( .C1(n20507), .C2(n20153), .A(n20101), .B(n20100), .ZN(
        P1_U3049) );
  AOI22_X1 U23035 ( .A1(n20145), .A2(n20457), .B1(n20508), .B2(n20115), .ZN(
        n20103) );
  AOI22_X1 U23036 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20118), .B1(
        n20509), .B2(n20117), .ZN(n20102) );
  OAI211_X1 U23037 ( .C1(n20460), .C2(n20114), .A(n20103), .B(n20102), .ZN(
        P1_U3050) );
  INV_X1 U23038 ( .A(n20519), .ZN(n20461) );
  AOI22_X1 U23039 ( .A1(n20145), .A2(n20461), .B1(n20514), .B2(n20115), .ZN(
        n20105) );
  AOI22_X1 U23040 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20118), .B1(
        n20515), .B2(n20117), .ZN(n20104) );
  OAI211_X1 U23041 ( .C1(n20464), .C2(n20114), .A(n20105), .B(n20104), .ZN(
        P1_U3051) );
  AOI22_X1 U23042 ( .A1(n20116), .A2(n20522), .B1(n20520), .B2(n20115), .ZN(
        n20107) );
  AOI22_X1 U23043 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20118), .B1(
        n20521), .B2(n20117), .ZN(n20106) );
  OAI211_X1 U23044 ( .C1(n20525), .C2(n20153), .A(n20107), .B(n20106), .ZN(
        P1_U3052) );
  AOI22_X1 U23045 ( .A1(n20145), .A2(n20469), .B1(n20526), .B2(n20115), .ZN(
        n20109) );
  AOI22_X1 U23046 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20118), .B1(
        n20527), .B2(n20117), .ZN(n20108) );
  OAI211_X1 U23047 ( .C1(n20472), .C2(n20114), .A(n20109), .B(n20108), .ZN(
        P1_U3053) );
  AOI22_X1 U23048 ( .A1(n20116), .A2(n20534), .B1(n20532), .B2(n20115), .ZN(
        n20111) );
  AOI22_X1 U23049 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20118), .B1(
        n20533), .B2(n20117), .ZN(n20110) );
  OAI211_X1 U23050 ( .C1(n20537), .C2(n20153), .A(n20111), .B(n20110), .ZN(
        P1_U3054) );
  AOI22_X1 U23051 ( .A1(n20145), .A2(n20477), .B1(n20538), .B2(n20115), .ZN(
        n20113) );
  AOI22_X1 U23052 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20118), .B1(
        n20539), .B2(n20117), .ZN(n20112) );
  OAI211_X1 U23053 ( .C1(n20480), .C2(n20114), .A(n20113), .B(n20112), .ZN(
        P1_U3055) );
  AOI22_X1 U23054 ( .A1(n20116), .A2(n20548), .B1(n20545), .B2(n20115), .ZN(
        n20120) );
  AOI22_X1 U23055 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20118), .B1(
        n20547), .B2(n20117), .ZN(n20119) );
  OAI211_X1 U23056 ( .C1(n20554), .C2(n20153), .A(n20120), .B(n20119), .ZN(
        P1_U3056) );
  INV_X1 U23057 ( .A(n20354), .ZN(n20121) );
  NOR2_X1 U23058 ( .A1(n20489), .A2(n20123), .ZN(n20148) );
  AOI22_X1 U23059 ( .A1(n20145), .A2(n20504), .B1(n20495), .B2(n20148), .ZN(
        n20134) );
  NOR2_X1 U23060 ( .A1(n20125), .A2(n20124), .ZN(n20490) );
  AOI21_X1 U23061 ( .B1(n20126), .B2(n20490), .A(n20148), .ZN(n20132) );
  AOI21_X1 U23062 ( .B1(n20127), .B2(n20641), .A(n20499), .ZN(n20131) );
  INV_X1 U23063 ( .A(n20131), .ZN(n20128) );
  AOI22_X1 U23064 ( .A1(n20132), .A2(n20128), .B1(n20646), .B2(n20130), .ZN(
        n20129) );
  NAND2_X1 U23065 ( .A1(n20501), .A2(n20129), .ZN(n20150) );
  OAI22_X1 U23066 ( .A1(n20132), .A2(n20131), .B1(n20417), .B2(n20130), .ZN(
        n20149) );
  AOI22_X1 U23067 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20150), .B1(
        n20496), .B2(n20149), .ZN(n20133) );
  OAI211_X1 U23068 ( .C1(n20507), .C2(n20178), .A(n20134), .B(n20133), .ZN(
        P1_U3057) );
  AOI22_X1 U23069 ( .A1(n20180), .A2(n20457), .B1(n20508), .B2(n20148), .ZN(
        n20136) );
  AOI22_X1 U23070 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20150), .B1(
        n20509), .B2(n20149), .ZN(n20135) );
  OAI211_X1 U23071 ( .C1(n20460), .C2(n20153), .A(n20136), .B(n20135), .ZN(
        P1_U3058) );
  AOI22_X1 U23072 ( .A1(n20180), .A2(n20461), .B1(n20514), .B2(n20148), .ZN(
        n20138) );
  AOI22_X1 U23073 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20150), .B1(
        n20515), .B2(n20149), .ZN(n20137) );
  OAI211_X1 U23074 ( .C1(n20464), .C2(n20153), .A(n20138), .B(n20137), .ZN(
        P1_U3059) );
  INV_X1 U23075 ( .A(n20525), .ZN(n20465) );
  AOI22_X1 U23076 ( .A1(n20180), .A2(n20465), .B1(n20520), .B2(n20148), .ZN(
        n20140) );
  AOI22_X1 U23077 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20150), .B1(
        n20521), .B2(n20149), .ZN(n20139) );
  OAI211_X1 U23078 ( .C1(n20468), .C2(n20153), .A(n20140), .B(n20139), .ZN(
        P1_U3060) );
  AOI22_X1 U23079 ( .A1(n20180), .A2(n20469), .B1(n20526), .B2(n20148), .ZN(
        n20142) );
  AOI22_X1 U23080 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20150), .B1(
        n20527), .B2(n20149), .ZN(n20141) );
  OAI211_X1 U23081 ( .C1(n20472), .C2(n20153), .A(n20142), .B(n20141), .ZN(
        P1_U3061) );
  AOI22_X1 U23082 ( .A1(n20180), .A2(n20473), .B1(n20532), .B2(n20148), .ZN(
        n20144) );
  AOI22_X1 U23083 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20150), .B1(
        n20533), .B2(n20149), .ZN(n20143) );
  OAI211_X1 U23084 ( .C1(n20476), .C2(n20153), .A(n20144), .B(n20143), .ZN(
        P1_U3062) );
  AOI22_X1 U23085 ( .A1(n20145), .A2(n20540), .B1(n20538), .B2(n20148), .ZN(
        n20147) );
  AOI22_X1 U23086 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20150), .B1(
        n20539), .B2(n20149), .ZN(n20146) );
  OAI211_X1 U23087 ( .C1(n20543), .C2(n20178), .A(n20147), .B(n20146), .ZN(
        P1_U3063) );
  INV_X1 U23088 ( .A(n20554), .ZN(n20483) );
  AOI22_X1 U23089 ( .A1(n20180), .A2(n20483), .B1(n20545), .B2(n20148), .ZN(
        n20152) );
  AOI22_X1 U23090 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20150), .B1(
        n20547), .B2(n20149), .ZN(n20151) );
  OAI211_X1 U23091 ( .C1(n20488), .C2(n20153), .A(n20152), .B(n20151), .ZN(
        P1_U3064) );
  NOR2_X1 U23092 ( .A1(n13568), .A2(n20157), .ZN(n20241) );
  NAND3_X1 U23093 ( .A1(n20241), .A2(n20641), .A3(n13646), .ZN(n20158) );
  OAI21_X1 U23094 ( .B1(n20159), .B2(n20444), .A(n20158), .ZN(n20179) );
  AOI22_X1 U23095 ( .A1(n20496), .A2(n20179), .B1(n20495), .B2(n9737), .ZN(
        n20165) );
  AOI21_X1 U23096 ( .B1(n20178), .B2(n20208), .A(n20640), .ZN(n20160) );
  AOI21_X1 U23097 ( .B1(n20241), .B2(n13646), .A(n20160), .ZN(n20161) );
  NOR2_X1 U23098 ( .A1(n20161), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20163) );
  AOI22_X1 U23099 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20181), .B1(
        n20180), .B2(n20504), .ZN(n20164) );
  OAI211_X1 U23100 ( .C1(n20507), .C2(n20208), .A(n20165), .B(n20164), .ZN(
        P1_U3065) );
  AOI22_X1 U23101 ( .A1(n20509), .A2(n20179), .B1(n20508), .B2(n9737), .ZN(
        n20167) );
  AOI22_X1 U23102 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20181), .B1(
        n20200), .B2(n20457), .ZN(n20166) );
  OAI211_X1 U23103 ( .C1(n20460), .C2(n20178), .A(n20167), .B(n20166), .ZN(
        P1_U3066) );
  AOI22_X1 U23104 ( .A1(n20515), .A2(n20179), .B1(n20514), .B2(n9737), .ZN(
        n20169) );
  AOI22_X1 U23105 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20181), .B1(
        n20200), .B2(n20461), .ZN(n20168) );
  OAI211_X1 U23106 ( .C1(n20464), .C2(n20178), .A(n20169), .B(n20168), .ZN(
        P1_U3067) );
  AOI22_X1 U23107 ( .A1(n20521), .A2(n20179), .B1(n20520), .B2(n9737), .ZN(
        n20171) );
  AOI22_X1 U23108 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20181), .B1(
        n20180), .B2(n20522), .ZN(n20170) );
  OAI211_X1 U23109 ( .C1(n20525), .C2(n20208), .A(n20171), .B(n20170), .ZN(
        P1_U3068) );
  AOI22_X1 U23110 ( .A1(n20527), .A2(n20179), .B1(n20526), .B2(n9737), .ZN(
        n20173) );
  AOI22_X1 U23111 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20181), .B1(
        n20200), .B2(n20469), .ZN(n20172) );
  OAI211_X1 U23112 ( .C1(n20472), .C2(n20178), .A(n20173), .B(n20172), .ZN(
        P1_U3069) );
  AOI22_X1 U23113 ( .A1(n20533), .A2(n20179), .B1(n20532), .B2(n9737), .ZN(
        n20175) );
  AOI22_X1 U23114 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20181), .B1(
        n20180), .B2(n20534), .ZN(n20174) );
  OAI211_X1 U23115 ( .C1(n20537), .C2(n20208), .A(n20175), .B(n20174), .ZN(
        P1_U3070) );
  AOI22_X1 U23116 ( .A1(n20539), .A2(n20179), .B1(n20538), .B2(n9737), .ZN(
        n20177) );
  AOI22_X1 U23117 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20181), .B1(
        n20200), .B2(n20477), .ZN(n20176) );
  OAI211_X1 U23118 ( .C1(n20480), .C2(n20178), .A(n20177), .B(n20176), .ZN(
        P1_U3071) );
  AOI22_X1 U23119 ( .A1(n20547), .A2(n20179), .B1(n20545), .B2(n9737), .ZN(
        n20183) );
  AOI22_X1 U23120 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20181), .B1(
        n20180), .B2(n20548), .ZN(n20182) );
  OAI211_X1 U23121 ( .C1(n20554), .C2(n20208), .A(n20183), .B(n20182), .ZN(
        P1_U3072) );
  NOR2_X1 U23122 ( .A1(n20209), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20187) );
  INV_X1 U23123 ( .A(n20187), .ZN(n20184) );
  NOR2_X1 U23124 ( .A1(n20415), .A2(n20184), .ZN(n20203) );
  AOI21_X1 U23125 ( .B1(n20241), .B2(n20416), .A(n20203), .ZN(n20185) );
  OAI22_X1 U23126 ( .A1(n20185), .A2(n20646), .B1(n20184), .B2(n20417), .ZN(
        n20204) );
  AOI22_X1 U23127 ( .A1(n20496), .A2(n20204), .B1(n20495), .B2(n20203), .ZN(
        n20189) );
  OAI211_X1 U23128 ( .C1(n20639), .C2(n20640), .A(n20641), .B(n20185), .ZN(
        n20186) );
  OAI211_X1 U23129 ( .C1(n20641), .C2(n20187), .A(n20501), .B(n20186), .ZN(
        n20205) );
  AOI22_X1 U23130 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20205), .B1(
        n20200), .B2(n20504), .ZN(n20188) );
  OAI211_X1 U23131 ( .C1(n20507), .C2(n20239), .A(n20189), .B(n20188), .ZN(
        P1_U3073) );
  AOI22_X1 U23132 ( .A1(n20509), .A2(n20204), .B1(n20508), .B2(n20203), .ZN(
        n20191) );
  AOI22_X1 U23133 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20205), .B1(
        n20200), .B2(n20510), .ZN(n20190) );
  OAI211_X1 U23134 ( .C1(n20513), .C2(n20239), .A(n20191), .B(n20190), .ZN(
        P1_U3074) );
  AOI22_X1 U23135 ( .A1(n20515), .A2(n20204), .B1(n20514), .B2(n20203), .ZN(
        n20193) );
  AOI22_X1 U23136 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20205), .B1(
        n20200), .B2(n20516), .ZN(n20192) );
  OAI211_X1 U23137 ( .C1(n20519), .C2(n20239), .A(n20193), .B(n20192), .ZN(
        P1_U3075) );
  AOI22_X1 U23138 ( .A1(n20521), .A2(n20204), .B1(n20520), .B2(n20203), .ZN(
        n20195) );
  AOI22_X1 U23139 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20205), .B1(
        n20200), .B2(n20522), .ZN(n20194) );
  OAI211_X1 U23140 ( .C1(n20525), .C2(n20239), .A(n20195), .B(n20194), .ZN(
        P1_U3076) );
  AOI22_X1 U23141 ( .A1(n20527), .A2(n20204), .B1(n20526), .B2(n20203), .ZN(
        n20197) );
  AOI22_X1 U23142 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20205), .B1(
        n20200), .B2(n20528), .ZN(n20196) );
  OAI211_X1 U23143 ( .C1(n20531), .C2(n20239), .A(n20197), .B(n20196), .ZN(
        P1_U3077) );
  AOI22_X1 U23144 ( .A1(n20533), .A2(n20204), .B1(n20532), .B2(n20203), .ZN(
        n20199) );
  AOI22_X1 U23145 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20205), .B1(
        n20200), .B2(n20534), .ZN(n20198) );
  OAI211_X1 U23146 ( .C1(n20537), .C2(n20239), .A(n20199), .B(n20198), .ZN(
        P1_U3078) );
  AOI22_X1 U23147 ( .A1(n20539), .A2(n20204), .B1(n20538), .B2(n20203), .ZN(
        n20202) );
  AOI22_X1 U23148 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20205), .B1(
        n20200), .B2(n20540), .ZN(n20201) );
  OAI211_X1 U23149 ( .C1(n20543), .C2(n20239), .A(n20202), .B(n20201), .ZN(
        P1_U3079) );
  AOI22_X1 U23150 ( .A1(n20547), .A2(n20204), .B1(n20545), .B2(n20203), .ZN(
        n20207) );
  INV_X1 U23151 ( .A(n20239), .ZN(n20229) );
  AOI22_X1 U23152 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20205), .B1(
        n20229), .B2(n20483), .ZN(n20206) );
  OAI211_X1 U23153 ( .C1(n20488), .C2(n20208), .A(n20207), .B(n20206), .ZN(
        P1_U3080) );
  NOR2_X1 U23154 ( .A1(n20493), .A2(n20209), .ZN(n20245) );
  NAND2_X1 U23155 ( .A1(n20415), .A2(n20245), .ZN(n20212) );
  AOI22_X1 U23156 ( .A1(n20495), .A2(n20234), .B1(n20258), .B2(n20453), .ZN(
        n20220) );
  NAND2_X1 U23157 ( .A1(n20267), .A2(n20239), .ZN(n20211) );
  AOI21_X1 U23158 ( .B1(n20211), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20646), 
        .ZN(n20215) );
  NAND2_X1 U23159 ( .A1(n20241), .A2(n20447), .ZN(n20217) );
  AOI22_X1 U23160 ( .A1(n20215), .A2(n20217), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20212), .ZN(n20214) );
  NAND3_X1 U23161 ( .A1(n20450), .A2(n20214), .A3(n20213), .ZN(n20236) );
  INV_X1 U23162 ( .A(n20215), .ZN(n20218) );
  OAI22_X1 U23163 ( .A1(n20218), .A2(n20217), .B1(n20216), .B2(n20444), .ZN(
        n20235) );
  AOI22_X1 U23164 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20236), .B1(
        n20496), .B2(n20235), .ZN(n20219) );
  OAI211_X1 U23165 ( .C1(n20456), .C2(n20239), .A(n20220), .B(n20219), .ZN(
        P1_U3081) );
  AOI22_X1 U23166 ( .A1(n20508), .A2(n20234), .B1(n20229), .B2(n20510), .ZN(
        n20222) );
  AOI22_X1 U23167 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20236), .B1(
        n20509), .B2(n20235), .ZN(n20221) );
  OAI211_X1 U23168 ( .C1(n20513), .C2(n20267), .A(n20222), .B(n20221), .ZN(
        P1_U3082) );
  AOI22_X1 U23169 ( .A1(n20514), .A2(n20234), .B1(n20229), .B2(n20516), .ZN(
        n20224) );
  AOI22_X1 U23170 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20236), .B1(
        n20515), .B2(n20235), .ZN(n20223) );
  OAI211_X1 U23171 ( .C1(n20519), .C2(n20267), .A(n20224), .B(n20223), .ZN(
        P1_U3083) );
  AOI22_X1 U23172 ( .A1(n20520), .A2(n20234), .B1(n20229), .B2(n20522), .ZN(
        n20226) );
  AOI22_X1 U23173 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20236), .B1(
        n20521), .B2(n20235), .ZN(n20225) );
  OAI211_X1 U23174 ( .C1(n20525), .C2(n20267), .A(n20226), .B(n20225), .ZN(
        P1_U3084) );
  AOI22_X1 U23175 ( .A1(n20526), .A2(n20234), .B1(n20258), .B2(n20469), .ZN(
        n20228) );
  AOI22_X1 U23176 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20236), .B1(
        n20527), .B2(n20235), .ZN(n20227) );
  OAI211_X1 U23177 ( .C1(n20472), .C2(n20239), .A(n20228), .B(n20227), .ZN(
        P1_U3085) );
  AOI22_X1 U23178 ( .A1(n20532), .A2(n20234), .B1(n20229), .B2(n20534), .ZN(
        n20231) );
  AOI22_X1 U23179 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20236), .B1(
        n20533), .B2(n20235), .ZN(n20230) );
  OAI211_X1 U23180 ( .C1(n20537), .C2(n20267), .A(n20231), .B(n20230), .ZN(
        P1_U3086) );
  AOI22_X1 U23181 ( .A1(n20538), .A2(n20234), .B1(n20258), .B2(n20477), .ZN(
        n20233) );
  AOI22_X1 U23182 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20236), .B1(
        n20539), .B2(n20235), .ZN(n20232) );
  OAI211_X1 U23183 ( .C1(n20480), .C2(n20239), .A(n20233), .B(n20232), .ZN(
        P1_U3087) );
  AOI22_X1 U23184 ( .A1(n20545), .A2(n20234), .B1(n20258), .B2(n20483), .ZN(
        n20238) );
  AOI22_X1 U23185 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20236), .B1(
        n20547), .B2(n20235), .ZN(n20237) );
  OAI211_X1 U23186 ( .C1(n20488), .C2(n20239), .A(n20238), .B(n20237), .ZN(
        P1_U3088) );
  INV_X1 U23187 ( .A(n20240), .ZN(n20262) );
  AOI21_X1 U23188 ( .B1(n20241), .B2(n20490), .A(n20262), .ZN(n20243) );
  INV_X1 U23189 ( .A(n20245), .ZN(n20242) );
  OAI22_X1 U23190 ( .A1(n20243), .A2(n20646), .B1(n20242), .B2(n12008), .ZN(
        n20263) );
  AOI22_X1 U23191 ( .A1(n20496), .A2(n20263), .B1(n20262), .B2(n20495), .ZN(
        n20247) );
  OAI211_X1 U23192 ( .C1(n20499), .C2(n20639), .A(n20641), .B(n20243), .ZN(
        n20244) );
  OAI211_X1 U23193 ( .C1(n20641), .C2(n20245), .A(n20501), .B(n20244), .ZN(
        n20264) );
  AOI22_X1 U23194 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20264), .B1(
        n20295), .B2(n20453), .ZN(n20246) );
  OAI211_X1 U23195 ( .C1(n20456), .C2(n20267), .A(n20247), .B(n20246), .ZN(
        P1_U3089) );
  AOI22_X1 U23196 ( .A1(n20509), .A2(n20263), .B1(n20262), .B2(n20508), .ZN(
        n20249) );
  AOI22_X1 U23197 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20264), .B1(
        n20295), .B2(n20457), .ZN(n20248) );
  OAI211_X1 U23198 ( .C1(n20460), .C2(n20267), .A(n20249), .B(n20248), .ZN(
        P1_U3090) );
  AOI22_X1 U23199 ( .A1(n20515), .A2(n20263), .B1(n20262), .B2(n20514), .ZN(
        n20251) );
  AOI22_X1 U23200 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20264), .B1(
        n20295), .B2(n20461), .ZN(n20250) );
  OAI211_X1 U23201 ( .C1(n20464), .C2(n20267), .A(n20251), .B(n20250), .ZN(
        P1_U3091) );
  AOI22_X1 U23202 ( .A1(n20521), .A2(n20263), .B1(n20262), .B2(n20520), .ZN(
        n20253) );
  AOI22_X1 U23203 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20264), .B1(
        n20295), .B2(n20465), .ZN(n20252) );
  OAI211_X1 U23204 ( .C1(n20468), .C2(n20267), .A(n20253), .B(n20252), .ZN(
        P1_U3092) );
  AOI22_X1 U23205 ( .A1(n20527), .A2(n20263), .B1(n20262), .B2(n20526), .ZN(
        n20255) );
  AOI22_X1 U23206 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20264), .B1(
        n20295), .B2(n20469), .ZN(n20254) );
  OAI211_X1 U23207 ( .C1(n20472), .C2(n20267), .A(n20255), .B(n20254), .ZN(
        P1_U3093) );
  AOI22_X1 U23208 ( .A1(n20533), .A2(n20263), .B1(n20262), .B2(n20532), .ZN(
        n20257) );
  AOI22_X1 U23209 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20264), .B1(
        n20258), .B2(n20534), .ZN(n20256) );
  OAI211_X1 U23210 ( .C1(n20537), .C2(n20261), .A(n20257), .B(n20256), .ZN(
        P1_U3094) );
  AOI22_X1 U23211 ( .A1(n20539), .A2(n20263), .B1(n20262), .B2(n20538), .ZN(
        n20260) );
  AOI22_X1 U23212 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20264), .B1(
        n20258), .B2(n20540), .ZN(n20259) );
  OAI211_X1 U23213 ( .C1(n20543), .C2(n20261), .A(n20260), .B(n20259), .ZN(
        P1_U3095) );
  AOI22_X1 U23214 ( .A1(n20547), .A2(n20263), .B1(n20262), .B2(n20545), .ZN(
        n20266) );
  AOI22_X1 U23215 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20264), .B1(
        n20295), .B2(n20483), .ZN(n20265) );
  OAI211_X1 U23216 ( .C1(n20488), .C2(n20267), .A(n20266), .B(n20265), .ZN(
        P1_U3096) );
  INV_X1 U23217 ( .A(n20268), .ZN(n20269) );
  INV_X1 U23218 ( .A(n20647), .ZN(n20271) );
  INV_X1 U23219 ( .A(n20272), .ZN(n20645) );
  NAND2_X1 U23220 ( .A1(n20274), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20355) );
  AOI21_X1 U23221 ( .B1(n20356), .B2(n13646), .A(n10080), .ZN(n20277) );
  NAND2_X1 U23222 ( .A1(n20275), .A2(n20326), .ZN(n20391) );
  OAI22_X1 U23223 ( .A1(n20277), .A2(n20646), .B1(n20330), .B2(n20391), .ZN(
        n20294) );
  AOI22_X1 U23224 ( .A1(n20496), .A2(n20294), .B1(n10080), .B2(n20495), .ZN(
        n20281) );
  INV_X1 U23225 ( .A(n20323), .ZN(n20276) );
  OAI21_X1 U23226 ( .B1(n20276), .B2(n20295), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20278) );
  NAND2_X1 U23227 ( .A1(n20278), .A2(n20277), .ZN(n20279) );
  AOI22_X1 U23228 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20296), .B1(
        n20295), .B2(n20504), .ZN(n20280) );
  OAI211_X1 U23229 ( .C1(n20507), .C2(n20323), .A(n20281), .B(n20280), .ZN(
        P1_U3097) );
  AOI22_X1 U23230 ( .A1(n20509), .A2(n20294), .B1(n10080), .B2(n20508), .ZN(
        n20283) );
  AOI22_X1 U23231 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20296), .B1(
        n20295), .B2(n20510), .ZN(n20282) );
  OAI211_X1 U23232 ( .C1(n20513), .C2(n20323), .A(n20283), .B(n20282), .ZN(
        P1_U3098) );
  AOI22_X1 U23233 ( .A1(n20515), .A2(n20294), .B1(n10080), .B2(n20514), .ZN(
        n20285) );
  AOI22_X1 U23234 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20296), .B1(
        n20295), .B2(n20516), .ZN(n20284) );
  OAI211_X1 U23235 ( .C1(n20519), .C2(n20323), .A(n20285), .B(n20284), .ZN(
        P1_U3099) );
  AOI22_X1 U23236 ( .A1(n20521), .A2(n20294), .B1(n10080), .B2(n20520), .ZN(
        n20287) );
  AOI22_X1 U23237 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20296), .B1(
        n20295), .B2(n20522), .ZN(n20286) );
  OAI211_X1 U23238 ( .C1(n20525), .C2(n20323), .A(n20287), .B(n20286), .ZN(
        P1_U3100) );
  AOI22_X1 U23239 ( .A1(n20527), .A2(n20294), .B1(n10080), .B2(n20526), .ZN(
        n20289) );
  AOI22_X1 U23240 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20296), .B1(
        n20295), .B2(n20528), .ZN(n20288) );
  OAI211_X1 U23241 ( .C1(n20531), .C2(n20323), .A(n20289), .B(n20288), .ZN(
        P1_U3101) );
  AOI22_X1 U23242 ( .A1(n20533), .A2(n20294), .B1(n10080), .B2(n20532), .ZN(
        n20291) );
  AOI22_X1 U23243 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20296), .B1(
        n20295), .B2(n20534), .ZN(n20290) );
  OAI211_X1 U23244 ( .C1(n20537), .C2(n20323), .A(n20291), .B(n20290), .ZN(
        P1_U3102) );
  AOI22_X1 U23245 ( .A1(n20539), .A2(n20294), .B1(n10080), .B2(n20538), .ZN(
        n20293) );
  AOI22_X1 U23246 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20296), .B1(
        n20295), .B2(n20540), .ZN(n20292) );
  OAI211_X1 U23247 ( .C1(n20543), .C2(n20323), .A(n20293), .B(n20292), .ZN(
        P1_U3103) );
  AOI22_X1 U23248 ( .A1(n20547), .A2(n20294), .B1(n10080), .B2(n20545), .ZN(
        n20298) );
  AOI22_X1 U23249 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20296), .B1(
        n20295), .B2(n20548), .ZN(n20297) );
  OAI211_X1 U23250 ( .C1(n20554), .C2(n20323), .A(n20298), .B(n20297), .ZN(
        P1_U3104) );
  NOR2_X1 U23251 ( .A1(n20355), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20302) );
  INV_X1 U23252 ( .A(n20302), .ZN(n20299) );
  NOR2_X1 U23253 ( .A1(n20415), .A2(n20299), .ZN(n20318) );
  AOI21_X1 U23254 ( .B1(n20356), .B2(n20416), .A(n20318), .ZN(n20300) );
  OAI22_X1 U23255 ( .A1(n20300), .A2(n20646), .B1(n20299), .B2(n12008), .ZN(
        n20319) );
  AOI22_X1 U23256 ( .A1(n20496), .A2(n20319), .B1(n20495), .B2(n20318), .ZN(
        n20305) );
  OAI211_X1 U23257 ( .C1(n20647), .C2(n20640), .A(n20503), .B(n20300), .ZN(
        n20301) );
  OAI211_X1 U23258 ( .C1(n20641), .C2(n20302), .A(n20501), .B(n20301), .ZN(
        n20320) );
  AOI22_X1 U23259 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20320), .B1(
        n20345), .B2(n20453), .ZN(n20304) );
  OAI211_X1 U23260 ( .C1(n20456), .C2(n20323), .A(n20305), .B(n20304), .ZN(
        P1_U3105) );
  AOI22_X1 U23261 ( .A1(n20509), .A2(n20319), .B1(n20508), .B2(n20318), .ZN(
        n20307) );
  AOI22_X1 U23262 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20320), .B1(
        n20345), .B2(n20457), .ZN(n20306) );
  OAI211_X1 U23263 ( .C1(n20460), .C2(n20323), .A(n20307), .B(n20306), .ZN(
        P1_U3106) );
  AOI22_X1 U23264 ( .A1(n20515), .A2(n20319), .B1(n20514), .B2(n20318), .ZN(
        n20309) );
  AOI22_X1 U23265 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20320), .B1(
        n20345), .B2(n20461), .ZN(n20308) );
  OAI211_X1 U23266 ( .C1(n20464), .C2(n20323), .A(n20309), .B(n20308), .ZN(
        P1_U3107) );
  AOI22_X1 U23267 ( .A1(n20521), .A2(n20319), .B1(n20520), .B2(n20318), .ZN(
        n20311) );
  AOI22_X1 U23268 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20320), .B1(
        n20345), .B2(n20465), .ZN(n20310) );
  OAI211_X1 U23269 ( .C1(n20468), .C2(n20323), .A(n20311), .B(n20310), .ZN(
        P1_U3108) );
  AOI22_X1 U23270 ( .A1(n20527), .A2(n20319), .B1(n20526), .B2(n20318), .ZN(
        n20313) );
  AOI22_X1 U23271 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20320), .B1(
        n20345), .B2(n20469), .ZN(n20312) );
  OAI211_X1 U23272 ( .C1(n20472), .C2(n20323), .A(n20313), .B(n20312), .ZN(
        P1_U3109) );
  AOI22_X1 U23273 ( .A1(n20533), .A2(n20319), .B1(n20532), .B2(n20318), .ZN(
        n20315) );
  AOI22_X1 U23274 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20320), .B1(
        n20345), .B2(n20473), .ZN(n20314) );
  OAI211_X1 U23275 ( .C1(n20476), .C2(n20323), .A(n20315), .B(n20314), .ZN(
        P1_U3110) );
  AOI22_X1 U23276 ( .A1(n20539), .A2(n20319), .B1(n20538), .B2(n20318), .ZN(
        n20317) );
  AOI22_X1 U23277 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20320), .B1(
        n20345), .B2(n20477), .ZN(n20316) );
  OAI211_X1 U23278 ( .C1(n20480), .C2(n20323), .A(n20317), .B(n20316), .ZN(
        P1_U3111) );
  AOI22_X1 U23279 ( .A1(n20547), .A2(n20319), .B1(n20545), .B2(n20318), .ZN(
        n20322) );
  AOI22_X1 U23280 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20320), .B1(
        n20345), .B2(n20483), .ZN(n20321) );
  OAI211_X1 U23281 ( .C1(n20488), .C2(n20323), .A(n20322), .B(n20321), .ZN(
        P1_U3112) );
  NOR2_X1 U23282 ( .A1(n20493), .A2(n20355), .ZN(n20360) );
  NAND2_X1 U23283 ( .A1(n20415), .A2(n20360), .ZN(n20325) );
  AOI22_X1 U23284 ( .A1(n20345), .A2(n20504), .B1(n20495), .B2(n20348), .ZN(
        n20334) );
  NAND2_X1 U23285 ( .A1(n20376), .A2(n20353), .ZN(n20324) );
  AOI21_X1 U23286 ( .B1(n20324), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20646), 
        .ZN(n20329) );
  NAND2_X1 U23287 ( .A1(n20356), .A2(n20447), .ZN(n20331) );
  AOI22_X1 U23288 ( .A1(n20329), .A2(n20331), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20325), .ZN(n20327) );
  OR2_X1 U23289 ( .A1(n20326), .A2(n20655), .ZN(n20443) );
  NAND2_X1 U23290 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20443), .ZN(n20449) );
  NAND3_X1 U23291 ( .A1(n20328), .A2(n20327), .A3(n20449), .ZN(n20350) );
  INV_X1 U23292 ( .A(n20329), .ZN(n20332) );
  AOI22_X1 U23293 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20350), .B1(
        n20496), .B2(n20349), .ZN(n20333) );
  OAI211_X1 U23294 ( .C1(n20507), .C2(n20376), .A(n20334), .B(n20333), .ZN(
        P1_U3113) );
  AOI22_X1 U23295 ( .A1(n20345), .A2(n20510), .B1(n20508), .B2(n20348), .ZN(
        n20336) );
  AOI22_X1 U23296 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20350), .B1(
        n20509), .B2(n20349), .ZN(n20335) );
  OAI211_X1 U23297 ( .C1(n20513), .C2(n20376), .A(n20336), .B(n20335), .ZN(
        P1_U3114) );
  AOI22_X1 U23298 ( .A1(n20379), .A2(n20461), .B1(n20514), .B2(n20348), .ZN(
        n20338) );
  AOI22_X1 U23299 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20350), .B1(
        n20515), .B2(n20349), .ZN(n20337) );
  OAI211_X1 U23300 ( .C1(n20464), .C2(n20353), .A(n20338), .B(n20337), .ZN(
        P1_U3115) );
  AOI22_X1 U23301 ( .A1(n20379), .A2(n20465), .B1(n20520), .B2(n20348), .ZN(
        n20340) );
  AOI22_X1 U23302 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20350), .B1(
        n20521), .B2(n20349), .ZN(n20339) );
  OAI211_X1 U23303 ( .C1(n20468), .C2(n20353), .A(n20340), .B(n20339), .ZN(
        P1_U3116) );
  AOI22_X1 U23304 ( .A1(n20345), .A2(n20528), .B1(n20526), .B2(n20348), .ZN(
        n20342) );
  AOI22_X1 U23305 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20350), .B1(
        n20527), .B2(n20349), .ZN(n20341) );
  OAI211_X1 U23306 ( .C1(n20531), .C2(n20376), .A(n20342), .B(n20341), .ZN(
        P1_U3117) );
  AOI22_X1 U23307 ( .A1(n20379), .A2(n20473), .B1(n20532), .B2(n20348), .ZN(
        n20344) );
  AOI22_X1 U23308 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20350), .B1(
        n20533), .B2(n20349), .ZN(n20343) );
  OAI211_X1 U23309 ( .C1(n20476), .C2(n20353), .A(n20344), .B(n20343), .ZN(
        P1_U3118) );
  AOI22_X1 U23310 ( .A1(n20345), .A2(n20540), .B1(n20538), .B2(n20348), .ZN(
        n20347) );
  AOI22_X1 U23311 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20350), .B1(
        n20539), .B2(n20349), .ZN(n20346) );
  OAI211_X1 U23312 ( .C1(n20543), .C2(n20376), .A(n20347), .B(n20346), .ZN(
        P1_U3119) );
  AOI22_X1 U23313 ( .A1(n20379), .A2(n20483), .B1(n20545), .B2(n20348), .ZN(
        n20352) );
  AOI22_X1 U23314 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20350), .B1(
        n20547), .B2(n20349), .ZN(n20351) );
  OAI211_X1 U23315 ( .C1(n20488), .C2(n20353), .A(n20352), .B(n20351), .ZN(
        P1_U3120) );
  NOR2_X1 U23316 ( .A1(n20489), .A2(n20355), .ZN(n20377) );
  AOI21_X1 U23317 ( .B1(n20356), .B2(n20490), .A(n20377), .ZN(n20358) );
  INV_X1 U23318 ( .A(n20360), .ZN(n20357) );
  OAI22_X1 U23319 ( .A1(n20358), .A2(n20646), .B1(n20357), .B2(n12008), .ZN(
        n20378) );
  AOI22_X1 U23320 ( .A1(n20496), .A2(n20378), .B1(n20495), .B2(n20377), .ZN(
        n20362) );
  OAI211_X1 U23321 ( .C1(n20647), .C2(n20499), .A(n20641), .B(n20358), .ZN(
        n20359) );
  OAI211_X1 U23322 ( .C1(n20641), .C2(n20360), .A(n20501), .B(n20359), .ZN(
        n20380) );
  AOI22_X1 U23323 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20380), .B1(
        n20379), .B2(n20504), .ZN(n20361) );
  OAI211_X1 U23324 ( .C1(n20507), .C2(n20412), .A(n20362), .B(n20361), .ZN(
        P1_U3121) );
  AOI22_X1 U23325 ( .A1(n20509), .A2(n20378), .B1(n20508), .B2(n20377), .ZN(
        n20364) );
  AOI22_X1 U23326 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20380), .B1(
        n20379), .B2(n20510), .ZN(n20363) );
  OAI211_X1 U23327 ( .C1(n20513), .C2(n20412), .A(n20364), .B(n20363), .ZN(
        P1_U3122) );
  AOI22_X1 U23328 ( .A1(n20515), .A2(n20378), .B1(n20514), .B2(n20377), .ZN(
        n20366) );
  AOI22_X1 U23329 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20380), .B1(
        n20379), .B2(n20516), .ZN(n20365) );
  OAI211_X1 U23330 ( .C1(n20519), .C2(n20412), .A(n20366), .B(n20365), .ZN(
        P1_U3123) );
  AOI22_X1 U23331 ( .A1(n20521), .A2(n20378), .B1(n20520), .B2(n20377), .ZN(
        n20368) );
  INV_X1 U23332 ( .A(n20412), .ZN(n20373) );
  AOI22_X1 U23333 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20380), .B1(
        n20373), .B2(n20465), .ZN(n20367) );
  OAI211_X1 U23334 ( .C1(n20468), .C2(n20376), .A(n20368), .B(n20367), .ZN(
        P1_U3124) );
  AOI22_X1 U23335 ( .A1(n20527), .A2(n20378), .B1(n20526), .B2(n20377), .ZN(
        n20370) );
  AOI22_X1 U23336 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20380), .B1(
        n20379), .B2(n20528), .ZN(n20369) );
  OAI211_X1 U23337 ( .C1(n20531), .C2(n20412), .A(n20370), .B(n20369), .ZN(
        P1_U3125) );
  AOI22_X1 U23338 ( .A1(n20533), .A2(n20378), .B1(n20532), .B2(n20377), .ZN(
        n20372) );
  AOI22_X1 U23339 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20380), .B1(
        n20373), .B2(n20473), .ZN(n20371) );
  OAI211_X1 U23340 ( .C1(n20476), .C2(n20376), .A(n20372), .B(n20371), .ZN(
        P1_U3126) );
  AOI22_X1 U23341 ( .A1(n20539), .A2(n20378), .B1(n20538), .B2(n20377), .ZN(
        n20375) );
  AOI22_X1 U23342 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20380), .B1(
        n20373), .B2(n20477), .ZN(n20374) );
  OAI211_X1 U23343 ( .C1(n20480), .C2(n20376), .A(n20375), .B(n20374), .ZN(
        P1_U3127) );
  AOI22_X1 U23344 ( .A1(n20547), .A2(n20378), .B1(n20545), .B2(n20377), .ZN(
        n20382) );
  AOI22_X1 U23345 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20380), .B1(
        n20379), .B2(n20548), .ZN(n20381) );
  OAI211_X1 U23346 ( .C1(n20554), .C2(n20412), .A(n20382), .B(n20381), .ZN(
        P1_U3128) );
  OR2_X1 U23347 ( .A1(n20498), .A2(n13601), .ZN(n20648) );
  NAND2_X1 U23348 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20492) );
  AOI22_X1 U23349 ( .A1(n20438), .A2(n20453), .B1(n20495), .B2(n9738), .ZN(
        n20395) );
  NAND2_X1 U23350 ( .A1(n20385), .A2(n20412), .ZN(n20386) );
  AOI21_X1 U23351 ( .B1(n20386), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20646), 
        .ZN(n20390) );
  NAND2_X1 U23352 ( .A1(n20491), .A2(n13646), .ZN(n20392) );
  AOI22_X1 U23353 ( .A1(n20390), .A2(n20392), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20391), .ZN(n20388) );
  OAI211_X1 U23354 ( .C1(n9738), .C2(n20389), .A(n20450), .B(n20388), .ZN(
        n20409) );
  INV_X1 U23355 ( .A(n20390), .ZN(n20393) );
  AOI22_X1 U23356 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20409), .B1(
        n20496), .B2(n20408), .ZN(n20394) );
  OAI211_X1 U23357 ( .C1(n20456), .C2(n20412), .A(n20395), .B(n20394), .ZN(
        P1_U3129) );
  AOI22_X1 U23358 ( .A1(n20438), .A2(n20457), .B1(n20508), .B2(n9738), .ZN(
        n20397) );
  AOI22_X1 U23359 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20409), .B1(
        n20509), .B2(n20408), .ZN(n20396) );
  OAI211_X1 U23360 ( .C1(n20460), .C2(n20412), .A(n20397), .B(n20396), .ZN(
        P1_U3130) );
  AOI22_X1 U23361 ( .A1(n20438), .A2(n20461), .B1(n20514), .B2(n9738), .ZN(
        n20399) );
  AOI22_X1 U23362 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20409), .B1(
        n20515), .B2(n20408), .ZN(n20398) );
  OAI211_X1 U23363 ( .C1(n20464), .C2(n20412), .A(n20399), .B(n20398), .ZN(
        P1_U3131) );
  AOI22_X1 U23364 ( .A1(n20438), .A2(n20465), .B1(n20520), .B2(n9738), .ZN(
        n20401) );
  AOI22_X1 U23365 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20409), .B1(
        n20521), .B2(n20408), .ZN(n20400) );
  OAI211_X1 U23366 ( .C1(n20468), .C2(n20412), .A(n20401), .B(n20400), .ZN(
        P1_U3132) );
  AOI22_X1 U23367 ( .A1(n20438), .A2(n20469), .B1(n20526), .B2(n9738), .ZN(
        n20403) );
  AOI22_X1 U23368 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20409), .B1(
        n20527), .B2(n20408), .ZN(n20402) );
  OAI211_X1 U23369 ( .C1(n20472), .C2(n20412), .A(n20403), .B(n20402), .ZN(
        P1_U3133) );
  AOI22_X1 U23370 ( .A1(n20438), .A2(n20473), .B1(n20532), .B2(n9738), .ZN(
        n20405) );
  AOI22_X1 U23371 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20409), .B1(
        n20533), .B2(n20408), .ZN(n20404) );
  OAI211_X1 U23372 ( .C1(n20476), .C2(n20412), .A(n20405), .B(n20404), .ZN(
        P1_U3134) );
  AOI22_X1 U23373 ( .A1(n20438), .A2(n20477), .B1(n20538), .B2(n9738), .ZN(
        n20407) );
  AOI22_X1 U23374 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20409), .B1(
        n20539), .B2(n20408), .ZN(n20406) );
  OAI211_X1 U23375 ( .C1(n20480), .C2(n20412), .A(n20407), .B(n20406), .ZN(
        P1_U3135) );
  AOI22_X1 U23376 ( .A1(n20438), .A2(n20483), .B1(n20545), .B2(n9738), .ZN(
        n20411) );
  AOI22_X1 U23377 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20409), .B1(
        n20547), .B2(n20408), .ZN(n20410) );
  OAI211_X1 U23378 ( .C1(n20488), .C2(n20412), .A(n20411), .B(n20410), .ZN(
        P1_U3136) );
  INV_X1 U23379 ( .A(n20498), .ZN(n20414) );
  NOR3_X2 U23380 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20415), .A3(
        n20492), .ZN(n20436) );
  AOI21_X1 U23381 ( .B1(n20491), .B2(n20416), .A(n20436), .ZN(n20419) );
  NOR2_X1 U23382 ( .A1(n20492), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20421) );
  INV_X1 U23383 ( .A(n20421), .ZN(n20418) );
  OAI22_X1 U23384 ( .A1(n20419), .A2(n20646), .B1(n20418), .B2(n20417), .ZN(
        n20437) );
  AOI22_X1 U23385 ( .A1(n20496), .A2(n20437), .B1(n20495), .B2(n20436), .ZN(
        n20423) );
  OAI211_X1 U23386 ( .C1(n20498), .C2(n20640), .A(n20503), .B(n20419), .ZN(
        n20420) );
  OAI211_X1 U23387 ( .C1(n20641), .C2(n20421), .A(n20501), .B(n20420), .ZN(
        n20439) );
  AOI22_X1 U23388 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20439), .B1(
        n20438), .B2(n20504), .ZN(n20422) );
  OAI211_X1 U23389 ( .C1(n20507), .C2(n20487), .A(n20423), .B(n20422), .ZN(
        P1_U3137) );
  AOI22_X1 U23390 ( .A1(n20509), .A2(n20437), .B1(n20508), .B2(n20436), .ZN(
        n20425) );
  AOI22_X1 U23391 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20439), .B1(
        n20438), .B2(n20510), .ZN(n20424) );
  OAI211_X1 U23392 ( .C1(n20513), .C2(n20487), .A(n20425), .B(n20424), .ZN(
        P1_U3138) );
  AOI22_X1 U23393 ( .A1(n20515), .A2(n20437), .B1(n20514), .B2(n20436), .ZN(
        n20427) );
  AOI22_X1 U23394 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20439), .B1(
        n20438), .B2(n20516), .ZN(n20426) );
  OAI211_X1 U23395 ( .C1(n20519), .C2(n20487), .A(n20427), .B(n20426), .ZN(
        P1_U3139) );
  AOI22_X1 U23396 ( .A1(n20521), .A2(n20437), .B1(n20520), .B2(n20436), .ZN(
        n20429) );
  AOI22_X1 U23397 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20439), .B1(
        n20438), .B2(n20522), .ZN(n20428) );
  OAI211_X1 U23398 ( .C1(n20525), .C2(n20487), .A(n20429), .B(n20428), .ZN(
        P1_U3140) );
  AOI22_X1 U23399 ( .A1(n20527), .A2(n20437), .B1(n20526), .B2(n20436), .ZN(
        n20431) );
  AOI22_X1 U23400 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20439), .B1(
        n20438), .B2(n20528), .ZN(n20430) );
  OAI211_X1 U23401 ( .C1(n20531), .C2(n20487), .A(n20431), .B(n20430), .ZN(
        P1_U3141) );
  AOI22_X1 U23402 ( .A1(n20533), .A2(n20437), .B1(n20532), .B2(n20436), .ZN(
        n20433) );
  AOI22_X1 U23403 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20439), .B1(
        n20438), .B2(n20534), .ZN(n20432) );
  OAI211_X1 U23404 ( .C1(n20537), .C2(n20487), .A(n20433), .B(n20432), .ZN(
        P1_U3142) );
  AOI22_X1 U23405 ( .A1(n20539), .A2(n20437), .B1(n20538), .B2(n20436), .ZN(
        n20435) );
  AOI22_X1 U23406 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20439), .B1(
        n20438), .B2(n20540), .ZN(n20434) );
  OAI211_X1 U23407 ( .C1(n20543), .C2(n20487), .A(n20435), .B(n20434), .ZN(
        P1_U3143) );
  AOI22_X1 U23408 ( .A1(n20547), .A2(n20437), .B1(n20545), .B2(n20436), .ZN(
        n20441) );
  AOI22_X1 U23409 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20439), .B1(
        n20438), .B2(n20548), .ZN(n20440) );
  OAI211_X1 U23410 ( .C1(n20554), .C2(n20487), .A(n20441), .B(n20440), .ZN(
        P1_U3144) );
  NAND3_X1 U23411 ( .A1(n20491), .A2(n20447), .A3(n20641), .ZN(n20442) );
  OAI21_X1 U23412 ( .B1(n20444), .B2(n20443), .A(n20442), .ZN(n20482) );
  NOR3_X2 U23413 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20493), .A3(
        n20492), .ZN(n20481) );
  AOI22_X1 U23414 ( .A1(n20496), .A2(n20482), .B1(n20495), .B2(n20481), .ZN(
        n20455) );
  AOI21_X1 U23415 ( .B1(n20487), .B2(n20452), .A(n20640), .ZN(n20446) );
  AOI21_X1 U23416 ( .B1(n20491), .B2(n20447), .A(n20446), .ZN(n20448) );
  NOR2_X1 U23417 ( .A1(n20448), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20451) );
  AOI22_X1 U23418 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20484), .B1(
        n20549), .B2(n20453), .ZN(n20454) );
  OAI211_X1 U23419 ( .C1(n20456), .C2(n20487), .A(n20455), .B(n20454), .ZN(
        P1_U3145) );
  AOI22_X1 U23420 ( .A1(n20509), .A2(n20482), .B1(n20508), .B2(n20481), .ZN(
        n20459) );
  AOI22_X1 U23421 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20484), .B1(
        n20549), .B2(n20457), .ZN(n20458) );
  OAI211_X1 U23422 ( .C1(n20460), .C2(n20487), .A(n20459), .B(n20458), .ZN(
        P1_U3146) );
  AOI22_X1 U23423 ( .A1(n20515), .A2(n20482), .B1(n20514), .B2(n20481), .ZN(
        n20463) );
  AOI22_X1 U23424 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20484), .B1(
        n20549), .B2(n20461), .ZN(n20462) );
  OAI211_X1 U23425 ( .C1(n20464), .C2(n20487), .A(n20463), .B(n20462), .ZN(
        P1_U3147) );
  AOI22_X1 U23426 ( .A1(n20521), .A2(n20482), .B1(n20520), .B2(n20481), .ZN(
        n20467) );
  AOI22_X1 U23427 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20484), .B1(
        n20549), .B2(n20465), .ZN(n20466) );
  OAI211_X1 U23428 ( .C1(n20468), .C2(n20487), .A(n20467), .B(n20466), .ZN(
        P1_U3148) );
  AOI22_X1 U23429 ( .A1(n20527), .A2(n20482), .B1(n20526), .B2(n20481), .ZN(
        n20471) );
  AOI22_X1 U23430 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20484), .B1(
        n20549), .B2(n20469), .ZN(n20470) );
  OAI211_X1 U23431 ( .C1(n20472), .C2(n20487), .A(n20471), .B(n20470), .ZN(
        P1_U3149) );
  AOI22_X1 U23432 ( .A1(n20533), .A2(n20482), .B1(n20532), .B2(n20481), .ZN(
        n20475) );
  AOI22_X1 U23433 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20484), .B1(
        n20549), .B2(n20473), .ZN(n20474) );
  OAI211_X1 U23434 ( .C1(n20476), .C2(n20487), .A(n20475), .B(n20474), .ZN(
        P1_U3150) );
  AOI22_X1 U23435 ( .A1(n20539), .A2(n20482), .B1(n20538), .B2(n20481), .ZN(
        n20479) );
  AOI22_X1 U23436 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20484), .B1(
        n20549), .B2(n20477), .ZN(n20478) );
  OAI211_X1 U23437 ( .C1(n20480), .C2(n20487), .A(n20479), .B(n20478), .ZN(
        P1_U3151) );
  AOI22_X1 U23438 ( .A1(n20547), .A2(n20482), .B1(n20545), .B2(n20481), .ZN(
        n20486) );
  AOI22_X1 U23439 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20484), .B1(
        n20549), .B2(n20483), .ZN(n20485) );
  OAI211_X1 U23440 ( .C1(n20488), .C2(n20487), .A(n20486), .B(n20485), .ZN(
        P1_U3152) );
  NOR2_X1 U23441 ( .A1(n20489), .A2(n20492), .ZN(n20544) );
  AOI21_X1 U23442 ( .B1(n20491), .B2(n20490), .A(n20544), .ZN(n20497) );
  NOR2_X1 U23443 ( .A1(n20493), .A2(n20492), .ZN(n20502) );
  INV_X1 U23444 ( .A(n20502), .ZN(n20494) );
  OAI22_X1 U23445 ( .A1(n20497), .A2(n20646), .B1(n20494), .B2(n12008), .ZN(
        n20546) );
  AOI22_X1 U23446 ( .A1(n20496), .A2(n20546), .B1(n20495), .B2(n20544), .ZN(
        n20506) );
  OAI211_X1 U23447 ( .C1(n20499), .C2(n20498), .A(n20641), .B(n20497), .ZN(
        n20500) );
  OAI211_X1 U23448 ( .C1(n20503), .C2(n20502), .A(n20501), .B(n20500), .ZN(
        n20550) );
  AOI22_X1 U23449 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20550), .B1(
        n20549), .B2(n20504), .ZN(n20505) );
  OAI211_X1 U23450 ( .C1(n20507), .C2(n20553), .A(n20506), .B(n20505), .ZN(
        P1_U3153) );
  AOI22_X1 U23451 ( .A1(n20509), .A2(n20546), .B1(n20508), .B2(n20544), .ZN(
        n20512) );
  AOI22_X1 U23452 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20550), .B1(
        n20549), .B2(n20510), .ZN(n20511) );
  OAI211_X1 U23453 ( .C1(n20513), .C2(n20553), .A(n20512), .B(n20511), .ZN(
        P1_U3154) );
  AOI22_X1 U23454 ( .A1(n20515), .A2(n20546), .B1(n20514), .B2(n20544), .ZN(
        n20518) );
  AOI22_X1 U23455 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20550), .B1(
        n20549), .B2(n20516), .ZN(n20517) );
  OAI211_X1 U23456 ( .C1(n20519), .C2(n20553), .A(n20518), .B(n20517), .ZN(
        P1_U3155) );
  AOI22_X1 U23457 ( .A1(n20521), .A2(n20546), .B1(n20520), .B2(n20544), .ZN(
        n20524) );
  AOI22_X1 U23458 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20550), .B1(
        n20549), .B2(n20522), .ZN(n20523) );
  OAI211_X1 U23459 ( .C1(n20525), .C2(n20553), .A(n20524), .B(n20523), .ZN(
        P1_U3156) );
  AOI22_X1 U23460 ( .A1(n20527), .A2(n20546), .B1(n20526), .B2(n20544), .ZN(
        n20530) );
  AOI22_X1 U23461 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20550), .B1(
        n20549), .B2(n20528), .ZN(n20529) );
  OAI211_X1 U23462 ( .C1(n20531), .C2(n20553), .A(n20530), .B(n20529), .ZN(
        P1_U3157) );
  AOI22_X1 U23463 ( .A1(n20533), .A2(n20546), .B1(n20532), .B2(n20544), .ZN(
        n20536) );
  AOI22_X1 U23464 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20550), .B1(
        n20549), .B2(n20534), .ZN(n20535) );
  OAI211_X1 U23465 ( .C1(n20537), .C2(n20553), .A(n20536), .B(n20535), .ZN(
        P1_U3158) );
  AOI22_X1 U23466 ( .A1(n20539), .A2(n20546), .B1(n20538), .B2(n20544), .ZN(
        n20542) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20550), .B1(
        n20549), .B2(n20540), .ZN(n20541) );
  OAI211_X1 U23468 ( .C1(n20543), .C2(n20553), .A(n20542), .B(n20541), .ZN(
        P1_U3159) );
  AOI22_X1 U23469 ( .A1(n20547), .A2(n20546), .B1(n20545), .B2(n20544), .ZN(
        n20552) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20550), .B1(
        n20549), .B2(n20548), .ZN(n20551) );
  OAI211_X1 U23471 ( .C1(n20554), .C2(n20553), .A(n20552), .B(n20551), .ZN(
        P1_U3160) );
  NOR2_X1 U23472 ( .A1(n20556), .A2(n20555), .ZN(n20559) );
  INV_X1 U23473 ( .A(n20557), .ZN(n20558) );
  OAI21_X1 U23474 ( .B1(n20559), .B2(n20417), .A(n20558), .ZN(P1_U3163) );
  AND2_X1 U23475 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20560), .ZN(
        P1_U3164) );
  AND2_X1 U23476 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20560), .ZN(
        P1_U3165) );
  AND2_X1 U23477 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20560), .ZN(
        P1_U3166) );
  AND2_X1 U23478 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20560), .ZN(
        P1_U3167) );
  AND2_X1 U23479 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20560), .ZN(
        P1_U3168) );
  AND2_X1 U23480 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20560), .ZN(
        P1_U3169) );
  AND2_X1 U23481 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20560), .ZN(
        P1_U3170) );
  AND2_X1 U23482 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20560), .ZN(
        P1_U3171) );
  AND2_X1 U23483 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20560), .ZN(
        P1_U3172) );
  AND2_X1 U23484 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20560), .ZN(
        P1_U3173) );
  AND2_X1 U23485 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20560), .ZN(
        P1_U3174) );
  AND2_X1 U23486 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20560), .ZN(
        P1_U3175) );
  AND2_X1 U23487 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20560), .ZN(
        P1_U3176) );
  AND2_X1 U23488 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20560), .ZN(
        P1_U3177) );
  AND2_X1 U23489 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20560), .ZN(
        P1_U3178) );
  AND2_X1 U23490 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20560), .ZN(
        P1_U3179) );
  AND2_X1 U23491 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20560), .ZN(
        P1_U3180) );
  AND2_X1 U23492 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20560), .ZN(
        P1_U3181) );
  AND2_X1 U23493 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20560), .ZN(
        P1_U3182) );
  AND2_X1 U23494 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20560), .ZN(
        P1_U3183) );
  AND2_X1 U23495 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20560), .ZN(
        P1_U3184) );
  AND2_X1 U23496 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20560), .ZN(
        P1_U3185) );
  AND2_X1 U23497 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20560), .ZN(P1_U3186) );
  AND2_X1 U23498 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20560), .ZN(P1_U3187) );
  AND2_X1 U23499 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20560), .ZN(P1_U3188) );
  AND2_X1 U23500 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20560), .ZN(P1_U3189) );
  INV_X1 U23501 ( .A(P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n20678) );
  NOR2_X1 U23502 ( .A1(n20632), .A2(n20678), .ZN(P1_U3190) );
  AND2_X1 U23503 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20560), .ZN(P1_U3191) );
  AND2_X1 U23504 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20560), .ZN(P1_U3192) );
  AND2_X1 U23505 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20560), .ZN(P1_U3193) );
  AOI21_X1 U23506 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20567), .A(n20564), 
        .ZN(n20570) );
  NOR2_X1 U23507 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20562) );
  OAI21_X1 U23508 ( .B1(n20562), .B2(n20561), .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20563) );
  AOI21_X1 U23509 ( .B1(NA), .B2(n20564), .A(n20563), .ZN(n20565) );
  OAI22_X1 U23510 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20570), .B1(n20666), 
        .B2(n20565), .ZN(P1_U3194) );
  NAND4_X1 U23511 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20567), .A3(
        P1_REQUESTPENDING_REG_SCAN_IN), .A4(n20566), .ZN(n20574) );
  NAND2_X1 U23512 ( .A1(n20567), .A2(n20566), .ZN(n20568) );
  OAI221_X1 U23513 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(
        P1_STATE_REG_1__SCAN_IN), .C1(P1_REQUESTPENDING_REG_SCAN_IN), .C2(
        n20568), .A(n20575), .ZN(n20569) );
  NAND3_X1 U23514 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(HOLD), .A3(n20569), .ZN(
        n20573) );
  AOI211_X1 U23515 ( .C1(n11362), .C2(NA), .A(n20575), .B(n20570), .ZN(n20571)
         );
  INV_X1 U23516 ( .A(n20571), .ZN(n20572) );
  OAI211_X1 U23517 ( .C1(n11362), .C2(n20574), .A(n20573), .B(n20572), .ZN(
        P1_U3196) );
  OR2_X1 U23518 ( .A1(n20664), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20623) );
  AOI222_X1 U23519 ( .A1(n20617), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20676), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20621), .ZN(n20576) );
  INV_X1 U23520 ( .A(n20576), .ZN(P1_U3197) );
  AOI22_X1 U23521 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20676), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n20617), .ZN(n20577) );
  OAI21_X1 U23522 ( .B1(n20578), .B2(n20619), .A(n20577), .ZN(P1_U3198) );
  AOI222_X1 U23523 ( .A1(n20621), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n20664), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20617), .ZN(n20579) );
  INV_X1 U23524 ( .A(n20579), .ZN(P1_U3199) );
  AOI222_X1 U23525 ( .A1(n20617), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20676), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20621), .ZN(n20580) );
  INV_X1 U23526 ( .A(n20580), .ZN(P1_U3200) );
  AOI222_X1 U23527 ( .A1(n20621), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20676), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20617), .ZN(n20581) );
  INV_X1 U23528 ( .A(n20581), .ZN(P1_U3201) );
  AOI222_X1 U23529 ( .A1(n20621), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20664), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20617), .ZN(n20582) );
  INV_X1 U23530 ( .A(n20582), .ZN(P1_U3202) );
  AOI222_X1 U23531 ( .A1(n20621), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20676), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20617), .ZN(n20583) );
  INV_X1 U23532 ( .A(n20583), .ZN(P1_U3203) );
  AOI222_X1 U23533 ( .A1(n20621), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20664), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n20617), .ZN(n20584) );
  INV_X1 U23534 ( .A(n20584), .ZN(P1_U3204) );
  AOI22_X1 U23535 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(n20676), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n20617), .ZN(n20585) );
  OAI21_X1 U23536 ( .B1(n20586), .B2(n20619), .A(n20585), .ZN(P1_U3205) );
  AOI22_X1 U23537 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n20676), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n20621), .ZN(n20587) );
  OAI21_X1 U23538 ( .B1(n20588), .B2(n20623), .A(n20587), .ZN(P1_U3206) );
  AOI222_X1 U23539 ( .A1(n20621), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20664), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20617), .ZN(n20589) );
  INV_X1 U23540 ( .A(n20589), .ZN(P1_U3207) );
  AOI222_X1 U23541 ( .A1(n20621), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20664), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20617), .ZN(n20590) );
  INV_X1 U23542 ( .A(n20590), .ZN(P1_U3208) );
  AOI22_X1 U23543 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20676), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20617), .ZN(n20591) );
  OAI21_X1 U23544 ( .B1(n20592), .B2(n20619), .A(n20591), .ZN(P1_U3209) );
  AOI22_X1 U23545 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20676), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20621), .ZN(n20593) );
  OAI21_X1 U23546 ( .B1(n20594), .B2(n20623), .A(n20593), .ZN(P1_U3210) );
  AOI222_X1 U23547 ( .A1(n20621), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20664), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20617), .ZN(n20595) );
  INV_X1 U23548 ( .A(n20595), .ZN(P1_U3211) );
  AOI22_X1 U23549 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20676), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20617), .ZN(n20596) );
  OAI21_X1 U23550 ( .B1(n20597), .B2(n20619), .A(n20596), .ZN(P1_U3212) );
  AOI22_X1 U23551 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20676), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20621), .ZN(n20598) );
  OAI21_X1 U23552 ( .B1(n20599), .B2(n20623), .A(n20598), .ZN(P1_U3213) );
  AOI222_X1 U23553 ( .A1(n20621), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20676), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20617), .ZN(n20600) );
  INV_X1 U23554 ( .A(n20600), .ZN(P1_U3214) );
  AOI22_X1 U23555 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20676), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20617), .ZN(n20601) );
  OAI21_X1 U23556 ( .B1(n20602), .B2(n20619), .A(n20601), .ZN(P1_U3215) );
  AOI22_X1 U23557 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20676), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20621), .ZN(n20603) );
  OAI21_X1 U23558 ( .B1(n20604), .B2(n20623), .A(n20603), .ZN(P1_U3216) );
  AOI222_X1 U23559 ( .A1(n20621), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20676), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20617), .ZN(n20605) );
  INV_X1 U23560 ( .A(n20605), .ZN(P1_U3217) );
  AOI222_X1 U23561 ( .A1(n20621), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20664), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20617), .ZN(n20606) );
  INV_X1 U23562 ( .A(n20606), .ZN(P1_U3218) );
  AOI22_X1 U23563 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n20617), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20664), .ZN(n20607) );
  OAI21_X1 U23564 ( .B1(n20608), .B2(n20619), .A(n20607), .ZN(P1_U3219) );
  AOI22_X1 U23565 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n20621), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20664), .ZN(n20609) );
  OAI21_X1 U23566 ( .B1(n20610), .B2(n20623), .A(n20609), .ZN(P1_U3220) );
  AOI222_X1 U23567 ( .A1(n20621), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20676), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20617), .ZN(n20611) );
  INV_X1 U23568 ( .A(n20611), .ZN(P1_U3221) );
  INV_X1 U23569 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20613) );
  AOI22_X1 U23570 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n20617), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20664), .ZN(n20612) );
  OAI21_X1 U23571 ( .B1(n20613), .B2(n20619), .A(n20612), .ZN(P1_U3222) );
  AOI22_X1 U23572 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n20621), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20664), .ZN(n20614) );
  OAI21_X1 U23573 ( .B1(n20615), .B2(n20623), .A(n20614), .ZN(P1_U3223) );
  AOI222_X1 U23574 ( .A1(n20621), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20664), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20617), .ZN(n20616) );
  INV_X1 U23575 ( .A(n20616), .ZN(P1_U3224) );
  AOI22_X1 U23576 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20617), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20664), .ZN(n20618) );
  OAI21_X1 U23577 ( .B1(n20620), .B2(n20619), .A(n20618), .ZN(P1_U3225) );
  AOI22_X1 U23578 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20621), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20664), .ZN(n20622) );
  OAI21_X1 U23579 ( .B1(n20624), .B2(n20623), .A(n20622), .ZN(P1_U3226) );
  OAI22_X1 U23580 ( .A1(n20664), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20666), .ZN(n20625) );
  INV_X1 U23581 ( .A(n20625), .ZN(P1_U3458) );
  OAI22_X1 U23582 ( .A1(n20676), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20666), .ZN(n20626) );
  INV_X1 U23583 ( .A(n20626), .ZN(P1_U3459) );
  OAI22_X1 U23584 ( .A1(n20664), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20666), .ZN(n20627) );
  INV_X1 U23585 ( .A(n20627), .ZN(P1_U3460) );
  OAI22_X1 U23586 ( .A1(n20676), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20666), .ZN(n20628) );
  INV_X1 U23587 ( .A(n20628), .ZN(P1_U3461) );
  OAI21_X1 U23588 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20632), .A(n20630), 
        .ZN(n20629) );
  INV_X1 U23589 ( .A(n20629), .ZN(P1_U3464) );
  OAI21_X1 U23590 ( .B1(n20632), .B2(n20631), .A(n20630), .ZN(P1_U3465) );
  OAI22_X1 U23591 ( .A1(n20636), .A2(n20635), .B1(n20634), .B2(n20633), .ZN(
        n20638) );
  MUX2_X1 U23592 ( .A(n20638), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n20637), .Z(P1_U3469) );
  INV_X1 U23593 ( .A(n20653), .ZN(n20656) );
  INV_X1 U23594 ( .A(n20639), .ZN(n20652) );
  NAND3_X1 U23595 ( .A1(n20642), .A2(n20641), .A3(n20640), .ZN(n20643) );
  OAI21_X1 U23596 ( .B1(n20645), .B2(n20644), .A(n20643), .ZN(n20650) );
  AOI21_X1 U23597 ( .B1(n20648), .B2(n20647), .A(n20646), .ZN(n20649) );
  AOI211_X1 U23598 ( .C1(n20652), .C2(n20651), .A(n20650), .B(n20649), .ZN(
        n20654) );
  AOI22_X1 U23599 ( .A1(n20656), .A2(n20655), .B1(n20654), .B2(n20653), .ZN(
        P1_U3475) );
  AOI211_X1 U23600 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_REIP_REG_1__SCAN_IN), .B(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20657) );
  AOI21_X1 U23601 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20657), .ZN(n20659) );
  INV_X1 U23602 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20658) );
  AOI22_X1 U23603 ( .A1(n20663), .A2(n20659), .B1(n20658), .B2(n20660), .ZN(
        P1_U3481) );
  NOR2_X1 U23604 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n20662) );
  INV_X1 U23605 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20661) );
  AOI22_X1 U23606 ( .A1(n20663), .A2(n20662), .B1(n20661), .B2(n20660), .ZN(
        P1_U3482) );
  AOI22_X1 U23607 ( .A1(n20666), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20665), 
        .B2(n20664), .ZN(P1_U3483) );
  AOI211_X1 U23608 ( .C1(n19930), .C2(n20669), .A(n20668), .B(n20667), .ZN(
        n20675) );
  OAI211_X1 U23609 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n11399), .A(n20670), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20672) );
  AOI21_X1 U23610 ( .B1(n20672), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n20671), 
        .ZN(n20674) );
  NAND2_X1 U23611 ( .A1(n20675), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20673) );
  OAI21_X1 U23612 ( .B1(n20675), .B2(n20674), .A(n20673), .ZN(P1_U3485) );
  MUX2_X1 U23613 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n20676), .Z(P1_U3486) );
  AOI22_X1 U23614 ( .A1(n20679), .A2(keyinput0), .B1(keyinput58), .B2(n20678), 
        .ZN(n20677) );
  OAI221_X1 U23615 ( .B1(n20679), .B2(keyinput0), .C1(n20678), .C2(keyinput58), 
        .A(n20677), .ZN(n20684) );
  XNOR2_X1 U23616 ( .A(n20680), .B(keyinput2), .ZN(n20683) );
  XOR2_X1 U23617 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B(keyinput63), .Z(
        n20682) );
  XNOR2_X1 U23618 ( .A(n9620), .B(keyinput61), .ZN(n20681) );
  OR4_X1 U23619 ( .A1(n20684), .A2(n20683), .A3(n20682), .A4(n20681), .ZN(
        n20691) );
  AOI22_X1 U23620 ( .A1(n20687), .A2(keyinput8), .B1(keyinput54), .B2(n20686), 
        .ZN(n20685) );
  OAI221_X1 U23621 ( .B1(n20687), .B2(keyinput8), .C1(n20686), .C2(keyinput54), 
        .A(n20685), .ZN(n20690) );
  XNOR2_X1 U23622 ( .A(n20688), .B(keyinput45), .ZN(n20689) );
  NOR3_X1 U23623 ( .A1(n20691), .A2(n20690), .A3(n20689), .ZN(n20736) );
  AOI22_X1 U23624 ( .A1(n20827), .A2(keyinput46), .B1(keyinput41), .B2(n20824), 
        .ZN(n20692) );
  OAI221_X1 U23625 ( .B1(n20827), .B2(keyinput46), .C1(n20824), .C2(keyinput41), .A(n20692), .ZN(n20701) );
  AOI22_X1 U23626 ( .A1(n11169), .A2(keyinput51), .B1(keyinput17), .B2(n20823), 
        .ZN(n20693) );
  OAI221_X1 U23627 ( .B1(n11169), .B2(keyinput51), .C1(n20823), .C2(keyinput17), .A(n20693), .ZN(n20700) );
  AOI22_X1 U23628 ( .A1(n20825), .A2(keyinput42), .B1(keyinput47), .B2(n20695), 
        .ZN(n20694) );
  OAI221_X1 U23629 ( .B1(n20825), .B2(keyinput42), .C1(n20695), .C2(keyinput47), .A(n20694), .ZN(n20699) );
  AOI22_X1 U23630 ( .A1(n20697), .A2(keyinput48), .B1(n12395), .B2(keyinput27), 
        .ZN(n20696) );
  OAI221_X1 U23631 ( .B1(n20697), .B2(keyinput48), .C1(n12395), .C2(keyinput27), .A(n20696), .ZN(n20698) );
  NOR4_X1 U23632 ( .A1(n20701), .A2(n20700), .A3(n20699), .A4(n20698), .ZN(
        n20735) );
  INV_X1 U23633 ( .A(DATAI_29_), .ZN(n20703) );
  AOI22_X1 U23634 ( .A1(n20704), .A2(keyinput35), .B1(n20703), .B2(keyinput19), 
        .ZN(n20702) );
  OAI221_X1 U23635 ( .B1(n20704), .B2(keyinput35), .C1(n20703), .C2(keyinput19), .A(n20702), .ZN(n20717) );
  INV_X1 U23636 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n20706) );
  AOI22_X1 U23637 ( .A1(n20707), .A2(keyinput59), .B1(n20706), .B2(keyinput7), 
        .ZN(n20705) );
  OAI221_X1 U23638 ( .B1(n20707), .B2(keyinput59), .C1(n20706), .C2(keyinput7), 
        .A(n20705), .ZN(n20716) );
  AOI22_X1 U23639 ( .A1(n20710), .A2(keyinput44), .B1(n20709), .B2(keyinput34), 
        .ZN(n20708) );
  OAI221_X1 U23640 ( .B1(n20710), .B2(keyinput44), .C1(n20709), .C2(keyinput34), .A(n20708), .ZN(n20715) );
  AOI22_X1 U23641 ( .A1(n20713), .A2(keyinput21), .B1(keyinput23), .B2(n20712), 
        .ZN(n20711) );
  OAI221_X1 U23642 ( .B1(n20713), .B2(keyinput21), .C1(n20712), .C2(keyinput23), .A(n20711), .ZN(n20714) );
  NOR4_X1 U23643 ( .A1(n20717), .A2(n20716), .A3(n20715), .A4(n20714), .ZN(
        n20734) );
  AOI22_X1 U23644 ( .A1(n20720), .A2(keyinput40), .B1(keyinput43), .B2(n20719), 
        .ZN(n20718) );
  OAI221_X1 U23645 ( .B1(n20720), .B2(keyinput40), .C1(n20719), .C2(keyinput43), .A(n20718), .ZN(n20732) );
  INV_X1 U23646 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n20723) );
  INV_X1 U23647 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n20722) );
  AOI22_X1 U23648 ( .A1(n20723), .A2(keyinput5), .B1(n20722), .B2(keyinput6), 
        .ZN(n20721) );
  OAI221_X1 U23649 ( .B1(n20723), .B2(keyinput5), .C1(n20722), .C2(keyinput6), 
        .A(n20721), .ZN(n20731) );
  AOI22_X1 U23650 ( .A1(n20726), .A2(keyinput14), .B1(n20725), .B2(keyinput13), 
        .ZN(n20724) );
  OAI221_X1 U23651 ( .B1(n20726), .B2(keyinput14), .C1(n20725), .C2(keyinput13), .A(n20724), .ZN(n20730) );
  AOI22_X1 U23652 ( .A1(n20728), .A2(keyinput32), .B1(n13655), .B2(keyinput20), 
        .ZN(n20727) );
  OAI221_X1 U23653 ( .B1(n20728), .B2(keyinput32), .C1(n13655), .C2(keyinput20), .A(n20727), .ZN(n20729) );
  NOR4_X1 U23654 ( .A1(n20732), .A2(n20731), .A3(n20730), .A4(n20729), .ZN(
        n20733) );
  NAND4_X1 U23655 ( .A1(n20736), .A2(n20735), .A3(n20734), .A4(n20733), .ZN(
        n20802) );
  AOI22_X1 U23656 ( .A1(n20739), .A2(keyinput50), .B1(keyinput60), .B2(n20738), 
        .ZN(n20737) );
  OAI221_X1 U23657 ( .B1(n20739), .B2(keyinput50), .C1(n20738), .C2(keyinput60), .A(n20737), .ZN(n20752) );
  INV_X1 U23658 ( .A(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n20741) );
  AOI22_X1 U23659 ( .A1(n20742), .A2(keyinput37), .B1(keyinput29), .B2(n20741), 
        .ZN(n20740) );
  OAI221_X1 U23660 ( .B1(n20742), .B2(keyinput37), .C1(n20741), .C2(keyinput29), .A(n20740), .ZN(n20751) );
  INV_X1 U23661 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n20745) );
  AOI22_X1 U23662 ( .A1(n20745), .A2(keyinput53), .B1(keyinput22), .B2(n20744), 
        .ZN(n20743) );
  OAI221_X1 U23663 ( .B1(n20745), .B2(keyinput53), .C1(n20744), .C2(keyinput22), .A(n20743), .ZN(n20750) );
  AOI22_X1 U23664 ( .A1(n20748), .A2(keyinput1), .B1(n20747), .B2(keyinput57), 
        .ZN(n20746) );
  OAI221_X1 U23665 ( .B1(n20748), .B2(keyinput1), .C1(n20747), .C2(keyinput57), 
        .A(n20746), .ZN(n20749) );
  NOR4_X1 U23666 ( .A1(n20752), .A2(n20751), .A3(n20750), .A4(n20749), .ZN(
        n20800) );
  AOI22_X1 U23667 ( .A1(n20755), .A2(keyinput30), .B1(keyinput4), .B2(n20754), 
        .ZN(n20753) );
  OAI221_X1 U23668 ( .B1(n20755), .B2(keyinput30), .C1(n20754), .C2(keyinput4), 
        .A(n20753), .ZN(n20767) );
  INV_X1 U23669 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n20757) );
  AOI22_X1 U23670 ( .A1(n20757), .A2(keyinput49), .B1(n10835), .B2(keyinput10), 
        .ZN(n20756) );
  OAI221_X1 U23671 ( .B1(n20757), .B2(keyinput49), .C1(n10835), .C2(keyinput10), .A(n20756), .ZN(n20766) );
  INV_X1 U23672 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n20759) );
  AOI22_X1 U23673 ( .A1(n20760), .A2(keyinput12), .B1(keyinput18), .B2(n20759), 
        .ZN(n20758) );
  OAI221_X1 U23674 ( .B1(n20760), .B2(keyinput12), .C1(n20759), .C2(keyinput18), .A(n20758), .ZN(n20765) );
  AOI22_X1 U23675 ( .A1(n20763), .A2(keyinput16), .B1(keyinput62), .B2(n20762), 
        .ZN(n20761) );
  OAI221_X1 U23676 ( .B1(n20763), .B2(keyinput16), .C1(n20762), .C2(keyinput62), .A(n20761), .ZN(n20764) );
  NOR4_X1 U23677 ( .A1(n20767), .A2(n20766), .A3(n20765), .A4(n20764), .ZN(
        n20799) );
  AOI22_X1 U23678 ( .A1(n20770), .A2(keyinput3), .B1(keyinput33), .B2(n20769), 
        .ZN(n20768) );
  OAI221_X1 U23679 ( .B1(n20770), .B2(keyinput3), .C1(n20769), .C2(keyinput33), 
        .A(n20768), .ZN(n20782) );
  AOI22_X1 U23680 ( .A1(n20773), .A2(keyinput36), .B1(n20772), .B2(keyinput31), 
        .ZN(n20771) );
  OAI221_X1 U23681 ( .B1(n20773), .B2(keyinput36), .C1(n20772), .C2(keyinput31), .A(n20771), .ZN(n20781) );
  AOI22_X1 U23682 ( .A1(n11134), .A2(keyinput52), .B1(keyinput9), .B2(n20775), 
        .ZN(n20774) );
  OAI221_X1 U23683 ( .B1(n11134), .B2(keyinput52), .C1(n20775), .C2(keyinput9), 
        .A(n20774), .ZN(n20780) );
  AOI22_X1 U23684 ( .A1(n20778), .A2(keyinput25), .B1(keyinput26), .B2(n20777), 
        .ZN(n20776) );
  OAI221_X1 U23685 ( .B1(n20778), .B2(keyinput25), .C1(n20777), .C2(keyinput26), .A(n20776), .ZN(n20779) );
  NOR4_X1 U23686 ( .A1(n20782), .A2(n20781), .A3(n20780), .A4(n20779), .ZN(
        n20798) );
  INV_X1 U23687 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n20784) );
  AOI22_X1 U23688 ( .A1(n20785), .A2(keyinput28), .B1(n20784), .B2(keyinput56), 
        .ZN(n20783) );
  OAI221_X1 U23689 ( .B1(n20785), .B2(keyinput28), .C1(n20784), .C2(keyinput56), .A(n20783), .ZN(n20796) );
  INV_X1 U23690 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n20787) );
  AOI22_X1 U23691 ( .A1(n20808), .A2(keyinput15), .B1(keyinput55), .B2(n20787), 
        .ZN(n20786) );
  OAI221_X1 U23692 ( .B1(n20808), .B2(keyinput15), .C1(n20787), .C2(keyinput55), .A(n20786), .ZN(n20795) );
  INV_X1 U23693 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n20826) );
  AOI22_X1 U23694 ( .A1(n20789), .A2(keyinput11), .B1(keyinput39), .B2(n20826), 
        .ZN(n20788) );
  OAI221_X1 U23695 ( .B1(n20789), .B2(keyinput11), .C1(n20826), .C2(keyinput39), .A(n20788), .ZN(n20794) );
  AOI22_X1 U23696 ( .A1(n20792), .A2(keyinput24), .B1(keyinput38), .B2(n20791), 
        .ZN(n20790) );
  OAI221_X1 U23697 ( .B1(n20792), .B2(keyinput24), .C1(n20791), .C2(keyinput38), .A(n20790), .ZN(n20793) );
  NOR4_X1 U23698 ( .A1(n20796), .A2(n20795), .A3(n20794), .A4(n20793), .ZN(
        n20797) );
  NAND4_X1 U23699 ( .A1(n20800), .A2(n20799), .A3(n20798), .A4(n20797), .ZN(
        n20801) );
  NOR2_X1 U23700 ( .A1(n20802), .A2(n20801), .ZN(n20839) );
  OAI22_X1 U23701 ( .A1(n20806), .A2(n20805), .B1(n20804), .B2(n20803), .ZN(
        n20807) );
  AOI21_X1 U23702 ( .B1(P3_LWORD_REG_6__SCAN_IN), .B2(n17454), .A(n20807), 
        .ZN(n20837) );
  NOR4_X1 U23703 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_7__4__SCAN_IN), .A3(P1_INSTQUEUE_REG_1__2__SCAN_IN), 
        .A4(BUF2_REG_27__SCAN_IN), .ZN(n20835) );
  NAND4_X1 U23704 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A3(P2_DATAO_REG_26__SCAN_IN), 
        .A4(P3_UWORD_REG_13__SCAN_IN), .ZN(n20812) );
  NAND4_X1 U23705 ( .A1(P2_ADDRESS_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(P3_BE_N_REG_2__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20811) );
  INV_X1 U23706 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n20809) );
  NAND4_X1 U23707 ( .A1(n20741), .A2(n20809), .A3(n20808), .A4(
        P2_DATAWIDTH_REG_13__SCAN_IN), .ZN(n20810) );
  NOR3_X1 U23708 ( .A1(n20812), .A2(n20811), .A3(n20810), .ZN(n20834) );
  NAND4_X1 U23709 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_12__SCAN_IN), 
        .A4(P3_UWORD_REG_14__SCAN_IN), .ZN(n20816) );
  NAND4_X1 U23710 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_REIP_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_DATAO_REG_19__SCAN_IN), .ZN(n20815)
         );
  NAND4_X1 U23711 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_5__6__SCAN_IN), .A3(P2_EBX_REG_19__SCAN_IN), .A4(
        P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n20814) );
  NAND4_X1 U23712 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_8__6__SCAN_IN), .A3(BUF1_REG_26__SCAN_IN), .A4(
        DATAI_29_), .ZN(n20813) );
  NOR4_X1 U23713 ( .A1(n20816), .A2(n20815), .A3(n20814), .A4(n20813), .ZN(
        n20833) );
  NOR4_X1 U23714 ( .A1(P2_EBX_REG_8__SCAN_IN), .A2(P2_REIP_REG_21__SCAN_IN), 
        .A3(P2_CODEFETCH_REG_SCAN_IN), .A4(P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(
        n20820) );
  NOR4_X1 U23715 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A3(P3_EAX_REG_13__SCAN_IN), .A4(
        P3_DATAO_REG_15__SCAN_IN), .ZN(n20819) );
  NOR4_X1 U23716 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(
        P3_EBX_REG_18__SCAN_IN), .A3(P3_EBX_REG_15__SCAN_IN), .A4(
        P3_REIP_REG_7__SCAN_IN), .ZN(n20818) );
  NOR4_X1 U23717 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_4__1__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A4(BUF2_REG_20__SCAN_IN), .ZN(
        n20817) );
  NAND4_X1 U23718 ( .A1(n20820), .A2(n20819), .A3(n20818), .A4(n20817), .ZN(
        n20831) );
  NOR4_X1 U23719 ( .A1(P2_ADDRESS_REG_25__SCAN_IN), .A2(P1_EBX_REG_25__SCAN_IN), .A3(P3_ADDRESS_REG_18__SCAN_IN), .A4(P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(
        n20821) );
  NAND4_X1 U23720 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .A3(n20822), .A4(n20821), .ZN(n20830)
         );
  NAND4_X1 U23721 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20825), .A3(
        n20824), .A4(n20823), .ZN(n20829) );
  NAND4_X1 U23722 ( .A1(n9620), .A2(n20827), .A3(n13655), .A4(n20826), .ZN(
        n20828) );
  NOR4_X1 U23723 ( .A1(n20831), .A2(n20830), .A3(n20829), .A4(n20828), .ZN(
        n20832) );
  NAND4_X1 U23724 ( .A1(n20835), .A2(n20834), .A3(n20833), .A4(n20832), .ZN(
        n20836) );
  XNOR2_X1 U23725 ( .A(n20837), .B(n20836), .ZN(n20838) );
  XNOR2_X1 U23726 ( .A(n20839), .B(n20838), .ZN(P3_U2789) );
  CLKBUF_X1 U11052 ( .A(n11496), .Z(n11441) );
  BUF_X2 U11042 ( .A(n11409), .Z(n9594) );
  CLKBUF_X1 U11072 ( .A(n11255), .Z(n11706) );
  AND2_X1 U11079 ( .A1(n10583), .A2(n13306), .ZN(n10610) );
  CLKBUF_X2 U11080 ( .A(n11255), .Z(n9643) );
  CLKBUF_X1 U11090 ( .A(n10488), .Z(n12587) );
  CLKBUF_X1 U11094 ( .A(n9629), .Z(n12623) );
  CLKBUF_X1 U11254 ( .A(n11376), .Z(n12917) );
  NAND4_X1 U11271 ( .A1(n10905), .A2(n10904), .A3(n10903), .A4(n10902), .ZN(
        n15220) );
  NAND2_X1 U11314 ( .A1(n13691), .A2(n10538), .ZN(n10546) );
  CLKBUF_X1 U11352 ( .A(n12657), .Z(n9616) );
  CLKBUF_X1 U11368 ( .A(n10619), .Z(n9607) );
  CLKBUF_X1 U11376 ( .A(n15288), .Z(n15289) );
  CLKBUF_X1 U11390 ( .A(n10587), .Z(n9617) );
  CLKBUF_X1 U11436 ( .A(n14404), .Z(n14405) );
  XNOR2_X1 U11442 ( .A(n12151), .B(n12152), .ZN(n13258) );
  CLKBUF_X1 U11469 ( .A(n13094), .Z(n13137) );
endmodule

