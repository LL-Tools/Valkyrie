

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2014, n2015, n2016, n2017, n2018, n2019, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828;

  OR2_X1 U2256 ( .A1(n3863), .A2(n3864), .ZN(n3861) );
  OR2_X1 U2257 ( .A1(n4319), .A2(n4320), .ZN(n4317) );
  XNOR2_X1 U2258 ( .A(n2409), .B(n3601), .ZN(n3598) );
  XNOR2_X1 U2259 ( .A(n2399), .B(n3274), .ZN(n3271) );
  CLKBUF_X2 U2260 ( .A(n3018), .Z(n3062) );
  INV_X1 U2261 ( .A(n3447), .ZN(n3466) );
  CLKBUF_X2 U2262 ( .A(n4076), .Z(n2016) );
  CLKBUF_X2 U2263 ( .A(n2479), .Z(n3695) );
  INV_X1 U2264 ( .A(n3066), .ZN(n3051) );
  INV_X1 U2265 ( .A(n3324), .ZN(n2823) );
  OAI21_X1 U2266 ( .B1(n2024), .B2(n2081), .A(n2445), .ZN(n3240) );
  AND2_X2 U2267 ( .A1(n4712), .A2(n4711), .ZN(n2468) );
  INV_X1 U2268 ( .A(n2439), .ZN(n4712) );
  AND2_X2 U2269 ( .A1(n2015), .A2(n3455), .ZN(n3018) );
  NAND2_X1 U2270 ( .A1(n3191), .A2(n2386), .ZN(n2387) );
  NAND2_X1 U2271 ( .A1(n4097), .A2(n2408), .ZN(n2409) );
  INV_X1 U2272 ( .A(n2475), .ZN(n3336) );
  INV_X1 U2273 ( .A(n3525), .ZN(n3672) );
  XNOR2_X1 U2275 ( .A(n2387), .B(n3147), .ZN(n3139) );
  INV_X1 U2276 ( .A(n4074), .ZN(n3541) );
  INV_X1 U2277 ( .A(n3344), .ZN(n3430) );
  OR2_X1 U2278 ( .A1(n4761), .A2(n4763), .ZN(n4760) );
  AND2_X1 U2279 ( .A1(n4298), .A2(n4301), .ZN(n4299) );
  INV_X1 U2280 ( .A(IR_REG_31__SCAN_IN), .ZN(n2080) );
  AOI21_X1 U2281 ( .B1(n4760), .B2(n4768), .A(n4767), .ZN(n4774) );
  AND2_X2 U2282 ( .A1(n2824), .A2(n2829), .ZN(n2015) );
  NOR2_X2 U2283 ( .A1(n3517), .A2(n2076), .ZN(n3524) );
  OAI22_X1 U2284 ( .A1(n2948), .A2(n2189), .B1(n2026), .B2(n2973), .ZN(n3774)
         );
  XNOR2_X2 U2285 ( .A(n2244), .B(IR_REG_2__SCAN_IN), .ZN(n2384) );
  INV_X1 U2286 ( .A(n2469), .ZN(n2607) );
  NAND2_X1 U2287 ( .A1(n2865), .A2(n2223), .ZN(n3386) );
  AOI21_X1 U2288 ( .B1(n3204), .B2(n2267), .A(n2053), .ZN(n2270) );
  INV_X2 U2289 ( .A(n2852), .ZN(n2022) );
  NAND4_X1 U2290 ( .A1(n2504), .A2(n2503), .A3(n2502), .A4(n2501), .ZN(n4075)
         );
  INV_X4 U2291 ( .A(n2983), .ZN(n2852) );
  NAND4_X1 U2292 ( .A1(n2508), .A2(n2507), .A3(n2506), .A4(n2505), .ZN(n4074)
         );
  INV_X1 U2293 ( .A(n2840), .ZN(n3323) );
  NAND4_X1 U2294 ( .A1(n2465), .A2(n2464), .A3(n2463), .A4(n2462), .ZN(n3344)
         );
  BUF_X4 U2296 ( .A(n2468), .Z(n2014) );
  NAND2_X1 U2297 ( .A1(n2437), .A2(n2436), .ZN(n2439) );
  CLKBUF_X1 U2298 ( .A(n2380), .Z(n4728) );
  INV_X2 U2299 ( .A(IR_REG_0__SCAN_IN), .ZN(n2081) );
  NAND2_X1 U2300 ( .A1(n3048), .A2(n3047), .ZN(n3885) );
  OAI21_X1 U2301 ( .B1(n2180), .B2(n2816), .A(n2183), .ZN(n2822) );
  NAND2_X1 U2302 ( .A1(n2211), .A2(n2210), .ZN(n3762) );
  NAND2_X1 U2303 ( .A1(n2130), .A2(n4107), .ZN(n4106) );
  AND2_X1 U2304 ( .A1(n2106), .A2(n2105), .ZN(n4104) );
  NAND2_X1 U2305 ( .A1(n2732), .A2(n2187), .ZN(n4168) );
  AND2_X1 U2306 ( .A1(n2791), .A2(n2790), .ZN(n2792) );
  XNOR2_X1 U2307 ( .A(n4117), .B(n4057), .ZN(n3708) );
  NOR2_X1 U2308 ( .A1(n4118), .A2(n4119), .ZN(n4117) );
  XNOR2_X1 U2309 ( .A(n2309), .B(n4739), .ZN(n4736) );
  OR2_X1 U2310 ( .A1(n3683), .A2(n4006), .ZN(n3681) );
  NAND2_X1 U2311 ( .A1(n4191), .A2(n2075), .ZN(n4174) );
  NAND2_X1 U2312 ( .A1(n2194), .A2(n2196), .ZN(n3493) );
  NAND2_X1 U2313 ( .A1(n4087), .A2(n2290), .ZN(n4090) );
  NAND2_X1 U2314 ( .A1(n2138), .A2(n2136), .ZN(n3557) );
  OR2_X1 U2315 ( .A1(n3522), .A2(n2532), .ZN(n2138) );
  AOI21_X1 U2316 ( .B1(n2177), .B2(n2179), .A(n2176), .ZN(n2175) );
  AND2_X1 U2317 ( .A1(n3638), .A2(n3855), .ZN(n3646) );
  INV_X1 U2318 ( .A(n2178), .ZN(n2177) );
  NOR2_X2 U2319 ( .A1(n3564), .A2(n3590), .ZN(n3638) );
  NAND2_X1 U2320 ( .A1(n2135), .A2(n2134), .ZN(n3452) );
  NAND2_X1 U2321 ( .A1(n2171), .A2(n2047), .ZN(n2170) );
  XNOR2_X1 U2322 ( .A(n2270), .B(n4721), .ZN(n3270) );
  OR2_X1 U2323 ( .A1(n3930), .A2(n2708), .ZN(n2710) );
  AND2_X1 U2324 ( .A1(n3918), .A2(n3915), .ZN(n3990) );
  AND4_X1 U2325 ( .A1(n2444), .A2(n2443), .A3(n2442), .A4(n2441), .ZN(n3324)
         );
  INV_X1 U2326 ( .A(n3313), .ZN(n2829) );
  AND2_X2 U2327 ( .A1(n2438), .A2(n2439), .ZN(n2461) );
  OAI21_X1 U2328 ( .B1(n3694), .B2(n2458), .A(n2457), .ZN(n3291) );
  NAND2_X1 U2329 ( .A1(n2741), .A2(n2740), .ZN(n4465) );
  OR2_X1 U2330 ( .A1(n3199), .A2(n4716), .ZN(n3455) );
  NAND2_X1 U2331 ( .A1(n2341), .A2(IR_REG_31__SCAN_IN), .ZN(n2342) );
  AND2_X1 U2332 ( .A1(n2694), .A2(n4715), .ZN(n3313) );
  AND2_X1 U2333 ( .A1(n2353), .A2(n2370), .ZN(n3118) );
  NAND2_X1 U2334 ( .A1(n2389), .A2(n2388), .ZN(n2390) );
  OR2_X1 U2336 ( .A1(n2023), .A2(n2447), .ZN(n2160) );
  XNOR2_X1 U2337 ( .A(n2692), .B(n2691), .ZN(n2694) );
  INV_X1 U2338 ( .A(n2074), .ZN(n2073) );
  XNOR2_X1 U2339 ( .A(n2362), .B(IR_REG_22__SCAN_IN), .ZN(n4714) );
  MUX2_X1 U2340 ( .A(IR_REG_31__SCAN_IN), .B(n2435), .S(IR_REG_29__SCAN_IN), 
        .Z(n2437) );
  MUX2_X1 U2341 ( .A(IR_REG_31__SCAN_IN), .B(n2359), .S(IR_REG_21__SCAN_IN), 
        .Z(n2360) );
  NAND2_X1 U2342 ( .A1(n2690), .A2(IR_REG_31__SCAN_IN), .ZN(n2692) );
  XNOR2_X1 U2343 ( .A(n2354), .B(IR_REG_26__SCAN_IN), .ZN(n3126) );
  OR2_X1 U2344 ( .A1(n2370), .A2(n2218), .ZN(n2434) );
  OAI21_X1 U2345 ( .B1(n2331), .B2(IR_REG_18__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2333) );
  NAND2_X2 U2346 ( .A1(n2352), .A2(n2351), .ZN(n2370) );
  NOR2_X1 U2347 ( .A1(n2350), .A2(n2349), .ZN(n2351) );
  NAND2_X1 U2348 ( .A1(n2235), .A2(n2234), .ZN(n2299) );
  NAND3_X1 U2349 ( .A1(n2079), .A2(n2078), .A3(n2077), .ZN(n2380) );
  NAND2_X1 U2350 ( .A1(n2243), .A2(IR_REG_31__SCAN_IN), .ZN(n2244) );
  AND2_X1 U2351 ( .A1(n2067), .A2(n2324), .ZN(n2338) );
  NOR2_X1 U2352 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2234)
         );
  NOR2_X1 U2353 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2066)
         );
  NOR2_X1 U2354 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2065)
         );
  NOR2_X1 U2355 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2064)
         );
  NOR2_X1 U2356 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2294)
         );
  NOR2_X1 U2357 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2295)
         );
  INV_X1 U2358 ( .A(IR_REG_24__SCAN_IN), .ZN(n2346) );
  NOR2_X1 U2359 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2296)
         );
  NAND2_X2 U2360 ( .A1(n2204), .A2(n3794), .ZN(n3747) );
  NOR2_X2 U2361 ( .A1(n4742), .A2(n4741), .ZN(n4740) );
  NAND2_X2 U2362 ( .A1(n3208), .A2(n2398), .ZN(n2399) );
  NOR2_X2 U2363 ( .A1(n3240), .A2(n2832), .ZN(n3239) );
  NAND2_X2 U2364 ( .A1(n2160), .A2(n2446), .ZN(n2832) );
  NAND2_X1 U2365 ( .A1(n3158), .A2(n2393), .ZN(n2394) );
  INV_X4 U2366 ( .A(n2852), .ZN(n3063) );
  OAI21_X2 U2367 ( .B1(n3493), .B2(n3495), .A(n3494), .ZN(n3548) );
  NOR2_X4 U2368 ( .A1(n2299), .A2(n2298), .ZN(n2352) );
  NAND2_X1 U2369 ( .A1(n2073), .A2(n2072), .ZN(n2017) );
  INV_X1 U2370 ( .A(n2017), .ZN(n2018) );
  NAND4_X2 U2371 ( .A1(n2452), .A2(n2451), .A3(n2450), .A4(n2449), .ZN(n2459)
         );
  AND2_X1 U2372 ( .A1(n2438), .A2(n2439), .ZN(n2019) );
  XNOR2_X2 U2373 ( .A(n2342), .B(IR_REG_24__SCAN_IN), .ZN(n2748) );
  NAND2_X1 U2374 ( .A1(n2073), .A2(n2072), .ZN(n2023) );
  NAND2_X1 U2375 ( .A1(n2073), .A2(n2072), .ZN(n2024) );
  INV_X1 U2376 ( .A(n2410), .ZN(n2122) );
  AND2_X1 U2377 ( .A1(n2150), .A2(n2155), .ZN(n2149) );
  NOR2_X1 U2378 ( .A1(n2680), .A2(n2156), .ZN(n2155) );
  NAND2_X1 U2379 ( .A1(n2153), .A2(n2151), .ZN(n2150) );
  INV_X1 U2380 ( .A(n2157), .ZN(n2156) );
  INV_X1 U2381 ( .A(n2153), .ZN(n2152) );
  OR2_X1 U2382 ( .A1(n2682), .A2(n2681), .ZN(n2697) );
  OR2_X1 U2383 ( .A1(n4387), .A2(n4177), .ZN(n4148) );
  AND2_X1 U2384 ( .A1(n2035), .A2(n2489), .ZN(n2134) );
  OR2_X1 U2385 ( .A1(n4143), .A2(n4129), .ZN(n3973) );
  NAND4_X1 U2386 ( .A1(n2297), .A2(n2296), .A3(n2295), .A4(n2294), .ZN(n2298)
         );
  NAND2_X1 U2387 ( .A1(n2063), .A2(n2656), .ZN(n2666) );
  NAND2_X1 U2388 ( .A1(n2062), .A2(REG3_REG_26__SCAN_IN), .ZN(n2682) );
  NOR2_X1 U2389 ( .A1(n3156), .A2(n2097), .ZN(n2260) );
  NOR2_X1 U2390 ( .A1(n3163), .A2(n2098), .ZN(n2097) );
  INV_X1 U2391 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2098) );
  NAND2_X1 U2392 ( .A1(n2282), .A2(n4719), .ZN(n2283) );
  NAND2_X1 U2393 ( .A1(n3474), .A2(REG1_REG_10__SCAN_IN), .ZN(n2284) );
  NAND2_X1 U2394 ( .A1(n2333), .A2(n2332), .ZN(n2690) );
  OAI22_X1 U2395 ( .A1(n2775), .A2(n2774), .B1(n4157), .B2(n4140), .ZN(n3734)
         );
  AND2_X1 U2396 ( .A1(n4039), .A2(n2733), .ZN(n2187) );
  INV_X1 U2397 ( .A(n4040), .ZN(n2733) );
  AND2_X2 U2398 ( .A1(n2438), .A2(n4712), .ZN(n2479) );
  NOR2_X1 U2399 ( .A1(n2809), .A2(n2182), .ZN(n2181) );
  INV_X1 U2400 ( .A(n2806), .ZN(n2182) );
  NOR2_X1 U2401 ( .A1(n2168), .A2(n2167), .ZN(n2166) );
  INV_X1 U2402 ( .A(n2047), .ZN(n2168) );
  NAND2_X1 U2403 ( .A1(n2219), .A2(n2372), .ZN(n2218) );
  INV_X1 U2404 ( .A(n2369), .ZN(n2219) );
  NAND2_X1 U2405 ( .A1(n2192), .A2(n2960), .ZN(n2189) );
  NAND2_X1 U2406 ( .A1(n2124), .A2(n2412), .ZN(n2413) );
  NAND2_X1 U2407 ( .A1(n2123), .A2(n2121), .ZN(n2124) );
  NOR2_X1 U2408 ( .A1(n2122), .A2(n2411), .ZN(n2121) );
  NAND2_X1 U2409 ( .A1(n2414), .A2(REG2_REG_14__SCAN_IN), .ZN(n2126) );
  INV_X1 U2410 ( .A(n2492), .ZN(n2490) );
  OR2_X1 U2411 ( .A1(n3565), .A2(n3566), .ZN(n3564) );
  AND2_X1 U2412 ( .A1(n2823), .A2(n3240), .ZN(n3232) );
  NAND2_X1 U2413 ( .A1(n3232), .A2(n3231), .ZN(n3287) );
  INV_X1 U2414 ( .A(n2218), .ZN(n2216) );
  INV_X1 U2415 ( .A(IR_REG_6__SCAN_IN), .ZN(n2262) );
  INV_X1 U2416 ( .A(IR_REG_2__SCAN_IN), .ZN(n2233) );
  NAND2_X1 U2417 ( .A1(n2203), .A2(n2202), .ZN(n2201) );
  INV_X1 U2418 ( .A(n3397), .ZN(n2202) );
  INV_X1 U2419 ( .A(n3396), .ZN(n2203) );
  INV_X1 U2420 ( .A(n3840), .ZN(n2213) );
  NOR2_X1 U2421 ( .A1(n3019), .A2(n2215), .ZN(n2214) );
  INV_X1 U2422 ( .A(n3842), .ZN(n2215) );
  OR2_X1 U2423 ( .A1(n3764), .A2(n3026), .ZN(n3019) );
  AND2_X1 U2424 ( .A1(n2201), .A2(n3439), .ZN(n2195) );
  NAND2_X1 U2425 ( .A1(n2513), .A2(n2512), .ZN(n2526) );
  AND2_X1 U2426 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2512) );
  INV_X1 U2427 ( .A(n2516), .ZN(n2513) );
  INV_X1 U2428 ( .A(n2604), .ZN(n2586) );
  OR2_X1 U2429 ( .A1(n2596), .A2(n3844), .ZN(n2630) );
  AND2_X1 U2430 ( .A1(n2926), .A2(n2927), .ZN(n3795) );
  NAND2_X1 U2431 ( .A1(n2207), .A2(n3616), .ZN(n2206) );
  AND2_X1 U2432 ( .A1(n2914), .A2(n2209), .ZN(n2208) );
  INV_X1 U2433 ( .A(n3617), .ZN(n2209) );
  NAND2_X1 U2434 ( .A1(n2480), .A2(REG3_REG_5__SCAN_IN), .ZN(n2492) );
  NAND2_X1 U2435 ( .A1(n2060), .A2(n2567), .ZN(n2579) );
  AND2_X1 U2436 ( .A1(REG3_REG_15__SCAN_IN), .A2(REG3_REG_14__SCAN_IN), .ZN(
        n2567) );
  INV_X1 U2437 ( .A(n2569), .ZN(n2060) );
  OAI21_X1 U2438 ( .B1(n3978), .B2(n4049), .A(n3977), .ZN(n4050) );
  AND2_X1 U2439 ( .A1(n3063), .A2(n3093), .ZN(n3100) );
  XNOR2_X1 U2440 ( .A(n2380), .B(n2241), .ZN(n4080) );
  OAI21_X1 U2441 ( .B1(n2384), .B2(n2245), .A(n2246), .ZN(n3185) );
  CLKBUF_X1 U2442 ( .A(n2299), .Z(n2236) );
  INV_X1 U2443 ( .A(n2391), .ZN(n2120) );
  AOI21_X1 U2444 ( .B1(n2391), .B2(n2119), .A(n2118), .ZN(n2116) );
  INV_X1 U2445 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2119) );
  NOR2_X1 U2446 ( .A1(n3477), .A2(n2114), .ZN(n2113) );
  NAND2_X1 U2447 ( .A1(n2404), .A2(n2403), .ZN(n2108) );
  NAND2_X1 U2448 ( .A1(n2052), .A2(n4718), .ZN(n2086) );
  AOI21_X1 U2449 ( .B1(n2091), .B2(REG1_REG_12__SCAN_IN), .A(n4718), .ZN(n2088) );
  NAND2_X1 U2450 ( .A1(n4090), .A2(n2087), .ZN(n2085) );
  INV_X1 U2451 ( .A(n2126), .ZN(n2125) );
  NAND2_X1 U2452 ( .A1(n4751), .A2(n2418), .ZN(n2130) );
  OAI21_X1 U2453 ( .B1(n2104), .B2(n2105), .A(n2221), .ZN(n2103) );
  INV_X1 U2454 ( .A(n2104), .ZN(n2101) );
  NAND2_X1 U2455 ( .A1(n4150), .A2(n2034), .ZN(n2798) );
  AND2_X1 U2456 ( .A1(n2697), .A2(n2683), .ZN(n4136) );
  INV_X1 U2457 ( .A(n3695), .ZN(n2701) );
  INV_X1 U2458 ( .A(n2468), .ZN(n2777) );
  NAND2_X1 U2459 ( .A1(n3738), .A2(n2698), .ZN(n3085) );
  OR2_X1 U2460 ( .A1(n4196), .A2(n4177), .ZN(n2157) );
  AND2_X1 U2461 ( .A1(n2159), .A2(n2041), .ZN(n2153) );
  NAND2_X1 U2462 ( .A1(n4185), .A2(n2665), .ZN(n2154) );
  NAND2_X1 U2463 ( .A1(n2628), .A2(REG3_REG_21__SCAN_IN), .ZN(n2641) );
  INV_X1 U2464 ( .A(n2630), .ZN(n2628) );
  INV_X1 U2465 ( .A(n2063), .ZN(n2655) );
  NAND2_X1 U2466 ( .A1(n2184), .A2(n4035), .ZN(n4238) );
  AND2_X1 U2467 ( .A1(n2024), .A2(DATAI_20_), .ZN(n4415) );
  INV_X1 U2468 ( .A(n2061), .ZN(n2612) );
  NAND2_X1 U2469 ( .A1(n4347), .A2(n3952), .ZN(n4326) );
  INV_X1 U2470 ( .A(n2577), .ZN(n2132) );
  INV_X1 U2471 ( .A(n2578), .ZN(n2133) );
  NOR2_X1 U2472 ( .A1(n3991), .A2(n2137), .ZN(n2136) );
  INV_X1 U2473 ( .A(n2533), .ZN(n2137) );
  AOI21_X1 U2474 ( .B1(n3452), .B2(n2231), .A(n2511), .ZN(n3538) );
  NAND2_X1 U2475 ( .A1(n2770), .A2(n2769), .ZN(n3517) );
  NAND2_X1 U2476 ( .A1(n3937), .A2(n2172), .ZN(n2171) );
  INV_X1 U2477 ( .A(n3305), .ZN(n3216) );
  NAND2_X1 U2478 ( .A1(n3324), .A2(n3240), .ZN(n3198) );
  NAND2_X1 U2479 ( .A1(n2788), .A2(n2068), .ZN(n4118) );
  NOR2_X1 U2480 ( .A1(n3965), .A2(n3068), .ZN(n2068) );
  OAI211_X1 U2481 ( .C1(n3734), .C2(n2813), .A(n2142), .B(n2815), .ZN(n2141)
         );
  INV_X1 U2482 ( .A(n2814), .ZN(n2815) );
  NAND2_X1 U2483 ( .A1(n3734), .A2(n2143), .ZN(n2142) );
  NAND2_X1 U2484 ( .A1(n2788), .A2(n4129), .ZN(n2817) );
  AND2_X1 U2485 ( .A1(n2771), .A2(n4140), .ZN(n2788) );
  NOR2_X2 U2486 ( .A1(n4174), .A2(n4154), .ZN(n2771) );
  NAND2_X1 U2487 ( .A1(n3524), .A2(n3572), .ZN(n3565) );
  INV_X1 U2488 ( .A(n3606), .ZN(n3543) );
  INV_X1 U2489 ( .A(n4727), .ZN(n2458) );
  NAND2_X1 U2490 ( .A1(n2024), .A2(DATAI_2_), .ZN(n2457) );
  NOR2_X1 U2491 ( .A1(n2751), .A2(n2752), .ZN(n3125) );
  XNOR2_X1 U2492 ( .A(n2433), .B(IR_REG_30__SCAN_IN), .ZN(n2440) );
  NAND2_X1 U2493 ( .A1(n2436), .A2(IR_REG_31__SCAN_IN), .ZN(n2433) );
  INV_X1 U2494 ( .A(IR_REG_23__SCAN_IN), .ZN(n2356) );
  INV_X1 U2495 ( .A(IR_REG_20__SCAN_IN), .ZN(n2691) );
  AND4_X1 U2496 ( .A1(n2325), .A2(n4497), .A3(n4496), .A4(n2324), .ZN(n2326)
         );
  OR2_X1 U2497 ( .A1(n2280), .A2(IR_REG_9__SCAN_IN), .ZN(n2285) );
  INV_X1 U2498 ( .A(IR_REG_7__SCAN_IN), .ZN(n2264) );
  NAND2_X1 U2499 ( .A1(n3396), .A2(n3397), .ZN(n2199) );
  AND2_X1 U2500 ( .A1(n2674), .A2(n2667), .ZN(n4175) );
  INV_X1 U2501 ( .A(n4414), .ZN(n3866) );
  NAND4_X1 U2502 ( .A1(n2561), .A2(n2560), .A3(n2559), .A4(n2558), .ZN(n4474)
         );
  XNOR2_X1 U2503 ( .A(n2390), .B(n3253), .ZN(n3249) );
  OAI21_X1 U2504 ( .B1(n3255), .B2(n2096), .A(n2094), .ZN(n3156) );
  NAND2_X1 U2505 ( .A1(n2095), .A2(REG1_REG_4__SCAN_IN), .ZN(n2096) );
  NAND2_X1 U2506 ( .A1(n3169), .A2(REG1_REG_6__SCAN_IN), .ZN(n3168) );
  NAND2_X1 U2507 ( .A1(n4090), .A2(n2093), .ZN(n2089) );
  OAI21_X1 U2508 ( .B1(n4107), .B2(n2130), .A(n4106), .ZN(n2129) );
  INV_X1 U2509 ( .A(n2128), .ZN(n2127) );
  AOI21_X1 U2510 ( .B1(n4765), .B2(ADDR_REG_17__SCAN_IN), .A(n4108), .ZN(n2128) );
  NAND2_X1 U2511 ( .A1(n2690), .A2(n2334), .ZN(n4063) );
  OR2_X1 U2512 ( .A1(n2333), .A2(n2332), .ZN(n2334) );
  NAND2_X1 U2513 ( .A1(n2807), .A2(n2048), .ZN(n2180) );
  INV_X1 U2514 ( .A(n2141), .ZN(n2816) );
  NAND2_X1 U2515 ( .A1(n4828), .A2(n4640), .ZN(n4484) );
  OR2_X1 U2516 ( .A1(n2947), .A2(n2191), .ZN(n2190) );
  INV_X1 U2517 ( .A(n2665), .ZN(n2151) );
  NAND2_X1 U2518 ( .A1(n3323), .A2(n3291), .ZN(n3912) );
  NAND2_X1 U2519 ( .A1(n3330), .A2(n2459), .ZN(n3909) );
  INV_X1 U2521 ( .A(n2546), .ZN(n2544) );
  NAND2_X1 U2522 ( .A1(n3183), .A2(n2247), .ZN(n2249) );
  NAND2_X1 U2523 ( .A1(n4727), .A2(REG1_REG_2__SCAN_IN), .ZN(n2247) );
  INV_X1 U2524 ( .A(n3160), .ZN(n2118) );
  NOR2_X1 U2525 ( .A1(n2049), .A2(n4499), .ZN(n2087) );
  INV_X1 U2526 ( .A(n2092), .ZN(n2090) );
  NAND2_X1 U2527 ( .A1(n4718), .A2(n2092), .ZN(n2091) );
  OR2_X1 U2528 ( .A1(n4137), .A2(n4159), .ZN(n2734) );
  AND2_X1 U2529 ( .A1(n3961), .A2(n2731), .ZN(n4036) );
  NOR2_X1 U2530 ( .A1(n2641), .A2(n4579), .ZN(n2063) );
  OR2_X1 U2531 ( .A1(n2620), .A2(n2619), .ZN(n2625) );
  NOR2_X1 U2532 ( .A1(n2610), .A2(n2609), .ZN(n2061) );
  INV_X1 U2533 ( .A(n3945), .ZN(n2176) );
  OAI21_X1 U2534 ( .B1(n2713), .B2(n2179), .A(n3943), .ZN(n2178) );
  INV_X1 U2535 ( .A(n3944), .ZN(n2179) );
  NAND2_X1 U2536 ( .A1(n2163), .A2(n3936), .ZN(n2162) );
  INV_X1 U2537 ( .A(n2170), .ZN(n2163) );
  NAND2_X1 U2538 ( .A1(n2448), .A2(n2832), .ZN(n3913) );
  AND2_X1 U2539 ( .A1(n3733), .A2(n2811), .ZN(n2143) );
  OR2_X1 U2540 ( .A1(n4431), .A2(n4352), .ZN(n4313) );
  NOR2_X1 U2541 ( .A1(n3685), .A2(n4449), .ZN(n3686) );
  NAND2_X1 U2542 ( .A1(n3916), .A2(n3912), .ZN(n3289) );
  NAND2_X1 U2543 ( .A1(n2366), .A2(IR_REG_28__SCAN_IN), .ZN(n2072) );
  OAI21_X1 U2544 ( .B1(n2366), .B2(IR_REG_27__SCAN_IN), .A(n2364), .ZN(n2074)
         );
  AND2_X1 U2545 ( .A1(n4715), .A2(n4714), .ZN(n3075) );
  INV_X1 U2546 ( .A(n3198), .ZN(n3911) );
  NAND2_X1 U2547 ( .A1(n2368), .A2(n2367), .ZN(n2369) );
  INV_X1 U2548 ( .A(IR_REG_27__SCAN_IN), .ZN(n2368) );
  AND2_X1 U2549 ( .A1(n2352), .A2(n2339), .ZN(n2357) );
  INV_X1 U2550 ( .A(IR_REG_17__SCAN_IN), .ZN(n4497) );
  INV_X1 U2551 ( .A(IR_REG_13__SCAN_IN), .ZN(n4496) );
  INV_X1 U2552 ( .A(IR_REG_11__SCAN_IN), .ZN(n2286) );
  AND2_X1 U2553 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2480) );
  OR2_X1 U2554 ( .A1(n2579), .A2(n4610), .ZN(n2610) );
  INV_X1 U2555 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2609) );
  INV_X1 U2556 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2555) );
  NAND2_X1 U2557 ( .A1(n2544), .A2(REG3_REG_12__SCAN_IN), .ZN(n2556) );
  NAND2_X1 U2558 ( .A1(n2525), .A2(REG3_REG_10__SCAN_IN), .ZN(n2534) );
  INV_X1 U2559 ( .A(n2526), .ZN(n2525) );
  OR2_X1 U2560 ( .A1(n2534), .A2(n4521), .ZN(n2546) );
  AOI22_X1 U2561 ( .A1(n3018), .A2(n2459), .B1(n2983), .B2(n2832), .ZN(n2836)
         );
  XNOR2_X1 U2562 ( .A(n2835), .B(n3066), .ZN(n2838) );
  NAND2_X1 U2563 ( .A1(n2490), .A2(REG3_REG_6__SCAN_IN), .ZN(n2499) );
  XNOR2_X1 U2564 ( .A(n2864), .B(n3066), .ZN(n2868) );
  NAND2_X1 U2565 ( .A1(n2544), .A2(n2059), .ZN(n2569) );
  NOR2_X1 U2566 ( .A1(n2555), .A2(n2545), .ZN(n2059) );
  NAND2_X1 U2567 ( .A1(n2019), .A2(REG0_REG_1__SCAN_IN), .ZN(n2449) );
  NAND2_X1 U2568 ( .A1(n2469), .A2(REG2_REG_1__SCAN_IN), .ZN(n2451) );
  NAND2_X1 U2569 ( .A1(n2479), .A2(REG1_REG_1__SCAN_IN), .ZN(n2450) );
  NAND2_X1 U2570 ( .A1(n4078), .A2(n2242), .ZN(n3184) );
  XNOR2_X1 U2571 ( .A(n2249), .B(n4726), .ZN(n3141) );
  NOR2_X1 U2572 ( .A1(n3141), .A2(n3142), .ZN(n3140) );
  NOR2_X1 U2573 ( .A1(n3140), .A2(n2250), .ZN(n2255) );
  AND2_X1 U2574 ( .A1(n2249), .A2(n4726), .ZN(n2250) );
  INV_X1 U2575 ( .A(n3487), .ZN(n2278) );
  AND2_X1 U2576 ( .A1(n2113), .A2(REG2_REG_10__SCAN_IN), .ZN(n2109) );
  NOR2_X1 U2577 ( .A1(n2052), .A2(n3601), .ZN(n2093) );
  NAND2_X1 U2578 ( .A1(n3660), .A2(n2307), .ZN(n2309) );
  NAND2_X1 U2579 ( .A1(n2084), .A2(n2082), .ZN(n2318) );
  NAND2_X1 U2580 ( .A1(n2083), .A2(n2046), .ZN(n2082) );
  NAND2_X1 U2581 ( .A1(n4736), .A2(n2050), .ZN(n2084) );
  NAND2_X1 U2582 ( .A1(n4745), .A2(n2313), .ZN(n2083) );
  INV_X1 U2583 ( .A(n4105), .ZN(n2105) );
  NAND2_X1 U2584 ( .A1(n2328), .A2(n4772), .ZN(n2104) );
  INV_X1 U2585 ( .A(IR_REG_19__SCAN_IN), .ZN(n2332) );
  NAND2_X1 U2586 ( .A1(n2032), .A2(n3972), .ZN(n2797) );
  NAND2_X1 U2587 ( .A1(n2148), .A2(n2147), .ZN(n2775) );
  AOI21_X1 U2588 ( .B1(n2149), .B2(n2152), .A(n2038), .ZN(n2147) );
  AND2_X1 U2589 ( .A1(n2033), .A2(n2577), .ZN(n2131) );
  NOR2_X1 U2590 ( .A1(n3955), .A2(n2186), .ZN(n2185) );
  NAND2_X1 U2591 ( .A1(n2061), .A2(REG3_REG_18__SCAN_IN), .ZN(n2604) );
  AOI21_X1 U2592 ( .B1(n2025), .B2(n2562), .A(n2051), .ZN(n2145) );
  NAND2_X1 U2593 ( .A1(n2490), .A2(n2037), .ZN(n2516) );
  INV_X1 U2594 ( .A(n3998), .ZN(n3924) );
  OR2_X1 U2595 ( .A1(n3453), .A2(n3924), .ZN(n3505) );
  NAND2_X1 U2596 ( .A1(n3374), .A2(n2488), .ZN(n2135) );
  NAND2_X1 U2597 ( .A1(n2461), .A2(REG0_REG_4__SCAN_IN), .ZN(n2471) );
  INV_X1 U2598 ( .A(n3919), .ZN(n2173) );
  INV_X1 U2599 ( .A(n4465), .ZN(n4327) );
  NAND2_X1 U2600 ( .A1(n2023), .A2(DATAI_0_), .ZN(n2445) );
  INV_X1 U2601 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4610) );
  NOR2_X1 U2602 ( .A1(n4386), .A2(n4377), .ZN(n2075) );
  NAND2_X1 U2603 ( .A1(n4191), .A2(n4195), .ZN(n4192) );
  INV_X1 U2604 ( .A(n4207), .ZN(n4216) );
  NAND2_X1 U2605 ( .A1(n4299), .A2(n2056), .ZN(n4244) );
  NAND2_X1 U2606 ( .A1(n4299), .A2(n4277), .ZN(n4273) );
  INV_X1 U2607 ( .A(n4291), .ZN(n4301) );
  NAND2_X1 U2608 ( .A1(n3646), .A2(n3756), .ZN(n3685) );
  INV_X1 U2609 ( .A(n3627), .ZN(n3855) );
  INV_X1 U2610 ( .A(n3668), .ZN(n3572) );
  NOR2_X1 U2611 ( .A1(n3517), .A2(n3516), .ZN(n3515) );
  NAND2_X1 U2612 ( .A1(n3543), .A2(n2707), .ZN(n2076) );
  OR2_X1 U2613 ( .A1(n4786), .A2(n4714), .ZN(n4644) );
  INV_X1 U2614 ( .A(n4458), .ZN(n4477) );
  INV_X1 U2615 ( .A(n4075), .ZN(n3510) );
  NAND2_X1 U2616 ( .A1(n3336), .A2(n2070), .ZN(n2069) );
  NAND2_X1 U2617 ( .A1(n2071), .A2(n3336), .ZN(n3369) );
  NAND2_X1 U2618 ( .A1(n3561), .A2(n4644), .ZN(n4482) );
  INV_X1 U2619 ( .A(n4462), .ZN(n4475) );
  INV_X1 U2620 ( .A(n3455), .ZN(n4640) );
  INV_X1 U2621 ( .A(n3126), .ZN(n2752) );
  INV_X1 U2622 ( .A(IR_REG_29__SCAN_IN), .ZN(n2432) );
  OR2_X1 U2623 ( .A1(n2275), .A2(n2274), .ZN(n2280) );
  NAND2_X1 U2624 ( .A1(n2239), .A2(n2238), .ZN(n2261) );
  INV_X1 U2625 ( .A(IR_REG_5__SCAN_IN), .ZN(n2238) );
  NAND2_X1 U2626 ( .A1(n2193), .A2(n2081), .ZN(n2243) );
  NAND2_X1 U2627 ( .A1(n2080), .A2(IR_REG_1__SCAN_IN), .ZN(n2079) );
  NAND3_X1 U2628 ( .A1(n2193), .A2(IR_REG_31__SCAN_IN), .A3(IR_REG_0__SCAN_IN), 
        .ZN(n2078) );
  NAND2_X1 U2629 ( .A1(n2081), .A2(IR_REG_1__SCAN_IN), .ZN(n2077) );
  NAND2_X1 U2630 ( .A1(n3399), .A2(n2201), .ZN(n2200) );
  AOI21_X1 U2631 ( .B1(n3885), .B2(n3882), .A(n3881), .ZN(n3725) );
  OR2_X1 U2632 ( .A1(n3710), .A2(n2214), .ZN(n2210) );
  NOR2_X1 U2633 ( .A1(n3710), .A2(n2213), .ZN(n2212) );
  INV_X1 U2634 ( .A(n2197), .ZN(n2196) );
  OAI21_X1 U2635 ( .B1(n2199), .B2(n2198), .A(n2887), .ZN(n2197) );
  NAND2_X1 U2636 ( .A1(n3838), .A2(n3842), .ZN(n3763) );
  INV_X1 U2637 ( .A(n4473), .ZN(n3799) );
  INV_X1 U2638 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3844) );
  INV_X1 U2639 ( .A(n3795), .ZN(n2205) );
  INV_X1 U2640 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4579) );
  OR2_X1 U2641 ( .A1(n3101), .A2(n4067), .ZN(n3865) );
  OR2_X1 U2642 ( .A1(n3101), .A2(n3099), .ZN(n3898) );
  NAND2_X1 U2643 ( .A1(n2682), .A2(n2675), .ZN(n4161) );
  INV_X1 U2644 ( .A(n3898), .ZN(n3890) );
  OR2_X1 U2645 ( .A1(n3101), .A2(n3079), .ZN(n3907) );
  INV_X1 U2646 ( .A(n3865), .ZN(n3902) );
  INV_X1 U2647 ( .A(n3886), .ZN(n3904) );
  MUX2_X1 U2648 ( .A(n4062), .B(n4061), .S(n4716), .Z(n4064) );
  NAND2_X1 U2649 ( .A1(n2688), .A2(n2687), .ZN(n4124) );
  NAND2_X1 U2650 ( .A1(n2672), .A2(n2671), .ZN(n4387) );
  NAND2_X1 U2651 ( .A1(n2662), .A2(n2661), .ZN(n4378) );
  OR2_X1 U2652 ( .A1(n3832), .A2(n2777), .ZN(n2662) );
  NAND2_X1 U2653 ( .A1(n2647), .A2(n2646), .ZN(n4247) );
  NAND2_X1 U2654 ( .A1(n2636), .A2(n2635), .ZN(n4414) );
  NAND2_X1 U2655 ( .A1(n2593), .A2(n2592), .ZN(n4405) );
  NAND2_X1 U2656 ( .A1(n2601), .A2(n2600), .ZN(n4416) );
  OAI211_X1 U2657 ( .C1(n4333), .C2(n2777), .A(n2614), .B(n2613), .ZN(n4441)
         );
  NAND4_X1 U2658 ( .A1(n2584), .A2(n2583), .A3(n2582), .A4(n2581), .ZN(n4432)
         );
  NAND4_X1 U2659 ( .A1(n2574), .A2(n2573), .A3(n2572), .A4(n2571), .ZN(n4440)
         );
  NAND2_X1 U2660 ( .A1(n2461), .A2(REG0_REG_3__SCAN_IN), .ZN(n2462) );
  XNOR2_X1 U2661 ( .A(n2380), .B(n3326), .ZN(n4082) );
  OR2_X1 U2662 ( .A1(n3255), .A2(n4826), .ZN(n2099) );
  NAND2_X1 U2663 ( .A1(n2117), .A2(n2391), .ZN(n3159) );
  NAND2_X1 U2664 ( .A1(n3249), .A2(REG2_REG_4__SCAN_IN), .ZN(n2117) );
  NAND2_X1 U2665 ( .A1(n3168), .A2(n2220), .ZN(n3204) );
  NAND2_X1 U2666 ( .A1(n2404), .A2(n2113), .ZN(n2112) );
  NAND2_X1 U2667 ( .A1(n2108), .A2(n3477), .ZN(n2115) );
  NAND2_X1 U2668 ( .A1(n3601), .A2(n2052), .ZN(n2092) );
  INV_X1 U2669 ( .A(n4088), .ZN(n2290) );
  NAND2_X1 U2670 ( .A1(n2123), .A2(n2410), .ZN(n3656) );
  NAND2_X1 U2671 ( .A1(n2029), .A2(n2414), .ZN(n4731) );
  XNOR2_X1 U2672 ( .A(n2318), .B(n2585), .ZN(n4757) );
  OR2_X1 U2673 ( .A1(n4104), .A2(n2104), .ZN(n4769) );
  OR2_X1 U2674 ( .A1(n3152), .A2(n4713), .ZN(n4775) );
  XNOR2_X1 U2675 ( .A(n2427), .B(n2426), .ZN(n2429) );
  NAND2_X1 U2676 ( .A1(n4760), .A2(n2423), .ZN(n2427) );
  INV_X1 U2677 ( .A(n2103), .ZN(n2102) );
  INV_X1 U2678 ( .A(n4113), .ZN(n4770) );
  NAND2_X1 U2679 ( .A1(n2807), .A2(n2806), .ZN(n3740) );
  INV_X1 U2680 ( .A(n2811), .ZN(n4027) );
  INV_X1 U2681 ( .A(n3968), .ZN(n4140) );
  NAND2_X1 U2682 ( .A1(n2704), .A2(n2703), .ZN(n4143) );
  OR2_X1 U2683 ( .A1(n3085), .A2(n2777), .ZN(n2704) );
  INV_X1 U2684 ( .A(n4337), .ZN(n4350) );
  NAND2_X1 U2685 ( .A1(n2158), .A2(n2157), .ZN(n4147) );
  NAND2_X1 U2686 ( .A1(n2154), .A2(n2153), .ZN(n2158) );
  INV_X1 U2687 ( .A(n4378), .ZN(n4210) );
  NAND2_X1 U2688 ( .A1(n2154), .A2(n2159), .ZN(n4172) );
  INV_X1 U2689 ( .A(n4415), .ZN(n4277) );
  INV_X1 U2690 ( .A(n4450), .ZN(n3854) );
  NAND2_X1 U2691 ( .A1(n2146), .A2(n2025), .ZN(n3644) );
  OR2_X1 U2692 ( .A1(n3636), .A2(n2562), .ZN(n2146) );
  NAND2_X1 U2693 ( .A1(n2138), .A2(n2533), .ZN(n3559) );
  NAND2_X1 U2694 ( .A1(n2714), .A2(n2713), .ZN(n3523) );
  NAND2_X1 U2695 ( .A1(n4323), .A2(n4640), .ZN(n4342) );
  OR2_X1 U2696 ( .A1(n4788), .A2(n3373), .ZN(n4361) );
  NAND2_X1 U2697 ( .A1(n2164), .A2(n2170), .ZN(n3407) );
  INV_X1 U2698 ( .A(n2832), .ZN(n3330) );
  OR2_X1 U2699 ( .A1(n4788), .A2(n4390), .ZN(n4356) );
  NAND2_X1 U2700 ( .A1(n3216), .A2(n3097), .ZN(n4792) );
  OR2_X1 U2701 ( .A1(n3125), .A2(n3305), .ZN(n4804) );
  INV_X1 U2702 ( .A(n3179), .ZN(n4713) );
  AND2_X1 U2703 ( .A1(n2363), .A2(STATE_REG_SCAN_IN), .ZN(n4805) );
  INV_X1 U2704 ( .A(n4063), .ZN(n4717) );
  INV_X1 U2705 ( .A(n3662), .ZN(n3659) );
  XNOR2_X1 U2706 ( .A(n2269), .B(IR_REG_8__SCAN_IN), .ZN(n4721) );
  AND2_X1 U2707 ( .A1(n2268), .A2(n2266), .ZN(n4722) );
  INV_X1 U2708 ( .A(IR_REG_3__SCAN_IN), .ZN(n2251) );
  AOI21_X1 U2710 ( .B1(n2129), .B2(n4096), .A(n2127), .ZN(n4112) );
  OR2_X1 U2711 ( .A1(n4828), .A2(REG1_REG_29__SCAN_IN), .ZN(n2183) );
  NAND2_X1 U2712 ( .A1(n2140), .A2(n2139), .ZN(n2820) );
  OR2_X1 U2713 ( .A1(n4824), .A2(REG0_REG_29__SCAN_IN), .ZN(n2139) );
  OR2_X1 U2714 ( .A1(n4123), .A2(n4706), .ZN(n2795) );
  NAND2_X1 U2715 ( .A1(n2648), .A2(n4222), .ZN(n4185) );
  AND2_X1 U2716 ( .A1(n2028), .A2(n3645), .ZN(n2025) );
  INV_X1 U2717 ( .A(n3157), .ZN(n2095) );
  AND2_X1 U2718 ( .A1(n2974), .A2(n2190), .ZN(n2026) );
  AND2_X1 U2719 ( .A1(n2185), .A2(n2728), .ZN(n2027) );
  INV_X1 U2720 ( .A(n4762), .ZN(n4096) );
  NAND2_X1 U2721 ( .A1(n3408), .A2(n3418), .ZN(n3409) );
  NAND2_X1 U2722 ( .A1(n4474), .A2(n3627), .ZN(n2028) );
  OR2_X1 U2723 ( .A1(n2413), .A2(n4739), .ZN(n2029) );
  NAND2_X1 U2724 ( .A1(n4736), .A2(REG1_REG_14__SCAN_IN), .ZN(n4735) );
  NOR2_X1 U2725 ( .A1(n4757), .A2(REG1_REG_16__SCAN_IN), .ZN(n4756) );
  AND2_X1 U2726 ( .A1(n2948), .A2(n2947), .ZN(n2030) );
  INV_X1 U2727 ( .A(n3464), .ZN(n2070) );
  NAND2_X1 U2728 ( .A1(n2732), .A2(n4039), .ZN(n4183) );
  OR2_X1 U2729 ( .A1(n4372), .A2(n4706), .ZN(n2031) );
  OR2_X1 U2730 ( .A1(n2736), .A2(n2689), .ZN(n2032) );
  NAND2_X1 U2731 ( .A1(n4347), .A2(n2185), .ZN(n4268) );
  NOR2_X1 U2732 ( .A1(n4357), .A2(n2627), .ZN(n2033) );
  NOR2_X1 U2733 ( .A1(n4756), .A2(n2319), .ZN(n4103) );
  NOR2_X1 U2734 ( .A1(n4045), .A2(n2783), .ZN(n2034) );
  NAND2_X1 U2735 ( .A1(n3447), .A2(n3411), .ZN(n2035) );
  INV_X1 U2736 ( .A(n3163), .ZN(n4724) );
  AND2_X1 U2737 ( .A1(n2795), .A2(n2794), .ZN(n2036) );
  NAND3_X1 U2738 ( .A1(n2193), .A2(n2081), .A3(n2233), .ZN(n2248) );
  NAND2_X1 U2739 ( .A1(n3485), .A2(n2222), .ZN(n2282) );
  AND2_X1 U2740 ( .A1(n3583), .A2(n3585), .ZN(n3991) );
  AND2_X1 U2741 ( .A1(REG3_REG_6__SCAN_IN), .A2(REG3_REG_7__SCAN_IN), .ZN(
        n2037) );
  NOR2_X1 U2742 ( .A1(n4137), .A2(n4154), .ZN(n2038) );
  AND2_X1 U2743 ( .A1(n2125), .A2(n2029), .ZN(n2039) );
  AND2_X1 U2744 ( .A1(n4214), .A2(n4216), .ZN(n4191) );
  NAND2_X1 U2745 ( .A1(n4753), .A2(n4752), .ZN(n4751) );
  INV_X1 U2746 ( .A(n2062), .ZN(n2674) );
  NOR2_X1 U2747 ( .A1(n2666), .A2(n3719), .ZN(n2062) );
  AND2_X1 U2748 ( .A1(n4210), .A2(n4195), .ZN(n2040) );
  INV_X1 U2749 ( .A(IR_REG_1__SCAN_IN), .ZN(n2193) );
  NOR2_X1 U2750 ( .A1(n4244), .A2(n4232), .ZN(n4214) );
  INV_X1 U2751 ( .A(n3439), .ZN(n2198) );
  OR2_X1 U2752 ( .A1(n4387), .A2(n4377), .ZN(n2041) );
  AND2_X1 U2753 ( .A1(n2807), .A2(n2181), .ZN(n2042) );
  NOR2_X1 U2754 ( .A1(n4719), .A2(n2111), .ZN(n2043) );
  AND2_X1 U2755 ( .A1(n2216), .A2(n2432), .ZN(n2044) );
  AND2_X1 U2756 ( .A1(n3838), .A2(n2214), .ZN(n2045) );
  INV_X1 U2757 ( .A(IR_REG_26__SCAN_IN), .ZN(n2367) );
  NAND2_X1 U2758 ( .A1(n3310), .A2(n4792), .ZN(n4334) );
  INV_X1 U2759 ( .A(n4334), .ZN(n4788) );
  CLKBUF_X1 U2760 ( .A(IR_REG_0__SCAN_IN), .Z(n4729) );
  OAI21_X1 U2761 ( .B1(n2714), .B2(n2179), .A(n2177), .ZN(n3556) );
  OR2_X1 U2762 ( .A1(n2315), .A2(n4748), .ZN(n2046) );
  NAND2_X1 U2763 ( .A1(n2016), .A2(n2070), .ZN(n2047) );
  XNOR2_X1 U2764 ( .A(n2282), .B(n3477), .ZN(n3474) );
  NAND2_X1 U2765 ( .A1(n2200), .A2(n2199), .ZN(n3438) );
  OAI211_X1 U2766 ( .C1(n4090), .C2(n4718), .A(n2089), .B(n2092), .ZN(n3597)
         );
  INV_X1 U2767 ( .A(n3936), .ZN(n2169) );
  INV_X1 U2768 ( .A(n3952), .ZN(n2186) );
  AND2_X1 U2769 ( .A1(n2181), .A2(n4828), .ZN(n2048) );
  NOR2_X1 U2770 ( .A1(n2093), .A2(n2090), .ZN(n2049) );
  NAND2_X1 U2771 ( .A1(n2284), .A2(n2283), .ZN(n4087) );
  AND2_X1 U2772 ( .A1(n2046), .A2(REG1_REG_14__SCAN_IN), .ZN(n2050) );
  INV_X1 U2773 ( .A(n2960), .ZN(n2191) );
  AND2_X1 U2774 ( .A1(n3854), .A2(n3756), .ZN(n2051) );
  AND2_X1 U2775 ( .A1(n2291), .A2(REG1_REG_11__SCAN_IN), .ZN(n2052) );
  AND2_X1 U2776 ( .A1(n4722), .A2(REG1_REG_7__SCAN_IN), .ZN(n2053) );
  INV_X1 U2777 ( .A(n2973), .ZN(n2192) );
  AND2_X1 U2778 ( .A1(n3686), .A2(n2226), .ZN(n4298) );
  AND2_X1 U2779 ( .A1(n2146), .A2(n2028), .ZN(n2054) );
  AND4_X1 U2780 ( .A1(n2473), .A2(n2472), .A3(n2471), .A4(n2470), .ZN(n3390)
         );
  NAND3_X1 U2781 ( .A1(n3287), .A2(n3289), .A3(n3286), .ZN(n3288) );
  AND2_X2 U2782 ( .A1(n2787), .A2(n3072), .ZN(n4828) );
  INV_X1 U2783 ( .A(n4828), .ZN(n4825) );
  AND2_X2 U2784 ( .A1(n2787), .A2(n3309), .ZN(n4824) );
  INV_X1 U2785 ( .A(IR_REG_15__SCAN_IN), .ZN(n2067) );
  NAND2_X1 U2786 ( .A1(n2188), .A2(IR_REG_31__SCAN_IN), .ZN(n2366) );
  OR2_X1 U2787 ( .A1(n2370), .A2(n2369), .ZN(n2055) );
  INV_X1 U2788 ( .A(n3068), .ZN(n4129) );
  AND2_X1 U2789 ( .A1(n4277), .A2(n4245), .ZN(n2056) );
  INV_X1 U2790 ( .A(n3409), .ZN(n2770) );
  INV_X1 U2791 ( .A(n3335), .ZN(n2071) );
  AND2_X1 U2792 ( .A1(n2047), .A2(n3921), .ZN(n2057) );
  INV_X1 U2793 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2111) );
  AND2_X1 U2794 ( .A1(n2099), .A2(n2257), .ZN(n2058) );
  NAND3_X1 U2795 ( .A1(n2798), .A2(n2797), .A3(n3964), .ZN(n2799) );
  OAI21_X2 U2796 ( .B1(n4161), .B2(n2777), .A(n2679), .ZN(n4137) );
  NAND4_X1 U2797 ( .A1(n2338), .A2(n2066), .A3(n2065), .A4(n2064), .ZN(n2350)
         );
  NOR2_X2 U2798 ( .A1(n3335), .A2(n2069), .ZN(n3408) );
  NAND2_X4 U2799 ( .A1(n2073), .A2(n2072), .ZN(n3694) );
  NAND2_X1 U2800 ( .A1(n2586), .A2(REG3_REG_19__SCAN_IN), .ZN(n2596) );
  INV_X1 U2801 ( .A(n3362), .ZN(n2768) );
  NAND2_X1 U2802 ( .A1(n3270), .A2(REG1_REG_8__SCAN_IN), .ZN(n2273) );
  NAND2_X1 U2803 ( .A1(n4080), .A2(n4079), .ZN(n4078) );
  OAI211_X1 U2804 ( .C1(n4090), .C2(n2088), .A(n2085), .B(n2086), .ZN(n2306)
         );
  INV_X1 U2805 ( .A(n2306), .ZN(n3658) );
  NAND2_X1 U2806 ( .A1(n2258), .A2(n2095), .ZN(n2094) );
  INV_X1 U2807 ( .A(n2099), .ZN(n3254) );
  INV_X1 U2808 ( .A(n4103), .ZN(n2106) );
  NAND2_X1 U2809 ( .A1(n2100), .A2(n2102), .ZN(n2337) );
  NAND2_X1 U2810 ( .A1(n4103), .A2(n2101), .ZN(n2100) );
  NOR2_X1 U2811 ( .A1(n4104), .A2(n2329), .ZN(n4771) );
  NAND2_X1 U2812 ( .A1(n2108), .A2(n2043), .ZN(n2107) );
  NAND3_X1 U2813 ( .A1(n2406), .A2(n2110), .A3(n2107), .ZN(n4099) );
  NAND2_X1 U2814 ( .A1(n2404), .A2(n2109), .ZN(n2110) );
  NAND2_X1 U2815 ( .A1(n2115), .A2(n2112), .ZN(n3475) );
  NAND2_X1 U2816 ( .A1(n2404), .A2(n2403), .ZN(n2405) );
  INV_X1 U2817 ( .A(n2403), .ZN(n2114) );
  OAI21_X1 U2818 ( .B1(n2120), .B2(n3249), .A(n2116), .ZN(n3158) );
  NAND2_X1 U2819 ( .A1(n3598), .A2(REG2_REG_12__SCAN_IN), .ZN(n2123) );
  AND2_X2 U2820 ( .A1(n2126), .A2(n2029), .ZN(n4742) );
  NAND2_X1 U2821 ( .A1(n2578), .A2(n2131), .ZN(n4241) );
  NAND2_X1 U2822 ( .A1(n4241), .A2(n2638), .ZN(n2640) );
  NOR2_X2 U2823 ( .A1(n2133), .A2(n2132), .ZN(n4360) );
  INV_X1 U2824 ( .A(n4360), .ZN(n4256) );
  AND2_X2 U2825 ( .A1(n2439), .A2(n2440), .ZN(n2469) );
  NAND2_X1 U2826 ( .A1(n2135), .A2(n2489), .ZN(n3406) );
  NAND3_X1 U2827 ( .A1(n2042), .A2(n4824), .A3(n2141), .ZN(n2140) );
  NAND2_X1 U2828 ( .A1(n3636), .A2(n2025), .ZN(n2144) );
  NAND2_X1 U2829 ( .A1(n2144), .A2(n2145), .ZN(n3684) );
  NAND2_X1 U2830 ( .A1(n4185), .A2(n2149), .ZN(n2148) );
  NOR2_X1 U2831 ( .A1(n2229), .A2(n2040), .ZN(n2159) );
  NAND2_X1 U2832 ( .A1(n3913), .A2(n3909), .ZN(n3231) );
  NAND2_X1 U2833 ( .A1(n2161), .A2(n3950), .ZN(n3683) );
  NAND2_X1 U2834 ( .A1(n3643), .A2(n3993), .ZN(n2161) );
  NAND3_X1 U2835 ( .A1(n2165), .A2(n3923), .A3(n2162), .ZN(n3445) );
  NAND2_X1 U2836 ( .A1(n3343), .A2(n2057), .ZN(n2164) );
  NAND2_X1 U2837 ( .A1(n3343), .A2(n2166), .ZN(n2165) );
  NAND2_X1 U2838 ( .A1(n3936), .A2(n3921), .ZN(n2167) );
  OAI21_X1 U2839 ( .B1(n3343), .B2(n2173), .A(n3921), .ZN(n3367) );
  NAND2_X1 U2840 ( .A1(n2173), .A2(n3921), .ZN(n2172) );
  NAND2_X1 U2841 ( .A1(n2714), .A2(n2177), .ZN(n2174) );
  NAND2_X1 U2842 ( .A1(n2174), .A2(n2175), .ZN(n2721) );
  NAND2_X1 U2843 ( .A1(n4347), .A2(n2027), .ZN(n2184) );
  INV_X1 U2844 ( .A(n4168), .ZN(n4150) );
  NAND3_X1 U2845 ( .A1(n2352), .A2(n2351), .A3(n2367), .ZN(n2188) );
  NAND2_X1 U2846 ( .A1(n3774), .A2(n2985), .ZN(n2995) );
  NAND2_X1 U2847 ( .A1(n3399), .A2(n2195), .ZN(n2194) );
  NAND2_X1 U2848 ( .A1(n3673), .A2(n2914), .ZN(n3619) );
  NAND2_X1 U2849 ( .A1(n2206), .A2(n2920), .ZN(n3793) );
  NAND3_X1 U2850 ( .A1(n2920), .A2(n2206), .A3(n2205), .ZN(n2204) );
  NAND2_X1 U2851 ( .A1(n3673), .A2(n2208), .ZN(n2207) );
  NAND2_X1 U2852 ( .A1(n3839), .A2(n2212), .ZN(n2211) );
  NAND2_X1 U2853 ( .A1(n3839), .A2(n3840), .ZN(n3838) );
  NAND2_X1 U2854 ( .A1(n2217), .A2(n2044), .ZN(n2436) );
  INV_X1 U2855 ( .A(n2370), .ZN(n2217) );
  NAND2_X1 U2856 ( .A1(n2413), .A2(n4739), .ZN(n2414) );
  AOI21_X1 U2857 ( .B1(n4761), .B2(n4763), .A(n4762), .ZN(n4768) );
  AOI21_X1 U2858 ( .B1(n4119), .B2(n4118), .A(n4117), .ZN(n4651) );
  NAND2_X1 U2859 ( .A1(n4118), .A2(n2818), .ZN(n3742) );
  OR2_X1 U2860 ( .A1(n4256), .A2(n4357), .ZN(n4358) );
  AND2_X1 U2861 ( .A1(n3694), .A2(DATAI_26_), .ZN(n4154) );
  AND2_X1 U2862 ( .A1(n3694), .A2(DATAI_25_), .ZN(n4377) );
  AND2_X1 U2863 ( .A1(n3694), .A2(DATAI_21_), .ZN(n4404) );
  NAND2_X1 U2864 ( .A1(n2023), .A2(DATAI_1_), .ZN(n2446) );
  AND4_X1 U2865 ( .A1(n2452), .A2(n2450), .A3(n2451), .A4(n2449), .ZN(n2448)
         );
  NOR2_X1 U2866 ( .A1(n4740), .A2(n2416), .ZN(n2417) );
  NAND2_X1 U2867 ( .A1(n2384), .A2(n2383), .ZN(n2382) );
  NAND2_X1 U2868 ( .A1(n2384), .A2(n2245), .ZN(n2246) );
  CLKBUF_X1 U2869 ( .A(n3774), .Z(n3874) );
  OR2_X1 U2870 ( .A1(n2260), .A2(n3170), .ZN(n2220) );
  NAND2_X1 U2871 ( .A1(n4106), .A2(n2421), .ZN(n4761) );
  OR2_X1 U2872 ( .A1(n4808), .A2(n4580), .ZN(n2221) );
  OR2_X1 U2873 ( .A1(n2279), .A2(n2277), .ZN(n2222) );
  INV_X1 U2874 ( .A(IR_REG_28__SCAN_IN), .ZN(n2372) );
  INV_X1 U2875 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2245) );
  NAND2_X1 U2876 ( .A1(n2344), .A2(IR_REG_31__SCAN_IN), .ZN(n2355) );
  NOR2_X1 U2877 ( .A1(n3433), .A2(n2873), .ZN(n2223) );
  AND2_X1 U2878 ( .A1(n2993), .A2(n2992), .ZN(n2224) );
  AND2_X1 U2879 ( .A1(n2798), .A2(n2797), .ZN(n2225) );
  NOR2_X1 U2880 ( .A1(n4308), .A2(n4313), .ZN(n2226) );
  NOR2_X1 U2881 ( .A1(n2990), .A2(n3872), .ZN(n2227) );
  AND2_X1 U2882 ( .A1(n3714), .A2(n3041), .ZN(n2228) );
  NAND2_X1 U2883 ( .A1(n2292), .A2(n2288), .ZN(n2542) );
  INV_X1 U2884 ( .A(n2542), .ZN(n2291) );
  NOR2_X1 U2885 ( .A1(n2664), .A2(n4187), .ZN(n2229) );
  AND2_X1 U2886 ( .A1(n3104), .A2(n3876), .ZN(n2230) );
  INV_X1 U2887 ( .A(n4052), .ZN(n2689) );
  INV_X1 U2888 ( .A(n3733), .ZN(n2776) );
  INV_X1 U2889 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2383) );
  INV_X1 U2890 ( .A(n4308), .ZN(n4315) );
  AND3_X1 U2891 ( .A1(n3998), .A2(n2509), .A3(n3451), .ZN(n2231) );
  NOR2_X1 U2892 ( .A1(n4349), .A2(n4352), .ZN(n2232) );
  INV_X1 U2893 ( .A(IR_REG_22__SCAN_IN), .ZN(n2347) );
  INV_X1 U2894 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2420) );
  OR2_X1 U2895 ( .A1(n3324), .A2(n3035), .ZN(n2827) );
  AND3_X1 U2896 ( .A1(n2970), .A2(n2969), .A3(n3817), .ZN(n2974) );
  AND2_X1 U2897 ( .A1(n2575), .A2(REG2_REG_15__SCAN_IN), .ZN(n2416) );
  NAND2_X1 U2898 ( .A1(n3293), .A2(n3912), .ZN(n3355) );
  NAND2_X1 U2899 ( .A1(n2705), .A2(n3927), .ZN(n3998) );
  OR2_X1 U2900 ( .A1(n2322), .A2(IR_REG_14__SCAN_IN), .ZN(n2310) );
  NOR2_X1 U2901 ( .A1(n2227), .A2(n2224), .ZN(n2994) );
  INV_X1 U2902 ( .A(n3676), .ZN(n2908) );
  NAND2_X1 U2903 ( .A1(n4082), .A2(n2381), .ZN(n3187) );
  NAND2_X1 U2904 ( .A1(n2608), .A2(REG2_REG_18__SCAN_IN), .ZN(n2423) );
  OR2_X1 U2905 ( .A1(n4247), .A2(n3867), .ZN(n4204) );
  NAND2_X1 U2906 ( .A1(n3557), .A2(n2543), .ZN(n3587) );
  OR2_X1 U2907 ( .A1(n2712), .A2(n2711), .ZN(n2713) );
  INV_X1 U2908 ( .A(n3289), .ZN(n3988) );
  INV_X1 U2909 ( .A(REG3_REG_11__SCAN_IN), .ZN(n4521) );
  NAND2_X1 U2910 ( .A1(n2372), .A2(IR_REG_27__SCAN_IN), .ZN(n2364) );
  INV_X1 U2911 ( .A(n3456), .ZN(n2769) );
  INV_X1 U2912 ( .A(IR_REG_21__SCAN_IN), .ZN(n4492) );
  OAI21_X1 U2913 ( .B1(n2285), .B2(IR_REG_10__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2287) );
  XNOR2_X1 U2914 ( .A(n2843), .B(n3051), .ZN(n2847) );
  INV_X1 U2915 ( .A(n4432), .ZN(n4452) );
  OR2_X1 U2916 ( .A1(n4248), .A2(n2777), .ZN(n2636) );
  AOI21_X1 U2917 ( .B1(n4765), .B2(ADDR_REG_18__SCAN_IN), .A(n4764), .ZN(n4766) );
  AND2_X1 U2918 ( .A1(n4003), .A2(n4202), .ZN(n4243) );
  INV_X1 U2919 ( .A(n4440), .ZN(n4463) );
  INV_X1 U2920 ( .A(n3621), .ZN(n3566) );
  INV_X1 U2921 ( .A(n3411), .ZN(n3418) );
  OR2_X1 U2922 ( .A1(n4788), .A2(n4477), .ZN(n4336) );
  AND2_X1 U2923 ( .A1(n3694), .A2(DATAI_22_), .ZN(n4232) );
  INV_X1 U2924 ( .A(n4261), .ZN(n4320) );
  NAND2_X1 U2925 ( .A1(n3075), .A2(n3179), .ZN(n4462) );
  NAND2_X1 U2926 ( .A1(n2357), .A2(n4492), .ZN(n2361) );
  OR2_X1 U2927 ( .A1(n2302), .A2(n2301), .ZN(n3662) );
  AND2_X1 U2928 ( .A1(n3105), .A2(n2230), .ZN(n3084) );
  INV_X1 U2929 ( .A(n3907), .ZN(n3876) );
  INV_X1 U2930 ( .A(n4356), .ZN(n4340) );
  NOR2_X1 U2931 ( .A1(n4365), .A2(n4717), .ZN(n4323) );
  AND2_X1 U2932 ( .A1(n4033), .A2(n3952), .ZN(n4357) );
  INV_X1 U2933 ( .A(n4361), .ZN(n4344) );
  INV_X1 U2934 ( .A(n4342), .ZN(n4779) );
  AOI21_X1 U2935 ( .B1(n3125), .B2(n3129), .A(n2766), .ZN(n3072) );
  INV_X1 U2936 ( .A(n3686), .ZN(n4349) );
  INV_X1 U2937 ( .A(n4459), .ZN(n3756) );
  AND3_X1 U2938 ( .A1(n2765), .A2(n2764), .A3(n3071), .ZN(n2787) );
  NAND2_X1 U2939 ( .A1(n2824), .A2(n4805), .ZN(n3305) );
  AND2_X1 U2940 ( .A1(n2312), .A2(n2316), .ZN(n2575) );
  AND2_X1 U2941 ( .A1(n2376), .A2(n2375), .ZN(n4765) );
  AND2_X1 U2942 ( .A1(n3098), .A2(n4792), .ZN(n3900) );
  AND2_X1 U2943 ( .A1(n3095), .A2(n3094), .ZN(n3886) );
  NAND2_X1 U2944 ( .A1(n2782), .A2(n2781), .ZN(n4125) );
  NAND2_X1 U2945 ( .A1(n2653), .A2(n2652), .ZN(n4224) );
  CLKBUF_X2 U2946 ( .A(U4043), .Z(n4077) );
  OR2_X1 U2947 ( .A1(n3152), .A2(n2428), .ZN(n4762) );
  OR2_X1 U2948 ( .A1(n3152), .A2(n4065), .ZN(n4113) );
  INV_X2 U2949 ( .A(n4334), .ZN(n4365) );
  OR2_X1 U2950 ( .A1(n3742), .A2(n4484), .ZN(n2821) );
  OR2_X1 U2951 ( .A1(n3742), .A2(n4706), .ZN(n2819) );
  INV_X1 U2952 ( .A(n4824), .ZN(n4822) );
  INV_X1 U2953 ( .A(n4804), .ZN(n4803) );
  INV_X1 U2954 ( .A(n2694), .ZN(n4716) );
  XNOR2_X1 U2955 ( .A(n2276), .B(IR_REG_9__SCAN_IN), .ZN(n4720) );
  OAI21_X1 U2956 ( .B1(n2796), .B2(n4825), .A(n2792), .ZN(U3546) );
  OAI21_X1 U2957 ( .B1(n2796), .B2(n4822), .A(n2036), .ZN(U3514) );
  INV_X2 U2958 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U2959 ( .A(n2248), .ZN(n2235) );
  NAND2_X1 U2960 ( .A1(n2236), .A2(IR_REG_31__SCAN_IN), .ZN(n2237) );
  MUX2_X1 U2961 ( .A(IR_REG_31__SCAN_IN), .B(n2237), .S(IR_REG_5__SCAN_IN), 
        .Z(n2240) );
  INV_X1 U2962 ( .A(n2236), .ZN(n2239) );
  NAND2_X1 U2963 ( .A1(n2240), .A2(n2261), .ZN(n3163) );
  INV_X1 U2964 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2241) );
  AND2_X1 U2965 ( .A1(n4729), .A2(REG1_REG_0__SCAN_IN), .ZN(n4079) );
  NAND2_X1 U2966 ( .A1(n4728), .A2(REG1_REG_1__SCAN_IN), .ZN(n2242) );
  NAND2_X1 U2967 ( .A1(n3184), .A2(n3185), .ZN(n3183) );
  NAND2_X1 U2968 ( .A1(n2248), .A2(IR_REG_31__SCAN_IN), .ZN(n2252) );
  XNOR2_X1 U2969 ( .A(n2252), .B(IR_REG_3__SCAN_IN), .ZN(n4726) );
  INV_X1 U2970 ( .A(n4726), .ZN(n3147) );
  INV_X1 U2971 ( .A(REG1_REG_3__SCAN_IN), .ZN(n3142) );
  NAND2_X1 U2972 ( .A1(n2252), .A2(n2251), .ZN(n2253) );
  NAND2_X1 U2973 ( .A1(n2253), .A2(IR_REG_31__SCAN_IN), .ZN(n2254) );
  XNOR2_X1 U2974 ( .A(n2254), .B(IR_REG_4__SCAN_IN), .ZN(n4725) );
  INV_X1 U2975 ( .A(n4725), .ZN(n3253) );
  XNOR2_X1 U2976 ( .A(n2255), .B(n3253), .ZN(n3255) );
  INV_X1 U2977 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4826) );
  INV_X1 U2978 ( .A(n2255), .ZN(n2256) );
  NAND2_X1 U2979 ( .A1(n2256), .A2(n4725), .ZN(n2257) );
  INV_X1 U2980 ( .A(n2257), .ZN(n2258) );
  XNOR2_X1 U2981 ( .A(n4724), .B(REG1_REG_5__SCAN_IN), .ZN(n3157) );
  NAND2_X1 U2982 ( .A1(n2261), .A2(IR_REG_31__SCAN_IN), .ZN(n2259) );
  XNOR2_X1 U2983 ( .A(n2259), .B(IR_REG_6__SCAN_IN), .ZN(n4723) );
  XNOR2_X1 U2984 ( .A(n2260), .B(n4723), .ZN(n3169) );
  INV_X1 U2985 ( .A(n4723), .ZN(n3170) );
  INV_X1 U2986 ( .A(n2261), .ZN(n2263) );
  NAND2_X1 U2987 ( .A1(n2263), .A2(n2262), .ZN(n2275) );
  NAND2_X1 U2988 ( .A1(n2275), .A2(IR_REG_31__SCAN_IN), .ZN(n2265) );
  NAND2_X1 U2989 ( .A1(n2265), .A2(n2264), .ZN(n2268) );
  OR2_X1 U2990 ( .A1(n2265), .A2(n2264), .ZN(n2266) );
  INV_X1 U2991 ( .A(n4722), .ZN(n3205) );
  INV_X1 U2992 ( .A(REG1_REG_7__SCAN_IN), .ZN(n3202) );
  NAND2_X1 U2993 ( .A1(n3205), .A2(n3202), .ZN(n2267) );
  NAND2_X1 U2994 ( .A1(n2268), .A2(IR_REG_31__SCAN_IN), .ZN(n2269) );
  INV_X1 U2995 ( .A(n2270), .ZN(n2271) );
  NAND2_X1 U2996 ( .A1(n2271), .A2(n4721), .ZN(n2272) );
  NAND2_X1 U2997 ( .A1(n2273), .A2(n2272), .ZN(n3484) );
  INV_X1 U2998 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2277) );
  NOR2_X2 U2999 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2297)
         );
  INV_X1 U3000 ( .A(n2297), .ZN(n2274) );
  NAND2_X1 U3001 ( .A1(n2280), .A2(IR_REG_31__SCAN_IN), .ZN(n2276) );
  MUX2_X1 U3002 ( .A(n2277), .B(REG1_REG_9__SCAN_IN), .S(n4720), .Z(n3487) );
  NAND2_X1 U3003 ( .A1(n3484), .A2(n2278), .ZN(n3485) );
  INV_X1 U3004 ( .A(n4720), .ZN(n2279) );
  NAND2_X1 U3005 ( .A1(n2285), .A2(IR_REG_31__SCAN_IN), .ZN(n2281) );
  XNOR2_X1 U3006 ( .A(n2281), .B(IR_REG_10__SCAN_IN), .ZN(n4719) );
  INV_X1 U3007 ( .A(n4719), .ZN(n3477) );
  INV_X1 U3008 ( .A(REG1_REG_11__SCAN_IN), .ZN(n2289) );
  NAND2_X1 U3009 ( .A1(n2287), .A2(n2286), .ZN(n2292) );
  OR2_X1 U3010 ( .A1(n2287), .A2(n2286), .ZN(n2288) );
  MUX2_X1 U3011 ( .A(REG1_REG_11__SCAN_IN), .B(n2289), .S(n2542), .Z(n4088) );
  NAND2_X1 U3012 ( .A1(n2292), .A2(IR_REG_31__SCAN_IN), .ZN(n2293) );
  XNOR2_X1 U3013 ( .A(n2293), .B(IR_REG_12__SCAN_IN), .ZN(n4718) );
  INV_X1 U3014 ( .A(n4718), .ZN(n3601) );
  NOR2_X1 U3015 ( .A1(n2352), .A2(n2080), .ZN(n2300) );
  MUX2_X1 U3016 ( .A(n2080), .B(n2300), .S(IR_REG_13__SCAN_IN), .Z(n2302) );
  NAND2_X1 U3017 ( .A1(n2352), .A2(n4496), .ZN(n2322) );
  INV_X1 U3018 ( .A(n2322), .ZN(n2301) );
  INV_X1 U3019 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4471) );
  NAND2_X1 U3020 ( .A1(n3662), .A2(n4471), .ZN(n2303) );
  OAI21_X1 U3021 ( .B1(n3662), .B2(n4471), .A(n2303), .ZN(n2304) );
  INV_X1 U3022 ( .A(n2304), .ZN(n2305) );
  NAND2_X1 U3023 ( .A1(n2306), .A2(n2305), .ZN(n3660) );
  NAND2_X1 U3024 ( .A1(n3659), .A2(REG1_REG_13__SCAN_IN), .ZN(n2307) );
  NAND2_X1 U3025 ( .A1(n2322), .A2(IR_REG_31__SCAN_IN), .ZN(n2308) );
  XNOR2_X1 U3026 ( .A(n2308), .B(IR_REG_14__SCAN_IN), .ZN(n4813) );
  INV_X1 U3027 ( .A(n4813), .ZN(n4739) );
  NAND2_X1 U3028 ( .A1(n4813), .A2(n2309), .ZN(n4745) );
  NAND2_X1 U3029 ( .A1(n2310), .A2(IR_REG_31__SCAN_IN), .ZN(n2311) );
  OR2_X1 U3030 ( .A1(n2311), .A2(n2067), .ZN(n2312) );
  NAND2_X1 U3031 ( .A1(n2311), .A2(n2067), .ZN(n2316) );
  NAND2_X1 U3032 ( .A1(REG1_REG_15__SCAN_IN), .A2(n2575), .ZN(n2313) );
  INV_X1 U3033 ( .A(n2313), .ZN(n2315) );
  INV_X1 U3034 ( .A(n2575), .ZN(n4812) );
  INV_X1 U3035 ( .A(REG1_REG_15__SCAN_IN), .ZN(n2314) );
  AOI22_X1 U3036 ( .A1(REG1_REG_15__SCAN_IN), .A2(n2575), .B1(n4812), .B2(
        n2314), .ZN(n4748) );
  NAND2_X1 U3037 ( .A1(n2316), .A2(IR_REG_31__SCAN_IN), .ZN(n2317) );
  XNOR2_X1 U3038 ( .A(n2317), .B(IR_REG_16__SCAN_IN), .ZN(n2585) );
  INV_X1 U3039 ( .A(n2585), .ZN(n4810) );
  NOR2_X1 U3040 ( .A1(n2585), .A2(n2318), .ZN(n2319) );
  INV_X1 U3041 ( .A(IR_REG_16__SCAN_IN), .ZN(n2320) );
  NAND2_X1 U3042 ( .A1(n2338), .A2(n2320), .ZN(n2321) );
  OAI21_X1 U3043 ( .B1(n2322), .B2(n2321), .A(IR_REG_31__SCAN_IN), .ZN(n2323)
         );
  MUX2_X1 U3044 ( .A(IR_REG_31__SCAN_IN), .B(n2323), .S(IR_REG_17__SCAN_IN), 
        .Z(n2327) );
  NOR2_X1 U3045 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2325)
         );
  INV_X1 U3046 ( .A(IR_REG_14__SCAN_IN), .ZN(n2324) );
  NAND2_X1 U3047 ( .A1(n2352), .A2(n2326), .ZN(n2331) );
  AND2_X1 U3048 ( .A1(n2327), .A2(n2331), .ZN(n4109) );
  INV_X1 U3049 ( .A(n4109), .ZN(n2419) );
  NOR2_X1 U3050 ( .A1(n4109), .A2(REG1_REG_17__SCAN_IN), .ZN(n2329) );
  INV_X1 U3051 ( .A(n2329), .ZN(n2328) );
  OAI21_X1 U3052 ( .B1(n4438), .B2(n2419), .A(n2328), .ZN(n4105) );
  NAND2_X1 U3053 ( .A1(n2331), .A2(IR_REG_31__SCAN_IN), .ZN(n2330) );
  XNOR2_X1 U3054 ( .A(n2330), .B(IR_REG_18__SCAN_IN), .ZN(n2608) );
  INV_X1 U3055 ( .A(n2608), .ZN(n4808) );
  INV_X1 U3056 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4580) );
  AOI22_X1 U3057 ( .A1(REG1_REG_18__SCAN_IN), .A2(n2608), .B1(n4808), .B2(
        n4580), .ZN(n4772) );
  INV_X1 U3058 ( .A(REG1_REG_19__SCAN_IN), .ZN(n2335) );
  MUX2_X1 U3059 ( .A(REG1_REG_19__SCAN_IN), .B(n2335), .S(n4063), .Z(n2336) );
  XNOR2_X1 U3060 ( .A(n2337), .B(n2336), .ZN(n2379) );
  INV_X1 U3061 ( .A(n2350), .ZN(n2339) );
  INV_X1 U3062 ( .A(n2361), .ZN(n2340) );
  NAND2_X1 U3063 ( .A1(n2340), .A2(n2347), .ZN(n2344) );
  NAND2_X1 U3064 ( .A1(n2355), .A2(n2356), .ZN(n2341) );
  NAND2_X1 U3065 ( .A1(n2356), .A2(n2346), .ZN(n2343) );
  OAI21_X1 U3066 ( .B1(n2344), .B2(n2343), .A(IR_REG_31__SCAN_IN), .ZN(n2345)
         );
  MUX2_X1 U3067 ( .A(IR_REG_31__SCAN_IN), .B(n2345), .S(IR_REG_25__SCAN_IN), 
        .Z(n2353) );
  NOR2_X1 U3068 ( .A1(IR_REG_23__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .ZN(n2348)
         );
  NAND4_X1 U3069 ( .A1(n2348), .A2(n2347), .A3(n2346), .A4(n4492), .ZN(n2349)
         );
  NAND2_X1 U3070 ( .A1(n2370), .A2(IR_REG_31__SCAN_IN), .ZN(n2354) );
  NAND3_X2 U3071 ( .A1(n2748), .A2(n3118), .A3(n3126), .ZN(n2824) );
  XNOR2_X1 U3072 ( .A(n2355), .B(n2356), .ZN(n2363) );
  OR2_X1 U3073 ( .A1(n2363), .A2(U3149), .ZN(n4070) );
  NAND2_X1 U3074 ( .A1(n3305), .A2(n4070), .ZN(n2376) );
  INV_X1 U3075 ( .A(n2357), .ZN(n2358) );
  NAND2_X1 U3076 ( .A1(n2358), .A2(IR_REG_31__SCAN_IN), .ZN(n2359) );
  NAND2_X1 U3077 ( .A1(n2360), .A2(n2361), .ZN(n2743) );
  INV_X1 U3078 ( .A(n2743), .ZN(n4715) );
  NAND2_X1 U3079 ( .A1(n2361), .A2(IR_REG_31__SCAN_IN), .ZN(n2362) );
  NAND2_X1 U3080 ( .A1(n3075), .A2(n2363), .ZN(n2365) );
  AND2_X1 U3081 ( .A1(n2365), .A2(n2024), .ZN(n2374) );
  NAND2_X1 U3082 ( .A1(n2376), .A2(n2374), .ZN(n3152) );
  XNOR2_X1 U3083 ( .A(n2366), .B(IR_REG_27__SCAN_IN), .ZN(n4065) );
  NAND2_X1 U3084 ( .A1(n2055), .A2(IR_REG_31__SCAN_IN), .ZN(n2371) );
  MUX2_X1 U3085 ( .A(n2371), .B(IR_REG_31__SCAN_IN), .S(n2372), .Z(n2373) );
  NAND2_X1 U3086 ( .A1(n2373), .A2(n2434), .ZN(n3179) );
  NAND2_X1 U3087 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3779) );
  INV_X1 U3088 ( .A(n2374), .ZN(n2375) );
  NAND2_X1 U3089 ( .A1(n4765), .A2(ADDR_REG_19__SCAN_IN), .ZN(n2377) );
  OAI211_X1 U3090 ( .C1(n4775), .C2(n4063), .A(n3779), .B(n2377), .ZN(n2378)
         );
  AOI21_X1 U3091 ( .B1(n2379), .B2(n4770), .A(n2378), .ZN(n2431) );
  INV_X1 U3092 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4732) );
  NAND2_X1 U3093 ( .A1(n4728), .A2(REG2_REG_1__SCAN_IN), .ZN(n3188) );
  INV_X1 U3094 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3326) );
  AND2_X1 U3095 ( .A1(n4729), .A2(REG2_REG_0__SCAN_IN), .ZN(n2381) );
  NAND2_X1 U3096 ( .A1(n3188), .A2(n3187), .ZN(n2385) );
  OAI21_X1 U3097 ( .B1(n2384), .B2(n2383), .A(n2382), .ZN(n3186) );
  NAND2_X1 U3098 ( .A1(n2385), .A2(n3186), .ZN(n3191) );
  NAND2_X1 U3099 ( .A1(n2384), .A2(REG2_REG_2__SCAN_IN), .ZN(n2386) );
  NAND2_X1 U3100 ( .A1(n3139), .A2(REG2_REG_3__SCAN_IN), .ZN(n2389) );
  NAND2_X1 U3101 ( .A1(n2387), .A2(n4726), .ZN(n2388) );
  NAND2_X1 U3102 ( .A1(n2390), .A2(n4725), .ZN(n2391) );
  INV_X1 U3103 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2392) );
  MUX2_X1 U3104 ( .A(n2392), .B(REG2_REG_5__SCAN_IN), .S(n3163), .Z(n3160) );
  NAND2_X1 U3105 ( .A1(n4724), .A2(REG2_REG_5__SCAN_IN), .ZN(n2393) );
  XNOR2_X1 U3106 ( .A(n2394), .B(n3170), .ZN(n3167) );
  NAND2_X1 U3107 ( .A1(n3167), .A2(REG2_REG_6__SCAN_IN), .ZN(n2396) );
  NAND2_X1 U3108 ( .A1(n2394), .A2(n4723), .ZN(n2395) );
  NAND2_X1 U3109 ( .A1(n2396), .A2(n2395), .ZN(n3210) );
  INV_X1 U3110 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2397) );
  MUX2_X1 U3111 ( .A(REG2_REG_7__SCAN_IN), .B(n2397), .S(n4722), .Z(n3209) );
  NAND2_X1 U3112 ( .A1(n3210), .A2(n3209), .ZN(n3208) );
  NAND2_X1 U3113 ( .A1(n4722), .A2(REG2_REG_7__SCAN_IN), .ZN(n2398) );
  INV_X1 U3114 ( .A(n4721), .ZN(n3274) );
  NAND2_X1 U3115 ( .A1(n3271), .A2(REG2_REG_8__SCAN_IN), .ZN(n2401) );
  NAND2_X1 U3116 ( .A1(n2399), .A2(n4721), .ZN(n2400) );
  NAND2_X1 U3117 ( .A1(n2401), .A2(n2400), .ZN(n3482) );
  INV_X1 U3118 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2402) );
  XNOR2_X1 U3119 ( .A(n4720), .B(n2402), .ZN(n3483) );
  NAND2_X1 U3120 ( .A1(n3482), .A2(n3483), .ZN(n2404) );
  NAND2_X1 U3121 ( .A1(n4720), .A2(REG2_REG_9__SCAN_IN), .ZN(n2403) );
  NAND2_X1 U3122 ( .A1(n2405), .A2(n4719), .ZN(n2406) );
  INV_X1 U3123 ( .A(REG2_REG_11__SCAN_IN), .ZN(n2407) );
  MUX2_X1 U3124 ( .A(n2407), .B(REG2_REG_11__SCAN_IN), .S(n2542), .Z(n4098) );
  NAND2_X1 U3125 ( .A1(n4099), .A2(n4098), .ZN(n4097) );
  NAND2_X1 U3126 ( .A1(n2291), .A2(REG2_REG_11__SCAN_IN), .ZN(n2408) );
  NAND2_X1 U3127 ( .A1(n2409), .A2(n4718), .ZN(n2410) );
  INV_X1 U3128 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3654) );
  NOR2_X1 U3129 ( .A1(n3662), .A2(n3654), .ZN(n2411) );
  NAND2_X1 U3130 ( .A1(n3662), .A2(n3654), .ZN(n2412) );
  NAND2_X1 U3131 ( .A1(REG2_REG_15__SCAN_IN), .A2(n2575), .ZN(n2415) );
  OAI21_X1 U3132 ( .B1(REG2_REG_15__SCAN_IN), .B2(n2575), .A(n2415), .ZN(n4741) );
  XNOR2_X1 U3133 ( .A(n2417), .B(n2585), .ZN(n4753) );
  INV_X1 U3134 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4752) );
  NAND2_X1 U3135 ( .A1(n2417), .A2(n4810), .ZN(n2418) );
  XNOR2_X1 U3136 ( .A(n2419), .B(REG2_REG_17__SCAN_IN), .ZN(n4107) );
  NAND2_X1 U3137 ( .A1(n2419), .A2(n2420), .ZN(n2421) );
  INV_X1 U3138 ( .A(REG2_REG_18__SCAN_IN), .ZN(n2422) );
  AOI22_X1 U3139 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4808), .B1(n2608), .B2(
        n2422), .ZN(n4763) );
  INV_X1 U3140 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2424) );
  MUX2_X1 U3141 ( .A(n2424), .B(REG2_REG_19__SCAN_IN), .S(n4063), .Z(n2425) );
  INV_X1 U3142 ( .A(n2425), .ZN(n2426) );
  NAND2_X1 U3143 ( .A1(n4713), .A2(n4065), .ZN(n2428) );
  NAND2_X1 U3144 ( .A1(n2429), .A2(n4096), .ZN(n2430) );
  NAND2_X1 U3145 ( .A1(n2431), .A2(n2430), .ZN(U3259) );
  INV_X1 U3146 ( .A(n2440), .ZN(n2438) );
  NAND2_X1 U3147 ( .A1(n2434), .A2(IR_REG_31__SCAN_IN), .ZN(n2435) );
  NAND2_X1 U31480 ( .A1(n2479), .A2(REG1_REG_0__SCAN_IN), .ZN(n2444) );
  NAND2_X1 U31490 ( .A1(n2461), .A2(REG0_REG_0__SCAN_IN), .ZN(n2443) );
  NAND2_X1 U3150 ( .A1(n2468), .A2(REG3_REG_0__SCAN_IN), .ZN(n2442) );
  NAND2_X1 U3151 ( .A1(n2469), .A2(REG2_REG_0__SCAN_IN), .ZN(n2441) );
  NAND2_X1 U3152 ( .A1(n2468), .A2(REG3_REG_1__SCAN_IN), .ZN(n2452) );
  INV_X1 U3153 ( .A(n4728), .ZN(n2447) );
  NAND2_X1 U3154 ( .A1(n2468), .A2(REG3_REG_2__SCAN_IN), .ZN(n2456) );
  NAND2_X1 U3155 ( .A1(n2469), .A2(REG2_REG_2__SCAN_IN), .ZN(n2455) );
  NAND2_X1 U3156 ( .A1(n2479), .A2(REG1_REG_2__SCAN_IN), .ZN(n2454) );
  NAND2_X1 U3157 ( .A1(n2461), .A2(REG0_REG_2__SCAN_IN), .ZN(n2453) );
  NAND4_X1 U3158 ( .A1(n2456), .A2(n2455), .A3(n2454), .A4(n2453), .ZN(n2840)
         );
  INV_X2 U3159 ( .A(n3291), .ZN(n3316) );
  NAND2_X1 U3160 ( .A1(n2840), .A2(n3316), .ZN(n3916) );
  NAND2_X1 U3161 ( .A1(n2459), .A2(n2832), .ZN(n3286) );
  MUX2_X1 U3162 ( .A(n4726), .B(DATAI_3_), .S(n2017), .Z(n3361) );
  INV_X1 U3163 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2460) );
  NAND2_X1 U3164 ( .A1(n2014), .A2(n2460), .ZN(n2465) );
  NAND2_X1 U3165 ( .A1(n2479), .A2(REG1_REG_3__SCAN_IN), .ZN(n2464) );
  NAND2_X1 U3166 ( .A1(n2469), .A2(REG2_REG_3__SCAN_IN), .ZN(n2463) );
  NAND2_X1 U3167 ( .A1(n3323), .A2(n3316), .ZN(n3337) );
  OAI21_X1 U3168 ( .B1(n3361), .B2(n3344), .A(n3337), .ZN(n2466) );
  INV_X1 U3169 ( .A(n2466), .ZN(n2474) );
  NAND2_X1 U3170 ( .A1(n2479), .A2(REG1_REG_4__SCAN_IN), .ZN(n2473) );
  INV_X1 U3171 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2467) );
  XNOR2_X1 U3172 ( .A(n2467), .B(REG3_REG_3__SCAN_IN), .ZN(n3436) );
  NAND2_X1 U3173 ( .A1(n2468), .A2(n3436), .ZN(n2472) );
  NAND2_X1 U3174 ( .A1(n2469), .A2(REG2_REG_4__SCAN_IN), .ZN(n2470) );
  NAND4_X1 U3175 ( .A1(n2473), .A2(n2472), .A3(n2471), .A4(n2470), .ZN(n2861)
         );
  MUX2_X1 U3176 ( .A(n4725), .B(DATAI_4_), .S(n3694), .Z(n2475) );
  NAND2_X1 U3177 ( .A1(n2861), .A2(n3336), .ZN(n3921) );
  NAND2_X1 U3178 ( .A1(n3390), .A2(n2475), .ZN(n3919) );
  NAND2_X1 U3179 ( .A1(n3921), .A2(n3919), .ZN(n3341) );
  NAND3_X1 U3180 ( .A1(n3288), .A2(n2474), .A3(n3341), .ZN(n2478) );
  AND2_X1 U3181 ( .A1(n3344), .A2(n3361), .ZN(n2476) );
  AOI22_X1 U3182 ( .A1(n3341), .A2(n2476), .B1(n2475), .B2(n2861), .ZN(n2477)
         );
  NAND2_X1 U3183 ( .A1(n2478), .A2(n2477), .ZN(n3374) );
  NAND2_X1 U3184 ( .A1(n3695), .A2(REG1_REG_5__SCAN_IN), .ZN(n2487) );
  INV_X1 U3185 ( .A(n2480), .ZN(n2482) );
  INV_X1 U3186 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2481) );
  NAND2_X1 U3187 ( .A1(n2482), .A2(n2481), .ZN(n2483) );
  AND2_X1 U3188 ( .A1(n2492), .A2(n2483), .ZN(n3382) );
  NAND2_X1 U3189 ( .A1(n2014), .A2(n3382), .ZN(n2486) );
  NAND2_X1 U3190 ( .A1(n2461), .A2(REG0_REG_5__SCAN_IN), .ZN(n2485) );
  INV_X2 U3191 ( .A(n2607), .ZN(n3696) );
  NAND2_X1 U3192 ( .A1(n3696), .A2(REG2_REG_5__SCAN_IN), .ZN(n2484) );
  NAND4_X1 U3193 ( .A1(n2487), .A2(n2486), .A3(n2485), .A4(n2484), .ZN(n4076)
         );
  INV_X1 U3194 ( .A(n2016), .ZN(n3402) );
  MUX2_X1 U3195 ( .A(n4724), .B(DATAI_5_), .S(n2017), .Z(n3464) );
  NAND2_X1 U3196 ( .A1(n3402), .A2(n2070), .ZN(n2488) );
  NAND2_X1 U3197 ( .A1(n2016), .A2(n3464), .ZN(n2489) );
  NAND2_X1 U3198 ( .A1(n3695), .A2(REG1_REG_6__SCAN_IN), .ZN(n2497) );
  INV_X1 U3199 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2491) );
  NAND2_X1 U3200 ( .A1(n2492), .A2(n2491), .ZN(n2493) );
  AND2_X1 U3201 ( .A1(n2499), .A2(n2493), .ZN(n3412) );
  NAND2_X1 U3202 ( .A1(n2014), .A2(n3412), .ZN(n2496) );
  NAND2_X1 U3203 ( .A1(n2461), .A2(REG0_REG_6__SCAN_IN), .ZN(n2495) );
  NAND2_X1 U3204 ( .A1(n3696), .A2(REG2_REG_6__SCAN_IN), .ZN(n2494) );
  NAND4_X1 U3205 ( .A1(n2497), .A2(n2496), .A3(n2495), .A4(n2494), .ZN(n3447)
         );
  MUX2_X1 U3206 ( .A(n4723), .B(DATAI_6_), .S(n3694), .Z(n3411) );
  NAND2_X1 U3207 ( .A1(n3695), .A2(REG1_REG_7__SCAN_IN), .ZN(n2504) );
  INV_X1 U3208 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2498) );
  NAND2_X1 U3209 ( .A1(n2499), .A2(n2498), .ZN(n2500) );
  AND2_X1 U32100 ( .A1(n2516), .A2(n2500), .ZN(n3458) );
  NAND2_X1 U32110 ( .A1(n2014), .A2(n3458), .ZN(n2503) );
  NAND2_X1 U32120 ( .A1(n2461), .A2(REG0_REG_7__SCAN_IN), .ZN(n2502) );
  NAND2_X1 U32130 ( .A1(n3696), .A2(REG2_REG_7__SCAN_IN), .ZN(n2501) );
  MUX2_X1 U32140 ( .A(n4722), .B(DATAI_7_), .S(n3694), .Z(n3456) );
  NAND2_X1 U32150 ( .A1(n3510), .A2(n3456), .ZN(n2705) );
  NAND2_X1 U32160 ( .A1(n4075), .A2(n2769), .ZN(n3927) );
  NAND2_X1 U32170 ( .A1(n3695), .A2(REG1_REG_8__SCAN_IN), .ZN(n2508) );
  XNOR2_X1 U32180 ( .A(n2516), .B(REG3_REG_8__SCAN_IN), .ZN(n3514) );
  NAND2_X1 U32190 ( .A1(n2014), .A2(n3514), .ZN(n2507) );
  NAND2_X1 U32200 ( .A1(n2461), .A2(REG0_REG_8__SCAN_IN), .ZN(n2506) );
  NAND2_X1 U32210 ( .A1(n3696), .A2(REG2_REG_8__SCAN_IN), .ZN(n2505) );
  MUX2_X1 U32220 ( .A(n4721), .B(DATAI_8_), .S(n3694), .Z(n3516) );
  INV_X1 U32230 ( .A(n3516), .ZN(n2707) );
  NAND2_X1 U32240 ( .A1(n3541), .A2(n2707), .ZN(n2509) );
  NAND2_X1 U32250 ( .A1(n3466), .A2(n3418), .ZN(n3451) );
  INV_X1 U32260 ( .A(n2509), .ZN(n2510) );
  NAND2_X1 U32270 ( .A1(n4075), .A2(n3456), .ZN(n3504) );
  OAI22_X1 U32280 ( .A1(n2510), .A2(n3504), .B1(n3541), .B2(n2707), .ZN(n2511)
         );
  NAND2_X1 U32290 ( .A1(n3695), .A2(REG1_REG_9__SCAN_IN), .ZN(n2521) );
  INV_X1 U32300 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2515) );
  INV_X1 U32310 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2514) );
  OAI21_X1 U32320 ( .B1(n2516), .B2(n2515), .A(n2514), .ZN(n2517) );
  AND2_X1 U32330 ( .A1(n2526), .A2(n2517), .ZN(n3553) );
  NAND2_X1 U32340 ( .A1(n2014), .A2(n3553), .ZN(n2520) );
  NAND2_X1 U32350 ( .A1(n2461), .A2(REG0_REG_9__SCAN_IN), .ZN(n2519) );
  NAND2_X1 U32360 ( .A1(n3696), .A2(REG2_REG_9__SCAN_IN), .ZN(n2518) );
  NAND4_X1 U32370 ( .A1(n2521), .A2(n2520), .A3(n2519), .A4(n2518), .ZN(n3525)
         );
  MUX2_X1 U32380 ( .A(n4720), .B(DATAI_9_), .S(n3694), .Z(n3606) );
  NAND2_X1 U32390 ( .A1(n3525), .A2(n3606), .ZN(n2522) );
  NAND2_X1 U32400 ( .A1(n3538), .A2(n2522), .ZN(n2524) );
  NAND2_X1 U32410 ( .A1(n3672), .A2(n3543), .ZN(n2523) );
  NAND2_X1 U32420 ( .A1(n2524), .A2(n2523), .ZN(n3522) );
  NAND2_X1 U32430 ( .A1(n3695), .A2(REG1_REG_10__SCAN_IN), .ZN(n2531) );
  INV_X1 U32440 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4498) );
  NAND2_X1 U32450 ( .A1(n2526), .A2(n4498), .ZN(n2527) );
  AND2_X1 U32460 ( .A1(n2534), .A2(n2527), .ZN(n3679) );
  NAND2_X1 U32470 ( .A1(n2014), .A2(n3679), .ZN(n2530) );
  NAND2_X1 U32480 ( .A1(n2461), .A2(REG0_REG_10__SCAN_IN), .ZN(n2529) );
  NAND2_X1 U32490 ( .A1(n3696), .A2(REG2_REG_10__SCAN_IN), .ZN(n2528) );
  NAND4_X1 U32500 ( .A1(n2531), .A2(n2530), .A3(n2529), .A4(n2528), .ZN(n4485)
         );
  MUX2_X1 U32510 ( .A(n4719), .B(DATAI_10_), .S(n3694), .Z(n3668) );
  NOR2_X1 U32520 ( .A1(n4485), .A2(n3668), .ZN(n2532) );
  NAND2_X1 U32530 ( .A1(n4485), .A2(n3668), .ZN(n2533) );
  NAND2_X1 U32540 ( .A1(n3695), .A2(REG1_REG_11__SCAN_IN), .ZN(n2540) );
  NAND2_X1 U32550 ( .A1(n2534), .A2(n4521), .ZN(n2535) );
  AND2_X1 U32560 ( .A1(n2546), .A2(n2535), .ZN(n3624) );
  NAND2_X1 U32570 ( .A1(n2014), .A2(n3624), .ZN(n2539) );
  NAND2_X1 U32580 ( .A1(n2461), .A2(REG0_REG_11__SCAN_IN), .ZN(n2538) );
  NAND2_X1 U32590 ( .A1(n3696), .A2(REG2_REG_11__SCAN_IN), .ZN(n2537) );
  NAND4_X1 U32600 ( .A1(n2540), .A2(n2539), .A3(n2538), .A4(n2537), .ZN(n4473)
         );
  INV_X1 U32610 ( .A(DATAI_11_), .ZN(n2541) );
  MUX2_X1 U32620 ( .A(n2542), .B(n2541), .S(n3694), .Z(n3621) );
  NAND2_X1 U32630 ( .A1(n3799), .A2(n3566), .ZN(n3583) );
  NAND2_X1 U32640 ( .A1(n4473), .A2(n3621), .ZN(n3585) );
  NAND2_X1 U32650 ( .A1(n3799), .A2(n3621), .ZN(n2543) );
  NAND2_X1 U32660 ( .A1(n3695), .A2(REG1_REG_12__SCAN_IN), .ZN(n2551) );
  INV_X1 U32670 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2545) );
  NAND2_X1 U32680 ( .A1(n2546), .A2(n2545), .ZN(n2547) );
  AND2_X1 U32690 ( .A1(n2556), .A2(n2547), .ZN(n3803) );
  NAND2_X1 U32700 ( .A1(n2014), .A2(n3803), .ZN(n2550) );
  NAND2_X1 U32710 ( .A1(n2536), .A2(REG0_REG_12__SCAN_IN), .ZN(n2549) );
  NAND2_X1 U32720 ( .A1(n3696), .A2(REG2_REG_12__SCAN_IN), .ZN(n2548) );
  NAND4_X1 U32730 ( .A1(n2551), .A2(n2550), .A3(n2549), .A4(n2548), .ZN(n4073)
         );
  MUX2_X1 U32740 ( .A(DATAI_12_), .B(n4718), .S(n2018), .Z(n3590) );
  NAND2_X1 U32750 ( .A1(n4073), .A2(n3590), .ZN(n2552) );
  NAND2_X1 U32760 ( .A1(n3587), .A2(n2552), .ZN(n2554) );
  INV_X1 U32770 ( .A(n4073), .ZN(n3853) );
  INV_X1 U32780 ( .A(n3590), .ZN(n4478) );
  NAND2_X1 U32790 ( .A1(n3853), .A2(n4478), .ZN(n2553) );
  NAND2_X1 U32800 ( .A1(n2554), .A2(n2553), .ZN(n3636) );
  NAND2_X1 U32810 ( .A1(n3695), .A2(REG1_REG_13__SCAN_IN), .ZN(n2561) );
  NAND2_X1 U32820 ( .A1(n2556), .A2(n2555), .ZN(n2557) );
  AND2_X1 U32830 ( .A1(n2569), .A2(n2557), .ZN(n3858) );
  NAND2_X1 U32840 ( .A1(n2014), .A2(n3858), .ZN(n2560) );
  NAND2_X1 U32850 ( .A1(n2461), .A2(REG0_REG_13__SCAN_IN), .ZN(n2559) );
  NAND2_X1 U32860 ( .A1(n3696), .A2(REG2_REG_13__SCAN_IN), .ZN(n2558) );
  MUX2_X1 U32870 ( .A(n3659), .B(DATAI_13_), .S(n3694), .Z(n3627) );
  NOR2_X1 U32880 ( .A1(n4474), .A2(n3627), .ZN(n2562) );
  NAND2_X1 U32890 ( .A1(n3695), .A2(REG1_REG_14__SCAN_IN), .ZN(n2566) );
  XNOR2_X1 U32900 ( .A(n2569), .B(REG3_REG_14__SCAN_IN), .ZN(n3759) );
  NAND2_X1 U32910 ( .A1(n2014), .A2(n3759), .ZN(n2565) );
  NAND2_X1 U32920 ( .A1(n2536), .A2(REG0_REG_14__SCAN_IN), .ZN(n2564) );
  NAND2_X1 U32930 ( .A1(n2469), .A2(REG2_REG_14__SCAN_IN), .ZN(n2563) );
  NAND4_X1 U32940 ( .A1(n2566), .A2(n2565), .A3(n2564), .A4(n2563), .ZN(n4450)
         );
  MUX2_X1 U32950 ( .A(n4813), .B(DATAI_14_), .S(n3694), .Z(n4459) );
  NAND2_X1 U32960 ( .A1(n3854), .A2(n4459), .ZN(n3950) );
  NAND2_X1 U32970 ( .A1(n4450), .A2(n3756), .ZN(n3932) );
  NAND2_X1 U32980 ( .A1(n3950), .A2(n3932), .ZN(n3645) );
  NAND2_X1 U32990 ( .A1(n3695), .A2(REG1_REG_15__SCAN_IN), .ZN(n2574) );
  INV_X1 U33000 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2568) );
  INV_X1 U33010 ( .A(REG3_REG_15__SCAN_IN), .ZN(n4547) );
  OAI21_X1 U33020 ( .B1(n2569), .B2(n2568), .A(n4547), .ZN(n2570) );
  AND2_X1 U33030 ( .A1(n2579), .A2(n2570), .ZN(n3903) );
  NAND2_X1 U33040 ( .A1(n2014), .A2(n3903), .ZN(n2573) );
  NAND2_X1 U33050 ( .A1(n2536), .A2(REG0_REG_15__SCAN_IN), .ZN(n2572) );
  NAND2_X1 U33060 ( .A1(n2469), .A2(REG2_REG_15__SCAN_IN), .ZN(n2571) );
  MUX2_X1 U33070 ( .A(n2575), .B(DATAI_15_), .S(n3694), .Z(n4449) );
  NAND2_X1 U33080 ( .A1(n4440), .A2(n4449), .ZN(n2576) );
  NAND2_X1 U33090 ( .A1(n3684), .A2(n2576), .ZN(n2578) );
  INV_X1 U33100 ( .A(n4449), .ZN(n3899) );
  NAND2_X1 U33110 ( .A1(n4463), .A2(n3899), .ZN(n2577) );
  NAND2_X1 U33120 ( .A1(n2579), .A2(n4610), .ZN(n2580) );
  AND2_X1 U33130 ( .A1(n2610), .A2(n2580), .ZN(n4353) );
  NAND2_X1 U33140 ( .A1(n4353), .A2(n2014), .ZN(n2584) );
  NAND2_X1 U33150 ( .A1(n2536), .A2(REG0_REG_16__SCAN_IN), .ZN(n2583) );
  NAND2_X1 U33160 ( .A1(n3695), .A2(REG1_REG_16__SCAN_IN), .ZN(n2582) );
  NAND2_X1 U33170 ( .A1(n2469), .A2(REG2_REG_16__SCAN_IN), .ZN(n2581) );
  MUX2_X1 U33180 ( .A(n2585), .B(DATAI_16_), .S(n2024), .Z(n4352) );
  NAND2_X1 U33190 ( .A1(n4452), .A2(n4352), .ZN(n4033) );
  INV_X1 U33200 ( .A(n4352), .ZN(n4443) );
  NAND2_X1 U33210 ( .A1(n4432), .A2(n4443), .ZN(n3952) );
  NAND2_X1 U33220 ( .A1(n2596), .A2(n3844), .ZN(n2587) );
  AND2_X1 U33230 ( .A1(n2630), .A2(n2587), .ZN(n4274) );
  NAND2_X1 U33240 ( .A1(n4274), .A2(n2014), .ZN(n2593) );
  INV_X1 U33250 ( .A(REG1_REG_20__SCAN_IN), .ZN(n2590) );
  NAND2_X1 U33260 ( .A1(n2536), .A2(REG0_REG_20__SCAN_IN), .ZN(n2589) );
  NAND2_X1 U33270 ( .A1(n2469), .A2(REG2_REG_20__SCAN_IN), .ZN(n2588) );
  OAI211_X1 U33280 ( .C1(n2701), .C2(n2590), .A(n2589), .B(n2588), .ZN(n2591)
         );
  INV_X1 U33290 ( .A(n2591), .ZN(n2592) );
  OR2_X1 U33300 ( .A1(n4405), .A2(n4415), .ZN(n4005) );
  INV_X1 U33310 ( .A(n4005), .ZN(n2620) );
  INV_X1 U33320 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2594) );
  NAND2_X1 U33330 ( .A1(n2604), .A2(n2594), .ZN(n2595) );
  NAND2_X1 U33340 ( .A1(n2596), .A2(n2595), .ZN(n3778) );
  OR2_X1 U33350 ( .A1(n3778), .A2(n2777), .ZN(n2601) );
  NAND2_X1 U33360 ( .A1(n2461), .A2(REG0_REG_19__SCAN_IN), .ZN(n2598) );
  NAND2_X1 U33370 ( .A1(n2469), .A2(REG2_REG_19__SCAN_IN), .ZN(n2597) );
  OAI211_X1 U33380 ( .C1(n2701), .C2(n2335), .A(n2598), .B(n2597), .ZN(n2599)
         );
  INV_X1 U33390 ( .A(n2599), .ZN(n2600) );
  MUX2_X1 U33400 ( .A(n4717), .B(DATAI_19_), .S(n3694), .Z(n4291) );
  OR2_X1 U33410 ( .A1(n4416), .A2(n4291), .ZN(n4264) );
  INV_X1 U33420 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2602) );
  NAND2_X1 U33430 ( .A1(n2612), .A2(n2602), .ZN(n2603) );
  NAND2_X1 U33440 ( .A1(n2604), .A2(n2603), .ZN(n4316) );
  OR2_X1 U33450 ( .A1(n4316), .A2(n2777), .ZN(n2606) );
  AOI22_X1 U33460 ( .A1(n3695), .A2(REG1_REG_18__SCAN_IN), .B1(n2536), .B2(
        REG0_REG_18__SCAN_IN), .ZN(n2605) );
  OAI211_X1 U33470 ( .C1(n2607), .C2(n2422), .A(n2606), .B(n2605), .ZN(n4292)
         );
  INV_X1 U33480 ( .A(n4292), .ZN(n4434) );
  MUX2_X1 U33490 ( .A(n2608), .B(DATAI_18_), .S(n3694), .Z(n4308) );
  NAND2_X1 U33500 ( .A1(n4434), .A2(n4315), .ZN(n4262) );
  AND2_X1 U33510 ( .A1(n4264), .A2(n4262), .ZN(n2621) );
  INV_X1 U33520 ( .A(n2621), .ZN(n2615) );
  NAND2_X1 U3353 ( .A1(n2610), .A2(n2609), .ZN(n2611) );
  NAND2_X1 U33540 ( .A1(n2612), .A2(n2611), .ZN(n4333) );
  AOI22_X1 U3355 ( .A1(n3695), .A2(REG1_REG_17__SCAN_IN), .B1(n2536), .B2(
        REG0_REG_17__SCAN_IN), .ZN(n2614) );
  NAND2_X1 U3356 ( .A1(n2469), .A2(REG2_REG_17__SCAN_IN), .ZN(n2613) );
  MUX2_X1 U3357 ( .A(n4109), .B(DATAI_17_), .S(n3694), .Z(n4431) );
  NAND2_X1 U3358 ( .A1(n4441), .A2(n4431), .ZN(n4259) );
  OR2_X1 U3359 ( .A1(n2615), .A2(n4259), .ZN(n2618) );
  NAND2_X1 U3360 ( .A1(n4434), .A2(n4308), .ZN(n4286) );
  NAND2_X1 U3361 ( .A1(n4292), .A2(n4315), .ZN(n4287) );
  NAND2_X1 U3362 ( .A1(n4286), .A2(n4287), .ZN(n4261) );
  NAND2_X1 U3363 ( .A1(n4416), .A2(n4291), .ZN(n4263) );
  NAND2_X1 U3364 ( .A1(n4405), .A2(n4415), .ZN(n4004) );
  OAI211_X1 U3365 ( .C1(n2615), .C2(n4261), .A(n4263), .B(n4004), .ZN(n2616)
         );
  INV_X1 U3366 ( .A(n2616), .ZN(n2617) );
  AND2_X1 U3367 ( .A1(n2618), .A2(n2617), .ZN(n2619) );
  INV_X1 U3368 ( .A(n2625), .ZN(n2624) );
  OR2_X1 U3369 ( .A1(n4441), .A2(n4431), .ZN(n4258) );
  AND2_X1 U3370 ( .A1(n4258), .A2(n2621), .ZN(n2622) );
  AND2_X1 U3371 ( .A1(n2622), .A2(n4005), .ZN(n2623) );
  NOR2_X1 U3372 ( .A1(n2624), .A2(n2623), .ZN(n2627) );
  NAND2_X1 U3373 ( .A1(n4432), .A2(n4352), .ZN(n4257) );
  AND2_X1 U3374 ( .A1(n4257), .A2(n2625), .ZN(n2626) );
  OR2_X1 U3375 ( .A1(n2627), .A2(n2626), .ZN(n4240) );
  INV_X1 U3376 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2629) );
  NAND2_X1 U3377 ( .A1(n2630), .A2(n2629), .ZN(n2631) );
  NAND2_X1 U3378 ( .A1(n2641), .A2(n2631), .ZN(n4248) );
  INV_X1 U3379 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4411) );
  NAND2_X1 U3380 ( .A1(n2536), .A2(REG0_REG_21__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U3381 ( .A1(n2469), .A2(REG2_REG_21__SCAN_IN), .ZN(n2632) );
  OAI211_X1 U3382 ( .C1(n2701), .C2(n4411), .A(n2633), .B(n2632), .ZN(n2634)
         );
  INV_X1 U3383 ( .A(n2634), .ZN(n2635) );
  NAND2_X1 U3384 ( .A1(n4414), .A2(n4404), .ZN(n2637) );
  AND2_X1 U3385 ( .A1(n4240), .A2(n2637), .ZN(n2638) );
  INV_X1 U3386 ( .A(n4404), .ZN(n4245) );
  NAND2_X1 U3387 ( .A1(n3866), .A2(n4245), .ZN(n2639) );
  NAND2_X1 U3388 ( .A1(n2640), .A2(n2639), .ZN(n4229) );
  INV_X1 U3389 ( .A(n4229), .ZN(n2648) );
  NAND2_X1 U3390 ( .A1(n2641), .A2(n4579), .ZN(n2642) );
  AND2_X1 U3391 ( .A1(n2655), .A2(n2642), .ZN(n4234) );
  NAND2_X1 U3392 ( .A1(n4234), .A2(n2014), .ZN(n2647) );
  INV_X1 U3393 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4402) );
  NAND2_X1 U3394 ( .A1(n2536), .A2(REG0_REG_22__SCAN_IN), .ZN(n2644) );
  NAND2_X1 U3395 ( .A1(n2469), .A2(REG2_REG_22__SCAN_IN), .ZN(n2643) );
  OAI211_X1 U3396 ( .C1(n2701), .C2(n4402), .A(n2644), .B(n2643), .ZN(n2645)
         );
  INV_X1 U3397 ( .A(n2645), .ZN(n2646) );
  INV_X1 U3398 ( .A(n4232), .ZN(n3867) );
  NAND2_X1 U3399 ( .A1(n4247), .A2(n3867), .ZN(n2730) );
  NAND2_X1 U3400 ( .A1(n4204), .A2(n2730), .ZN(n4222) );
  INV_X1 U3401 ( .A(n4222), .ZN(n4230) );
  NAND2_X1 U3402 ( .A1(n4247), .A2(n4232), .ZN(n4211) );
  XNOR2_X1 U3403 ( .A(n2655), .B(REG3_REG_23__SCAN_IN), .ZN(n4217) );
  NAND2_X1 U3404 ( .A1(n4217), .A2(n2014), .ZN(n2653) );
  INV_X1 U3405 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4397) );
  NAND2_X1 U3406 ( .A1(n2536), .A2(REG0_REG_23__SCAN_IN), .ZN(n2650) );
  NAND2_X1 U3407 ( .A1(n2469), .A2(REG2_REG_23__SCAN_IN), .ZN(n2649) );
  OAI211_X1 U3408 ( .C1(n2701), .C2(n4397), .A(n2650), .B(n2649), .ZN(n2651)
         );
  INV_X1 U3409 ( .A(n2651), .ZN(n2652) );
  AND2_X1 U3410 ( .A1(n2024), .A2(DATAI_23_), .ZN(n4207) );
  NAND2_X1 U3411 ( .A1(n4224), .A2(n4207), .ZN(n2654) );
  AND2_X1 U3412 ( .A1(n4211), .A2(n2654), .ZN(n4186) );
  INV_X1 U3413 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4535) );
  INV_X1 U3414 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3833) );
  OAI21_X1 U3415 ( .B1(n2655), .B2(n4535), .A(n3833), .ZN(n2657) );
  AND2_X1 U3416 ( .A1(REG3_REG_23__SCAN_IN), .A2(REG3_REG_24__SCAN_IN), .ZN(
        n2656) );
  NAND2_X1 U3417 ( .A1(n2657), .A2(n2666), .ZN(n3832) );
  INV_X1 U3418 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4565) );
  NAND2_X1 U3419 ( .A1(n2536), .A2(REG0_REG_24__SCAN_IN), .ZN(n2659) );
  NAND2_X1 U3420 ( .A1(n2469), .A2(REG2_REG_24__SCAN_IN), .ZN(n2658) );
  OAI211_X1 U3421 ( .C1(n2701), .C2(n4565), .A(n2659), .B(n2658), .ZN(n2660)
         );
  INV_X1 U3422 ( .A(n2660), .ZN(n2661) );
  NAND2_X1 U3423 ( .A1(n3694), .A2(DATAI_24_), .ZN(n4195) );
  INV_X1 U3424 ( .A(n4195), .ZN(n4386) );
  AND2_X1 U3425 ( .A1(n4378), .A2(n4386), .ZN(n2664) );
  INV_X1 U3426 ( .A(n2664), .ZN(n2663) );
  AND2_X1 U3427 ( .A1(n4186), .A2(n2663), .ZN(n2665) );
  OR2_X1 U3428 ( .A1(n4224), .A2(n4207), .ZN(n4187) );
  INV_X1 U3429 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3719) );
  NAND2_X1 U3430 ( .A1(n2666), .A2(n3719), .ZN(n2667) );
  NAND2_X1 U3431 ( .A1(n4175), .A2(n2014), .ZN(n2672) );
  INV_X1 U3432 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4384) );
  NAND2_X1 U3433 ( .A1(n2536), .A2(REG0_REG_25__SCAN_IN), .ZN(n2669) );
  NAND2_X1 U3434 ( .A1(n3696), .A2(REG2_REG_25__SCAN_IN), .ZN(n2668) );
  OAI211_X1 U3435 ( .C1(n2701), .C2(n4384), .A(n2669), .B(n2668), .ZN(n2670)
         );
  INV_X1 U3436 ( .A(n2670), .ZN(n2671) );
  INV_X1 U3437 ( .A(n4387), .ZN(n4196) );
  INV_X1 U3438 ( .A(n4377), .ZN(n4177) );
  INV_X1 U3439 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2673) );
  NAND2_X1 U3440 ( .A1(n2674), .A2(n2673), .ZN(n2675) );
  INV_X1 U3441 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4375) );
  NAND2_X1 U3442 ( .A1(n2536), .A2(REG0_REG_26__SCAN_IN), .ZN(n2677) );
  NAND2_X1 U3443 ( .A1(n3696), .A2(REG2_REG_26__SCAN_IN), .ZN(n2676) );
  OAI211_X1 U3444 ( .C1(n2701), .C2(n4375), .A(n2677), .B(n2676), .ZN(n2678)
         );
  INV_X1 U3445 ( .A(n2678), .ZN(n2679) );
  AND2_X1 U3446 ( .A1(n4137), .A2(n4154), .ZN(n2680) );
  INV_X1 U3447 ( .A(REG3_REG_27__SCAN_IN), .ZN(n2681) );
  NAND2_X1 U3448 ( .A1(n2682), .A2(n2681), .ZN(n2683) );
  NAND2_X1 U3449 ( .A1(n4136), .A2(n2014), .ZN(n2688) );
  INV_X1 U3450 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4369) );
  NAND2_X1 U3451 ( .A1(n3696), .A2(REG2_REG_27__SCAN_IN), .ZN(n2685) );
  NAND2_X1 U3452 ( .A1(n2536), .A2(REG0_REG_27__SCAN_IN), .ZN(n2684) );
  OAI211_X1 U3453 ( .C1(n2701), .C2(n4369), .A(n2685), .B(n2684), .ZN(n2686)
         );
  INV_X1 U3454 ( .A(n2686), .ZN(n2687) );
  AND2_X1 U3455 ( .A1(n3694), .A2(DATAI_27_), .ZN(n3968) );
  XNOR2_X1 U3456 ( .A(n4124), .B(n3968), .ZN(n4052) );
  XNOR2_X1 U3457 ( .A(n2775), .B(n2689), .ZN(n4135) );
  INV_X1 U34580 ( .A(n4714), .ZN(n2744) );
  XNOR2_X1 U34590 ( .A(n3313), .B(n2744), .ZN(n2693) );
  NAND2_X1 U3460 ( .A1(n2693), .A2(n4063), .ZN(n3561) );
  NAND2_X1 U3461 ( .A1(n2694), .A2(n4717), .ZN(n4786) );
  INV_X1 U3462 ( .A(n2697), .ZN(n2695) );
  NAND2_X1 U3463 ( .A1(n2695), .A2(REG3_REG_28__SCAN_IN), .ZN(n3738) );
  INV_X1 U3464 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2696) );
  NAND2_X1 U3465 ( .A1(n2697), .A2(n2696), .ZN(n2698) );
  INV_X1 U3466 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2789) );
  NAND2_X1 U34670 ( .A1(n2536), .A2(REG0_REG_28__SCAN_IN), .ZN(n2700) );
  NAND2_X1 U3468 ( .A1(n3696), .A2(REG2_REG_28__SCAN_IN), .ZN(n2699) );
  OAI211_X1 U34690 ( .C1(n2701), .C2(n2789), .A(n2700), .B(n2699), .ZN(n2702)
         );
  INV_X1 U3470 ( .A(n2702), .ZN(n2703) );
  INV_X1 U34710 ( .A(n4143), .ZN(n2746) );
  NAND2_X1 U3472 ( .A1(n3989), .A2(n3911), .ZN(n3234) );
  NAND2_X1 U34730 ( .A1(n3234), .A2(n3913), .ZN(n3294) );
  NAND2_X1 U3474 ( .A1(n3294), .A2(n3988), .ZN(n3293) );
  NAND2_X1 U34750 ( .A1(n3430), .A2(n3361), .ZN(n3918) );
  INV_X1 U3476 ( .A(n3361), .ZN(n3338) );
  NAND2_X1 U34770 ( .A1(n3344), .A2(n3338), .ZN(n3915) );
  NAND2_X1 U3478 ( .A1(n3355), .A2(n3990), .ZN(n3354) );
  NAND2_X1 U34790 ( .A1(n3354), .A2(n3918), .ZN(n3343) );
  NAND2_X1 U3480 ( .A1(n3402), .A2(n3464), .ZN(n3937) );
  NAND2_X1 U34810 ( .A1(n3447), .A2(n3418), .ZN(n3936) );
  NAND2_X1 U3482 ( .A1(n3466), .A2(n3411), .ZN(n3923) );
  INV_X1 U34830 ( .A(n3445), .ZN(n2706) );
  NAND2_X1 U3484 ( .A1(n2706), .A2(n2705), .ZN(n3503) );
  NAND2_X1 U34850 ( .A1(n3672), .A2(n3606), .ZN(n3532) );
  INV_X1 U3486 ( .A(n3532), .ZN(n3930) );
  NAND2_X1 U34870 ( .A1(n4074), .A2(n2707), .ZN(n3926) );
  AND2_X1 U3488 ( .A1(n3525), .A2(n3543), .ZN(n3938) );
  INV_X1 U34890 ( .A(n3938), .ZN(n3533) );
  AND2_X1 U3490 ( .A1(n3926), .A2(n3533), .ZN(n2708) );
  AND2_X1 U34910 ( .A1(n3927), .A2(n2710), .ZN(n2709) );
  NAND2_X1 U3492 ( .A1(n3503), .A2(n2709), .ZN(n2714) );
  INV_X1 U34930 ( .A(n2710), .ZN(n2712) );
  NAND2_X1 U3494 ( .A1(n3541), .A2(n3516), .ZN(n3928) );
  AND2_X1 U34950 ( .A1(n3928), .A2(n3532), .ZN(n2711) );
  NAND2_X1 U3496 ( .A1(n4485), .A2(n3572), .ZN(n3944) );
  INV_X1 U34970 ( .A(n4485), .ZN(n3620) );
  NAND2_X1 U3498 ( .A1(n3620), .A2(n3668), .ZN(n3943) );
  NAND2_X1 U34990 ( .A1(n4478), .A2(n4073), .ZN(n3628) );
  NAND2_X1 U3500 ( .A1(n4474), .A2(n3855), .ZN(n2715) );
  NAND2_X1 U35010 ( .A1(n3628), .A2(n2715), .ZN(n2717) );
  INV_X1 U3502 ( .A(n3585), .ZN(n2716) );
  NOR2_X1 U35030 ( .A1(n2717), .A2(n2716), .ZN(n3945) );
  INV_X1 U3504 ( .A(n2717), .ZN(n2720) );
  NAND2_X1 U35050 ( .A1(n3853), .A2(n3590), .ZN(n3630) );
  NAND2_X1 U35060 ( .A1(n3583), .A2(n3630), .ZN(n2719) );
  NOR2_X1 U35070 ( .A1(n4474), .A2(n3855), .ZN(n2718) );
  AOI21_X1 U35080 ( .B1(n2720), .B2(n2719), .A(n2718), .ZN(n3948) );
  NAND2_X1 U35090 ( .A1(n2721), .A2(n3948), .ZN(n3643) );
  INV_X1 U35100 ( .A(n3645), .ZN(n3993) );
  NAND2_X1 U35110 ( .A1(n4463), .A2(n4449), .ZN(n3949) );
  NAND2_X1 U35120 ( .A1(n4440), .A2(n3899), .ZN(n3933) );
  NAND2_X1 U35130 ( .A1(n3949), .A2(n3933), .ZN(n4006) );
  NAND2_X1 U35140 ( .A1(n3681), .A2(n3933), .ZN(n4348) );
  NAND2_X1 U35150 ( .A1(n4348), .A2(n4357), .ZN(n4347) );
  NAND2_X1 U35160 ( .A1(n4416), .A2(n4301), .ZN(n2722) );
  AND2_X1 U35170 ( .A1(n2722), .A2(n4287), .ZN(n2724) );
  INV_X1 U35180 ( .A(n4431), .ZN(n4335) );
  NAND2_X1 U35190 ( .A1(n4441), .A2(n4335), .ZN(n4283) );
  NAND2_X1 U35200 ( .A1(n2724), .A2(n4283), .ZN(n3955) );
  NAND2_X1 U35210 ( .A1(n4405), .A2(n4277), .ZN(n2728) );
  INV_X1 U35220 ( .A(n2728), .ZN(n3956) );
  OR2_X1 U35230 ( .A1(n4441), .A2(n4335), .ZN(n4284) );
  NAND2_X1 U35240 ( .A1(n4286), .A2(n4284), .ZN(n2723) );
  NAND2_X1 U35250 ( .A1(n2724), .A2(n2723), .ZN(n2726) );
  OR2_X1 U35260 ( .A1(n4416), .A2(n4301), .ZN(n2725) );
  NAND2_X1 U35270 ( .A1(n2726), .A2(n2725), .ZN(n4269) );
  NOR2_X1 U35280 ( .A1(n4405), .A2(n4277), .ZN(n2727) );
  OR2_X1 U35290 ( .A1(n4269), .A2(n2727), .ZN(n2729) );
  NAND2_X1 U35300 ( .A1(n2729), .A2(n2728), .ZN(n4035) );
  NAND2_X1 U35310 ( .A1(n4224), .A2(n4216), .ZN(n4020) );
  AND2_X1 U35320 ( .A1(n4020), .A2(n2730), .ZN(n3961) );
  AND2_X1 U35330 ( .A1(n4414), .A2(n4245), .ZN(n4002) );
  NAND2_X1 U35340 ( .A1(n4204), .A2(n4002), .ZN(n2731) );
  NAND2_X1 U35350 ( .A1(n4238), .A2(n4036), .ZN(n2732) );
  NAND2_X1 U35360 ( .A1(n3866), .A2(n4404), .ZN(n4202) );
  NAND2_X1 U35370 ( .A1(n4204), .A2(n4202), .ZN(n3962) );
  NOR2_X1 U35380 ( .A1(n4224), .A2(n4216), .ZN(n4022) );
  AOI21_X1 U35390 ( .B1(n4036), .B2(n3962), .A(n4022), .ZN(n4039) );
  NOR2_X1 U35400 ( .A1(n4378), .A2(n4195), .ZN(n4040) );
  INV_X1 U35410 ( .A(n4154), .ZN(n4159) );
  NAND2_X1 U35420 ( .A1(n2734), .A2(n4148), .ZN(n4045) );
  NOR2_X1 U35430 ( .A1(n4168), .A2(n4045), .ZN(n2737) );
  INV_X1 U35440 ( .A(n4045), .ZN(n2735) );
  NAND2_X1 U35450 ( .A1(n4387), .A2(n4177), .ZN(n4019) );
  NAND2_X1 U35460 ( .A1(n4378), .A2(n4195), .ZN(n4167) );
  NAND2_X1 U35470 ( .A1(n4019), .A2(n4167), .ZN(n4149) );
  AND2_X1 U35480 ( .A1(n4137), .A2(n4159), .ZN(n4048) );
  AOI21_X1 U35490 ( .B1(n2735), .B2(n4149), .A(n4048), .ZN(n3967) );
  INV_X1 U35500 ( .A(n3967), .ZN(n2736) );
  NOR2_X1 U35510 ( .A1(n2737), .A2(n2736), .ZN(n2739) );
  OR2_X1 U35520 ( .A1(n2737), .A2(n2032), .ZN(n2738) );
  OAI21_X1 U35530 ( .B1(n4052), .B2(n2739), .A(n2738), .ZN(n2742) );
  OR2_X1 U35540 ( .A1(n2743), .A2(n2694), .ZN(n2741) );
  NAND2_X1 U35550 ( .A1(n4717), .A2(n4714), .ZN(n2740) );
  NAND2_X1 U35560 ( .A1(n2742), .A2(n4465), .ZN(n4146) );
  AND2_X2 U35570 ( .A1(n4713), .A2(n3075), .ZN(n4486) );
  NAND2_X1 U35580 ( .A1(n2744), .A2(n2743), .ZN(n3199) );
  INV_X1 U35590 ( .A(n3199), .ZN(n3073) );
  AND2_X2 U35600 ( .A1(n3073), .A2(n4716), .ZN(n4458) );
  AOI22_X1 U35610 ( .A1(n4137), .A2(n4486), .B1(n3968), .B2(n4458), .ZN(n2745)
         );
  OAI211_X1 U35620 ( .C1(n2746), .C2(n4462), .A(n4146), .B(n2745), .ZN(n2747)
         );
  AOI21_X1 U35630 ( .B1(n4135), .B2(n4482), .A(n2747), .ZN(n4370) );
  INV_X1 U35640 ( .A(REG0_REG_27__SCAN_IN), .ZN(n2767) );
  INV_X1 U35650 ( .A(B_REG_SCAN_IN), .ZN(n2749) );
  NOR2_X1 U35660 ( .A1(n3118), .A2(n2749), .ZN(n2750) );
  MUX2_X1 U35670 ( .A(n2750), .B(n2749), .S(n2748), .Z(n2751) );
  INV_X1 U35680 ( .A(D_REG_1__SCAN_IN), .ZN(n3132) );
  NAND2_X1 U35690 ( .A1(n3125), .A2(n3132), .ZN(n3306) );
  INV_X1 U35700 ( .A(n3118), .ZN(n2753) );
  NAND2_X1 U35710 ( .A1(n2753), .A2(n2752), .ZN(n3130) );
  NAND2_X1 U35720 ( .A1(n3306), .A2(n3130), .ZN(n2765) );
  NOR2_X1 U35730 ( .A1(n4644), .A2(n4715), .ZN(n3097) );
  NAND2_X1 U35740 ( .A1(n2694), .A2(n4063), .ZN(n3074) );
  NAND2_X1 U35750 ( .A1(n3074), .A2(n3075), .ZN(n3088) );
  INV_X1 U35760 ( .A(n3088), .ZN(n3304) );
  OR2_X1 U35770 ( .A1(n3097), .A2(n3304), .ZN(n2754) );
  NOR2_X1 U35780 ( .A1(n2754), .A2(n3305), .ZN(n2764) );
  NOR4_X1 U35790 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_18__SCAN_IN), .ZN(n2758) );
  NOR4_X1 U35800 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2757) );
  NOR4_X1 U35810 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_26__SCAN_IN), .ZN(n2756) );
  NOR4_X1 U3582 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2755) );
  NAND4_X1 U3583 ( .A1(n2758), .A2(n2757), .A3(n2756), .A4(n2755), .ZN(n2763)
         );
  NOR4_X1 U3584 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n4508) );
  NOR2_X1 U3585 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .ZN(n2761)
         );
  NOR4_X1 U3586 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2760) );
  NOR4_X1 U3587 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n2759) );
  NAND4_X1 U3588 ( .A1(n4508), .A2(n2761), .A3(n2760), .A4(n2759), .ZN(n2762)
         );
  OAI21_X1 U3589 ( .B1(n2763), .B2(n2762), .A(n3125), .ZN(n3071) );
  INV_X1 U3590 ( .A(D_REG_0__SCAN_IN), .ZN(n3129) );
  NOR2_X1 U3591 ( .A1(n2748), .A2(n3126), .ZN(n2766) );
  INV_X1 U3592 ( .A(n3072), .ZN(n3309) );
  MUX2_X1 U3593 ( .A(n4370), .B(n2767), .S(n4822), .Z(n2773) );
  NAND2_X1 U3594 ( .A1(n3239), .A2(n3316), .ZN(n3362) );
  NAND2_X1 U3595 ( .A1(n2768), .A2(n3338), .ZN(n3335) );
  NOR2_X1 U3596 ( .A1(n2771), .A2(n4140), .ZN(n2772) );
  OR2_X1 U3597 ( .A1(n2788), .A2(n2772), .ZN(n4372) );
  NAND2_X1 U3598 ( .A1(n4824), .A2(n4640), .ZN(n4706) );
  NAND2_X1 U3599 ( .A1(n2773), .A2(n2031), .ZN(U3513) );
  NOR2_X1 U3600 ( .A1(n4124), .A2(n3968), .ZN(n2774) );
  INV_X1 U3601 ( .A(n4124), .ZN(n4157) );
  AND2_X1 U3602 ( .A1(n3694), .A2(DATAI_28_), .ZN(n3068) );
  NAND2_X1 U3603 ( .A1(n4143), .A2(n4129), .ZN(n3964) );
  NAND2_X1 U3604 ( .A1(n3973), .A2(n3964), .ZN(n3733) );
  XNOR2_X1 U3605 ( .A(n3734), .B(n2776), .ZN(n4122) );
  OR2_X1 U3606 ( .A1(n3738), .A2(n2777), .ZN(n2782) );
  NAND2_X1 U3607 ( .A1(n3695), .A2(REG1_REG_29__SCAN_IN), .ZN(n2780) );
  NAND2_X1 U3608 ( .A1(n3696), .A2(REG2_REG_29__SCAN_IN), .ZN(n2779) );
  NAND2_X1 U3609 ( .A1(n2536), .A2(REG0_REG_29__SCAN_IN), .ZN(n2778) );
  AND3_X1 U3610 ( .A1(n2780), .A2(n2779), .A3(n2778), .ZN(n2781) );
  INV_X1 U3611 ( .A(n4125), .ZN(n3966) );
  OR2_X1 U3612 ( .A1(n4124), .A2(n4140), .ZN(n3972) );
  INV_X1 U3613 ( .A(n3972), .ZN(n2783) );
  XNOR2_X1 U3614 ( .A(n2225), .B(n2776), .ZN(n2784) );
  NAND2_X1 U3615 ( .A1(n2784), .A2(n4465), .ZN(n4134) );
  AOI22_X1 U3616 ( .A1(n4124), .A2(n4486), .B1(n3068), .B2(n4458), .ZN(n2785)
         );
  OAI211_X1 U3617 ( .C1(n3966), .C2(n4462), .A(n4134), .B(n2785), .ZN(n2786)
         );
  AOI21_X1 U3618 ( .B1(n4122), .B2(n4482), .A(n2786), .ZN(n2796) );
  OAI21_X1 U3619 ( .B1(n2788), .B2(n4129), .A(n2817), .ZN(n4123) );
  OR2_X1 U3620 ( .A1(n4123), .A2(n4484), .ZN(n2791) );
  OR2_X1 U3621 ( .A1(n4828), .A2(n2789), .ZN(n2790) );
  INV_X1 U3622 ( .A(REG0_REG_28__SCAN_IN), .ZN(n2793) );
  OR2_X1 U3623 ( .A1(n4824), .A2(n2793), .ZN(n2794) );
  NAND2_X1 U3624 ( .A1(n2799), .A2(n3973), .ZN(n2800) );
  NAND2_X1 U3625 ( .A1(n3694), .A2(DATAI_29_), .ZN(n3974) );
  XNOR2_X1 U3626 ( .A(n4125), .B(n3974), .ZN(n2811) );
  XNOR2_X1 U3627 ( .A(n2800), .B(n4027), .ZN(n2801) );
  NAND2_X1 U3628 ( .A1(n2801), .A2(n4465), .ZN(n2807) );
  NAND2_X1 U3629 ( .A1(n3695), .A2(REG1_REG_30__SCAN_IN), .ZN(n2804) );
  NAND2_X1 U3630 ( .A1(n3696), .A2(REG2_REG_30__SCAN_IN), .ZN(n2803) );
  NAND2_X1 U3631 ( .A1(n2536), .A2(REG0_REG_30__SCAN_IN), .ZN(n2802) );
  NAND3_X1 U3632 ( .A1(n2804), .A2(n2803), .A3(n2802), .ZN(n3980) );
  AND2_X1 U3633 ( .A1(n4065), .A2(B_REG_SCAN_IN), .ZN(n2805) );
  NOR2_X1 U3634 ( .A1(n4462), .A2(n2805), .ZN(n3700) );
  NAND2_X1 U3635 ( .A1(n3980), .A2(n3700), .ZN(n2806) );
  NAND2_X1 U3636 ( .A1(n4143), .A2(n4486), .ZN(n2808) );
  OAI21_X1 U3637 ( .B1(n3974), .B2(n4477), .A(n2808), .ZN(n2809) );
  NAND2_X1 U3638 ( .A1(n4143), .A2(n3068), .ZN(n2810) );
  NAND2_X1 U3639 ( .A1(n4027), .A2(n2810), .ZN(n2813) );
  INV_X1 U3640 ( .A(n2810), .ZN(n3732) );
  NAND2_X1 U3641 ( .A1(n3732), .A2(n2811), .ZN(n2812) );
  OAI211_X1 U3642 ( .C1(n2813), .C2(n3733), .A(n4482), .B(n2812), .ZN(n2814)
         );
  INV_X1 U3643 ( .A(n3974), .ZN(n3965) );
  NAND2_X1 U3644 ( .A1(n2817), .A2(n3965), .ZN(n2818) );
  NAND2_X1 U3645 ( .A1(n2820), .A2(n2819), .ZN(U3515) );
  NAND2_X1 U3646 ( .A1(n2822), .A2(n2821), .ZN(U3547) );
  NAND2_X1 U3647 ( .A1(n3018), .A2(n2823), .ZN(n2826) );
  AND2_X2 U3648 ( .A1(n2824), .A2(n3313), .ZN(n2983) );
  INV_X1 U3649 ( .A(n2824), .ZN(n3090) );
  AOI22_X1 U3650 ( .A1(n2983), .A2(n3240), .B1(n3090), .B2(n4729), .ZN(n2825)
         );
  NAND2_X1 U3651 ( .A1(n2826), .A2(n2825), .ZN(n3178) );
  INV_X1 U3652 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2828) );
  NAND2_X1 U3653 ( .A1(n2015), .A2(n3240), .ZN(n2830) );
  OAI211_X1 U3654 ( .C1(n2828), .C2(n2824), .A(n2827), .B(n2830), .ZN(n3177)
         );
  NAND2_X1 U3655 ( .A1(n3178), .A2(n3177), .ZN(n3176) );
  NAND2_X1 U3656 ( .A1(n4714), .A2(n4063), .ZN(n3091) );
  NAND2_X4 U3657 ( .A1(n2829), .A2(n3091), .ZN(n3066) );
  NAND2_X1 U3658 ( .A1(n2830), .A2(n3051), .ZN(n2831) );
  NAND2_X1 U3659 ( .A1(n3176), .A2(n2831), .ZN(n3225) );
  NAND2_X1 U3660 ( .A1(n2459), .A2(n2983), .ZN(n2834) );
  NAND2_X1 U3661 ( .A1(n2015), .A2(n2832), .ZN(n2833) );
  NAND2_X1 U3662 ( .A1(n2834), .A2(n2833), .ZN(n2835) );
  XNOR2_X1 U3663 ( .A(n2836), .B(n2838), .ZN(n3226) );
  NAND2_X1 U3664 ( .A1(n3225), .A2(n3226), .ZN(n3224) );
  INV_X1 U3665 ( .A(n2836), .ZN(n2837) );
  NAND2_X1 U3666 ( .A1(n2838), .A2(n2837), .ZN(n2839) );
  NAND2_X1 U3667 ( .A1(n3224), .A2(n2839), .ZN(n3263) );
  INV_X1 U3668 ( .A(n3263), .ZN(n2845) );
  AOI22_X1 U3669 ( .A1(n3018), .A2(n2840), .B1(n2022), .B2(n3291), .ZN(n2846)
         );
  NAND2_X1 U3670 ( .A1(n2840), .A2(n2983), .ZN(n2842) );
  NAND2_X1 U3671 ( .A1(n2015), .A2(n3291), .ZN(n2841) );
  NAND2_X1 U3672 ( .A1(n2842), .A2(n2841), .ZN(n2843) );
  XNOR2_X1 U3673 ( .A(n2846), .B(n2847), .ZN(n3264) );
  INV_X1 U3674 ( .A(n3264), .ZN(n2844) );
  NAND2_X1 U3675 ( .A1(n2845), .A2(n2844), .ZN(n3261) );
  NAND2_X1 U3676 ( .A1(n2847), .A2(n2846), .ZN(n2848) );
  NAND2_X1 U3677 ( .A1(n3261), .A2(n2848), .ZN(n3281) );
  NAND2_X1 U3678 ( .A1(n3344), .A2(n2022), .ZN(n2850) );
  NAND2_X1 U3679 ( .A1(n2015), .A2(n3361), .ZN(n2849) );
  NAND2_X1 U3680 ( .A1(n2850), .A2(n2849), .ZN(n2851) );
  XNOR2_X1 U3681 ( .A(n2851), .B(n3066), .ZN(n2853) );
  AOI22_X1 U3682 ( .A1(n3018), .A2(n3344), .B1(n3063), .B2(n3361), .ZN(n2854)
         );
  XNOR2_X1 U3683 ( .A(n2853), .B(n2854), .ZN(n3282) );
  NAND2_X1 U3684 ( .A1(n3281), .A2(n3282), .ZN(n2857) );
  INV_X1 U3685 ( .A(n2853), .ZN(n2855) );
  NAND2_X1 U3686 ( .A1(n2855), .A2(n2854), .ZN(n2856) );
  NAND2_X1 U3687 ( .A1(n2857), .A2(n2856), .ZN(n3383) );
  INV_X1 U3688 ( .A(n3383), .ZN(n2865) );
  NAND2_X1 U3689 ( .A1(n2861), .A2(n3063), .ZN(n2859) );
  NAND2_X1 U3690 ( .A1(n2015), .A2(n2475), .ZN(n2858) );
  NAND2_X1 U3691 ( .A1(n2859), .A2(n2858), .ZN(n2860) );
  XNOR2_X1 U3692 ( .A(n2860), .B(n3051), .ZN(n2869) );
  AOI22_X1 U3693 ( .A1(n3018), .A2(n2861), .B1(n3063), .B2(n2475), .ZN(n2870)
         );
  XNOR2_X1 U3694 ( .A(n2869), .B(n2870), .ZN(n3433) );
  NAND2_X1 U3695 ( .A1(n2016), .A2(n3063), .ZN(n2863) );
  NAND2_X1 U3696 ( .A1(n2015), .A2(n3464), .ZN(n2862) );
  NAND2_X1 U3697 ( .A1(n2863), .A2(n2862), .ZN(n2864) );
  AOI22_X1 U3698 ( .A1(n3062), .A2(n2016), .B1(n3063), .B2(n3464), .ZN(n2866)
         );
  XNOR2_X1 U3699 ( .A(n2868), .B(n2866), .ZN(n3388) );
  INV_X1 U3700 ( .A(n3388), .ZN(n2873) );
  INV_X1 U3701 ( .A(n2866), .ZN(n2867) );
  NAND2_X1 U3702 ( .A1(n2868), .A2(n2867), .ZN(n2874) );
  INV_X1 U3703 ( .A(n2869), .ZN(n2872) );
  INV_X1 U3704 ( .A(n2870), .ZN(n2871) );
  NAND2_X1 U3705 ( .A1(n2872), .A2(n2871), .ZN(n3384) );
  OR2_X1 U3706 ( .A1(n2873), .A2(n3384), .ZN(n3385) );
  AND2_X1 U3707 ( .A1(n2874), .A2(n3385), .ZN(n2875) );
  NAND2_X2 U3708 ( .A1(n3386), .A2(n2875), .ZN(n3399) );
  NAND2_X1 U3709 ( .A1(n3062), .A2(n3447), .ZN(n2877) );
  NAND2_X1 U3710 ( .A1(n3063), .A2(n3411), .ZN(n2876) );
  NAND2_X1 U3711 ( .A1(n2877), .A2(n2876), .ZN(n3397) );
  NAND2_X1 U3712 ( .A1(n3447), .A2(n3063), .ZN(n2879) );
  NAND2_X1 U3713 ( .A1(n2015), .A2(n3411), .ZN(n2878) );
  NAND2_X1 U3714 ( .A1(n2879), .A2(n2878), .ZN(n2880) );
  XNOR2_X1 U3715 ( .A(n2880), .B(n3066), .ZN(n3396) );
  NAND2_X1 U3716 ( .A1(n4075), .A2(n3063), .ZN(n2882) );
  NAND2_X1 U3717 ( .A1(n2015), .A2(n3456), .ZN(n2881) );
  NAND2_X1 U3718 ( .A1(n2882), .A2(n2881), .ZN(n2883) );
  XNOR2_X1 U3719 ( .A(n2883), .B(n3066), .ZN(n2886) );
  AOI22_X1 U3720 ( .A1(n3018), .A2(n4075), .B1(n3063), .B2(n3456), .ZN(n2884)
         );
  XNOR2_X1 U3721 ( .A(n2886), .B(n2884), .ZN(n3439) );
  INV_X1 U3722 ( .A(n2884), .ZN(n2885) );
  NAND2_X1 U3723 ( .A1(n2886), .A2(n2885), .ZN(n2887) );
  NAND2_X1 U3724 ( .A1(n4074), .A2(n3063), .ZN(n2889) );
  NAND2_X1 U3725 ( .A1(n3013), .A2(n3516), .ZN(n2888) );
  NAND2_X1 U3726 ( .A1(n2889), .A2(n2888), .ZN(n2890) );
  XNOR2_X1 U3727 ( .A(n2890), .B(n3066), .ZN(n2893) );
  NAND2_X1 U3728 ( .A1(n3062), .A2(n4074), .ZN(n2892) );
  NAND2_X1 U3729 ( .A1(n3063), .A2(n3516), .ZN(n2891) );
  NAND2_X1 U3730 ( .A1(n2892), .A2(n2891), .ZN(n2894) );
  AND2_X1 U3731 ( .A1(n2893), .A2(n2894), .ZN(n3495) );
  INV_X1 U3732 ( .A(n2893), .ZN(n2896) );
  INV_X1 U3733 ( .A(n2894), .ZN(n2895) );
  NAND2_X1 U3734 ( .A1(n2896), .A2(n2895), .ZN(n3494) );
  NAND2_X1 U3735 ( .A1(n3525), .A2(n2022), .ZN(n2898) );
  NAND2_X1 U3736 ( .A1(n3013), .A2(n3606), .ZN(n2897) );
  NAND2_X1 U3737 ( .A1(n2898), .A2(n2897), .ZN(n2899) );
  XNOR2_X1 U3738 ( .A(n2899), .B(n3066), .ZN(n2900) );
  AOI22_X1 U3739 ( .A1(n3018), .A2(n3525), .B1(n3063), .B2(n3606), .ZN(n2901)
         );
  XNOR2_X1 U3740 ( .A(n2900), .B(n2901), .ZN(n3549) );
  NAND2_X1 U3741 ( .A1(n3548), .A2(n3549), .ZN(n2904) );
  INV_X1 U3742 ( .A(n2900), .ZN(n2902) );
  NAND2_X1 U3743 ( .A1(n2902), .A2(n2901), .ZN(n2903) );
  NAND2_X1 U3744 ( .A1(n2904), .A2(n2903), .ZN(n3675) );
  INV_X1 U3745 ( .A(n3675), .ZN(n2909) );
  NAND2_X1 U3746 ( .A1(n4485), .A2(n2022), .ZN(n2906) );
  NAND2_X1 U3747 ( .A1(n3013), .A2(n3668), .ZN(n2905) );
  NAND2_X1 U3748 ( .A1(n2906), .A2(n2905), .ZN(n2907) );
  XNOR2_X1 U3749 ( .A(n2907), .B(n3051), .ZN(n2910) );
  AOI22_X1 U3750 ( .A1(n3018), .A2(n4485), .B1(n3063), .B2(n3668), .ZN(n2911)
         );
  XNOR2_X1 U3751 ( .A(n2910), .B(n2911), .ZN(n3676) );
  NAND2_X2 U3752 ( .A1(n2909), .A2(n2908), .ZN(n3673) );
  INV_X1 U3753 ( .A(n2910), .ZN(n2913) );
  INV_X1 U3754 ( .A(n2911), .ZN(n2912) );
  NAND2_X1 U3755 ( .A1(n2913), .A2(n2912), .ZN(n2914) );
  NAND2_X1 U3756 ( .A1(n3062), .A2(n4473), .ZN(n2916) );
  NAND2_X1 U3757 ( .A1(n3566), .A2(n2022), .ZN(n2915) );
  NAND2_X1 U3758 ( .A1(n2916), .A2(n2915), .ZN(n3617) );
  NAND2_X1 U3759 ( .A1(n4473), .A2(n3063), .ZN(n2918) );
  NAND2_X1 U3760 ( .A1(n3566), .A2(n3013), .ZN(n2917) );
  NAND2_X1 U3761 ( .A1(n2918), .A2(n2917), .ZN(n2919) );
  XNOR2_X1 U3762 ( .A(n2919), .B(n3066), .ZN(n3616) );
  NAND2_X1 U3763 ( .A1(n3619), .A2(n3617), .ZN(n2920) );
  NAND2_X1 U3764 ( .A1(n4073), .A2(n3063), .ZN(n2922) );
  NAND2_X1 U3765 ( .A1(n3590), .A2(n3013), .ZN(n2921) );
  NAND2_X1 U3766 ( .A1(n2922), .A2(n2921), .ZN(n2923) );
  XNOR2_X1 U3767 ( .A(n2923), .B(n3066), .ZN(n2926) );
  NAND2_X1 U3768 ( .A1(n3062), .A2(n4073), .ZN(n2925) );
  NAND2_X1 U3769 ( .A1(n3590), .A2(n2022), .ZN(n2924) );
  NAND2_X1 U3770 ( .A1(n2925), .A2(n2924), .ZN(n2927) );
  INV_X1 U3771 ( .A(n2926), .ZN(n2929) );
  INV_X1 U3772 ( .A(n2927), .ZN(n2928) );
  NAND2_X1 U3773 ( .A1(n2929), .A2(n2928), .ZN(n3794) );
  NAND2_X1 U3774 ( .A1(n4450), .A2(n2022), .ZN(n2931) );
  NAND2_X1 U3775 ( .A1(n3013), .A2(n4459), .ZN(n2930) );
  NAND2_X1 U3776 ( .A1(n2931), .A2(n2930), .ZN(n2932) );
  XNOR2_X1 U3777 ( .A(n2932), .B(n3066), .ZN(n2942) );
  NAND2_X1 U3778 ( .A1(n3018), .A2(n4450), .ZN(n2934) );
  NAND2_X1 U3779 ( .A1(n3063), .A2(n4459), .ZN(n2933) );
  NAND2_X1 U3780 ( .A1(n2934), .A2(n2933), .ZN(n2943) );
  NAND2_X1 U3781 ( .A1(n2942), .A2(n2943), .ZN(n3753) );
  NAND2_X1 U3782 ( .A1(n4474), .A2(n2022), .ZN(n2936) );
  NAND2_X1 U3783 ( .A1(n3013), .A2(n3627), .ZN(n2935) );
  NAND2_X1 U3784 ( .A1(n2936), .A2(n2935), .ZN(n2937) );
  XNOR2_X1 U3785 ( .A(n2937), .B(n3066), .ZN(n3850) );
  NAND2_X1 U3786 ( .A1(n3062), .A2(n4474), .ZN(n2939) );
  NAND2_X1 U3787 ( .A1(n3063), .A2(n3627), .ZN(n2938) );
  NAND2_X1 U3788 ( .A1(n2939), .A2(n2938), .ZN(n3849) );
  NAND2_X1 U3789 ( .A1(n3850), .A2(n3849), .ZN(n2940) );
  AND2_X1 U3790 ( .A1(n3753), .A2(n2940), .ZN(n2941) );
  NAND2_X1 U3791 ( .A1(n3747), .A2(n2941), .ZN(n2948) );
  INV_X1 U3792 ( .A(n3849), .ZN(n3748) );
  INV_X1 U3793 ( .A(n3850), .ZN(n3749) );
  NAND3_X1 U3794 ( .A1(n3753), .A2(n3748), .A3(n3749), .ZN(n2946) );
  INV_X1 U3795 ( .A(n2942), .ZN(n2945) );
  INV_X1 U3796 ( .A(n2943), .ZN(n2944) );
  NAND2_X1 U3797 ( .A1(n2945), .A2(n2944), .ZN(n3752) );
  AND2_X1 U3798 ( .A1(n2946), .A2(n3752), .ZN(n2947) );
  NAND2_X1 U3799 ( .A1(n4432), .A2(n3063), .ZN(n2950) );
  NAND2_X1 U3800 ( .A1(n3013), .A2(n4352), .ZN(n2949) );
  NAND2_X1 U3801 ( .A1(n2950), .A2(n2949), .ZN(n2951) );
  XNOR2_X1 U3802 ( .A(n2951), .B(n3066), .ZN(n3808) );
  NAND2_X1 U3803 ( .A1(n4432), .A2(n3062), .ZN(n2953) );
  NAND2_X1 U3804 ( .A1(n3063), .A2(n4352), .ZN(n2952) );
  NAND2_X1 U3805 ( .A1(n2953), .A2(n2952), .ZN(n2967) );
  NAND2_X1 U3806 ( .A1(n3808), .A2(n2967), .ZN(n2962) );
  NAND2_X1 U3807 ( .A1(n4440), .A2(n3063), .ZN(n2955) );
  NAND2_X1 U3808 ( .A1(n3013), .A2(n4449), .ZN(n2954) );
  NAND2_X1 U3809 ( .A1(n2955), .A2(n2954), .ZN(n2956) );
  XNOR2_X1 U3810 ( .A(n2956), .B(n3066), .ZN(n3806) );
  NAND2_X1 U3811 ( .A1(n3018), .A2(n4440), .ZN(n2958) );
  NAND2_X1 U3812 ( .A1(n3063), .A2(n4449), .ZN(n2957) );
  NAND2_X1 U3813 ( .A1(n2958), .A2(n2957), .ZN(n3896) );
  NAND2_X1 U3814 ( .A1(n3806), .A2(n3896), .ZN(n2959) );
  AND2_X1 U3815 ( .A1(n2962), .A2(n2959), .ZN(n2960) );
  INV_X1 U3816 ( .A(n3896), .ZN(n3816) );
  INV_X1 U3817 ( .A(n3806), .ZN(n2961) );
  NAND3_X1 U3818 ( .A1(n2962), .A2(n3816), .A3(n2961), .ZN(n2970) );
  NAND2_X1 U3819 ( .A1(n4441), .A2(n2022), .ZN(n2964) );
  NAND2_X1 U3820 ( .A1(n3013), .A2(n4431), .ZN(n2963) );
  NAND2_X1 U3821 ( .A1(n2964), .A2(n2963), .ZN(n2965) );
  XNOR2_X1 U3822 ( .A(n2965), .B(n3051), .ZN(n3820) );
  NOR2_X1 U3823 ( .A1(n2852), .A2(n4335), .ZN(n2966) );
  AOI21_X1 U3824 ( .B1(n4441), .B2(n3018), .A(n2966), .ZN(n2971) );
  NAND2_X1 U3825 ( .A1(n3820), .A2(n2971), .ZN(n2969) );
  INV_X1 U3826 ( .A(n3808), .ZN(n2968) );
  INV_X1 U3827 ( .A(n2967), .ZN(n3807) );
  NAND2_X1 U3828 ( .A1(n2968), .A2(n3807), .ZN(n3817) );
  INV_X1 U3829 ( .A(n3820), .ZN(n2972) );
  INV_X1 U3830 ( .A(n2971), .ZN(n3819) );
  AND2_X1 U3831 ( .A1(n2972), .A2(n3819), .ZN(n2973) );
  NAND2_X1 U3832 ( .A1(n4292), .A2(n2022), .ZN(n2976) );
  NAND2_X1 U3833 ( .A1(n3013), .A2(n4308), .ZN(n2975) );
  NAND2_X1 U3834 ( .A1(n2976), .A2(n2975), .ZN(n2977) );
  XNOR2_X1 U3835 ( .A(n2977), .B(n3066), .ZN(n2986) );
  NAND2_X1 U3836 ( .A1(n4292), .A2(n3062), .ZN(n2979) );
  NAND2_X1 U3837 ( .A1(n3063), .A2(n4308), .ZN(n2978) );
  NAND2_X1 U3838 ( .A1(n2979), .A2(n2978), .ZN(n2987) );
  NAND2_X1 U3839 ( .A1(n2986), .A2(n2987), .ZN(n3873) );
  NAND2_X1 U3840 ( .A1(n4416), .A2(n3063), .ZN(n2981) );
  NAND2_X1 U3841 ( .A1(n3013), .A2(n4291), .ZN(n2980) );
  NAND2_X1 U3842 ( .A1(n2981), .A2(n2980), .ZN(n2982) );
  XNOR2_X1 U3843 ( .A(n2982), .B(n3066), .ZN(n2991) );
  INV_X1 U3844 ( .A(n2983), .ZN(n3035) );
  NOR2_X1 U3845 ( .A1(n2852), .A2(n4301), .ZN(n2984) );
  AOI21_X1 U3846 ( .B1(n4416), .B2(n3062), .A(n2984), .ZN(n2992) );
  XNOR2_X1 U3847 ( .A(n2991), .B(n2992), .ZN(n3777) );
  AND2_X1 U3848 ( .A1(n3873), .A2(n3777), .ZN(n2985) );
  INV_X1 U3849 ( .A(n3777), .ZN(n2990) );
  INV_X1 U3850 ( .A(n2986), .ZN(n2989) );
  INV_X1 U3851 ( .A(n2987), .ZN(n2988) );
  NAND2_X1 U3852 ( .A1(n2989), .A2(n2988), .ZN(n3872) );
  INV_X1 U3853 ( .A(n2991), .ZN(n2993) );
  NAND2_X1 U3854 ( .A1(n2995), .A2(n2994), .ZN(n3839) );
  NAND2_X1 U3855 ( .A1(n4405), .A2(n3063), .ZN(n2997) );
  NAND2_X1 U3856 ( .A1(n3013), .A2(n4415), .ZN(n2996) );
  NAND2_X1 U3857 ( .A1(n2997), .A2(n2996), .ZN(n2998) );
  XNOR2_X1 U3858 ( .A(n2998), .B(n3066), .ZN(n3001) );
  NAND2_X1 U3859 ( .A1(n4405), .A2(n3062), .ZN(n3000) );
  NAND2_X1 U3860 ( .A1(n2022), .A2(n4415), .ZN(n2999) );
  NAND2_X1 U3861 ( .A1(n3000), .A2(n2999), .ZN(n3002) );
  NAND2_X1 U3862 ( .A1(n3001), .A2(n3002), .ZN(n3840) );
  INV_X1 U3863 ( .A(n3001), .ZN(n3004) );
  INV_X1 U3864 ( .A(n3002), .ZN(n3003) );
  NAND2_X1 U3865 ( .A1(n3004), .A2(n3003), .ZN(n3842) );
  NAND2_X1 U3866 ( .A1(n4414), .A2(n3063), .ZN(n3006) );
  NAND2_X1 U3867 ( .A1(n3013), .A2(n4404), .ZN(n3005) );
  NAND2_X1 U3868 ( .A1(n3006), .A2(n3005), .ZN(n3007) );
  XNOR2_X1 U3869 ( .A(n3007), .B(n3051), .ZN(n3785) );
  NOR2_X1 U3870 ( .A1(n2852), .A2(n4245), .ZN(n3008) );
  AOI21_X1 U3871 ( .B1(n4414), .B2(n3062), .A(n3008), .ZN(n3022) );
  AND2_X1 U3872 ( .A1(n3785), .A2(n3022), .ZN(n3764) );
  NAND2_X1 U3873 ( .A1(n4224), .A2(n3063), .ZN(n3010) );
  NAND2_X1 U3874 ( .A1(n3013), .A2(n4207), .ZN(n3009) );
  NAND2_X1 U3875 ( .A1(n3010), .A2(n3009), .ZN(n3011) );
  XNOR2_X1 U3876 ( .A(n3011), .B(n3066), .ZN(n3034) );
  NOR2_X1 U3877 ( .A1(n2852), .A2(n4216), .ZN(n3012) );
  AOI21_X1 U3878 ( .B1(n4224), .B2(n3062), .A(n3012), .ZN(n3032) );
  XNOR2_X1 U3879 ( .A(n3034), .B(n3032), .ZN(n3767) );
  NAND2_X1 U3880 ( .A1(n4247), .A2(n3063), .ZN(n3015) );
  NAND2_X1 U3881 ( .A1(n3013), .A2(n4232), .ZN(n3014) );
  NAND2_X1 U3882 ( .A1(n3015), .A2(n3014), .ZN(n3016) );
  XNOR2_X1 U3883 ( .A(n3016), .B(n3051), .ZN(n3021) );
  NOR2_X1 U3884 ( .A1(n2852), .A2(n3867), .ZN(n3017) );
  AOI21_X1 U3885 ( .B1(n4247), .B2(n3018), .A(n3017), .ZN(n3020) );
  NAND2_X1 U3886 ( .A1(n3021), .A2(n3020), .ZN(n3768) );
  NAND2_X1 U3887 ( .A1(n3767), .A2(n3768), .ZN(n3026) );
  XNOR2_X1 U3888 ( .A(n3021), .B(n3020), .ZN(n3864) );
  INV_X1 U3889 ( .A(n3864), .ZN(n3024) );
  INV_X1 U3890 ( .A(n3785), .ZN(n3023) );
  INV_X1 U3891 ( .A(n3022), .ZN(n3784) );
  NAND2_X1 U3892 ( .A1(n3023), .A2(n3784), .ZN(n3765) );
  AND2_X1 U3893 ( .A1(n3024), .A2(n3765), .ZN(n3025) );
  NOR2_X1 U3894 ( .A1(n3026), .A2(n3025), .ZN(n3710) );
  NAND2_X1 U3895 ( .A1(n4387), .A2(n3063), .ZN(n3028) );
  NAND2_X1 U3896 ( .A1(n3013), .A2(n4377), .ZN(n3027) );
  NAND2_X1 U3897 ( .A1(n3028), .A2(n3027), .ZN(n3029) );
  XNOR2_X1 U3898 ( .A(n3029), .B(n3066), .ZN(n3716) );
  NAND2_X1 U3899 ( .A1(n4387), .A2(n3062), .ZN(n3031) );
  NAND2_X1 U3900 ( .A1(n3063), .A2(n4377), .ZN(n3030) );
  NAND2_X1 U3901 ( .A1(n3031), .A2(n3030), .ZN(n3715) );
  NAND2_X1 U3902 ( .A1(n3716), .A2(n3715), .ZN(n3714) );
  INV_X1 U3903 ( .A(n3032), .ZN(n3033) );
  NAND2_X1 U3904 ( .A1(n3034), .A2(n3033), .ZN(n3713) );
  NOR2_X1 U3905 ( .A1(n2852), .A2(n4195), .ZN(n3036) );
  AOI21_X1 U3906 ( .B1(n4378), .B2(n3062), .A(n3036), .ZN(n3712) );
  NAND2_X1 U3907 ( .A1(n3713), .A2(n3712), .ZN(n3709) );
  NAND2_X1 U3908 ( .A1(n4378), .A2(n3063), .ZN(n3038) );
  NAND2_X1 U3909 ( .A1(n3013), .A2(n4386), .ZN(n3037) );
  NAND2_X1 U3910 ( .A1(n3038), .A2(n3037), .ZN(n3039) );
  XNOR2_X1 U3911 ( .A(n3039), .B(n3051), .ZN(n3044) );
  NAND2_X1 U3912 ( .A1(n3713), .A2(n3044), .ZN(n3040) );
  NAND2_X1 U3913 ( .A1(n3709), .A2(n3040), .ZN(n3041) );
  NAND2_X1 U3914 ( .A1(n3762), .A2(n2228), .ZN(n3048) );
  INV_X1 U3915 ( .A(n3044), .ZN(n3830) );
  INV_X1 U3916 ( .A(n3712), .ZN(n3042) );
  OAI21_X1 U3917 ( .B1(n3830), .B2(n3042), .A(n3715), .ZN(n3046) );
  INV_X1 U3918 ( .A(n3716), .ZN(n3045) );
  NOR2_X1 U3919 ( .A1(n3715), .A2(n3042), .ZN(n3043) );
  AOI22_X1 U3920 ( .A1(n3046), .A2(n3045), .B1(n3044), .B2(n3043), .ZN(n3047)
         );
  NAND2_X1 U3921 ( .A1(n4137), .A2(n3063), .ZN(n3050) );
  NAND2_X1 U3922 ( .A1(n3013), .A2(n4154), .ZN(n3049) );
  NAND2_X1 U3923 ( .A1(n3050), .A2(n3049), .ZN(n3052) );
  XNOR2_X1 U3924 ( .A(n3052), .B(n3051), .ZN(n3057) );
  INV_X1 U3925 ( .A(n3057), .ZN(n3055) );
  NOR2_X1 U3926 ( .A1(n2852), .A2(n4159), .ZN(n3053) );
  AOI21_X1 U3927 ( .B1(n4137), .B2(n3062), .A(n3053), .ZN(n3056) );
  INV_X1 U3928 ( .A(n3056), .ZN(n3054) );
  NAND2_X1 U3929 ( .A1(n3055), .A2(n3054), .ZN(n3882) );
  AND2_X1 U3930 ( .A1(n3057), .A2(n3056), .ZN(n3881) );
  NAND2_X1 U3931 ( .A1(n4124), .A2(n3063), .ZN(n3059) );
  NAND2_X1 U3932 ( .A1(n3013), .A2(n3968), .ZN(n3058) );
  NAND2_X1 U3933 ( .A1(n3059), .A2(n3058), .ZN(n3060) );
  XNOR2_X1 U3934 ( .A(n3060), .B(n3066), .ZN(n3083) );
  NOR2_X1 U3935 ( .A1(n2852), .A2(n4140), .ZN(n3061) );
  AOI21_X1 U3936 ( .B1(n4124), .B2(n3062), .A(n3061), .ZN(n3081) );
  XNOR2_X1 U3937 ( .A(n3083), .B(n3081), .ZN(n3724) );
  NAND2_X1 U3938 ( .A1(n3725), .A2(n3724), .ZN(n3111) );
  NAND2_X1 U3939 ( .A1(n4143), .A2(n3062), .ZN(n3065) );
  NAND2_X1 U3940 ( .A1(n3063), .A2(n3068), .ZN(n3064) );
  NAND2_X1 U3941 ( .A1(n3065), .A2(n3064), .ZN(n3067) );
  XNOR2_X1 U3942 ( .A(n3067), .B(n3066), .ZN(n3070) );
  AOI22_X1 U3943 ( .A1(n4143), .A2(n2022), .B1(n3013), .B2(n3068), .ZN(n3069)
         );
  XNOR2_X1 U3944 ( .A(n3070), .B(n3069), .ZN(n3105) );
  INV_X1 U3945 ( .A(n3105), .ZN(n3080) );
  AND2_X1 U3946 ( .A1(n3071), .A2(n3130), .ZN(n3308) );
  NAND3_X1 U3947 ( .A1(n3308), .A2(n3072), .A3(n3306), .ZN(n3101) );
  NAND2_X1 U3948 ( .A1(n3074), .A2(n3073), .ZN(n3077) );
  INV_X1 U3949 ( .A(n3075), .ZN(n3076) );
  NAND2_X1 U3950 ( .A1(n3077), .A2(n3076), .ZN(n3086) );
  INV_X1 U3951 ( .A(n3086), .ZN(n3078) );
  NAND2_X1 U3952 ( .A1(n3216), .A2(n3078), .ZN(n3079) );
  NAND2_X1 U3953 ( .A1(n3080), .A2(n3876), .ZN(n3110) );
  INV_X1 U3954 ( .A(n3081), .ZN(n3082) );
  NAND2_X1 U3955 ( .A1(n3083), .A2(n3082), .ZN(n3104) );
  NAND2_X1 U3956 ( .A1(n3111), .A2(n3084), .ZN(n3109) );
  INV_X1 U3957 ( .A(n3085), .ZN(n4126) );
  NAND2_X1 U3958 ( .A1(n3086), .A2(n4477), .ZN(n3087) );
  NAND2_X1 U3959 ( .A1(n3101), .A2(n3087), .ZN(n3089) );
  NAND2_X1 U3960 ( .A1(n3089), .A2(n3088), .ZN(n3214) );
  OAI21_X1 U3961 ( .B1(n3214), .B2(n3090), .A(STATE_REG_SCAN_IN), .ZN(n3095)
         );
  INV_X1 U3962 ( .A(n3091), .ZN(n3092) );
  AND2_X1 U3963 ( .A1(n4805), .A2(n3092), .ZN(n3093) );
  NAND2_X1 U3964 ( .A1(n3101), .A2(n3100), .ZN(n3215) );
  AND2_X1 U3965 ( .A1(n3215), .A2(n4070), .ZN(n3094) );
  NAND2_X1 U3966 ( .A1(n3216), .A2(n4458), .ZN(n3096) );
  OR2_X1 U3967 ( .A1(n3101), .A2(n3096), .ZN(n3098) );
  NAND2_X1 U3968 ( .A1(n3100), .A2(n3179), .ZN(n3099) );
  NAND2_X1 U3969 ( .A1(n3100), .A2(n4713), .ZN(n4067) );
  AOI22_X1 U3970 ( .A1(n3890), .A2(n4125), .B1(n4124), .B2(n3902), .ZN(n3103)
         );
  NAND2_X1 U3971 ( .A1(U3149), .A2(REG3_REG_28__SCAN_IN), .ZN(n3102) );
  OAI211_X1 U3972 ( .C1(n3900), .C2(n4129), .A(n3103), .B(n3102), .ZN(n3107)
         );
  NOR3_X1 U3973 ( .A1(n3105), .A2(n3907), .A3(n3104), .ZN(n3106) );
  AOI211_X1 U3974 ( .C1(n4126), .C2(n3904), .A(n3107), .B(n3106), .ZN(n3108)
         );
  OAI211_X1 U3975 ( .C1(n3111), .C2(n3110), .A(n3109), .B(n3108), .ZN(U3217)
         );
  INV_X1 U3976 ( .A(n4805), .ZN(n3127) );
  NOR2_X1 U3977 ( .A1(n2824), .A2(n3127), .ZN(U4043) );
  INV_X1 U3978 ( .A(DATAI_26_), .ZN(n3113) );
  NAND2_X1 U3979 ( .A1(n3126), .A2(STATE_REG_SCAN_IN), .ZN(n3112) );
  OAI21_X1 U3980 ( .B1(STATE_REG_SCAN_IN), .B2(n3113), .A(n3112), .ZN(U3326)
         );
  INV_X1 U3981 ( .A(DATAI_17_), .ZN(n4623) );
  NAND2_X1 U3982 ( .A1(n4109), .A2(STATE_REG_SCAN_IN), .ZN(n3114) );
  OAI21_X1 U3983 ( .B1(STATE_REG_SCAN_IN), .B2(n4623), .A(n3114), .ZN(U3335)
         );
  INV_X1 U3984 ( .A(DATAI_13_), .ZN(n4559) );
  NAND2_X1 U3985 ( .A1(n3659), .A2(STATE_REG_SCAN_IN), .ZN(n3115) );
  OAI21_X1 U3986 ( .B1(STATE_REG_SCAN_IN), .B2(n4559), .A(n3115), .ZN(U3339)
         );
  INV_X1 U3987 ( .A(DATAI_27_), .ZN(n3117) );
  NAND2_X1 U3988 ( .A1(n4065), .A2(STATE_REG_SCAN_IN), .ZN(n3116) );
  OAI21_X1 U3989 ( .B1(STATE_REG_SCAN_IN), .B2(n3117), .A(n3116), .ZN(U3325)
         );
  INV_X1 U3990 ( .A(DATAI_25_), .ZN(n3120) );
  NAND2_X1 U3991 ( .A1(n3118), .A2(STATE_REG_SCAN_IN), .ZN(n3119) );
  OAI21_X1 U3992 ( .B1(STATE_REG_SCAN_IN), .B2(n3120), .A(n3119), .ZN(U3327)
         );
  INV_X1 U3993 ( .A(DATAI_24_), .ZN(n3122) );
  NAND2_X1 U3994 ( .A1(n2748), .A2(STATE_REG_SCAN_IN), .ZN(n3121) );
  OAI21_X1 U3995 ( .B1(STATE_REG_SCAN_IN), .B2(n3122), .A(n3121), .ZN(U3328)
         );
  INV_X1 U3996 ( .A(DATAI_31_), .ZN(n3124) );
  OR4_X1 U3997 ( .A1(n2436), .A2(IR_REG_30__SCAN_IN), .A3(U3149), .A4(n2080), 
        .ZN(n3123) );
  OAI21_X1 U3998 ( .B1(STATE_REG_SCAN_IN), .B2(n3124), .A(n3123), .ZN(U3321)
         );
  NOR3_X1 U3999 ( .A1(n3127), .A2(n2748), .A3(n3126), .ZN(n3128) );
  AOI21_X1 U4000 ( .B1(n4804), .B2(n3129), .A(n3128), .ZN(U3458) );
  INV_X1 U4001 ( .A(n3130), .ZN(n3131) );
  AOI22_X1 U4002 ( .A1(n4804), .A2(n3132), .B1(n3131), .B2(n4805), .ZN(U3459)
         );
  NOR2_X1 U4003 ( .A1(n4765), .A2(U4043), .ZN(U3148) );
  INV_X1 U4004 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n4622) );
  NAND2_X1 U4005 ( .A1(n3344), .A2(U4043), .ZN(n3134) );
  OAI21_X1 U4006 ( .B1(n4077), .B2(n4622), .A(n3134), .ZN(U3553) );
  INV_X1 U4007 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4552) );
  NAND2_X1 U4008 ( .A1(n3980), .A2(U4043), .ZN(n3135) );
  OAI21_X1 U4009 ( .B1(n4077), .B2(n4552), .A(n3135), .ZN(U3580) );
  INV_X1 U4010 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n4615) );
  NAND2_X1 U4011 ( .A1(n3447), .A2(n4077), .ZN(n3136) );
  OAI21_X1 U4012 ( .B1(n4615), .B2(U4043), .A(n3136), .ZN(U3556) );
  INV_X1 U4013 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n4601) );
  NAND2_X1 U4014 ( .A1(n3525), .A2(n4077), .ZN(n3137) );
  OAI21_X1 U4015 ( .B1(n4601), .B2(U4043), .A(n3137), .ZN(U3559) );
  INV_X1 U4016 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n4574) );
  NAND2_X1 U4017 ( .A1(n4440), .A2(U4043), .ZN(n3138) );
  OAI21_X1 U4018 ( .B1(n4077), .B2(n4574), .A(n3138), .ZN(U3565) );
  XOR2_X1 U4019 ( .A(n3139), .B(REG2_REG_3__SCAN_IN), .Z(n3144) );
  AOI211_X1 U4020 ( .C1(n3142), .C2(n3141), .A(n3140), .B(n4113), .ZN(n3143)
         );
  AOI21_X1 U4021 ( .B1(n4096), .B2(n3144), .A(n3143), .ZN(n3146) );
  NOR2_X1 U4022 ( .A1(STATE_REG_SCAN_IN), .A2(n2460), .ZN(n3280) );
  AOI21_X1 U4023 ( .B1(n4765), .B2(ADDR_REG_3__SCAN_IN), .A(n3280), .ZN(n3145)
         );
  OAI211_X1 U4024 ( .C1(n3147), .C2(n4775), .A(n3146), .B(n3145), .ZN(U3243)
         );
  INV_X1 U4025 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3148) );
  AOI21_X1 U4026 ( .B1(n4065), .B2(n3148), .A(n3179), .ZN(n3182) );
  OAI21_X1 U4027 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4065), .A(n3182), .ZN(n3149)
         );
  MUX2_X1 U4028 ( .A(n3149), .B(n3182), .S(n4729), .Z(n3151) );
  INV_X1 U4029 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3150) );
  OAI22_X1 U4030 ( .A1(n3152), .A2(n3151), .B1(STATE_REG_SCAN_IN), .B2(n3150), 
        .ZN(n3154) );
  NOR3_X1 U4031 ( .A1(n4113), .A2(REG1_REG_0__SCAN_IN), .A3(n2081), .ZN(n3153)
         );
  AOI211_X1 U4032 ( .C1(n4765), .C2(ADDR_REG_0__SCAN_IN), .A(n3154), .B(n3153), 
        .ZN(n3155) );
  INV_X1 U4033 ( .A(n3155), .ZN(U3240) );
  AOI211_X1 U4034 ( .C1(n2058), .C2(n3157), .A(n4113), .B(n3156), .ZN(n3165)
         );
  OAI211_X1 U4035 ( .C1(n3160), .C2(n3159), .A(n4096), .B(n3158), .ZN(n3162)
         );
  AND2_X1 U4036 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3392) );
  AOI21_X1 U4037 ( .B1(n4765), .B2(ADDR_REG_5__SCAN_IN), .A(n3392), .ZN(n3161)
         );
  OAI211_X1 U4038 ( .C1(n4775), .C2(n3163), .A(n3162), .B(n3161), .ZN(n3164)
         );
  OR2_X1 U4039 ( .A1(n3165), .A2(n3164), .ZN(U3245) );
  INV_X1 U4040 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n4620) );
  NAND2_X1 U4041 ( .A1(n4414), .A2(U4043), .ZN(n3166) );
  OAI21_X1 U4042 ( .B1(n4077), .B2(n4620), .A(n3166), .ZN(U3571) );
  XNOR2_X1 U40430 ( .A(n3167), .B(REG2_REG_6__SCAN_IN), .ZN(n3175) );
  OAI211_X1 U4044 ( .C1(n3169), .C2(REG1_REG_6__SCAN_IN), .A(n3168), .B(n4770), 
        .ZN(n3174) );
  NAND2_X1 U4045 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3400) );
  INV_X1 U4046 ( .A(n3400), .ZN(n3172) );
  NOR2_X1 U4047 ( .A1(n4775), .A2(n3170), .ZN(n3171) );
  AOI211_X1 U4048 ( .C1(n4765), .C2(ADDR_REG_6__SCAN_IN), .A(n3172), .B(n3171), 
        .ZN(n3173) );
  OAI211_X1 U4049 ( .C1(n3175), .C2(n4762), .A(n3174), .B(n3173), .ZN(U3246)
         );
  OAI21_X1 U4050 ( .B1(n3178), .B2(n3177), .A(n3176), .ZN(n3218) );
  NAND2_X1 U4051 ( .A1(n4729), .A2(REG2_REG_0__SCAN_IN), .ZN(n4081) );
  AOI21_X1 U4052 ( .B1(n4065), .B2(n4081), .A(n3179), .ZN(n3180) );
  OAI21_X1 U4053 ( .B1(n3218), .B2(n4065), .A(n3180), .ZN(n3181) );
  OAI211_X1 U4054 ( .C1(n4729), .C2(n3182), .A(n3181), .B(U4043), .ZN(n3252)
         );
  INV_X1 U4055 ( .A(n3252), .ZN(n3197) );
  OAI211_X1 U4056 ( .C1(n3185), .C2(n3184), .A(n4770), .B(n3183), .ZN(n3195)
         );
  INV_X1 U4057 ( .A(n3186), .ZN(n3189) );
  NAND3_X1 U4058 ( .A1(n3189), .A2(n3187), .A3(n3188), .ZN(n3190) );
  NAND3_X1 U4059 ( .A1(n4096), .A2(n3191), .A3(n3190), .ZN(n3194) );
  INV_X1 U4060 ( .A(n4775), .ZN(n4110) );
  NAND2_X1 U4061 ( .A1(n4110), .A2(n4727), .ZN(n3193) );
  AOI22_X1 U4062 ( .A1(n4765), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3192) );
  NAND4_X1 U4063 ( .A1(n3195), .A2(n3194), .A3(n3193), .A4(n3192), .ZN(n3196)
         );
  OR2_X1 U4064 ( .A1(n3197), .A2(n3196), .ZN(U3242) );
  INV_X1 U4065 ( .A(n4644), .ZN(n4821) );
  INV_X1 U4066 ( .A(n3240), .ZN(n3222) );
  NAND2_X1 U4067 ( .A1(n2823), .A2(n3222), .ZN(n3910) );
  NAND2_X1 U4068 ( .A1(n3198), .A2(n3910), .ZN(n4783) );
  NOR2_X1 U4069 ( .A1(n3222), .A2(n3199), .ZN(n4787) );
  INV_X1 U4070 ( .A(n2459), .ZN(n3312) );
  INV_X1 U4071 ( .A(n3561), .ZN(n3507) );
  OAI21_X1 U4072 ( .B1(n3507), .B2(n4465), .A(n4783), .ZN(n3200) );
  OAI21_X1 U4073 ( .B1(n3312), .B2(n4462), .A(n3200), .ZN(n4785) );
  AOI211_X1 U4074 ( .C1(n4821), .C2(n4783), .A(n4787), .B(n4785), .ZN(n4816)
         );
  NAND2_X1 U4075 ( .A1(n4825), .A2(REG1_REG_0__SCAN_IN), .ZN(n3201) );
  OAI21_X1 U4076 ( .B1(n4816), .B2(n4825), .A(n3201), .ZN(U3518) );
  XNOR2_X1 U4077 ( .A(n4722), .B(n3202), .ZN(n3203) );
  XNOR2_X1 U4078 ( .A(n3204), .B(n3203), .ZN(n3213) );
  NAND2_X1 U4079 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3440) );
  INV_X1 U4080 ( .A(n3440), .ZN(n3207) );
  NOR2_X1 U4081 ( .A1(n4775), .A2(n3205), .ZN(n3206) );
  AOI211_X1 U4082 ( .C1(n4765), .C2(ADDR_REG_7__SCAN_IN), .A(n3207), .B(n3206), 
        .ZN(n3212) );
  OAI211_X1 U4083 ( .C1(n3210), .C2(n3209), .A(n3208), .B(n4096), .ZN(n3211)
         );
  OAI211_X1 U4084 ( .C1(n3213), .C2(n4113), .A(n3212), .B(n3211), .ZN(U3247)
         );
  INV_X1 U4085 ( .A(n3214), .ZN(n3217) );
  NAND3_X1 U4086 ( .A1(n3217), .A2(n3216), .A3(n3215), .ZN(n3267) );
  NAND2_X1 U4087 ( .A1(n3267), .A2(REG3_REG_0__SCAN_IN), .ZN(n3221) );
  INV_X1 U4088 ( .A(n3218), .ZN(n3219) );
  AOI22_X1 U4089 ( .A1(n3876), .A2(n3219), .B1(n3890), .B2(n2459), .ZN(n3220)
         );
  OAI211_X1 U4090 ( .C1(n3900), .C2(n3222), .A(n3221), .B(n3220), .ZN(U3229)
         );
  INV_X1 U4091 ( .A(n3267), .ZN(n3230) );
  INV_X1 U4092 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3229) );
  INV_X1 U4093 ( .A(n3900), .ZN(n3669) );
  OAI22_X1 U4094 ( .A1(n3324), .A2(n3865), .B1(n3898), .B2(n3323), .ZN(n3223)
         );
  AOI21_X1 U4095 ( .B1(n2832), .B2(n3669), .A(n3223), .ZN(n3228) );
  OAI211_X1 U4096 ( .C1(n3226), .C2(n3225), .A(n3224), .B(n3876), .ZN(n3227)
         );
  OAI211_X1 U4097 ( .C1(n3230), .C2(n3229), .A(n3228), .B(n3227), .ZN(U3219)
         );
  OR2_X1 U4098 ( .A1(n3231), .A2(n3232), .ZN(n3233) );
  AND2_X1 U4099 ( .A1(n3287), .A2(n3233), .ZN(n3325) );
  INV_X1 U4100 ( .A(n3231), .ZN(n3989) );
  OAI21_X1 U4101 ( .B1(n3989), .B2(n3911), .A(n3234), .ZN(n3235) );
  AOI22_X1 U4102 ( .A1(n3507), .A2(n3325), .B1(n3235), .B2(n4465), .ZN(n3327)
         );
  AOI22_X1 U4103 ( .A1(n2840), .A2(n4475), .B1(n4458), .B2(n2832), .ZN(n3238)
         );
  NAND2_X1 U4104 ( .A1(n2823), .A2(n4486), .ZN(n3237) );
  NAND2_X1 U4105 ( .A1(n3325), .A2(n4821), .ZN(n3236) );
  NAND4_X1 U4106 ( .A1(n3327), .A2(n3238), .A3(n3237), .A4(n3236), .ZN(n3247)
         );
  AND2_X1 U4107 ( .A1(n2832), .A2(n3240), .ZN(n3241) );
  NOR2_X1 U4108 ( .A1(n3239), .A2(n3241), .ZN(n3333) );
  INV_X1 U4109 ( .A(n3333), .ZN(n3245) );
  OAI22_X1 U4110 ( .A1(n4484), .A2(n3245), .B1(n4828), .B2(n2241), .ZN(n3242)
         );
  AOI21_X1 U4111 ( .B1(n3247), .B2(n4828), .A(n3242), .ZN(n3243) );
  INV_X1 U4112 ( .A(n3243), .ZN(U3519) );
  INV_X1 U4113 ( .A(REG0_REG_1__SCAN_IN), .ZN(n3244) );
  OAI22_X1 U4114 ( .A1(n4706), .A2(n3245), .B1(n4824), .B2(n3244), .ZN(n3246)
         );
  AOI21_X1 U4115 ( .B1(n3247), .B2(n4824), .A(n3246), .ZN(n3248) );
  INV_X1 U4116 ( .A(n3248), .ZN(U3469) );
  XOR2_X1 U4117 ( .A(n3249), .B(REG2_REG_4__SCAN_IN), .Z(n3258) );
  NAND2_X1 U4118 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3428) );
  INV_X1 U4119 ( .A(n3428), .ZN(n3250) );
  AOI21_X1 U4120 ( .B1(n4765), .B2(ADDR_REG_4__SCAN_IN), .A(n3250), .ZN(n3251)
         );
  OAI211_X1 U4121 ( .C1(n4775), .C2(n3253), .A(n3252), .B(n3251), .ZN(n3257)
         );
  AOI211_X1 U4122 ( .C1(n4826), .C2(n3255), .A(n4113), .B(n3254), .ZN(n3256)
         );
  AOI211_X1 U4123 ( .C1(n4096), .C2(n3258), .A(n3257), .B(n3256), .ZN(n3259)
         );
  INV_X1 U4124 ( .A(n3259), .ZN(U3244) );
  INV_X1 U4125 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4537) );
  NAND2_X1 U4126 ( .A1(n4387), .A2(U4043), .ZN(n3260) );
  OAI21_X1 U4127 ( .B1(n4077), .B2(n4537), .A(n3260), .ZN(U3575) );
  INV_X1 U4128 ( .A(n3261), .ZN(n3262) );
  AOI21_X1 U4129 ( .B1(n3264), .B2(n3263), .A(n3262), .ZN(n3269) );
  AOI22_X1 U4130 ( .A1(n3890), .A2(n3344), .B1(n3902), .B2(n2459), .ZN(n3265)
         );
  OAI21_X1 U4131 ( .B1(n3900), .B2(n3316), .A(n3265), .ZN(n3266) );
  AOI21_X1 U4132 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3267), .A(n3266), .ZN(n3268)
         );
  OAI21_X1 U4133 ( .B1(n3269), .B2(n3907), .A(n3268), .ZN(U3234) );
  XNOR2_X1 U4134 ( .A(n3270), .B(REG1_REG_8__SCAN_IN), .ZN(n3278) );
  XOR2_X1 U4135 ( .A(n3271), .B(REG2_REG_8__SCAN_IN), .Z(n3272) );
  NAND2_X1 U4136 ( .A1(n4096), .A2(n3272), .ZN(n3273) );
  NAND2_X1 U4137 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3498) );
  NAND2_X1 U4138 ( .A1(n3273), .A2(n3498), .ZN(n3276) );
  NOR2_X1 U4139 ( .A1(n4775), .A2(n3274), .ZN(n3275) );
  AOI211_X1 U4140 ( .C1(n4765), .C2(ADDR_REG_8__SCAN_IN), .A(n3276), .B(n3275), 
        .ZN(n3277) );
  OAI21_X1 U4141 ( .B1(n3278), .B2(n4113), .A(n3277), .ZN(U3248) );
  OAI22_X1 U4142 ( .A1(n3900), .A2(n3338), .B1(n3390), .B2(n3898), .ZN(n3279)
         );
  AOI211_X1 U4143 ( .C1(n3902), .C2(n2840), .A(n3280), .B(n3279), .ZN(n3285)
         );
  XNOR2_X1 U4144 ( .A(n3281), .B(n3282), .ZN(n3283) );
  NAND2_X1 U4145 ( .A1(n3283), .A2(n3876), .ZN(n3284) );
  OAI211_X1 U4146 ( .C1(REG3_REG_3__SCAN_IN), .C2(n3886), .A(n3285), .B(n3284), 
        .ZN(U3215) );
  AND2_X1 U4147 ( .A1(n3287), .A2(n3286), .ZN(n3290) );
  OAI21_X1 U4148 ( .B1(n3290), .B2(n3289), .A(n3288), .ZN(n3314) );
  INV_X1 U4149 ( .A(n4486), .ZN(n4390) );
  AOI22_X1 U4150 ( .A1(n3344), .A2(n4475), .B1(n3291), .B2(n4458), .ZN(n3292)
         );
  OAI21_X1 U4151 ( .B1(n3312), .B2(n4390), .A(n3292), .ZN(n3297) );
  OAI21_X1 U4152 ( .B1(n3988), .B2(n3294), .A(n3293), .ZN(n3295) );
  AOI22_X1 U4153 ( .A1(n3314), .A2(n3507), .B1(n3295), .B2(n4465), .ZN(n3320)
         );
  INV_X1 U4154 ( .A(n3320), .ZN(n3296) );
  AOI211_X1 U4155 ( .C1(n4821), .C2(n3314), .A(n3297), .B(n3296), .ZN(n3302)
         );
  XNOR2_X1 U4156 ( .A(n3239), .B(n3316), .ZN(n3311) );
  INV_X1 U4157 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3298) );
  OAI22_X1 U4158 ( .A1(n4706), .A2(n3311), .B1(n4824), .B2(n3298), .ZN(n3299)
         );
  INV_X1 U4159 ( .A(n3299), .ZN(n3300) );
  OAI21_X1 U4160 ( .B1(n3302), .B2(n4822), .A(n3300), .ZN(U3471) );
  INV_X1 U4161 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n4549) );
  NAND2_X1 U4162 ( .A1(n4137), .A2(U4043), .ZN(n3301) );
  OAI21_X1 U4163 ( .B1(n4077), .B2(n4549), .A(n3301), .ZN(U3576) );
  MUX2_X1 U4164 ( .A(n2245), .B(n3302), .S(n4828), .Z(n3303) );
  OAI21_X1 U4165 ( .B1(n3311), .B2(n4484), .A(n3303), .ZN(U3520) );
  NOR2_X1 U4166 ( .A1(n3305), .A2(n3304), .ZN(n3307) );
  NAND4_X1 U4167 ( .A1(n3309), .A2(n3308), .A3(n3307), .A4(n3306), .ZN(n3310)
         );
  INV_X1 U4168 ( .A(n3311), .ZN(n3319) );
  OR2_X1 U4169 ( .A1(n4788), .A2(n4462), .ZN(n4337) );
  OAI22_X1 U4170 ( .A1(n3430), .A2(n4337), .B1(n4356), .B2(n3312), .ZN(n3318)
         );
  NAND2_X1 U4171 ( .A1(n3313), .A2(n4717), .ZN(n3372) );
  NOR2_X1 U4172 ( .A1(n4365), .A2(n3372), .ZN(n4784) );
  INV_X2 U4173 ( .A(n4792), .ZN(n4776) );
  AOI22_X1 U4174 ( .A1(n4784), .A2(n3314), .B1(REG3_REG_2__SCAN_IN), .B2(n4776), .ZN(n3315) );
  OAI21_X1 U4175 ( .B1(n3316), .B2(n4336), .A(n3315), .ZN(n3317) );
  AOI211_X1 U4176 ( .C1(n4779), .C2(n3319), .A(n3318), .B(n3317), .ZN(n3322)
         );
  MUX2_X1 U4177 ( .A(n2383), .B(n3320), .S(n4334), .Z(n3321) );
  NAND2_X1 U4178 ( .A1(n3322), .A2(n3321), .ZN(U3288) );
  OAI22_X1 U4179 ( .A1(n3324), .A2(n4356), .B1(n4337), .B2(n3323), .ZN(n3332)
         );
  AOI22_X1 U4180 ( .A1(n4784), .A2(n3325), .B1(REG3_REG_1__SCAN_IN), .B2(n4776), .ZN(n3329) );
  MUX2_X1 U4181 ( .A(n3327), .B(n3326), .S(n4788), .Z(n3328) );
  OAI211_X1 U4182 ( .C1(n4336), .C2(n3330), .A(n3329), .B(n3328), .ZN(n3331)
         );
  AOI211_X1 U4183 ( .C1(n4779), .C2(n3333), .A(n3332), .B(n3331), .ZN(n3334)
         );
  INV_X1 U4184 ( .A(n3334), .ZN(U3289) );
  OAI211_X1 U4185 ( .C1(n2071), .C2(n3336), .A(n4640), .B(n3369), .ZN(n4817)
         );
  NOR2_X1 U4186 ( .A1(n4817), .A2(n4717), .ZN(n3349) );
  NAND2_X1 U4187 ( .A1(n3288), .A2(n3337), .ZN(n3339) );
  INV_X1 U4188 ( .A(n3339), .ZN(n3353) );
  OAI21_X1 U4189 ( .B1(n3339), .B2(n3338), .A(n3430), .ZN(n3340) );
  OAI21_X1 U4190 ( .B1(n3353), .B2(n3361), .A(n3340), .ZN(n3342) );
  INV_X1 U4191 ( .A(n3341), .ZN(n3992) );
  XNOR2_X1 U4192 ( .A(n3342), .B(n3992), .ZN(n3350) );
  XNOR2_X1 U4193 ( .A(n3343), .B(n3992), .ZN(n3347) );
  AOI22_X1 U4194 ( .A1(n3344), .A2(n4486), .B1(n2475), .B2(n4458), .ZN(n3345)
         );
  OAI21_X1 U4195 ( .B1(n3402), .B2(n4462), .A(n3345), .ZN(n3346) );
  AOI21_X1 U4196 ( .B1(n3347), .B2(n4465), .A(n3346), .ZN(n3348) );
  OAI21_X1 U4197 ( .B1(n3350), .B2(n3561), .A(n3348), .ZN(n4818) );
  AOI211_X1 U4198 ( .C1(n4776), .C2(n3436), .A(n3349), .B(n4818), .ZN(n3352)
         );
  INV_X1 U4199 ( .A(n3350), .ZN(n4820) );
  AOI22_X1 U4200 ( .A1(n4820), .A2(n4784), .B1(REG2_REG_4__SCAN_IN), .B2(n4365), .ZN(n3351) );
  OAI21_X1 U4201 ( .B1(n3352), .B2(n4365), .A(n3351), .ZN(U3286) );
  XNOR2_X1 U4202 ( .A(n3353), .B(n3990), .ZN(n4777) );
  OAI21_X1 U4203 ( .B1(n3990), .B2(n3355), .A(n3354), .ZN(n3356) );
  NAND2_X1 U4204 ( .A1(n3356), .A2(n4465), .ZN(n3358) );
  AOI22_X1 U4205 ( .A1(n2840), .A2(n4486), .B1(n4458), .B2(n3361), .ZN(n3357)
         );
  OAI211_X1 U4206 ( .C1(n3390), .C2(n4462), .A(n3358), .B(n3357), .ZN(n3359)
         );
  AOI21_X1 U4207 ( .B1(n3507), .B2(n4777), .A(n3359), .ZN(n4782) );
  INV_X1 U4208 ( .A(n4782), .ZN(n3360) );
  AOI21_X1 U4209 ( .B1(n4821), .B2(n4777), .A(n3360), .ZN(n3366) );
  INV_X1 U4210 ( .A(n4484), .ZN(n4366) );
  NAND2_X1 U4211 ( .A1(n3362), .A2(n3361), .ZN(n3363) );
  AND2_X1 U4212 ( .A1(n3335), .A2(n3363), .ZN(n4778) );
  AOI22_X1 U4213 ( .A1(n4366), .A2(n4778), .B1(REG1_REG_3__SCAN_IN), .B2(n4825), .ZN(n3364) );
  OAI21_X1 U4214 ( .B1(n3366), .B2(n4825), .A(n3364), .ZN(U3521) );
  INV_X1 U4215 ( .A(n4706), .ZN(n4650) );
  AOI22_X1 U4216 ( .A1(n4650), .A2(n4778), .B1(REG0_REG_3__SCAN_IN), .B2(n4822), .ZN(n3365) );
  OAI21_X1 U4217 ( .B1(n3366), .B2(n4822), .A(n3365), .ZN(U3473) );
  AND2_X1 U4218 ( .A1(n2047), .A2(n3937), .ZN(n3987) );
  XNOR2_X1 U4219 ( .A(n3367), .B(n3987), .ZN(n3368) );
  NOR2_X1 U4220 ( .A1(n3368), .A2(n4327), .ZN(n3467) );
  INV_X1 U4221 ( .A(n3467), .ZN(n3381) );
  AND2_X1 U4222 ( .A1(n3369), .A2(n3464), .ZN(n3370) );
  NOR2_X1 U4223 ( .A1(n3408), .A2(n3370), .ZN(n3471) );
  INV_X1 U4224 ( .A(n3471), .ZN(n3371) );
  NOR2_X1 U4225 ( .A1(n4342), .A2(n3371), .ZN(n3379) );
  OAI22_X1 U4226 ( .A1(n3466), .A2(n4337), .B1(n4336), .B2(n2070), .ZN(n3378)
         );
  AND2_X1 U4227 ( .A1(n3561), .A2(n3372), .ZN(n3373) );
  XNOR2_X1 U4228 ( .A(n3374), .B(n3987), .ZN(n3469) );
  AND2_X1 U4229 ( .A1(n4344), .A2(n3469), .ZN(n3377) );
  AOI22_X1 U4230 ( .A1(n4365), .A2(REG2_REG_5__SCAN_IN), .B1(n3382), .B2(n4776), .ZN(n3375) );
  OAI21_X1 U4231 ( .B1(n4356), .B2(n3390), .A(n3375), .ZN(n3376) );
  NOR4_X1 U4232 ( .A1(n3379), .A2(n3378), .A3(n3377), .A4(n3376), .ZN(n3380)
         );
  OAI21_X1 U4233 ( .B1(n3381), .B2(n4365), .A(n3380), .ZN(U3285) );
  INV_X1 U4234 ( .A(n3382), .ZN(n3395) );
  OR2_X1 U4235 ( .A1(n3383), .A2(n3433), .ZN(n3431) );
  NAND2_X1 U4236 ( .A1(n3431), .A2(n3384), .ZN(n3389) );
  AND2_X1 U4237 ( .A1(n3386), .A2(n3385), .ZN(n3387) );
  OAI211_X1 U4238 ( .C1(n3389), .C2(n3388), .A(n3387), .B(n3876), .ZN(n3394)
         );
  OAI22_X1 U4239 ( .A1(n3900), .A2(n2070), .B1(n3466), .B2(n3898), .ZN(n3391)
         );
  AOI211_X1 U4240 ( .C1(n3902), .C2(n2861), .A(n3392), .B(n3391), .ZN(n3393)
         );
  OAI211_X1 U4241 ( .C1(n3886), .C2(n3395), .A(n3394), .B(n3393), .ZN(U3224)
         );
  XOR2_X1 U4242 ( .A(n3397), .B(n3396), .Z(n3398) );
  XNOR2_X1 U4243 ( .A(n3399), .B(n3398), .ZN(n3405) );
  AOI22_X1 U4244 ( .A1(n3669), .A2(n3411), .B1(n3890), .B2(n4075), .ZN(n3401)
         );
  OAI211_X1 U4245 ( .C1(n3402), .C2(n3865), .A(n3401), .B(n3400), .ZN(n3403)
         );
  AOI21_X1 U4246 ( .B1(n3412), .B2(n3904), .A(n3403), .ZN(n3404) );
  OAI21_X1 U4247 ( .B1(n3405), .B2(n3907), .A(n3404), .ZN(U3236) );
  NAND2_X1 U4248 ( .A1(n3923), .A2(n3936), .ZN(n3997) );
  XNOR2_X1 U4249 ( .A(n3406), .B(n3997), .ZN(n3421) );
  XOR2_X1 U4250 ( .A(n3407), .B(n3997), .Z(n3423) );
  NOR2_X1 U4251 ( .A1(n4365), .A2(n4327), .ZN(n4280) );
  NAND2_X1 U4252 ( .A1(n3423), .A2(n4280), .ZN(n3417) );
  INV_X1 U4253 ( .A(n3408), .ZN(n3410) );
  AOI21_X1 U4254 ( .B1(n3411), .B2(n3410), .A(n2770), .ZN(n3425) );
  AOI22_X1 U4255 ( .A1(n4350), .A2(n4075), .B1(n4340), .B2(n2016), .ZN(n3414)
         );
  AOI22_X1 U4256 ( .A1(n4365), .A2(REG2_REG_6__SCAN_IN), .B1(n3412), .B2(n4776), .ZN(n3413) );
  OAI211_X1 U4257 ( .C1(n3418), .C2(n4336), .A(n3414), .B(n3413), .ZN(n3415)
         );
  AOI21_X1 U4258 ( .B1(n4779), .B2(n3425), .A(n3415), .ZN(n3416) );
  OAI211_X1 U4259 ( .C1(n4361), .C2(n3421), .A(n3417), .B(n3416), .ZN(U3284)
         );
  INV_X1 U4260 ( .A(n4482), .ZN(n4649) );
  OAI22_X1 U4261 ( .A1(n3510), .A2(n4462), .B1(n3418), .B2(n4477), .ZN(n3419)
         );
  AOI21_X1 U4262 ( .B1(n4486), .B2(n2016), .A(n3419), .ZN(n3420) );
  OAI21_X1 U4263 ( .B1(n3421), .B2(n4649), .A(n3420), .ZN(n3422) );
  AOI21_X1 U4264 ( .B1(n3423), .B2(n4465), .A(n3422), .ZN(n3427) );
  AOI22_X1 U4265 ( .A1(n3425), .A2(n4650), .B1(REG0_REG_6__SCAN_IN), .B2(n4822), .ZN(n3424) );
  OAI21_X1 U4266 ( .B1(n3427), .B2(n4822), .A(n3424), .ZN(U3479) );
  AOI22_X1 U4267 ( .A1(n3425), .A2(n4366), .B1(REG1_REG_6__SCAN_IN), .B2(n4825), .ZN(n3426) );
  OAI21_X1 U4268 ( .B1(n3427), .B2(n4825), .A(n3426), .ZN(U3524) );
  AOI22_X1 U4269 ( .A1(n3669), .A2(n2475), .B1(n3890), .B2(n2016), .ZN(n3429)
         );
  OAI211_X1 U4270 ( .C1(n3430), .C2(n3865), .A(n3429), .B(n3428), .ZN(n3435)
         );
  INV_X1 U4271 ( .A(n3431), .ZN(n3432) );
  AOI211_X1 U4272 ( .C1(n3433), .C2(n3383), .A(n3907), .B(n3432), .ZN(n3434)
         );
  AOI211_X1 U4273 ( .C1(n3436), .C2(n3904), .A(n3435), .B(n3434), .ZN(n3437)
         );
  INV_X1 U4274 ( .A(n3437), .ZN(U3227) );
  XNOR2_X1 U4275 ( .A(n3438), .B(n3439), .ZN(n3444) );
  AOI22_X1 U4276 ( .A1(n3669), .A2(n3456), .B1(n3902), .B2(n3447), .ZN(n3441)
         );
  OAI211_X1 U4277 ( .C1(n3541), .C2(n3898), .A(n3441), .B(n3440), .ZN(n3442)
         );
  AOI21_X1 U4278 ( .B1(n3458), .B2(n3904), .A(n3442), .ZN(n3443) );
  OAI21_X1 U4279 ( .B1(n3444), .B2(n3907), .A(n3443), .ZN(U3210) );
  XNOR2_X1 U4280 ( .A(n3445), .B(n3924), .ZN(n3446) );
  NAND2_X1 U4281 ( .A1(n3446), .A2(n4465), .ZN(n3449) );
  AOI22_X1 U4282 ( .A1(n3447), .A2(n4486), .B1(n4458), .B2(n3456), .ZN(n3448)
         );
  OAI211_X1 U4283 ( .C1(n3541), .C2(n4462), .A(n3449), .B(n3448), .ZN(n3450)
         );
  INV_X1 U4284 ( .A(n3450), .ZN(n4647) );
  NAND2_X1 U4285 ( .A1(n3452), .A2(n3451), .ZN(n3453) );
  NAND2_X1 U4286 ( .A1(n3453), .A2(n3924), .ZN(n3454) );
  NAND2_X1 U4287 ( .A1(n3505), .A2(n3454), .ZN(n4648) );
  INV_X1 U4288 ( .A(n4648), .ZN(n3462) );
  INV_X1 U4289 ( .A(n4323), .ZN(n3460) );
  AOI21_X1 U4290 ( .B1(n3409), .B2(n3456), .A(n3455), .ZN(n3457) );
  NAND2_X1 U4291 ( .A1(n3457), .A2(n3517), .ZN(n4646) );
  AOI22_X1 U4292 ( .A1(n4365), .A2(REG2_REG_7__SCAN_IN), .B1(n3458), .B2(n4776), .ZN(n3459) );
  OAI21_X1 U4293 ( .B1(n3460), .B2(n4646), .A(n3459), .ZN(n3461) );
  AOI21_X1 U4294 ( .B1(n3462), .B2(n4344), .A(n3461), .ZN(n3463) );
  OAI21_X1 U4295 ( .B1(n4647), .B2(n4365), .A(n3463), .ZN(U3283) );
  AOI22_X1 U4296 ( .A1(n2861), .A2(n4486), .B1(n4458), .B2(n3464), .ZN(n3465)
         );
  OAI21_X1 U4297 ( .B1(n3466), .B2(n4462), .A(n3465), .ZN(n3468) );
  AOI211_X1 U4298 ( .C1(n3469), .C2(n4482), .A(n3468), .B(n3467), .ZN(n3473)
         );
  AOI22_X1 U4299 ( .A1(n4366), .A2(n3471), .B1(REG1_REG_5__SCAN_IN), .B2(n4825), .ZN(n3470) );
  OAI21_X1 U4300 ( .B1(n3473), .B2(n4825), .A(n3470), .ZN(U3523) );
  AOI22_X1 U4301 ( .A1(n4650), .A2(n3471), .B1(REG0_REG_5__SCAN_IN), .B2(n4822), .ZN(n3472) );
  OAI21_X1 U4302 ( .B1(n3473), .B2(n4822), .A(n3472), .ZN(U3477) );
  XNOR2_X1 U4303 ( .A(n3474), .B(REG1_REG_10__SCAN_IN), .ZN(n3481) );
  XOR2_X1 U4304 ( .A(n3475), .B(REG2_REG_10__SCAN_IN), .Z(n3479) );
  NAND2_X1 U4305 ( .A1(U3149), .A2(REG3_REG_10__SCAN_IN), .ZN(n3670) );
  NAND2_X1 U4306 ( .A1(n4765), .A2(ADDR_REG_10__SCAN_IN), .ZN(n3476) );
  OAI211_X1 U4307 ( .C1(n4775), .C2(n3477), .A(n3670), .B(n3476), .ZN(n3478)
         );
  AOI21_X1 U4308 ( .B1(n3479), .B2(n4096), .A(n3478), .ZN(n3480) );
  OAI21_X1 U4309 ( .B1(n3481), .B2(n4113), .A(n3480), .ZN(U3250) );
  XNOR2_X1 U4310 ( .A(n3482), .B(n3483), .ZN(n3492) );
  INV_X1 U4311 ( .A(n4765), .ZN(n4094) );
  NAND2_X1 U4312 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n3550) );
  OAI21_X1 U4313 ( .B1(n4094), .B2(n4585), .A(n3550), .ZN(n3490) );
  INV_X1 U4314 ( .A(n3484), .ZN(n3488) );
  INV_X1 U4315 ( .A(n3485), .ZN(n3486) );
  AOI211_X1 U4316 ( .C1(n3488), .C2(n3487), .A(n4113), .B(n3486), .ZN(n3489)
         );
  AOI211_X1 U4317 ( .C1(n4110), .C2(n4720), .A(n3490), .B(n3489), .ZN(n3491)
         );
  OAI21_X1 U4318 ( .B1(n3492), .B2(n4762), .A(n3491), .ZN(U3249) );
  INV_X1 U4319 ( .A(n3494), .ZN(n3496) );
  NOR2_X1 U4320 ( .A1(n3496), .A2(n3495), .ZN(n3497) );
  XNOR2_X1 U4321 ( .A(n3493), .B(n3497), .ZN(n3502) );
  AOI22_X1 U4322 ( .A1(n3669), .A2(n3516), .B1(n3902), .B2(n4075), .ZN(n3499)
         );
  OAI211_X1 U4323 ( .C1(n3672), .C2(n3898), .A(n3499), .B(n3498), .ZN(n3500)
         );
  AOI21_X1 U4324 ( .B1(n3514), .B2(n3904), .A(n3500), .ZN(n3501) );
  OAI21_X1 U4325 ( .B1(n3502), .B2(n3907), .A(n3501), .ZN(U3218) );
  NAND2_X1 U4326 ( .A1(n3503), .A2(n3927), .ZN(n3534) );
  AND2_X1 U4327 ( .A1(n3928), .A2(n3926), .ZN(n3986) );
  XOR2_X1 U4328 ( .A(n3534), .B(n3986), .Z(n3512) );
  NAND2_X1 U4329 ( .A1(n3505), .A2(n3504), .ZN(n3506) );
  XNOR2_X1 U4330 ( .A(n3506), .B(n3986), .ZN(n3513) );
  NAND2_X1 U4331 ( .A1(n3513), .A2(n3507), .ZN(n3509) );
  AOI22_X1 U4332 ( .A1(n3525), .A2(n4475), .B1(n3516), .B2(n4458), .ZN(n3508)
         );
  OAI211_X1 U4333 ( .C1(n3510), .C2(n4390), .A(n3509), .B(n3508), .ZN(n3511)
         );
  AOI21_X1 U4334 ( .B1(n3512), .B2(n4465), .A(n3511), .ZN(n4643) );
  INV_X1 U4335 ( .A(n3513), .ZN(n4645) );
  INV_X1 U4336 ( .A(n4784), .ZN(n3568) );
  AOI22_X1 U4337 ( .A1(n4365), .A2(REG2_REG_8__SCAN_IN), .B1(n3514), .B2(n4776), .ZN(n3519) );
  INV_X1 U4338 ( .A(n3515), .ZN(n4641) );
  NAND2_X1 U4339 ( .A1(n3517), .A2(n3516), .ZN(n4639) );
  NAND3_X1 U4340 ( .A1(n4779), .A2(n4641), .A3(n4639), .ZN(n3518) );
  OAI211_X1 U4341 ( .C1(n4645), .C2(n3568), .A(n3519), .B(n3518), .ZN(n3520)
         );
  INV_X1 U4342 ( .A(n3520), .ZN(n3521) );
  OAI21_X1 U4343 ( .B1(n4643), .B2(n4365), .A(n3521), .ZN(U3282) );
  NAND2_X1 U4344 ( .A1(n3943), .A2(n3944), .ZN(n4010) );
  XOR2_X1 U4345 ( .A(n3522), .B(n4010), .Z(n3575) );
  XOR2_X1 U4346 ( .A(n3523), .B(n4010), .Z(n3577) );
  NAND2_X1 U4347 ( .A1(n3577), .A2(n4280), .ZN(n3531) );
  OAI21_X1 U4348 ( .B1(n3524), .B2(n3572), .A(n3565), .ZN(n3582) );
  INV_X1 U4349 ( .A(n3582), .ZN(n3529) );
  AOI22_X1 U4350 ( .A1(n4340), .A2(n3525), .B1(n4350), .B2(n4473), .ZN(n3527)
         );
  AOI22_X1 U4351 ( .A1(n4365), .A2(REG2_REG_10__SCAN_IN), .B1(n3679), .B2(
        n4776), .ZN(n3526) );
  OAI211_X1 U4352 ( .C1(n3572), .C2(n4336), .A(n3527), .B(n3526), .ZN(n3528)
         );
  AOI21_X1 U4353 ( .B1(n3529), .B2(n4779), .A(n3528), .ZN(n3530) );
  OAI211_X1 U4354 ( .C1(n4361), .C2(n3575), .A(n3531), .B(n3530), .ZN(U3280)
         );
  NAND2_X1 U4355 ( .A1(n3533), .A2(n3532), .ZN(n3996) );
  NAND2_X1 U4356 ( .A1(n3534), .A2(n3928), .ZN(n3535) );
  NAND2_X1 U4357 ( .A1(n3535), .A2(n3926), .ZN(n3536) );
  XOR2_X1 U4358 ( .A(n3996), .B(n3536), .Z(n3537) );
  NOR2_X1 U4359 ( .A1(n3537), .A2(n4327), .ZN(n3608) );
  INV_X1 U4360 ( .A(n3608), .ZN(n3547) );
  XNOR2_X1 U4361 ( .A(n3538), .B(n3996), .ZN(n3610) );
  INV_X1 U4362 ( .A(n4336), .ZN(n4351) );
  AOI22_X1 U4363 ( .A1(n4351), .A2(n3606), .B1(n4350), .B2(n4485), .ZN(n3540)
         );
  AOI22_X1 U4364 ( .A1(n4788), .A2(REG2_REG_9__SCAN_IN), .B1(n3553), .B2(n4776), .ZN(n3539) );
  OAI211_X1 U4365 ( .C1(n3541), .C2(n4356), .A(n3540), .B(n3539), .ZN(n3545)
         );
  INV_X1 U4366 ( .A(n3524), .ZN(n3542) );
  OAI21_X1 U4367 ( .B1(n3515), .B2(n3543), .A(n3542), .ZN(n3615) );
  NOR2_X1 U4368 ( .A1(n3615), .A2(n4342), .ZN(n3544) );
  AOI211_X1 U4369 ( .C1(n3610), .C2(n4344), .A(n3545), .B(n3544), .ZN(n3546)
         );
  OAI21_X1 U4370 ( .B1(n3547), .B2(n4788), .A(n3546), .ZN(U3281) );
  XOR2_X1 U4371 ( .A(n3548), .B(n3549), .Z(n3555) );
  AOI22_X1 U4372 ( .A1(n3669), .A2(n3606), .B1(n3902), .B2(n4074), .ZN(n3551)
         );
  OAI211_X1 U4373 ( .C1(n3620), .C2(n3898), .A(n3551), .B(n3550), .ZN(n3552)
         );
  AOI21_X1 U4374 ( .B1(n3553), .B2(n3904), .A(n3552), .ZN(n3554) );
  OAI21_X1 U4375 ( .B1(n3555), .B2(n3907), .A(n3554), .ZN(U3228) );
  XNOR2_X1 U4376 ( .A(n3556), .B(n3991), .ZN(n3563) );
  INV_X1 U4377 ( .A(n3557), .ZN(n3558) );
  AOI21_X1 U4378 ( .B1(n3991), .B2(n3559), .A(n3558), .ZN(n4490) );
  AOI22_X1 U4379 ( .A1(n4073), .A2(n4475), .B1(n4458), .B2(n3566), .ZN(n3560)
         );
  OAI21_X1 U4380 ( .B1(n4490), .B2(n3561), .A(n3560), .ZN(n3562) );
  AOI21_X1 U4381 ( .B1(n3563), .B2(n4465), .A(n3562), .ZN(n4489) );
  INV_X1 U4382 ( .A(n3564), .ZN(n3589) );
  AOI21_X1 U4383 ( .B1(n3566), .B2(n3565), .A(n3589), .ZN(n4487) );
  AOI22_X1 U4384 ( .A1(n4365), .A2(REG2_REG_11__SCAN_IN), .B1(n3624), .B2(
        n4776), .ZN(n3567) );
  OAI21_X1 U4385 ( .B1(n4356), .B2(n3620), .A(n3567), .ZN(n3570) );
  NOR2_X1 U4386 ( .A1(n4490), .A2(n3568), .ZN(n3569) );
  AOI211_X1 U4387 ( .C1(n4487), .C2(n4779), .A(n3570), .B(n3569), .ZN(n3571)
         );
  OAI21_X1 U4388 ( .B1(n4489), .B2(n4365), .A(n3571), .ZN(U3279) );
  OAI22_X1 U4389 ( .A1(n3672), .A2(n4390), .B1(n3572), .B2(n4477), .ZN(n3573)
         );
  AOI21_X1 U4390 ( .B1(n4475), .B2(n4473), .A(n3573), .ZN(n3574) );
  OAI21_X1 U4391 ( .B1(n3575), .B2(n4649), .A(n3574), .ZN(n3576) );
  AOI21_X1 U4392 ( .B1(n3577), .B2(n4465), .A(n3576), .ZN(n3580) );
  INV_X1 U4393 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3578) );
  MUX2_X1 U4394 ( .A(n3580), .B(n3578), .S(n4825), .Z(n3579) );
  OAI21_X1 U4395 ( .B1(n4484), .B2(n3582), .A(n3579), .ZN(U3528) );
  INV_X1 U4396 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4567) );
  MUX2_X1 U4397 ( .A(n3580), .B(n4567), .S(n4822), .Z(n3581) );
  OAI21_X1 U4398 ( .B1(n3582), .B2(n4706), .A(n3581), .ZN(U3487) );
  INV_X1 U4399 ( .A(n3583), .ZN(n3584) );
  AOI21_X1 U4400 ( .B1(n3556), .B2(n3585), .A(n3584), .ZN(n3631) );
  AND2_X1 U4401 ( .A1(n3630), .A2(n3628), .ZN(n4000) );
  XNOR2_X1 U4402 ( .A(n3631), .B(n4000), .ZN(n3586) );
  NOR2_X1 U4403 ( .A1(n3586), .A2(n4327), .ZN(n4479) );
  INV_X1 U4404 ( .A(n4479), .ZN(n3596) );
  XOR2_X1 U4405 ( .A(n4000), .B(n3587), .Z(n4481) );
  INV_X1 U4406 ( .A(n3638), .ZN(n3588) );
  OAI21_X1 U4407 ( .B1(n3589), .B2(n4478), .A(n3588), .ZN(n4707) );
  NOR2_X1 U4408 ( .A1(n4707), .A2(n4342), .ZN(n3594) );
  AOI22_X1 U4409 ( .A1(n3590), .A2(n4351), .B1(n4350), .B2(n4474), .ZN(n3592)
         );
  AOI22_X1 U4410 ( .A1(n4365), .A2(REG2_REG_12__SCAN_IN), .B1(n3803), .B2(
        n4776), .ZN(n3591) );
  OAI211_X1 U4411 ( .C1(n3799), .C2(n4356), .A(n3592), .B(n3591), .ZN(n3593)
         );
  AOI211_X1 U4412 ( .C1(n4481), .C2(n4344), .A(n3594), .B(n3593), .ZN(n3595)
         );
  OAI21_X1 U4413 ( .B1(n3596), .B2(n4365), .A(n3595), .ZN(U3278) );
  XNOR2_X1 U4414 ( .A(n3597), .B(REG1_REG_12__SCAN_IN), .ZN(n3605) );
  XOR2_X1 U4415 ( .A(REG2_REG_12__SCAN_IN), .B(n3598), .Z(n3599) );
  NAND2_X1 U4416 ( .A1(n4096), .A2(n3599), .ZN(n3600) );
  NAND2_X1 U4417 ( .A1(U3149), .A2(REG3_REG_12__SCAN_IN), .ZN(n3798) );
  NAND2_X1 U4418 ( .A1(n3600), .A2(n3798), .ZN(n3603) );
  NOR2_X1 U4419 ( .A1(n4775), .A2(n3601), .ZN(n3602) );
  AOI211_X1 U4420 ( .C1(n4765), .C2(ADDR_REG_12__SCAN_IN), .A(n3603), .B(n3602), .ZN(n3604) );
  OAI21_X1 U4421 ( .B1(n3605), .B2(n4113), .A(n3604), .ZN(U3252) );
  AOI22_X1 U4422 ( .A1(n4074), .A2(n4486), .B1(n4458), .B2(n3606), .ZN(n3607)
         );
  OAI21_X1 U4423 ( .B1(n3620), .B2(n4462), .A(n3607), .ZN(n3609) );
  AOI211_X1 U4424 ( .C1(n3610), .C2(n4482), .A(n3609), .B(n3608), .ZN(n3612)
         );
  MUX2_X1 U4425 ( .A(n2277), .B(n3612), .S(n4828), .Z(n3611) );
  OAI21_X1 U4426 ( .B1(n4484), .B2(n3615), .A(n3611), .ZN(U3527) );
  INV_X1 U4427 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3613) );
  MUX2_X1 U4428 ( .A(n3613), .B(n3612), .S(n4824), .Z(n3614) );
  OAI21_X1 U4429 ( .B1(n3615), .B2(n4706), .A(n3614), .ZN(U3485) );
  XOR2_X1 U4430 ( .A(n3617), .B(n3616), .Z(n3618) );
  XNOR2_X1 U4431 ( .A(n3619), .B(n3618), .ZN(n3626) );
  NAND2_X1 U4432 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4092) );
  OAI21_X1 U4433 ( .B1(n3865), .B2(n3620), .A(n4092), .ZN(n3623) );
  OAI22_X1 U4434 ( .A1(n3900), .A2(n3621), .B1(n3853), .B2(n3898), .ZN(n3622)
         );
  AOI211_X1 U4435 ( .C1(n3904), .C2(n3624), .A(n3623), .B(n3622), .ZN(n3625)
         );
  OAI21_X1 U4436 ( .B1(n3626), .B2(n3907), .A(n3625), .ZN(U3233) );
  XNOR2_X1 U4437 ( .A(n4474), .B(n3627), .ZN(n4015) );
  INV_X1 U4438 ( .A(n3628), .ZN(n3629) );
  AOI21_X1 U4439 ( .B1(n3631), .B2(n3630), .A(n3629), .ZN(n3632) );
  XOR2_X1 U4440 ( .A(n4015), .B(n3632), .Z(n3635) );
  OAI22_X1 U4441 ( .A1(n3853), .A2(n4390), .B1(n4477), .B2(n3855), .ZN(n3633)
         );
  AOI21_X1 U4442 ( .B1(n4475), .B2(n4450), .A(n3633), .ZN(n3634) );
  OAI21_X1 U4443 ( .B1(n3635), .B2(n4327), .A(n3634), .ZN(n4469) );
  INV_X1 U4444 ( .A(n4469), .ZN(n3642) );
  XOR2_X1 U4445 ( .A(n4015), .B(n3636), .Z(n4470) );
  INV_X1 U4446 ( .A(n3646), .ZN(n3637) );
  OAI21_X1 U4447 ( .B1(n3638), .B2(n3855), .A(n3637), .ZN(n4702) );
  AOI22_X1 U4448 ( .A1(n4365), .A2(REG2_REG_13__SCAN_IN), .B1(n3858), .B2(
        n4776), .ZN(n3639) );
  OAI21_X1 U4449 ( .B1(n4702), .B2(n4342), .A(n3639), .ZN(n3640) );
  AOI21_X1 U4450 ( .B1(n4470), .B2(n4344), .A(n3640), .ZN(n3641) );
  OAI21_X1 U4451 ( .B1(n3642), .B2(n4365), .A(n3641), .ZN(U3277) );
  XNOR2_X1 U4452 ( .A(n3643), .B(n3993), .ZN(n4466) );
  INV_X1 U4453 ( .A(n4466), .ZN(n3653) );
  INV_X1 U4454 ( .A(n4280), .ZN(n3652) );
  OAI21_X1 U4455 ( .B1(n2054), .B2(n3645), .A(n3644), .ZN(n4457) );
  OAI21_X1 U4456 ( .B1(n3646), .B2(n3756), .A(n3685), .ZN(n4699) );
  NOR2_X1 U4457 ( .A1(n4699), .A2(n4342), .ZN(n3650) );
  AOI22_X1 U4458 ( .A1(n4350), .A2(n4440), .B1(n4340), .B2(n4474), .ZN(n3648)
         );
  AOI22_X1 U4459 ( .A1(n4788), .A2(REG2_REG_14__SCAN_IN), .B1(n3759), .B2(
        n4776), .ZN(n3647) );
  OAI211_X1 U4460 ( .C1(n3756), .C2(n4336), .A(n3648), .B(n3647), .ZN(n3649)
         );
  AOI211_X1 U4461 ( .C1(n4457), .C2(n4344), .A(n3650), .B(n3649), .ZN(n3651)
         );
  OAI21_X1 U4462 ( .B1(n3653), .B2(n3652), .A(n3651), .ZN(U3276) );
  XNOR2_X1 U4463 ( .A(n3659), .B(n3654), .ZN(n3655) );
  XNOR2_X1 U4464 ( .A(n3656), .B(n3655), .ZN(n3667) );
  NAND2_X1 U4465 ( .A1(n3659), .A2(n4471), .ZN(n3657) );
  OAI211_X1 U4466 ( .C1(n3659), .C2(n4471), .A(n3658), .B(n3657), .ZN(n3661)
         );
  NAND3_X1 U4467 ( .A1(n3661), .A2(n4770), .A3(n3660), .ZN(n3666) );
  NAND2_X1 U4468 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n3852) );
  INV_X1 U4469 ( .A(n3852), .ZN(n3664) );
  NOR2_X1 U4470 ( .A1(n4775), .A2(n3662), .ZN(n3663) );
  AOI211_X1 U4471 ( .C1(n4765), .C2(ADDR_REG_13__SCAN_IN), .A(n3664), .B(n3663), .ZN(n3665) );
  OAI211_X1 U4472 ( .C1(n3667), .C2(n4762), .A(n3666), .B(n3665), .ZN(U3253)
         );
  AOI22_X1 U4473 ( .A1(n3669), .A2(n3668), .B1(n3890), .B2(n4473), .ZN(n3671)
         );
  OAI211_X1 U4474 ( .C1(n3672), .C2(n3865), .A(n3671), .B(n3670), .ZN(n3678)
         );
  INV_X1 U4475 ( .A(n3673), .ZN(n3674) );
  AOI211_X1 U4476 ( .C1(n3676), .C2(n3675), .A(n3907), .B(n3674), .ZN(n3677)
         );
  AOI211_X1 U4477 ( .C1(n3679), .C2(n3904), .A(n3678), .B(n3677), .ZN(n3680)
         );
  INV_X1 U4478 ( .A(n3680), .ZN(U3214) );
  INV_X1 U4479 ( .A(n3681), .ZN(n3682) );
  AOI211_X1 U4480 ( .C1(n3683), .C2(n4006), .A(n4327), .B(n3682), .ZN(n4453)
         );
  INV_X1 U4481 ( .A(n4453), .ZN(n3693) );
  XNOR2_X1 U4482 ( .A(n3684), .B(n4006), .ZN(n4455) );
  INV_X1 U4483 ( .A(n3685), .ZN(n3687) );
  OAI21_X1 U4484 ( .B1(n3687), .B2(n3899), .A(n4349), .ZN(n4695) );
  NOR2_X1 U4485 ( .A1(n4695), .A2(n4342), .ZN(n3691) );
  AOI22_X1 U4486 ( .A1(n4351), .A2(n4449), .B1(n4350), .B2(n4432), .ZN(n3689)
         );
  AOI22_X1 U4487 ( .A1(n4788), .A2(REG2_REG_15__SCAN_IN), .B1(n3903), .B2(
        n4776), .ZN(n3688) );
  OAI211_X1 U4488 ( .C1(n3854), .C2(n4356), .A(n3689), .B(n3688), .ZN(n3690)
         );
  AOI211_X1 U4489 ( .C1(n4455), .C2(n4344), .A(n3691), .B(n3690), .ZN(n3692)
         );
  OAI21_X1 U4490 ( .B1(n3693), .B2(n4365), .A(n3692), .ZN(U3275) );
  AND2_X1 U4491 ( .A1(n3694), .A2(DATAI_30_), .ZN(n4119) );
  NAND2_X1 U4492 ( .A1(n3694), .A2(DATAI_31_), .ZN(n4057) );
  NAND2_X1 U4493 ( .A1(n3695), .A2(REG1_REG_31__SCAN_IN), .ZN(n3699) );
  NAND2_X1 U4494 ( .A1(n3696), .A2(REG2_REG_31__SCAN_IN), .ZN(n3698) );
  NAND2_X1 U4495 ( .A1(n2536), .A2(REG0_REG_31__SCAN_IN), .ZN(n3697) );
  NAND3_X1 U4496 ( .A1(n3699), .A2(n3698), .A3(n3697), .ZN(n4072) );
  NAND2_X1 U4497 ( .A1(n4072), .A2(n3700), .ZN(n4115) );
  OAI21_X1 U4498 ( .B1(n4057), .B2(n4477), .A(n4115), .ZN(n3705) );
  NAND2_X1 U4499 ( .A1(n4334), .A2(n3705), .ZN(n3702) );
  NAND2_X1 U4500 ( .A1(n4788), .A2(REG2_REG_31__SCAN_IN), .ZN(n3701) );
  OAI211_X1 U4501 ( .C1(n3708), .C2(n4342), .A(n3702), .B(n3701), .ZN(U3260)
         );
  NAND2_X1 U4502 ( .A1(n4828), .A2(n3705), .ZN(n3704) );
  NAND2_X1 U4503 ( .A1(n4825), .A2(REG1_REG_31__SCAN_IN), .ZN(n3703) );
  OAI211_X1 U4504 ( .C1(n3708), .C2(n4484), .A(n3704), .B(n3703), .ZN(U3549)
         );
  NAND2_X1 U4505 ( .A1(n4824), .A2(n3705), .ZN(n3707) );
  NAND2_X1 U4506 ( .A1(n4822), .A2(REG0_REG_31__SCAN_IN), .ZN(n3706) );
  OAI211_X1 U4507 ( .C1(n3708), .C2(n4706), .A(n3707), .B(n3706), .ZN(U3517)
         );
  OR2_X1 U4508 ( .A1(n3710), .A2(n3709), .ZN(n3711) );
  OR2_X1 U4509 ( .A1(n2045), .A2(n3711), .ZN(n3827) );
  AOI21_X1 U4510 ( .B1(n3762), .B2(n3713), .A(n3712), .ZN(n3829) );
  AOI21_X2 U4511 ( .B1(n3830), .B2(n3827), .A(n3829), .ZN(n3718) );
  OAI21_X1 U4512 ( .B1(n3716), .B2(n3715), .A(n3714), .ZN(n3717) );
  XNOR2_X1 U4513 ( .A(n3718), .B(n3717), .ZN(n3723) );
  OAI22_X1 U4514 ( .A1(n4210), .A2(n3865), .B1(STATE_REG_SCAN_IN), .B2(n3719), 
        .ZN(n3721) );
  INV_X1 U4515 ( .A(n4137), .ZN(n4381) );
  OAI22_X1 U4516 ( .A1(n4381), .A2(n3898), .B1(n3900), .B2(n4177), .ZN(n3720)
         );
  AOI211_X1 U4517 ( .C1(n4175), .C2(n3904), .A(n3721), .B(n3720), .ZN(n3722)
         );
  OAI21_X1 U4518 ( .B1(n3723), .B2(n3907), .A(n3722), .ZN(U3222) );
  XNOR2_X1 U4519 ( .A(n3725), .B(n3724), .ZN(n3731) );
  INV_X1 U4520 ( .A(n4136), .ZN(n3726) );
  NOR2_X1 U4521 ( .A1(n3726), .A2(n3886), .ZN(n3729) );
  AOI22_X1 U4522 ( .A1(n4137), .A2(n3902), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3727) );
  OAI21_X1 U4523 ( .B1(n3900), .B2(n4140), .A(n3727), .ZN(n3728) );
  AOI211_X1 U4524 ( .C1(n3890), .C2(n4143), .A(n3729), .B(n3728), .ZN(n3730)
         );
  OAI21_X1 U4525 ( .B1(n3731), .B2(n3907), .A(n3730), .ZN(U3211) );
  AOI21_X1 U4526 ( .B1(n3734), .B2(n3733), .A(n3732), .ZN(n3735) );
  XNOR2_X1 U4527 ( .A(n3735), .B(n4027), .ZN(n3746) );
  INV_X1 U4528 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3736) );
  OAI22_X1 U4529 ( .A1(n3974), .A2(n4336), .B1(n4334), .B2(n3736), .ZN(n3737)
         );
  AOI21_X1 U4530 ( .B1(n4143), .B2(n4340), .A(n3737), .ZN(n3745) );
  NOR2_X1 U4531 ( .A1(n3738), .A2(n4792), .ZN(n3739) );
  NOR2_X1 U4532 ( .A1(n3740), .A2(n3739), .ZN(n3741) );
  OAI21_X1 U4533 ( .B1(n3742), .B2(n4342), .A(n3741), .ZN(n3743) );
  NAND2_X1 U4534 ( .A1(n3743), .A2(n4334), .ZN(n3744) );
  OAI211_X1 U4535 ( .C1(n3746), .C2(n4361), .A(n3745), .B(n3744), .ZN(U3354)
         );
  INV_X1 U4536 ( .A(n3747), .ZN(n3751) );
  AOI21_X1 U4537 ( .B1(n3747), .B2(n3749), .A(n3748), .ZN(n3750) );
  AOI21_X1 U4538 ( .B1(n3751), .B2(n3850), .A(n3750), .ZN(n3755) );
  NAND2_X1 U4539 ( .A1(n3753), .A2(n3752), .ZN(n3754) );
  XNOR2_X1 U4540 ( .A(n3755), .B(n3754), .ZN(n3761) );
  INV_X1 U4541 ( .A(n4474), .ZN(n3800) );
  NAND2_X1 U4542 ( .A1(U3149), .A2(REG3_REG_14__SCAN_IN), .ZN(n4730) );
  OAI21_X1 U4543 ( .B1(n3865), .B2(n3800), .A(n4730), .ZN(n3758) );
  OAI22_X1 U4544 ( .A1(n3900), .A2(n3756), .B1(n4463), .B2(n3898), .ZN(n3757)
         );
  AOI211_X1 U4545 ( .C1(n3904), .C2(n3759), .A(n3758), .B(n3757), .ZN(n3760)
         );
  OAI21_X1 U4546 ( .B1(n3761), .B2(n3907), .A(n3760), .ZN(U3212) );
  NAND2_X1 U4547 ( .A1(n3762), .A2(n3876), .ZN(n3773) );
  OR2_X2 U4548 ( .A1(n3763), .A2(n3764), .ZN(n3766) );
  NAND2_X1 U4549 ( .A1(n3766), .A2(n3765), .ZN(n3863) );
  AOI21_X1 U4550 ( .B1(n3861), .B2(n3768), .A(n3767), .ZN(n3772) );
  INV_X1 U4551 ( .A(n4247), .ZN(n4407) );
  OAI22_X1 U4552 ( .A1(n4407), .A2(n3865), .B1(n3900), .B2(n4216), .ZN(n3770)
         );
  OAI22_X1 U4553 ( .A1(n4210), .A2(n3898), .B1(STATE_REG_SCAN_IN), .B2(n4535), 
        .ZN(n3769) );
  AOI211_X1 U4554 ( .C1(n4217), .C2(n3904), .A(n3770), .B(n3769), .ZN(n3771)
         );
  OAI21_X1 U4555 ( .B1(n3773), .B2(n3772), .A(n3771), .ZN(U3213) );
  NAND2_X1 U4556 ( .A1(n3874), .A2(n3873), .ZN(n3775) );
  NAND2_X1 U4557 ( .A1(n3775), .A2(n3872), .ZN(n3776) );
  XOR2_X1 U4558 ( .A(n3777), .B(n3776), .Z(n3783) );
  INV_X1 U4559 ( .A(n3778), .ZN(n4302) );
  INV_X1 U4560 ( .A(n4405), .ZN(n4295) );
  OAI21_X1 U4561 ( .B1(n4295), .B2(n3898), .A(n3779), .ZN(n3781) );
  OAI22_X1 U4562 ( .A1(n3900), .A2(n4301), .B1(n4434), .B2(n3865), .ZN(n3780)
         );
  AOI211_X1 U4563 ( .C1(n3904), .C2(n4302), .A(n3781), .B(n3780), .ZN(n3782)
         );
  OAI21_X1 U4564 ( .B1(n3783), .B2(n3907), .A(n3782), .ZN(U3216) );
  XNOR2_X1 U4565 ( .A(n3785), .B(n3784), .ZN(n3786) );
  XNOR2_X1 U4566 ( .A(n3763), .B(n3786), .ZN(n3791) );
  AOI22_X1 U4567 ( .A1(n4247), .A2(n3890), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3789) );
  OAI22_X1 U4568 ( .A1(n3900), .A2(n4245), .B1(n4295), .B2(n3865), .ZN(n3787)
         );
  INV_X1 U4569 ( .A(n3787), .ZN(n3788) );
  OAI211_X1 U4570 ( .C1(n3886), .C2(n4248), .A(n3789), .B(n3788), .ZN(n3790)
         );
  AOI21_X1 U4571 ( .B1(n3791), .B2(n3876), .A(n3790), .ZN(n3792) );
  INV_X1 U4572 ( .A(n3792), .ZN(U3220) );
  INV_X1 U4573 ( .A(n3794), .ZN(n3796) );
  NOR2_X1 U4574 ( .A1(n3796), .A2(n3795), .ZN(n3797) );
  XNOR2_X1 U4575 ( .A(n3793), .B(n3797), .ZN(n3805) );
  OAI21_X1 U4576 ( .B1(n3865), .B2(n3799), .A(n3798), .ZN(n3802) );
  OAI22_X1 U4577 ( .A1(n3900), .A2(n4478), .B1(n3800), .B2(n3898), .ZN(n3801)
         );
  AOI211_X1 U4578 ( .C1(n3904), .C2(n3803), .A(n3802), .B(n3801), .ZN(n3804)
         );
  OAI21_X1 U4579 ( .B1(n3805), .B2(n3907), .A(n3804), .ZN(U3221) );
  NAND2_X1 U4580 ( .A1(n2030), .A2(n3806), .ZN(n3893) );
  NOR2_X1 U4581 ( .A1(n2030), .A2(n3806), .ZN(n3895) );
  AOI21_X1 U4582 ( .B1(n3816), .B2(n3893), .A(n3895), .ZN(n3809) );
  XNOR2_X1 U4583 ( .A(n3808), .B(n3807), .ZN(n3815) );
  XNOR2_X1 U4584 ( .A(n3809), .B(n3815), .ZN(n3814) );
  NOR2_X1 U4585 ( .A1(n4610), .A2(STATE_REG_SCAN_IN), .ZN(n4755) );
  INV_X1 U4586 ( .A(n4441), .ZN(n3810) );
  OAI22_X1 U4587 ( .A1(n3900), .A2(n4443), .B1(n3810), .B2(n3898), .ZN(n3811)
         );
  AOI211_X1 U4588 ( .C1(n3902), .C2(n4440), .A(n4755), .B(n3811), .ZN(n3813)
         );
  NAND2_X1 U4589 ( .A1(n3904), .A2(n4353), .ZN(n3812) );
  OAI211_X1 U4590 ( .C1(n3814), .C2(n3907), .A(n3813), .B(n3812), .ZN(U3223)
         );
  OAI211_X1 U4591 ( .C1(n3895), .C2(n3816), .A(n3815), .B(n3893), .ZN(n3818)
         );
  NAND2_X1 U4592 ( .A1(n3818), .A2(n3817), .ZN(n3822) );
  XNOR2_X1 U4593 ( .A(n3820), .B(n3819), .ZN(n3821) );
  XNOR2_X1 U4594 ( .A(n3822), .B(n3821), .ZN(n3823) );
  NAND2_X1 U4595 ( .A1(n3823), .A2(n3876), .ZN(n3826) );
  AND2_X1 U4596 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4108) );
  OAI22_X1 U4597 ( .A1(n3900), .A2(n4335), .B1(n4434), .B2(n3898), .ZN(n3824)
         );
  AOI211_X1 U4598 ( .C1(n3902), .C2(n4432), .A(n4108), .B(n3824), .ZN(n3825)
         );
  OAI211_X1 U4599 ( .C1(n3886), .C2(n4333), .A(n3826), .B(n3825), .ZN(U3225)
         );
  INV_X1 U4600 ( .A(n3827), .ZN(n3828) );
  NOR2_X1 U4601 ( .A1(n3829), .A2(n3828), .ZN(n3831) );
  XNOR2_X1 U4602 ( .A(n3831), .B(n3830), .ZN(n3837) );
  INV_X1 U4603 ( .A(n3832), .ZN(n4193) );
  INV_X1 U4604 ( .A(n4224), .ZN(n4391) );
  OAI22_X1 U4605 ( .A1(n4391), .A2(n3865), .B1(n3900), .B2(n4195), .ZN(n3835)
         );
  OAI22_X1 U4606 ( .A1(n4196), .A2(n3898), .B1(STATE_REG_SCAN_IN), .B2(n3833), 
        .ZN(n3834) );
  AOI211_X1 U4607 ( .C1(n4193), .C2(n3904), .A(n3835), .B(n3834), .ZN(n3836)
         );
  OAI21_X1 U4608 ( .B1(n3837), .B2(n3907), .A(n3836), .ZN(U3226) );
  INV_X1 U4609 ( .A(n3838), .ZN(n3843) );
  AOI21_X1 U4610 ( .B1(n3842), .B2(n3840), .A(n3839), .ZN(n3841) );
  AOI21_X1 U4611 ( .B1(n3843), .B2(n3842), .A(n3841), .ZN(n3848) );
  INV_X1 U4612 ( .A(n4416), .ZN(n4310) );
  OAI22_X1 U4613 ( .A1(n3900), .A2(n4277), .B1(n4310), .B2(n3865), .ZN(n3846)
         );
  OAI22_X1 U4614 ( .A1(n3866), .A2(n3898), .B1(STATE_REG_SCAN_IN), .B2(n3844), 
        .ZN(n3845) );
  AOI211_X1 U4615 ( .C1(n3904), .C2(n4274), .A(n3846), .B(n3845), .ZN(n3847)
         );
  OAI21_X1 U4616 ( .B1(n3848), .B2(n3907), .A(n3847), .ZN(U3230) );
  XNOR2_X1 U4617 ( .A(n3850), .B(n3849), .ZN(n3851) );
  XNOR2_X1 U4618 ( .A(n3747), .B(n3851), .ZN(n3860) );
  OAI21_X1 U4619 ( .B1(n3865), .B2(n3853), .A(n3852), .ZN(n3857) );
  OAI22_X1 U4620 ( .A1(n3900), .A2(n3855), .B1(n3854), .B2(n3898), .ZN(n3856)
         );
  AOI211_X1 U4621 ( .C1(n3904), .C2(n3858), .A(n3857), .B(n3856), .ZN(n3859)
         );
  OAI21_X1 U4622 ( .B1(n3860), .B2(n3907), .A(n3859), .ZN(U3231) );
  INV_X1 U4623 ( .A(n3861), .ZN(n3862) );
  AOI21_X1 U4624 ( .B1(n3864), .B2(n3863), .A(n3862), .ZN(n3871) );
  OAI22_X1 U4625 ( .A1(n3866), .A2(n3865), .B1(STATE_REG_SCAN_IN), .B2(n4579), 
        .ZN(n3869) );
  OAI22_X1 U4626 ( .A1(n4391), .A2(n3898), .B1(n3900), .B2(n3867), .ZN(n3868)
         );
  AOI211_X1 U4627 ( .C1(n4234), .C2(n3904), .A(n3869), .B(n3868), .ZN(n3870)
         );
  OAI21_X1 U4628 ( .B1(n3871), .B2(n3907), .A(n3870), .ZN(U3232) );
  NAND2_X1 U4629 ( .A1(n3873), .A2(n3872), .ZN(n3875) );
  XOR2_X1 U4630 ( .A(n3875), .B(n3874), .Z(n3877) );
  NAND2_X1 U4631 ( .A1(n3877), .A2(n3876), .ZN(n3880) );
  AND2_X1 U4632 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4764) );
  OAI22_X1 U4633 ( .A1(n3900), .A2(n4315), .B1(n4310), .B2(n3898), .ZN(n3878)
         );
  AOI211_X1 U4634 ( .C1(n3902), .C2(n4441), .A(n4764), .B(n3878), .ZN(n3879)
         );
  OAI211_X1 U4635 ( .C1(n3886), .C2(n4316), .A(n3880), .B(n3879), .ZN(U3235)
         );
  INV_X1 U4636 ( .A(n3881), .ZN(n3883) );
  NAND2_X1 U4637 ( .A1(n3883), .A2(n3882), .ZN(n3884) );
  XNOR2_X1 U4638 ( .A(n3885), .B(n3884), .ZN(n3892) );
  NOR2_X1 U4639 ( .A1(n4161), .A2(n3886), .ZN(n3889) );
  AOI22_X1 U4640 ( .A1(n4387), .A2(n3902), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3887) );
  OAI21_X1 U4641 ( .B1(n3900), .B2(n4159), .A(n3887), .ZN(n3888) );
  AOI211_X1 U4642 ( .C1(n3890), .C2(n4124), .A(n3889), .B(n3888), .ZN(n3891)
         );
  OAI21_X1 U4643 ( .B1(n3892), .B2(n3907), .A(n3891), .ZN(U3237) );
  INV_X1 U4644 ( .A(n3893), .ZN(n3894) );
  NOR2_X1 U4645 ( .A1(n3895), .A2(n3894), .ZN(n3897) );
  XNOR2_X1 U4646 ( .A(n3897), .B(n3896), .ZN(n3908) );
  NOR2_X1 U4647 ( .A1(n4547), .A2(STATE_REG_SCAN_IN), .ZN(n4744) );
  OAI22_X1 U4648 ( .A1(n3900), .A2(n3899), .B1(n4452), .B2(n3898), .ZN(n3901)
         );
  AOI211_X1 U4649 ( .C1(n3902), .C2(n4450), .A(n4744), .B(n3901), .ZN(n3906)
         );
  NAND2_X1 U4650 ( .A1(n3904), .A2(n3903), .ZN(n3905) );
  OAI211_X1 U4651 ( .C1(n3908), .C2(n3907), .A(n3906), .B(n3905), .ZN(U3238)
         );
  OAI211_X1 U4652 ( .C1(n3911), .C2(n4715), .A(n3910), .B(n3909), .ZN(n3914)
         );
  NAND3_X1 U4653 ( .A1(n3914), .A2(n3913), .A3(n3912), .ZN(n3917) );
  NAND3_X1 U4654 ( .A1(n3917), .A2(n3916), .A3(n3915), .ZN(n3920) );
  NAND3_X1 U4655 ( .A1(n3920), .A2(n3919), .A3(n3918), .ZN(n3922) );
  NAND4_X1 U4656 ( .A1(n3922), .A2(n3921), .A3(n3936), .A4(n2047), .ZN(n3925)
         );
  NAND3_X1 U4657 ( .A1(n3925), .A2(n3924), .A3(n3923), .ZN(n3931) );
  AND2_X1 U4658 ( .A1(n3927), .A2(n3926), .ZN(n3935) );
  INV_X1 U4659 ( .A(n3928), .ZN(n3929) );
  AOI211_X1 U4660 ( .C1(n3931), .C2(n3935), .A(n3930), .B(n3929), .ZN(n3934)
         );
  NAND2_X1 U4661 ( .A1(n3933), .A2(n3932), .ZN(n3940) );
  NOR3_X1 U4662 ( .A1(n3934), .A2(n3938), .A3(n3940), .ZN(n3947) );
  INV_X1 U4663 ( .A(n3935), .ZN(n3939) );
  OR4_X1 U4664 ( .A1(n3939), .A2(n3938), .A3(n2169), .A4(n3937), .ZN(n3942) );
  NAND2_X1 U4665 ( .A1(n3940), .A2(n3949), .ZN(n4030) );
  INV_X1 U4666 ( .A(n4030), .ZN(n3941) );
  AOI21_X1 U4667 ( .B1(n3943), .B2(n3942), .A(n3941), .ZN(n3946) );
  OAI211_X1 U4668 ( .C1(n3947), .C2(n3946), .A(n3945), .B(n3944), .ZN(n3954)
         );
  INV_X1 U4669 ( .A(n3948), .ZN(n3951) );
  NAND2_X1 U4670 ( .A1(n3950), .A2(n3949), .ZN(n4031) );
  OAI21_X1 U4671 ( .B1(n3951), .B2(n4031), .A(n4030), .ZN(n3953) );
  AOI21_X1 U4672 ( .B1(n3954), .B2(n3953), .A(n2186), .ZN(n3959) );
  INV_X1 U4673 ( .A(n4033), .ZN(n3958) );
  OR2_X1 U4674 ( .A1(n3956), .A2(n3955), .ZN(n4032) );
  INV_X1 U4675 ( .A(n4032), .ZN(n3957) );
  OAI21_X1 U4676 ( .B1(n3959), .B2(n3958), .A(n3957), .ZN(n3960) );
  AOI21_X1 U4677 ( .B1(n3960), .B2(n4035), .A(n4002), .ZN(n3963) );
  OAI21_X1 U4678 ( .B1(n3963), .B2(n3962), .A(n3961), .ZN(n3971) );
  NOR3_X1 U4679 ( .A1(n4045), .A2(n4040), .A3(n4022), .ZN(n3970) );
  OAI21_X1 U4680 ( .B1(n3966), .B2(n3965), .A(n3964), .ZN(n4049) );
  OAI21_X1 U4681 ( .B1(n4157), .B2(n3968), .A(n3967), .ZN(n3969) );
  AOI211_X1 U4682 ( .C1(n3971), .C2(n3970), .A(n4049), .B(n3969), .ZN(n3984)
         );
  NAND2_X1 U4683 ( .A1(n3973), .A2(n3972), .ZN(n4046) );
  INV_X1 U4684 ( .A(n4046), .ZN(n3978) );
  OR2_X1 U4685 ( .A1(n4125), .A2(n3974), .ZN(n3976) );
  INV_X1 U4686 ( .A(n4119), .ZN(n4053) );
  NAND2_X1 U4687 ( .A1(n4072), .A2(n4057), .ZN(n3979) );
  OAI21_X1 U4688 ( .B1(n3980), .B2(n4053), .A(n3979), .ZN(n4008) );
  INV_X1 U4689 ( .A(n4008), .ZN(n3975) );
  NAND2_X1 U4690 ( .A1(n3976), .A2(n3975), .ZN(n4044) );
  INV_X1 U4691 ( .A(n4044), .ZN(n3977) );
  INV_X1 U4692 ( .A(n3979), .ZN(n3983) );
  AND2_X1 U4693 ( .A1(n3980), .A2(n4053), .ZN(n4029) );
  INV_X1 U4694 ( .A(n4029), .ZN(n3981) );
  OAI21_X1 U4695 ( .B1(n4072), .B2(n4057), .A(n3981), .ZN(n4009) );
  INV_X1 U4696 ( .A(n4009), .ZN(n3982) );
  OAI22_X1 U4697 ( .A1(n3984), .A2(n4050), .B1(n3983), .B2(n3982), .ZN(n4062)
         );
  INV_X1 U4698 ( .A(n4167), .ZN(n3985) );
  NOR2_X1 U4699 ( .A1(n4040), .A2(n3985), .ZN(n4189) );
  NAND4_X1 U4700 ( .A1(n3989), .A2(n3988), .A3(n3987), .A4(n3986), .ZN(n3995)
         );
  NAND4_X1 U4701 ( .A1(n3993), .A2(n3992), .A3(n3991), .A4(n3990), .ZN(n3994)
         );
  NOR2_X1 U4702 ( .A1(n3995), .A2(n3994), .ZN(n4001) );
  NOR4_X1 U4703 ( .A1(n4261), .A2(n3998), .A3(n3997), .A4(n3996), .ZN(n3999)
         );
  NAND4_X1 U4704 ( .A1(n4230), .A2(n4001), .A3(n4000), .A4(n3999), .ZN(n4017)
         );
  INV_X1 U4705 ( .A(n4002), .ZN(n4003) );
  NAND2_X1 U4706 ( .A1(n4005), .A2(n4004), .ZN(n4271) );
  NOR2_X1 U4707 ( .A1(n4783), .A2(n4006), .ZN(n4007) );
  AND2_X1 U4708 ( .A1(n4271), .A2(n4007), .ZN(n4014) );
  NAND2_X1 U4709 ( .A1(n4264), .A2(n4263), .ZN(n4296) );
  NOR2_X1 U4710 ( .A1(n4009), .A2(n4008), .ZN(n4012) );
  NAND2_X1 U4711 ( .A1(n4284), .A2(n4283), .ZN(n4329) );
  NOR2_X1 U4712 ( .A1(n4329), .A2(n4010), .ZN(n4011) );
  AND4_X1 U4713 ( .A1(n4296), .A2(n4012), .A3(n4357), .A4(n4011), .ZN(n4013)
         );
  NAND4_X1 U4714 ( .A1(n4243), .A2(n4015), .A3(n4014), .A4(n4013), .ZN(n4016)
         );
  NOR2_X1 U4715 ( .A1(n4017), .A2(n4016), .ZN(n4018) );
  AND2_X1 U4716 ( .A1(n4189), .A2(n4018), .ZN(n4025) );
  XNOR2_X1 U4717 ( .A(n4137), .B(n4154), .ZN(n4151) );
  NAND2_X1 U4718 ( .A1(n4148), .A2(n4019), .ZN(n4171) );
  INV_X1 U4719 ( .A(n4171), .ZN(n4024) );
  INV_X1 U4720 ( .A(n4020), .ZN(n4021) );
  OR2_X1 U4721 ( .A1(n4022), .A2(n4021), .ZN(n4212) );
  INV_X1 U4722 ( .A(n4212), .ZN(n4023) );
  AND4_X1 U4723 ( .A1(n4025), .A2(n4151), .A3(n4024), .A4(n4023), .ZN(n4026)
         );
  NAND4_X1 U4724 ( .A1(n2776), .A2(n4052), .A3(n4027), .A4(n4026), .ZN(n4060)
         );
  INV_X1 U4725 ( .A(n4072), .ZN(n4028) );
  NOR2_X1 U4726 ( .A1(n4029), .A2(n4028), .ZN(n4058) );
  OAI21_X1 U4727 ( .B1(n3643), .B2(n4031), .A(n4030), .ZN(n4034) );
  AOI211_X1 U4728 ( .C1(n4034), .C2(n4033), .A(n2186), .B(n4032), .ZN(n4038)
         );
  INV_X1 U4729 ( .A(n4035), .ZN(n4037) );
  OAI21_X1 U4730 ( .B1(n4038), .B2(n4037), .A(n4036), .ZN(n4043) );
  INV_X1 U4731 ( .A(n4039), .ZN(n4041) );
  NOR2_X1 U4732 ( .A1(n4041), .A2(n4040), .ZN(n4042) );
  AOI21_X1 U4733 ( .B1(n4043), .B2(n4042), .A(n4149), .ZN(n4047) );
  NOR4_X1 U4734 ( .A1(n4047), .A2(n4046), .A3(n4045), .A4(n4044), .ZN(n4055)
         );
  NOR2_X1 U4735 ( .A1(n4049), .A2(n4048), .ZN(n4051) );
  AOI21_X1 U4736 ( .B1(n4052), .B2(n4051), .A(n4050), .ZN(n4054) );
  OAI22_X1 U4737 ( .A1(n4055), .A2(n4054), .B1(n4072), .B2(n4053), .ZN(n4056)
         );
  OAI21_X1 U4738 ( .B1(n4058), .B2(n4057), .A(n4056), .ZN(n4059) );
  MUX2_X1 U4739 ( .A(n4060), .B(n4059), .S(n4715), .Z(n4061) );
  XNOR2_X1 U4740 ( .A(n4064), .B(n4063), .ZN(n4071) );
  INV_X1 U4741 ( .A(n4065), .ZN(n4066) );
  NOR2_X1 U4742 ( .A1(n4067), .A2(n4066), .ZN(n4069) );
  OAI21_X1 U4743 ( .B1(n4070), .B2(n4714), .A(B_REG_SCAN_IN), .ZN(n4068) );
  OAI22_X1 U4744 ( .A1(n4071), .A2(n4070), .B1(n4069), .B2(n4068), .ZN(U3239)
         );
  MUX2_X1 U4745 ( .A(DATAO_REG_31__SCAN_IN), .B(n4072), .S(n4077), .Z(U3581)
         );
  MUX2_X1 U4746 ( .A(DATAO_REG_29__SCAN_IN), .B(n4125), .S(n4077), .Z(U3579)
         );
  MUX2_X1 U4747 ( .A(DATAO_REG_28__SCAN_IN), .B(n4143), .S(n4077), .Z(U3578)
         );
  MUX2_X1 U4748 ( .A(DATAO_REG_27__SCAN_IN), .B(n4124), .S(n4077), .Z(U3577)
         );
  MUX2_X1 U4749 ( .A(DATAO_REG_24__SCAN_IN), .B(n4378), .S(n4077), .Z(U3574)
         );
  MUX2_X1 U4750 ( .A(DATAO_REG_23__SCAN_IN), .B(n4224), .S(n4077), .Z(U3573)
         );
  MUX2_X1 U4751 ( .A(DATAO_REG_22__SCAN_IN), .B(n4247), .S(n4077), .Z(U3572)
         );
  MUX2_X1 U4752 ( .A(DATAO_REG_20__SCAN_IN), .B(n4405), .S(n4077), .Z(U3570)
         );
  MUX2_X1 U4753 ( .A(DATAO_REG_19__SCAN_IN), .B(n4416), .S(n4077), .Z(U3569)
         );
  MUX2_X1 U4754 ( .A(DATAO_REG_18__SCAN_IN), .B(n4292), .S(n4077), .Z(U3568)
         );
  MUX2_X1 U4755 ( .A(DATAO_REG_17__SCAN_IN), .B(n4441), .S(n4077), .Z(U3567)
         );
  MUX2_X1 U4756 ( .A(DATAO_REG_16__SCAN_IN), .B(n4432), .S(n4077), .Z(U3566)
         );
  MUX2_X1 U4757 ( .A(DATAO_REG_14__SCAN_IN), .B(n4450), .S(n4077), .Z(U3564)
         );
  MUX2_X1 U4758 ( .A(DATAO_REG_13__SCAN_IN), .B(n4474), .S(n4077), .Z(U3563)
         );
  MUX2_X1 U4759 ( .A(DATAO_REG_12__SCAN_IN), .B(n4073), .S(n4077), .Z(U3562)
         );
  MUX2_X1 U4760 ( .A(DATAO_REG_11__SCAN_IN), .B(n4473), .S(n4077), .Z(U3561)
         );
  MUX2_X1 U4761 ( .A(DATAO_REG_10__SCAN_IN), .B(n4485), .S(n4077), .Z(U3560)
         );
  MUX2_X1 U4762 ( .A(DATAO_REG_8__SCAN_IN), .B(n4074), .S(n4077), .Z(U3558) );
  MUX2_X1 U4763 ( .A(DATAO_REG_7__SCAN_IN), .B(n4075), .S(n4077), .Z(U3557) );
  MUX2_X1 U4764 ( .A(DATAO_REG_5__SCAN_IN), .B(n2016), .S(n4077), .Z(U3555) );
  MUX2_X1 U4765 ( .A(DATAO_REG_4__SCAN_IN), .B(n2861), .S(n4077), .Z(U3554) );
  MUX2_X1 U4766 ( .A(DATAO_REG_2__SCAN_IN), .B(n2840), .S(n4077), .Z(U3552) );
  MUX2_X1 U4767 ( .A(DATAO_REG_1__SCAN_IN), .B(n2459), .S(n4077), .Z(U3551) );
  MUX2_X1 U4768 ( .A(DATAO_REG_0__SCAN_IN), .B(n2823), .S(n4077), .Z(U3550) );
  OAI211_X1 U4769 ( .C1(n4080), .C2(n4079), .A(n4770), .B(n4078), .ZN(n4086)
         );
  OAI211_X1 U4770 ( .C1(n2381), .C2(n4082), .A(n4096), .B(n3187), .ZN(n4085)
         );
  AOI22_X1 U4771 ( .A1(n4765), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4084) );
  NAND2_X1 U4772 ( .A1(n4110), .A2(n4728), .ZN(n4083) );
  NAND4_X1 U4773 ( .A1(n4086), .A2(n4085), .A3(n4084), .A4(n4083), .ZN(U3241)
         );
  INV_X1 U4774 ( .A(n4087), .ZN(n4089) );
  AOI21_X1 U4775 ( .B1(n4089), .B2(n4088), .A(n4113), .ZN(n4091) );
  NAND2_X1 U4776 ( .A1(n4091), .A2(n4090), .ZN(n4102) );
  INV_X1 U4777 ( .A(ADDR_REG_11__SCAN_IN), .ZN(n4093) );
  OAI21_X1 U4778 ( .B1(n4094), .B2(n4093), .A(n4092), .ZN(n4095) );
  AOI21_X1 U4779 ( .B1(n2291), .B2(n4110), .A(n4095), .ZN(n4101) );
  OAI211_X1 U4780 ( .C1(n4099), .C2(n4098), .A(n4097), .B(n4096), .ZN(n4100)
         );
  NAND3_X1 U4781 ( .A1(n4102), .A2(n4101), .A3(n4100), .ZN(U3251) );
  AOI21_X1 U4782 ( .B1(n4103), .B2(n4105), .A(n4104), .ZN(n4114) );
  NAND2_X1 U4783 ( .A1(n4110), .A2(n4109), .ZN(n4111) );
  OAI211_X1 U4784 ( .C1(n4114), .C2(n4113), .A(n4112), .B(n4111), .ZN(U3257)
         );
  INV_X1 U4785 ( .A(n4115), .ZN(n4116) );
  AOI21_X1 U4786 ( .B1(n4119), .B2(n4458), .A(n4116), .ZN(n4654) );
  NAND2_X1 U4787 ( .A1(n4651), .A2(n4779), .ZN(n4121) );
  NAND2_X1 U4788 ( .A1(n4365), .A2(REG2_REG_30__SCAN_IN), .ZN(n4120) );
  OAI211_X1 U4789 ( .C1(n4788), .C2(n4654), .A(n4121), .B(n4120), .ZN(U3261)
         );
  NAND2_X1 U4790 ( .A1(n4122), .A2(n4344), .ZN(n4133) );
  INV_X1 U4791 ( .A(n4123), .ZN(n4131) );
  AOI22_X1 U4792 ( .A1(n4350), .A2(n4125), .B1(n4124), .B2(n4340), .ZN(n4128)
         );
  AOI22_X1 U4793 ( .A1(n4126), .A2(n4776), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4788), .ZN(n4127) );
  OAI211_X1 U4794 ( .C1(n4129), .C2(n4336), .A(n4128), .B(n4127), .ZN(n4130)
         );
  AOI21_X1 U4795 ( .B1(n4131), .B2(n4779), .A(n4130), .ZN(n4132) );
  OAI211_X1 U4796 ( .C1(n4365), .C2(n4134), .A(n4133), .B(n4132), .ZN(U3262)
         );
  NAND2_X1 U4797 ( .A1(n4135), .A2(n4344), .ZN(n4145) );
  AOI22_X1 U4798 ( .A1(n4136), .A2(n4776), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4788), .ZN(n4139) );
  NAND2_X1 U4799 ( .A1(n4137), .A2(n4340), .ZN(n4138) );
  OAI211_X1 U4800 ( .C1(n4336), .C2(n4140), .A(n4139), .B(n4138), .ZN(n4142)
         );
  NOR2_X1 U4801 ( .A1(n4372), .A2(n4342), .ZN(n4141) );
  AOI211_X1 U4802 ( .C1(n4350), .C2(n4143), .A(n4142), .B(n4141), .ZN(n4144)
         );
  OAI211_X1 U4803 ( .C1(n4365), .C2(n4146), .A(n4145), .B(n4144), .ZN(U3263)
         );
  XNOR2_X1 U4804 ( .A(n4147), .B(n4151), .ZN(n4374) );
  INV_X1 U4805 ( .A(n4374), .ZN(n4166) );
  OAI21_X1 U4806 ( .B1(n4150), .B2(n4149), .A(n4148), .ZN(n4152) );
  XNOR2_X1 U4807 ( .A(n4152), .B(n4151), .ZN(n4153) );
  NAND2_X1 U4808 ( .A1(n4153), .A2(n4465), .ZN(n4156) );
  AOI22_X1 U4809 ( .A1(n4387), .A2(n4486), .B1(n4154), .B2(n4458), .ZN(n4155)
         );
  OAI211_X1 U4810 ( .C1(n4157), .C2(n4462), .A(n4156), .B(n4155), .ZN(n4373)
         );
  INV_X1 U4811 ( .A(n4174), .ZN(n4160) );
  INV_X1 U4812 ( .A(n2771), .ZN(n4158) );
  OAI21_X1 U4813 ( .B1(n4160), .B2(n4159), .A(n4158), .ZN(n4658) );
  INV_X1 U4814 ( .A(n4161), .ZN(n4162) );
  AOI22_X1 U4815 ( .A1(n4162), .A2(n4776), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4365), .ZN(n4163) );
  OAI21_X1 U4816 ( .B1(n4658), .B2(n4342), .A(n4163), .ZN(n4164) );
  AOI21_X1 U4817 ( .B1(n4373), .B2(n4334), .A(n4164), .ZN(n4165) );
  OAI21_X1 U4818 ( .B1(n4166), .B2(n4361), .A(n4165), .ZN(U3264) );
  NAND2_X1 U4819 ( .A1(n4168), .A2(n4167), .ZN(n4169) );
  XNOR2_X1 U4820 ( .A(n4169), .B(n4171), .ZN(n4170) );
  NAND2_X1 U4821 ( .A1(n4170), .A2(n4465), .ZN(n4380) );
  XNOR2_X1 U4822 ( .A(n4172), .B(n4171), .ZN(n4383) );
  NAND2_X1 U4823 ( .A1(n4383), .A2(n4344), .ZN(n4182) );
  NAND2_X1 U4824 ( .A1(n4192), .A2(n4377), .ZN(n4173) );
  NAND2_X1 U4825 ( .A1(n4174), .A2(n4173), .ZN(n4662) );
  INV_X1 U4826 ( .A(n4662), .ZN(n4180) );
  AOI22_X1 U4827 ( .A1(n4175), .A2(n4776), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4788), .ZN(n4176) );
  OAI21_X1 U4828 ( .B1(n4210), .B2(n4356), .A(n4176), .ZN(n4179) );
  OAI22_X1 U4829 ( .A1(n4381), .A2(n4337), .B1(n4336), .B2(n4177), .ZN(n4178)
         );
  AOI211_X1 U4830 ( .C1(n4180), .C2(n4779), .A(n4179), .B(n4178), .ZN(n4181)
         );
  OAI211_X1 U4831 ( .C1(n4788), .C2(n4380), .A(n4182), .B(n4181), .ZN(U3265)
         );
  XNOR2_X1 U4832 ( .A(n4183), .B(n4189), .ZN(n4184) );
  NAND2_X1 U4833 ( .A1(n4184), .A2(n4465), .ZN(n4389) );
  NAND2_X1 U4834 ( .A1(n4185), .A2(n4186), .ZN(n4188) );
  AND2_X1 U4835 ( .A1(n4188), .A2(n4187), .ZN(n4190) );
  XNOR2_X1 U4836 ( .A(n4190), .B(n4189), .ZN(n4393) );
  NAND2_X1 U4837 ( .A1(n4393), .A2(n4344), .ZN(n4201) );
  OAI21_X1 U4838 ( .B1(n4191), .B2(n4195), .A(n4192), .ZN(n4666) );
  INV_X1 U4839 ( .A(n4666), .ZN(n4199) );
  AOI22_X1 U4840 ( .A1(n4193), .A2(n4776), .B1(REG2_REG_24__SCAN_IN), .B2(
        n4788), .ZN(n4194) );
  OAI21_X1 U4841 ( .B1(n4391), .B2(n4356), .A(n4194), .ZN(n4198) );
  OAI22_X1 U4842 ( .A1(n4196), .A2(n4337), .B1(n4195), .B2(n4336), .ZN(n4197)
         );
  AOI211_X1 U4843 ( .C1(n4199), .C2(n4779), .A(n4198), .B(n4197), .ZN(n4200)
         );
  OAI211_X1 U4844 ( .C1(n4365), .C2(n4389), .A(n4201), .B(n4200), .ZN(U3266)
         );
  INV_X1 U4845 ( .A(n4202), .ZN(n4203) );
  AOI21_X1 U4846 ( .B1(n4238), .B2(n4243), .A(n4203), .ZN(n4223) );
  OAI21_X1 U4847 ( .B1(n4223), .B2(n4222), .A(n4204), .ZN(n4205) );
  XOR2_X1 U4848 ( .A(n4212), .B(n4205), .Z(n4206) );
  NAND2_X1 U4849 ( .A1(n4206), .A2(n4465), .ZN(n4209) );
  AOI22_X1 U4850 ( .A1(n4247), .A2(n4486), .B1(n4458), .B2(n4207), .ZN(n4208)
         );
  OAI211_X1 U4851 ( .C1(n4210), .C2(n4462), .A(n4209), .B(n4208), .ZN(n4395)
         );
  INV_X1 U4852 ( .A(n4395), .ZN(n4221) );
  NAND2_X1 U4853 ( .A1(n4185), .A2(n4211), .ZN(n4213) );
  XOR2_X1 U4854 ( .A(n4213), .B(n4212), .Z(n4396) );
  INV_X1 U4855 ( .A(n4191), .ZN(n4215) );
  OAI21_X1 U4856 ( .B1(n4214), .B2(n4216), .A(n4215), .ZN(n4670) );
  AOI22_X1 U4857 ( .A1(n4217), .A2(n4776), .B1(n4365), .B2(
        REG2_REG_23__SCAN_IN), .ZN(n4218) );
  OAI21_X1 U4858 ( .B1(n4670), .B2(n4342), .A(n4218), .ZN(n4219) );
  AOI21_X1 U4859 ( .B1(n4396), .B2(n4344), .A(n4219), .ZN(n4220) );
  OAI21_X1 U4860 ( .B1(n4221), .B2(n4365), .A(n4220), .ZN(U3267) );
  XNOR2_X1 U4861 ( .A(n4223), .B(n4222), .ZN(n4228) );
  NAND2_X1 U4862 ( .A1(n4224), .A2(n4475), .ZN(n4226) );
  AOI22_X1 U4863 ( .A1(n4414), .A2(n4486), .B1(n4232), .B2(n4458), .ZN(n4225)
         );
  NAND2_X1 U4864 ( .A1(n4226), .A2(n4225), .ZN(n4227) );
  AOI21_X1 U4865 ( .B1(n4228), .B2(n4465), .A(n4227), .ZN(n4401) );
  NAND2_X1 U4866 ( .A1(n4229), .A2(n4230), .ZN(n4231) );
  AND2_X1 U4867 ( .A1(n4185), .A2(n4231), .ZN(n4399) );
  AND2_X1 U4868 ( .A1(n4244), .A2(n4232), .ZN(n4233) );
  OR2_X1 U4869 ( .A1(n4233), .A2(n4214), .ZN(n4674) );
  AOI22_X1 U4870 ( .A1(n4234), .A2(n4776), .B1(n4365), .B2(
        REG2_REG_22__SCAN_IN), .ZN(n4235) );
  OAI21_X1 U4871 ( .B1(n4674), .B2(n4342), .A(n4235), .ZN(n4236) );
  AOI21_X1 U4872 ( .B1(n4399), .B2(n4344), .A(n4236), .ZN(n4237) );
  OAI21_X1 U4873 ( .B1(n4401), .B2(n4365), .A(n4237), .ZN(U3268) );
  XOR2_X1 U4874 ( .A(n4238), .B(n4243), .Z(n4239) );
  NOR2_X1 U4875 ( .A1(n4239), .A2(n4327), .ZN(n4408) );
  INV_X1 U4876 ( .A(n4408), .ZN(n4255) );
  AND2_X1 U4877 ( .A1(n4241), .A2(n4240), .ZN(n4242) );
  XOR2_X1 U4878 ( .A(n4243), .B(n4242), .Z(n4410) );
  INV_X1 U4879 ( .A(n4273), .ZN(n4246) );
  OAI21_X1 U4880 ( .B1(n4246), .B2(n4245), .A(n4244), .ZN(n4678) );
  NOR2_X1 U4881 ( .A1(n4678), .A2(n4342), .ZN(n4253) );
  AOI22_X1 U4882 ( .A1(n4351), .A2(n4404), .B1(n4350), .B2(n4247), .ZN(n4251)
         );
  INV_X1 U4883 ( .A(n4248), .ZN(n4249) );
  AOI22_X1 U4884 ( .A1(n4365), .A2(REG2_REG_21__SCAN_IN), .B1(n4249), .B2(
        n4776), .ZN(n4250) );
  OAI211_X1 U4885 ( .C1(n4295), .C2(n4356), .A(n4251), .B(n4250), .ZN(n4252)
         );
  AOI211_X1 U4886 ( .C1(n4410), .C2(n4344), .A(n4253), .B(n4252), .ZN(n4254)
         );
  OAI21_X1 U4887 ( .B1(n4255), .B2(n4365), .A(n4254), .ZN(U3269) );
  NAND2_X1 U4888 ( .A1(n4358), .A2(n4257), .ZN(n4330) );
  NAND2_X1 U4889 ( .A1(n4330), .A2(n4258), .ZN(n4260) );
  NAND2_X1 U4890 ( .A1(n4260), .A2(n4259), .ZN(n4319) );
  NAND2_X1 U4891 ( .A1(n4317), .A2(n4262), .ZN(n4297) );
  NAND2_X1 U4892 ( .A1(n4297), .A2(n4263), .ZN(n4265) );
  NAND2_X1 U4893 ( .A1(n4265), .A2(n4264), .ZN(n4267) );
  INV_X1 U4894 ( .A(n4271), .ZN(n4266) );
  XNOR2_X1 U4895 ( .A(n4267), .B(n4266), .ZN(n4413) );
  INV_X1 U4896 ( .A(n4413), .ZN(n4282) );
  INV_X1 U4897 ( .A(n4269), .ZN(n4270) );
  NAND2_X1 U4898 ( .A1(n4268), .A2(n4270), .ZN(n4272) );
  XNOR2_X1 U4899 ( .A(n4272), .B(n4271), .ZN(n4420) );
  OAI21_X1 U4900 ( .B1(n4299), .B2(n4277), .A(n4273), .ZN(n4682) );
  NOR2_X1 U4901 ( .A1(n4682), .A2(n4342), .ZN(n4279) );
  AOI22_X1 U4902 ( .A1(n4340), .A2(n4416), .B1(n4350), .B2(n4414), .ZN(n4276)
         );
  AOI22_X1 U4903 ( .A1(n4365), .A2(REG2_REG_20__SCAN_IN), .B1(n4274), .B2(
        n4776), .ZN(n4275) );
  OAI211_X1 U4904 ( .C1(n4277), .C2(n4336), .A(n4276), .B(n4275), .ZN(n4278)
         );
  AOI211_X1 U4905 ( .C1(n4420), .C2(n4280), .A(n4279), .B(n4278), .ZN(n4281)
         );
  OAI21_X1 U4906 ( .B1(n4282), .B2(n4361), .A(n4281), .ZN(U3270) );
  INV_X1 U4907 ( .A(n4283), .ZN(n4285) );
  OAI21_X1 U4908 ( .B1(n4326), .B2(n4285), .A(n4284), .ZN(n4307) );
  INV_X1 U4909 ( .A(n4286), .ZN(n4288) );
  OAI21_X1 U4910 ( .B1(n4307), .B2(n4288), .A(n4287), .ZN(n4289) );
  XOR2_X1 U4911 ( .A(n4296), .B(n4289), .Z(n4290) );
  NAND2_X1 U4912 ( .A1(n4290), .A2(n4465), .ZN(n4294) );
  AOI22_X1 U4913 ( .A1(n4292), .A2(n4486), .B1(n4458), .B2(n4291), .ZN(n4293)
         );
  OAI211_X1 U4914 ( .C1(n4295), .C2(n4462), .A(n4294), .B(n4293), .ZN(n4425)
         );
  INV_X1 U4915 ( .A(n4425), .ZN(n4306) );
  XOR2_X1 U4916 ( .A(n4297), .B(n4296), .Z(n4426) );
  INV_X1 U4917 ( .A(n4299), .ZN(n4300) );
  OAI21_X1 U4918 ( .B1(n4298), .B2(n4301), .A(n4300), .ZN(n4685) );
  AOI22_X1 U4919 ( .A1(n4365), .A2(REG2_REG_19__SCAN_IN), .B1(n4302), .B2(
        n4776), .ZN(n4303) );
  OAI21_X1 U4920 ( .B1(n4685), .B2(n4342), .A(n4303), .ZN(n4304) );
  AOI21_X1 U4921 ( .B1(n4426), .B2(n4344), .A(n4304), .ZN(n4305) );
  OAI21_X1 U4922 ( .B1(n4306), .B2(n4365), .A(n4305), .ZN(U3271) );
  XNOR2_X1 U4923 ( .A(n4307), .B(n4320), .ZN(n4312) );
  AOI22_X1 U4924 ( .A1(n4441), .A2(n4486), .B1(n4308), .B2(n4458), .ZN(n4309)
         );
  OAI21_X1 U4925 ( .B1(n4310), .B2(n4462), .A(n4309), .ZN(n4311) );
  AOI21_X1 U4926 ( .B1(n4312), .B2(n4465), .A(n4311), .ZN(n4429) );
  NOR2_X1 U4927 ( .A1(n4349), .A2(n4313), .ZN(n4331) );
  INV_X1 U4928 ( .A(n4298), .ZN(n4314) );
  OAI211_X1 U4929 ( .C1(n4331), .C2(n4315), .A(n4314), .B(n4640), .ZN(n4428)
         );
  INV_X1 U4930 ( .A(n4428), .ZN(n4324) );
  OAI22_X1 U4931 ( .A1(n4334), .A2(n2422), .B1(n4316), .B2(n4792), .ZN(n4322)
         );
  INV_X1 U4932 ( .A(n4317), .ZN(n4318) );
  AOI21_X1 U4933 ( .B1(n4320), .B2(n4319), .A(n4318), .ZN(n4430) );
  NOR2_X1 U4934 ( .A1(n4430), .A2(n4361), .ZN(n4321) );
  AOI211_X1 U4935 ( .C1(n4324), .C2(n4323), .A(n4322), .B(n4321), .ZN(n4325)
         );
  OAI21_X1 U4936 ( .B1(n4365), .B2(n4429), .A(n4325), .ZN(U3272) );
  XOR2_X1 U4937 ( .A(n4329), .B(n4326), .Z(n4328) );
  NOR2_X1 U4938 ( .A1(n4328), .A2(n4327), .ZN(n4435) );
  INV_X1 U4939 ( .A(n4435), .ZN(n4346) );
  XOR2_X1 U4940 ( .A(n4330), .B(n4329), .Z(n4437) );
  INV_X1 U4941 ( .A(n4331), .ZN(n4332) );
  OAI21_X1 U4942 ( .B1(n2232), .B2(n4335), .A(n4332), .ZN(n4690) );
  OAI22_X1 U4943 ( .A1(n4334), .A2(n2420), .B1(n4333), .B2(n4792), .ZN(n4339)
         );
  OAI22_X1 U4944 ( .A1(n4434), .A2(n4337), .B1(n4336), .B2(n4335), .ZN(n4338)
         );
  AOI211_X1 U4945 ( .C1(n4340), .C2(n4432), .A(n4339), .B(n4338), .ZN(n4341)
         );
  OAI21_X1 U4946 ( .B1(n4690), .B2(n4342), .A(n4341), .ZN(n4343) );
  AOI21_X1 U4947 ( .B1(n4437), .B2(n4344), .A(n4343), .ZN(n4345) );
  OAI21_X1 U4948 ( .B1(n4346), .B2(n4365), .A(n4345), .ZN(U3273) );
  OAI211_X1 U4949 ( .C1(n4348), .C2(n4357), .A(n4347), .B(n4465), .ZN(n4447)
         );
  AOI21_X1 U4950 ( .B1(n4352), .B2(n4349), .A(n2232), .ZN(n4445) );
  AOI22_X1 U4951 ( .A1(n4352), .A2(n4351), .B1(n4350), .B2(n4441), .ZN(n4355)
         );
  AOI22_X1 U4952 ( .A1(n4365), .A2(REG2_REG_16__SCAN_IN), .B1(n4353), .B2(
        n4776), .ZN(n4354) );
  OAI211_X1 U4953 ( .C1(n4463), .C2(n4356), .A(n4355), .B(n4354), .ZN(n4363)
         );
  INV_X1 U4954 ( .A(n4357), .ZN(n4359) );
  OAI21_X1 U4955 ( .B1(n4360), .B2(n4359), .A(n4358), .ZN(n4448) );
  NOR2_X1 U4956 ( .A1(n4448), .A2(n4361), .ZN(n4362) );
  AOI211_X1 U4957 ( .C1(n4445), .C2(n4779), .A(n4363), .B(n4362), .ZN(n4364)
         );
  OAI21_X1 U4958 ( .B1(n4365), .B2(n4447), .A(n4364), .ZN(U3274) );
  NAND2_X1 U4959 ( .A1(n4651), .A2(n4366), .ZN(n4368) );
  NAND2_X1 U4960 ( .A1(n4825), .A2(REG1_REG_30__SCAN_IN), .ZN(n4367) );
  OAI211_X1 U4961 ( .C1(n4654), .C2(n4825), .A(n4368), .B(n4367), .ZN(U3548)
         );
  MUX2_X1 U4962 ( .A(n4370), .B(n4369), .S(n4825), .Z(n4371) );
  OAI21_X1 U4963 ( .B1(n4484), .B2(n4372), .A(n4371), .ZN(U3545) );
  AOI21_X1 U4964 ( .B1(n4374), .B2(n4482), .A(n4373), .ZN(n4655) );
  MUX2_X1 U4965 ( .A(n4375), .B(n4655), .S(n4828), .Z(n4376) );
  OAI21_X1 U4966 ( .B1(n4484), .B2(n4658), .A(n4376), .ZN(U3544) );
  AOI22_X1 U4967 ( .A1(n4378), .A2(n4486), .B1(n4458), .B2(n4377), .ZN(n4379)
         );
  OAI211_X1 U4968 ( .C1(n4381), .C2(n4462), .A(n4380), .B(n4379), .ZN(n4382)
         );
  AOI21_X1 U4969 ( .B1(n4383), .B2(n4482), .A(n4382), .ZN(n4660) );
  MUX2_X1 U4970 ( .A(n4660), .B(n4384), .S(n4825), .Z(n4385) );
  OAI21_X1 U4971 ( .B1(n4484), .B2(n4662), .A(n4385), .ZN(U3543) );
  AOI22_X1 U4972 ( .A1(n4387), .A2(n4475), .B1(n4386), .B2(n4458), .ZN(n4388)
         );
  OAI211_X1 U4973 ( .C1(n4391), .C2(n4390), .A(n4389), .B(n4388), .ZN(n4392)
         );
  AOI21_X1 U4974 ( .B1(n4393), .B2(n4482), .A(n4392), .ZN(n4663) );
  MUX2_X1 U4975 ( .A(n4565), .B(n4663), .S(n4828), .Z(n4394) );
  OAI21_X1 U4976 ( .B1(n4484), .B2(n4666), .A(n4394), .ZN(U3542) );
  AOI21_X1 U4977 ( .B1(n4396), .B2(n4482), .A(n4395), .ZN(n4667) );
  MUX2_X1 U4978 ( .A(n4397), .B(n4667), .S(n4828), .Z(n4398) );
  OAI21_X1 U4979 ( .B1(n4484), .B2(n4670), .A(n4398), .ZN(U3541) );
  NAND2_X1 U4980 ( .A1(n4399), .A2(n4482), .ZN(n4400) );
  AND2_X1 U4981 ( .A1(n4401), .A2(n4400), .ZN(n4671) );
  MUX2_X1 U4982 ( .A(n4402), .B(n4671), .S(n4828), .Z(n4403) );
  OAI21_X1 U4983 ( .B1(n4484), .B2(n4674), .A(n4403), .ZN(U3540) );
  AOI22_X1 U4984 ( .A1(n4405), .A2(n4486), .B1(n4404), .B2(n4458), .ZN(n4406)
         );
  OAI21_X1 U4985 ( .B1(n4407), .B2(n4462), .A(n4406), .ZN(n4409) );
  AOI211_X1 U4986 ( .C1(n4482), .C2(n4410), .A(n4409), .B(n4408), .ZN(n4675)
         );
  MUX2_X1 U4987 ( .A(n4411), .B(n4675), .S(n4828), .Z(n4412) );
  OAI21_X1 U4988 ( .B1(n4484), .B2(n4678), .A(n4412), .ZN(U3539) );
  NAND2_X1 U4989 ( .A1(n4413), .A2(n4482), .ZN(n4422) );
  NAND2_X1 U4990 ( .A1(n4414), .A2(n4475), .ZN(n4418) );
  AOI22_X1 U4991 ( .A1(n4416), .A2(n4486), .B1(n4415), .B2(n4458), .ZN(n4417)
         );
  NAND2_X1 U4992 ( .A1(n4418), .A2(n4417), .ZN(n4419) );
  AOI21_X1 U4993 ( .B1(n4420), .B2(n4465), .A(n4419), .ZN(n4421) );
  NAND2_X1 U4994 ( .A1(n4422), .A2(n4421), .ZN(n4679) );
  MUX2_X1 U4995 ( .A(REG1_REG_20__SCAN_IN), .B(n4679), .S(n4828), .Z(n4423) );
  INV_X1 U4996 ( .A(n4423), .ZN(n4424) );
  OAI21_X1 U4997 ( .B1(n4484), .B2(n4682), .A(n4424), .ZN(U3538) );
  AOI21_X1 U4998 ( .B1(n4426), .B2(n4482), .A(n4425), .ZN(n4683) );
  MUX2_X1 U4999 ( .A(n2335), .B(n4683), .S(n4828), .Z(n4427) );
  OAI21_X1 U5000 ( .B1(n4484), .B2(n4685), .A(n4427), .ZN(U3537) );
  OAI211_X1 U5001 ( .C1(n4649), .C2(n4430), .A(n4429), .B(n4428), .ZN(n4686)
         );
  MUX2_X1 U5002 ( .A(REG1_REG_18__SCAN_IN), .B(n4686), .S(n4828), .Z(U3536) );
  INV_X1 U5003 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4438) );
  AOI22_X1 U5004 ( .A1(n4432), .A2(n4486), .B1(n4458), .B2(n4431), .ZN(n4433)
         );
  OAI21_X1 U5005 ( .B1(n4434), .B2(n4462), .A(n4433), .ZN(n4436) );
  AOI211_X1 U5006 ( .C1(n4437), .C2(n4482), .A(n4436), .B(n4435), .ZN(n4687)
         );
  MUX2_X1 U5007 ( .A(n4438), .B(n4687), .S(n4828), .Z(n4439) );
  OAI21_X1 U5008 ( .B1(n4484), .B2(n4690), .A(n4439), .ZN(U3535) );
  AOI22_X1 U5009 ( .A1(n4441), .A2(n4475), .B1(n4486), .B2(n4440), .ZN(n4442)
         );
  OAI21_X1 U5010 ( .B1(n4443), .B2(n4477), .A(n4442), .ZN(n4444) );
  AOI21_X1 U5011 ( .B1(n4445), .B2(n4640), .A(n4444), .ZN(n4446) );
  OAI211_X1 U5012 ( .C1(n4649), .C2(n4448), .A(n4447), .B(n4446), .ZN(n4691)
         );
  MUX2_X1 U5013 ( .A(n4691), .B(REG1_REG_16__SCAN_IN), .S(n4825), .Z(U3534) );
  AOI22_X1 U5014 ( .A1(n4450), .A2(n4486), .B1(n4458), .B2(n4449), .ZN(n4451)
         );
  OAI21_X1 U5015 ( .B1(n4452), .B2(n4462), .A(n4451), .ZN(n4454) );
  AOI211_X1 U5016 ( .C1(n4482), .C2(n4455), .A(n4454), .B(n4453), .ZN(n4692)
         );
  MUX2_X1 U5017 ( .A(n2314), .B(n4692), .S(n4828), .Z(n4456) );
  OAI21_X1 U5018 ( .B1(n4484), .B2(n4695), .A(n4456), .ZN(U3533) );
  INV_X1 U5019 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4467) );
  NAND2_X1 U5020 ( .A1(n4457), .A2(n4482), .ZN(n4461) );
  AOI22_X1 U5021 ( .A1(n4474), .A2(n4486), .B1(n4459), .B2(n4458), .ZN(n4460)
         );
  OAI211_X1 U5022 ( .C1(n4463), .C2(n4462), .A(n4461), .B(n4460), .ZN(n4464)
         );
  AOI21_X1 U5023 ( .B1(n4466), .B2(n4465), .A(n4464), .ZN(n4696) );
  MUX2_X1 U5024 ( .A(n4467), .B(n4696), .S(n4828), .Z(n4468) );
  OAI21_X1 U5025 ( .B1(n4484), .B2(n4699), .A(n4468), .ZN(U3532) );
  AOI21_X1 U5026 ( .B1(n4482), .B2(n4470), .A(n4469), .ZN(n4700) );
  MUX2_X1 U5027 ( .A(n4471), .B(n4700), .S(n4828), .Z(n4472) );
  OAI21_X1 U5028 ( .B1(n4484), .B2(n4702), .A(n4472), .ZN(U3531) );
  INV_X1 U5029 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4499) );
  AOI22_X1 U5030 ( .A1(n4475), .A2(n4474), .B1(n4473), .B2(n4486), .ZN(n4476)
         );
  OAI21_X1 U5031 ( .B1(n4478), .B2(n4477), .A(n4476), .ZN(n4480) );
  AOI211_X1 U5032 ( .C1(n4482), .C2(n4481), .A(n4480), .B(n4479), .ZN(n4703)
         );
  MUX2_X1 U5033 ( .A(n4499), .B(n4703), .S(n4828), .Z(n4483) );
  OAI21_X1 U5034 ( .B1(n4484), .B2(n4707), .A(n4483), .ZN(U3530) );
  AOI22_X1 U5035 ( .A1(n4487), .A2(n4640), .B1(n4486), .B2(n4485), .ZN(n4488)
         );
  OAI211_X1 U5036 ( .C1(n4490), .C2(n4644), .A(n4489), .B(n4488), .ZN(n4708)
         );
  MUX2_X1 U5037 ( .A(REG1_REG_11__SCAN_IN), .B(n4708), .S(n4828), .Z(n4638) );
  NAND3_X1 U5038 ( .A1(REG3_REG_11__SCAN_IN), .A2(DATAI_30_), .A3(
        REG2_REG_31__SCAN_IN), .ZN(n4491) );
  NOR4_X1 U5039 ( .A1(n4492), .A2(IR_REG_1__SCAN_IN), .A3(IR_REG_4__SCAN_IN), 
        .A4(n4491), .ZN(n4493) );
  NAND3_X1 U5040 ( .A1(n4493), .A2(DATAO_REG_9__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .ZN(n4495) );
  NAND4_X1 U5041 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        REG0_REG_6__SCAN_IN), .A4(DATAO_REG_25__SCAN_IN), .ZN(n4494) );
  NOR2_X1 U5042 ( .A1(n4495), .A2(n4494), .ZN(n4505) );
  NOR4_X1 U5043 ( .A1(n4497), .A2(n4496), .A3(IR_REG_8__SCAN_IN), .A4(
        REG3_REG_23__SCAN_IN), .ZN(n4504) );
  NOR4_X1 U5044 ( .A1(n4499), .A2(n4498), .A3(REG2_REG_3__SCAN_IN), .A4(
        DATAI_19_), .ZN(n4503) );
  NAND3_X1 U5045 ( .A1(REG3_REG_27__SCAN_IN), .A2(ADDR_REG_18__SCAN_IN), .A3(
        DATAO_REG_26__SCAN_IN), .ZN(n4501) );
  INV_X1 U5046 ( .A(DATAI_21_), .ZN(n4576) );
  NAND2_X1 U5047 ( .A1(n4576), .A2(DATAI_23_), .ZN(n4500) );
  NOR4_X1 U5048 ( .A1(n4501), .A2(n4500), .A3(DATAO_REG_21__SCAN_IN), .A4(
        DATAO_REG_30__SCAN_IN), .ZN(n4502) );
  NAND4_X1 U5049 ( .A1(n4505), .A2(n4504), .A3(n4503), .A4(n4502), .ZN(n4512)
         );
  NOR4_X1 U5050 ( .A1(REG2_REG_7__SCAN_IN), .A2(REG2_REG_5__SCAN_IN), .A3(
        ADDR_REG_1__SCAN_IN), .A4(n2383), .ZN(n4507) );
  NOR3_X1 U5051 ( .A1(REG1_REG_23__SCAN_IN), .A2(REG0_REG_19__SCAN_IN), .A3(
        REG0_REG_13__SCAN_IN), .ZN(n4506) );
  NAND4_X1 U5052 ( .A1(n4508), .A2(DATAI_13_), .A3(n4507), .A4(n4506), .ZN(
        n4511) );
  NAND4_X1 U5053 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        DATAO_REG_3__SCAN_IN), .A4(n4623), .ZN(n4510) );
  INV_X1 U5054 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n4564) );
  NAND4_X1 U5055 ( .A1(REG0_REG_10__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        n4565), .A4(n4564), .ZN(n4509) );
  NOR4_X1 U5056 ( .A1(n4512), .A2(n4511), .A3(n4510), .A4(n4509), .ZN(n4518)
         );
  NAND4_X1 U5057 ( .A1(REG2_REG_6__SCAN_IN), .A2(REG3_REG_2__SCAN_IN), .A3(
        REG1_REG_18__SCAN_IN), .A4(n4579), .ZN(n4515) );
  NAND3_X1 U5058 ( .A1(IR_REG_31__SCAN_IN), .A2(REG2_REG_8__SCAN_IN), .A3(
        ADDR_REG_9__SCAN_IN), .ZN(n4514) );
  INV_X1 U5059 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4546) );
  NAND4_X1 U5060 ( .A1(REG3_REG_15__SCAN_IN), .A2(REG3_REG_21__SCAN_IN), .A3(
        ADDR_REG_0__SCAN_IN), .A4(n4546), .ZN(n4513) );
  NOR4_X1 U5061 ( .A1(ADDR_REG_11__SCAN_IN), .A2(n4515), .A3(n4514), .A4(n4513), .ZN(n4517) );
  INV_X1 U5062 ( .A(DATAI_10_), .ZN(n4573) );
  NOR4_X1 U5063 ( .A1(DATAI_15_), .A2(DATAO_REG_15__SCAN_IN), .A3(n4610), .A4(
        n4573), .ZN(n4516) );
  AND3_X1 U5064 ( .A1(n4518), .A2(n4517), .A3(n4516), .ZN(n4519) );
  OAI21_X1 U5065 ( .B1(n4519), .B2(keyinput31), .A(n4615), .ZN(n4636) );
  INV_X1 U5066 ( .A(DATAI_30_), .ZN(n4522) );
  AOI22_X1 U5067 ( .A1(n4522), .A2(keyinput55), .B1(n4521), .B2(keyinput43), 
        .ZN(n4520) );
  OAI221_X1 U5068 ( .B1(n4522), .B2(keyinput55), .C1(n4521), .C2(keyinput43), 
        .A(n4520), .ZN(n4532) );
  INV_X1 U5069 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4525) );
  INV_X1 U5070 ( .A(REG2_REG_3__SCAN_IN), .ZN(n4524) );
  AOI22_X1 U5071 ( .A1(n4525), .A2(keyinput11), .B1(n4524), .B2(keyinput18), 
        .ZN(n4523) );
  OAI221_X1 U5072 ( .B1(n4525), .B2(keyinput11), .C1(n4524), .C2(keyinput18), 
        .A(n4523), .ZN(n4531) );
  INV_X1 U5073 ( .A(ADDR_REG_1__SCAN_IN), .ZN(n4527) );
  AOI22_X1 U5074 ( .A1(n4527), .A2(keyinput8), .B1(n2383), .B2(keyinput39), 
        .ZN(n4526) );
  OAI221_X1 U5075 ( .B1(n4527), .B2(keyinput8), .C1(n2383), .C2(keyinput39), 
        .A(n4526), .ZN(n4530) );
  AOI22_X1 U5076 ( .A1(n2392), .A2(keyinput35), .B1(n2397), .B2(keyinput63), 
        .ZN(n4528) );
  OAI221_X1 U5077 ( .B1(n2392), .B2(keyinput35), .C1(n2397), .C2(keyinput63), 
        .A(n4528), .ZN(n4529) );
  NOR4_X1 U5078 ( .A1(n4532), .A2(n4531), .A3(n4530), .A4(n4529), .ZN(n4635)
         );
  INV_X1 U5079 ( .A(D_REG_6__SCAN_IN), .ZN(n4801) );
  INV_X1 U5080 ( .A(D_REG_5__SCAN_IN), .ZN(n4802) );
  AOI22_X1 U5081 ( .A1(n4801), .A2(keyinput30), .B1(keyinput22), .B2(n4802), 
        .ZN(n4533) );
  OAI221_X1 U5082 ( .B1(n4801), .B2(keyinput30), .C1(n4802), .C2(keyinput22), 
        .A(n4533), .ZN(n4543) );
  INV_X1 U5083 ( .A(DATAI_23_), .ZN(n4806) );
  AOI22_X1 U5084 ( .A1(n4806), .A2(keyinput26), .B1(n4535), .B2(keyinput29), 
        .ZN(n4534) );
  OAI221_X1 U5085 ( .B1(n4806), .B2(keyinput26), .C1(n4535), .C2(keyinput29), 
        .A(n4534), .ZN(n4542) );
  INV_X1 U5086 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4538) );
  AOI22_X1 U5087 ( .A1(n4538), .A2(keyinput40), .B1(keyinput32), .B2(n4537), 
        .ZN(n4536) );
  OAI221_X1 U5088 ( .B1(n4538), .B2(keyinput40), .C1(n4537), .C2(keyinput32), 
        .A(n4536), .ZN(n4541) );
  INV_X1 U5089 ( .A(D_REG_31__SCAN_IN), .ZN(n4793) );
  INV_X1 U5090 ( .A(D_REG_11__SCAN_IN), .ZN(n4799) );
  AOI22_X1 U5091 ( .A1(n4793), .A2(keyinput24), .B1(keyinput41), .B2(n4799), 
        .ZN(n4539) );
  OAI221_X1 U5092 ( .B1(n4793), .B2(keyinput24), .C1(n4799), .C2(keyinput41), 
        .A(n4539), .ZN(n4540) );
  NOR4_X1 U5093 ( .A1(n4543), .A2(n4542), .A3(n4541), .A4(n4540), .ZN(n4633)
         );
  INV_X1 U5094 ( .A(D_REG_14__SCAN_IN), .ZN(n4798) );
  AOI22_X1 U5095 ( .A1(n2629), .A2(keyinput28), .B1(n4798), .B2(keyinput48), 
        .ZN(n4544) );
  OAI221_X1 U5096 ( .B1(n2629), .B2(keyinput28), .C1(n4798), .C2(keyinput48), 
        .A(n4544), .ZN(n4557) );
  AOI22_X1 U5097 ( .A1(n4547), .A2(keyinput44), .B1(keyinput20), .B2(n4546), 
        .ZN(n4545) );
  OAI221_X1 U5098 ( .B1(n4547), .B2(keyinput44), .C1(n4546), .C2(keyinput20), 
        .A(n4545), .ZN(n4556) );
  INV_X1 U5099 ( .A(ADDR_REG_18__SCAN_IN), .ZN(n4550) );
  AOI22_X1 U5100 ( .A1(n4550), .A2(keyinput42), .B1(keyinput45), .B2(n4549), 
        .ZN(n4548) );
  OAI221_X1 U5101 ( .B1(n4550), .B2(keyinput42), .C1(n4549), .C2(keyinput45), 
        .A(n4548), .ZN(n4555) );
  INV_X1 U5102 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n4553) );
  AOI22_X1 U5103 ( .A1(n4553), .A2(keyinput50), .B1(keyinput53), .B2(n4552), 
        .ZN(n4551) );
  OAI221_X1 U5104 ( .B1(n4553), .B2(keyinput50), .C1(n4552), .C2(keyinput53), 
        .A(n4551), .ZN(n4554) );
  NOR4_X1 U5105 ( .A1(n4557), .A2(n4556), .A3(n4555), .A4(n4554), .ZN(n4632)
         );
  INV_X1 U5106 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4560) );
  AOI22_X1 U5107 ( .A1(n4560), .A2(keyinput17), .B1(keyinput10), .B2(n4559), 
        .ZN(n4558) );
  OAI221_X1 U5108 ( .B1(n4560), .B2(keyinput17), .C1(n4559), .C2(keyinput10), 
        .A(n4558), .ZN(n4571) );
  INV_X1 U5109 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4562) );
  AOI22_X1 U5110 ( .A1(n4562), .A2(keyinput51), .B1(n4397), .B2(keyinput59), 
        .ZN(n4561) );
  OAI221_X1 U5111 ( .B1(n4562), .B2(keyinput51), .C1(n4397), .C2(keyinput59), 
        .A(n4561), .ZN(n4570) );
  AOI22_X1 U5112 ( .A1(n4565), .A2(keyinput1), .B1(keyinput21), .B2(n4564), 
        .ZN(n4563) );
  OAI221_X1 U5113 ( .B1(n4565), .B2(keyinput1), .C1(n4564), .C2(keyinput21), 
        .A(n4563), .ZN(n4569) );
  INV_X1 U5114 ( .A(D_REG_17__SCAN_IN), .ZN(n4796) );
  AOI22_X1 U5115 ( .A1(n4567), .A2(keyinput16), .B1(n4796), .B2(keyinput12), 
        .ZN(n4566) );
  OAI221_X1 U5116 ( .B1(n4567), .B2(keyinput16), .C1(n4796), .C2(keyinput12), 
        .A(n4566), .ZN(n4568) );
  NOR4_X1 U5117 ( .A1(n4571), .A2(n4570), .A3(n4569), .A4(n4568), .ZN(n4631)
         );
  AOI22_X1 U5118 ( .A1(n4574), .A2(keyinput47), .B1(n4573), .B2(keyinput27), 
        .ZN(n4572) );
  OAI221_X1 U5119 ( .B1(n4574), .B2(keyinput47), .C1(n4573), .C2(keyinput27), 
        .A(n4572), .ZN(n4583) );
  INV_X1 U5120 ( .A(DATAI_19_), .ZN(n4577) );
  AOI22_X1 U5121 ( .A1(n4577), .A2(keyinput61), .B1(n4576), .B2(keyinput60), 
        .ZN(n4575) );
  OAI221_X1 U5122 ( .B1(n4577), .B2(keyinput61), .C1(n4576), .C2(keyinput60), 
        .A(n4575), .ZN(n4582) );
  AOI22_X1 U5123 ( .A1(n4580), .A2(keyinput38), .B1(n4579), .B2(keyinput62), 
        .ZN(n4578) );
  OAI221_X1 U5124 ( .B1(n4580), .B2(keyinput38), .C1(n4579), .C2(keyinput62), 
        .A(n4578), .ZN(n4581) );
  NOR3_X1 U5125 ( .A1(n4583), .A2(n4582), .A3(n4581), .ZN(n4629) );
  INV_X1 U5126 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4586) );
  INV_X1 U5127 ( .A(ADDR_REG_9__SCAN_IN), .ZN(n4585) );
  AOI22_X1 U5128 ( .A1(n4586), .A2(keyinput33), .B1(keyinput36), .B2(n4585), 
        .ZN(n4584) );
  OAI221_X1 U5129 ( .B1(n4586), .B2(keyinput33), .C1(n4585), .C2(keyinput36), 
        .A(n4584), .ZN(n4587) );
  INV_X1 U5130 ( .A(n4587), .ZN(n4607) );
  XNOR2_X1 U5131 ( .A(REG3_REG_2__SCAN_IN), .B(keyinput25), .ZN(n4591) );
  XNOR2_X1 U5132 ( .A(IR_REG_4__SCAN_IN), .B(keyinput56), .ZN(n4590) );
  XNOR2_X1 U5133 ( .A(IR_REG_13__SCAN_IN), .B(keyinput57), .ZN(n4589) );
  XNOR2_X1 U5134 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput15), .ZN(n4588) );
  NAND4_X1 U5135 ( .A1(n4591), .A2(n4590), .A3(n4589), .A4(n4588), .ZN(n4597)
         );
  XNOR2_X1 U5136 ( .A(REG1_REG_12__SCAN_IN), .B(keyinput3), .ZN(n4595) );
  XNOR2_X1 U5137 ( .A(IR_REG_8__SCAN_IN), .B(keyinput7), .ZN(n4594) );
  XNOR2_X1 U5138 ( .A(IR_REG_1__SCAN_IN), .B(keyinput0), .ZN(n4593) );
  XNOR2_X1 U5139 ( .A(IR_REG_17__SCAN_IN), .B(keyinput2), .ZN(n4592) );
  NAND4_X1 U5140 ( .A1(n4595), .A2(n4594), .A3(n4593), .A4(n4592), .ZN(n4596)
         );
  NOR2_X1 U5141 ( .A1(n4597), .A2(n4596), .ZN(n4606) );
  INV_X1 U5142 ( .A(REG2_REG_6__SCAN_IN), .ZN(n4598) );
  XNOR2_X1 U5143 ( .A(keyinput49), .B(n4598), .ZN(n4600) );
  XNOR2_X1 U5144 ( .A(keyinput34), .B(n4093), .ZN(n4599) );
  NOR2_X1 U5145 ( .A1(n4600), .A2(n4599), .ZN(n4605) );
  INV_X1 U5146 ( .A(D_REG_28__SCAN_IN), .ZN(n4794) );
  XNOR2_X1 U5147 ( .A(keyinput5), .B(n4794), .ZN(n4603) );
  XNOR2_X1 U5148 ( .A(keyinput6), .B(n4601), .ZN(n4602) );
  NOR2_X1 U5149 ( .A1(n4603), .A2(n4602), .ZN(n4604) );
  AND4_X1 U5150 ( .A1(n4607), .A2(n4606), .A3(n4605), .A4(n4604), .ZN(n4628)
         );
  INV_X1 U5151 ( .A(D_REG_16__SCAN_IN), .ZN(n4797) );
  INV_X1 U5152 ( .A(D_REG_25__SCAN_IN), .ZN(n4795) );
  AOI22_X1 U5153 ( .A1(n4797), .A2(keyinput14), .B1(keyinput13), .B2(n4795), 
        .ZN(n4608) );
  OAI221_X1 U5154 ( .B1(n4797), .B2(keyinput14), .C1(n4795), .C2(keyinput13), 
        .A(n4608), .ZN(n4618) );
  INV_X1 U5155 ( .A(DATAI_15_), .ZN(n4811) );
  AOI22_X1 U5156 ( .A1(n4610), .A2(keyinput19), .B1(keyinput23), .B2(n4811), 
        .ZN(n4609) );
  OAI221_X1 U5157 ( .B1(n4610), .B2(keyinput19), .C1(n4811), .C2(keyinput23), 
        .A(n4609), .ZN(n4617) );
  XNOR2_X1 U5158 ( .A(REG3_REG_27__SCAN_IN), .B(keyinput46), .ZN(n4612) );
  XNOR2_X1 U5159 ( .A(IR_REG_21__SCAN_IN), .B(keyinput58), .ZN(n4611) );
  AND2_X1 U5160 ( .A1(n4612), .A2(n4611), .ZN(n4614) );
  XNOR2_X1 U5161 ( .A(IR_REG_31__SCAN_IN), .B(keyinput37), .ZN(n4613) );
  OAI211_X1 U5162 ( .C1(n4615), .C2(keyinput31), .A(n4614), .B(n4613), .ZN(
        n4616) );
  NOR3_X1 U5163 ( .A1(n4618), .A2(n4617), .A3(n4616), .ZN(n4627) );
  INV_X1 U5164 ( .A(D_REG_7__SCAN_IN), .ZN(n4800) );
  AOI22_X1 U5165 ( .A1(n4800), .A2(keyinput52), .B1(keyinput54), .B2(n4620), 
        .ZN(n4619) );
  OAI221_X1 U5166 ( .B1(n4800), .B2(keyinput52), .C1(n4620), .C2(keyinput54), 
        .A(n4619), .ZN(n4625) );
  AOI22_X1 U5167 ( .A1(n4623), .A2(keyinput9), .B1(keyinput4), .B2(n4622), 
        .ZN(n4621) );
  OAI221_X1 U5168 ( .B1(n4623), .B2(keyinput9), .C1(n4622), .C2(keyinput4), 
        .A(n4621), .ZN(n4624) );
  NOR2_X1 U5169 ( .A1(n4625), .A2(n4624), .ZN(n4626) );
  AND4_X1 U5170 ( .A1(n4629), .A2(n4628), .A3(n4627), .A4(n4626), .ZN(n4630)
         );
  AND4_X1 U5171 ( .A1(n4633), .A2(n4632), .A3(n4631), .A4(n4630), .ZN(n4634)
         );
  NAND3_X1 U5172 ( .A1(n4636), .A2(n4635), .A3(n4634), .ZN(n4637) );
  XNOR2_X1 U5173 ( .A(n4638), .B(n4637), .ZN(U3529) );
  NAND3_X1 U5174 ( .A1(n4641), .A2(n4640), .A3(n4639), .ZN(n4642) );
  OAI211_X1 U5175 ( .C1(n4645), .C2(n4644), .A(n4643), .B(n4642), .ZN(n4709)
         );
  MUX2_X1 U5176 ( .A(REG1_REG_8__SCAN_IN), .B(n4709), .S(n4828), .Z(U3526) );
  OAI211_X1 U5177 ( .C1(n4649), .C2(n4648), .A(n4647), .B(n4646), .ZN(n4710)
         );
  MUX2_X1 U5178 ( .A(REG1_REG_7__SCAN_IN), .B(n4710), .S(n4828), .Z(U3525) );
  NAND2_X1 U5179 ( .A1(n4651), .A2(n4650), .ZN(n4653) );
  NAND2_X1 U5180 ( .A1(n4822), .A2(REG0_REG_30__SCAN_IN), .ZN(n4652) );
  OAI211_X1 U5181 ( .C1(n4654), .C2(n4822), .A(n4653), .B(n4652), .ZN(U3516)
         );
  INV_X1 U5182 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4656) );
  MUX2_X1 U5183 ( .A(n4656), .B(n4655), .S(n4824), .Z(n4657) );
  OAI21_X1 U5184 ( .B1(n4658), .B2(n4706), .A(n4657), .ZN(U3512) );
  INV_X1 U5185 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4659) );
  MUX2_X1 U5186 ( .A(n4660), .B(n4659), .S(n4822), .Z(n4661) );
  OAI21_X1 U5187 ( .B1(n4662), .B2(n4706), .A(n4661), .ZN(U3511) );
  INV_X1 U5188 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4664) );
  MUX2_X1 U5189 ( .A(n4664), .B(n4663), .S(n4824), .Z(n4665) );
  OAI21_X1 U5190 ( .B1(n4666), .B2(n4706), .A(n4665), .ZN(U3510) );
  INV_X1 U5191 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4668) );
  MUX2_X1 U5192 ( .A(n4668), .B(n4667), .S(n4824), .Z(n4669) );
  OAI21_X1 U5193 ( .B1(n4670), .B2(n4706), .A(n4669), .ZN(U3509) );
  INV_X1 U5194 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4672) );
  MUX2_X1 U5195 ( .A(n4672), .B(n4671), .S(n4824), .Z(n4673) );
  OAI21_X1 U5196 ( .B1(n4674), .B2(n4706), .A(n4673), .ZN(U3508) );
  INV_X1 U5197 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4676) );
  MUX2_X1 U5198 ( .A(n4676), .B(n4675), .S(n4824), .Z(n4677) );
  OAI21_X1 U5199 ( .B1(n4678), .B2(n4706), .A(n4677), .ZN(U3507) );
  MUX2_X1 U5200 ( .A(REG0_REG_20__SCAN_IN), .B(n4679), .S(n4824), .Z(n4680) );
  INV_X1 U5201 ( .A(n4680), .ZN(n4681) );
  OAI21_X1 U5202 ( .B1(n4682), .B2(n4706), .A(n4681), .ZN(U3506) );
  MUX2_X1 U5203 ( .A(n4562), .B(n4683), .S(n4824), .Z(n4684) );
  OAI21_X1 U5204 ( .B1(n4685), .B2(n4706), .A(n4684), .ZN(U3505) );
  MUX2_X1 U5205 ( .A(REG0_REG_18__SCAN_IN), .B(n4686), .S(n4824), .Z(U3503) );
  INV_X1 U5206 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4688) );
  MUX2_X1 U5207 ( .A(n4688), .B(n4687), .S(n4824), .Z(n4689) );
  OAI21_X1 U5208 ( .B1(n4690), .B2(n4706), .A(n4689), .ZN(U3501) );
  MUX2_X1 U5209 ( .A(n4691), .B(REG0_REG_16__SCAN_IN), .S(n4822), .Z(U3499) );
  INV_X1 U5210 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4693) );
  MUX2_X1 U5211 ( .A(n4693), .B(n4692), .S(n4824), .Z(n4694) );
  OAI21_X1 U5212 ( .B1(n4695), .B2(n4706), .A(n4694), .ZN(U3497) );
  INV_X1 U5213 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4697) );
  MUX2_X1 U5214 ( .A(n4697), .B(n4696), .S(n4824), .Z(n4698) );
  OAI21_X1 U5215 ( .B1(n4699), .B2(n4706), .A(n4698), .ZN(U3495) );
  MUX2_X1 U5216 ( .A(n4560), .B(n4700), .S(n4824), .Z(n4701) );
  OAI21_X1 U5217 ( .B1(n4702), .B2(n4706), .A(n4701), .ZN(U3493) );
  INV_X1 U5218 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4704) );
  MUX2_X1 U5219 ( .A(n4704), .B(n4703), .S(n4824), .Z(n4705) );
  OAI21_X1 U5220 ( .B1(n4707), .B2(n4706), .A(n4705), .ZN(U3491) );
  MUX2_X1 U5221 ( .A(REG0_REG_11__SCAN_IN), .B(n4708), .S(n4824), .Z(U3489) );
  MUX2_X1 U5222 ( .A(REG0_REG_8__SCAN_IN), .B(n4709), .S(n4824), .Z(U3483) );
  MUX2_X1 U5223 ( .A(REG0_REG_7__SCAN_IN), .B(n4710), .S(n4824), .Z(U3481) );
  MUX2_X1 U5224 ( .A(n4711), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U5225 ( .A(n4712), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5226 ( .A(n4713), .B(DATAI_28_), .S(U3149), .Z(U3324) );
  MUX2_X1 U5227 ( .A(DATAI_22_), .B(n4714), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U5228 ( .A(n4715), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5229 ( .A(DATAI_20_), .B(n4716), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5230 ( .A(n4717), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5231 ( .A(DATAI_12_), .B(n4718), .S(STATE_REG_SCAN_IN), .Z(U3340)
         );
  MUX2_X1 U5232 ( .A(n2291), .B(DATAI_11_), .S(U3149), .Z(U3341) );
  MUX2_X1 U5233 ( .A(n4719), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U5234 ( .A(n4720), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U5235 ( .A(DATAI_8_), .B(n4721), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U5236 ( .A(n4722), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5237 ( .A(DATAI_6_), .B(n4723), .S(STATE_REG_SCAN_IN), .Z(U3346) );
  MUX2_X1 U5238 ( .A(n4724), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5239 ( .A(DATAI_4_), .B(n4725), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5240 ( .A(DATAI_3_), .B(n4726), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U5241 ( .A(n4727), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5242 ( .A(n4728), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U5243 ( .A(DATAI_0_), .B(n4729), .S(STATE_REG_SCAN_IN), .Z(U3352) );
  INV_X1 U5244 ( .A(n4730), .ZN(n4734) );
  AOI211_X1 U5245 ( .C1(n4732), .C2(n4731), .A(n2039), .B(n4762), .ZN(n4733)
         );
  AOI211_X1 U5246 ( .C1(n4765), .C2(ADDR_REG_14__SCAN_IN), .A(n4734), .B(n4733), .ZN(n4738) );
  OAI211_X1 U5247 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4736), .A(n4770), .B(n4735), .ZN(n4737) );
  OAI211_X1 U5248 ( .C1(n4775), .C2(n4739), .A(n4738), .B(n4737), .ZN(U3254)
         );
  AOI211_X1 U5249 ( .C1(n4742), .C2(n4741), .A(n4740), .B(n4762), .ZN(n4743)
         );
  AOI211_X1 U5250 ( .C1(n4765), .C2(ADDR_REG_15__SCAN_IN), .A(n4744), .B(n4743), .ZN(n4750) );
  NAND2_X1 U5251 ( .A1(n4745), .A2(n4735), .ZN(n4747) );
  NAND2_X1 U5252 ( .A1(n4748), .A2(n4747), .ZN(n4746) );
  OAI211_X1 U5253 ( .C1(n4748), .C2(n4747), .A(n4770), .B(n4746), .ZN(n4749)
         );
  OAI211_X1 U5254 ( .C1(n4775), .C2(n4812), .A(n4750), .B(n4749), .ZN(U3255)
         );
  AOI221_X1 U5255 ( .B1(n4753), .B2(n4751), .C1(n4752), .C2(n4751), .A(n4762), 
        .ZN(n4754) );
  AOI211_X1 U5256 ( .C1(n4765), .C2(ADDR_REG_16__SCAN_IN), .A(n4755), .B(n4754), .ZN(n4759) );
  OAI221_X1 U5257 ( .B1(n4756), .B2(REG1_REG_16__SCAN_IN), .C1(n4756), .C2(
        n4757), .A(n4770), .ZN(n4758) );
  OAI211_X1 U5258 ( .C1(n4775), .C2(n4810), .A(n4759), .B(n4758), .ZN(U3256)
         );
  INV_X1 U5259 ( .A(n4766), .ZN(n4767) );
  OAI211_X1 U5260 ( .C1(n4772), .C2(n4771), .A(n4770), .B(n4769), .ZN(n4773)
         );
  OAI211_X1 U5261 ( .C1(n4775), .C2(n4808), .A(n4774), .B(n4773), .ZN(U3258)
         );
  AOI22_X1 U5262 ( .A1(n4788), .A2(REG2_REG_3__SCAN_IN), .B1(n4776), .B2(n2460), .ZN(n4781) );
  AOI22_X1 U5263 ( .A1(n4779), .A2(n4778), .B1(n4777), .B2(n4784), .ZN(n4780)
         );
  OAI211_X1 U5264 ( .C1(n4788), .C2(n4782), .A(n4781), .B(n4780), .ZN(U3287)
         );
  AOI22_X1 U5265 ( .A1(n4784), .A2(n4783), .B1(REG2_REG_0__SCAN_IN), .B2(n4365), .ZN(n4791) );
  AOI21_X1 U5266 ( .B1(n4787), .B2(n4786), .A(n4785), .ZN(n4789) );
  OR2_X1 U5267 ( .A1(n4789), .A2(n4788), .ZN(n4790) );
  OAI211_X1 U5268 ( .C1(n4792), .C2(n3150), .A(n4791), .B(n4790), .ZN(U3290)
         );
  NOR2_X1 U5269 ( .A1(n4803), .A2(n4793), .ZN(U3291) );
  AND2_X1 U5270 ( .A1(D_REG_30__SCAN_IN), .A2(n4804), .ZN(U3292) );
  AND2_X1 U5271 ( .A1(D_REG_29__SCAN_IN), .A2(n4804), .ZN(U3293) );
  NOR2_X1 U5272 ( .A1(n4803), .A2(n4794), .ZN(U3294) );
  AND2_X1 U5273 ( .A1(D_REG_27__SCAN_IN), .A2(n4804), .ZN(U3295) );
  AND2_X1 U5274 ( .A1(D_REG_26__SCAN_IN), .A2(n4804), .ZN(U3296) );
  NOR2_X1 U5275 ( .A1(n4803), .A2(n4795), .ZN(U3297) );
  AND2_X1 U5276 ( .A1(D_REG_24__SCAN_IN), .A2(n4804), .ZN(U3298) );
  AND2_X1 U5277 ( .A1(D_REG_23__SCAN_IN), .A2(n4804), .ZN(U3299) );
  AND2_X1 U5278 ( .A1(D_REG_22__SCAN_IN), .A2(n4804), .ZN(U3300) );
  AND2_X1 U5279 ( .A1(D_REG_21__SCAN_IN), .A2(n4804), .ZN(U3301) );
  AND2_X1 U5280 ( .A1(D_REG_20__SCAN_IN), .A2(n4804), .ZN(U3302) );
  AND2_X1 U5281 ( .A1(D_REG_19__SCAN_IN), .A2(n4804), .ZN(U3303) );
  AND2_X1 U5282 ( .A1(D_REG_18__SCAN_IN), .A2(n4804), .ZN(U3304) );
  NOR2_X1 U5283 ( .A1(n4803), .A2(n4796), .ZN(U3305) );
  NOR2_X1 U5284 ( .A1(n4803), .A2(n4797), .ZN(U3306) );
  AND2_X1 U5285 ( .A1(D_REG_15__SCAN_IN), .A2(n4804), .ZN(U3307) );
  NOR2_X1 U5286 ( .A1(n4803), .A2(n4798), .ZN(U3308) );
  AND2_X1 U5287 ( .A1(D_REG_13__SCAN_IN), .A2(n4804), .ZN(U3309) );
  AND2_X1 U5288 ( .A1(D_REG_12__SCAN_IN), .A2(n4804), .ZN(U3310) );
  NOR2_X1 U5289 ( .A1(n4803), .A2(n4799), .ZN(U3311) );
  AND2_X1 U5290 ( .A1(D_REG_10__SCAN_IN), .A2(n4804), .ZN(U3312) );
  AND2_X1 U5291 ( .A1(D_REG_9__SCAN_IN), .A2(n4804), .ZN(U3313) );
  AND2_X1 U5292 ( .A1(D_REG_8__SCAN_IN), .A2(n4804), .ZN(U3314) );
  NOR2_X1 U5293 ( .A1(n4803), .A2(n4800), .ZN(U3315) );
  NOR2_X1 U5294 ( .A1(n4803), .A2(n4801), .ZN(U3316) );
  NOR2_X1 U5295 ( .A1(n4803), .A2(n4802), .ZN(U3317) );
  AND2_X1 U5296 ( .A1(D_REG_4__SCAN_IN), .A2(n4804), .ZN(U3318) );
  AND2_X1 U5297 ( .A1(D_REG_3__SCAN_IN), .A2(n4804), .ZN(U3319) );
  AND2_X1 U5298 ( .A1(D_REG_2__SCAN_IN), .A2(n4804), .ZN(U3320) );
  AOI21_X1 U5299 ( .B1(U3149), .B2(n4806), .A(n4805), .ZN(U3329) );
  INV_X1 U5300 ( .A(DATAI_18_), .ZN(n4807) );
  AOI22_X1 U5301 ( .A1(STATE_REG_SCAN_IN), .A2(n4808), .B1(n4807), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U5302 ( .A(DATAI_16_), .ZN(n4809) );
  AOI22_X1 U5303 ( .A1(STATE_REG_SCAN_IN), .A2(n4810), .B1(n4809), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5304 ( .A1(STATE_REG_SCAN_IN), .A2(n4812), .B1(n4811), .B2(U3149), 
        .ZN(U3337) );
  OAI22_X1 U5305 ( .A1(U3149), .A2(n4813), .B1(DATAI_14_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4814) );
  INV_X1 U5306 ( .A(n4814), .ZN(U3338) );
  INV_X1 U5307 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4815) );
  AOI22_X1 U5308 ( .A1(n4824), .A2(n4816), .B1(n4815), .B2(n4822), .ZN(U3467)
         );
  INV_X1 U5309 ( .A(n4817), .ZN(n4819) );
  AOI211_X1 U5310 ( .C1(n4821), .C2(n4820), .A(n4819), .B(n4818), .ZN(n4827)
         );
  INV_X1 U5311 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4823) );
  AOI22_X1 U5312 ( .A1(n4824), .A2(n4827), .B1(n4823), .B2(n4822), .ZN(U3475)
         );
  AOI22_X1 U5313 ( .A1(n4828), .A2(n4827), .B1(n4826), .B2(n4825), .ZN(U3522)
         );
  CLKBUF_X1 U2274 ( .A(n2015), .Z(n3013) );
  CLKBUF_X1 U2295 ( .A(n2461), .Z(n2536) );
  CLKBUF_X1 U2335 ( .A(n2440), .Z(n4711) );
  CLKBUF_X1 U2520 ( .A(n2384), .Z(n4727) );
endmodule

