

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput127, keyinput126,
         keyinput125, keyinput124, keyinput123, keyinput122, keyinput121,
         keyinput120, keyinput119, keyinput118, keyinput117, keyinput116,
         keyinput115, keyinput114, keyinput113, keyinput112, keyinput111,
         keyinput110, keyinput109, keyinput108, keyinput107, keyinput106,
         keyinput105, keyinput104, keyinput103, keyinput102, keyinput101,
         keyinput100, keyinput99, keyinput98, keyinput97, keyinput96,
         keyinput95, keyinput94, keyinput93, keyinput92, keyinput91,
         keyinput90, keyinput89, keyinput88, keyinput87, keyinput86,
         keyinput85, keyinput84, keyinput83, keyinput82, keyinput81,
         keyinput80, keyinput79, keyinput78, keyinput77, keyinput76,
         keyinput75, keyinput74, keyinput73, keyinput72, keyinput71,
         keyinput70, keyinput69, keyinput68, keyinput67, keyinput66,
         keyinput65, keyinput64, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049;

  INV_X1 U3580 ( .A(n6361), .ZN(n6347) );
  NAND2_X1 U3581 ( .A1(n5461), .A2(n5460), .ZN(n5459) );
  INV_X2 U3582 ( .A(n6434), .ZN(n3952) );
  NAND2_X1 U3583 ( .A1(n5716), .A2(n5700), .ZN(n5802) );
  CLKBUF_X2 U3585 ( .A(n3830), .Z(n3138) );
  CLKBUF_X2 U3586 ( .A(n4089), .Z(n4172) );
  CLKBUF_X2 U3587 ( .A(n3475), .Z(n4162) );
  CLKBUF_X2 U3588 ( .A(n3242), .Z(n3137) );
  CLKBUF_X1 U3589 ( .A(n3330), .Z(n4805) );
  INV_X2 U3590 ( .A(n3960), .ZN(n4683) );
  AND4_X1 U3591 ( .A1(n3280), .A2(n3279), .A3(n3278), .A4(n3277), .ZN(n3291)
         );
  AND4_X1 U3592 ( .A1(n3260), .A2(n3259), .A3(n3258), .A4(n3257), .ZN(n3271)
         );
  AND4_X1 U3593 ( .A1(n3264), .A2(n3263), .A3(n3262), .A4(n3261), .ZN(n3270)
         );
  AND2_X1 U3595 ( .A1(n3171), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5557)
         );
  AOI22_X1 U3596 ( .A1(n6835), .A2(keyinput93), .B1(n6984), .B2(keyinput108), 
        .ZN(n6834) );
  OAI221_X1 U3597 ( .B1(n6835), .B2(keyinput93), .C1(n6984), .C2(keyinput108), 
        .A(n6834), .ZN(n6836) );
  AND2_X1 U3598 ( .A1(n3176), .A2(n3177), .ZN(n4089) );
  AND2_X2 U3599 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4627) );
  NAND2_X1 U3600 ( .A1(n4931), .A2(n4004), .ZN(n4337) );
  BUF_X1 U3601 ( .A(n3299), .Z(n5493) );
  INV_X1 U3602 ( .A(n4154), .ZN(n4193) );
  NAND2_X1 U3603 ( .A1(n3563), .A2(n3562), .ZN(n4206) );
  BUF_X1 U3605 ( .A(n5291), .Z(n3146) );
  NOR2_X1 U3606 ( .A1(n5569), .A2(n5568), .ZN(n4349) );
  AND4_X1 U3607 ( .A1(n3288), .A2(n3287), .A3(n3286), .A4(n3285), .ZN(n3289)
         );
  NOR2_X1 U3608 ( .A1(n4583), .A2(n4952), .ZN(n4950) );
  CLKBUF_X3 U3610 ( .A(n4216), .Z(n4640) );
  XNOR2_X1 U3611 ( .A(n3372), .B(n3371), .ZN(n5763) );
  MUX2_X1 U3612 ( .A(n3448), .B(n3447), .S(n3446), .Z(n5379) );
  INV_X1 U3613 ( .A(n6220), .ZN(n6171) );
  INV_X1 U3614 ( .A(n6196), .ZN(n6258) );
  AOI211_X1 U3615 ( .C1(n5576), .C2(n5575), .A(n5574), .B(n5573), .ZN(n5577)
         );
  INV_X1 U3616 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4622) );
  AND2_X1 U3617 ( .A1(n4699), .A2(n3473), .ZN(n3132) );
  NAND2_X2 U3618 ( .A1(n4412), .A2(n5613), .ZN(n5853) );
  AND2_X4 U3619 ( .A1(n5557), .A2(n4627), .ZN(n4121) );
  NOR2_X4 U3620 ( .A1(n4304), .A2(n4302), .ZN(n4442) );
  AND2_X2 U3621 ( .A1(n5505), .A2(n5506), .ZN(n4304) );
  AND2_X1 U3622 ( .A1(n3176), .A2(n5551), .ZN(n3133) );
  AND2_X1 U3623 ( .A1(n3176), .A2(n5551), .ZN(n3134) );
  AND2_X1 U3624 ( .A1(n3176), .A2(n5551), .ZN(n3390) );
  AOI211_X2 U3626 ( .C1(n6336), .C2(n5856), .A(n5855), .B(n5854), .ZN(n5857)
         );
  INV_X1 U3627 ( .A(n3132), .ZN(n3135) );
  NOR2_X1 U3628 ( .A1(n5578), .A2(n5521), .ZN(n5520) );
  OAI21_X1 U3629 ( .B1(n5902), .B2(n4296), .A(n4295), .ZN(n5858) );
  INV_X1 U3630 ( .A(n5459), .ZN(n3142) );
  NAND2_X1 U3631 ( .A1(n4573), .A2(n4582), .ZN(n4583) );
  CLKBUF_X1 U3632 ( .A(n4639), .Z(n6012) );
  CLKBUF_X1 U3633 ( .A(n4614), .Z(n6014) );
  NAND2_X1 U3634 ( .A1(n3421), .A2(n4207), .ZN(n3439) );
  AND2_X1 U3635 ( .A1(n3341), .A2(n3319), .ZN(n3370) );
  OAI21_X1 U3636 ( .B1(n4602), .B2(n3309), .A(n4355), .ZN(n3310) );
  NOR2_X1 U3637 ( .A1(n3312), .A2(n3311), .ZN(n3892) );
  OR2_X2 U3638 ( .A1(n4321), .A2(n4689), .ZN(n4602) );
  AND2_X1 U3639 ( .A1(n3306), .A2(n3297), .ZN(n4364) );
  INV_X2 U3640 ( .A(n3983), .ZN(n3979) );
  NAND2_X1 U3641 ( .A1(n4213), .A2(n4662), .ZN(n4359) );
  BUF_X1 U3642 ( .A(n3304), .Z(n3365) );
  INV_X2 U3643 ( .A(n3299), .ZN(n4800) );
  INV_X2 U3644 ( .A(n4213), .ZN(n3136) );
  AND4_X1 U3645 ( .A1(n3284), .A2(n3283), .A3(n3282), .A4(n3281), .ZN(n3290)
         );
  AND4_X1 U3646 ( .A1(n3276), .A2(n3275), .A3(n3274), .A4(n3273), .ZN(n3292)
         );
  BUF_X2 U3648 ( .A(n3390), .Z(n3407) );
  BUF_X2 U3649 ( .A(n3208), .Z(n4166) );
  CLKBUF_X2 U3650 ( .A(n4121), .Z(n4173) );
  CLKBUF_X1 U3651 ( .A(n3156), .Z(n3139) );
  AND2_X2 U3652 ( .A1(n3177), .A2(n4627), .ZN(n3475) );
  AOI211_X1 U3653 ( .C1(n5566), .C2(n5575), .A(n5565), .B(n5564), .ZN(n5588)
         );
  INV_X1 U3654 ( .A(n6041), .ZN(n5772) );
  AND2_X1 U3655 ( .A1(n5642), .A2(n5641), .ZN(n6041) );
  NAND2_X1 U3656 ( .A1(n5517), .A2(n5516), .ZN(n5562) );
  NOR2_X2 U3657 ( .A1(n5850), .A2(n5930), .ZN(n5566) );
  XNOR2_X1 U3658 ( .A(n5520), .B(n4194), .ZN(n5818) );
  NAND2_X1 U3659 ( .A1(n5578), .A2(n5581), .ZN(n5603) );
  AND2_X1 U3660 ( .A1(n5889), .A2(n5890), .ZN(n5865) );
  OR2_X1 U3661 ( .A1(n4439), .A2(n4409), .ZN(n4412) );
  NAND2_X1 U3662 ( .A1(n5579), .A2(n5580), .ZN(n5578) );
  AOI21_X1 U3663 ( .B1(n5991), .B2(n5863), .A(n5862), .ZN(n5889) );
  CLKBUF_X1 U3664 ( .A(n5666), .Z(n5667) );
  AND2_X2 U3665 ( .A1(n5666), .A2(n3819), .ZN(n4411) );
  AND2_X1 U3666 ( .A1(n5861), .A2(n5860), .ZN(n5991) );
  CLKBUF_X1 U3668 ( .A(n5902), .Z(n6061) );
  INV_X1 U3669 ( .A(n5799), .ZN(n5786) );
  CLKBUF_X1 U3670 ( .A(n5903), .Z(n5916) );
  XNOR2_X1 U3671 ( .A(n4354), .B(n4353), .ZN(n5513) );
  CLKBUF_X1 U3672 ( .A(n5315), .Z(n5330) );
  INV_X1 U3673 ( .A(n5182), .ZN(n5280) );
  NAND2_X2 U3674 ( .A1(n4206), .A2(n4208), .ZN(n5880) );
  AND2_X1 U3675 ( .A1(n5754), .A2(n3959), .ZN(n6220) );
  AOI21_X1 U3676 ( .B1(n4257), .B2(n3695), .A(n3559), .ZN(n4952) );
  INV_X1 U3677 ( .A(n6090), .ZN(n6414) );
  CLKBUF_X1 U3678 ( .A(n4638), .Z(n4730) );
  NAND2_X1 U3679 ( .A1(n4539), .A2(n3461), .ZN(n4576) );
  OR2_X1 U3680 ( .A1(n4375), .A2(n4697), .ZN(n5147) );
  NAND2_X1 U3681 ( .A1(n4541), .A2(n4540), .ZN(n4539) );
  NAND2_X1 U3682 ( .A1(n5438), .A2(n5437), .ZN(n5454) );
  NAND2_X1 U3683 ( .A1(n4380), .A2(n6576), .ZN(n6415) );
  NAND2_X1 U3684 ( .A1(n4326), .A2(n4325), .ZN(n4380) );
  NAND2_X1 U3685 ( .A1(n3445), .A2(n3444), .ZN(n4541) );
  AND2_X1 U3686 ( .A1(n3430), .A2(n3429), .ZN(n3434) );
  CLKBUF_X1 U3687 ( .A(n4585), .Z(n6439) );
  XNOR2_X1 U3688 ( .A(n4631), .B(n4897), .ZN(n4585) );
  NOR2_X1 U3689 ( .A1(n5344), .A2(n5343), .ZN(n4007) );
  NAND2_X1 U3690 ( .A1(n3467), .A2(n3350), .ZN(n4614) );
  NAND2_X1 U3691 ( .A1(n3384), .A2(n3385), .ZN(n3388) );
  NAND2_X1 U3692 ( .A1(n3325), .A2(n3324), .ZN(n3384) );
  CLKBUF_X1 U3693 ( .A(n3892), .Z(n4461) );
  CLKBUF_X1 U3694 ( .A(n4321), .Z(n4586) );
  OR2_X1 U3695 ( .A1(n3296), .A2(n3249), .ZN(n4315) );
  OR2_X1 U3696 ( .A1(n3332), .A2(n3331), .ZN(n4617) );
  INV_X1 U3697 ( .A(n3972), .ZN(n4010) );
  NOR2_X1 U3698 ( .A1(n4359), .A2(n3305), .ZN(n3307) );
  INV_X1 U3699 ( .A(n3704), .ZN(n4196) );
  INV_X1 U3700 ( .A(n4705), .ZN(n5815) );
  AND2_X2 U3701 ( .A1(n4683), .A2(n3154), .ZN(n4456) );
  AND4_X2 U3702 ( .A1(n3161), .A2(n3237), .A3(n3236), .A4(n3235), .ZN(n4662)
         );
  INV_X1 U3703 ( .A(n4564), .ZN(n3330) );
  OR2_X1 U3704 ( .A1(n3248), .A2(n3247), .ZN(n4705) );
  INV_X2 U3705 ( .A(n3962), .ZN(n4689) );
  NAND4_X2 U3706 ( .A1(n3292), .A2(n3291), .A3(n3290), .A4(n3289), .ZN(n3962)
         );
  OR2_X2 U3707 ( .A1(n3187), .A2(n3186), .ZN(n4213) );
  NAND2_X2 U3708 ( .A1(n3218), .A2(n3217), .ZN(n3249) );
  AND4_X1 U3709 ( .A1(n3230), .A2(n3229), .A3(n3228), .A4(n3227), .ZN(n3236)
         );
  AND4_X1 U3710 ( .A1(n3226), .A2(n3225), .A3(n3224), .A4(n3223), .ZN(n3237)
         );
  AND4_X1 U3711 ( .A1(n3212), .A2(n3211), .A3(n3210), .A4(n3209), .ZN(n3218)
         );
  AND4_X1 U3712 ( .A1(n3216), .A2(n3215), .A3(n3214), .A4(n3213), .ZN(n3217)
         );
  AND4_X1 U3713 ( .A1(n3256), .A2(n3255), .A3(n3254), .A4(n3253), .ZN(n3272)
         );
  BUF_X2 U3714 ( .A(n3351), .Z(n4163) );
  BUF_X2 U3715 ( .A(n3358), .Z(n4165) );
  INV_X2 U3716 ( .A(n3474), .ZN(n3408) );
  BUF_X2 U3717 ( .A(n3406), .Z(n4171) );
  INV_X2 U3718 ( .A(n6741), .ZN(n6727) );
  AND2_X1 U3719 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4593) );
  NOR2_X2 U3720 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6442) );
  CLKBUF_X1 U3721 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n6988) );
  NAND2_X1 U3722 ( .A1(n4544), .A2(n4225), .ZN(n6344) );
  NOR2_X1 U3723 ( .A1(n5785), .A2(n5778), .ZN(n3140) );
  AND2_X1 U3724 ( .A1(n3140), .A2(n3141), .ZN(n5579) );
  AND2_X1 U3725 ( .A1(n4137), .A2(n3819), .ZN(n3141) );
  AND2_X1 U3726 ( .A1(n3718), .A2(n3702), .ZN(n3143) );
  AND2_X1 U3727 ( .A1(n3142), .A2(n3702), .ZN(n5728) );
  NOR2_X1 U3728 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3181) );
  AND2_X2 U3729 ( .A1(n3179), .A2(n3177), .ZN(n3351) );
  NAND3_X1 U3730 ( .A1(n3329), .A2(n3252), .A3(n3251), .ZN(n3312) );
  NOR2_X4 U3731 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3177) );
  AND2_X2 U3732 ( .A1(n3330), .A2(n3299), .ZN(n3704) );
  AND2_X1 U3733 ( .A1(n4593), .A2(n3181), .ZN(n3144) );
  AND2_X2 U3734 ( .A1(n4593), .A2(n3181), .ZN(n4164) );
  AND2_X1 U3735 ( .A1(n3176), .A2(n3177), .ZN(n3145) );
  AND2_X1 U3736 ( .A1(n4411), .A2(n3890), .ZN(n4438) );
  NOR2_X4 U3737 ( .A1(n4947), .A2(n4940), .ZN(n4942) );
  OR2_X1 U3738 ( .A1(n5579), .A2(n5580), .ZN(n5581) );
  OR2_X2 U3739 ( .A1(n4945), .A2(n4944), .ZN(n4947) );
  AND2_X2 U3740 ( .A1(n4552), .A2(n4553), .ZN(n4551) );
  NOR2_X1 U3741 ( .A1(n3960), .A2(n3151), .ZN(n5291) );
  AND2_X1 U3742 ( .A1(n4627), .A2(n5551), .ZN(n3147) );
  AND2_X1 U3743 ( .A1(n4627), .A2(n5551), .ZN(n3148) );
  NOR2_X4 U3744 ( .A1(n5654), .A2(n5644), .ZN(n5643) );
  AND2_X2 U3745 ( .A1(n4593), .A2(n3181), .ZN(n3149) );
  AND2_X2 U3746 ( .A1(n3178), .A2(n5551), .ZN(n3155) );
  OR2_X2 U3747 ( .A1(n5651), .A2(n5652), .ZN(n5654) );
  NOR2_X4 U3748 ( .A1(n5346), .A2(n5307), .ZN(n5357) );
  AND2_X2 U3749 ( .A1(n4551), .A2(n4574), .ZN(n4573) );
  NOR2_X4 U3750 ( .A1(n5051), .A2(n5050), .ZN(n5222) );
  NAND4_X1 U3751 ( .A1(n3292), .A2(n3291), .A3(n3290), .A4(n3289), .ZN(n3150)
         );
  NAND4_X1 U3752 ( .A1(n3292), .A2(n3291), .A3(n3290), .A4(n3289), .ZN(n3151)
         );
  INV_X1 U3753 ( .A(n3972), .ZN(n3152) );
  OAI21_X2 U3754 ( .B1(n3449), .B2(STATE2_REG_0__SCAN_IN), .A(n3448), .ZN(
        n3447) );
  NAND4_X1 U3755 ( .A1(n3292), .A2(n3291), .A3(n3290), .A4(n3289), .ZN(n3153)
         );
  NAND4_X1 U3756 ( .A1(n3292), .A2(n3291), .A3(n3290), .A4(n3289), .ZN(n3154)
         );
  AND2_X1 U3757 ( .A1(n3178), .A2(n5551), .ZN(n3156) );
  AND2_X1 U3758 ( .A1(n3178), .A2(n5551), .ZN(n3357) );
  AND2_X2 U3759 ( .A1(n3170), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3176)
         );
  AND2_X1 U3760 ( .A1(n4114), .A2(n5655), .ZN(n4410) );
  INV_X1 U3761 ( .A(n4191), .ZN(n4185) );
  AND2_X1 U3762 ( .A1(n4364), .A2(n4197), .ZN(n4327) );
  NOR2_X1 U3763 ( .A1(n4588), .A2(n4369), .ZN(n4374) );
  NOR2_X1 U3764 ( .A1(n4699), .A2(n3401), .ZN(n3420) );
  NAND3_X1 U3765 ( .A1(n3249), .A2(STATE2_REG_0__SCAN_IN), .A3(n3962), .ZN(
        n3944) );
  AND2_X1 U3766 ( .A1(n4450), .A2(n4451), .ZN(n4056) );
  NOR2_X1 U3767 ( .A1(n4056), .A2(n4059), .ZN(n4054) );
  OR2_X1 U3768 ( .A1(n4473), .A2(n4683), .ZN(n6316) );
  AND2_X1 U3769 ( .A1(n4407), .A2(n5655), .ZN(n4408) );
  NAND2_X1 U3770 ( .A1(n6601), .A2(n6606), .ZN(n4472) );
  NOR2_X1 U3771 ( .A1(n5562), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5565)
         );
  NOR2_X1 U3772 ( .A1(n3944), .A2(n4270), .ZN(n3935) );
  CLKBUF_X1 U3773 ( .A(n3480), .Z(n4084) );
  NAND2_X1 U3774 ( .A1(n3512), .A2(n3513), .ZN(n3539) );
  INV_X1 U3775 ( .A(n4188), .ZN(n4156) );
  OR2_X1 U3776 ( .A1(n3400), .A2(n3399), .ZN(n4275) );
  XNOR2_X1 U3777 ( .A(n3369), .B(n3368), .ZN(n3433) );
  OAI22_X1 U3778 ( .A1(n4614), .A2(STATE2_REG_0__SCAN_IN), .B1(n4228), .B2(
        n4699), .ZN(n3369) );
  INV_X1 U3779 ( .A(n4640), .ZN(n4839) );
  INV_X1 U3780 ( .A(n6012), .ZN(n5066) );
  NOR2_X1 U3781 ( .A1(n3157), .A2(n3234), .ZN(n3235) );
  AND2_X1 U3782 ( .A1(n6502), .A2(n3346), .ZN(n4711) );
  OAI21_X1 U3783 ( .B1(n6736), .B2(n4647), .A(n6705), .ZN(n4661) );
  NAND2_X1 U3784 ( .A1(n4056), .A2(n3954), .ZN(n5754) );
  NAND2_X1 U3785 ( .A1(n3365), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4699) );
  INV_X1 U3786 ( .A(n4472), .ZN(n4568) );
  AND2_X1 U3787 ( .A1(n4410), .A2(n4136), .ZN(n4137) );
  NAND2_X1 U3788 ( .A1(n4411), .A2(n4410), .ZN(n5613) );
  NAND2_X1 U3789 ( .A1(n3868), .A2(n3867), .ZN(n5642) );
  INV_X1 U3790 ( .A(n5711), .ZN(n3718) );
  INV_X1 U3791 ( .A(n5281), .ZN(n3589) );
  INV_X1 U3792 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6977) );
  NAND2_X1 U3793 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3495), .ZN(n3521)
         );
  NOR2_X1 U3794 ( .A1(n6774), .A2(n3521), .ZN(n3541) );
  NOR4_X1 U3795 ( .A1(n5504), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n5515), .ZN(n4306) );
  AND2_X1 U3796 ( .A1(n5880), .A2(n6073), .ZN(n4302) );
  NAND2_X1 U3797 ( .A1(n6415), .A2(n4379), .ZN(n6090) );
  XNOR2_X1 U3798 ( .A(n3441), .B(n3440), .ZN(n4216) );
  XNOR2_X1 U3799 ( .A(n3439), .B(n3438), .ZN(n3441) );
  AND2_X1 U3800 ( .A1(n4613), .A2(n4612), .ZN(n6582) );
  NOR2_X1 U3801 ( .A1(n4713), .A2(n4640), .ZN(n4772) );
  NOR2_X1 U3802 ( .A1(n4713), .A2(n4839), .ZN(n4660) );
  AND2_X1 U3803 ( .A1(n5381), .A2(n4839), .ZN(n4845) );
  INV_X1 U3804 ( .A(n5379), .ZN(n4964) );
  AND2_X1 U3805 ( .A1(n6709), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4565) );
  OAI22_X1 U3806 ( .A1(n3939), .A2(n3938), .B1(n3937), .B2(n3936), .ZN(n3941)
         );
  OR2_X1 U3807 ( .A1(n3909), .A2(n3908), .ZN(n3911) );
  AND2_X1 U3808 ( .A1(n6590), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3908)
         );
  NAND2_X1 U3809 ( .A1(n4054), .A2(n3961), .ZN(n6257) );
  OR2_X1 U3810 ( .A1(n4438), .A2(n4437), .ZN(n4441) );
  INV_X1 U3811 ( .A(n4439), .ZN(n4440) );
  AND2_X1 U3812 ( .A1(n5816), .A2(n5495), .ZN(n6271) );
  INV_X1 U3813 ( .A(n5816), .ZN(n6743) );
  AND2_X1 U3814 ( .A1(n5816), .A2(n4572), .ZN(n6742) );
  INV_X1 U3815 ( .A(n4445), .ZN(n4446) );
  NAND2_X1 U3816 ( .A1(n6355), .A2(n4200), .ZN(n6342) );
  INV_X1 U3817 ( .A(n6352), .ZN(n6336) );
  NAND2_X1 U3818 ( .A1(n6342), .A2(n6357), .ZN(n6352) );
  AOI21_X1 U3819 ( .B1(n5526), .B2(n5615), .A(n5525), .ZN(n5531) );
  XNOR2_X1 U3820 ( .A(n5519), .B(n5518), .ZN(n5539) );
  NAND2_X1 U3821 ( .A1(n4380), .A2(n4331), .ZN(n6425) );
  INV_X1 U3822 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n7014) );
  NAND2_X1 U3823 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6601), .ZN(n6705) );
  NAND2_X1 U3824 ( .A1(n4213), .A2(n4196), .ZN(n3329) );
  INV_X1 U3825 ( .A(n3538), .ZN(n3536) );
  OR2_X1 U3826 ( .A1(n3553), .A2(n3552), .ZN(n4266) );
  OR2_X1 U3827 ( .A1(n3509), .A2(n3508), .ZN(n4247) );
  OR2_X1 U3828 ( .A1(n3382), .A2(n3381), .ZN(n4217) );
  INV_X1 U3829 ( .A(n3296), .ZN(n3306) );
  OR2_X1 U3830 ( .A1(n3486), .A2(n3485), .ZN(n4210) );
  OAI211_X1 U3831 ( .C1(n3320), .C2(n5560), .A(n3316), .B(n3315), .ZN(n3341)
         );
  AND2_X1 U3832 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n3956), .ZN(n4108)
         );
  NAND2_X1 U3833 ( .A1(n3704), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4188) );
  INV_X1 U3834 ( .A(n5364), .ZN(n3652) );
  AND2_X1 U3835 ( .A1(n5495), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3493) );
  NAND2_X1 U3836 ( .A1(n4285), .A2(n5371), .ZN(n5352) );
  NAND2_X1 U3837 ( .A1(n4281), .A2(n4280), .ZN(n5315) );
  NAND2_X1 U3838 ( .A1(n3489), .A2(n3490), .ZN(n3515) );
  NAND2_X1 U3839 ( .A1(n4198), .A2(n3979), .ZN(n4587) );
  INV_X1 U3840 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6579) );
  AOI21_X1 U3841 ( .B1(n3935), .B2(n3934), .A(n3933), .ZN(n3938) );
  INV_X1 U3842 ( .A(n4456), .ZN(n6735) );
  NOR2_X1 U3843 ( .A1(n5679), .A2(n4061), .ZN(n4416) );
  AND2_X1 U3844 ( .A1(n6018), .A2(REIP_REG_17__SCAN_IN), .ZN(n6027) );
  AND2_X1 U3845 ( .A1(n3606), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3631)
         );
  OR2_X1 U3846 ( .A1(n5789), .A2(n4038), .ZN(n5686) );
  NAND2_X1 U3847 ( .A1(n4374), .A2(n4373), .ZN(n4697) );
  OR2_X1 U3848 ( .A1(n4138), .A2(n5583), .ZN(n4160) );
  NOR2_X1 U3849 ( .A1(n3860), .A2(n5659), .ZN(n3886) );
  AND2_X1 U3850 ( .A1(n5658), .A2(n4185), .ZN(n3844) );
  NOR2_X1 U3851 ( .A1(n5668), .A2(n5669), .ZN(n3819) );
  AND2_X1 U3852 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3815), .ZN(n3816)
         );
  NAND2_X1 U3853 ( .A1(n3816), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3860)
         );
  NOR2_X1 U3854 ( .A1(n3768), .A2(n5898), .ZN(n3769) );
  NAND2_X1 U3855 ( .A1(n3769), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3814)
         );
  NOR2_X1 U3856 ( .A1(n3735), .A2(n3720), .ZN(n3736) );
  NAND2_X1 U3857 ( .A1(n3736), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3768)
         );
  CLKBUF_X1 U3858 ( .A(n5698), .Z(n5798) );
  NAND2_X1 U3859 ( .A1(n3703), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3719)
         );
  INV_X1 U3860 ( .A(n5729), .ZN(n3702) );
  NAND2_X1 U3861 ( .A1(n3654), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3655)
         );
  OR2_X1 U3862 ( .A1(n6981), .A2(n3655), .ZN(n3671) );
  INV_X1 U3863 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6981) );
  AND2_X1 U3864 ( .A1(n3635), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3654)
         );
  CLKBUF_X1 U3865 ( .A(n5304), .Z(n5305) );
  CLKBUF_X1 U3866 ( .A(n5363), .Z(n5436) );
  AND2_X1 U3867 ( .A1(n3631), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3635)
         );
  AND2_X1 U3868 ( .A1(n3588), .A2(n3587), .ZN(n5281) );
  AND3_X1 U3869 ( .A1(n3586), .A2(n3585), .A3(n3584), .ZN(n3587) );
  NAND2_X1 U3870 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n3541), .ZN(n3554)
         );
  NOR2_X1 U3871 ( .A1(n6890), .A2(n3554), .ZN(n3566) );
  OR2_X1 U3872 ( .A1(n6715), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6728) );
  NAND2_X1 U3873 ( .A1(n3517), .A2(n3695), .ZN(n3525) );
  NAND2_X1 U3874 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3494) );
  CLKBUF_X1 U3875 ( .A(n4413), .Z(n5628) );
  AND2_X1 U3876 ( .A1(n4045), .A2(n4044), .ZN(n5644) );
  NOR2_X2 U3877 ( .A1(n5686), .A2(n5685), .ZN(n5687) );
  CLKBUF_X1 U3878 ( .A(n5651), .Z(n5674) );
  AND2_X1 U3879 ( .A1(n4026), .A2(n4025), .ZN(n5700) );
  AND2_X1 U3880 ( .A1(n4018), .A2(n4017), .ZN(n5453) );
  AND2_X1 U3881 ( .A1(n4288), .A2(n5467), .ZN(n5442) );
  AND2_X1 U3882 ( .A1(n4016), .A2(n4015), .ZN(n5437) );
  CLKBUF_X1 U3883 ( .A(n5352), .Z(n5464) );
  XNOR2_X1 U3884 ( .A(n4236), .B(n7003), .ZN(n4556) );
  OR2_X1 U3885 ( .A1(n6416), .A2(n4386), .ZN(n5447) );
  INV_X1 U3886 ( .A(n3416), .ZN(n3448) );
  AND2_X1 U3887 ( .A1(n4840), .A2(n6442), .ZN(n4842) );
  AND2_X1 U3888 ( .A1(n5382), .A2(n6442), .ZN(n5387) );
  AND2_X1 U3889 ( .A1(n5383), .A2(n6439), .ZN(n6507) );
  OAI21_X1 U3890 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6702), .A(n5000), 
        .ZN(n6508) );
  NOR2_X1 U3891 ( .A1(n4730), .A2(n5066), .ZN(n5381) );
  OR3_X1 U3892 ( .A1(n6012), .A2(n4642), .A3(n4640), .ZN(n4674) );
  NAND2_X1 U3893 ( .A1(n5542), .A2(n4661), .ZN(n4806) );
  OR2_X1 U3894 ( .A1(n6012), .A2(n4957), .ZN(n4965) );
  INV_X2 U3895 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6935) );
  NOR2_X1 U3896 ( .A1(n6935), .A2(n6709), .ZN(n4647) );
  INV_X1 U3897 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6975) );
  INV_X1 U3898 ( .A(n6616), .ZN(n6736) );
  AND2_X1 U3899 ( .A1(n5754), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6239) );
  AND2_X1 U3900 ( .A1(n6732), .A2(n4060), .ZN(n6246) );
  INV_X1 U3901 ( .A(n6239), .ZN(n6253) );
  NAND2_X1 U3902 ( .A1(n4058), .A2(n4428), .ZN(n6264) );
  INV_X1 U3903 ( .A(n6257), .ZN(n6155) );
  INV_X1 U3904 ( .A(n5878), .ZN(n5829) );
  CLKBUF_X1 U3905 ( .A(n5494), .Z(n6273) );
  AOI22_X1 U3906 ( .A1(n4569), .A2(n4568), .B1(n4567), .B2(n4566), .ZN(n4570)
         );
  INV_X1 U3907 ( .A(n6742), .ZN(n5481) );
  AND2_X1 U3908 ( .A1(n4523), .A2(n6627), .ZN(n6298) );
  INV_X1 U3909 ( .A(n6730), .ZN(n6305) );
  INV_X1 U3910 ( .A(n6298), .ZN(n6307) );
  AND2_X1 U3911 ( .A1(n4473), .A2(n6329), .ZN(n6327) );
  INV_X1 U3912 ( .A(n6329), .ZN(n6330) );
  INV_X1 U3913 ( .A(n6316), .ZN(n6331) );
  INV_X1 U3914 ( .A(n6327), .ZN(n6333) );
  INV_X1 U3915 ( .A(n6017), .ZN(n6054) );
  INV_X1 U3916 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6890) );
  INV_X1 U3917 ( .A(n6342), .ZN(n6358) );
  INV_X1 U3918 ( .A(n4306), .ZN(n4307) );
  OR2_X1 U3919 ( .A1(n6087), .A2(n4393), .ZN(n5979) );
  OAI21_X1 U3920 ( .B1(n6399), .B2(n5474), .A(n5446), .ZN(n6366) );
  OR2_X1 U3921 ( .A1(n5226), .A2(n5225), .ZN(n6384) );
  AND2_X1 U3922 ( .A1(n6415), .A2(n5447), .ZN(n6399) );
  INV_X1 U3923 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4838) );
  INV_X1 U3924 ( .A(n6442), .ZN(n6729) );
  INV_X1 U3925 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6590) );
  AND3_X1 U3926 ( .A1(n4649), .A2(n6571), .A3(n6122), .ZN(n4637) );
  INV_X1 U3927 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5560) );
  INV_X1 U3928 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3171) );
  NAND2_X1 U3929 ( .A1(n6702), .A2(n6709), .ZN(n6715) );
  INV_X1 U3930 ( .A(n6713), .ZN(n6707) );
  CLKBUF_X1 U3931 ( .A(n4329), .Z(n6108) );
  INV_X1 U3932 ( .A(n5164), .ZN(n5212) );
  INV_X1 U3933 ( .A(n5165), .ZN(n5211) );
  NOR2_X1 U3934 ( .A1(n4737), .A2(n5379), .ZN(n5002) );
  NOR2_X1 U3935 ( .A1(n4737), .A2(n4964), .ZN(n5164) );
  INV_X1 U3936 ( .A(n5003), .ZN(n5101) );
  INV_X1 U3937 ( .A(n4719), .ZN(n5100) );
  OR3_X1 U3938 ( .A1(n6449), .A2(n6448), .A3(n6447), .ZN(n6479) );
  AND2_X1 U3939 ( .A1(n4845), .A2(n4964), .ZN(n5431) );
  INV_X1 U3940 ( .A(n4895), .ZN(n4925) );
  NOR2_X1 U3941 ( .A1(n4674), .A2(n4964), .ZN(n4895) );
  INV_X1 U3942 ( .A(n6520), .ZN(n5425) );
  INV_X1 U3943 ( .A(n6526), .ZN(n5409) );
  INV_X1 U3944 ( .A(n6532), .ZN(n5414) );
  INV_X1 U3945 ( .A(n6538), .ZN(n5420) );
  INV_X1 U3946 ( .A(n6551), .ZN(n5404) );
  INV_X1 U3947 ( .A(n5113), .ZN(n5139) );
  OAI211_X1 U3948 ( .C1(n5142), .C2(n6702), .A(n5118), .B(n5117), .ZN(n5143)
         );
  INV_X1 U3949 ( .A(n6561), .ZN(n5394) );
  NOR2_X1 U3950 ( .A1(n4690), .A2(n4900), .ZN(n6514) );
  NOR2_X1 U3951 ( .A1(n4655), .A2(n4900), .ZN(n6526) );
  NOR2_X1 U3952 ( .A1(n4678), .A2(n4900), .ZN(n6532) );
  NOR2_X1 U3953 ( .A1(n6918), .A2(n4900), .ZN(n6538) );
  NOR2_X1 U3954 ( .A1(n4799), .A2(n4900), .ZN(n6544) );
  NOR2_X1 U3955 ( .A1(n5039), .A2(n4900), .ZN(n6551) );
  NOR2_X1 U3956 ( .A1(n4965), .A2(n5379), .ZN(n5165) );
  NOR2_X1 U3957 ( .A1(n4965), .A2(n4964), .ZN(n5114) );
  NOR2_X1 U3958 ( .A1(n5049), .A2(n4900), .ZN(n6561) );
  NAND2_X1 U3959 ( .A1(n3935), .A2(n3947), .ZN(n3950) );
  INV_X1 U3960 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6709) );
  INV_X1 U3961 ( .A(n6606), .ZN(n6612) );
  INV_X1 U3962 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6974) );
  INV_X1 U3963 ( .A(n6683), .ZN(n6689) );
  INV_X1 U3964 ( .A(n4434), .ZN(n4435) );
  INV_X1 U3965 ( .A(n5586), .ZN(n5587) );
  AOI21_X1 U3966 ( .B1(n6336), .B2(n5606), .A(n5584), .ZN(n5585) );
  INV_X1 U3967 ( .A(n4447), .ZN(n4448) );
  OAI21_X1 U3968 ( .B1(n5955), .B2(n6355), .A(n4446), .ZN(n4447) );
  AOI21_X1 U3969 ( .B1(n5601), .B2(n6390), .A(n5537), .ZN(n5538) );
  NAND2_X1 U3970 ( .A1(n5536), .A2(n5535), .ZN(n5537) );
  AOI21_X1 U3971 ( .B1(n5534), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5533), 
        .ZN(n5535) );
  NAND2_X1 U3972 ( .A1(n4942), .A2(n4937), .ZN(n4706) );
  AND2_X1 U3973 ( .A1(n4089), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3157) );
  NAND2_X1 U3974 ( .A1(n3143), .A2(n3142), .ZN(n5697) );
  NAND2_X1 U3975 ( .A1(n4380), .A2(n4356), .ZN(n6424) );
  NAND2_X1 U3976 ( .A1(n4805), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3648) );
  INV_X1 U3977 ( .A(n3648), .ZN(n3695) );
  INV_X1 U3978 ( .A(n4270), .ZN(n4314) );
  NAND2_X1 U3979 ( .A1(n3488), .A2(n3487), .ZN(n3490) );
  INV_X1 U3980 ( .A(n4706), .ZN(n3991) );
  INV_X1 U3981 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3170) );
  INV_X1 U3982 ( .A(n3983), .ZN(n5780) );
  NAND2_X1 U3983 ( .A1(n4213), .A2(n3960), .ZN(n3983) );
  OR2_X1 U3984 ( .A1(n3317), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3158)
         );
  OR2_X1 U3985 ( .A1(n6569), .A2(n4472), .ZN(n6355) );
  INV_X1 U3986 ( .A(n6355), .ZN(n4310) );
  INV_X1 U3987 ( .A(n5834), .ZN(n6744) );
  OR2_X1 U3988 ( .A1(n5631), .A2(REIP_REG_25__SCAN_IN), .ZN(n3159) );
  AND2_X1 U3989 ( .A1(n3767), .A2(n3766), .ZN(n3160) );
  AND2_X1 U3990 ( .A1(n4411), .A2(n4408), .ZN(n4439) );
  AND4_X1 U3991 ( .A1(n3222), .A2(n3221), .A3(n3220), .A4(n3219), .ZN(n3161)
         );
  OR2_X1 U3992 ( .A1(n6253), .A2(n5852), .ZN(n3162) );
  AND2_X1 U3993 ( .A1(n5880), .A2(n5443), .ZN(n3163) );
  NOR2_X1 U3994 ( .A1(n5880), .A2(n5443), .ZN(n3164) );
  NAND2_X1 U3995 ( .A1(n5880), .A2(n7012), .ZN(n3165) );
  NOR2_X1 U3996 ( .A1(n5329), .A2(n4282), .ZN(n3166) );
  AND2_X1 U3997 ( .A1(n4003), .A2(n4002), .ZN(n3167) );
  INV_X1 U3998 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6835) );
  INV_X1 U3999 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5518) );
  INV_X1 U4000 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6774) );
  AND2_X1 U4001 ( .A1(n5814), .A2(n4705), .ZN(n5810) );
  AND2_X1 U4002 ( .A1(n5534), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n3168)
         );
  AOI21_X1 U4003 ( .B1(n5642), .B2(n3891), .A(n4438), .ZN(n5498) );
  INV_X1 U4004 ( .A(n3567), .ZN(n4154) );
  NAND2_X1 U4005 ( .A1(n6442), .A2(n6709), .ZN(n3169) );
  NAND2_X2 U4006 ( .A1(n4704), .A2(n4703), .ZN(n5814) );
  INV_X1 U4007 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3921) );
  AOI21_X1 U4008 ( .B1(n4683), .B2(n5493), .A(n3146), .ZN(n3937) );
  AND2_X1 U4009 ( .A1(n4364), .A2(n3298), .ZN(n3337) );
  AND2_X1 U4010 ( .A1(n3295), .A2(n4587), .ZN(n3328) );
  AND2_X1 U4011 ( .A1(n4838), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3920)
         );
  OR2_X1 U4012 ( .A1(n3364), .A2(n3363), .ZN(n3366) );
  OR3_X1 U4013 ( .A1(n3909), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(n6590), 
        .ZN(n3907) );
  INV_X1 U4014 ( .A(n4217), .ZN(n3425) );
  OR2_X1 U4015 ( .A1(n3535), .A2(n3534), .ZN(n4250) );
  INV_X1 U4016 ( .A(n3366), .ZN(n4228) );
  OR2_X1 U4017 ( .A1(n3962), .A2(n6609), .ZN(n3473) );
  NAND2_X1 U4018 ( .A1(n3303), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3320) );
  NOR2_X1 U4019 ( .A1(n4705), .A2(n6935), .ZN(n3567) );
  INV_X1 U4020 ( .A(n3944), .ZN(n3916) );
  INV_X1 U4021 ( .A(n4662), .ZN(n4361) );
  AOI21_X1 U4022 ( .B1(n3294), .B2(n4361), .A(n5815), .ZN(n3252) );
  INV_X1 U4023 ( .A(n4275), .ZN(n3401) );
  INV_X1 U4024 ( .A(n3979), .ZN(n4004) );
  NOR2_X1 U4025 ( .A1(n4107), .A2(n5852), .ZN(n4115) );
  INV_X1 U4026 ( .A(n3814), .ZN(n3815) );
  OAI21_X1 U4027 ( .B1(n4271), .B2(n4270), .A(n4269), .ZN(n4272) );
  OR3_X1 U4028 ( .A1(n5989), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n5931), 
        .ZN(n5515) );
  INV_X1 U4029 ( .A(n5442), .ZN(n4289) );
  AND2_X1 U4030 ( .A1(n3996), .A2(n3995), .ZN(n4755) );
  NAND2_X1 U4031 ( .A1(n4640), .A2(n4314), .ZN(n4223) );
  AOI21_X1 U4032 ( .B1(n3343), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3347), 
        .ZN(n3348) );
  OR2_X1 U4033 ( .A1(n3414), .A2(n3413), .ZN(n4218) );
  AND2_X1 U4034 ( .A1(n3911), .A2(n3910), .ZN(n3947) );
  INV_X1 U4035 ( .A(n4707), .ZN(n3990) );
  NAND2_X1 U4036 ( .A1(n4010), .A2(n4004), .ZN(n4796) );
  INV_X1 U4037 ( .A(n3861), .ZN(n4192) );
  NAND2_X1 U4038 ( .A1(n4115), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4138)
         );
  AOI21_X1 U4039 ( .B1(n3846), .B2(n3845), .A(n3844), .ZN(n5655) );
  OR2_X1 U4040 ( .A1(n3719), .A2(n5723), .ZN(n3735) );
  OR2_X1 U4041 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4191) );
  INV_X1 U4042 ( .A(n3494), .ZN(n3495) );
  INV_X1 U4043 ( .A(n5515), .ZN(n5516) );
  OR2_X1 U4044 ( .A1(n5858), .A2(n4300), .ZN(n5838) );
  NOR2_X1 U4045 ( .A1(n3163), .A2(n4289), .ZN(n4290) );
  NAND2_X1 U4046 ( .A1(n4283), .A2(n3166), .ZN(n5369) );
  NAND2_X1 U4047 ( .A1(n5493), .A2(n4357), .ZN(n4270) );
  OAI21_X1 U4048 ( .B1(n6344), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .A(n6343), 
        .ZN(n4235) );
  AND2_X1 U4049 ( .A1(n4732), .A2(n6442), .ZN(n4734) );
  INV_X1 U4050 ( .A(n4900), .ZN(n5000) );
  INV_X1 U4051 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6586) );
  INV_X1 U4052 ( .A(n3490), .ZN(n4642) );
  NAND2_X1 U4053 ( .A1(n3472), .A2(n3471), .ZN(n4897) );
  AND2_X1 U4054 ( .A1(n6439), .A2(n6575), .ZN(n4956) );
  OR2_X1 U4055 ( .A1(n4602), .A2(n4472), .ZN(n4451) );
  AND2_X1 U4056 ( .A1(n5632), .A2(REIP_REG_27__SCAN_IN), .ZN(n4420) );
  INV_X1 U4057 ( .A(n4931), .ZN(n4352) );
  INV_X1 U4058 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5723) );
  NOR2_X1 U4059 ( .A1(n3573), .A2(n6977), .ZN(n3606) );
  AND2_X1 U4060 ( .A1(n4204), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4053) );
  INV_X1 U4061 ( .A(n6264), .ZN(n6180) );
  AND2_X1 U4062 ( .A1(n4006), .A2(n4005), .ZN(n5343) );
  NAND2_X1 U4063 ( .A1(n3465), .A2(n3464), .ZN(n4552) );
  XNOR2_X1 U4064 ( .A(n3958), .B(n4427), .ZN(n4204) );
  NAND2_X1 U4065 ( .A1(n4108), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4107)
         );
  NOR2_X1 U4066 ( .A1(n6835), .A2(n3671), .ZN(n3703) );
  INV_X1 U4067 ( .A(n5181), .ZN(n3605) );
  INV_X1 U4068 ( .A(n5864), .ZN(n5989) );
  AND2_X1 U4069 ( .A1(n4382), .A2(n4381), .ZN(n5355) );
  INV_X1 U4071 ( .A(n5002), .ZN(n5033) );
  NAND2_X1 U4072 ( .A1(n4772), .A2(n4964), .ZN(n6450) );
  OR2_X1 U4073 ( .A1(n6012), .A2(n3490), .ZN(n4713) );
  INV_X1 U4074 ( .A(n6508), .ZN(n4959) );
  INV_X1 U4075 ( .A(n5114), .ZN(n5140) );
  NAND2_X1 U4076 ( .A1(n3950), .A2(n3949), .ZN(n6601) );
  OR2_X1 U4077 ( .A1(n4455), .A2(n6612), .ZN(n4450) );
  OAI21_X1 U4078 ( .B1(n5513), .B2(n6257), .A(n4433), .ZN(n4434) );
  AOI21_X1 U4079 ( .B1(n5618), .B2(n6680), .A(n4420), .ZN(n4421) );
  NAND2_X1 U4080 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n3566), .ZN(n3573)
         );
  AND2_X1 U4081 ( .A1(n5754), .A2(n4053), .ZN(n6196) );
  INV_X1 U4082 ( .A(n5754), .ZN(n6236) );
  NAND2_X1 U4083 ( .A1(n5224), .A2(n3167), .ZN(n5344) );
  INV_X1 U4084 ( .A(n5808), .ZN(n5811) );
  OR2_X1 U4085 ( .A1(n4697), .A2(n4696), .ZN(n4704) );
  INV_X1 U4086 ( .A(n6301), .ZN(n6304) );
  OR2_X1 U4087 ( .A1(n4586), .A2(n6735), .ZN(n6595) );
  OAI21_X1 U4088 ( .B1(n5603), .B2(n6361), .A(n5585), .ZN(n5586) );
  AND2_X1 U4089 ( .A1(n5639), .A2(n5656), .ZN(n5878) );
  OR2_X1 U4090 ( .A1(n4402), .A2(n3168), .ZN(n4403) );
  NOR2_X1 U4091 ( .A1(n6001), .A2(n5993), .ZN(n5984) );
  INV_X1 U4092 ( .A(n6424), .ZN(n6390) );
  CLKBUF_X1 U4093 ( .A(n4750), .Z(n4751) );
  INV_X1 U4094 ( .A(n6425), .ZN(n6420) );
  INV_X1 U4095 ( .A(n5763), .ZN(n6010) );
  NAND2_X1 U4096 ( .A1(n6609), .A2(n4661), .ZN(n4900) );
  OAI21_X1 U4097 ( .B1(n5163), .B2(n5162), .A(n5161), .ZN(n5210) );
  OAI21_X1 U4098 ( .B1(n5001), .B2(n5035), .A(n5389), .ZN(n5032) );
  OAI21_X1 U4099 ( .B1(n5079), .B2(n5078), .A(n5077), .ZN(n5104) );
  INV_X1 U4100 ( .A(n6439), .ZN(n6254) );
  INV_X1 U4101 ( .A(n6450), .ZN(n6477) );
  AND2_X1 U4102 ( .A1(n4660), .A2(n4964), .ZN(n6495) );
  INV_X1 U4103 ( .A(n6565), .ZN(n6549) );
  INV_X1 U4104 ( .A(n6554), .ZN(n6557) );
  OR2_X1 U4105 ( .A1(n4902), .A2(n4901), .ZN(n4924) );
  NOR2_X1 U4106 ( .A1(n4674), .A2(n5379), .ZN(n5113) );
  NOR2_X1 U4107 ( .A1(n4684), .A2(n4900), .ZN(n6520) );
  AND2_X1 U4108 ( .A1(n4565), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6606) );
  AND2_X1 U4109 ( .A1(n6600), .A2(n6599), .ZN(n6698) );
  INV_X1 U4110 ( .A(n6689), .ZN(n6675) );
  NOR2_X1 U4111 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6727), .ZN(n6683) );
  INV_X1 U4112 ( .A(n4056), .ZN(n6732) );
  OR2_X1 U4113 ( .A1(n4069), .A2(n4068), .ZN(n4070) );
  AND2_X1 U4114 ( .A1(n6171), .A2(n5292), .ZN(n6260) );
  NAND2_X1 U4115 ( .A1(n4441), .A2(n4440), .ZN(n6037) );
  NAND2_X1 U4116 ( .A1(n5814), .A2(n5815), .ZN(n5808) );
  OAI211_X2 U4117 ( .C1(n4608), .C2(n6612), .A(n4570), .B(n6316), .ZN(n5816)
         );
  OR2_X1 U4118 ( .A1(n6298), .A2(n6305), .ZN(n6301) );
  OR2_X1 U4119 ( .A1(n6595), .A2(n4472), .ZN(n6329) );
  NOR2_X1 U4120 ( .A1(n4404), .A2(n4403), .ZN(n4405) );
  INV_X1 U4121 ( .A(n5230), .ZN(n6388) );
  OAI21_X1 U4122 ( .B1(n6699), .B2(n4637), .A(n4900), .ZN(n6435) );
  INV_X1 U4123 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6113) );
  INV_X1 U4124 ( .A(n4771), .ZN(n4814) );
  NAND2_X1 U4125 ( .A1(n4660), .A2(n5379), .ZN(n6501) );
  AOI21_X1 U4126 ( .B1(n5241), .B2(n5239), .A(n5238), .ZN(n5277) );
  NAND2_X1 U4127 ( .A1(n4845), .A2(n5379), .ZN(n5272) );
  AOI21_X1 U4128 ( .B1(n5387), .B2(n6507), .A(n5385), .ZN(n5434) );
  NAND2_X1 U4129 ( .A1(n5381), .A2(n4894), .ZN(n6554) );
  INV_X1 U4130 ( .A(n6514), .ZN(n5433) );
  INV_X1 U4131 ( .A(n6544), .ZN(n5399) );
  INV_X1 U4132 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6609) );
  INV_X1 U4133 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6702) );
  INV_X1 U4134 ( .A(n6687), .ZN(n6685) );
  OR2_X1 U4135 ( .A1(n4424), .A2(n4423), .ZN(U2800) );
  NOR2_X2 U4136 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n4622), .ZN(n3179)
         );
  AND2_X4 U4137 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5551) );
  AOI22_X1 U4138 ( .A1(n3351), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3175) );
  AND2_X2 U4139 ( .A1(n3921), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3180)
         );
  NOR2_X4 U4140 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3178) );
  AND2_X4 U4141 ( .A1(n3180), .A2(n3178), .ZN(n4174) );
  AOI22_X1 U4142 ( .A1(n4174), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4089), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3174) );
  AND2_X2 U4143 ( .A1(n5557), .A2(n3178), .ZN(n3406) );
  AOI22_X1 U4144 ( .A1(n3406), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3173) );
  AOI22_X1 U4145 ( .A1(n4121), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3172) );
  NAND4_X1 U4146 ( .A1(n3175), .A2(n3174), .A3(n3173), .A4(n3172), .ZN(n3187)
         );
  AND2_X2 U4147 ( .A1(n3180), .A2(n3176), .ZN(n3480) );
  AND2_X2 U4148 ( .A1(n3179), .A2(n5557), .ZN(n3208) );
  AOI22_X1 U4149 ( .A1(n3480), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3185) );
  AND2_X2 U4150 ( .A1(n5557), .A2(n3176), .ZN(n3242) );
  AND2_X2 U4151 ( .A1(n3178), .A2(n3177), .ZN(n3830) );
  AOI22_X1 U4152 ( .A1(n3242), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3830), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3184) );
  AND2_X4 U4153 ( .A1(n3179), .A2(n5551), .ZN(n4161) );
  AOI22_X1 U4154 ( .A1(n4161), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3357), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3183) );
  AND2_X2 U4155 ( .A1(n3180), .A2(n4627), .ZN(n3358) );
  AOI22_X1 U4156 ( .A1(n3358), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4164), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3182) );
  NAND4_X1 U4157 ( .A1(n3185), .A2(n3184), .A3(n3183), .A4(n3182), .ZN(n3186)
         );
  AOI22_X1 U4158 ( .A1(n3480), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3191) );
  AOI22_X1 U4159 ( .A1(n3242), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3830), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3190) );
  AOI22_X1 U4160 ( .A1(n4161), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3155), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3189) );
  AOI22_X1 U4161 ( .A1(n3358), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4164), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3188) );
  NAND4_X1 U4162 ( .A1(n3191), .A2(n3190), .A3(n3189), .A4(n3188), .ZN(n3197)
         );
  AOI22_X1 U4163 ( .A1(n3351), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3195) );
  AOI22_X1 U4164 ( .A1(n4174), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3194) );
  AOI22_X1 U4165 ( .A1(n3406), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3148), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3193) );
  AOI22_X1 U4166 ( .A1(n4121), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3192) );
  NAND4_X1 U4167 ( .A1(n3195), .A2(n3194), .A3(n3193), .A4(n3192), .ZN(n3196)
         );
  AOI22_X1 U4169 ( .A1(n3480), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3201) );
  AOI22_X1 U4170 ( .A1(n3208), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4089), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3200) );
  AOI22_X1 U4171 ( .A1(n3830), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3144), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3199) );
  AOI22_X1 U4172 ( .A1(n3351), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3198) );
  NAND4_X1 U4173 ( .A1(n3201), .A2(n3200), .A3(n3199), .A4(n3198), .ZN(n3207)
         );
  AOI22_X1 U4174 ( .A1(n3242), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3205) );
  AOI22_X1 U4175 ( .A1(n4161), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4121), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3204) );
  AOI22_X1 U4176 ( .A1(n3358), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3147), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3203) );
  AOI22_X1 U4177 ( .A1(n3406), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3155), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3202) );
  NAND4_X1 U4178 ( .A1(n3205), .A2(n3204), .A3(n3203), .A4(n3202), .ZN(n3206)
         );
  OR2_X2 U4179 ( .A1(n3207), .A2(n3206), .ZN(n3299) );
  AOI22_X1 U4180 ( .A1(n3242), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3830), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3212) );
  AOI22_X1 U4181 ( .A1(n3480), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3211) );
  AOI22_X1 U4182 ( .A1(n4161), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3155), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3210) );
  AOI22_X1 U4183 ( .A1(n3358), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4164), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3209) );
  AOI22_X1 U4184 ( .A1(n3351), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3216) );
  AOI22_X1 U4185 ( .A1(n4174), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3215) );
  AOI22_X1 U4186 ( .A1(n3406), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3214) );
  AOI22_X1 U4187 ( .A1(n4121), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3213) );
  INV_X1 U4188 ( .A(n3249), .ZN(n3304) );
  NAND2_X1 U4189 ( .A1(n3304), .A2(n3299), .ZN(n3294) );
  NAND2_X1 U4190 ( .A1(n3358), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3222)
         );
  NAND2_X1 U4191 ( .A1(n3242), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3221) );
  NAND2_X1 U4192 ( .A1(n3480), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3220)
         );
  NAND2_X1 U4193 ( .A1(n4121), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3219)
         );
  NAND2_X1 U4194 ( .A1(n3134), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3226)
         );
  NAND2_X1 U4195 ( .A1(n3351), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3225) );
  NAND2_X1 U4196 ( .A1(n3406), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3224) );
  NAND2_X1 U4197 ( .A1(n3475), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3223)
         );
  NAND2_X1 U4198 ( .A1(n4174), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3230) );
  NAND2_X1 U4199 ( .A1(n4161), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3229) );
  NAND2_X1 U4200 ( .A1(n3830), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3228) );
  NAND2_X1 U4201 ( .A1(n3352), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3227)
         );
  NAND2_X1 U4202 ( .A1(n3208), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3233) );
  NAND2_X1 U4203 ( .A1(n4164), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3232) );
  NAND2_X1 U4204 ( .A1(n3156), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3231) );
  NAND3_X1 U4205 ( .A1(n3233), .A2(n3232), .A3(n3231), .ZN(n3234) );
  AOI22_X1 U4206 ( .A1(n3351), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3241) );
  AOI22_X1 U4207 ( .A1(n4174), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4089), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3240) );
  AOI22_X1 U4208 ( .A1(n3406), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3239) );
  AOI22_X1 U4209 ( .A1(n4121), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3238) );
  NAND4_X1 U4210 ( .A1(n3241), .A2(n3240), .A3(n3239), .A4(n3238), .ZN(n3248)
         );
  AOI22_X1 U4211 ( .A1(n3242), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3830), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3246) );
  AOI22_X1 U4212 ( .A1(n3480), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3245) );
  AOI22_X1 U4213 ( .A1(n4161), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3155), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3244) );
  AOI22_X1 U4214 ( .A1(n3358), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4164), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3243) );
  NAND4_X1 U4215 ( .A1(n3246), .A2(n3245), .A3(n3244), .A4(n3243), .ZN(n3247)
         );
  NAND2_X1 U4216 ( .A1(n4662), .A2(n3299), .ZN(n3250) );
  MUX2_X1 U4217 ( .A(n3249), .B(n3250), .S(n4564), .Z(n3251) );
  NAND2_X1 U4218 ( .A1(n4121), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3256)
         );
  NAND2_X1 U4219 ( .A1(n3208), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3255) );
  NAND2_X1 U4220 ( .A1(n3242), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3254) );
  NAND2_X1 U4221 ( .A1(n3133), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3253)
         );
  NAND2_X1 U4222 ( .A1(n3480), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3260)
         );
  NAND2_X1 U4223 ( .A1(n3351), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3259) );
  NAND2_X1 U4224 ( .A1(n4161), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3258) );
  NAND2_X1 U4225 ( .A1(n3352), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3257)
         );
  NAND2_X1 U4226 ( .A1(n3358), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3264)
         );
  NAND2_X1 U4227 ( .A1(n3145), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3263) );
  NAND2_X1 U4228 ( .A1(n3830), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3262) );
  NAND2_X1 U4229 ( .A1(n4164), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3261) );
  NAND2_X1 U4230 ( .A1(n4174), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3268) );
  NAND2_X1 U4231 ( .A1(n3406), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3267) );
  NAND2_X1 U4232 ( .A1(n3155), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3266) );
  NAND2_X1 U4233 ( .A1(n3475), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3265)
         );
  NAND4_X4 U4235 ( .A1(n3272), .A2(n3271), .A3(n3270), .A4(n3269), .ZN(n3960)
         );
  NAND2_X1 U4236 ( .A1(n3208), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3276) );
  NAND2_X1 U4237 ( .A1(n3480), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3275)
         );
  NAND2_X1 U4238 ( .A1(n3242), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3274) );
  NAND2_X1 U4239 ( .A1(n3144), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3273) );
  NAND2_X1 U4240 ( .A1(n3358), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3280)
         );
  NAND2_X1 U4241 ( .A1(n4161), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3279) );
  NAND2_X1 U4242 ( .A1(n4121), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3278)
         );
  NAND2_X1 U4243 ( .A1(n3830), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3277) );
  NAND2_X1 U4244 ( .A1(n3390), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3284)
         );
  NAND2_X1 U4245 ( .A1(n3351), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3283) );
  NAND2_X1 U4246 ( .A1(n4089), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3282) );
  NAND2_X1 U4247 ( .A1(n3352), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3281)
         );
  NAND2_X1 U4248 ( .A1(n4174), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3288) );
  NAND2_X1 U4249 ( .A1(n3406), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3287) );
  NAND2_X1 U4250 ( .A1(n3156), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3286) );
  NAND2_X1 U4251 ( .A1(n3475), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3285)
         );
  NAND2_X1 U4252 ( .A1(n3312), .A2(n3146), .ZN(n3327) );
  NAND2_X1 U4253 ( .A1(n4800), .A2(n4564), .ZN(n3293) );
  NAND2_X1 U4254 ( .A1(n3293), .A2(n4705), .ZN(n3296) );
  NAND2_X1 U4255 ( .A1(n4315), .A2(n4456), .ZN(n3295) );
  INV_X1 U4256 ( .A(n3294), .ZN(n4198) );
  NAND2_X1 U4257 ( .A1(n3704), .A2(n3365), .ZN(n3297) );
  NAND2_X1 U4258 ( .A1(n4196), .A2(n3249), .ZN(n3298) );
  NAND2_X1 U4259 ( .A1(n4689), .A2(n4357), .ZN(n4358) );
  NAND2_X1 U4260 ( .A1(n4358), .A2(n5493), .ZN(n3301) );
  XNOR2_X1 U4261 ( .A(n6975), .B(STATE_REG_1__SCAN_IN), .ZN(n4055) );
  NOR2_X1 U4262 ( .A1(n4357), .A2(n4055), .ZN(n3309) );
  INV_X1 U4263 ( .A(n3309), .ZN(n3300) );
  AOI21_X1 U4264 ( .B1(n3301), .B2(n3300), .A(n4359), .ZN(n3302) );
  NAND4_X1 U4265 ( .A1(n3327), .A2(n3328), .A3(n3337), .A4(n3302), .ZN(n3303)
         );
  NAND2_X1 U4266 ( .A1(n4800), .A2(n3304), .ZN(n3305) );
  NAND2_X1 U4267 ( .A1(n3307), .A2(n3306), .ZN(n4321) );
  NAND2_X1 U4268 ( .A1(n3136), .A2(n4662), .ZN(n3308) );
  NOR2_X2 U4269 ( .A1(n3308), .A2(n5493), .ZN(n4701) );
  NAND2_X1 U4270 ( .A1(n4701), .A2(n3146), .ZN(n4563) );
  NAND2_X1 U4271 ( .A1(n4564), .A2(n4705), .ZN(n4360) );
  OR2_X2 U4272 ( .A1(n4563), .A2(n4360), .ZN(n4355) );
  INV_X1 U4273 ( .A(n3310), .ZN(n3313) );
  NAND2_X1 U4274 ( .A1(n4198), .A2(n4689), .ZN(n3311) );
  NAND2_X1 U4275 ( .A1(n3892), .A2(n4683), .ZN(n4329) );
  NAND2_X1 U4276 ( .A1(n3313), .A2(n4329), .ZN(n3314) );
  NAND2_X1 U4277 ( .A1(n3314), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3316) );
  XNOR2_X1 U4278 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5384) );
  OAI22_X1 U4279 ( .A1(n6728), .A2(n5384), .B1(n4565), .B2(n6579), .ZN(n3317)
         );
  INV_X1 U4280 ( .A(n3317), .ZN(n3315) );
  INV_X1 U4281 ( .A(n3316), .ZN(n3318) );
  NAND2_X1 U4282 ( .A1(n3318), .A2(n3158), .ZN(n3319) );
  INV_X1 U4283 ( .A(n3320), .ZN(n3343) );
  NAND2_X1 U4284 ( .A1(n3343), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3325) );
  INV_X1 U4285 ( .A(n4565), .ZN(n3322) );
  INV_X1 U4286 ( .A(n6728), .ZN(n3321) );
  MUX2_X1 U4287 ( .A(n3322), .B(n3321), .S(n4838), .Z(n3323) );
  INV_X1 U4288 ( .A(n3323), .ZN(n3324) );
  INV_X1 U4289 ( .A(n4358), .ZN(n5295) );
  AOI22_X1 U4290 ( .A1(n5295), .A2(n3294), .B1(n3962), .B2(n4361), .ZN(n3326)
         );
  AND2_X1 U4291 ( .A1(n3327), .A2(n3326), .ZN(n4368) );
  INV_X1 U4292 ( .A(n3328), .ZN(n3336) );
  NAND2_X1 U4293 ( .A1(n3329), .A2(n4456), .ZN(n3334) );
  NAND3_X1 U4294 ( .A1(n4662), .A2(n4805), .A3(n3249), .ZN(n3332) );
  NAND2_X1 U4295 ( .A1(n3136), .A2(n4705), .ZN(n3331) );
  OR2_X1 U4296 ( .A1(n6715), .A2(n6609), .ZN(n6611) );
  INV_X1 U4297 ( .A(n6611), .ZN(n3333) );
  NAND3_X1 U4298 ( .A1(n3334), .A2(n4617), .A3(n3333), .ZN(n3335) );
  NOR2_X1 U4299 ( .A1(n3336), .A2(n3335), .ZN(n3340) );
  INV_X1 U4300 ( .A(n3337), .ZN(n3338) );
  OAI21_X1 U4301 ( .B1(n3338), .B2(n3136), .A(n4357), .ZN(n3339) );
  NAND3_X1 U4302 ( .A1(n4368), .A2(n3340), .A3(n3339), .ZN(n3385) );
  NAND2_X1 U4303 ( .A1(n3370), .A2(n3388), .ZN(n3342) );
  NAND2_X1 U4304 ( .A1(n3342), .A2(n3341), .ZN(n3349) );
  AND2_X1 U4305 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3344) );
  NAND2_X1 U4306 ( .A1(n3344), .A2(n6586), .ZN(n6502) );
  INV_X1 U4307 ( .A(n3344), .ZN(n3345) );
  NAND2_X1 U4308 ( .A1(n3345), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3346) );
  OAI22_X1 U4309 ( .A1(n4711), .A2(n6728), .B1(n4565), .B2(n6586), .ZN(n3347)
         );
  OR2_X2 U4310 ( .A1(n3349), .A2(n3348), .ZN(n3467) );
  NAND2_X1 U4311 ( .A1(n3349), .A2(n3348), .ZN(n3350) );
  AOI22_X1 U4312 ( .A1(n4163), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3356) );
  INV_X1 U4313 ( .A(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n7023) );
  AOI22_X1 U4314 ( .A1(n4174), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3355) );
  INV_X1 U4315 ( .A(n3352), .ZN(n3474) );
  AOI22_X1 U4316 ( .A1(n4171), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3354) );
  AOI22_X1 U4317 ( .A1(n4173), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3353) );
  NAND4_X1 U4318 ( .A1(n3356), .A2(n3355), .A3(n3354), .A4(n3353), .ZN(n3364)
         );
  AOI22_X1 U4319 ( .A1(n4084), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4166), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3362) );
  AOI22_X1 U4320 ( .A1(n3137), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3361) );
  AOI22_X1 U4321 ( .A1(n4146), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3155), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4322 ( .A1(n4165), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3359) );
  NAND4_X1 U4323 ( .A1(n3362), .A2(n3361), .A3(n3360), .A4(n3359), .ZN(n3363)
         );
  INV_X1 U4324 ( .A(n3473), .ZN(n3367) );
  AOI22_X1 U4325 ( .A1(n3916), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3367), 
        .B2(n3366), .ZN(n3368) );
  INV_X1 U4326 ( .A(n3433), .ZN(n3432) );
  INV_X1 U4327 ( .A(n3388), .ZN(n3372) );
  INV_X1 U4328 ( .A(n3370), .ZN(n3371) );
  AOI22_X1 U4329 ( .A1(n4084), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4163), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U4330 ( .A1(n3137), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3375) );
  AOI22_X1 U4331 ( .A1(n3139), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3144), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4332 ( .A1(n4172), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3373) );
  NAND4_X1 U4333 ( .A1(n3376), .A2(n3375), .A3(n3374), .A4(n3373), .ZN(n3382)
         );
  AOI22_X1 U4334 ( .A1(n4165), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4161), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3380) );
  AOI22_X1 U4335 ( .A1(n4166), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3379) );
  AOI22_X1 U4336 ( .A1(n4173), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4337 ( .A1(n4174), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3377) );
  NAND4_X1 U4338 ( .A1(n3380), .A2(n3379), .A3(n3378), .A4(n3377), .ZN(n3381)
         );
  NOR2_X1 U4339 ( .A1(n4699), .A2(n3425), .ZN(n3383) );
  INV_X1 U4340 ( .A(n3384), .ZN(n3387) );
  INV_X1 U4341 ( .A(n3385), .ZN(n3386) );
  NAND2_X1 U4342 ( .A1(n3387), .A2(n3386), .ZN(n3389) );
  NAND2_X1 U4343 ( .A1(n3389), .A2(n3388), .ZN(n3449) );
  AOI22_X1 U4344 ( .A1(n3137), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4166), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4345 ( .A1(n4146), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3393) );
  AOI22_X1 U4346 ( .A1(n4172), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3392) );
  BUF_X1 U4347 ( .A(n4174), .Z(n4120) );
  AOI22_X1 U4348 ( .A1(n4120), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3391) );
  NAND4_X1 U4349 ( .A1(n3394), .A2(n3393), .A3(n3392), .A4(n3391), .ZN(n3400)
         );
  AOI22_X1 U4350 ( .A1(n4165), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3480), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3398) );
  AOI22_X1 U4351 ( .A1(n3138), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4164), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3397) );
  AOI22_X1 U4352 ( .A1(n4173), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3357), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3396) );
  AOI22_X1 U4353 ( .A1(n4163), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3395) );
  NAND4_X1 U4354 ( .A1(n3398), .A2(n3397), .A3(n3396), .A4(n3395), .ZN(n3399)
         );
  NOR2_X1 U4355 ( .A1(n4699), .A2(n4275), .ZN(n3422) );
  AOI22_X1 U4356 ( .A1(n4120), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4166), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3405) );
  AOI22_X1 U4357 ( .A1(n3137), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3404) );
  AOI22_X1 U4358 ( .A1(n4165), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4164), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3403) );
  AOI22_X1 U4359 ( .A1(n4163), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3402) );
  NAND4_X1 U4360 ( .A1(n3405), .A2(n3404), .A3(n3403), .A4(n3402), .ZN(n3414)
         );
  AOI22_X1 U4361 ( .A1(n4141), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3412) );
  AOI22_X1 U4362 ( .A1(n4146), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3411) );
  AOI22_X1 U4363 ( .A1(n3133), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3410) );
  AOI22_X1 U4364 ( .A1(n3155), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3409) );
  NAND4_X1 U4365 ( .A1(n3412), .A2(n3411), .A3(n3410), .A4(n3409), .ZN(n3413)
         );
  INV_X1 U4366 ( .A(n4218), .ZN(n3415) );
  MUX2_X1 U4367 ( .A(n3422), .B(n3420), .S(n3415), .Z(n3416) );
  INV_X1 U4368 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3419) );
  AOI21_X1 U4369 ( .B1(n3365), .B2(n4275), .A(n6609), .ZN(n3418) );
  NAND2_X1 U4370 ( .A1(n4689), .A2(n4218), .ZN(n3417) );
  OAI211_X1 U4371 ( .C1(n3944), .C2(n3419), .A(n3418), .B(n3417), .ZN(n3446)
         );
  NAND2_X1 U4372 ( .A1(n3447), .A2(n3446), .ZN(n3421) );
  INV_X1 U4373 ( .A(n3420), .ZN(n4207) );
  INV_X1 U4374 ( .A(n3422), .ZN(n3424) );
  NAND2_X1 U4375 ( .A1(n3916), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3423) );
  OAI211_X1 U4376 ( .C1(n3425), .C2(n3473), .A(n3424), .B(n3423), .ZN(n3427)
         );
  NAND2_X1 U4377 ( .A1(n3439), .A2(n3427), .ZN(n3426) );
  NAND2_X1 U4378 ( .A1(n3440), .A2(n3426), .ZN(n3430) );
  INV_X1 U4379 ( .A(n3439), .ZN(n3428) );
  INV_X1 U4380 ( .A(n3427), .ZN(n3438) );
  NAND2_X1 U4381 ( .A1(n3428), .A2(n3438), .ZN(n3429) );
  INV_X1 U4382 ( .A(n3434), .ZN(n3431) );
  NAND2_X1 U4383 ( .A1(n3432), .A2(n3431), .ZN(n3435) );
  NAND2_X1 U4384 ( .A1(n3434), .A2(n3433), .ZN(n3466) );
  BUF_X2 U4385 ( .A(n3466), .Z(n3491) );
  NAND2_X1 U4386 ( .A1(n3435), .A2(n3491), .ZN(n4639) );
  INV_X1 U4387 ( .A(n4639), .ZN(n3436) );
  NAND2_X1 U4388 ( .A1(n3436), .A2(n3695), .ZN(n3437) );
  NAND2_X1 U4389 ( .A1(n6935), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3861) );
  NAND2_X1 U4390 ( .A1(n3437), .A2(n3861), .ZN(n4577) );
  NAND2_X1 U4391 ( .A1(n4216), .A2(n3695), .ZN(n3445) );
  AOI22_X1 U4392 ( .A1(n4193), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6935), .ZN(n3443) );
  INV_X1 U4393 ( .A(n4360), .ZN(n5495) );
  NAND2_X1 U4394 ( .A1(n3493), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3442) );
  AND2_X1 U4395 ( .A1(n3443), .A2(n3442), .ZN(n3444) );
  AOI21_X1 U4396 ( .B1(n5379), .B2(n4805), .A(n6935), .ZN(n4581) );
  OR2_X1 U4397 ( .A1(n5297), .A2(n3648), .ZN(n3453) );
  AOI22_X1 U4398 ( .A1(n4193), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6935), .ZN(n3451) );
  NAND2_X1 U4399 ( .A1(n3493), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3450) );
  AND2_X1 U4400 ( .A1(n3451), .A2(n3450), .ZN(n3452) );
  NAND2_X1 U4401 ( .A1(n3453), .A2(n3452), .ZN(n4580) );
  NAND2_X1 U4402 ( .A1(n4581), .A2(n4580), .ZN(n4579) );
  INV_X1 U4403 ( .A(n4580), .ZN(n3454) );
  NAND2_X1 U4404 ( .A1(n3454), .A2(n4185), .ZN(n3455) );
  NAND2_X1 U4405 ( .A1(n4579), .A2(n3455), .ZN(n4540) );
  NAND2_X1 U4406 ( .A1(n3493), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3460) );
  OAI21_X1 U4407 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3494), .ZN(n6351) );
  NAND2_X1 U4408 ( .A1(n6351), .A2(n4185), .ZN(n3457) );
  NAND2_X1 U4409 ( .A1(n4192), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3456)
         );
  NAND2_X1 U4410 ( .A1(n3457), .A2(n3456), .ZN(n3458) );
  AOI21_X1 U4411 ( .B1(n4193), .B2(EAX_REG_2__SCAN_IN), .A(n3458), .ZN(n3459)
         );
  AND2_X1 U4412 ( .A1(n3460), .A2(n3459), .ZN(n3461) );
  NAND2_X1 U4413 ( .A1(n4577), .A2(n4576), .ZN(n3465) );
  INV_X1 U4414 ( .A(n4539), .ZN(n3463) );
  INV_X1 U4415 ( .A(n3461), .ZN(n3462) );
  NAND2_X1 U4416 ( .A1(n3463), .A2(n3462), .ZN(n3464) );
  INV_X1 U4417 ( .A(n3466), .ZN(n3489) );
  NAND2_X1 U4418 ( .A1(n3343), .A2(n6988), .ZN(n3472) );
  NAND3_X1 U4419 ( .A1(n7014), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6441) );
  INV_X1 U4420 ( .A(n6441), .ZN(n3468) );
  NAND2_X1 U4421 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3468), .ZN(n5041) );
  NAND2_X1 U4422 ( .A1(n7014), .A2(n5041), .ZN(n3469) );
  NAND3_X1 U4423 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5110) );
  INV_X1 U4424 ( .A(n5110), .ZN(n4960) );
  NAND2_X1 U4425 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4960), .ZN(n4955) );
  NAND2_X1 U4426 ( .A1(n3469), .A2(n4955), .ZN(n4710) );
  OAI22_X1 U4427 ( .A1(n6728), .A2(n4710), .B1(n4565), .B2(n7014), .ZN(n3470)
         );
  INV_X1 U4428 ( .A(n3470), .ZN(n3471) );
  NAND2_X1 U4429 ( .A1(n4585), .A2(n6609), .ZN(n3488) );
  AOI22_X1 U4430 ( .A1(n4163), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3479) );
  AOI22_X1 U4431 ( .A1(n4120), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3478) );
  AOI22_X1 U4432 ( .A1(n4171), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3477) );
  AOI22_X1 U4433 ( .A1(n4173), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3476) );
  NAND4_X1 U4434 ( .A1(n3479), .A2(n3478), .A3(n3477), .A4(n3476), .ZN(n3486)
         );
  AOI22_X1 U4435 ( .A1(n4084), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4166), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3484) );
  AOI22_X1 U4436 ( .A1(n3137), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3483) );
  AOI22_X1 U4437 ( .A1(n4146), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3155), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3482) );
  AOI22_X1 U4438 ( .A1(n4165), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3481) );
  NAND4_X1 U4439 ( .A1(n3484), .A2(n3483), .A3(n3482), .A4(n3481), .ZN(n3485)
         );
  AOI22_X1 U4440 ( .A1(n3135), .A2(n4210), .B1(INSTQUEUE_REG_0__3__SCAN_IN), 
        .B2(n3916), .ZN(n3487) );
  NAND2_X1 U4441 ( .A1(n3491), .A2(n4642), .ZN(n3492) );
  NAND2_X1 U4442 ( .A1(n3515), .A2(n3492), .ZN(n4638) );
  INV_X1 U4443 ( .A(n3493), .ZN(n3520) );
  INV_X1 U4444 ( .A(n6988), .ZN(n4592) );
  OAI21_X1 U4445 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3495), .A(n3521), 
        .ZN(n6259) );
  AOI22_X1 U4446 ( .A1(n6259), .A2(n4185), .B1(n4192), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3497) );
  NAND2_X1 U4447 ( .A1(n4193), .A2(EAX_REG_3__SCAN_IN), .ZN(n3496) );
  OAI211_X1 U4448 ( .C1(n3520), .C2(n4592), .A(n3497), .B(n3496), .ZN(n3498)
         );
  INV_X1 U4449 ( .A(n3498), .ZN(n3499) );
  OAI21_X1 U4450 ( .B1(n4638), .B2(n3648), .A(n3499), .ZN(n4553) );
  INV_X1 U4451 ( .A(n3515), .ZN(n3512) );
  AOI22_X1 U4452 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4163), .B1(n3407), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3503) );
  AOI22_X1 U4453 ( .A1(n3137), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3502) );
  AOI22_X1 U4454 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n4173), .B1(n4172), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3501) );
  AOI22_X1 U4455 ( .A1(n4120), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3500) );
  NAND4_X1 U4456 ( .A1(n3503), .A2(n3502), .A3(n3501), .A4(n3500), .ZN(n3509)
         );
  AOI22_X1 U4457 ( .A1(n4165), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3155), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3507) );
  AOI22_X1 U4458 ( .A1(n4146), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3506) );
  AOI22_X1 U4459 ( .A1(n4084), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3505) );
  AOI22_X1 U4460 ( .A1(n4166), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3504) );
  NAND4_X1 U4461 ( .A1(n3507), .A2(n3506), .A3(n3505), .A4(n3504), .ZN(n3508)
         );
  NAND2_X1 U4462 ( .A1(n3135), .A2(n4247), .ZN(n3511) );
  NAND2_X1 U4463 ( .A1(n3916), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3510) );
  NAND2_X1 U4464 ( .A1(n3511), .A2(n3510), .ZN(n3513) );
  INV_X1 U4465 ( .A(n3513), .ZN(n3514) );
  NAND2_X1 U4466 ( .A1(n3515), .A2(n3514), .ZN(n3516) );
  NAND2_X1 U4467 ( .A1(n3539), .A2(n3516), .ZN(n4241) );
  INV_X1 U4468 ( .A(n4241), .ZN(n3517) );
  INV_X1 U4469 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6121) );
  OAI21_X1 U4470 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n6121), .A(n6935), 
        .ZN(n3519) );
  NAND2_X1 U4471 ( .A1(n4193), .A2(EAX_REG_4__SCAN_IN), .ZN(n3518) );
  OAI211_X1 U4472 ( .C1(n3520), .C2(n6113), .A(n3519), .B(n3518), .ZN(n3523)
         );
  AOI21_X1 U4473 ( .B1(n6774), .B2(n3521), .A(n3541), .ZN(n6240) );
  NAND2_X1 U4474 ( .A1(n6240), .A2(n4185), .ZN(n3522) );
  NAND2_X1 U4475 ( .A1(n3523), .A2(n3522), .ZN(n3524) );
  NAND2_X1 U4476 ( .A1(n3525), .A2(n3524), .ZN(n4574) );
  INV_X1 U4477 ( .A(n3539), .ZN(n3537) );
  AOI22_X1 U4478 ( .A1(n4163), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3529) );
  AOI22_X1 U4479 ( .A1(n4120), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3528) );
  AOI22_X1 U4480 ( .A1(n4171), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3527) );
  AOI22_X1 U4481 ( .A1(n4173), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3526) );
  NAND4_X1 U4482 ( .A1(n3529), .A2(n3528), .A3(n3527), .A4(n3526), .ZN(n3535)
         );
  AOI22_X1 U4483 ( .A1(n4084), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4166), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3533) );
  AOI22_X1 U4484 ( .A1(n3137), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3532) );
  INV_X1 U4485 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n6980) );
  AOI22_X1 U4486 ( .A1(n4146), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3531) );
  AOI22_X1 U4487 ( .A1(n4165), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3530) );
  NAND4_X1 U4488 ( .A1(n3533), .A2(n3532), .A3(n3531), .A4(n3530), .ZN(n3534)
         );
  AOI22_X1 U4489 ( .A1(n3135), .A2(n4250), .B1(INSTQUEUE_REG_0__5__SCAN_IN), 
        .B2(n3916), .ZN(n3538) );
  NAND2_X1 U4490 ( .A1(n3537), .A2(n3536), .ZN(n3560) );
  NAND2_X1 U4491 ( .A1(n3539), .A2(n3538), .ZN(n3540) );
  NAND2_X1 U4492 ( .A1(n3560), .A2(n3540), .ZN(n4245) );
  AOI22_X1 U4493 ( .A1(n4193), .A2(EAX_REG_5__SCAN_IN), .B1(n4192), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3543) );
  OAI21_X1 U4494 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n3541), .A(n3554), 
        .ZN(n6232) );
  NAND2_X1 U4495 ( .A1(n6232), .A2(n4185), .ZN(n3542) );
  OAI211_X1 U4496 ( .C1(n4245), .C2(n3648), .A(n3543), .B(n3542), .ZN(n4582)
         );
  AOI22_X1 U4497 ( .A1(n4165), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3547) );
  AOI22_X1 U4498 ( .A1(n4146), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4163), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3546) );
  AOI22_X1 U4499 ( .A1(n4084), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3545) );
  AOI22_X1 U4500 ( .A1(n4171), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3544) );
  NAND4_X1 U4501 ( .A1(n3547), .A2(n3546), .A3(n3545), .A4(n3544), .ZN(n3553)
         );
  AOI22_X1 U4502 ( .A1(n4166), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3551) );
  AOI22_X1 U4503 ( .A1(n3407), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4504 ( .A1(n3138), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U4505 ( .A1(n4120), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3548) );
  NAND4_X1 U4506 ( .A1(n3551), .A2(n3550), .A3(n3549), .A4(n3548), .ZN(n3552)
         );
  AOI22_X1 U4507 ( .A1(n3135), .A2(n4266), .B1(n3916), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3561) );
  NAND2_X1 U4508 ( .A1(n3560), .A2(n3561), .ZN(n4257) );
  NAND2_X1 U4509 ( .A1(n4193), .A2(EAX_REG_6__SCAN_IN), .ZN(n3558) );
  NAND2_X1 U4510 ( .A1(n3554), .A2(n6890), .ZN(n3556) );
  INV_X1 U4511 ( .A(n3566), .ZN(n3555) );
  NAND2_X1 U4512 ( .A1(n3556), .A2(n3555), .ZN(n6335) );
  NAND2_X1 U4513 ( .A1(n6335), .A2(n4185), .ZN(n3557) );
  OAI211_X1 U4514 ( .C1(n3861), .C2(n6890), .A(n3558), .B(n3557), .ZN(n3559)
         );
  INV_X1 U4515 ( .A(n3560), .ZN(n3563) );
  INV_X1 U4516 ( .A(n3561), .ZN(n3562) );
  INV_X1 U4517 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n6986) );
  NAND2_X1 U4518 ( .A1(n3135), .A2(n4275), .ZN(n3564) );
  OAI21_X1 U4519 ( .B1(n6986), .B2(n3944), .A(n3564), .ZN(n3565) );
  XNOR2_X1 U4520 ( .A(n4206), .B(n3565), .ZN(n4264) );
  NAND2_X1 U4521 ( .A1(n4264), .A2(n3695), .ZN(n3572) );
  OAI21_X1 U4522 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n3566), .A(n3573), 
        .ZN(n6214) );
  INV_X1 U4523 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3569) );
  INV_X1 U4524 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3568) );
  OAI22_X1 U4525 ( .A1(n4154), .A2(n3569), .B1(n3861), .B2(n3568), .ZN(n3570)
         );
  AOI21_X1 U4526 ( .B1(n6214), .B2(n4185), .A(n3570), .ZN(n3571) );
  NAND2_X1 U4527 ( .A1(n3572), .A2(n3571), .ZN(n5046) );
  NAND2_X1 U4528 ( .A1(n4950), .A2(n5046), .ZN(n5047) );
  INV_X1 U4529 ( .A(n5047), .ZN(n3590) );
  AOI21_X1 U4530 ( .B1(n3573), .B2(n6977), .A(n3606), .ZN(n6195) );
  OR2_X1 U4531 ( .A1(n6195), .A2(n4191), .ZN(n3588) );
  AOI22_X1 U4532 ( .A1(n4165), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3577) );
  AOI22_X1 U4533 ( .A1(n4120), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3576) );
  AOI22_X1 U4534 ( .A1(n4084), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3575) );
  AOI22_X1 U4535 ( .A1(n4166), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3574) );
  NAND4_X1 U4536 ( .A1(n3577), .A2(n3576), .A3(n3575), .A4(n3574), .ZN(n3583)
         );
  AOI22_X1 U4537 ( .A1(n3137), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4538 ( .A1(n4146), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4539 ( .A1(n4163), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3579) );
  AOI22_X1 U4540 ( .A1(n4173), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3578) );
  NAND4_X1 U4541 ( .A1(n3581), .A2(n3580), .A3(n3579), .A4(n3578), .ZN(n3582)
         );
  OAI21_X1 U4542 ( .B1(n3583), .B2(n3582), .A(n3695), .ZN(n3586) );
  NAND2_X1 U4543 ( .A1(n3567), .A2(EAX_REG_8__SCAN_IN), .ZN(n3585) );
  NAND2_X1 U4544 ( .A1(n4192), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3584)
         );
  NAND2_X1 U4545 ( .A1(n3590), .A2(n3589), .ZN(n5182) );
  XNOR2_X1 U4546 ( .A(n3606), .B(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5317) );
  AOI22_X1 U4547 ( .A1(n3137), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3594) );
  AOI22_X1 U4548 ( .A1(n4120), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3593) );
  AOI22_X1 U4549 ( .A1(n4165), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3592) );
  AOI22_X1 U4550 ( .A1(n4163), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3591) );
  NAND4_X1 U4551 ( .A1(n3594), .A2(n3593), .A3(n3592), .A4(n3591), .ZN(n3600)
         );
  AOI22_X1 U4552 ( .A1(n4166), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4161), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4553 ( .A1(n4084), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4554 ( .A1(n4173), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4555 ( .A1(n4172), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3595) );
  NAND4_X1 U4556 ( .A1(n3598), .A2(n3597), .A3(n3596), .A4(n3595), .ZN(n3599)
         );
  OAI21_X1 U4557 ( .B1(n3600), .B2(n3599), .A(n3695), .ZN(n3603) );
  NAND2_X1 U4558 ( .A1(n3567), .A2(EAX_REG_9__SCAN_IN), .ZN(n3602) );
  NAND2_X1 U4559 ( .A1(n4192), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3601)
         );
  NAND3_X1 U4560 ( .A1(n3603), .A2(n3602), .A3(n3601), .ZN(n3604) );
  AOI21_X1 U4561 ( .B1(n5317), .B2(n4185), .A(n3604), .ZN(n5181) );
  NAND2_X1 U4562 ( .A1(n5280), .A2(n3605), .ZN(n5312) );
  XOR2_X1 U4563 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3631), .Z(n6187) );
  INV_X1 U4564 ( .A(n6187), .ZN(n5337) );
  AOI22_X1 U4565 ( .A1(n4166), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3610) );
  AOI22_X1 U4566 ( .A1(n4173), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3609) );
  AOI22_X1 U4567 ( .A1(n4163), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3608) );
  AOI22_X1 U4568 ( .A1(n3138), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3607) );
  NAND4_X1 U4569 ( .A1(n3610), .A2(n3609), .A3(n3608), .A4(n3607), .ZN(n3616)
         );
  AOI22_X1 U4570 ( .A1(n4165), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4571 ( .A1(n4084), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4161), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3613) );
  AOI22_X1 U4572 ( .A1(n4172), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4573 ( .A1(n4120), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3611) );
  NAND4_X1 U4574 ( .A1(n3614), .A2(n3613), .A3(n3612), .A4(n3611), .ZN(n3615)
         );
  OAI21_X1 U4575 ( .B1(n3616), .B2(n3615), .A(n3695), .ZN(n3619) );
  NAND2_X1 U4576 ( .A1(n3567), .A2(EAX_REG_10__SCAN_IN), .ZN(n3618) );
  NAND2_X1 U4577 ( .A1(n4192), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3617)
         );
  NAND3_X1 U4578 ( .A1(n3619), .A2(n3618), .A3(n3617), .ZN(n3620) );
  AOI21_X1 U4579 ( .B1(n5337), .B2(n4185), .A(n3620), .ZN(n5311) );
  NOR2_X2 U4580 ( .A1(n5312), .A2(n5311), .ZN(n5302) );
  AOI22_X1 U4581 ( .A1(n4084), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4582 ( .A1(n4146), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3623) );
  AOI22_X1 U4583 ( .A1(n4165), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4584 ( .A1(n4172), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3621) );
  NAND4_X1 U4585 ( .A1(n3624), .A2(n3623), .A3(n3622), .A4(n3621), .ZN(n3630)
         );
  AOI22_X1 U4586 ( .A1(n4166), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4163), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3628) );
  AOI22_X1 U4587 ( .A1(n4120), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3627) );
  AOI22_X1 U4588 ( .A1(n4171), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4589 ( .A1(n3407), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3625) );
  NAND4_X1 U4590 ( .A1(n3628), .A2(n3627), .A3(n3626), .A4(n3625), .ZN(n3629)
         );
  NOR2_X1 U4591 ( .A1(n3630), .A2(n3629), .ZN(n3634) );
  XNOR2_X1 U4592 ( .A(n3635), .B(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5741)
         );
  NAND2_X1 U4593 ( .A1(n5741), .A2(n4185), .ZN(n3633) );
  AOI22_X1 U4594 ( .A1(n4193), .A2(EAX_REG_11__SCAN_IN), .B1(n4192), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3632) );
  OAI211_X1 U4595 ( .C1(n3634), .C2(n3648), .A(n3633), .B(n3632), .ZN(n5306)
         );
  NAND2_X1 U4596 ( .A1(n5302), .A2(n5306), .ZN(n5304) );
  INV_X1 U4597 ( .A(n5304), .ZN(n3653) );
  XOR2_X1 U4598 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3654), .Z(n6169) );
  NAND2_X1 U4599 ( .A1(n6169), .A2(n4185), .ZN(n3651) );
  INV_X1 U4600 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5367) );
  OAI21_X1 U4601 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6121), .A(n6935), 
        .ZN(n3636) );
  OAI21_X1 U4602 ( .B1(n4154), .B2(n5367), .A(n3636), .ZN(n3650) );
  AOI22_X1 U4603 ( .A1(n4165), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4604 ( .A1(n3137), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4605 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n4173), .B1(n3138), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3638) );
  AOI22_X1 U4606 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n4171), .B1(n4162), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3637) );
  NAND4_X1 U4607 ( .A1(n3640), .A2(n3639), .A3(n3638), .A4(n3637), .ZN(n3646)
         );
  AOI22_X1 U4608 ( .A1(n4084), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4163), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4609 ( .A1(n4166), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4610 ( .A1(n3357), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4611 ( .A1(n4172), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3641) );
  NAND4_X1 U4612 ( .A1(n3644), .A2(n3643), .A3(n3642), .A4(n3641), .ZN(n3645)
         );
  NOR2_X1 U4613 ( .A1(n3646), .A2(n3645), .ZN(n3647) );
  NOR2_X1 U4614 ( .A1(n3648), .A2(n3647), .ZN(n3649) );
  AOI21_X1 U4615 ( .B1(n3651), .B2(n3650), .A(n3649), .ZN(n5364) );
  NAND2_X1 U4616 ( .A1(n3653), .A2(n3652), .ZN(n5363) );
  NAND2_X1 U4617 ( .A1(n3655), .A2(n6981), .ZN(n3656) );
  NAND2_X1 U4618 ( .A1(n3656), .A2(n3671), .ZN(n6158) );
  AOI22_X1 U4619 ( .A1(n4120), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3660) );
  AOI22_X1 U4620 ( .A1(n4084), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3659) );
  AOI22_X1 U4621 ( .A1(n4173), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4622 ( .A1(n4172), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3657) );
  NAND4_X1 U4623 ( .A1(n3660), .A2(n3659), .A3(n3658), .A4(n3657), .ZN(n3666)
         );
  AOI22_X1 U4624 ( .A1(n4165), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4166), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3664) );
  AOI22_X1 U4625 ( .A1(n4146), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4626 ( .A1(n4163), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U4627 ( .A1(n3138), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3661) );
  NAND4_X1 U4628 ( .A1(n3664), .A2(n3663), .A3(n3662), .A4(n3661), .ZN(n3665)
         );
  OAI21_X1 U4629 ( .B1(n3666), .B2(n3665), .A(n3695), .ZN(n3669) );
  NAND2_X1 U4630 ( .A1(n4193), .A2(EAX_REG_13__SCAN_IN), .ZN(n3668) );
  NAND2_X1 U4631 ( .A1(n4192), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3667)
         );
  NAND3_X1 U4632 ( .A1(n3669), .A2(n3668), .A3(n3667), .ZN(n3670) );
  AOI21_X1 U4633 ( .B1(n6158), .B2(n4185), .A(n3670), .ZN(n5435) );
  NOR2_X2 U4634 ( .A1(n5363), .A2(n5435), .ZN(n5461) );
  AOI21_X1 U4635 ( .B1(n6835), .B2(n3671), .A(n3703), .ZN(n6148) );
  OR2_X1 U4636 ( .A1(n6148), .A2(n4191), .ZN(n3686) );
  AOI22_X1 U4637 ( .A1(n3137), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3675) );
  AOI22_X1 U4638 ( .A1(n4084), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3674) );
  AOI22_X1 U4639 ( .A1(n4165), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3673) );
  AOI22_X1 U4640 ( .A1(n4146), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3672) );
  NAND4_X1 U4641 ( .A1(n3675), .A2(n3674), .A3(n3673), .A4(n3672), .ZN(n3681)
         );
  AOI22_X1 U4642 ( .A1(n4166), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3679) );
  AOI22_X1 U4643 ( .A1(n4120), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3678) );
  AOI22_X1 U4644 ( .A1(n4173), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3677) );
  AOI22_X1 U4645 ( .A1(n4163), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3676) );
  NAND4_X1 U4646 ( .A1(n3679), .A2(n3678), .A3(n3677), .A4(n3676), .ZN(n3680)
         );
  OAI21_X1 U4647 ( .B1(n3681), .B2(n3680), .A(n3695), .ZN(n3684) );
  NAND2_X1 U4648 ( .A1(n4193), .A2(EAX_REG_14__SCAN_IN), .ZN(n3683) );
  NAND2_X1 U4649 ( .A1(n4192), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3682)
         );
  AND3_X1 U4650 ( .A1(n3684), .A2(n3683), .A3(n3682), .ZN(n3685) );
  NAND2_X1 U4651 ( .A1(n3686), .A2(n3685), .ZN(n5460) );
  XNOR2_X1 U4652 ( .A(n3703), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5920)
         );
  AOI22_X1 U4653 ( .A1(n3137), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4161), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4654 ( .A1(n4120), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4655 ( .A1(n4165), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4656 ( .A1(n3407), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3687) );
  NAND4_X1 U4657 ( .A1(n3690), .A2(n3689), .A3(n3688), .A4(n3687), .ZN(n3697)
         );
  AOI22_X1 U4658 ( .A1(n4163), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3694) );
  AOI22_X1 U4659 ( .A1(n4171), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3693) );
  AOI22_X1 U4660 ( .A1(n4166), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4661 ( .A1(n4084), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3691) );
  NAND4_X1 U4662 ( .A1(n3694), .A2(n3693), .A3(n3692), .A4(n3691), .ZN(n3696)
         );
  OAI21_X1 U4663 ( .B1(n3697), .B2(n3696), .A(n3695), .ZN(n3700) );
  NAND2_X1 U4664 ( .A1(n4193), .A2(EAX_REG_15__SCAN_IN), .ZN(n3699) );
  NAND2_X1 U4665 ( .A1(n4192), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3698)
         );
  NAND3_X1 U4666 ( .A1(n3700), .A2(n3699), .A3(n3698), .ZN(n3701) );
  AOI21_X1 U4667 ( .B1(n5920), .B2(n4185), .A(n3701), .ZN(n5729) );
  XOR2_X1 U4668 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3719), .Z(n5913) );
  AOI22_X1 U4669 ( .A1(n4141), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3708) );
  AOI22_X1 U4670 ( .A1(n4165), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4161), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3707) );
  AOI22_X1 U4671 ( .A1(n4120), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4672 ( .A1(n4163), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3705) );
  NAND4_X1 U4673 ( .A1(n3708), .A2(n3707), .A3(n3706), .A4(n3705), .ZN(n3714)
         );
  AOI22_X1 U4674 ( .A1(n3137), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3712) );
  AOI22_X1 U4675 ( .A1(n4171), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3711) );
  AOI22_X1 U4676 ( .A1(n4172), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4677 ( .A1(n4166), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3709) );
  NAND4_X1 U4678 ( .A1(n3712), .A2(n3711), .A3(n3710), .A4(n3709), .ZN(n3713)
         );
  NOR2_X1 U4679 ( .A1(n3714), .A2(n3713), .ZN(n3716) );
  AOI22_X1 U4680 ( .A1(n4193), .A2(EAX_REG_16__SCAN_IN), .B1(n4192), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3715) );
  OAI21_X1 U4681 ( .B1(n4188), .B2(n3716), .A(n3715), .ZN(n3717) );
  AOI21_X1 U4682 ( .B1(n5913), .B2(n4185), .A(n3717), .ZN(n5711) );
  INV_X1 U4683 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3720) );
  XNOR2_X1 U4684 ( .A(n3735), .B(n3720), .ZN(n5907) );
  AOI22_X1 U4685 ( .A1(n4165), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4686 ( .A1(n4120), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4687 ( .A1(n4166), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4688 ( .A1(n4173), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3721) );
  NAND4_X1 U4689 ( .A1(n3724), .A2(n3723), .A3(n3722), .A4(n3721), .ZN(n3730)
         );
  AOI22_X1 U4690 ( .A1(n4146), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3728) );
  AOI22_X1 U4691 ( .A1(n4172), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3727) );
  AOI22_X1 U4692 ( .A1(n4141), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4693 ( .A1(n4163), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3725) );
  NAND4_X1 U4694 ( .A1(n3728), .A2(n3727), .A3(n3726), .A4(n3725), .ZN(n3729)
         );
  NOR2_X1 U4695 ( .A1(n3730), .A2(n3729), .ZN(n3731) );
  NOR2_X1 U4696 ( .A1(n4188), .A2(n3731), .ZN(n3734) );
  INV_X1 U4697 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4513) );
  NAND2_X1 U4698 ( .A1(n6935), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3732)
         );
  OAI211_X1 U4699 ( .C1(n4154), .C2(n4513), .A(n4191), .B(n3732), .ZN(n3733)
         );
  OAI22_X1 U4700 ( .A1(n5907), .A2(n4191), .B1(n3734), .B2(n3733), .ZN(n5699)
         );
  NOR2_X2 U4701 ( .A1(n5697), .A2(n5699), .ZN(n5698) );
  OR2_X1 U4702 ( .A1(n3736), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3737)
         );
  NAND2_X1 U4703 ( .A1(n3737), .A2(n3768), .ZN(n6138) );
  INV_X1 U4704 ( .A(n6138), .ZN(n3752) );
  AOI22_X1 U4705 ( .A1(n4141), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3741) );
  AOI22_X1 U4706 ( .A1(n4146), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4707 ( .A1(n4165), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4708 ( .A1(n4172), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3738) );
  NAND4_X1 U4709 ( .A1(n3741), .A2(n3740), .A3(n3739), .A4(n3738), .ZN(n3747)
         );
  AOI22_X1 U4710 ( .A1(n4166), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4163), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3745) );
  AOI22_X1 U4711 ( .A1(n4120), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3744) );
  AOI22_X1 U4712 ( .A1(n4171), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U4713 ( .A1(n3407), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3742) );
  NAND4_X1 U4714 ( .A1(n3745), .A2(n3744), .A3(n3743), .A4(n3742), .ZN(n3746)
         );
  OR2_X1 U4715 ( .A1(n3747), .A2(n3746), .ZN(n3750) );
  INV_X1 U4716 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4506) );
  NAND2_X1 U4717 ( .A1(n6935), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3748)
         );
  OAI211_X1 U4718 ( .C1(n4154), .C2(n4506), .A(n4191), .B(n3748), .ZN(n3749)
         );
  AOI21_X1 U4719 ( .B1(n4156), .B2(n3750), .A(n3749), .ZN(n3751) );
  AOI21_X1 U4720 ( .B1(n3752), .B2(n4185), .A(n3751), .ZN(n5797) );
  NAND2_X1 U4721 ( .A1(n5698), .A2(n5797), .ZN(n5799) );
  AOI22_X1 U4722 ( .A1(n4163), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4723 ( .A1(n4120), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4724 ( .A1(n4171), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3754) );
  AOI22_X1 U4725 ( .A1(n4173), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3753) );
  NAND4_X1 U4726 ( .A1(n3756), .A2(n3755), .A3(n3754), .A4(n3753), .ZN(n3762)
         );
  AOI22_X1 U4727 ( .A1(n4141), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4166), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4728 ( .A1(n3137), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3759) );
  AOI22_X1 U4729 ( .A1(n4146), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3758) );
  AOI22_X1 U4730 ( .A1(n4165), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3757) );
  NAND4_X1 U4731 ( .A1(n3760), .A2(n3759), .A3(n3758), .A4(n3757), .ZN(n3761)
         );
  NOR2_X1 U4732 ( .A1(n3762), .A2(n3761), .ZN(n3765) );
  INV_X1 U4733 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5898) );
  AOI21_X1 U4734 ( .B1(n5898), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3763) );
  AOI21_X1 U4735 ( .B1(n3567), .B2(EAX_REG_19__SCAN_IN), .A(n3763), .ZN(n3764)
         );
  OAI21_X1 U4736 ( .B1(n4188), .B2(n3765), .A(n3764), .ZN(n3767) );
  XNOR2_X1 U4737 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n3768), .ZN(n6028)
         );
  NAND2_X1 U4738 ( .A1(n6028), .A2(n4185), .ZN(n3766) );
  NAND2_X1 U4739 ( .A1(n5786), .A2(n3160), .ZN(n5785) );
  OR2_X1 U4740 ( .A1(n3769), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3770)
         );
  NAND2_X1 U4741 ( .A1(n3770), .A2(n3814), .ZN(n6058) );
  AOI22_X1 U4742 ( .A1(n4141), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4163), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4743 ( .A1(n4166), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4744 ( .A1(n3138), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4745 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4172), .B1(n4162), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3771) );
  NAND4_X1 U4746 ( .A1(n3774), .A2(n3773), .A3(n3772), .A4(n3771), .ZN(n3780)
         );
  AOI22_X1 U4747 ( .A1(n3137), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4748 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n4173), .B1(n4171), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4749 ( .A1(n4165), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4750 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4120), .B1(n3139), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3775) );
  NAND4_X1 U4751 ( .A1(n3778), .A2(n3777), .A3(n3776), .A4(n3775), .ZN(n3779)
         );
  NOR2_X1 U4752 ( .A1(n3780), .A2(n3779), .ZN(n3781) );
  NOR2_X1 U4753 ( .A1(n4188), .A2(n3781), .ZN(n3784) );
  INV_X1 U4754 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4504) );
  NAND2_X1 U4755 ( .A1(n6935), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3782)
         );
  OAI211_X1 U4756 ( .C1(n4154), .C2(n4504), .A(n4191), .B(n3782), .ZN(n3783)
         );
  OAI22_X1 U4757 ( .A1(n6058), .A2(n4191), .B1(n3784), .B2(n3783), .ZN(n5778)
         );
  NOR2_X2 U4758 ( .A1(n5785), .A2(n5778), .ZN(n5666) );
  AOI22_X1 U4759 ( .A1(n3137), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4760 ( .A1(n4141), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4163), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4761 ( .A1(n4120), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4762 ( .A1(n3139), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3785) );
  NAND4_X1 U4763 ( .A1(n3788), .A2(n3787), .A3(n3786), .A4(n3785), .ZN(n3794)
         );
  AOI22_X1 U4764 ( .A1(n4166), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4765 ( .A1(n4165), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4766 ( .A1(n3138), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4767 ( .A1(n4173), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3789) );
  NAND4_X1 U4768 ( .A1(n3792), .A2(n3791), .A3(n3790), .A4(n3789), .ZN(n3793)
         );
  NOR2_X1 U4769 ( .A1(n3794), .A2(n3793), .ZN(n3797) );
  INV_X1 U4770 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5891) );
  OAI21_X1 U4771 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5891), .A(n4191), .ZN(
        n3795) );
  AOI21_X1 U4772 ( .B1(n3567), .B2(EAX_REG_21__SCAN_IN), .A(n3795), .ZN(n3796)
         );
  OAI21_X1 U4773 ( .B1(n4188), .B2(n3797), .A(n3796), .ZN(n3799) );
  XNOR2_X1 U4774 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n3814), .ZN(n5893)
         );
  NAND2_X1 U4775 ( .A1(n4185), .A2(n5893), .ZN(n3798) );
  NAND2_X1 U4776 ( .A1(n3799), .A2(n3798), .ZN(n5668) );
  AOI22_X1 U4777 ( .A1(n4165), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4778 ( .A1(n4172), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4779 ( .A1(n4174), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4780 ( .A1(n3407), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3800) );
  NAND4_X1 U4781 ( .A1(n3803), .A2(n3802), .A3(n3801), .A4(n3800), .ZN(n3809)
         );
  AOI22_X1 U4782 ( .A1(n4166), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4161), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4783 ( .A1(n4163), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4784 ( .A1(n3139), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4785 ( .A1(n4141), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3804) );
  NAND4_X1 U4786 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(n3808)
         );
  NOR2_X1 U4787 ( .A1(n3809), .A2(n3808), .ZN(n3813) );
  NAND2_X1 U4788 ( .A1(n6935), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3810)
         );
  NAND2_X1 U4789 ( .A1(n4191), .A2(n3810), .ZN(n3811) );
  AOI21_X1 U4790 ( .B1(n3567), .B2(EAX_REG_22__SCAN_IN), .A(n3811), .ZN(n3812)
         );
  OAI21_X1 U4791 ( .B1(n4188), .B2(n3813), .A(n3812), .ZN(n3818) );
  OAI21_X1 U4792 ( .B1(n3816), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n3860), 
        .ZN(n5885) );
  OR2_X1 U4793 ( .A1(n5885), .A2(n4191), .ZN(n3817) );
  NAND2_X1 U4794 ( .A1(n3818), .A2(n3817), .ZN(n5669) );
  AOI22_X1 U4795 ( .A1(n3137), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4166), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4796 ( .A1(n4084), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4797 ( .A1(n3138), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4798 ( .A1(n4172), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3820) );
  NAND4_X1 U4799 ( .A1(n3823), .A2(n3822), .A3(n3821), .A4(n3820), .ZN(n3829)
         );
  AOI22_X1 U4800 ( .A1(n4165), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4801 ( .A1(n4163), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4802 ( .A1(n4161), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4803 ( .A1(n4174), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3824) );
  NAND4_X1 U4804 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), .ZN(n3828)
         );
  NOR2_X1 U4805 ( .A1(n3829), .A2(n3828), .ZN(n3847) );
  AOI22_X1 U4806 ( .A1(n4146), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4807 ( .A1(n4165), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4808 ( .A1(n4084), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4809 ( .A1(n4121), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3831) );
  NAND4_X1 U4810 ( .A1(n3834), .A2(n3833), .A3(n3832), .A4(n3831), .ZN(n3840)
         );
  AOI22_X1 U4811 ( .A1(n3137), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4163), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4812 ( .A1(n4174), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4813 ( .A1(n4166), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4814 ( .A1(n4171), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3835) );
  NAND4_X1 U4815 ( .A1(n3838), .A2(n3837), .A3(n3836), .A4(n3835), .ZN(n3839)
         );
  NOR2_X1 U4816 ( .A1(n3840), .A2(n3839), .ZN(n3848) );
  XOR2_X1 U4817 ( .A(n3847), .B(n3848), .Z(n3841) );
  NAND2_X1 U4818 ( .A1(n3841), .A2(n4156), .ZN(n3846) );
  NAND2_X1 U4819 ( .A1(n6935), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3842)
         );
  NAND2_X1 U4820 ( .A1(n4191), .A2(n3842), .ZN(n3843) );
  AOI21_X1 U4821 ( .B1(n3567), .B2(EAX_REG_23__SCAN_IN), .A(n3843), .ZN(n3845)
         );
  XNOR2_X1 U4822 ( .A(n3860), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5658)
         );
  NAND2_X1 U4823 ( .A1(n4411), .A2(n5655), .ZN(n5639) );
  INV_X1 U4824 ( .A(n5639), .ZN(n3868) );
  OR2_X1 U4825 ( .A1(n3848), .A2(n3847), .ZN(n3880) );
  AOI22_X1 U4826 ( .A1(n3137), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4166), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4827 ( .A1(n4141), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4828 ( .A1(n4165), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4163), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4829 ( .A1(n4121), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3849) );
  NAND4_X1 U4830 ( .A1(n3852), .A2(n3851), .A3(n3850), .A4(n3849), .ZN(n3858)
         );
  AOI22_X1 U4831 ( .A1(n4171), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3856) );
  INV_X1 U4832 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n7009) );
  AOI22_X1 U4833 ( .A1(n3407), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4834 ( .A1(n4174), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4835 ( .A1(n4172), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3853) );
  NAND4_X1 U4836 ( .A1(n3856), .A2(n3855), .A3(n3854), .A4(n3853), .ZN(n3857)
         );
  NOR2_X1 U4837 ( .A1(n3858), .A2(n3857), .ZN(n3879) );
  INV_X1 U4838 ( .A(n3879), .ZN(n3859) );
  XNOR2_X1 U4839 ( .A(n3880), .B(n3859), .ZN(n3866) );
  INV_X1 U4840 ( .A(EAX_REG_24__SCAN_IN), .ZN(n3864) );
  INV_X1 U4841 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5659) );
  XNOR2_X1 U4842 ( .A(n3886), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5869)
         );
  INV_X1 U4843 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5645) );
  NOR2_X1 U4844 ( .A1(n3861), .A2(n5645), .ZN(n3862) );
  AOI21_X1 U4845 ( .B1(n5869), .B2(n4185), .A(n3862), .ZN(n3863) );
  OAI21_X1 U4846 ( .B1(n4154), .B2(n3864), .A(n3863), .ZN(n3865) );
  AOI21_X1 U4847 ( .B1(n3866), .B2(n4156), .A(n3865), .ZN(n5640) );
  INV_X1 U4848 ( .A(n5640), .ZN(n3867) );
  AOI22_X1 U4849 ( .A1(n4165), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4850 ( .A1(n4146), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4851 ( .A1(n4166), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4852 ( .A1(n4141), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3869) );
  NAND4_X1 U4853 ( .A1(n3872), .A2(n3871), .A3(n3870), .A4(n3869), .ZN(n3878)
         );
  AOI22_X1 U4854 ( .A1(n4120), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4855 ( .A1(n4173), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4856 ( .A1(n4163), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4857 ( .A1(n4171), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3873) );
  NAND4_X1 U4858 ( .A1(n3876), .A2(n3875), .A3(n3874), .A4(n3873), .ZN(n3877)
         );
  NOR2_X1 U4859 ( .A1(n3878), .A2(n3877), .ZN(n4073) );
  OR2_X1 U4860 ( .A1(n3880), .A2(n3879), .ZN(n4072) );
  XOR2_X1 U4861 ( .A(n4073), .B(n4072), .Z(n3884) );
  INV_X1 U4862 ( .A(EAX_REG_25__SCAN_IN), .ZN(n3882) );
  NAND2_X1 U4863 ( .A1(n6935), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3881)
         );
  OAI211_X1 U4864 ( .C1(n4154), .C2(n3882), .A(n4191), .B(n3881), .ZN(n3883)
         );
  AOI21_X1 U4865 ( .B1(n3884), .B2(n4156), .A(n3883), .ZN(n3885) );
  INV_X1 U4866 ( .A(n3885), .ZN(n3888) );
  NAND2_X1 U4867 ( .A1(n3886), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3955)
         );
  XNOR2_X1 U4868 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .B(n3955), .ZN(n5507)
         );
  NAND2_X1 U4869 ( .A1(n5507), .A2(n4185), .ZN(n3887) );
  NAND2_X1 U4870 ( .A1(n3888), .A2(n3887), .ZN(n3891) );
  OR2_X1 U4871 ( .A1(n3891), .A2(n5640), .ZN(n4112) );
  INV_X1 U4872 ( .A(n4112), .ZN(n3889) );
  AND2_X1 U4873 ( .A1(n5655), .A2(n3889), .ZN(n3890) );
  INV_X1 U4874 ( .A(n5498), .ZN(n4052) );
  XNOR2_X1 U4875 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3896) );
  NAND2_X1 U4876 ( .A1(n3920), .A2(n3896), .ZN(n3894) );
  NAND2_X1 U4877 ( .A1(n6579), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3893) );
  NAND2_X1 U4878 ( .A1(n3894), .A2(n3893), .ZN(n3898) );
  XNOR2_X1 U4879 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3897) );
  INV_X1 U4880 ( .A(n3897), .ZN(n3895) );
  XNOR2_X1 U4881 ( .A(n3898), .B(n3895), .ZN(n3917) );
  XOR2_X1 U4882 ( .A(n3920), .B(n3896), .Z(n3924) );
  NAND2_X1 U4883 ( .A1(n3917), .A2(n3924), .ZN(n3913) );
  NAND2_X1 U4884 ( .A1(n3898), .A2(n3897), .ZN(n3900) );
  NAND2_X1 U4885 ( .A1(n6586), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3899) );
  NAND2_X1 U4886 ( .A1(n3900), .A2(n3899), .ZN(n3905) );
  XNOR2_X1 U4887 ( .A(n6988), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3903)
         );
  NAND2_X1 U4888 ( .A1(n3905), .A2(n3903), .ZN(n3902) );
  NAND2_X1 U4889 ( .A1(n7014), .A2(n6988), .ZN(n3901) );
  NAND2_X1 U4890 ( .A1(n3902), .A2(n3901), .ZN(n3909) );
  INV_X1 U4891 ( .A(n3903), .ZN(n3904) );
  XNOR2_X1 U4892 ( .A(n3905), .B(n3904), .ZN(n3906) );
  NAND2_X1 U4893 ( .A1(n3907), .A2(n3906), .ZN(n3940) );
  NAND2_X1 U4894 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6113), .ZN(n3910) );
  INV_X1 U4895 ( .A(n3947), .ZN(n3912) );
  OAI21_X1 U4896 ( .B1(n3913), .B2(n3940), .A(n3912), .ZN(n4460) );
  INV_X1 U4897 ( .A(n4460), .ZN(n3914) );
  NAND2_X1 U4898 ( .A1(n4461), .A2(n3914), .ZN(n4455) );
  INV_X1 U4899 ( .A(n3917), .ZN(n3915) );
  NAND2_X1 U4900 ( .A1(n3916), .A2(n3915), .ZN(n3918) );
  NAND2_X1 U4901 ( .A1(n3917), .A2(n3135), .ZN(n3936) );
  AND3_X1 U4902 ( .A1(n3937), .A2(n3918), .A3(n3936), .ZN(n3939) );
  INV_X1 U4903 ( .A(n3924), .ZN(n3919) );
  NOR2_X1 U4904 ( .A1(n3919), .A2(n6609), .ZN(n3926) );
  OAI21_X1 U4905 ( .B1(n3132), .B2(n4683), .A(n5493), .ZN(n3925) );
  AOI21_X1 U4906 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n3921), .A(n3920), 
        .ZN(n3929) );
  AOI21_X1 U4907 ( .B1(n3929), .B2(n3294), .A(n4689), .ZN(n3923) );
  INV_X1 U4908 ( .A(n3937), .ZN(n3922) );
  OAI22_X1 U4909 ( .A1(n3926), .A2(n3925), .B1(n3923), .B2(n3922), .ZN(n3927)
         );
  NAND2_X1 U4910 ( .A1(n3924), .A2(n3927), .ZN(n3934) );
  INV_X1 U4911 ( .A(n3925), .ZN(n3932) );
  INV_X1 U4912 ( .A(n3926), .ZN(n3931) );
  INV_X1 U4913 ( .A(n3927), .ZN(n3928) );
  NAND3_X1 U4914 ( .A1(n3929), .A2(n3928), .A3(n3135), .ZN(n3930) );
  OAI21_X1 U4915 ( .B1(n3932), .B2(n3931), .A(n3930), .ZN(n3933) );
  AOI21_X1 U4916 ( .B1(n4314), .B2(n3940), .A(n3941), .ZN(n3945) );
  INV_X1 U4917 ( .A(n3940), .ZN(n3942) );
  AOI22_X1 U4918 ( .A1(n3942), .A2(n3941), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6609), .ZN(n3943) );
  OAI21_X1 U4919 ( .B1(n3945), .B2(n3944), .A(n3943), .ZN(n3946) );
  AOI21_X1 U4920 ( .B1(n3135), .B2(n3947), .A(n3946), .ZN(n3948) );
  INV_X1 U4921 ( .A(n3948), .ZN(n3949) );
  NOR2_X1 U4922 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6619) );
  INV_X1 U4923 ( .A(n6619), .ZN(n3951) );
  NOR3_X1 U4924 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n3951), .A3(n6709), .ZN(
        n6615) );
  NAND2_X1 U4925 ( .A1(n6935), .A2(n6709), .ZN(n6616) );
  NOR3_X1 U4926 ( .A1(n6609), .A2(n6702), .A3(n6616), .ZN(n6604) );
  OR2_X2 U4927 ( .A1(n6715), .A2(n3951), .ZN(n6434) );
  OR2_X1 U4928 ( .A1(n6604), .A2(n3952), .ZN(n3953) );
  NOR2_X1 U4929 ( .A1(n6615), .A2(n3953), .ZN(n3954) );
  INV_X1 U4930 ( .A(n3955), .ZN(n3956) );
  INV_X1 U4931 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5852) );
  INV_X1 U4932 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5583) );
  INV_X1 U4933 ( .A(n4160), .ZN(n3957) );
  NAND2_X1 U4934 ( .A1(n3957), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n3958)
         );
  INV_X1 U4935 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4427) );
  NOR2_X1 U4936 ( .A1(n4204), .A2(n6709), .ZN(n3959) );
  NOR2_X1 U4937 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4059) );
  AND2_X4 U4938 ( .A1(n3150), .A2(n3960), .ZN(n4931) );
  INV_X1 U4939 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5514) );
  NOR2_X1 U4940 ( .A1(n4352), .A2(n5514), .ZN(n3961) );
  INV_X1 U4941 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3965) );
  NAND2_X1 U4942 ( .A1(n4931), .A2(n3965), .ZN(n3964) );
  NAND2_X1 U4943 ( .A1(n3136), .A2(n3153), .ZN(n3971) );
  INV_X1 U4944 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6900) );
  NAND2_X1 U4945 ( .A1(n3971), .A2(n6900), .ZN(n3963) );
  NAND3_X1 U4946 ( .A1(n3964), .A2(n3963), .A3(n3983), .ZN(n3967) );
  NAND2_X1 U4947 ( .A1(n3979), .A2(n3965), .ZN(n3966) );
  NAND2_X1 U4948 ( .A1(n3967), .A2(n3966), .ZN(n3970) );
  NAND2_X1 U4949 ( .A1(n3971), .A2(EBX_REG_0__SCAN_IN), .ZN(n3969) );
  INV_X1 U4950 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U4951 ( .A1(n3983), .A2(n5293), .ZN(n3968) );
  NAND2_X1 U4952 ( .A1(n3969), .A2(n3968), .ZN(n4797) );
  XNOR2_X1 U4953 ( .A(n3970), .B(n4797), .ZN(n4932) );
  NAND2_X1 U4954 ( .A1(n4932), .A2(n4931), .ZN(n4934) );
  NAND2_X1 U4955 ( .A1(n4934), .A2(n3970), .ZN(n4945) );
  INV_X1 U4956 ( .A(n3971), .ZN(n3972) );
  INV_X1 U4957 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3973) );
  NAND2_X1 U4958 ( .A1(n3152), .A2(n3973), .ZN(n3975) );
  INV_X1 U4959 ( .A(n3979), .ZN(n3980) );
  INV_X1 U4960 ( .A(EBX_REG_2__SCAN_IN), .ZN(n3976) );
  NAND2_X1 U4961 ( .A1(n4931), .A2(n3976), .ZN(n3974) );
  NAND3_X1 U4962 ( .A1(n3975), .A2(n3980), .A3(n3974), .ZN(n3978) );
  NAND2_X1 U4963 ( .A1(n3979), .A2(n3976), .ZN(n3977) );
  AND2_X1 U4964 ( .A1(n3978), .A2(n3977), .ZN(n4944) );
  NAND2_X1 U4965 ( .A1(n3980), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3981)
         );
  OAI211_X1 U4966 ( .C1(n4352), .C2(EBX_REG_3__SCAN_IN), .A(n4010), .B(n3981), 
        .ZN(n3982) );
  OAI21_X1 U4967 ( .B1(n4337), .B2(EBX_REG_3__SCAN_IN), .A(n3982), .ZN(n4940)
         );
  INV_X1 U4968 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6749) );
  NAND2_X1 U4969 ( .A1(n4010), .A2(n6749), .ZN(n3985) );
  INV_X1 U4970 ( .A(EBX_REG_4__SCAN_IN), .ZN(n3986) );
  NAND2_X1 U4971 ( .A1(n4931), .A2(n3986), .ZN(n3984) );
  NAND3_X1 U4972 ( .A1(n3985), .A2(n3980), .A3(n3984), .ZN(n3988) );
  NAND2_X1 U4973 ( .A1(n3979), .A2(n3986), .ZN(n3987) );
  NAND2_X1 U4974 ( .A1(n3988), .A2(n3987), .ZN(n4937) );
  MUX2_X1 U4975 ( .A(n4337), .B(n4004), .S(EBX_REG_5__SCAN_IN), .Z(n3989) );
  OAI21_X1 U4976 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4796), .A(n3989), 
        .ZN(n4707) );
  NAND2_X1 U4977 ( .A1(n3991), .A2(n3990), .ZN(n4708) );
  INV_X1 U4978 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4759) );
  NAND2_X1 U4979 ( .A1(n4010), .A2(n4759), .ZN(n3993) );
  INV_X1 U4980 ( .A(EBX_REG_6__SCAN_IN), .ZN(n3994) );
  NAND2_X1 U4981 ( .A1(n4931), .A2(n3994), .ZN(n3992) );
  NAND3_X1 U4982 ( .A1(n3993), .A2(n4004), .A3(n3992), .ZN(n3996) );
  NAND2_X1 U4983 ( .A1(n5780), .A2(n3994), .ZN(n3995) );
  OR2_X2 U4984 ( .A1(n4708), .A2(n4755), .ZN(n5051) );
  MUX2_X1 U4985 ( .A(n4337), .B(n4004), .S(EBX_REG_7__SCAN_IN), .Z(n3997) );
  OAI21_X1 U4986 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n4796), .A(n3997), 
        .ZN(n5050) );
  INV_X1 U4987 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U4988 ( .A1(n4010), .A2(n5227), .ZN(n3999) );
  INV_X1 U4989 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6913) );
  NAND2_X1 U4990 ( .A1(n4931), .A2(n6913), .ZN(n3998) );
  NAND3_X1 U4991 ( .A1(n3999), .A2(n4004), .A3(n3998), .ZN(n4001) );
  NAND2_X1 U4992 ( .A1(n5780), .A2(n6913), .ZN(n4000) );
  NAND2_X1 U4993 ( .A1(n4001), .A2(n4000), .ZN(n5221) );
  AND2_X2 U4994 ( .A1(n5222), .A2(n5221), .ZN(n5224) );
  MUX2_X1 U4995 ( .A(n4337), .B(n4004), .S(EBX_REG_9__SCAN_IN), .Z(n4003) );
  OR2_X1 U4996 ( .A1(n4796), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4002)
         );
  MUX2_X1 U4997 ( .A(n4004), .B(n4010), .S(EBX_REG_10__SCAN_IN), .Z(n4006) );
  NAND2_X1 U4998 ( .A1(n4352), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4005) );
  INV_X1 U4999 ( .A(n4007), .ZN(n5346) );
  NAND2_X1 U5000 ( .A1(n4004), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4008) );
  OAI211_X1 U5001 ( .C1(n4352), .C2(EBX_REG_11__SCAN_IN), .A(n4010), .B(n4008), 
        .ZN(n4009) );
  OAI21_X1 U5002 ( .B1(n4337), .B2(EBX_REG_11__SCAN_IN), .A(n4009), .ZN(n5307)
         );
  MUX2_X1 U5003 ( .A(n3980), .B(n4010), .S(EBX_REG_12__SCAN_IN), .Z(n4012) );
  NAND2_X1 U5004 ( .A1(n4352), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4011) );
  NAND2_X1 U5005 ( .A1(n4012), .A2(n4011), .ZN(n5356) );
  AND2_X2 U5006 ( .A1(n5357), .A2(n5356), .ZN(n5438) );
  INV_X1 U5007 ( .A(n4337), .ZN(n4046) );
  INV_X1 U5008 ( .A(EBX_REG_13__SCAN_IN), .ZN(n4013) );
  NAND2_X1 U5009 ( .A1(n4046), .A2(n4013), .ZN(n4016) );
  NAND2_X1 U5010 ( .A1(n4004), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4014) );
  OAI211_X1 U5011 ( .C1(n4352), .C2(EBX_REG_13__SCAN_IN), .A(n4010), .B(n4014), 
        .ZN(n4015) );
  MUX2_X1 U5012 ( .A(n4004), .B(n4010), .S(EBX_REG_14__SCAN_IN), .Z(n4018) );
  NAND2_X1 U5013 ( .A1(n4352), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4017) );
  OR2_X2 U5014 ( .A1(n5454), .A2(n5453), .ZN(n5731) );
  NAND2_X1 U5015 ( .A1(n3980), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4019) );
  OAI211_X1 U5016 ( .C1(n4352), .C2(EBX_REG_15__SCAN_IN), .A(n4010), .B(n4019), 
        .ZN(n4020) );
  OAI21_X1 U5017 ( .B1(n4337), .B2(EBX_REG_15__SCAN_IN), .A(n4020), .ZN(n5730)
         );
  NOR2_X4 U5018 ( .A1(n5731), .A2(n5730), .ZN(n5733) );
  MUX2_X1 U5019 ( .A(n4004), .B(n4010), .S(EBX_REG_16__SCAN_IN), .Z(n4022) );
  NAND2_X1 U5020 ( .A1(n4352), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4021) );
  NAND2_X1 U5021 ( .A1(n4022), .A2(n4021), .ZN(n5714) );
  AND2_X2 U5022 ( .A1(n5733), .A2(n5714), .ZN(n5716) );
  INV_X1 U5023 ( .A(EBX_REG_17__SCAN_IN), .ZN(n4023) );
  NAND2_X1 U5024 ( .A1(n4046), .A2(n4023), .ZN(n4026) );
  NAND2_X1 U5025 ( .A1(n4004), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4024) );
  OAI211_X1 U5026 ( .C1(n4352), .C2(EBX_REG_17__SCAN_IN), .A(n4010), .B(n4024), 
        .ZN(n4025) );
  INV_X1 U5027 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6897) );
  NAND2_X1 U5028 ( .A1(n4010), .A2(n6897), .ZN(n4028) );
  INV_X1 U5029 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6957) );
  NAND2_X1 U5030 ( .A1(n4931), .A2(n6957), .ZN(n4027) );
  NAND3_X1 U5031 ( .A1(n4028), .A2(n3980), .A3(n4027), .ZN(n4030) );
  NAND2_X1 U5032 ( .A1(n5780), .A2(n6957), .ZN(n4029) );
  AND2_X1 U5033 ( .A1(n4030), .A2(n4029), .ZN(n5790) );
  OR2_X2 U5034 ( .A1(n5802), .A2(n5790), .ZN(n5789) );
  NAND2_X1 U5035 ( .A1(n4796), .A2(EBX_REG_18__SCAN_IN), .ZN(n4032) );
  NAND2_X1 U5036 ( .A1(n4352), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4031) );
  NAND2_X1 U5037 ( .A1(n4032), .A2(n4031), .ZN(n5781) );
  OR2_X1 U5038 ( .A1(n5781), .A2(n4004), .ZN(n5788) );
  OR2_X1 U5039 ( .A1(n4796), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4034)
         );
  INV_X1 U5040 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5784) );
  NAND2_X1 U5041 ( .A1(n4931), .A2(n5784), .ZN(n4033) );
  NAND2_X1 U5042 ( .A1(n4034), .A2(n4033), .ZN(n4035) );
  NAND2_X1 U5043 ( .A1(n5788), .A2(n4035), .ZN(n4037) );
  NAND2_X1 U5044 ( .A1(n5781), .A2(n4004), .ZN(n5787) );
  INV_X1 U5045 ( .A(n4035), .ZN(n5782) );
  NAND2_X1 U5046 ( .A1(n5787), .A2(n5782), .ZN(n4036) );
  NAND2_X1 U5047 ( .A1(n4037), .A2(n4036), .ZN(n4038) );
  MUX2_X1 U5048 ( .A(n4337), .B(n4004), .S(EBX_REG_21__SCAN_IN), .Z(n4039) );
  OAI21_X1 U5049 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n4796), .A(n4039), 
        .ZN(n5685) );
  MUX2_X1 U5050 ( .A(n3980), .B(n4010), .S(EBX_REG_22__SCAN_IN), .Z(n4041) );
  NAND2_X1 U5051 ( .A1(n4352), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4040) );
  NAND2_X1 U5052 ( .A1(n4041), .A2(n4040), .ZN(n5672) );
  NAND2_X1 U5053 ( .A1(n5687), .A2(n5672), .ZN(n5651) );
  NAND2_X1 U5054 ( .A1(n4004), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4042) );
  OAI211_X1 U5055 ( .C1(n4352), .C2(EBX_REG_23__SCAN_IN), .A(n4010), .B(n4042), 
        .ZN(n4043) );
  OAI21_X1 U5056 ( .B1(n4337), .B2(EBX_REG_23__SCAN_IN), .A(n4043), .ZN(n5652)
         );
  MUX2_X1 U5057 ( .A(n4004), .B(n4010), .S(EBX_REG_24__SCAN_IN), .Z(n4045) );
  NAND2_X1 U5058 ( .A1(n4352), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4044) );
  INV_X1 U5059 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U5060 ( .A1(n4046), .A2(n5501), .ZN(n4049) );
  NAND2_X1 U5061 ( .A1(n4004), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4047) );
  OAI211_X1 U5062 ( .C1(n4352), .C2(EBX_REG_25__SCAN_IN), .A(n4010), .B(n4047), 
        .ZN(n4048) );
  AND2_X1 U5063 ( .A1(n4049), .A2(n4048), .ZN(n4050) );
  AND2_X2 U5064 ( .A1(n5643), .A2(n4050), .ZN(n4336) );
  NOR2_X1 U5065 ( .A1(n5643), .A2(n4050), .ZN(n4051) );
  OR2_X1 U5066 ( .A1(n4336), .A2(n4051), .ZN(n6068) );
  OAI22_X1 U5067 ( .A1(n4052), .A2(n6171), .B1(n6257), .B2(n6068), .ZN(n4071)
         );
  NAND2_X1 U5068 ( .A1(n6196), .A2(n5507), .ZN(n4063) );
  NAND3_X1 U5069 ( .A1(n4054), .A2(n3962), .A3(n5514), .ZN(n4058) );
  INV_X1 U5070 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6628) );
  NAND2_X1 U5071 ( .A1(n4055), .A2(n6628), .ZN(n6596) );
  INV_X1 U5072 ( .A(n4059), .ZN(n4057) );
  OAI211_X1 U5073 ( .C1(n6596), .C2(n4057), .A(n6732), .B(n4456), .ZN(n4428)
         );
  AOI22_X1 U5074 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6264), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6239), .ZN(n4062) );
  NAND2_X1 U5075 ( .A1(n4683), .A2(n6596), .ZN(n4322) );
  AND3_X1 U5076 ( .A1(n4322), .A2(n4059), .A3(n3962), .ZN(n4060) );
  INV_X1 U5077 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6670) );
  INV_X1 U5078 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6664) );
  INV_X1 U5079 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6662) );
  INV_X1 U5080 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6653) );
  INV_X1 U5081 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6641) );
  NAND3_X1 U5082 ( .A1(REIP_REG_3__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        REIP_REG_1__SCAN_IN), .ZN(n6244) );
  NOR2_X1 U5083 ( .A1(n6641), .A2(n6244), .ZN(n6222) );
  NAND2_X1 U5084 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6222), .ZN(n5187) );
  INV_X1 U5085 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6649) );
  INV_X1 U5086 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6647) );
  INV_X1 U5087 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6645) );
  NOR3_X1 U5088 ( .A1(n6649), .A2(n6647), .A3(n6645), .ZN(n5191) );
  NAND2_X1 U5089 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5191), .ZN(n6184) );
  NOR3_X1 U5090 ( .A1(n6653), .A2(n5187), .A3(n6184), .ZN(n5745) );
  NAND2_X1 U5091 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5745), .ZN(n5718) );
  NAND3_X1 U5092 ( .A1(REIP_REG_12__SCAN_IN), .A2(REIP_REG_14__SCAN_IN), .A3(
        REIP_REG_13__SCAN_IN), .ZN(n5719) );
  NOR2_X1 U5093 ( .A1(n5718), .A2(n5719), .ZN(n5717) );
  NAND2_X1 U5094 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5717), .ZN(n5703) );
  NOR3_X1 U5095 ( .A1(n6664), .A2(n6662), .A3(n5703), .ZN(n5705) );
  NAND4_X1 U5096 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5705), .A3(
        REIP_REG_19__SCAN_IN), .A4(REIP_REG_18__SCAN_IN), .ZN(n5690) );
  NOR2_X1 U5097 ( .A1(n6670), .A2(n5690), .ZN(n4065) );
  NAND2_X1 U5098 ( .A1(n6246), .A2(n4065), .ZN(n5679) );
  INV_X1 U5099 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6674) );
  INV_X1 U5100 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6955) );
  NOR2_X1 U5101 ( .A1(n6674), .A2(n6955), .ZN(n4064) );
  INV_X1 U5102 ( .A(n4064), .ZN(n4061) );
  NAND2_X1 U5103 ( .A1(REIP_REG_24__SCAN_IN), .A2(n4416), .ZN(n5631) );
  NAND3_X1 U5104 ( .A1(n4063), .A2(n4062), .A3(n3159), .ZN(n4069) );
  NAND2_X1 U5105 ( .A1(n4065), .A2(n4064), .ZN(n4066) );
  NAND2_X1 U5106 ( .A1(n6246), .A2(n4066), .ZN(n4067) );
  AND2_X1 U5107 ( .A1(n4067), .A2(n5754), .ZN(n5657) );
  INV_X1 U5108 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6677) );
  NAND2_X1 U5109 ( .A1(n4416), .A2(n6677), .ZN(n5649) );
  INV_X1 U5110 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6846) );
  AOI21_X1 U5111 ( .B1(n5657), .B2(n5649), .A(n6846), .ZN(n4068) );
  OR2_X1 U5112 ( .A1(n4071), .A2(n4070), .ZN(U2802) );
  NOR2_X1 U5113 ( .A1(n4073), .A2(n4072), .ZN(n4103) );
  AOI22_X1 U5114 ( .A1(n4163), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U5115 ( .A1(n4174), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U5116 ( .A1(n4171), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4075) );
  AOI22_X1 U5117 ( .A1(n4121), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4074) );
  NAND4_X1 U5118 ( .A1(n4077), .A2(n4076), .A3(n4075), .A4(n4074), .ZN(n4083)
         );
  AOI22_X1 U5119 ( .A1(n4141), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4166), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4081) );
  AOI22_X1 U5120 ( .A1(n3137), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4080) );
  AOI22_X1 U5121 ( .A1(n4161), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4079) );
  AOI22_X1 U5122 ( .A1(n4165), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4078) );
  NAND4_X1 U5123 ( .A1(n4081), .A2(n4080), .A3(n4079), .A4(n4078), .ZN(n4082)
         );
  OR2_X1 U5124 ( .A1(n4083), .A2(n4082), .ZN(n4101) );
  NAND2_X1 U5125 ( .A1(n4103), .A2(n4101), .ZN(n4118) );
  AOI22_X1 U5126 ( .A1(n4165), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4088) );
  AOI22_X1 U5127 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n4084), .B1(n4174), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4087) );
  AOI22_X1 U5128 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4171), .B1(n4173), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4086) );
  AOI22_X1 U5129 ( .A1(n4166), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4085) );
  NAND4_X1 U5130 ( .A1(n4088), .A2(n4087), .A3(n4086), .A4(n4085), .ZN(n4095)
         );
  AOI22_X1 U5131 ( .A1(n4163), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4093) );
  AOI22_X1 U5132 ( .A1(n3137), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4092) );
  AOI22_X1 U5133 ( .A1(n4146), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U5134 ( .A1(n4162), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4090) );
  NAND4_X1 U5135 ( .A1(n4093), .A2(n4092), .A3(n4091), .A4(n4090), .ZN(n4094)
         );
  NOR2_X1 U5136 ( .A1(n4095), .A2(n4094), .ZN(n4119) );
  XOR2_X1 U5137 ( .A(n4118), .B(n4119), .Z(n4096) );
  NAND2_X1 U5138 ( .A1(n4096), .A2(n4156), .ZN(n4100) );
  OAI21_X1 U5139 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5852), .A(n4191), .ZN(
        n4097) );
  AOI21_X1 U5140 ( .B1(n3567), .B2(EAX_REG_27__SCAN_IN), .A(n4097), .ZN(n4099)
         );
  XNOR2_X1 U5141 ( .A(n4107), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5856)
         );
  AND2_X1 U5142 ( .A1(n5856), .A2(n4185), .ZN(n4098) );
  AOI21_X1 U5143 ( .B1(n4100), .B2(n4099), .A(n4098), .ZN(n4409) );
  INV_X1 U5144 ( .A(n4101), .ZN(n4102) );
  XNOR2_X1 U5145 ( .A(n4103), .B(n4102), .ZN(n4104) );
  NAND2_X1 U5146 ( .A1(n4104), .A2(n4156), .ZN(n4111) );
  INV_X1 U5147 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4105) );
  AOI21_X1 U5148 ( .B1(n4105), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4106) );
  AOI21_X1 U5149 ( .B1(n3567), .B2(EAX_REG_26__SCAN_IN), .A(n4106), .ZN(n4110)
         );
  OAI21_X1 U5150 ( .B1(n4108), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n4107), 
        .ZN(n5629) );
  NOR2_X1 U5151 ( .A1(n5629), .A2(n4191), .ZN(n4109) );
  AOI21_X1 U5152 ( .B1(n4111), .B2(n4110), .A(n4109), .ZN(n4437) );
  INV_X1 U5153 ( .A(n4437), .ZN(n4113) );
  NOR2_X1 U5154 ( .A1(n4113), .A2(n4112), .ZN(n4407) );
  AND2_X1 U5155 ( .A1(n4409), .A2(n4407), .ZN(n4114) );
  INV_X1 U5156 ( .A(n4115), .ZN(n4116) );
  INV_X1 U5157 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U5158 ( .A1(n4116), .A2(n5619), .ZN(n4117) );
  NAND2_X1 U5159 ( .A1(n4138), .A2(n4117), .ZN(n5845) );
  NOR2_X1 U5160 ( .A1(n4119), .A2(n4118), .ZN(n4140) );
  AOI22_X1 U5161 ( .A1(n4163), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5162 ( .A1(n4120), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5163 ( .A1(n4171), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4123) );
  AOI22_X1 U5164 ( .A1(n4121), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4122) );
  NAND4_X1 U5165 ( .A1(n4125), .A2(n4124), .A3(n4123), .A4(n4122), .ZN(n4131)
         );
  AOI22_X1 U5166 ( .A1(n4141), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4166), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U5167 ( .A1(n3137), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4128) );
  AOI22_X1 U5168 ( .A1(n4146), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4127) );
  AOI22_X1 U5169 ( .A1(n4165), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4126) );
  NAND4_X1 U5170 ( .A1(n4129), .A2(n4128), .A3(n4127), .A4(n4126), .ZN(n4130)
         );
  OR2_X1 U5171 ( .A1(n4131), .A2(n4130), .ZN(n4139) );
  XNOR2_X1 U5172 ( .A(n4140), .B(n4139), .ZN(n4134) );
  AOI21_X1 U5173 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6935), .A(n4185), 
        .ZN(n4133) );
  NAND2_X1 U5174 ( .A1(n4193), .A2(EAX_REG_28__SCAN_IN), .ZN(n4132) );
  OAI211_X1 U5175 ( .C1(n4134), .C2(n4188), .A(n4133), .B(n4132), .ZN(n4135)
         );
  OAI21_X1 U5176 ( .B1(n4191), .B2(n5845), .A(n4135), .ZN(n5614) );
  INV_X1 U5177 ( .A(n5614), .ZN(n4136) );
  XNOR2_X1 U5178 ( .A(n4138), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5606)
         );
  NAND2_X1 U5179 ( .A1(n4140), .A2(n4139), .ZN(n4181) );
  AOI22_X1 U5180 ( .A1(n4166), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4163), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4145) );
  AOI22_X1 U5181 ( .A1(n4173), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4144) );
  AOI22_X1 U5182 ( .A1(n4141), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4143) );
  AOI22_X1 U5183 ( .A1(n4172), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4142) );
  NAND4_X1 U5184 ( .A1(n4145), .A2(n4144), .A3(n4143), .A4(n4142), .ZN(n4152)
         );
  AOI22_X1 U5185 ( .A1(n4165), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U5186 ( .A1(n4146), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U5187 ( .A1(n4174), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U5188 ( .A1(n3138), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4147) );
  NAND4_X1 U5189 ( .A1(n4150), .A2(n4149), .A3(n4148), .A4(n4147), .ZN(n4151)
         );
  NOR2_X1 U5190 ( .A1(n4152), .A2(n4151), .ZN(n4182) );
  XOR2_X1 U5191 ( .A(n4181), .B(n4182), .Z(n4157) );
  INV_X1 U5192 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4508) );
  AOI21_X1 U5193 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6935), .A(n4185), 
        .ZN(n4153) );
  OAI21_X1 U5194 ( .B1(n4154), .B2(n4508), .A(n4153), .ZN(n4155) );
  AOI21_X1 U5195 ( .B1(n4157), .B2(n4156), .A(n4155), .ZN(n4158) );
  AOI21_X1 U5196 ( .B1(n4185), .B2(n5606), .A(n4158), .ZN(n5580) );
  INV_X1 U5197 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4159) );
  XNOR2_X1 U5198 ( .A(n4160), .B(n4159), .ZN(n5596) );
  AOI22_X1 U5199 ( .A1(n3137), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4161), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4170) );
  AOI22_X1 U5200 ( .A1(n4163), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4162), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U5201 ( .A1(n4165), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U5202 ( .A1(n4166), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4167) );
  NAND4_X1 U5203 ( .A1(n4170), .A2(n4169), .A3(n4168), .A4(n4167), .ZN(n4180)
         );
  AOI22_X1 U5204 ( .A1(n4141), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4178) );
  AOI22_X1 U5205 ( .A1(n4172), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4177) );
  AOI22_X1 U5206 ( .A1(n4174), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4176) );
  AOI22_X1 U5207 ( .A1(n3138), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4175) );
  NAND4_X1 U5208 ( .A1(n4178), .A2(n4177), .A3(n4176), .A4(n4175), .ZN(n4179)
         );
  NOR2_X1 U5209 ( .A1(n4180), .A2(n4179), .ZN(n4184) );
  NOR2_X1 U5210 ( .A1(n4182), .A2(n4181), .ZN(n4183) );
  XOR2_X1 U5211 ( .A(n4184), .B(n4183), .Z(n4189) );
  AOI21_X1 U5212 ( .B1(PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6935), .A(n4185), 
        .ZN(n4187) );
  NAND2_X1 U5213 ( .A1(n4193), .A2(EAX_REG_30__SCAN_IN), .ZN(n4186) );
  OAI211_X1 U5214 ( .C1(n4189), .C2(n4188), .A(n4187), .B(n4186), .ZN(n4190)
         );
  OAI21_X1 U5215 ( .B1(n4191), .B2(n5596), .A(n4190), .ZN(n5521) );
  AOI22_X1 U5216 ( .A1(n4193), .A2(EAX_REG_31__SCAN_IN), .B1(n4192), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4194) );
  NAND3_X1 U5217 ( .A1(n6609), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6617) );
  INV_X1 U5218 ( .A(n6617), .ZN(n4195) );
  NAND2_X2 U5219 ( .A1(n4195), .A2(n6442), .ZN(n6361) );
  AOI21_X1 U5220 ( .B1(n4689), .B2(n4196), .A(n4359), .ZN(n4197) );
  NAND2_X1 U5221 ( .A1(n4327), .A2(n4198), .ZN(n6569) );
  NAND2_X1 U5222 ( .A1(n6729), .A2(n6728), .ZN(n4199) );
  NAND2_X1 U5223 ( .A1(n4199), .A2(n6609), .ZN(n4200) );
  NAND2_X1 U5224 ( .A1(n6609), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4202) );
  NAND2_X1 U5225 ( .A1(n6121), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4201) );
  NAND2_X1 U5226 ( .A1(n4202), .A2(n4201), .ZN(n6357) );
  NAND2_X1 U5227 ( .A1(n3952), .A2(REIP_REG_31__SCAN_IN), .ZN(n4377) );
  NAND2_X1 U5228 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4203)
         );
  OAI211_X1 U5229 ( .C1(n6352), .C2(n4204), .A(n4377), .B(n4203), .ZN(n4205)
         );
  AOI21_X1 U5230 ( .B1(n5818), .B2(n6347), .A(n4205), .ZN(n4313) );
  NOR2_X1 U5231 ( .A1(n4207), .A2(n4270), .ZN(n4208) );
  INV_X1 U5232 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4286) );
  NOR2_X1 U5233 ( .A1(n5880), .A2(n4286), .ZN(n5463) );
  XNOR2_X1 U5234 ( .A(n5880), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5470)
         );
  INV_X1 U5235 ( .A(n5470), .ZN(n4287) );
  OR2_X1 U5236 ( .A1(n5463), .A2(n4287), .ZN(n5441) );
  INV_X1 U5237 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5443) );
  OR2_X1 U5238 ( .A1(n5441), .A2(n3164), .ZN(n4291) );
  INV_X1 U5239 ( .A(n4638), .ZN(n4209) );
  NAND2_X1 U5240 ( .A1(n4209), .A2(n4314), .ZN(n4212) );
  NAND2_X1 U5241 ( .A1(n4217), .A2(n4218), .ZN(n4227) );
  NAND2_X1 U5242 ( .A1(n4227), .A2(n4228), .ZN(n4226) );
  NAND2_X1 U5243 ( .A1(n4226), .A2(n4210), .ZN(n4249) );
  OAI211_X1 U5244 ( .C1(n4210), .C2(n4226), .A(n4249), .B(n4456), .ZN(n4211)
         );
  NAND2_X1 U5245 ( .A1(n4212), .A2(n4211), .ZN(n4236) );
  INV_X1 U5246 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n7003) );
  NAND2_X1 U5247 ( .A1(n4689), .A2(n4213), .ZN(n4229) );
  OAI21_X1 U5248 ( .B1(n6735), .B2(n4218), .A(n4229), .ZN(n4214) );
  INV_X1 U5249 ( .A(n4214), .ZN(n4215) );
  OAI21_X1 U5250 ( .B1(n5379), .B2(n4270), .A(n4215), .ZN(n6354) );
  NAND2_X1 U5251 ( .A1(n6354), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6353)
         );
  XNOR2_X1 U5252 ( .A(n6353), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4543)
         );
  OAI21_X1 U5253 ( .B1(n4218), .B2(n4217), .A(n4227), .ZN(n4220) );
  INV_X1 U5254 ( .A(n4359), .ZN(n4219) );
  OAI211_X1 U5255 ( .C1(n4220), .C2(n6735), .A(n4219), .B(n5493), .ZN(n4221)
         );
  INV_X1 U5256 ( .A(n4221), .ZN(n4222) );
  NAND2_X1 U5257 ( .A1(n4223), .A2(n4222), .ZN(n4542) );
  NAND2_X1 U5258 ( .A1(n4543), .A2(n4542), .ZN(n4544) );
  INV_X1 U5259 ( .A(n6353), .ZN(n4224) );
  NAND2_X1 U5260 ( .A1(n4224), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4225)
         );
  OR2_X1 U5261 ( .A1(n4639), .A2(n4270), .ZN(n4233) );
  OAI21_X1 U5262 ( .B1(n4228), .B2(n4227), .A(n4226), .ZN(n4231) );
  INV_X1 U5263 ( .A(n4229), .ZN(n4230) );
  AOI21_X1 U5264 ( .B1(n4231), .B2(n4456), .A(n4230), .ZN(n4232) );
  NAND2_X1 U5265 ( .A1(n4233), .A2(n4232), .ZN(n6343) );
  NAND2_X1 U5266 ( .A1(n6344), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4234)
         );
  NAND2_X1 U5267 ( .A1(n4235), .A2(n4234), .ZN(n4555) );
  NAND2_X1 U5268 ( .A1(n4556), .A2(n4555), .ZN(n4238) );
  NAND2_X1 U5269 ( .A1(n4236), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4237)
         );
  NAND2_X1 U5270 ( .A1(n4238), .A2(n4237), .ZN(n4723) );
  XNOR2_X1 U5271 ( .A(n4249), .B(n4247), .ZN(n4239) );
  NAND2_X1 U5272 ( .A1(n4239), .A2(n4456), .ZN(n4240) );
  OAI21_X1 U5273 ( .B1(n4241), .B2(n4270), .A(n4240), .ZN(n4242) );
  XNOR2_X1 U5274 ( .A(n4242), .B(n6749), .ZN(n4724) );
  NAND2_X1 U5275 ( .A1(n4723), .A2(n4724), .ZN(n4244) );
  NAND2_X1 U5276 ( .A1(n4242), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4243)
         );
  NAND2_X1 U5277 ( .A1(n4244), .A2(n4243), .ZN(n4827) );
  INV_X1 U5278 ( .A(n4245), .ZN(n4246) );
  NAND2_X1 U5279 ( .A1(n4246), .A2(n4314), .ZN(n4253) );
  INV_X1 U5280 ( .A(n4247), .ZN(n4248) );
  NOR2_X1 U5281 ( .A1(n4249), .A2(n4248), .ZN(n4251) );
  NAND2_X1 U5282 ( .A1(n4251), .A2(n4250), .ZN(n4265) );
  OAI211_X1 U5283 ( .C1(n4251), .C2(n4250), .A(n4265), .B(n4456), .ZN(n4252)
         );
  NAND2_X1 U5284 ( .A1(n4253), .A2(n4252), .ZN(n4254) );
  INV_X1 U5285 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4384) );
  XNOR2_X1 U5286 ( .A(n4254), .B(n4384), .ZN(n4828) );
  NAND2_X1 U5287 ( .A1(n4827), .A2(n4828), .ZN(n4256) );
  NAND2_X1 U5288 ( .A1(n4254), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4255)
         );
  NAND2_X1 U5289 ( .A1(n4256), .A2(n4255), .ZN(n4750) );
  NAND3_X1 U5290 ( .A1(n4206), .A2(n4314), .A3(n4257), .ZN(n4260) );
  XNOR2_X1 U5291 ( .A(n4265), .B(n4266), .ZN(n4258) );
  NAND2_X1 U5292 ( .A1(n4258), .A2(n4456), .ZN(n4259) );
  NAND2_X1 U5293 ( .A1(n4260), .A2(n4259), .ZN(n4261) );
  XNOR2_X1 U5294 ( .A(n4261), .B(n4759), .ZN(n4752) );
  NAND2_X1 U5295 ( .A1(n4750), .A2(n4752), .ZN(n4263) );
  NAND2_X1 U5296 ( .A1(n4261), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4262)
         );
  NAND2_X1 U5297 ( .A1(n4263), .A2(n4262), .ZN(n5200) );
  INV_X1 U5298 ( .A(n4264), .ZN(n4271) );
  INV_X1 U5299 ( .A(n4265), .ZN(n4267) );
  NAND2_X1 U5300 ( .A1(n4267), .A2(n4266), .ZN(n4277) );
  XNOR2_X1 U5301 ( .A(n4277), .B(n4275), .ZN(n4268) );
  NAND2_X1 U5302 ( .A1(n4268), .A2(n4456), .ZN(n4269) );
  INV_X1 U5303 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6387) );
  XNOR2_X1 U5304 ( .A(n4272), .B(n6387), .ZN(n5201) );
  NAND2_X1 U5305 ( .A1(n5200), .A2(n5201), .ZN(n4274) );
  NAND2_X1 U5306 ( .A1(n4272), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4273)
         );
  NAND2_X1 U5307 ( .A1(n4274), .A2(n4273), .ZN(n5218) );
  NAND2_X1 U5308 ( .A1(n4456), .A2(n4275), .ZN(n4276) );
  OR2_X1 U5309 ( .A1(n4277), .A2(n4276), .ZN(n4278) );
  NAND2_X1 U5310 ( .A1(n5880), .A2(n4278), .ZN(n4279) );
  XNOR2_X1 U5311 ( .A(n4279), .B(n5227), .ZN(n5219) );
  NAND2_X1 U5312 ( .A1(n5218), .A2(n5219), .ZN(n4281) );
  NAND2_X1 U5313 ( .A1(n4279), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4280)
         );
  INV_X1 U5314 ( .A(n5315), .ZN(n4283) );
  INV_X1 U5315 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6377) );
  NOR2_X1 U5316 ( .A1(n5880), .A2(n6377), .ZN(n5329) );
  INV_X1 U5317 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n7012) );
  OR2_X1 U5318 ( .A1(n5880), .A2(n7012), .ZN(n5333) );
  INV_X1 U5319 ( .A(n5333), .ZN(n4282) );
  INV_X1 U5320 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6365) );
  NAND2_X1 U5321 ( .A1(n5880), .A2(n6365), .ZN(n5370) );
  NAND2_X1 U5322 ( .A1(n5880), .A2(n6377), .ZN(n5331) );
  AND2_X1 U5323 ( .A1(n3165), .A2(n5331), .ZN(n5368) );
  AND2_X1 U5324 ( .A1(n5370), .A2(n5368), .ZN(n4284) );
  NAND2_X1 U5325 ( .A1(n5369), .A2(n4284), .ZN(n4285) );
  OR2_X1 U5326 ( .A1(n5880), .A2(n6365), .ZN(n5371) );
  INV_X1 U5327 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6758) );
  NAND2_X1 U5328 ( .A1(n5880), .A2(n6758), .ZN(n4288) );
  NAND2_X1 U5329 ( .A1(n5880), .A2(n4286), .ZN(n5465) );
  OR2_X1 U5330 ( .A1(n4287), .A2(n5465), .ZN(n5467) );
  OAI21_X1 U5331 ( .B1(n4291), .B2(n5352), .A(n4290), .ZN(n5918) );
  INV_X1 U5332 ( .A(n5880), .ZN(n5864) );
  XNOR2_X1 U5333 ( .A(n5989), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5917)
         );
  NAND2_X1 U5334 ( .A1(n5918), .A2(n5917), .ZN(n5903) );
  INV_X1 U5335 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n7010) );
  NAND2_X1 U5336 ( .A1(n5880), .A2(n7010), .ZN(n4292) );
  NAND2_X1 U5337 ( .A1(n5903), .A2(n4292), .ZN(n5902) );
  AND2_X1 U5338 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U5339 ( .A1(n6059), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4293) );
  AND2_X1 U5340 ( .A1(n5880), .A2(n4293), .ZN(n4296) );
  NOR3_X1 U5341 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(INSTADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n4294) );
  OR2_X1 U5342 ( .A1(n5880), .A2(n4294), .ZN(n4295) );
  NOR2_X1 U5343 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4298) );
  NOR2_X1 U5344 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4297) );
  INV_X1 U5345 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5987) );
  AND4_X1 U5346 ( .A1(n4298), .A2(n4297), .A3(n5987), .A4(n6897), .ZN(n4299)
         );
  NOR2_X1 U5347 ( .A1(n5989), .A2(n4299), .ZN(n4300) );
  AND2_X1 U5348 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4391) );
  AND2_X1 U5349 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4394) );
  NAND2_X1 U5350 ( .A1(n4391), .A2(n4394), .ZN(n5873) );
  NAND2_X1 U5351 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4397) );
  OAI21_X1 U5352 ( .B1(n5873), .B2(n4397), .A(n5989), .ZN(n4301) );
  NAND2_X1 U5353 ( .A1(n5838), .A2(n4301), .ZN(n5505) );
  XNOR2_X1 U5354 ( .A(n5880), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5506)
         );
  INV_X1 U5355 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6073) );
  AND2_X1 U5356 ( .A1(n5989), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4303)
         );
  NAND2_X1 U5357 ( .A1(n4442), .A2(n4303), .ZN(n5850) );
  NAND2_X1 U5358 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5930) );
  AND2_X1 U5359 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4401) );
  NAND2_X1 U5360 ( .A1(n5566), .A2(n4401), .ZN(n4308) );
  INV_X1 U5361 ( .A(n4304), .ZN(n5504) );
  INV_X1 U5362 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4339) );
  INV_X1 U5363 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4305) );
  NAND2_X1 U5364 ( .A1(n4339), .A2(n4305), .ZN(n5931) );
  NAND2_X1 U5365 ( .A1(n4308), .A2(n4307), .ZN(n4309) );
  XNOR2_X1 U5366 ( .A(n4309), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4406)
         );
  INV_X1 U5367 ( .A(n4406), .ZN(n4311) );
  NAND2_X1 U5368 ( .A1(n4311), .A2(n4310), .ZN(n4312) );
  NAND2_X1 U5369 ( .A1(n4313), .A2(n4312), .ZN(U2955) );
  INV_X1 U5370 ( .A(n4461), .ZN(n4317) );
  NAND2_X1 U5371 ( .A1(n4314), .A2(n4805), .ZN(n4372) );
  OAI211_X1 U5372 ( .C1(n4315), .C2(n3704), .A(n3962), .B(n4372), .ZN(n4366)
         );
  NAND2_X1 U5373 ( .A1(n4327), .A2(n4366), .ZN(n4316) );
  NAND2_X1 U5374 ( .A1(n4317), .A2(n4316), .ZN(n4610) );
  OR3_X1 U5375 ( .A1(n6601), .A2(n4196), .A3(n4683), .ZN(n4319) );
  INV_X1 U5376 ( .A(n6596), .ZN(n6627) );
  NOR2_X1 U5377 ( .A1(READY_N), .A2(n4460), .ZN(n4561) );
  OAI211_X1 U5378 ( .C1(n4683), .C2(n6627), .A(n4361), .B(n4561), .ZN(n4318)
         );
  NAND3_X1 U5379 ( .A1(n4610), .A2(n4319), .A3(n4318), .ZN(n4320) );
  NAND2_X1 U5380 ( .A1(n4320), .A2(n6606), .ZN(n4326) );
  INV_X1 U5381 ( .A(READY_N), .ZN(n6630) );
  NAND2_X1 U5382 ( .A1(n4322), .A2(n6630), .ZN(n4323) );
  OR2_X1 U5383 ( .A1(n4586), .A2(n4323), .ZN(n4603) );
  NAND3_X1 U5384 ( .A1(n4603), .A2(n3962), .A3(n4360), .ZN(n4324) );
  NAND3_X1 U5385 ( .A1(n4568), .A2(n4662), .A3(n4324), .ZN(n4325) );
  AND2_X1 U5386 ( .A1(n4327), .A2(n3146), .ZN(n4569) );
  INV_X1 U5387 ( .A(n4569), .ZN(n4601) );
  OAI22_X1 U5388 ( .A1(n4602), .A2(n4683), .B1(n4355), .B2(n3365), .ZN(n4328)
         );
  INV_X1 U5389 ( .A(n4328), .ZN(n4330) );
  NAND4_X1 U5390 ( .A1(n4601), .A2(n4330), .A3(n6108), .A4(n6569), .ZN(n4331)
         );
  INV_X1 U5391 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5841) );
  NAND2_X1 U5392 ( .A1(n4010), .A2(n5841), .ZN(n4333) );
  INV_X1 U5393 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5768) );
  NAND2_X1 U5394 ( .A1(n4931), .A2(n5768), .ZN(n4332) );
  NAND3_X1 U5395 ( .A1(n4333), .A2(n4004), .A3(n4332), .ZN(n4335) );
  NAND2_X1 U5396 ( .A1(n5780), .A2(n5768), .ZN(n4334) );
  NAND2_X1 U5397 ( .A1(n4335), .A2(n4334), .ZN(n5626) );
  NAND2_X1 U5398 ( .A1(n4336), .A2(n5626), .ZN(n4413) );
  MUX2_X1 U5399 ( .A(n4337), .B(n4004), .S(EBX_REG_27__SCAN_IN), .Z(n4338) );
  OAI21_X1 U5400 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n4796), .A(n4338), 
        .ZN(n4414) );
  OR2_X2 U5401 ( .A1(n4413), .A2(n4414), .ZN(n5616) );
  NAND2_X1 U5402 ( .A1(n4010), .A2(n4339), .ZN(n4341) );
  INV_X1 U5403 ( .A(EBX_REG_28__SCAN_IN), .ZN(n4342) );
  NAND2_X1 U5404 ( .A1(n4931), .A2(n4342), .ZN(n4340) );
  NAND3_X1 U5405 ( .A1(n4341), .A2(n4004), .A3(n4340), .ZN(n4344) );
  NAND2_X1 U5406 ( .A1(n5780), .A2(n4342), .ZN(n4343) );
  AND2_X1 U5407 ( .A1(n4344), .A2(n4343), .ZN(n5617) );
  NOR2_X2 U5408 ( .A1(n5616), .A2(n5617), .ZN(n4348) );
  OR2_X1 U5409 ( .A1(n4796), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4346)
         );
  INV_X1 U5410 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U5411 ( .A1(n4931), .A2(n5592), .ZN(n4345) );
  NAND2_X1 U5412 ( .A1(n4346), .A2(n4345), .ZN(n5570) );
  INV_X1 U5413 ( .A(n5570), .ZN(n4347) );
  AND2_X2 U5414 ( .A1(n4348), .A2(n4347), .ZN(n5527) );
  INV_X1 U5415 ( .A(n4348), .ZN(n5569) );
  NAND2_X1 U5416 ( .A1(n5780), .A2(n5592), .ZN(n5568) );
  AOI21_X1 U5417 ( .B1(n5527), .B2(n3980), .A(n4349), .ZN(n5572) );
  NAND2_X1 U5418 ( .A1(n4796), .A2(EBX_REG_30__SCAN_IN), .ZN(n4351) );
  NAND2_X1 U5419 ( .A1(n4352), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4350) );
  NAND2_X1 U5420 ( .A1(n4351), .A2(n4350), .ZN(n5528) );
  INV_X1 U5421 ( .A(n5527), .ZN(n5526) );
  NAND2_X2 U5422 ( .A1(n5526), .A2(n4004), .ZN(n5530) );
  OAI21_X2 U5423 ( .B1(n5572), .B2(n5528), .A(n5530), .ZN(n4354) );
  AOI22_X1 U5424 ( .A1(n4796), .A2(EBX_REG_31__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4352), .ZN(n4353) );
  OAI21_X1 U5425 ( .B1(n4355), .B2(n3249), .A(n6595), .ZN(n4356) );
  NOR2_X1 U5426 ( .A1(n5513), .A2(n6424), .ZN(n4404) );
  INV_X1 U5427 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4376) );
  INV_X1 U5428 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6100) );
  NAND3_X1 U5429 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5452) );
  NOR2_X1 U5430 ( .A1(n5443), .A2(n5452), .ZN(n6092) );
  NAND2_X1 U5431 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n6092), .ZN(n6093) );
  NOR2_X1 U5432 ( .A1(n6100), .A2(n6093), .ZN(n4390) );
  AND2_X1 U5433 ( .A1(n4461), .A2(n4357), .ZN(n6576) );
  INV_X1 U5434 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6416) );
  NOR2_X1 U5435 ( .A1(n4358), .A2(n4361), .ZN(n4607) );
  OAI21_X1 U5436 ( .B1(n4607), .B2(n4796), .A(n4359), .ZN(n4363) );
  NAND2_X1 U5437 ( .A1(n4361), .A2(n4360), .ZN(n4362) );
  OAI211_X1 U5438 ( .C1(n4364), .C2(n4004), .A(n4363), .B(n4362), .ZN(n4365)
         );
  INV_X1 U5439 ( .A(n4365), .ZN(n4367) );
  NAND3_X1 U5440 ( .A1(n4368), .A2(n4367), .A3(n4366), .ZN(n4588) );
  OAI21_X1 U5441 ( .B1(n4587), .B2(n3962), .A(n4617), .ZN(n4369) );
  INV_X1 U5442 ( .A(n4374), .ZN(n4370) );
  NAND2_X1 U5443 ( .A1(n4370), .A2(n4380), .ZN(n4386) );
  NAND2_X1 U5444 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U5445 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5341) );
  NOR2_X1 U5446 ( .A1(n5340), .A2(n5341), .ZN(n4389) );
  NAND2_X1 U5447 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4371) );
  NOR2_X1 U5448 ( .A1(n3973), .A2(n6900), .ZN(n4753) );
  NAND3_X1 U5449 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n4753), .ZN(n4830) );
  NOR2_X1 U5450 ( .A1(n4371), .A2(n4830), .ZN(n4385) );
  NAND2_X1 U5451 ( .A1(n4389), .A2(n4385), .ZN(n5474) );
  INV_X1 U5452 ( .A(n4380), .ZN(n4375) );
  INV_X1 U5453 ( .A(n4372), .ZN(n4373) );
  OAI21_X1 U5454 ( .B1(n6900), .B2(n6416), .A(n3973), .ZN(n6401) );
  NAND3_X1 U5455 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n6401), .ZN(n4383) );
  NOR2_X1 U5456 ( .A1(n5147), .A2(n4383), .ZN(n4832) );
  NAND4_X1 U5457 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n4832), .A4(n4389), .ZN(n5446) );
  NAND2_X1 U5458 ( .A1(n4390), .A2(n6366), .ZN(n5992) );
  NOR2_X1 U5459 ( .A1(n4376), .A2(n5992), .ZN(n6077) );
  NAND2_X1 U5460 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n6077), .ZN(n6001) );
  INV_X1 U5461 ( .A(n4391), .ZN(n5993) );
  NAND2_X1 U5462 ( .A1(n5984), .A2(n4394), .ZN(n5965) );
  NOR2_X1 U5463 ( .A1(n5965), .A2(n4397), .ZN(n6074) );
  AND2_X1 U5464 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5947) );
  NAND2_X1 U5465 ( .A1(n6074), .A2(n5947), .ZN(n5941) );
  NOR2_X1 U5466 ( .A1(n5941), .A2(n5930), .ZN(n5576) );
  NAND3_X1 U5467 ( .A1(n5576), .A2(n4401), .A3(n5544), .ZN(n4378) );
  NAND2_X1 U5468 ( .A1(n4378), .A2(n4377), .ZN(n4402) );
  NAND2_X1 U5469 ( .A1(n5147), .A2(n4386), .ZN(n6429) );
  INV_X1 U5470 ( .A(n6429), .ZN(n4379) );
  OR2_X1 U5471 ( .A1(n4386), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4382)
         );
  OR2_X1 U5472 ( .A1(n4380), .A2(n3952), .ZN(n4381) );
  INV_X1 U5473 ( .A(n5147), .ZN(n6413) );
  NOR2_X1 U5474 ( .A1(n4384), .A2(n4383), .ZN(n4760) );
  NAND2_X1 U5475 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4760), .ZN(n5226)
         );
  INV_X1 U5476 ( .A(n4385), .ZN(n4387) );
  NAND2_X1 U5477 ( .A1(n6415), .A2(n4386), .ZN(n4754) );
  AOI22_X1 U5478 ( .A1(n6413), .A2(n5226), .B1(n4387), .B2(n4754), .ZN(n4388)
         );
  NAND2_X1 U5479 ( .A1(n5355), .A2(n4388), .ZN(n5230) );
  OAI21_X1 U5480 ( .B1(n4389), .B2(n6414), .A(n6388), .ZN(n6367) );
  INV_X1 U5481 ( .A(n6367), .ZN(n5450) );
  OAI21_X1 U5482 ( .B1(n4390), .B2(n6414), .A(n5450), .ZN(n6087) );
  NAND3_X1 U5483 ( .A1(n4391), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4392) );
  AND2_X1 U5484 ( .A1(n6090), .A2(n4392), .ZN(n4393) );
  INV_X1 U5485 ( .A(n4394), .ZN(n4395) );
  AND2_X1 U5486 ( .A1(n6090), .A2(n4395), .ZN(n4396) );
  NOR2_X1 U5487 ( .A1(n5979), .A2(n4396), .ZN(n5962) );
  NAND2_X1 U5488 ( .A1(n6399), .A2(n5147), .ZN(n4398) );
  NAND2_X1 U5489 ( .A1(n4398), .A2(n4397), .ZN(n4399) );
  NAND2_X1 U5490 ( .A1(n5962), .A2(n4399), .ZN(n6072) );
  INV_X1 U5491 ( .A(n6072), .ZN(n4400) );
  OAI21_X1 U5492 ( .B1(n6414), .B2(n5947), .A(n4400), .ZN(n5944) );
  AOI21_X1 U5493 ( .B1(n5930), .B2(n6090), .A(n5944), .ZN(n5567) );
  OAI21_X1 U5494 ( .B1(n4401), .B2(n6414), .A(n5567), .ZN(n5534) );
  OAI21_X1 U5495 ( .B1(n4406), .B2(n6425), .A(n4405), .ZN(U2987) );
  NAND2_X1 U5496 ( .A1(n5628), .A2(n4414), .ZN(n4415) );
  NAND2_X1 U5497 ( .A1(n5616), .A2(n4415), .ZN(n5940) );
  OAI22_X1 U5498 ( .A1(n5853), .A2(n6171), .B1(n5940), .B2(n6257), .ZN(n4424)
         );
  AOI22_X1 U5499 ( .A1(EBX_REG_27__SCAN_IN), .A2(n6264), .B1(n5856), .B2(n6196), .ZN(n4422) );
  AND3_X1 U5500 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4417) );
  NAND2_X1 U5501 ( .A1(n4416), .A2(n4417), .ZN(n4425) );
  INV_X1 U5502 ( .A(n4425), .ZN(n5618) );
  INV_X1 U5503 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6680) );
  INV_X1 U5504 ( .A(n4417), .ZN(n4418) );
  NAND2_X1 U5505 ( .A1(n6246), .A2(n4418), .ZN(n4419) );
  NAND2_X1 U5506 ( .A1(n5657), .A2(n4419), .ZN(n5632) );
  NAND3_X1 U5507 ( .A1(n4422), .A2(n3162), .A3(n4421), .ZN(n4423) );
  NAND2_X1 U5508 ( .A1(n5818), .A2(n6220), .ZN(n4436) );
  NAND2_X1 U5509 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4426) );
  OR2_X1 U5510 ( .A1(n4425), .A2(n4426), .ZN(n5608) );
  AND2_X1 U5511 ( .A1(REIP_REG_30__SCAN_IN), .A2(REIP_REG_29__SCAN_IN), .ZN(
        n4429) );
  AOI21_X1 U5512 ( .B1(n6246), .B2(n4426), .A(n5632), .ZN(n5622) );
  OAI21_X1 U5513 ( .B1(n5608), .B2(n4429), .A(n5622), .ZN(n5594) );
  OAI22_X1 U5514 ( .A1(n5514), .A2(n4428), .B1(n6253), .B2(n4427), .ZN(n4432)
         );
  INV_X1 U5515 ( .A(n4429), .ZN(n4430) );
  NOR3_X1 U5516 ( .A1(n5608), .A2(REIP_REG_31__SCAN_IN), .A3(n4430), .ZN(n4431) );
  AOI211_X1 U5517 ( .C1(REIP_REG_31__SCAN_IN), .C2(n5594), .A(n4432), .B(n4431), .ZN(n4433) );
  NAND2_X1 U5518 ( .A1(n4436), .A2(n4435), .ZN(U2796) );
  INV_X1 U5519 ( .A(n6037), .ZN(n5637) );
  NAND2_X1 U5520 ( .A1(n5637), .A2(n6347), .ZN(n4449) );
  XNOR2_X1 U5521 ( .A(n5989), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4443)
         );
  XNOR2_X1 U5522 ( .A(n4442), .B(n4443), .ZN(n5955) );
  NAND2_X1 U5523 ( .A1(n3952), .A2(REIP_REG_26__SCAN_IN), .ZN(n5950) );
  NAND2_X1 U5524 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4444)
         );
  OAI211_X1 U5525 ( .C1(n6352), .C2(n5629), .A(n5950), .B(n4444), .ZN(n4445)
         );
  NAND2_X1 U5526 ( .A1(n4449), .A2(n4448), .ZN(U2960) );
  INV_X1 U5527 ( .A(n4450), .ZN(n4468) );
  INV_X1 U5528 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n4453) );
  NAND2_X1 U5529 ( .A1(n4451), .A2(n3169), .ZN(n4467) );
  INV_X1 U5530 ( .A(n4467), .ZN(n4452) );
  OAI21_X1 U5531 ( .B1(n4468), .B2(n4453), .A(n4452), .ZN(U2788) );
  NOR2_X1 U5532 ( .A1(n6601), .A2(n3146), .ZN(n4454) );
  AOI21_X1 U5533 ( .B1(n4455), .B2(n4602), .A(n4454), .ZN(n6115) );
  OR2_X1 U5534 ( .A1(n5295), .A2(n4456), .ZN(n4470) );
  NAND2_X1 U5535 ( .A1(n4470), .A2(n6596), .ZN(n4457) );
  NAND2_X1 U5536 ( .A1(n4457), .A2(n6630), .ZN(n6733) );
  AND2_X1 U5537 ( .A1(n6115), .A2(n6733), .ZN(n6567) );
  NOR2_X1 U5538 ( .A1(n6567), .A2(n6612), .ZN(n6123) );
  INV_X1 U5539 ( .A(MORE_REG_SCAN_IN), .ZN(n4466) );
  NAND2_X1 U5540 ( .A1(n6569), .A2(n4602), .ZN(n4458) );
  NOR2_X1 U5541 ( .A1(n4458), .A2(n4569), .ZN(n4459) );
  MUX2_X1 U5542 ( .A(n4459), .B(n4697), .S(n6601), .Z(n4463) );
  NAND2_X1 U5543 ( .A1(n4461), .A2(n4460), .ZN(n4462) );
  AND2_X1 U5544 ( .A1(n4463), .A2(n4462), .ZN(n6570) );
  INV_X1 U5545 ( .A(n6570), .ZN(n4464) );
  NAND2_X1 U5546 ( .A1(n4464), .A2(n6123), .ZN(n4465) );
  OAI21_X1 U5547 ( .B1(n6123), .B2(n4466), .A(n4465), .ZN(U3471) );
  NOR3_X1 U5548 ( .A1(n4468), .A2(READREQUEST_REG_SCAN_IN), .A3(n4467), .ZN(
        n4469) );
  AOI21_X1 U5549 ( .B1(n6732), .B2(n4470), .A(n4469), .ZN(U3474) );
  NOR2_X1 U5550 ( .A1(n4602), .A2(READY_N), .ZN(n4471) );
  NAND2_X1 U5551 ( .A1(n4568), .A2(n4471), .ZN(n4473) );
  INV_X1 U5552 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n4475) );
  INV_X1 U5553 ( .A(DATAI_0_), .ZN(n4690) );
  NOR2_X1 U5554 ( .A1(n6316), .A2(n4690), .ZN(n4476) );
  AOI21_X1 U5555 ( .B1(n6330), .B2(EAX_REG_0__SCAN_IN), .A(n4476), .ZN(n4474)
         );
  OAI21_X1 U5556 ( .B1(n6333), .B2(n4475), .A(n4474), .ZN(U2939) );
  INV_X1 U5557 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n4478) );
  AOI21_X1 U5558 ( .B1(n6330), .B2(EAX_REG_16__SCAN_IN), .A(n4476), .ZN(n4477)
         );
  OAI21_X1 U5559 ( .B1(n6333), .B2(n4478), .A(n4477), .ZN(U2924) );
  INV_X1 U5560 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n4480) );
  INV_X1 U5561 ( .A(DATAI_7_), .ZN(n5049) );
  NOR2_X1 U5562 ( .A1(n6316), .A2(n5049), .ZN(n4498) );
  AOI21_X1 U5563 ( .B1(n6330), .B2(EAX_REG_7__SCAN_IN), .A(n4498), .ZN(n4479)
         );
  OAI21_X1 U5564 ( .B1(n6333), .B2(n4480), .A(n4479), .ZN(U2946) );
  INV_X1 U5565 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n4482) );
  INV_X1 U5566 ( .A(DATAI_6_), .ZN(n5039) );
  NOR2_X1 U5567 ( .A1(n6316), .A2(n5039), .ZN(n4492) );
  AOI21_X1 U5568 ( .B1(n6330), .B2(EAX_REG_6__SCAN_IN), .A(n4492), .ZN(n4481)
         );
  OAI21_X1 U5569 ( .B1(n6333), .B2(n4482), .A(n4481), .ZN(U2945) );
  INV_X1 U5570 ( .A(LWORD_REG_11__SCAN_IN), .ZN(n4484) );
  INV_X1 U5571 ( .A(DATAI_11_), .ZN(n6844) );
  NOR2_X1 U5572 ( .A1(n6316), .A2(n6844), .ZN(n4485) );
  AOI21_X1 U5573 ( .B1(n6330), .B2(EAX_REG_11__SCAN_IN), .A(n4485), .ZN(n4483)
         );
  OAI21_X1 U5574 ( .B1(n6333), .B2(n4484), .A(n4483), .ZN(U2950) );
  INV_X1 U5575 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n4487) );
  AOI21_X1 U5576 ( .B1(n6330), .B2(EAX_REG_27__SCAN_IN), .A(n4485), .ZN(n4486)
         );
  OAI21_X1 U5577 ( .B1(n6333), .B2(n4487), .A(n4486), .ZN(U2935) );
  INV_X1 U5578 ( .A(LWORD_REG_3__SCAN_IN), .ZN(n4489) );
  INV_X1 U5579 ( .A(DATAI_3_), .ZN(n4678) );
  NOR2_X1 U5580 ( .A1(n6316), .A2(n4678), .ZN(n4495) );
  AOI21_X1 U5581 ( .B1(n6330), .B2(EAX_REG_3__SCAN_IN), .A(n4495), .ZN(n4488)
         );
  OAI21_X1 U5582 ( .B1(n6333), .B2(n4489), .A(n4488), .ZN(U2942) );
  INV_X1 U5583 ( .A(UWORD_REG_5__SCAN_IN), .ZN(n4491) );
  INV_X1 U5584 ( .A(DATAI_5_), .ZN(n4799) );
  NOR2_X1 U5585 ( .A1(n6316), .A2(n4799), .ZN(n4501) );
  AOI21_X1 U5586 ( .B1(n6330), .B2(EAX_REG_21__SCAN_IN), .A(n4501), .ZN(n4490)
         );
  OAI21_X1 U5587 ( .B1(n6333), .B2(n4491), .A(n4490), .ZN(U2929) );
  INV_X1 U5588 ( .A(UWORD_REG_6__SCAN_IN), .ZN(n4494) );
  AOI21_X1 U5589 ( .B1(n6330), .B2(EAX_REG_22__SCAN_IN), .A(n4492), .ZN(n4493)
         );
  OAI21_X1 U5590 ( .B1(n6333), .B2(n4494), .A(n4493), .ZN(U2930) );
  INV_X1 U5591 ( .A(UWORD_REG_3__SCAN_IN), .ZN(n4497) );
  AOI21_X1 U5592 ( .B1(n6330), .B2(EAX_REG_19__SCAN_IN), .A(n4495), .ZN(n4496)
         );
  OAI21_X1 U5593 ( .B1(n6333), .B2(n4497), .A(n4496), .ZN(U2927) );
  INV_X1 U5594 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n4500) );
  AOI21_X1 U5595 ( .B1(n6330), .B2(EAX_REG_23__SCAN_IN), .A(n4498), .ZN(n4499)
         );
  OAI21_X1 U5596 ( .B1(n6333), .B2(n4500), .A(n4499), .ZN(U2931) );
  AOI21_X1 U5597 ( .B1(n6330), .B2(EAX_REG_5__SCAN_IN), .A(n4501), .ZN(n4502)
         );
  OAI21_X1 U5598 ( .B1(n6333), .B2(n6297), .A(n4502), .ZN(U2944) );
  NAND2_X1 U5599 ( .A1(n6331), .A2(DATAI_4_), .ZN(n4517) );
  NAND2_X1 U5600 ( .A1(n6327), .A2(UWORD_REG_4__SCAN_IN), .ZN(n4503) );
  OAI211_X1 U5601 ( .C1(n6329), .C2(n4504), .A(n4517), .B(n4503), .ZN(U2928)
         );
  NAND2_X1 U5602 ( .A1(n6331), .A2(DATAI_2_), .ZN(n4520) );
  NAND2_X1 U5603 ( .A1(n6327), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4505) );
  OAI211_X1 U5604 ( .C1(n6329), .C2(n4506), .A(n4520), .B(n4505), .ZN(U2926)
         );
  NAND2_X1 U5605 ( .A1(n6331), .A2(DATAI_13_), .ZN(n4515) );
  NAND2_X1 U5606 ( .A1(n6327), .A2(UWORD_REG_13__SCAN_IN), .ZN(n4507) );
  OAI211_X1 U5607 ( .C1(n6329), .C2(n4508), .A(n4515), .B(n4507), .ZN(U2937)
         );
  INV_X1 U5608 ( .A(EAX_REG_1__SCAN_IN), .ZN(n4510) );
  NAND2_X1 U5609 ( .A1(n6331), .A2(DATAI_1_), .ZN(n4512) );
  NAND2_X1 U5610 ( .A1(n6327), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4509) );
  OAI211_X1 U5611 ( .C1(n6329), .C2(n4510), .A(n4512), .B(n4509), .ZN(U2940)
         );
  NAND2_X1 U5612 ( .A1(n6327), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4511) );
  OAI211_X1 U5613 ( .C1(n6329), .C2(n4513), .A(n4512), .B(n4511), .ZN(U2925)
         );
  INV_X1 U5614 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5482) );
  NAND2_X1 U5615 ( .A1(n6327), .A2(LWORD_REG_13__SCAN_IN), .ZN(n4514) );
  OAI211_X1 U5616 ( .C1(n6329), .C2(n5482), .A(n4515), .B(n4514), .ZN(U2952)
         );
  INV_X1 U5617 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n4518) );
  NAND2_X1 U5618 ( .A1(n6330), .A2(EAX_REG_4__SCAN_IN), .ZN(n4516) );
  OAI211_X1 U5619 ( .C1(n6333), .C2(n4518), .A(n4517), .B(n4516), .ZN(U2943)
         );
  INV_X1 U5620 ( .A(LWORD_REG_2__SCAN_IN), .ZN(n4521) );
  NAND2_X1 U5621 ( .A1(n6330), .A2(EAX_REG_2__SCAN_IN), .ZN(n4519) );
  OAI211_X1 U5622 ( .C1(n6333), .C2(n4521), .A(n4520), .B(n4519), .ZN(U2941)
         );
  NAND2_X1 U5623 ( .A1(n6576), .A2(n4568), .ZN(n4522) );
  NAND2_X1 U5624 ( .A1(n4522), .A2(n6329), .ZN(n4523) );
  NAND2_X1 U5625 ( .A1(n6609), .A2(n4647), .ZN(n6730) );
  INV_X1 U5626 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n6757) );
  NAND2_X1 U5627 ( .A1(n6298), .A2(n3962), .ZN(n6276) );
  INV_X1 U5628 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4524) );
  OAI222_X1 U5629 ( .A1(n6301), .A2(n6757), .B1(n6276), .B2(n4524), .C1(n4491), 
        .C2(n6730), .ZN(U2902) );
  INV_X1 U5630 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6313) );
  INV_X1 U5631 ( .A(UWORD_REG_10__SCAN_IN), .ZN(n4525) );
  INV_X1 U5632 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n6943) );
  OAI222_X1 U5633 ( .A1(n6276), .A2(n6313), .B1(n6730), .B2(n4525), .C1(n6301), 
        .C2(n6943), .ZN(U2897) );
  INV_X1 U5634 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6849) );
  AOI22_X1 U5635 ( .A1(n6305), .A2(UWORD_REG_14__SCAN_IN), .B1(n6304), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4526) );
  OAI21_X1 U5636 ( .B1(n6849), .B2(n6276), .A(n4526), .ZN(U2893) );
  INV_X1 U5637 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4528) );
  AOI22_X1 U5638 ( .A1(n6305), .A2(UWORD_REG_0__SCAN_IN), .B1(n6304), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4527) );
  OAI21_X1 U5639 ( .B1(n4528), .B2(n6276), .A(n4527), .ZN(U2907) );
  AOI22_X1 U5640 ( .A1(n6305), .A2(UWORD_REG_1__SCAN_IN), .B1(n6304), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4529) );
  OAI21_X1 U5641 ( .B1(n4513), .B2(n6276), .A(n4529), .ZN(U2906) );
  INV_X1 U5642 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4531) );
  AOI22_X1 U5643 ( .A1(n6305), .A2(UWORD_REG_3__SCAN_IN), .B1(n6304), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4530) );
  OAI21_X1 U5644 ( .B1(n4531), .B2(n6276), .A(n4530), .ZN(U2904) );
  INV_X1 U5645 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6814) );
  AOI22_X1 U5646 ( .A1(n6305), .A2(UWORD_REG_6__SCAN_IN), .B1(n6304), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4532) );
  OAI21_X1 U5647 ( .B1(n6814), .B2(n6276), .A(n4532), .ZN(U2901) );
  INV_X1 U5648 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4534) );
  AOI22_X1 U5649 ( .A1(n6305), .A2(UWORD_REG_7__SCAN_IN), .B1(n6304), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4533) );
  OAI21_X1 U5650 ( .B1(n4534), .B2(n6276), .A(n4533), .ZN(U2900) );
  AOI22_X1 U5651 ( .A1(n6305), .A2(UWORD_REG_8__SCAN_IN), .B1(n6304), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4535) );
  OAI21_X1 U5652 ( .B1(n3864), .B2(n6276), .A(n4535), .ZN(U2899) );
  AOI22_X1 U5653 ( .A1(n6305), .A2(UWORD_REG_9__SCAN_IN), .B1(n6304), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4536) );
  OAI21_X1 U5654 ( .B1(n3882), .B2(n6276), .A(n4536), .ZN(U2898) );
  INV_X1 U5655 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4538) );
  AOI22_X1 U5656 ( .A1(n6305), .A2(UWORD_REG_12__SCAN_IN), .B1(n6304), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4537) );
  OAI21_X1 U5657 ( .B1(n4538), .B2(n6276), .A(n4537), .ZN(U2895) );
  OAI21_X1 U5658 ( .B1(n4541), .B2(n4540), .A(n4539), .ZN(n5760) );
  OR2_X1 U5659 ( .A1(n4543), .A2(n4542), .ZN(n4545) );
  AND2_X1 U5660 ( .A1(n4545), .A2(n4544), .ZN(n6421) );
  AOI22_X1 U5661 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n3952), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4548) );
  INV_X1 U5662 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4546) );
  NAND2_X1 U5663 ( .A1(n6336), .A2(n4546), .ZN(n4547) );
  NAND2_X1 U5664 ( .A1(n4548), .A2(n4547), .ZN(n4549) );
  AOI21_X1 U5665 ( .B1(n6421), .B2(n4310), .A(n4549), .ZN(n4550) );
  OAI21_X1 U5666 ( .B1(n6361), .B2(n5760), .A(n4550), .ZN(U2985) );
  NOR2_X1 U5667 ( .A1(n4552), .A2(n4553), .ZN(n4554) );
  OR2_X1 U5668 ( .A1(n4551), .A2(n4554), .ZN(n6261) );
  XOR2_X1 U5669 ( .A(n4556), .B(n4555), .Z(n6396) );
  NAND2_X1 U5670 ( .A1(n6396), .A2(n4310), .ZN(n4560) );
  NAND2_X1 U5671 ( .A1(n3952), .A2(REIP_REG_3__SCAN_IN), .ZN(n6392) );
  INV_X1 U5672 ( .A(n6392), .ZN(n4558) );
  NOR2_X1 U5673 ( .A1(n6352), .A2(n6259), .ZN(n4557) );
  AOI211_X1 U5674 ( .C1(n6358), .C2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4558), 
        .B(n4557), .ZN(n4559) );
  OAI211_X1 U5675 ( .C1(n6361), .C2(n6261), .A(n4560), .B(n4559), .ZN(U2983)
         );
  INV_X1 U5676 ( .A(n4561), .ZN(n4562) );
  OR2_X1 U5677 ( .A1(n6108), .A2(n4562), .ZN(n4608) );
  INV_X1 U5678 ( .A(n4563), .ZN(n4567) );
  NAND3_X1 U5679 ( .A1(n5815), .A2(n4565), .A3(n4564), .ZN(n4698) );
  NOR2_X1 U5680 ( .A1(n4698), .A2(n4699), .ZN(n4566) );
  NAND2_X1 U5681 ( .A1(n4196), .A2(n4705), .ZN(n4571) );
  NAND2_X2 U5682 ( .A1(n5816), .A2(n4571), .ZN(n5834) );
  INV_X1 U5683 ( .A(n4571), .ZN(n4572) );
  INV_X1 U5684 ( .A(DATAI_1_), .ZN(n4684) );
  OAI222_X1 U5685 ( .A1(n5760), .A2(n5834), .B1(n5481), .B2(n4684), .C1(n5816), 
        .C2(n4510), .ZN(U2890) );
  NOR2_X1 U5686 ( .A1(n4551), .A2(n4574), .ZN(n4575) );
  OR2_X1 U5687 ( .A1(n4573), .A2(n4575), .ZN(n6242) );
  INV_X1 U5688 ( .A(DATAI_4_), .ZN(n6918) );
  INV_X1 U5689 ( .A(EAX_REG_4__SCAN_IN), .ZN(n7013) );
  OAI222_X1 U5690 ( .A1(n6242), .A2(n5834), .B1(n5481), .B2(n6918), .C1(n5816), 
        .C2(n7013), .ZN(U2887) );
  INV_X1 U5691 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6300) );
  OAI222_X1 U5692 ( .A1(n6261), .A2(n5834), .B1(n5481), .B2(n4678), .C1(n5816), 
        .C2(n6300), .ZN(U2888) );
  NOR2_X1 U5693 ( .A1(n4577), .A2(n4576), .ZN(n4578) );
  OR2_X1 U5694 ( .A1(n4552), .A2(n4578), .ZN(n6346) );
  INV_X1 U5695 ( .A(DATAI_2_), .ZN(n4655) );
  INV_X1 U5696 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6953) );
  OAI222_X1 U5697 ( .A1(n6346), .A2(n5834), .B1(n5481), .B2(n4655), .C1(n5816), 
        .C2(n6953), .ZN(U2889) );
  OAI21_X1 U5698 ( .B1(n4581), .B2(n4580), .A(n4579), .ZN(n6362) );
  INV_X1 U5699 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6308) );
  OAI222_X1 U5700 ( .A1(n6362), .A2(n5834), .B1(n5481), .B2(n4690), .C1(n5816), 
        .C2(n6308), .ZN(U2891) );
  OR2_X1 U5701 ( .A1(n4573), .A2(n4582), .ZN(n4584) );
  NAND2_X1 U5702 ( .A1(n4584), .A2(n4583), .ZN(n6228) );
  INV_X1 U5703 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6296) );
  OAI222_X1 U5704 ( .A1(n6228), .A2(n5834), .B1(n5481), .B2(n4799), .C1(n5816), 
        .C2(n6296), .ZN(U2886) );
  NAND2_X1 U5705 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4647), .ZN(n6699) );
  NAND4_X1 U5706 ( .A1(n4587), .A2(n6108), .A3(n4586), .A4(n4563), .ZN(n4589)
         );
  NOR2_X1 U5707 ( .A1(n4589), .A2(n4588), .ZN(n5554) );
  INV_X1 U5708 ( .A(n5554), .ZN(n6574) );
  NAND2_X1 U5709 ( .A1(n6439), .A2(n6574), .ZN(n4599) );
  NAND2_X1 U5710 ( .A1(n4697), .A2(n4601), .ZN(n4620) );
  MUX2_X1 U5711 ( .A(n3178), .B(n6988), .S(n5551), .Z(n4590) );
  NOR2_X1 U5712 ( .A1(n4590), .A2(n4627), .ZN(n4597) );
  INV_X1 U5713 ( .A(n3178), .ZN(n4591) );
  OAI211_X1 U5714 ( .C1(n6988), .C2(n5551), .A(n3474), .B(n4591), .ZN(n6704)
         );
  XNOR2_X1 U5715 ( .A(n4593), .B(n4592), .ZN(n4594) );
  NAND2_X1 U5716 ( .A1(n6576), .A2(n4594), .ZN(n4595) );
  OAI21_X1 U5717 ( .B1(n6704), .B2(n4617), .A(n4595), .ZN(n4596) );
  AOI21_X1 U5718 ( .B1(n4620), .B2(n4597), .A(n4596), .ZN(n4598) );
  NAND2_X1 U5719 ( .A1(n4599), .A2(n4598), .ZN(n6703) );
  INV_X1 U5720 ( .A(n6601), .ZN(n4600) );
  MUX2_X1 U5721 ( .A(n4601), .B(n4697), .S(n4600), .Z(n4613) );
  INV_X1 U5722 ( .A(n4602), .ZN(n4606) );
  NAND2_X1 U5723 ( .A1(n6576), .A2(n6630), .ZN(n4604) );
  NAND2_X1 U5724 ( .A1(n4604), .A2(n4603), .ZN(n4605) );
  OAI211_X1 U5725 ( .C1(n4606), .C2(n6627), .A(n4605), .B(n6601), .ZN(n4611)
         );
  INV_X1 U5726 ( .A(n4607), .ZN(n4609) );
  AND4_X1 U5727 ( .A1(n4611), .A2(n4610), .A3(n4609), .A4(n4608), .ZN(n4612)
         );
  MUX2_X1 U5728 ( .A(n6703), .B(n6988), .S(n6582), .Z(n6592) );
  XNOR2_X1 U5729 ( .A(n5551), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4619)
         );
  XNOR2_X1 U5730 ( .A(n5560), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4615)
         );
  NAND2_X1 U5731 ( .A1(n6576), .A2(n4615), .ZN(n4616) );
  OAI21_X1 U5732 ( .B1(n4619), .B2(n4617), .A(n4616), .ZN(n4618) );
  AOI21_X1 U5733 ( .B1(n4620), .B2(n4619), .A(n4618), .ZN(n4621) );
  OAI21_X1 U5734 ( .B1(n6014), .B2(n5554), .A(n4621), .ZN(n5547) );
  OR2_X1 U5735 ( .A1(n5547), .A2(n6582), .ZN(n4624) );
  NAND2_X1 U5736 ( .A1(n6582), .A2(n4622), .ZN(n4623) );
  NAND2_X1 U5737 ( .A1(n4624), .A2(n4623), .ZN(n6584) );
  NOR2_X1 U5738 ( .A1(n6584), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4625) );
  NAND2_X1 U5739 ( .A1(n6592), .A2(n4625), .ZN(n4629) );
  INV_X1 U5740 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6122) );
  NAND2_X1 U5741 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6122), .ZN(n4633) );
  INV_X1 U5742 ( .A(n4633), .ZN(n4626) );
  NAND2_X1 U5743 ( .A1(n4627), .A2(n4626), .ZN(n4628) );
  NAND2_X1 U5744 ( .A1(n4629), .A2(n4628), .ZN(n6573) );
  INV_X1 U5745 ( .A(n3177), .ZN(n4630) );
  NAND2_X1 U5746 ( .A1(n6573), .A2(n4630), .ZN(n4649) );
  INV_X1 U5747 ( .A(n4897), .ZN(n4654) );
  NOR2_X1 U5748 ( .A1(n4631), .A2(n4654), .ZN(n4632) );
  XNOR2_X1 U5749 ( .A(n4632), .B(n6113), .ZN(n6234) );
  NOR2_X1 U5750 ( .A1(n6108), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4636) );
  NAND2_X1 U5751 ( .A1(n6582), .A2(n6709), .ZN(n4634) );
  AOI21_X1 U5752 ( .B1(n4634), .B2(n4633), .A(n6113), .ZN(n4635) );
  AOI21_X1 U5753 ( .B1(n6234), .B2(n4636), .A(n4635), .ZN(n6571) );
  INV_X1 U5754 ( .A(n5381), .ZN(n6506) );
  INV_X1 U5755 ( .A(n4674), .ZN(n4641) );
  NAND2_X1 U5756 ( .A1(n4641), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4670) );
  NAND2_X1 U5757 ( .A1(n6506), .A2(n4670), .ZN(n5067) );
  INV_X1 U5758 ( .A(n5067), .ZN(n4643) );
  NAND2_X1 U5759 ( .A1(n4640), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6505) );
  OR2_X1 U5760 ( .A1(n4713), .A2(n6505), .ZN(n4653) );
  AOI21_X1 U5761 ( .B1(n4643), .B2(n4653), .A(n6729), .ZN(n4645) );
  NAND2_X1 U5762 ( .A1(n6442), .A2(n6121), .ZN(n6444) );
  AND2_X1 U5763 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6702), .ZN(n6013) );
  OAI22_X1 U5764 ( .A1(n4730), .A2(n6444), .B1(n6254), .B2(n6013), .ZN(n4644)
         );
  OAI21_X1 U5765 ( .B1(n4645), .B2(n4644), .A(n6435), .ZN(n4646) );
  OAI21_X1 U5766 ( .B1(n6435), .B2(n7014), .A(n4646), .ZN(U3462) );
  AND2_X1 U5767 ( .A1(n6571), .A2(n4647), .ZN(n4648) );
  NAND2_X1 U5768 ( .A1(n4649), .A2(n4648), .ZN(n6608) );
  INV_X1 U5769 ( .A(n6608), .ZN(n4651) );
  OAI22_X1 U5770 ( .A1(n5379), .A2(n6729), .B1(n5297), .B2(n6013), .ZN(n4650)
         );
  OAI21_X1 U5771 ( .B1(n4651), .B2(n4650), .A(n6435), .ZN(n4652) );
  OAI21_X1 U5772 ( .B1(n6435), .B2(n4838), .A(n4652), .ZN(U3465) );
  NAND2_X1 U5773 ( .A1(n4653), .A2(n6442), .ZN(n4659) );
  NOR2_X1 U5774 ( .A1(n6014), .A2(n6010), .ZN(n5112) );
  AND2_X1 U5775 ( .A1(n5112), .A2(n4654), .ZN(n6443) );
  INV_X1 U5776 ( .A(n5297), .ZN(n6575) );
  INV_X1 U5777 ( .A(n5041), .ZN(n6496) );
  AOI21_X1 U5778 ( .B1(n6443), .B2(n6575), .A(n6496), .ZN(n4656) );
  OAI22_X1 U5779 ( .A1(n4659), .A2(n4656), .B1(n6441), .B2(n6935), .ZN(n6497)
         );
  INV_X1 U5780 ( .A(n6497), .ZN(n5045) );
  INV_X1 U5781 ( .A(n4656), .ZN(n4658) );
  AOI21_X1 U5782 ( .B1(n6729), .B2(n6441), .A(n6508), .ZN(n4657) );
  OAI21_X1 U5783 ( .B1(n4659), .B2(n4658), .A(n4657), .ZN(n6498) );
  INV_X1 U5784 ( .A(n6495), .ZN(n5233) );
  INV_X1 U5785 ( .A(DATAI_18_), .ZN(n6901) );
  OR2_X1 U5786 ( .A1(n6361), .A2(n6901), .ZN(n6462) );
  INV_X1 U5787 ( .A(DATAI_26_), .ZN(n6035) );
  OR2_X1 U5788 ( .A1(n6361), .A2(n6035), .ZN(n6529) );
  OAI22_X1 U5789 ( .A1(n5233), .A2(n6462), .B1(n6529), .B2(n6501), .ZN(n4664)
         );
  NOR2_X1 U5790 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6702), .ZN(n5542) );
  NOR2_X2 U5791 ( .A1(n4806), .A2(n4662), .ZN(n6525) );
  INV_X1 U5792 ( .A(n6525), .ZN(n5406) );
  NOR2_X1 U5793 ( .A1(n5406), .A2(n5041), .ZN(n4663) );
  AOI211_X1 U5794 ( .C1(INSTQUEUE_REG_7__2__SCAN_IN), .C2(n6498), .A(n4664), 
        .B(n4663), .ZN(n4665) );
  OAI21_X1 U5795 ( .B1(n5045), .B2(n5409), .A(n4665), .ZN(U3078) );
  NOR2_X2 U5796 ( .A1(n4806), .A2(n5815), .ZN(n6559) );
  INV_X1 U5797 ( .A(n6559), .ZN(n5391) );
  NAND3_X1 U5798 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6579), .ZN(n4899) );
  NOR2_X1 U5799 ( .A1(n4838), .A2(n4899), .ZN(n4667) );
  INV_X1 U5800 ( .A(n4667), .ZN(n4880) );
  INV_X1 U5801 ( .A(n4899), .ZN(n4669) );
  INV_X1 U5802 ( .A(n6014), .ZN(n4666) );
  NAND2_X1 U5803 ( .A1(n4666), .A2(n6010), .ZN(n4716) );
  INV_X1 U5804 ( .A(n4716), .ZN(n4898) );
  AOI21_X1 U5805 ( .B1(n4898), .B2(n4956), .A(n4667), .ZN(n4672) );
  NAND3_X1 U5806 ( .A1(n6442), .A2(n4672), .A3(n4670), .ZN(n4668) );
  OAI211_X1 U5807 ( .C1(n6442), .C2(n4669), .A(n4959), .B(n4668), .ZN(n4877)
         );
  NAND2_X1 U5808 ( .A1(n6442), .A2(n4670), .ZN(n4671) );
  OAI22_X1 U5809 ( .A1(n4672), .A2(n4671), .B1(n6935), .B2(n4899), .ZN(n4876)
         );
  AOI22_X1 U5810 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4877), .B1(n6561), 
        .B2(n4876), .ZN(n4677) );
  INV_X1 U5811 ( .A(DATAI_31_), .ZN(n4673) );
  OR2_X1 U5812 ( .A1(n6361), .A2(n4673), .ZN(n6566) );
  INV_X1 U5813 ( .A(n6566), .ZN(n6478) );
  INV_X1 U5814 ( .A(DATAI_23_), .ZN(n4675) );
  OR2_X1 U5815 ( .A1(n6361), .A2(n4675), .ZN(n6482) );
  INV_X1 U5816 ( .A(n6482), .ZN(n6556) );
  AOI22_X1 U5817 ( .A1(n6478), .A2(n4895), .B1(n5113), .B2(n6556), .ZN(n4676)
         );
  OAI211_X1 U5818 ( .C1(n5391), .C2(n4880), .A(n4677), .B(n4676), .ZN(U3131)
         );
  NOR2_X2 U5819 ( .A1(n4806), .A2(n3136), .ZN(n6531) );
  INV_X1 U5820 ( .A(n6531), .ZN(n5411) );
  AOI22_X1 U5821 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4877), .B1(n6532), 
        .B2(n4876), .ZN(n4682) );
  INV_X1 U5822 ( .A(DATAI_27_), .ZN(n4679) );
  OR2_X1 U5823 ( .A1(n6361), .A2(n4679), .ZN(n6535) );
  INV_X1 U5824 ( .A(n6535), .ZN(n6463) );
  INV_X1 U5825 ( .A(DATAI_19_), .ZN(n4680) );
  OR2_X1 U5826 ( .A1(n6361), .A2(n4680), .ZN(n6466) );
  INV_X1 U5827 ( .A(n6466), .ZN(n6530) );
  AOI22_X1 U5828 ( .A1(n6463), .A2(n4895), .B1(n5113), .B2(n6530), .ZN(n4681)
         );
  OAI211_X1 U5829 ( .C1(n5411), .C2(n4880), .A(n4682), .B(n4681), .ZN(U3127)
         );
  NOR2_X2 U5830 ( .A1(n4806), .A2(n4683), .ZN(n6519) );
  INV_X1 U5831 ( .A(n6519), .ZN(n5422) );
  AOI22_X1 U5832 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4877), .B1(n6520), 
        .B2(n4876), .ZN(n4688) );
  INV_X1 U5833 ( .A(DATAI_25_), .ZN(n4685) );
  OR2_X1 U5834 ( .A1(n6361), .A2(n4685), .ZN(n6523) );
  INV_X1 U5835 ( .A(n6523), .ZN(n6455) );
  INV_X1 U5836 ( .A(DATAI_17_), .ZN(n4686) );
  OR2_X1 U5837 ( .A1(n6361), .A2(n4686), .ZN(n6458) );
  INV_X1 U5838 ( .A(n6458), .ZN(n6518) );
  AOI22_X1 U5839 ( .A1(n6455), .A2(n4895), .B1(n5113), .B2(n6518), .ZN(n4687)
         );
  OAI211_X1 U5840 ( .C1(n5422), .C2(n4880), .A(n4688), .B(n4687), .ZN(U3125)
         );
  NOR2_X2 U5841 ( .A1(n4806), .A2(n4689), .ZN(n6504) );
  INV_X1 U5842 ( .A(n6504), .ZN(n5429) );
  AOI22_X1 U5843 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4877), .B1(n6514), 
        .B2(n4876), .ZN(n4693) );
  INV_X1 U5844 ( .A(DATAI_24_), .ZN(n4691) );
  OR2_X1 U5845 ( .A1(n6361), .A2(n4691), .ZN(n6517) );
  INV_X1 U5846 ( .A(n6517), .ZN(n6451) );
  INV_X1 U5847 ( .A(DATAI_16_), .ZN(n6817) );
  OR2_X1 U5848 ( .A1(n6361), .A2(n6817), .ZN(n6454) );
  INV_X1 U5849 ( .A(n6454), .ZN(n6503) );
  AOI22_X1 U5850 ( .A1(n6451), .A2(n4895), .B1(n5113), .B2(n6503), .ZN(n4692)
         );
  OAI211_X1 U5851 ( .C1(n5429), .C2(n4880), .A(n4693), .B(n4692), .ZN(U3124)
         );
  AOI22_X1 U5852 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4877), .B1(n6526), 
        .B2(n4876), .ZN(n4695) );
  INV_X1 U5853 ( .A(n6529), .ZN(n6459) );
  INV_X1 U5854 ( .A(n6462), .ZN(n6524) );
  AOI22_X1 U5855 ( .A1(n6459), .A2(n4895), .B1(n5113), .B2(n6524), .ZN(n4694)
         );
  OAI211_X1 U5856 ( .C1(n5406), .C2(n4880), .A(n4695), .B(n4694), .ZN(U3126)
         );
  OR2_X1 U5857 ( .A1(n6601), .A2(n6612), .ZN(n4696) );
  INV_X1 U5858 ( .A(n4698), .ZN(n4702) );
  INV_X1 U5859 ( .A(n4699), .ZN(n4700) );
  NAND4_X1 U5860 ( .A1(n4702), .A2(n4701), .A3(n4700), .A4(n4931), .ZN(n4703)
         );
  INV_X2 U5861 ( .A(n5810), .ZN(n5796) );
  INV_X1 U5862 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4709) );
  CLKBUF_X1 U5863 ( .A(n4708), .Z(n4756) );
  OAI21_X1 U5864 ( .B1(n3991), .B2(n3990), .A(n4756), .ZN(n6225) );
  OAI222_X1 U5865 ( .A1(n6228), .A2(n5796), .B1(n5814), .B2(n4709), .C1(n6225), 
        .C2(n5808), .ZN(U2854) );
  NOR2_X1 U5866 ( .A1(n4716), .A2(n6729), .ZN(n4893) );
  NOR2_X1 U5867 ( .A1(n4711), .A2(n6935), .ZN(n6437) );
  INV_X1 U5868 ( .A(n4710), .ZN(n4891) );
  INV_X1 U5869 ( .A(n5384), .ZN(n6436) );
  NOR2_X1 U5870 ( .A1(n4891), .A2(n6436), .ZN(n5155) );
  AOI22_X1 U5871 ( .A1(n4893), .A2(n6254), .B1(n6437), .B2(n5155), .ZN(n4890)
         );
  NAND3_X1 U5872 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n7014), .A3(n6579), .ZN(n4774) );
  NOR2_X1 U5873 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4774), .ZN(n4887)
         );
  INV_X1 U5874 ( .A(n4887), .ZN(n4712) );
  AND2_X1 U5875 ( .A1(n4711), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5154) );
  OAI21_X1 U5876 ( .B1(n5155), .B2(n6935), .A(n5000), .ZN(n5159) );
  AOI211_X1 U5877 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4712), .A(n5154), .B(
        n5159), .ZN(n4718) );
  AOI21_X1 U5878 ( .B1(n4772), .B2(STATEBS16_REG_SCAN_IN), .A(n6729), .ZN(
        n4776) );
  AND2_X1 U5879 ( .A1(n6012), .A2(n4640), .ZN(n4714) );
  AND2_X1 U5880 ( .A1(n4714), .A2(n4730), .ZN(n4998) );
  AND2_X1 U5881 ( .A1(n4998), .A2(n4964), .ZN(n4719) );
  NAND2_X1 U5882 ( .A1(n4719), .A2(n6444), .ZN(n4715) );
  OAI211_X1 U5883 ( .C1(n4897), .C2(n4716), .A(n4776), .B(n4715), .ZN(n4717)
         );
  NAND2_X1 U5884 ( .A1(n4718), .A2(n4717), .ZN(n4884) );
  NAND2_X1 U5885 ( .A1(n4884), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4722) );
  NAND2_X1 U5886 ( .A1(n4772), .A2(n5379), .ZN(n4885) );
  OAI22_X1 U5887 ( .A1(n4885), .A2(n6454), .B1(n5100), .B2(n6517), .ZN(n4720)
         );
  AOI21_X1 U5888 ( .B1(n6504), .B2(n4887), .A(n4720), .ZN(n4721) );
  OAI211_X1 U5889 ( .C1(n4890), .C2(n5433), .A(n4722), .B(n4721), .ZN(U3052)
         );
  CLKBUF_X1 U5890 ( .A(n4723), .Z(n4725) );
  XNOR2_X1 U5891 ( .A(n4725), .B(n4724), .ZN(n5153) );
  OAI22_X1 U5892 ( .A1(n6342), .A2(n6774), .B1(n6434), .B2(n6641), .ZN(n4727)
         );
  NOR2_X1 U5893 ( .A1(n6242), .A2(n6361), .ZN(n4726) );
  AOI211_X1 U5894 ( .C1(n6336), .C2(n6240), .A(n4727), .B(n4726), .ZN(n4728)
         );
  OAI21_X1 U5895 ( .B1(n6355), .B2(n5153), .A(n4728), .ZN(U2982) );
  NAND3_X1 U5896 ( .A1(n7014), .A2(n6586), .A3(n6579), .ZN(n5158) );
  NOR2_X1 U5897 ( .A1(n4838), .A2(n5158), .ZN(n4729) );
  INV_X1 U5898 ( .A(n4729), .ZN(n4875) );
  NAND2_X1 U5899 ( .A1(n6014), .A2(n6010), .ZN(n4837) );
  NOR2_X1 U5900 ( .A1(n6439), .A2(n4837), .ZN(n5163) );
  AOI21_X1 U5901 ( .B1(n5163), .B2(n6575), .A(n4729), .ZN(n4736) );
  AND2_X1 U5902 ( .A1(n6012), .A2(n4839), .ZN(n4731) );
  NAND2_X1 U5903 ( .A1(n4731), .A2(n4730), .ZN(n4737) );
  OR2_X1 U5904 ( .A1(n4737), .A2(n6121), .ZN(n4732) );
  AOI22_X1 U5905 ( .A1(n4736), .A2(n4734), .B1(n6729), .B2(n5158), .ZN(n4733)
         );
  NAND2_X1 U5906 ( .A1(n4959), .A2(n4733), .ZN(n4872) );
  INV_X1 U5907 ( .A(n4734), .ZN(n4735) );
  OAI22_X1 U5908 ( .A1(n4736), .A2(n4735), .B1(n6935), .B2(n5158), .ZN(n4871)
         );
  AOI22_X1 U5909 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4872), .B1(n6532), 
        .B2(n4871), .ZN(n4739) );
  AOI22_X1 U5910 ( .A1(n6463), .A2(n5164), .B1(n5002), .B2(n6530), .ZN(n4738)
         );
  OAI211_X1 U5911 ( .C1(n5411), .C2(n4875), .A(n4739), .B(n4738), .ZN(U3031)
         );
  AOI22_X1 U5912 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4872), .B1(n6520), 
        .B2(n4871), .ZN(n4741) );
  AOI22_X1 U5913 ( .A1(n6455), .A2(n5164), .B1(n5002), .B2(n6518), .ZN(n4740)
         );
  OAI211_X1 U5914 ( .C1(n5422), .C2(n4875), .A(n4741), .B(n4740), .ZN(U3029)
         );
  AOI22_X1 U5915 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4872), .B1(n6561), 
        .B2(n4871), .ZN(n4743) );
  AOI22_X1 U5916 ( .A1(n6478), .A2(n5164), .B1(n5002), .B2(n6556), .ZN(n4742)
         );
  OAI211_X1 U5917 ( .C1(n5391), .C2(n4875), .A(n4743), .B(n4742), .ZN(U3035)
         );
  AOI22_X1 U5918 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4872), .B1(n6514), 
        .B2(n4871), .ZN(n4745) );
  AOI22_X1 U5919 ( .A1(n6451), .A2(n5164), .B1(n5002), .B2(n6503), .ZN(n4744)
         );
  OAI211_X1 U5920 ( .C1(n5429), .C2(n4875), .A(n4745), .B(n4744), .ZN(U3028)
         );
  NOR2_X2 U5921 ( .A1(n4806), .A2(n3365), .ZN(n6537) );
  INV_X1 U5922 ( .A(n6537), .ZN(n5417) );
  AOI22_X1 U5923 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4877), .B1(n6538), 
        .B2(n4876), .ZN(n4749) );
  INV_X1 U5924 ( .A(DATAI_28_), .ZN(n4746) );
  OR2_X1 U5925 ( .A1(n6361), .A2(n4746), .ZN(n5196) );
  INV_X1 U5926 ( .A(n5196), .ZN(n6536) );
  INV_X1 U5927 ( .A(DATAI_20_), .ZN(n4747) );
  OR2_X1 U5928 ( .A1(n6361), .A2(n4747), .ZN(n6541) );
  INV_X1 U5929 ( .A(n6541), .ZN(n5415) );
  AOI22_X1 U5930 ( .A1(n6536), .A2(n4895), .B1(n5113), .B2(n5415), .ZN(n4748)
         );
  OAI211_X1 U5931 ( .C1(n5417), .C2(n4880), .A(n4749), .B(n4748), .ZN(U3128)
         );
  XNOR2_X1 U5932 ( .A(n4752), .B(n4751), .ZN(n6334) );
  INV_X1 U5933 ( .A(n4753), .ZN(n6402) );
  INV_X1 U5934 ( .A(n5355), .ZN(n6412) );
  AOI21_X1 U5935 ( .B1(n6402), .B2(n4754), .A(n6412), .ZN(n6410) );
  OAI21_X1 U5936 ( .B1(n4760), .B2(n6414), .A(n6410), .ZN(n4831) );
  NAND2_X1 U5937 ( .A1(n4756), .A2(n4755), .ZN(n4757) );
  NAND2_X1 U5938 ( .A1(n5051), .A2(n4757), .ZN(n6215) );
  NOR2_X1 U5939 ( .A1(n6215), .A2(n6424), .ZN(n4763) );
  OR2_X1 U5940 ( .A1(n6399), .A2(n6402), .ZN(n4758) );
  NAND2_X1 U5941 ( .A1(n4758), .A2(n5147), .ZN(n5148) );
  INV_X1 U5942 ( .A(n5148), .ZN(n5225) );
  NAND2_X1 U5943 ( .A1(n4760), .A2(n4759), .ZN(n4761) );
  NAND2_X1 U5944 ( .A1(n3952), .A2(REIP_REG_6__SCAN_IN), .ZN(n6340) );
  OAI21_X1 U5945 ( .B1(n5225), .B2(n4761), .A(n6340), .ZN(n4762) );
  AOI211_X1 U5946 ( .C1(n4831), .C2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n4763), 
        .B(n4762), .ZN(n4764) );
  OAI21_X1 U5947 ( .B1(n6425), .B2(n6334), .A(n4764), .ZN(U3012) );
  AOI22_X1 U5948 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4872), .B1(n6538), 
        .B2(n4871), .ZN(n4766) );
  AOI22_X1 U5949 ( .A1(n6536), .A2(n5164), .B1(n5002), .B2(n5415), .ZN(n4765)
         );
  OAI211_X1 U5950 ( .C1(n5417), .C2(n4875), .A(n4766), .B(n4765), .ZN(U3032)
         );
  AOI22_X1 U5951 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4872), .B1(n6526), 
        .B2(n4871), .ZN(n4768) );
  AOI22_X1 U5952 ( .A1(n6459), .A2(n5164), .B1(n5002), .B2(n6524), .ZN(n4767)
         );
  OAI211_X1 U5953 ( .C1(n5406), .C2(n4875), .A(n4768), .B(n4767), .ZN(U3030)
         );
  INV_X1 U5954 ( .A(n4776), .ZN(n4770) );
  NOR2_X1 U5955 ( .A1(n5297), .A2(n4897), .ZN(n4769) );
  NOR2_X1 U5956 ( .A1(n4838), .A2(n4774), .ZN(n4810) );
  AOI21_X1 U5957 ( .B1(n4898), .B2(n4769), .A(n4810), .ZN(n4775) );
  OAI22_X1 U5958 ( .A1(n4770), .A2(n4775), .B1(n4774), .B2(n6935), .ZN(n4771)
         );
  OAI22_X1 U5959 ( .A1(n5196), .A2(n4885), .B1(n6450), .B2(n6541), .ZN(n4773)
         );
  AOI21_X1 U5960 ( .B1(n6537), .B2(n4810), .A(n4773), .ZN(n4780) );
  INV_X1 U5961 ( .A(n4774), .ZN(n4778) );
  NAND2_X1 U5962 ( .A1(n4776), .A2(n4775), .ZN(n4777) );
  OAI211_X1 U5963 ( .C1(n6442), .C2(n4778), .A(n4777), .B(n4959), .ZN(n4811)
         );
  NAND2_X1 U5964 ( .A1(n4811), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4779) );
  OAI211_X1 U5965 ( .C1(n4814), .C2(n5420), .A(n4780), .B(n4779), .ZN(U3064)
         );
  OAI22_X1 U5966 ( .A1(n6566), .A2(n4885), .B1(n6450), .B2(n6482), .ZN(n4781)
         );
  AOI21_X1 U5967 ( .B1(n6559), .B2(n4810), .A(n4781), .ZN(n4783) );
  NAND2_X1 U5968 ( .A1(n4811), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4782) );
  OAI211_X1 U5969 ( .C1(n4814), .C2(n5394), .A(n4783), .B(n4782), .ZN(U3067)
         );
  OAI22_X1 U5970 ( .A1(n6535), .A2(n4885), .B1(n6450), .B2(n6466), .ZN(n4784)
         );
  AOI21_X1 U5971 ( .B1(n6531), .B2(n4810), .A(n4784), .ZN(n4786) );
  NAND2_X1 U5972 ( .A1(n4811), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4785) );
  OAI211_X1 U5973 ( .C1(n4814), .C2(n5414), .A(n4786), .B(n4785), .ZN(U3063)
         );
  OAI22_X1 U5974 ( .A1(n6517), .A2(n4885), .B1(n6450), .B2(n6454), .ZN(n4787)
         );
  AOI21_X1 U5975 ( .B1(n6504), .B2(n4810), .A(n4787), .ZN(n4789) );
  NAND2_X1 U5976 ( .A1(n4811), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4788) );
  OAI211_X1 U5977 ( .C1(n4814), .C2(n5433), .A(n4789), .B(n4788), .ZN(U3060)
         );
  OAI22_X1 U5978 ( .A1(n6523), .A2(n4885), .B1(n6450), .B2(n6458), .ZN(n4790)
         );
  AOI21_X1 U5979 ( .B1(n6519), .B2(n4810), .A(n4790), .ZN(n4792) );
  NAND2_X1 U5980 ( .A1(n4811), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4791) );
  OAI211_X1 U5981 ( .C1(n4814), .C2(n5425), .A(n4792), .B(n4791), .ZN(U3061)
         );
  OAI22_X1 U5982 ( .A1(n6529), .A2(n4885), .B1(n6450), .B2(n6462), .ZN(n4793)
         );
  AOI21_X1 U5983 ( .B1(n6525), .B2(n4810), .A(n4793), .ZN(n4795) );
  NAND2_X1 U5984 ( .A1(n4811), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4794) );
  OAI211_X1 U5985 ( .C1(n4814), .C2(n5409), .A(n4795), .B(n4794), .ZN(U3062)
         );
  OR2_X1 U5986 ( .A1(n4796), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4798)
         );
  AND2_X1 U5987 ( .A1(n4798), .A2(n4797), .ZN(n5299) );
  INV_X1 U5988 ( .A(n5299), .ZN(n6423) );
  OAI222_X1 U5989 ( .A1(n6423), .A2(n5808), .B1(n5814), .B2(n5293), .C1(n6362), 
        .C2(n5796), .ZN(U2859) );
  NOR2_X2 U5990 ( .A1(n4806), .A2(n4800), .ZN(n6543) );
  INV_X1 U5991 ( .A(DATAI_29_), .ZN(n4801) );
  OR2_X1 U5992 ( .A1(n6361), .A2(n4801), .ZN(n6547) );
  INV_X1 U5993 ( .A(DATAI_21_), .ZN(n6823) );
  OR2_X1 U5994 ( .A1(n6361), .A2(n6823), .ZN(n6472) );
  OAI22_X1 U5995 ( .A1(n6547), .A2(n4885), .B1(n6450), .B2(n6472), .ZN(n4802)
         );
  AOI21_X1 U5996 ( .B1(n6543), .B2(n4810), .A(n4802), .ZN(n4804) );
  NAND2_X1 U5997 ( .A1(n4811), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4803) );
  OAI211_X1 U5998 ( .C1(n4814), .C2(n5399), .A(n4804), .B(n4803), .ZN(U3065)
         );
  NOR2_X2 U5999 ( .A1(n4806), .A2(n4805), .ZN(n6550) );
  INV_X1 U6000 ( .A(DATAI_30_), .ZN(n4807) );
  OR2_X1 U6001 ( .A1(n6361), .A2(n4807), .ZN(n6494) );
  INV_X1 U6002 ( .A(DATAI_22_), .ZN(n4808) );
  OR2_X1 U6003 ( .A1(n6361), .A2(n4808), .ZN(n6555) );
  OAI22_X1 U6004 ( .A1(n6494), .A2(n4885), .B1(n6450), .B2(n6555), .ZN(n4809)
         );
  AOI21_X1 U6005 ( .B1(n6550), .B2(n4810), .A(n4809), .ZN(n4813) );
  NAND2_X1 U6006 ( .A1(n4811), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4812) );
  OAI211_X1 U6007 ( .C1(n4814), .C2(n5404), .A(n4813), .B(n4812), .ZN(U3066)
         );
  NAND2_X1 U6008 ( .A1(n4884), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4817) );
  OAI22_X1 U6009 ( .A1(n5100), .A2(n6566), .B1(n6482), .B2(n4885), .ZN(n4815)
         );
  AOI21_X1 U6010 ( .B1(n6559), .B2(n4887), .A(n4815), .ZN(n4816) );
  OAI211_X1 U6011 ( .C1(n4890), .C2(n5394), .A(n4817), .B(n4816), .ZN(U3059)
         );
  NAND2_X1 U6012 ( .A1(n4884), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4820) );
  OAI22_X1 U6013 ( .A1(n5100), .A2(n6523), .B1(n6458), .B2(n4885), .ZN(n4818)
         );
  AOI21_X1 U6014 ( .B1(n6519), .B2(n4887), .A(n4818), .ZN(n4819) );
  OAI211_X1 U6015 ( .C1(n4890), .C2(n5425), .A(n4820), .B(n4819), .ZN(U3053)
         );
  NAND2_X1 U6016 ( .A1(n4884), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4823) );
  OAI22_X1 U6017 ( .A1(n5100), .A2(n6535), .B1(n6466), .B2(n4885), .ZN(n4821)
         );
  AOI21_X1 U6018 ( .B1(n6531), .B2(n4887), .A(n4821), .ZN(n4822) );
  OAI211_X1 U6019 ( .C1(n4890), .C2(n5414), .A(n4823), .B(n4822), .ZN(U3055)
         );
  NAND2_X1 U6020 ( .A1(n4884), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4826) );
  OAI22_X1 U6021 ( .A1(n5100), .A2(n6529), .B1(n6462), .B2(n4885), .ZN(n4824)
         );
  AOI21_X1 U6022 ( .B1(n6525), .B2(n4887), .A(n4824), .ZN(n4825) );
  OAI211_X1 U6023 ( .C1(n4890), .C2(n5409), .A(n4826), .B(n4825), .ZN(U3054)
         );
  CLKBUF_X1 U6024 ( .A(n4827), .Z(n4829) );
  XOR2_X1 U6025 ( .A(n4829), .B(n4828), .Z(n4861) );
  NOR3_X1 U6026 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6399), .A3(n4830), 
        .ZN(n4835) );
  OAI21_X1 U6027 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4832), .A(n4831), 
        .ZN(n4833) );
  NAND2_X1 U6028 ( .A1(n3952), .A2(REIP_REG_5__SCAN_IN), .ZN(n4862) );
  OAI211_X1 U6029 ( .C1(n6424), .C2(n6225), .A(n4833), .B(n4862), .ZN(n4834)
         );
  AOI211_X1 U6030 ( .C1(n4861), .C2(n6420), .A(n4835), .B(n4834), .ZN(n4836)
         );
  INV_X1 U6031 ( .A(n4836), .ZN(U3013) );
  INV_X1 U6032 ( .A(n4837), .ZN(n5232) );
  NAND3_X1 U6033 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6586), .A3(n6579), .ZN(n5235) );
  NOR2_X1 U6034 ( .A1(n4838), .A2(n5235), .ZN(n5023) );
  AOI21_X1 U6035 ( .B1(n4956), .B2(n5232), .A(n5023), .ZN(n4843) );
  NAND3_X1 U6036 ( .A1(n5381), .A2(n4839), .A3(STATEBS16_REG_SCAN_IN), .ZN(
        n4840) );
  AOI22_X1 U6037 ( .A1(n4843), .A2(n4842), .B1(n6729), .B2(n5235), .ZN(n4841)
         );
  NAND2_X1 U6038 ( .A1(n4959), .A2(n4841), .ZN(n5022) );
  INV_X1 U6039 ( .A(n4842), .ZN(n4844) );
  OAI22_X1 U6040 ( .A1(n4844), .A2(n4843), .B1(n6935), .B2(n5235), .ZN(n5021)
         );
  AOI22_X1 U6041 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5022), .B1(n6532), 
        .B2(n5021), .ZN(n4847) );
  AOI22_X1 U6042 ( .A1(n5431), .A2(n6530), .B1(n6531), .B2(n5023), .ZN(n4846)
         );
  OAI211_X1 U6043 ( .C1(n5272), .C2(n6535), .A(n4847), .B(n4846), .ZN(U3095)
         );
  AOI22_X1 U6044 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5022), .B1(n6514), 
        .B2(n5021), .ZN(n4849) );
  AOI22_X1 U6045 ( .A1(n5431), .A2(n6503), .B1(n6504), .B2(n5023), .ZN(n4848)
         );
  OAI211_X1 U6046 ( .C1(n5272), .C2(n6517), .A(n4849), .B(n4848), .ZN(U3092)
         );
  AOI22_X1 U6047 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5022), .B1(n6561), 
        .B2(n5021), .ZN(n4851) );
  AOI22_X1 U6048 ( .A1(n5431), .A2(n6556), .B1(n6559), .B2(n5023), .ZN(n4850)
         );
  OAI211_X1 U6049 ( .C1(n5272), .C2(n6566), .A(n4851), .B(n4850), .ZN(U3099)
         );
  AOI22_X1 U6050 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5022), .B1(n6520), 
        .B2(n5021), .ZN(n4853) );
  AOI22_X1 U6051 ( .A1(n5431), .A2(n6518), .B1(n6519), .B2(n5023), .ZN(n4852)
         );
  OAI211_X1 U6052 ( .C1(n5272), .C2(n6523), .A(n4853), .B(n4852), .ZN(U3093)
         );
  AOI22_X1 U6053 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5022), .B1(n6526), 
        .B2(n5021), .ZN(n4855) );
  AOI22_X1 U6054 ( .A1(n5431), .A2(n6524), .B1(n6525), .B2(n5023), .ZN(n4854)
         );
  OAI211_X1 U6055 ( .C1(n5272), .C2(n6529), .A(n4855), .B(n4854), .ZN(U3094)
         );
  AOI22_X1 U6056 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5022), .B1(n6538), 
        .B2(n5021), .ZN(n4857) );
  AOI22_X1 U6057 ( .A1(n5431), .A2(n5415), .B1(n6537), .B2(n5023), .ZN(n4856)
         );
  OAI211_X1 U6058 ( .C1(n5272), .C2(n5196), .A(n4857), .B(n4856), .ZN(U3096)
         );
  NAND2_X1 U6059 ( .A1(n4884), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4860) );
  OAI22_X1 U6060 ( .A1(n5100), .A2(n5196), .B1(n6541), .B2(n4885), .ZN(n4858)
         );
  AOI21_X1 U6061 ( .B1(n6537), .B2(n4887), .A(n4858), .ZN(n4859) );
  OAI211_X1 U6062 ( .C1(n4890), .C2(n5420), .A(n4860), .B(n4859), .ZN(U3056)
         );
  NAND2_X1 U6063 ( .A1(n4861), .A2(n4310), .ZN(n4866) );
  INV_X1 U6064 ( .A(n4862), .ZN(n4864) );
  NOR2_X1 U6065 ( .A1(n6352), .A2(n6232), .ZN(n4863) );
  AOI211_X1 U6066 ( .C1(n6358), .C2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4864), 
        .B(n4863), .ZN(n4865) );
  OAI211_X1 U6067 ( .C1(n6361), .C2(n6228), .A(n4866), .B(n4865), .ZN(U2981)
         );
  INV_X1 U6068 ( .A(n6543), .ZN(n5396) );
  AOI22_X1 U6069 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4877), .B1(n6544), 
        .B2(n4876), .ZN(n4868) );
  INV_X1 U6070 ( .A(n6547), .ZN(n6469) );
  INV_X1 U6071 ( .A(n6472), .ZN(n6542) );
  AOI22_X1 U6072 ( .A1(n6469), .A2(n4895), .B1(n5113), .B2(n6542), .ZN(n4867)
         );
  OAI211_X1 U6073 ( .C1(n5396), .C2(n4880), .A(n4868), .B(n4867), .ZN(U3129)
         );
  INV_X1 U6074 ( .A(n6550), .ZN(n5401) );
  AOI22_X1 U6075 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4872), .B1(n6551), 
        .B2(n4871), .ZN(n4870) );
  INV_X1 U6076 ( .A(n6494), .ZN(n6548) );
  INV_X1 U6077 ( .A(n6555), .ZN(n6491) );
  AOI22_X1 U6078 ( .A1(n6548), .A2(n5164), .B1(n5002), .B2(n6491), .ZN(n4869)
         );
  OAI211_X1 U6079 ( .C1(n5401), .C2(n4875), .A(n4870), .B(n4869), .ZN(U3034)
         );
  AOI22_X1 U6080 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4872), .B1(n6544), 
        .B2(n4871), .ZN(n4874) );
  AOI22_X1 U6081 ( .A1(n6469), .A2(n5164), .B1(n5002), .B2(n6542), .ZN(n4873)
         );
  OAI211_X1 U6082 ( .C1(n5396), .C2(n4875), .A(n4874), .B(n4873), .ZN(U3033)
         );
  AOI22_X1 U6083 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4877), .B1(n6551), 
        .B2(n4876), .ZN(n4879) );
  AOI22_X1 U6084 ( .A1(n6548), .A2(n4895), .B1(n5113), .B2(n6491), .ZN(n4878)
         );
  OAI211_X1 U6085 ( .C1(n5401), .C2(n4880), .A(n4879), .B(n4878), .ZN(U3130)
         );
  NAND2_X1 U6086 ( .A1(n4884), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4883) );
  OAI22_X1 U6087 ( .A1(n5100), .A2(n6494), .B1(n6555), .B2(n4885), .ZN(n4881)
         );
  AOI21_X1 U6088 ( .B1(n6550), .B2(n4887), .A(n4881), .ZN(n4882) );
  OAI211_X1 U6089 ( .C1(n4890), .C2(n5404), .A(n4883), .B(n4882), .ZN(U3058)
         );
  NAND2_X1 U6090 ( .A1(n4884), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4889) );
  OAI22_X1 U6091 ( .A1(n5100), .A2(n6547), .B1(n6472), .B2(n4885), .ZN(n4886)
         );
  AOI21_X1 U6092 ( .B1(n6543), .B2(n4887), .A(n4886), .ZN(n4888) );
  OAI211_X1 U6093 ( .C1(n4890), .C2(n5399), .A(n4889), .B(n4888), .ZN(U3057)
         );
  NAND2_X1 U6094 ( .A1(n4891), .A2(n5384), .ZN(n5240) );
  INV_X1 U6095 ( .A(n5240), .ZN(n4892) );
  AOI22_X1 U6096 ( .A1(n4893), .A2(n6439), .B1(n4892), .B2(n6437), .ZN(n4930)
         );
  AND2_X1 U6097 ( .A1(n4640), .A2(n4964), .ZN(n4894) );
  AOI21_X1 U6098 ( .B1(n6554), .B2(n4925), .A(n6121), .ZN(n4896) );
  AOI211_X1 U6099 ( .C1(n4898), .C2(n4897), .A(n6729), .B(n4896), .ZN(n4902)
         );
  NOR2_X1 U6100 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4899), .ZN(n4927)
         );
  INV_X1 U6101 ( .A(n5154), .ZN(n6446) );
  AOI21_X1 U6102 ( .B1(n5240), .B2(STATE2_REG_2__SCAN_IN), .A(n4900), .ZN(
        n5236) );
  OAI211_X1 U6103 ( .C1(n6702), .C2(n4927), .A(n6446), .B(n5236), .ZN(n4901)
         );
  NAND2_X1 U6104 ( .A1(n4924), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4905)
         );
  OAI22_X1 U6105 ( .A1(n6554), .A2(n6529), .B1(n4925), .B2(n6462), .ZN(n4903)
         );
  AOI21_X1 U6106 ( .B1(n6525), .B2(n4927), .A(n4903), .ZN(n4904) );
  OAI211_X1 U6107 ( .C1(n4930), .C2(n5409), .A(n4905), .B(n4904), .ZN(U3118)
         );
  NAND2_X1 U6108 ( .A1(n4924), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4908)
         );
  OAI22_X1 U6109 ( .A1(n6554), .A2(n6517), .B1(n4925), .B2(n6454), .ZN(n4906)
         );
  AOI21_X1 U6110 ( .B1(n6504), .B2(n4927), .A(n4906), .ZN(n4907) );
  OAI211_X1 U6111 ( .C1(n4930), .C2(n5433), .A(n4908), .B(n4907), .ZN(U3116)
         );
  NAND2_X1 U6112 ( .A1(n4924), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4911)
         );
  OAI22_X1 U6113 ( .A1(n6554), .A2(n6535), .B1(n4925), .B2(n6466), .ZN(n4909)
         );
  AOI21_X1 U6114 ( .B1(n6531), .B2(n4927), .A(n4909), .ZN(n4910) );
  OAI211_X1 U6115 ( .C1(n4930), .C2(n5414), .A(n4911), .B(n4910), .ZN(U3119)
         );
  NAND2_X1 U6116 ( .A1(n4924), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4914)
         );
  OAI22_X1 U6117 ( .A1(n6554), .A2(n6494), .B1(n4925), .B2(n6555), .ZN(n4912)
         );
  AOI21_X1 U6118 ( .B1(n6550), .B2(n4927), .A(n4912), .ZN(n4913) );
  OAI211_X1 U6119 ( .C1(n4930), .C2(n5404), .A(n4914), .B(n4913), .ZN(U3122)
         );
  NAND2_X1 U6120 ( .A1(n4924), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4917)
         );
  OAI22_X1 U6121 ( .A1(n6554), .A2(n6566), .B1(n4925), .B2(n6482), .ZN(n4915)
         );
  AOI21_X1 U6122 ( .B1(n6559), .B2(n4927), .A(n4915), .ZN(n4916) );
  OAI211_X1 U6123 ( .C1(n4930), .C2(n5394), .A(n4917), .B(n4916), .ZN(U3123)
         );
  NAND2_X1 U6124 ( .A1(n4924), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4920)
         );
  OAI22_X1 U6125 ( .A1(n6554), .A2(n6547), .B1(n4925), .B2(n6472), .ZN(n4918)
         );
  AOI21_X1 U6126 ( .B1(n6543), .B2(n4927), .A(n4918), .ZN(n4919) );
  OAI211_X1 U6127 ( .C1(n4930), .C2(n5399), .A(n4920), .B(n4919), .ZN(U3121)
         );
  NAND2_X1 U6128 ( .A1(n4924), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4923)
         );
  OAI22_X1 U6129 ( .A1(n6554), .A2(n6523), .B1(n4925), .B2(n6458), .ZN(n4921)
         );
  AOI21_X1 U6130 ( .B1(n6519), .B2(n4927), .A(n4921), .ZN(n4922) );
  OAI211_X1 U6131 ( .C1(n4930), .C2(n5425), .A(n4923), .B(n4922), .ZN(U3117)
         );
  NAND2_X1 U6132 ( .A1(n4924), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4929)
         );
  OAI22_X1 U6133 ( .A1(n6554), .A2(n5196), .B1(n4925), .B2(n6541), .ZN(n4926)
         );
  AOI21_X1 U6134 ( .B1(n6537), .B2(n4927), .A(n4926), .ZN(n4928) );
  OAI211_X1 U6135 ( .C1(n4930), .C2(n5420), .A(n4929), .B(n4928), .ZN(U3120)
         );
  OR2_X1 U6136 ( .A1(n4932), .A2(n4931), .ZN(n4933) );
  AND2_X1 U6137 ( .A1(n4934), .A2(n4933), .ZN(n6417) );
  INV_X1 U6138 ( .A(n6417), .ZN(n4935) );
  INV_X1 U6139 ( .A(n5814), .ZN(n5805) );
  AOI22_X1 U6140 ( .A1(n5811), .A2(n4935), .B1(n5805), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4936) );
  OAI21_X1 U6141 ( .B1(n5760), .B2(n5796), .A(n4936), .ZN(U2858) );
  OAI21_X1 U6142 ( .B1(n4942), .B2(n4937), .A(n4706), .ZN(n6237) );
  INV_X1 U6143 ( .A(n6237), .ZN(n4938) );
  AOI22_X1 U6144 ( .A1(n5811), .A2(n4938), .B1(n5805), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4939) );
  OAI21_X1 U6145 ( .B1(n6242), .B2(n5796), .A(n4939), .ZN(U2855) );
  AND2_X1 U6146 ( .A1(n4947), .A2(n4940), .ZN(n4941) );
  NOR2_X1 U6147 ( .A1(n4942), .A2(n4941), .ZN(n6391) );
  AOI22_X1 U6148 ( .A1(n5811), .A2(n6391), .B1(n5805), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4943) );
  OAI21_X1 U6149 ( .B1(n6261), .B2(n5796), .A(n4943), .ZN(U2856) );
  NAND2_X1 U6150 ( .A1(n4945), .A2(n4944), .ZN(n4946) );
  NAND2_X1 U6151 ( .A1(n4947), .A2(n4946), .ZN(n6406) );
  INV_X1 U6152 ( .A(n6406), .ZN(n4948) );
  AOI22_X1 U6153 ( .A1(n5811), .A2(n4948), .B1(n5805), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4949) );
  OAI21_X1 U6154 ( .B1(n6346), .B2(n5796), .A(n4949), .ZN(U2857) );
  CLKBUF_X1 U6155 ( .A(n4950), .Z(n4951) );
  AOI21_X1 U6156 ( .B1(n4952), .B2(n4583), .A(n4951), .ZN(n6338) );
  INV_X1 U6157 ( .A(n6338), .ZN(n5040) );
  INV_X1 U6158 ( .A(n6215), .ZN(n4953) );
  AOI22_X1 U6159 ( .A1(n4953), .A2(n5811), .B1(n5805), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4954) );
  OAI21_X1 U6160 ( .B1(n5040), .B2(n5796), .A(n4954), .ZN(U2853) );
  INV_X1 U6161 ( .A(n4955), .ZN(n5059) );
  AOI21_X1 U6162 ( .B1(n4956), .B2(n5112), .A(n5059), .ZN(n4962) );
  OAI22_X1 U6163 ( .A1(n4962), .A2(n6729), .B1(n5110), .B2(n6935), .ZN(n5064)
         );
  NAND2_X1 U6164 ( .A1(n3490), .A2(n4640), .ZN(n4957) );
  NAND2_X1 U6165 ( .A1(n4965), .A2(n6347), .ZN(n4958) );
  NAND2_X1 U6166 ( .A1(n4958), .A2(n6444), .ZN(n4963) );
  OAI21_X1 U6167 ( .B1(n6442), .B2(n4960), .A(n4959), .ZN(n4961) );
  AOI21_X1 U6168 ( .B1(n4963), .B2(n4962), .A(n4961), .ZN(n5062) );
  INV_X1 U6169 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4968) );
  NAND2_X1 U6170 ( .A1(n6519), .A2(n5059), .ZN(n4967) );
  AOI22_X1 U6171 ( .A1(n6455), .A2(n5114), .B1(n5165), .B2(n6518), .ZN(n4966)
         );
  OAI211_X1 U6172 ( .C1(n5062), .C2(n4968), .A(n4967), .B(n4966), .ZN(n4969)
         );
  AOI21_X1 U6173 ( .B1(n6520), .B2(n5064), .A(n4969), .ZN(n4970) );
  INV_X1 U6174 ( .A(n4970), .ZN(U3141) );
  INV_X1 U6175 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4973) );
  NAND2_X1 U6176 ( .A1(n6525), .A2(n5059), .ZN(n4972) );
  AOI22_X1 U6177 ( .A1(n6459), .A2(n5114), .B1(n5165), .B2(n6524), .ZN(n4971)
         );
  OAI211_X1 U6178 ( .C1(n5062), .C2(n4973), .A(n4972), .B(n4971), .ZN(n4974)
         );
  AOI21_X1 U6179 ( .B1(n6526), .B2(n5064), .A(n4974), .ZN(n4975) );
  INV_X1 U6180 ( .A(n4975), .ZN(U3142) );
  INV_X1 U6181 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4978) );
  NAND2_X1 U6182 ( .A1(n6504), .A2(n5059), .ZN(n4977) );
  AOI22_X1 U6183 ( .A1(n6451), .A2(n5114), .B1(n5165), .B2(n6503), .ZN(n4976)
         );
  OAI211_X1 U6184 ( .C1(n5062), .C2(n4978), .A(n4977), .B(n4976), .ZN(n4979)
         );
  AOI21_X1 U6185 ( .B1(n6514), .B2(n5064), .A(n4979), .ZN(n4980) );
  INV_X1 U6186 ( .A(n4980), .ZN(U3140) );
  INV_X1 U6187 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4983) );
  NAND2_X1 U6188 ( .A1(n6559), .A2(n5059), .ZN(n4982) );
  AOI22_X1 U6189 ( .A1(n6478), .A2(n5114), .B1(n5165), .B2(n6556), .ZN(n4981)
         );
  OAI211_X1 U6190 ( .C1(n5062), .C2(n4983), .A(n4982), .B(n4981), .ZN(n4984)
         );
  AOI21_X1 U6191 ( .B1(n6561), .B2(n5064), .A(n4984), .ZN(n4985) );
  INV_X1 U6192 ( .A(n4985), .ZN(U3147) );
  INV_X1 U6193 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4988) );
  NAND2_X1 U6194 ( .A1(n6537), .A2(n5059), .ZN(n4987) );
  AOI22_X1 U6195 ( .A1(n6536), .A2(n5114), .B1(n5165), .B2(n5415), .ZN(n4986)
         );
  OAI211_X1 U6196 ( .C1(n5062), .C2(n4988), .A(n4987), .B(n4986), .ZN(n4989)
         );
  AOI21_X1 U6197 ( .B1(n6538), .B2(n5064), .A(n4989), .ZN(n4990) );
  INV_X1 U6198 ( .A(n4990), .ZN(U3144) );
  INV_X1 U6199 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4993) );
  NAND2_X1 U6200 ( .A1(n6531), .A2(n5059), .ZN(n4992) );
  AOI22_X1 U6201 ( .A1(n6463), .A2(n5114), .B1(n5165), .B2(n6530), .ZN(n4991)
         );
  OAI211_X1 U6202 ( .C1(n5062), .C2(n4993), .A(n4992), .B(n4991), .ZN(n4994)
         );
  AOI21_X1 U6203 ( .B1(n6532), .B2(n5064), .A(n4994), .ZN(n4995) );
  INV_X1 U6204 ( .A(n4995), .ZN(U3143) );
  AND2_X1 U6205 ( .A1(n6014), .A2(n5763), .ZN(n5383) );
  NAND2_X1 U6206 ( .A1(n6254), .A2(n5383), .ZN(n5069) );
  INV_X1 U6207 ( .A(n5069), .ZN(n4997) );
  NOR3_X1 U6208 ( .A1(n6446), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n5384), 
        .ZN(n4996) );
  AOI21_X1 U6209 ( .B1(n4997), .B2(n6442), .A(n4996), .ZN(n5038) );
  AND2_X1 U6210 ( .A1(n4998), .A2(n5379), .ZN(n5003) );
  OAI21_X1 U6211 ( .B1(n5002), .B2(n5003), .A(n6444), .ZN(n4999) );
  AOI21_X1 U6212 ( .B1(n4999), .B2(n5069), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n5001) );
  NAND3_X1 U6213 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n7014), .A3(n6586), .ZN(n5076) );
  NOR2_X1 U6214 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5076), .ZN(n5035)
         );
  OAI21_X1 U6215 ( .B1(n6436), .B2(n6935), .A(n5000), .ZN(n6449) );
  NOR2_X1 U6216 ( .A1(n6437), .A2(n6449), .ZN(n5389) );
  NAND2_X1 U6217 ( .A1(n5032), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5006) );
  OAI22_X1 U6218 ( .A1(n6523), .A2(n5033), .B1(n5101), .B2(n6458), .ZN(n5004)
         );
  AOI21_X1 U6219 ( .B1(n6519), .B2(n5035), .A(n5004), .ZN(n5005) );
  OAI211_X1 U6220 ( .C1(n5038), .C2(n5425), .A(n5006), .B(n5005), .ZN(U3037)
         );
  NAND2_X1 U6221 ( .A1(n5032), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5009) );
  OAI22_X1 U6222 ( .A1(n6566), .A2(n5033), .B1(n5101), .B2(n6482), .ZN(n5007)
         );
  AOI21_X1 U6223 ( .B1(n6559), .B2(n5035), .A(n5007), .ZN(n5008) );
  OAI211_X1 U6224 ( .C1(n5038), .C2(n5394), .A(n5009), .B(n5008), .ZN(U3043)
         );
  NAND2_X1 U6225 ( .A1(n5032), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5012) );
  OAI22_X1 U6226 ( .A1(n6529), .A2(n5033), .B1(n5101), .B2(n6462), .ZN(n5010)
         );
  AOI21_X1 U6227 ( .B1(n6525), .B2(n5035), .A(n5010), .ZN(n5011) );
  OAI211_X1 U6228 ( .C1(n5038), .C2(n5409), .A(n5012), .B(n5011), .ZN(U3038)
         );
  NAND2_X1 U6229 ( .A1(n5032), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5015) );
  OAI22_X1 U6230 ( .A1(n5033), .A2(n6517), .B1(n6454), .B2(n5101), .ZN(n5013)
         );
  AOI21_X1 U6231 ( .B1(n6504), .B2(n5035), .A(n5013), .ZN(n5014) );
  OAI211_X1 U6232 ( .C1(n5038), .C2(n5433), .A(n5015), .B(n5014), .ZN(U3036)
         );
  NAND2_X1 U6233 ( .A1(n5032), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5018) );
  OAI22_X1 U6234 ( .A1(n6535), .A2(n5033), .B1(n5101), .B2(n6466), .ZN(n5016)
         );
  AOI21_X1 U6235 ( .B1(n6531), .B2(n5035), .A(n5016), .ZN(n5017) );
  OAI211_X1 U6236 ( .C1(n5038), .C2(n5414), .A(n5018), .B(n5017), .ZN(U3039)
         );
  AOI22_X1 U6237 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5022), .B1(n6544), 
        .B2(n5021), .ZN(n5020) );
  AOI22_X1 U6238 ( .A1(n5431), .A2(n6542), .B1(n6543), .B2(n5023), .ZN(n5019)
         );
  OAI211_X1 U6239 ( .C1(n5272), .C2(n6547), .A(n5020), .B(n5019), .ZN(U3097)
         );
  AOI22_X1 U6240 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5022), .B1(n6551), 
        .B2(n5021), .ZN(n5025) );
  AOI22_X1 U6241 ( .A1(n5431), .A2(n6491), .B1(n6550), .B2(n5023), .ZN(n5024)
         );
  OAI211_X1 U6242 ( .C1(n5272), .C2(n6494), .A(n5025), .B(n5024), .ZN(U3098)
         );
  NAND2_X1 U6243 ( .A1(n5032), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5028) );
  OAI22_X1 U6244 ( .A1(n5196), .A2(n5033), .B1(n5101), .B2(n6541), .ZN(n5026)
         );
  AOI21_X1 U6245 ( .B1(n6537), .B2(n5035), .A(n5026), .ZN(n5027) );
  OAI211_X1 U6246 ( .C1(n5038), .C2(n5420), .A(n5028), .B(n5027), .ZN(U3040)
         );
  NAND2_X1 U6247 ( .A1(n5032), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5031) );
  OAI22_X1 U6248 ( .A1(n6494), .A2(n5033), .B1(n5101), .B2(n6555), .ZN(n5029)
         );
  AOI21_X1 U6249 ( .B1(n6550), .B2(n5035), .A(n5029), .ZN(n5030) );
  OAI211_X1 U6250 ( .C1(n5038), .C2(n5404), .A(n5031), .B(n5030), .ZN(U3042)
         );
  NAND2_X1 U6251 ( .A1(n5032), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5037) );
  OAI22_X1 U6252 ( .A1(n6547), .A2(n5033), .B1(n5101), .B2(n6472), .ZN(n5034)
         );
  AOI21_X1 U6253 ( .B1(n6543), .B2(n5035), .A(n5034), .ZN(n5036) );
  OAI211_X1 U6254 ( .C1(n5038), .C2(n5399), .A(n5037), .B(n5036), .ZN(U3041)
         );
  INV_X1 U6255 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6295) );
  OAI222_X1 U6256 ( .A1(n5040), .A2(n5834), .B1(n5481), .B2(n5039), .C1(n5816), 
        .C2(n6295), .ZN(U2885) );
  OAI22_X1 U6257 ( .A1(n5233), .A2(n6541), .B1(n5196), .B2(n6501), .ZN(n5043)
         );
  NOR2_X1 U6258 ( .A1(n5417), .A2(n5041), .ZN(n5042) );
  AOI211_X1 U6259 ( .C1(INSTQUEUE_REG_7__4__SCAN_IN), .C2(n6498), .A(n5043), 
        .B(n5042), .ZN(n5044) );
  OAI21_X1 U6260 ( .B1(n5045), .B2(n5420), .A(n5044), .ZN(U3080) );
  CLKBUF_X1 U6261 ( .A(n5047), .Z(n5048) );
  OAI21_X1 U6262 ( .B1(n4951), .B2(n5046), .A(n5048), .ZN(n6203) );
  OAI222_X1 U6263 ( .A1(n6203), .A2(n5834), .B1(n5481), .B2(n5049), .C1(n5816), 
        .C2(n3569), .ZN(U2884) );
  INV_X1 U6264 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5053) );
  AND2_X1 U6265 ( .A1(n5051), .A2(n5050), .ZN(n5052) );
  NOR2_X1 U6266 ( .A1(n5222), .A2(n5052), .ZN(n6380) );
  INV_X1 U6267 ( .A(n6380), .ZN(n6209) );
  OAI222_X1 U6268 ( .A1(n6203), .A2(n5796), .B1(n5814), .B2(n5053), .C1(n6209), 
        .C2(n5808), .ZN(U2852) );
  INV_X1 U6269 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5056) );
  NAND2_X1 U6270 ( .A1(n6543), .A2(n5059), .ZN(n5055) );
  AOI22_X1 U6271 ( .A1(n6469), .A2(n5114), .B1(n5165), .B2(n6542), .ZN(n5054)
         );
  OAI211_X1 U6272 ( .C1(n5062), .C2(n5056), .A(n5055), .B(n5054), .ZN(n5057)
         );
  AOI21_X1 U6273 ( .B1(n6544), .B2(n5064), .A(n5057), .ZN(n5058) );
  INV_X1 U6274 ( .A(n5058), .ZN(U3145) );
  NAND2_X1 U6275 ( .A1(n6550), .A2(n5059), .ZN(n5061) );
  AOI22_X1 U6276 ( .A1(n6548), .A2(n5114), .B1(n5165), .B2(n6491), .ZN(n5060)
         );
  OAI211_X1 U6277 ( .C1(n5062), .C2(n6806), .A(n5061), .B(n5060), .ZN(n5063)
         );
  AOI21_X1 U6278 ( .B1(n6551), .B2(n5064), .A(n5063), .ZN(n5065) );
  INV_X1 U6279 ( .A(n5065), .ZN(U3146) );
  NOR3_X1 U6280 ( .A1(n5067), .A2(n5066), .A3(n6505), .ZN(n5068) );
  NOR2_X1 U6281 ( .A1(n5068), .A2(n6729), .ZN(n5075) );
  OR2_X1 U6282 ( .A1(n5069), .A2(n5297), .ZN(n5071) );
  INV_X1 U6283 ( .A(n6502), .ZN(n5070) );
  NAND2_X1 U6284 ( .A1(n5070), .A2(n7014), .ZN(n5073) );
  NAND2_X1 U6285 ( .A1(n5071), .A2(n5073), .ZN(n5078) );
  INV_X1 U6286 ( .A(n5076), .ZN(n5072) );
  AOI22_X1 U6287 ( .A1(n5075), .A2(n5078), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5072), .ZN(n5107) );
  INV_X1 U6288 ( .A(n5073), .ZN(n5103) );
  OAI22_X1 U6289 ( .A1(n6566), .A2(n5101), .B1(n5100), .B2(n6482), .ZN(n5074)
         );
  AOI21_X1 U6290 ( .B1(n6559), .B2(n5103), .A(n5074), .ZN(n5081) );
  INV_X1 U6291 ( .A(n5075), .ZN(n5079) );
  AOI21_X1 U6292 ( .B1(n6729), .B2(n5076), .A(n6508), .ZN(n5077) );
  NAND2_X1 U6293 ( .A1(n5104), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5080) );
  OAI211_X1 U6294 ( .C1(n5107), .C2(n5394), .A(n5081), .B(n5080), .ZN(U3051)
         );
  OAI22_X1 U6295 ( .A1(n6494), .A2(n5101), .B1(n5100), .B2(n6555), .ZN(n5082)
         );
  AOI21_X1 U6296 ( .B1(n6550), .B2(n5103), .A(n5082), .ZN(n5084) );
  NAND2_X1 U6297 ( .A1(n5104), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5083) );
  OAI211_X1 U6298 ( .C1(n5107), .C2(n5404), .A(n5084), .B(n5083), .ZN(U3050)
         );
  OAI22_X1 U6299 ( .A1(n6523), .A2(n5101), .B1(n5100), .B2(n6458), .ZN(n5085)
         );
  AOI21_X1 U6300 ( .B1(n6519), .B2(n5103), .A(n5085), .ZN(n5087) );
  NAND2_X1 U6301 ( .A1(n5104), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n5086) );
  OAI211_X1 U6302 ( .C1(n5107), .C2(n5425), .A(n5087), .B(n5086), .ZN(U3045)
         );
  OAI22_X1 U6303 ( .A1(n6547), .A2(n5101), .B1(n5100), .B2(n6472), .ZN(n5088)
         );
  AOI21_X1 U6304 ( .B1(n6543), .B2(n5103), .A(n5088), .ZN(n5090) );
  NAND2_X1 U6305 ( .A1(n5104), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5089) );
  OAI211_X1 U6306 ( .C1(n5107), .C2(n5399), .A(n5090), .B(n5089), .ZN(U3049)
         );
  OAI22_X1 U6307 ( .A1(n5196), .A2(n5101), .B1(n5100), .B2(n6541), .ZN(n5091)
         );
  AOI21_X1 U6308 ( .B1(n6537), .B2(n5103), .A(n5091), .ZN(n5093) );
  NAND2_X1 U6309 ( .A1(n5104), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5092) );
  OAI211_X1 U6310 ( .C1(n5107), .C2(n5420), .A(n5093), .B(n5092), .ZN(U3048)
         );
  OAI22_X1 U6311 ( .A1(n6535), .A2(n5101), .B1(n5100), .B2(n6466), .ZN(n5094)
         );
  AOI21_X1 U6312 ( .B1(n6531), .B2(n5103), .A(n5094), .ZN(n5096) );
  NAND2_X1 U6313 ( .A1(n5104), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5095) );
  OAI211_X1 U6314 ( .C1(n5107), .C2(n5414), .A(n5096), .B(n5095), .ZN(U3047)
         );
  OAI22_X1 U6315 ( .A1(n6529), .A2(n5101), .B1(n5100), .B2(n6462), .ZN(n5097)
         );
  AOI21_X1 U6316 ( .B1(n6525), .B2(n5103), .A(n5097), .ZN(n5099) );
  NAND2_X1 U6317 ( .A1(n5104), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n5098) );
  OAI211_X1 U6318 ( .C1(n5107), .C2(n5409), .A(n5099), .B(n5098), .ZN(U3046)
         );
  OAI22_X1 U6319 ( .A1(n6517), .A2(n5101), .B1(n5100), .B2(n6454), .ZN(n5102)
         );
  AOI21_X1 U6320 ( .B1(n6504), .B2(n5103), .A(n5102), .ZN(n5106) );
  NAND2_X1 U6321 ( .A1(n5104), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n5105) );
  OAI211_X1 U6322 ( .C1(n5107), .C2(n5433), .A(n5106), .B(n5105), .ZN(U3044)
         );
  NAND2_X1 U6323 ( .A1(n5112), .A2(n6442), .ZN(n6440) );
  INV_X1 U6324 ( .A(n6440), .ZN(n5109) );
  INV_X1 U6325 ( .A(n6437), .ZN(n5237) );
  NOR3_X1 U6326 ( .A1(n5237), .A2(n7014), .A3(n5384), .ZN(n5108) );
  AOI21_X1 U6327 ( .B1(n5109), .B2(n6439), .A(n5108), .ZN(n5146) );
  NOR2_X1 U6328 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5110), .ZN(n5142)
         );
  OAI22_X1 U6329 ( .A1(n6466), .A2(n5140), .B1(n5139), .B2(n6535), .ZN(n5111)
         );
  AOI21_X1 U6330 ( .B1(n6531), .B2(n5142), .A(n5111), .ZN(n5120) );
  INV_X1 U6331 ( .A(n5112), .ZN(n5116) );
  OAI21_X1 U6332 ( .B1(n5114), .B2(n5113), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5115) );
  NAND3_X1 U6333 ( .A1(n5116), .A2(n6442), .A3(n5115), .ZN(n5118) );
  NOR3_X1 U6334 ( .A1(n6449), .A2(n7014), .A3(n5154), .ZN(n5117) );
  NAND2_X1 U6335 ( .A1(n5143), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5119)
         );
  OAI211_X1 U6336 ( .C1(n5414), .C2(n5146), .A(n5120), .B(n5119), .ZN(U3135)
         );
  OAI22_X1 U6337 ( .A1(n6541), .A2(n5140), .B1(n5139), .B2(n5196), .ZN(n5121)
         );
  AOI21_X1 U6338 ( .B1(n6537), .B2(n5142), .A(n5121), .ZN(n5123) );
  NAND2_X1 U6339 ( .A1(n5143), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5122)
         );
  OAI211_X1 U6340 ( .C1(n5420), .C2(n5146), .A(n5123), .B(n5122), .ZN(U3136)
         );
  OAI22_X1 U6341 ( .A1(n5139), .A2(n6517), .B1(n6454), .B2(n5140), .ZN(n5124)
         );
  AOI21_X1 U6342 ( .B1(n6504), .B2(n5142), .A(n5124), .ZN(n5126) );
  NAND2_X1 U6343 ( .A1(n5143), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5125)
         );
  OAI211_X1 U6344 ( .C1(n5433), .C2(n5146), .A(n5126), .B(n5125), .ZN(U3132)
         );
  OAI22_X1 U6345 ( .A1(n6458), .A2(n5140), .B1(n5139), .B2(n6523), .ZN(n5127)
         );
  AOI21_X1 U6346 ( .B1(n6519), .B2(n5142), .A(n5127), .ZN(n5129) );
  NAND2_X1 U6347 ( .A1(n5143), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5128)
         );
  OAI211_X1 U6348 ( .C1(n5425), .C2(n5146), .A(n5129), .B(n5128), .ZN(U3133)
         );
  OAI22_X1 U6349 ( .A1(n6462), .A2(n5140), .B1(n5139), .B2(n6529), .ZN(n5130)
         );
  AOI21_X1 U6350 ( .B1(n6525), .B2(n5142), .A(n5130), .ZN(n5132) );
  NAND2_X1 U6351 ( .A1(n5143), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5131)
         );
  OAI211_X1 U6352 ( .C1(n5409), .C2(n5146), .A(n5132), .B(n5131), .ZN(U3134)
         );
  OAI22_X1 U6353 ( .A1(n6482), .A2(n5140), .B1(n5139), .B2(n6566), .ZN(n5133)
         );
  AOI21_X1 U6354 ( .B1(n6559), .B2(n5142), .A(n5133), .ZN(n5135) );
  NAND2_X1 U6355 ( .A1(n5143), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5134)
         );
  OAI211_X1 U6356 ( .C1(n5394), .C2(n5146), .A(n5135), .B(n5134), .ZN(U3139)
         );
  OAI22_X1 U6357 ( .A1(n6555), .A2(n5140), .B1(n5139), .B2(n6494), .ZN(n5136)
         );
  AOI21_X1 U6358 ( .B1(n6550), .B2(n5142), .A(n5136), .ZN(n5138) );
  NAND2_X1 U6359 ( .A1(n5143), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5137)
         );
  OAI211_X1 U6360 ( .C1(n5404), .C2(n5146), .A(n5138), .B(n5137), .ZN(U3138)
         );
  OAI22_X1 U6361 ( .A1(n6472), .A2(n5140), .B1(n5139), .B2(n6547), .ZN(n5141)
         );
  AOI21_X1 U6362 ( .B1(n6543), .B2(n5142), .A(n5141), .ZN(n5145) );
  NAND2_X1 U6363 ( .A1(n5143), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5144)
         );
  OAI211_X1 U6364 ( .C1(n5399), .C2(n5146), .A(n5145), .B(n5144), .ZN(U3137)
         );
  OAI21_X1 U6365 ( .B1(n5147), .B2(n6401), .A(n6410), .ZN(n6389) );
  NAND2_X1 U6366 ( .A1(n5148), .A2(n6401), .ZN(n6394) );
  AOI221_X1 U6367 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n7003), .C2(n6749), .A(n6394), 
        .ZN(n5149) );
  AOI21_X1 U6368 ( .B1(n3952), .B2(REIP_REG_4__SCAN_IN), .A(n5149), .ZN(n5150)
         );
  OAI21_X1 U6369 ( .B1(n6237), .B2(n6424), .A(n5150), .ZN(n5151) );
  AOI21_X1 U6370 ( .B1(n6389), .B2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n5151), 
        .ZN(n5152) );
  OAI21_X1 U6371 ( .B1(n6425), .B2(n5153), .A(n5152), .ZN(U3014) );
  AOI22_X1 U6372 ( .A1(n5163), .A2(n6442), .B1(n5155), .B2(n5154), .ZN(n5217)
         );
  NOR3_X1 U6373 ( .A1(n5164), .A2(n5165), .A3(n6729), .ZN(n5157) );
  INV_X1 U6374 ( .A(n6444), .ZN(n5156) );
  NOR2_X1 U6375 ( .A1(n5157), .A2(n5156), .ZN(n5162) );
  NOR2_X1 U6376 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5158), .ZN(n5214)
         );
  INV_X1 U6377 ( .A(n5214), .ZN(n5160) );
  AOI211_X1 U6378 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5160), .A(n6437), .B(
        n5159), .ZN(n5161) );
  NAND2_X1 U6379 ( .A1(n5210), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5168) );
  OAI22_X1 U6380 ( .A1(n5212), .A2(n6462), .B1(n6529), .B2(n5211), .ZN(n5166)
         );
  AOI21_X1 U6381 ( .B1(n6525), .B2(n5214), .A(n5166), .ZN(n5167) );
  OAI211_X1 U6382 ( .C1(n5217), .C2(n5409), .A(n5168), .B(n5167), .ZN(U3022)
         );
  NAND2_X1 U6383 ( .A1(n5210), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5171) );
  OAI22_X1 U6384 ( .A1(n5212), .A2(n6458), .B1(n6523), .B2(n5211), .ZN(n5169)
         );
  AOI21_X1 U6385 ( .B1(n6519), .B2(n5214), .A(n5169), .ZN(n5170) );
  OAI211_X1 U6386 ( .C1(n5217), .C2(n5425), .A(n5171), .B(n5170), .ZN(U3021)
         );
  NAND2_X1 U6387 ( .A1(n5210), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5174) );
  OAI22_X1 U6388 ( .A1(n5212), .A2(n6454), .B1(n6517), .B2(n5211), .ZN(n5172)
         );
  AOI21_X1 U6389 ( .B1(n6504), .B2(n5214), .A(n5172), .ZN(n5173) );
  OAI211_X1 U6390 ( .C1(n5217), .C2(n5433), .A(n5174), .B(n5173), .ZN(U3020)
         );
  NAND2_X1 U6391 ( .A1(n5210), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5177) );
  OAI22_X1 U6392 ( .A1(n5212), .A2(n6466), .B1(n6535), .B2(n5211), .ZN(n5175)
         );
  AOI21_X1 U6393 ( .B1(n6531), .B2(n5214), .A(n5175), .ZN(n5176) );
  OAI211_X1 U6394 ( .C1(n5217), .C2(n5414), .A(n5177), .B(n5176), .ZN(U3023)
         );
  NAND2_X1 U6395 ( .A1(n5210), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5180) );
  OAI22_X1 U6396 ( .A1(n5212), .A2(n6482), .B1(n6566), .B2(n5211), .ZN(n5178)
         );
  AOI21_X1 U6397 ( .B1(n6559), .B2(n5214), .A(n5178), .ZN(n5179) );
  OAI211_X1 U6398 ( .C1(n5217), .C2(n5394), .A(n5180), .B(n5179), .ZN(U3027)
         );
  NAND2_X1 U6399 ( .A1(n5182), .A2(n5181), .ZN(n5183) );
  NAND2_X1 U6400 ( .A1(n5312), .A2(n5183), .ZN(n5321) );
  AOI22_X1 U6401 ( .A1(n6742), .A2(DATAI_9_), .B1(n6743), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n5184) );
  OAI21_X1 U6402 ( .B1(n5321), .B2(n5834), .A(n5184), .ZN(U2882) );
  INV_X1 U6403 ( .A(n5317), .ZN(n5194) );
  INV_X1 U6404 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5186) );
  OAI21_X1 U6405 ( .B1(n5224), .B2(n3167), .A(n5344), .ZN(n5279) );
  INV_X1 U6406 ( .A(n5279), .ZN(n6372) );
  AOI22_X1 U6407 ( .A1(n6155), .A2(n6372), .B1(EBX_REG_9__SCAN_IN), .B2(n6264), 
        .ZN(n5185) );
  OAI211_X1 U6408 ( .C1(n6253), .C2(n5186), .A(n5185), .B(n6434), .ZN(n5193)
         );
  INV_X1 U6409 ( .A(n5191), .ZN(n5189) );
  INV_X1 U6410 ( .A(n5187), .ZN(n5190) );
  AND2_X1 U6411 ( .A1(n5754), .A2(n5190), .ZN(n6204) );
  INV_X1 U6412 ( .A(n6204), .ZN(n5188) );
  NOR2_X1 U6413 ( .A1(n6246), .A2(n6236), .ZN(n6205) );
  INV_X1 U6414 ( .A(n6205), .ZN(n6235) );
  OAI21_X1 U6415 ( .B1(n5189), .B2(n5188), .A(n6235), .ZN(n6200) );
  INV_X1 U6416 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6651) );
  AND2_X1 U6417 ( .A1(n6246), .A2(n5190), .ZN(n6206) );
  NAND3_X1 U6418 ( .A1(n5191), .A2(n6206), .A3(n6651), .ZN(n6183) );
  OAI21_X1 U6419 ( .B1(n6200), .B2(n6651), .A(n6183), .ZN(n5192) );
  AOI211_X1 U6420 ( .C1(n6196), .C2(n5194), .A(n5193), .B(n5192), .ZN(n5195)
         );
  OAI21_X1 U6421 ( .B1(n6171), .B2(n5321), .A(n5195), .ZN(U2818) );
  NAND2_X1 U6422 ( .A1(n5210), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5199) );
  OAI22_X1 U6423 ( .A1(n5212), .A2(n6541), .B1(n5196), .B2(n5211), .ZN(n5197)
         );
  AOI21_X1 U6424 ( .B1(n6537), .B2(n5214), .A(n5197), .ZN(n5198) );
  OAI211_X1 U6425 ( .C1(n5217), .C2(n5420), .A(n5199), .B(n5198), .ZN(U3024)
         );
  CLKBUF_X1 U6426 ( .A(n5200), .Z(n5203) );
  INV_X1 U6427 ( .A(n5201), .ZN(n5202) );
  XNOR2_X1 U6428 ( .A(n5203), .B(n5202), .ZN(n6381) );
  NAND2_X1 U6429 ( .A1(n6381), .A2(n4310), .ZN(n5206) );
  NOR2_X1 U6430 ( .A1(n6434), .A2(n6647), .ZN(n6379) );
  NOR2_X1 U6431 ( .A1(n6352), .A2(n6214), .ZN(n5204) );
  AOI211_X1 U6432 ( .C1(n6358), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6379), 
        .B(n5204), .ZN(n5205) );
  OAI211_X1 U6433 ( .C1(n6361), .C2(n6203), .A(n5206), .B(n5205), .ZN(U2979)
         );
  NAND2_X1 U6434 ( .A1(n5210), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5209) );
  OAI22_X1 U6435 ( .A1(n5212), .A2(n6555), .B1(n6494), .B2(n5211), .ZN(n5207)
         );
  AOI21_X1 U6436 ( .B1(n6550), .B2(n5214), .A(n5207), .ZN(n5208) );
  OAI211_X1 U6437 ( .C1(n5217), .C2(n5404), .A(n5209), .B(n5208), .ZN(U3026)
         );
  NAND2_X1 U6438 ( .A1(n5210), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5216) );
  OAI22_X1 U6439 ( .A1(n5212), .A2(n6472), .B1(n6547), .B2(n5211), .ZN(n5213)
         );
  AOI21_X1 U6440 ( .B1(n6543), .B2(n5214), .A(n5213), .ZN(n5215) );
  OAI211_X1 U6441 ( .C1(n5217), .C2(n5399), .A(n5216), .B(n5215), .ZN(U3025)
         );
  CLKBUF_X1 U6442 ( .A(n5218), .Z(n5220) );
  XNOR2_X1 U6443 ( .A(n5220), .B(n5219), .ZN(n5290) );
  NOR2_X1 U6444 ( .A1(n5222), .A2(n5221), .ZN(n5223) );
  OR2_X1 U6445 ( .A1(n5224), .A2(n5223), .ZN(n6193) );
  OAI22_X1 U6446 ( .A1(n6193), .A2(n6424), .B1(n6649), .B2(n6434), .ZN(n5229)
         );
  INV_X1 U6447 ( .A(n5340), .ZN(n5342) );
  AOI211_X1 U6448 ( .C1(n6387), .C2(n5227), .A(n5342), .B(n6384), .ZN(n5228)
         );
  AOI211_X1 U6449 ( .C1(INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n5230), .A(n5229), 
        .B(n5228), .ZN(n5231) );
  OAI21_X1 U6450 ( .B1(n6425), .B2(n5290), .A(n5231), .ZN(U3010) );
  NAND2_X1 U6451 ( .A1(n5232), .A2(n6439), .ZN(n5241) );
  NAND3_X1 U6452 ( .A1(n5272), .A2(n6442), .A3(n5233), .ZN(n5234) );
  NAND2_X1 U6453 ( .A1(n5234), .A2(n6444), .ZN(n5239) );
  NOR2_X1 U6454 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5235), .ZN(n5270)
         );
  OAI211_X1 U6455 ( .C1(n6702), .C2(n5270), .A(n5237), .B(n5236), .ZN(n5238)
         );
  INV_X1 U6456 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5245) );
  OAI22_X1 U6457 ( .A1(n5241), .A2(n6729), .B1(n6446), .B2(n5240), .ZN(n5274)
         );
  AOI22_X1 U6458 ( .A1(n6525), .A2(n5270), .B1(n6459), .B2(n6495), .ZN(n5242)
         );
  OAI21_X1 U6459 ( .B1(n5272), .B2(n6462), .A(n5242), .ZN(n5243) );
  AOI21_X1 U6460 ( .B1(n6526), .B2(n5274), .A(n5243), .ZN(n5244) );
  OAI21_X1 U6461 ( .B1(n5277), .B2(n5245), .A(n5244), .ZN(U3086) );
  INV_X1 U6462 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5249) );
  AOI22_X1 U6463 ( .A1(n6537), .A2(n5270), .B1(n6536), .B2(n6495), .ZN(n5246)
         );
  OAI21_X1 U6464 ( .B1(n5272), .B2(n6541), .A(n5246), .ZN(n5247) );
  AOI21_X1 U6465 ( .B1(n6538), .B2(n5274), .A(n5247), .ZN(n5248) );
  OAI21_X1 U6466 ( .B1(n5277), .B2(n5249), .A(n5248), .ZN(U3088) );
  INV_X1 U6467 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5253) );
  AOI22_X1 U6468 ( .A1(n6550), .A2(n5270), .B1(n6548), .B2(n6495), .ZN(n5250)
         );
  OAI21_X1 U6469 ( .B1(n5272), .B2(n6555), .A(n5250), .ZN(n5251) );
  AOI21_X1 U6470 ( .B1(n6551), .B2(n5274), .A(n5251), .ZN(n5252) );
  OAI21_X1 U6471 ( .B1(n5277), .B2(n5253), .A(n5252), .ZN(U3090) );
  INV_X1 U6472 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5257) );
  AOI22_X1 U6473 ( .A1(n6519), .A2(n5270), .B1(n6455), .B2(n6495), .ZN(n5254)
         );
  OAI21_X1 U6474 ( .B1(n5272), .B2(n6458), .A(n5254), .ZN(n5255) );
  AOI21_X1 U6475 ( .B1(n6520), .B2(n5274), .A(n5255), .ZN(n5256) );
  OAI21_X1 U6476 ( .B1(n5277), .B2(n5257), .A(n5256), .ZN(U3085) );
  INV_X1 U6477 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5261) );
  AOI22_X1 U6478 ( .A1(n6559), .A2(n5270), .B1(n6478), .B2(n6495), .ZN(n5258)
         );
  OAI21_X1 U6479 ( .B1(n5272), .B2(n6482), .A(n5258), .ZN(n5259) );
  AOI21_X1 U6480 ( .B1(n6561), .B2(n5274), .A(n5259), .ZN(n5260) );
  OAI21_X1 U6481 ( .B1(n5277), .B2(n5261), .A(n5260), .ZN(U3091) );
  INV_X1 U6482 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5265) );
  AOI22_X1 U6483 ( .A1(n6543), .A2(n5270), .B1(n6469), .B2(n6495), .ZN(n5262)
         );
  OAI21_X1 U6484 ( .B1(n5272), .B2(n6472), .A(n5262), .ZN(n5263) );
  AOI21_X1 U6485 ( .B1(n6544), .B2(n5274), .A(n5263), .ZN(n5264) );
  OAI21_X1 U6486 ( .B1(n5277), .B2(n5265), .A(n5264), .ZN(U3089) );
  INV_X1 U6487 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5269) );
  AOI22_X1 U6488 ( .A1(n6504), .A2(n5270), .B1(n6451), .B2(n6495), .ZN(n5266)
         );
  OAI21_X1 U6489 ( .B1(n5272), .B2(n6454), .A(n5266), .ZN(n5267) );
  AOI21_X1 U6490 ( .B1(n6514), .B2(n5274), .A(n5267), .ZN(n5268) );
  OAI21_X1 U6491 ( .B1(n5277), .B2(n5269), .A(n5268), .ZN(U3084) );
  INV_X1 U6492 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5276) );
  AOI22_X1 U6493 ( .A1(n6531), .A2(n5270), .B1(n6463), .B2(n6495), .ZN(n5271)
         );
  OAI21_X1 U6494 ( .B1(n5272), .B2(n6466), .A(n5271), .ZN(n5273) );
  AOI21_X1 U6495 ( .B1(n6532), .B2(n5274), .A(n5273), .ZN(n5275) );
  OAI21_X1 U6496 ( .B1(n5277), .B2(n5276), .A(n5275), .ZN(U3087) );
  INV_X1 U6497 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5278) );
  OAI222_X1 U6498 ( .A1(n5279), .A2(n5808), .B1(n5278), .B2(n5814), .C1(n5796), 
        .C2(n5321), .ZN(U2850) );
  AOI21_X1 U6499 ( .B1(n5281), .B2(n5048), .A(n5280), .ZN(n6197) );
  INV_X1 U6500 ( .A(n6197), .ZN(n5283) );
  AOI22_X1 U6501 ( .A1(n6742), .A2(DATAI_8_), .B1(n6743), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n5282) );
  OAI21_X1 U6502 ( .B1(n5283), .B2(n5834), .A(n5282), .ZN(U2883) );
  OAI22_X1 U6503 ( .A1(n6193), .A2(n5808), .B1(n6913), .B2(n5814), .ZN(n5284)
         );
  AOI21_X1 U6504 ( .B1(n6197), .B2(n5810), .A(n5284), .ZN(n5285) );
  INV_X1 U6505 ( .A(n5285), .ZN(U2851) );
  INV_X1 U6506 ( .A(n6195), .ZN(n5287) );
  AOI22_X1 U6507 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n3952), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n5286) );
  OAI21_X1 U6508 ( .B1(n6352), .B2(n5287), .A(n5286), .ZN(n5288) );
  AOI21_X1 U6509 ( .B1(n6197), .B2(n6347), .A(n5288), .ZN(n5289) );
  OAI21_X1 U6510 ( .B1(n6355), .B2(n5290), .A(n5289), .ZN(U2978) );
  NAND2_X1 U6511 ( .A1(n6732), .A2(n3146), .ZN(n5292) );
  INV_X1 U6512 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6724) );
  OAI22_X1 U6513 ( .A1(n6180), .A2(n5293), .B1(n6205), .B2(n6724), .ZN(n5294)
         );
  INV_X1 U6514 ( .A(n5294), .ZN(n5301) );
  NAND2_X1 U6515 ( .A1(n6732), .A2(n5295), .ZN(n6255) );
  OAI21_X1 U6516 ( .B1(n6239), .B2(n6196), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5296) );
  OAI21_X1 U6517 ( .B1(n6255), .B2(n5297), .A(n5296), .ZN(n5298) );
  AOI21_X1 U6518 ( .B1(n6155), .B2(n5299), .A(n5298), .ZN(n5300) );
  OAI211_X1 U6519 ( .C1(n6260), .C2(n6362), .A(n5301), .B(n5300), .ZN(U2827)
         );
  CLKBUF_X1 U6520 ( .A(n5302), .Z(n5303) );
  OAI21_X1 U6521 ( .B1(n5303), .B2(n5306), .A(n5305), .ZN(n5751) );
  AND2_X1 U6522 ( .A1(n5346), .A2(n5307), .ZN(n5308) );
  NOR2_X1 U6523 ( .A1(n5357), .A2(n5308), .ZN(n6363) );
  INV_X1 U6524 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5747) );
  NOR2_X1 U6525 ( .A1(n5814), .A2(n5747), .ZN(n5309) );
  AOI21_X1 U6526 ( .B1(n6363), .B2(n5811), .A(n5309), .ZN(n5310) );
  OAI21_X1 U6527 ( .B1(n5751), .B2(n5796), .A(n5310), .ZN(U2848) );
  INV_X1 U6528 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6287) );
  OAI222_X1 U6529 ( .A1(n5751), .A2(n5834), .B1(n5481), .B2(n6844), .C1(n5816), 
        .C2(n6287), .ZN(U2880) );
  AND2_X1 U6530 ( .A1(n5312), .A2(n5311), .ZN(n5313) );
  NOR2_X1 U6531 ( .A1(n5303), .A2(n5313), .ZN(n6188) );
  INV_X1 U6532 ( .A(n6188), .ZN(n5351) );
  AOI22_X1 U6533 ( .A1(n6742), .A2(DATAI_10_), .B1(n6743), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5314) );
  OAI21_X1 U6534 ( .B1(n5351), .B2(n5834), .A(n5314), .ZN(U2881) );
  XNOR2_X1 U6535 ( .A(n5880), .B(n6377), .ZN(n5316) );
  XNOR2_X1 U6536 ( .A(n5330), .B(n5316), .ZN(n6373) );
  NAND2_X1 U6537 ( .A1(n6373), .A2(n4310), .ZN(n5320) );
  NOR2_X1 U6538 ( .A1(n6434), .A2(n6651), .ZN(n6371) );
  NOR2_X1 U6539 ( .A1(n6352), .A2(n5317), .ZN(n5318) );
  AOI211_X1 U6540 ( .C1(n6358), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6371), 
        .B(n5318), .ZN(n5319) );
  OAI211_X1 U6541 ( .C1(n6361), .C2(n5321), .A(n5320), .B(n5319), .ZN(U2977)
         );
  INV_X1 U6542 ( .A(n6351), .ZN(n5322) );
  AOI22_X1 U6543 ( .A1(n6239), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n6196), 
        .B2(n5322), .ZN(n5324) );
  INV_X1 U6544 ( .A(REIP_REG_2__SCAN_IN), .ZN(n5325) );
  NAND3_X1 U6545 ( .A1(n6246), .A2(REIP_REG_1__SCAN_IN), .A3(n5325), .ZN(n5323) );
  OAI211_X1 U6546 ( .C1(n6257), .C2(n6406), .A(n5324), .B(n5323), .ZN(n5327)
         );
  INV_X1 U6547 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5755) );
  AND2_X1 U6548 ( .A1(n6246), .A2(n5755), .ZN(n5757) );
  NOR2_X1 U6549 ( .A1(n5757), .A2(n6236), .ZN(n6251) );
  OAI22_X1 U6550 ( .A1(n6251), .A2(n5325), .B1(n6014), .B2(n6255), .ZN(n5326)
         );
  AOI211_X1 U6551 ( .C1(EBX_REG_2__SCAN_IN), .C2(n6264), .A(n5327), .B(n5326), 
        .ZN(n5328) );
  OAI21_X1 U6552 ( .B1(n6346), .B2(n6260), .A(n5328), .ZN(U2825) );
  OR2_X1 U6553 ( .A1(n5330), .A2(n5329), .ZN(n5332) );
  NAND2_X1 U6554 ( .A1(n5332), .A2(n5331), .ZN(n5335) );
  NAND2_X1 U6555 ( .A1(n3165), .A2(n5333), .ZN(n5334) );
  XNOR2_X1 U6556 ( .A(n5335), .B(n5334), .ZN(n5350) );
  AOI22_X1 U6557 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n3952), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5336) );
  OAI21_X1 U6558 ( .B1(n6352), .B2(n5337), .A(n5336), .ZN(n5338) );
  AOI21_X1 U6559 ( .B1(n6188), .B2(n6347), .A(n5338), .ZN(n5339) );
  OAI21_X1 U6560 ( .B1(n5350), .B2(n6355), .A(n5339), .ZN(U2976) );
  NOR2_X1 U6561 ( .A1(n5340), .A2(n6384), .ZN(n6374) );
  OAI211_X1 U6562 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6374), .B(n5341), .ZN(n5349) );
  OAI21_X1 U6563 ( .B1(n5342), .B2(n6414), .A(n6388), .ZN(n6370) );
  NAND2_X1 U6564 ( .A1(n5344), .A2(n5343), .ZN(n5345) );
  NAND2_X1 U6565 ( .A1(n5346), .A2(n5345), .ZN(n6181) );
  OAI22_X1 U6566 ( .A1(n6181), .A2(n6424), .B1(n6653), .B2(n6434), .ZN(n5347)
         );
  AOI21_X1 U6567 ( .B1(n6370), .B2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n5347), 
        .ZN(n5348) );
  OAI211_X1 U6568 ( .C1(n5350), .C2(n6425), .A(n5349), .B(n5348), .ZN(U3008)
         );
  INV_X1 U6569 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6179) );
  OAI222_X1 U6570 ( .A1(n6181), .A2(n5808), .B1(n6179), .B2(n5814), .C1(n5351), 
        .C2(n5796), .ZN(U2849) );
  INV_X1 U6571 ( .A(n5465), .ZN(n5353) );
  NOR2_X1 U6572 ( .A1(n5463), .A2(n5353), .ZN(n5354) );
  XNOR2_X1 U6573 ( .A(n5464), .B(n5354), .ZN(n5492) );
  AOI22_X1 U6574 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n5450), .B1(n5355), .B2(n6414), .ZN(n5361) );
  NOR2_X1 U6575 ( .A1(n5357), .A2(n5356), .ZN(n5358) );
  OR2_X1 U6576 ( .A1(n5438), .A2(n5358), .ZN(n6166) );
  INV_X1 U6577 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6808) );
  OAI22_X1 U6578 ( .A1(n6166), .A2(n6424), .B1(n6808), .B2(n6434), .ZN(n5360)
         );
  INV_X1 U6579 ( .A(n6366), .ZN(n6094) );
  NOR3_X1 U6580 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6094), .A3(n6365), 
        .ZN(n5359) );
  AOI211_X1 U6581 ( .C1(n5361), .C2(INSTADDRPOINTER_REG_12__SCAN_IN), .A(n5360), .B(n5359), .ZN(n5362) );
  OAI21_X1 U6582 ( .B1(n5492), .B2(n6425), .A(n5362), .ZN(U3006) );
  NAND2_X1 U6583 ( .A1(n5305), .A2(n5364), .ZN(n5365) );
  NAND2_X1 U6584 ( .A1(n5436), .A2(n5365), .ZN(n6172) );
  INV_X1 U6585 ( .A(DATAI_12_), .ZN(n5366) );
  OAI222_X1 U6586 ( .A1(n6172), .A2(n5834), .B1(n5816), .B2(n5367), .C1(n5366), 
        .C2(n5481), .ZN(U2879) );
  AND2_X1 U6587 ( .A1(n5369), .A2(n5368), .ZN(n5373) );
  NAND2_X1 U6588 ( .A1(n5371), .A2(n5370), .ZN(n5372) );
  XNOR2_X1 U6589 ( .A(n5373), .B(n5372), .ZN(n6364) );
  INV_X1 U6590 ( .A(n6364), .ZN(n5378) );
  INV_X1 U6591 ( .A(n5751), .ZN(n5376) );
  AOI22_X1 U6592 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .B1(n3952), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n5374) );
  OAI21_X1 U6593 ( .B1(n5741), .B2(n6352), .A(n5374), .ZN(n5375) );
  AOI21_X1 U6594 ( .B1(n5376), .B2(n6347), .A(n5375), .ZN(n5377) );
  OAI21_X1 U6595 ( .B1(n5378), .B2(n6355), .A(n5377), .ZN(U2975) );
  INV_X1 U6596 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6165) );
  OAI222_X1 U6597 ( .A1(n6166), .A2(n5808), .B1(n6165), .B2(n5814), .C1(n6172), 
        .C2(n5796), .ZN(U2847) );
  AND2_X1 U6598 ( .A1(n4640), .A2(n5379), .ZN(n5380) );
  NAND2_X1 U6599 ( .A1(n5381), .A2(n5380), .ZN(n6565) );
  OAI21_X1 U6600 ( .B1(n5431), .B2(n6549), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5382) );
  NOR3_X1 U6601 ( .A1(n6446), .A2(n7014), .A3(n5384), .ZN(n5385) );
  NAND3_X1 U6602 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6586), .ZN(n6511) );
  OR2_X1 U6603 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6511), .ZN(n5428)
         );
  INV_X1 U6604 ( .A(n6507), .ZN(n5386) );
  AOI22_X1 U6605 ( .A1(n5387), .A2(n5386), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5428), .ZN(n5388) );
  OAI211_X1 U6606 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6935), .A(n5389), .B(n5388), .ZN(n5426) );
  AOI22_X1 U6607 ( .A1(n6549), .A2(n6556), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5426), .ZN(n5390) );
  OAI21_X1 U6608 ( .B1(n5391), .B2(n5428), .A(n5390), .ZN(n5392) );
  AOI21_X1 U6609 ( .B1(n5431), .B2(n6478), .A(n5392), .ZN(n5393) );
  OAI21_X1 U6610 ( .B1(n5434), .B2(n5394), .A(n5393), .ZN(U3107) );
  AOI22_X1 U6611 ( .A1(n6549), .A2(n6542), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5426), .ZN(n5395) );
  OAI21_X1 U6612 ( .B1(n5396), .B2(n5428), .A(n5395), .ZN(n5397) );
  AOI21_X1 U6613 ( .B1(n5431), .B2(n6469), .A(n5397), .ZN(n5398) );
  OAI21_X1 U6614 ( .B1(n5434), .B2(n5399), .A(n5398), .ZN(U3105) );
  AOI22_X1 U6615 ( .A1(n6549), .A2(n6491), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5426), .ZN(n5400) );
  OAI21_X1 U6616 ( .B1(n5401), .B2(n5428), .A(n5400), .ZN(n5402) );
  AOI21_X1 U6617 ( .B1(n5431), .B2(n6548), .A(n5402), .ZN(n5403) );
  OAI21_X1 U6618 ( .B1(n5434), .B2(n5404), .A(n5403), .ZN(U3106) );
  AOI22_X1 U6619 ( .A1(n6549), .A2(n6524), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5426), .ZN(n5405) );
  OAI21_X1 U6620 ( .B1(n5406), .B2(n5428), .A(n5405), .ZN(n5407) );
  AOI21_X1 U6621 ( .B1(n5431), .B2(n6459), .A(n5407), .ZN(n5408) );
  OAI21_X1 U6622 ( .B1(n5434), .B2(n5409), .A(n5408), .ZN(U3102) );
  AOI22_X1 U6623 ( .A1(n6549), .A2(n6530), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5426), .ZN(n5410) );
  OAI21_X1 U6624 ( .B1(n5411), .B2(n5428), .A(n5410), .ZN(n5412) );
  AOI21_X1 U6625 ( .B1(n5431), .B2(n6463), .A(n5412), .ZN(n5413) );
  OAI21_X1 U6626 ( .B1(n5434), .B2(n5414), .A(n5413), .ZN(U3103) );
  AOI22_X1 U6627 ( .A1(n6549), .A2(n5415), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5426), .ZN(n5416) );
  OAI21_X1 U6628 ( .B1(n5417), .B2(n5428), .A(n5416), .ZN(n5418) );
  AOI21_X1 U6629 ( .B1(n5431), .B2(n6536), .A(n5418), .ZN(n5419) );
  OAI21_X1 U6630 ( .B1(n5434), .B2(n5420), .A(n5419), .ZN(U3104) );
  AOI22_X1 U6631 ( .A1(n6549), .A2(n6518), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5426), .ZN(n5421) );
  OAI21_X1 U6632 ( .B1(n5422), .B2(n5428), .A(n5421), .ZN(n5423) );
  AOI21_X1 U6633 ( .B1(n5431), .B2(n6455), .A(n5423), .ZN(n5424) );
  OAI21_X1 U6634 ( .B1(n5434), .B2(n5425), .A(n5424), .ZN(U3101) );
  AOI22_X1 U6635 ( .A1(n6549), .A2(n6503), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5426), .ZN(n5427) );
  OAI21_X1 U6636 ( .B1(n5429), .B2(n5428), .A(n5427), .ZN(n5430) );
  AOI21_X1 U6637 ( .B1(n6451), .B2(n5431), .A(n5430), .ZN(n5432) );
  OAI21_X1 U6638 ( .B1(n5434), .B2(n5433), .A(n5432), .ZN(U3100) );
  XNOR2_X1 U6639 ( .A(n5436), .B(n5435), .ZN(n6159) );
  OAI21_X1 U6640 ( .B1(n5438), .B2(n5437), .A(n5454), .ZN(n5439) );
  INV_X1 U6641 ( .A(n5439), .ZN(n6156) );
  AOI22_X1 U6642 ( .A1(n6156), .A2(n5811), .B1(n5805), .B2(EBX_REG_13__SCAN_IN), .ZN(n5440) );
  OAI21_X1 U6643 ( .B1(n6159), .B2(n5796), .A(n5440), .ZN(U2846) );
  OR2_X1 U6644 ( .A1(n5464), .A2(n5441), .ZN(n5468) );
  NAND2_X1 U6645 ( .A1(n5468), .A2(n5442), .ZN(n5445) );
  XNOR2_X1 U6646 ( .A(n5989), .B(n5443), .ZN(n5444) );
  XNOR2_X1 U6647 ( .A(n5445), .B(n5444), .ZN(n5928) );
  NAND3_X1 U6648 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n6758), .ZN(n5475) );
  AOI221_X1 U6649 ( .B1(n5447), .B2(n5446), .C1(n5474), .C2(n5446), .A(n5475), 
        .ZN(n5472) );
  INV_X1 U6650 ( .A(n6415), .ZN(n6431) );
  NAND2_X1 U6651 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5448) );
  AOI22_X1 U6652 ( .A1(n6431), .A2(n5452), .B1(n5448), .B2(n6429), .ZN(n5449)
         );
  NAND2_X1 U6653 ( .A1(n5450), .A2(n5449), .ZN(n5473) );
  OAI21_X1 U6654 ( .B1(n5472), .B2(n5473), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5451) );
  INV_X1 U6655 ( .A(n5451), .ZN(n5457) );
  NOR3_X1 U6656 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6094), .A3(n5452), 
        .ZN(n5456) );
  XNOR2_X1 U6657 ( .A(n5454), .B(n5453), .ZN(n6145) );
  INV_X1 U6658 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6659) );
  OAI22_X1 U6659 ( .A1(n6145), .A2(n6424), .B1(n6659), .B2(n6434), .ZN(n5455)
         );
  NOR3_X1 U6660 ( .A1(n5457), .A2(n5456), .A3(n5455), .ZN(n5458) );
  OAI21_X1 U6661 ( .B1(n5928), .B2(n6425), .A(n5458), .ZN(U3004) );
  OAI21_X1 U6662 ( .B1(n5461), .B2(n5460), .A(n5459), .ZN(n6147) );
  INV_X1 U6663 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5462) );
  OAI222_X1 U6664 ( .A1(n6147), .A2(n5796), .B1(n5808), .B2(n6145), .C1(n5462), 
        .C2(n5814), .ZN(U2845) );
  OR2_X1 U6665 ( .A1(n5464), .A2(n5463), .ZN(n5466) );
  NAND2_X1 U6666 ( .A1(n5466), .A2(n5465), .ZN(n5471) );
  AND2_X1 U6667 ( .A1(n5468), .A2(n5467), .ZN(n5469) );
  OAI21_X1 U6668 ( .B1(n5471), .B2(n5470), .A(n5469), .ZN(n5483) );
  INV_X1 U6669 ( .A(n5483), .ZN(n5480) );
  AOI21_X1 U6670 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5473), .A(n5472), 
        .ZN(n5479) );
  INV_X1 U6671 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6657) );
  NOR2_X1 U6672 ( .A1(n6434), .A2(n6657), .ZN(n5477) );
  NOR3_X1 U6673 ( .A1(n6415), .A2(n5475), .A3(n5474), .ZN(n5476) );
  AOI211_X1 U6674 ( .C1(n6156), .C2(n6390), .A(n5477), .B(n5476), .ZN(n5478)
         );
  OAI211_X1 U6675 ( .C1(n5480), .C2(n6425), .A(n5479), .B(n5478), .ZN(U3005)
         );
  INV_X1 U6676 ( .A(DATAI_13_), .ZN(n6822) );
  OAI222_X1 U6677 ( .A1(n5816), .A2(n5482), .B1(n5481), .B2(n6822), .C1(n5834), 
        .C2(n6159), .ZN(U2878) );
  NAND2_X1 U6678 ( .A1(n5483), .A2(n4310), .ZN(n5487) );
  INV_X1 U6679 ( .A(n6158), .ZN(n5485) );
  OAI22_X1 U6680 ( .A1(n6342), .A2(n6981), .B1(n6434), .B2(n6657), .ZN(n5484)
         );
  AOI21_X1 U6681 ( .B1(n5485), .B2(n6336), .A(n5484), .ZN(n5486) );
  OAI211_X1 U6682 ( .C1(n6159), .C2(n6361), .A(n5487), .B(n5486), .ZN(U2973)
         );
  INV_X1 U6683 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5488) );
  OAI22_X1 U6684 ( .A1(n6342), .A2(n5488), .B1(n6434), .B2(n6808), .ZN(n5490)
         );
  NOR2_X1 U6685 ( .A1(n6172), .A2(n6361), .ZN(n5489) );
  AOI211_X1 U6686 ( .C1(n6336), .C2(n6169), .A(n5490), .B(n5489), .ZN(n5491)
         );
  OAI21_X1 U6687 ( .B1(n5492), .B2(n6355), .A(n5491), .ZN(U2974) );
  NOR3_X1 U6688 ( .A1(n6743), .A2(n5815), .A3(n5493), .ZN(n5494) );
  AOI22_X1 U6689 ( .A1(n6273), .A2(DATAI_11_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6743), .ZN(n5497) );
  NAND2_X1 U6690 ( .A1(n6271), .A2(DATAI_27_), .ZN(n5496) );
  OAI211_X1 U6691 ( .C1(n5853), .C2(n5834), .A(n5497), .B(n5496), .ZN(U2864)
         );
  AOI22_X1 U6692 ( .A1(n6273), .A2(DATAI_9_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6743), .ZN(n5500) );
  NAND2_X1 U6693 ( .A1(n6271), .A2(DATAI_25_), .ZN(n5499) );
  OAI211_X1 U6694 ( .C1(n4052), .C2(n5834), .A(n5500), .B(n5499), .ZN(U2866)
         );
  OAI22_X1 U6695 ( .A1(n6068), .A2(n5808), .B1(n5501), .B2(n5814), .ZN(n5502)
         );
  INV_X1 U6696 ( .A(n5502), .ZN(n5503) );
  OAI21_X1 U6697 ( .B1(n4052), .B2(n5796), .A(n5503), .ZN(U2834) );
  OAI21_X1 U6698 ( .B1(n5506), .B2(n5505), .A(n5504), .ZN(n6070) );
  INV_X1 U6699 ( .A(n6070), .ZN(n5512) );
  INV_X1 U6700 ( .A(n5507), .ZN(n5509) );
  AOI22_X1 U6701 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .B1(n3952), 
        .B2(REIP_REG_25__SCAN_IN), .ZN(n5508) );
  OAI21_X1 U6702 ( .B1(n5509), .B2(n6352), .A(n5508), .ZN(n5510) );
  AOI21_X1 U6703 ( .B1(n5498), .B2(n6347), .A(n5510), .ZN(n5511) );
  OAI21_X1 U6704 ( .B1(n5512), .B2(n6355), .A(n5511), .ZN(U2961) );
  OAI22_X1 U6705 ( .A1(n5513), .A2(n5808), .B1(n5514), .B2(n5814), .ZN(U2828)
         );
  INV_X1 U6706 ( .A(n4442), .ZN(n5517) );
  AOI21_X1 U6707 ( .B1(n5566), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5565), 
        .ZN(n5519) );
  AOI21_X1 U6708 ( .B1(n5521), .B2(n5578), .A(n5520), .ZN(n5593) );
  NAND2_X1 U6709 ( .A1(n3952), .A2(REIP_REG_30__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U6710 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5522)
         );
  OAI211_X1 U6711 ( .C1(n6352), .C2(n5596), .A(n5532), .B(n5522), .ZN(n5523)
         );
  AOI21_X1 U6712 ( .B1(n5593), .B2(n6347), .A(n5523), .ZN(n5524) );
  OAI21_X1 U6713 ( .B1(n5539), .B2(n6355), .A(n5524), .ZN(U2956) );
  INV_X1 U6714 ( .A(n5569), .ZN(n5615) );
  INV_X1 U6715 ( .A(n5528), .ZN(n5525) );
  AOI211_X1 U6716 ( .C1(n5780), .C2(n5569), .A(n5528), .B(n5527), .ZN(n5529)
         );
  AOI21_X1 U6717 ( .B1(n5531), .B2(n5530), .A(n5529), .ZN(n5601) );
  INV_X1 U6718 ( .A(n5601), .ZN(n5765) );
  NAND3_X1 U6719 ( .A1(n5576), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5518), .ZN(n5536) );
  INV_X1 U6720 ( .A(n5532), .ZN(n5533) );
  OAI21_X1 U6721 ( .B1(n5539), .B2(n6425), .A(n5538), .ZN(U2988) );
  INV_X1 U6722 ( .A(n5551), .ZN(n5543) );
  INV_X1 U6723 ( .A(n6705), .ZN(n5558) );
  INV_X1 U6724 ( .A(n6582), .ZN(n5541) );
  NOR2_X1 U6725 ( .A1(n6122), .A2(n6699), .ZN(n5540) );
  AOI21_X1 U6726 ( .B1(n5541), .B2(n6606), .A(n5540), .ZN(n6107) );
  INV_X1 U6727 ( .A(n5542), .ZN(n6700) );
  NAND2_X1 U6728 ( .A1(n6107), .A2(n6700), .ZN(n6713) );
  AOI21_X1 U6729 ( .B1(n5543), .B2(n5558), .A(n6707), .ZN(n5549) );
  INV_X1 U6730 ( .A(n6715), .ZN(n6109) );
  INV_X1 U6731 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5544) );
  AOI22_X1 U6732 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5544), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6900), .ZN(n5556) );
  NAND2_X1 U6733 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5550) );
  NAND3_X1 U6734 ( .A1(n5551), .A2(n3170), .A3(n5558), .ZN(n5545) );
  OAI21_X1 U6735 ( .B1(n5556), .B2(n5550), .A(n5545), .ZN(n5546) );
  AOI21_X1 U6736 ( .B1(n5547), .B2(n6109), .A(n5546), .ZN(n5548) );
  OAI22_X1 U6737 ( .A1(n5549), .A2(n4622), .B1(n5548), .B2(n6707), .ZN(U3459)
         );
  OAI21_X1 U6738 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6705), .A(n6713), 
        .ZN(n6711) );
  INV_X1 U6739 ( .A(n6711), .ZN(n5561) );
  INV_X1 U6740 ( .A(n5550), .ZN(n5555) );
  NOR3_X1 U6741 ( .A1(n4196), .A2(n3177), .A3(n5551), .ZN(n5552) );
  AOI21_X1 U6742 ( .B1(n6576), .B2(n5560), .A(n5552), .ZN(n5553) );
  OAI21_X1 U6743 ( .B1(n6010), .B2(n5554), .A(n5553), .ZN(n6577) );
  AOI222_X1 U6744 ( .A1(n5558), .A2(n5557), .B1(n5556), .B2(n5555), .C1(n6577), 
        .C2(n6109), .ZN(n5559) );
  OAI22_X1 U6745 ( .A1(n5561), .A2(n5560), .B1(n6707), .B2(n5559), .ZN(U3460)
         );
  INV_X1 U6746 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5575) );
  INV_X1 U6747 ( .A(n5562), .ZN(n5563) );
  NOR3_X1 U6748 ( .A1(n5566), .A2(n5563), .A3(n5575), .ZN(n5564) );
  NOR2_X1 U6749 ( .A1(n5567), .A2(n5575), .ZN(n5574) );
  OAI211_X1 U6750 ( .C1(n5780), .C2(n5570), .A(n5569), .B(n5568), .ZN(n5571)
         );
  NAND2_X1 U6751 ( .A1(n5572), .A2(n5571), .ZN(n5591) );
  NAND2_X1 U6752 ( .A1(n3952), .A2(REIP_REG_29__SCAN_IN), .ZN(n5582) );
  OAI21_X1 U6753 ( .B1(n5591), .B2(n6424), .A(n5582), .ZN(n5573) );
  OAI21_X1 U6754 ( .B1(n5588), .B2(n6425), .A(n5577), .ZN(U2989) );
  OAI21_X1 U6755 ( .B1(n6342), .B2(n5583), .A(n5582), .ZN(n5584) );
  OAI21_X1 U6756 ( .B1(n5588), .B2(n6355), .A(n5587), .ZN(U2957) );
  AOI22_X1 U6757 ( .A1(n6271), .A2(DATAI_29_), .B1(n6743), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5590) );
  NAND2_X1 U6758 ( .A1(n6273), .A2(DATAI_13_), .ZN(n5589) );
  OAI211_X1 U6759 ( .C1(n5603), .C2(n5834), .A(n5590), .B(n5589), .ZN(U2862)
         );
  OAI222_X1 U6760 ( .A1(n5796), .A2(n5603), .B1(n5814), .B2(n5592), .C1(n5591), 
        .C2(n5808), .ZN(U2830) );
  INV_X1 U6761 ( .A(n5593), .ZN(n5823) );
  INV_X1 U6762 ( .A(EBX_REG_30__SCAN_IN), .ZN(n6871) );
  INV_X1 U6763 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6686) );
  NOR2_X1 U6764 ( .A1(n5608), .A2(n6686), .ZN(n5595) );
  OAI21_X1 U6765 ( .B1(n5595), .B2(REIP_REG_30__SCAN_IN), .A(n5594), .ZN(n5599) );
  INV_X1 U6766 ( .A(n5596), .ZN(n5597) );
  AOI22_X1 U6767 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n6239), .B1(n6196), 
        .B2(n5597), .ZN(n5598) );
  OAI211_X1 U6768 ( .C1(n6180), .C2(n6871), .A(n5599), .B(n5598), .ZN(n5600)
         );
  AOI21_X1 U6769 ( .B1(n5601), .B2(n6155), .A(n5600), .ZN(n5602) );
  OAI21_X1 U6770 ( .B1(n5823), .B2(n6171), .A(n5602), .ZN(U2797) );
  INV_X1 U6771 ( .A(n5603), .ZN(n5604) );
  NAND2_X1 U6772 ( .A1(n5604), .A2(n6220), .ZN(n5612) );
  AOI22_X1 U6773 ( .A1(EBX_REG_29__SCAN_IN), .A2(n6264), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6239), .ZN(n5605) );
  OAI21_X1 U6774 ( .B1(n5622), .B2(n6686), .A(n5605), .ZN(n5610) );
  INV_X1 U6775 ( .A(n5606), .ZN(n5607) );
  OAI22_X1 U6776 ( .A1(n5608), .A2(REIP_REG_29__SCAN_IN), .B1(n5607), .B2(
        n6258), .ZN(n5609) );
  NOR2_X1 U6777 ( .A1(n5610), .A2(n5609), .ZN(n5611) );
  OAI211_X1 U6778 ( .C1(n6257), .C2(n5591), .A(n5612), .B(n5611), .ZN(U2798)
         );
  AOI21_X1 U6779 ( .B1(n5614), .B2(n5613), .A(n5579), .ZN(n5847) );
  INV_X1 U6780 ( .A(n5847), .ZN(n5826) );
  AOI21_X1 U6781 ( .B1(n5617), .B2(n5616), .A(n5615), .ZN(n5929) );
  AOI21_X1 U6782 ( .B1(n5618), .B2(REIP_REG_27__SCAN_IN), .A(
        REIP_REG_28__SCAN_IN), .ZN(n5623) );
  OAI22_X1 U6783 ( .A1(n5619), .A2(n6253), .B1(n6258), .B2(n5845), .ZN(n5620)
         );
  AOI21_X1 U6784 ( .B1(EBX_REG_28__SCAN_IN), .B2(n6264), .A(n5620), .ZN(n5621)
         );
  OAI21_X1 U6785 ( .B1(n5623), .B2(n5622), .A(n5621), .ZN(n5624) );
  AOI21_X1 U6786 ( .B1(n5929), .B2(n6155), .A(n5624), .ZN(n5625) );
  OAI21_X1 U6787 ( .B1(n5826), .B2(n6171), .A(n5625), .ZN(U2799) );
  OR2_X1 U6788 ( .A1(n4336), .A2(n5626), .ZN(n5627) );
  NAND2_X1 U6789 ( .A1(n5628), .A2(n5627), .ZN(n5952) );
  OAI22_X1 U6790 ( .A1(n6180), .A2(n5768), .B1(n5629), .B2(n6258), .ZN(n5630)
         );
  AOI21_X1 U6791 ( .B1(n6239), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5630), 
        .ZN(n5635) );
  INV_X1 U6792 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6679) );
  OAI21_X1 U6793 ( .B1(n6846), .B2(n5631), .A(n6679), .ZN(n5633) );
  NAND2_X1 U6794 ( .A1(n5633), .A2(n5632), .ZN(n5634) );
  OAI211_X1 U6795 ( .C1(n5952), .C2(n6257), .A(n5635), .B(n5634), .ZN(n5636)
         );
  AOI21_X1 U6796 ( .B1(n5637), .B2(n6220), .A(n5636), .ZN(n5638) );
  INV_X1 U6797 ( .A(n5638), .ZN(U2801) );
  NAND2_X1 U6798 ( .A1(n5639), .A2(n5640), .ZN(n5641) );
  AOI21_X1 U6799 ( .B1(n5644), .B2(n5654), .A(n5643), .ZN(n5957) );
  OAI22_X1 U6800 ( .A1(n5657), .A2(n6677), .B1(n5645), .B2(n6253), .ZN(n5648)
         );
  INV_X1 U6801 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5646) );
  OAI22_X1 U6802 ( .A1(n6180), .A2(n5646), .B1(n5869), .B2(n6258), .ZN(n5647)
         );
  AOI211_X1 U6803 ( .C1(n5957), .C2(n6155), .A(n5648), .B(n5647), .ZN(n5650)
         );
  OAI211_X1 U6804 ( .C1(n5772), .C2(n6171), .A(n5650), .B(n5649), .ZN(U2803)
         );
  NAND2_X1 U6805 ( .A1(n5674), .A2(n5652), .ZN(n5653) );
  NAND2_X1 U6806 ( .A1(n5654), .A2(n5653), .ZN(n5964) );
  OR2_X1 U6807 ( .A1(n4411), .A2(n5655), .ZN(n5656) );
  NAND2_X1 U6808 ( .A1(n5878), .A2(n6220), .ZN(n5665) );
  INV_X1 U6809 ( .A(n5657), .ZN(n5663) );
  OAI21_X1 U6810 ( .B1(n6955), .B2(n5679), .A(n6674), .ZN(n5662) );
  INV_X1 U6811 ( .A(n5658), .ZN(n5876) );
  NOR2_X1 U6812 ( .A1(n6258), .A2(n5876), .ZN(n5661) );
  INV_X1 U6813 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5773) );
  OAI22_X1 U6814 ( .A1(n6180), .A2(n5773), .B1(n5659), .B2(n6253), .ZN(n5660)
         );
  AOI211_X1 U6815 ( .C1(n5663), .C2(n5662), .A(n5661), .B(n5660), .ZN(n5664)
         );
  OAI211_X1 U6816 ( .C1(n6257), .C2(n5964), .A(n5665), .B(n5664), .ZN(U2804)
         );
  INV_X1 U6817 ( .A(n5668), .ZN(n5684) );
  INV_X1 U6818 ( .A(n5669), .ZN(n5670) );
  AOI21_X1 U6819 ( .B1(n5667), .B2(n5684), .A(n5670), .ZN(n5671) );
  OR2_X1 U6820 ( .A1(n4411), .A2(n5671), .ZN(n5883) );
  OR2_X1 U6821 ( .A1(n5687), .A2(n5672), .ZN(n5673) );
  NAND2_X1 U6822 ( .A1(n5674), .A2(n5673), .ZN(n5975) );
  INV_X1 U6823 ( .A(n5975), .ZN(n5682) );
  INV_X1 U6824 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5776) );
  INV_X1 U6825 ( .A(n5885), .ZN(n5676) );
  OAI21_X1 U6826 ( .B1(n6236), .B2(n5690), .A(n6235), .ZN(n6020) );
  NAND2_X1 U6827 ( .A1(n6246), .A2(n6670), .ZN(n5689) );
  AOI21_X1 U6828 ( .B1(n6020), .B2(n5689), .A(n6955), .ZN(n5675) );
  AOI21_X1 U6829 ( .B1(n6196), .B2(n5676), .A(n5675), .ZN(n5677) );
  OAI21_X1 U6830 ( .B1(n6180), .B2(n5776), .A(n5677), .ZN(n5681) );
  INV_X1 U6831 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5678) );
  OAI22_X1 U6832 ( .A1(REIP_REG_22__SCAN_IN), .A2(n5679), .B1(n5678), .B2(
        n6253), .ZN(n5680) );
  AOI211_X1 U6833 ( .C1(n6155), .C2(n5682), .A(n5681), .B(n5680), .ZN(n5683)
         );
  OAI21_X1 U6834 ( .B1(n5883), .B2(n6171), .A(n5683), .ZN(U2805) );
  XNOR2_X1 U6835 ( .A(n5667), .B(n5684), .ZN(n6047) );
  AND2_X1 U6836 ( .A1(n5686), .A2(n5685), .ZN(n5688) );
  OR2_X1 U6837 ( .A1(n5688), .A2(n5687), .ZN(n5982) );
  OAI22_X1 U6838 ( .A1(n6020), .A2(n6670), .B1(n5891), .B2(n6253), .ZN(n5692)
         );
  NOR2_X1 U6839 ( .A1(n5690), .A2(n5689), .ZN(n5691) );
  AOI211_X1 U6840 ( .C1(n6196), .C2(n5893), .A(n5692), .B(n5691), .ZN(n5694)
         );
  NAND2_X1 U6841 ( .A1(n6264), .A2(EBX_REG_21__SCAN_IN), .ZN(n5693) );
  OAI211_X1 U6842 ( .C1(n5982), .C2(n6257), .A(n5694), .B(n5693), .ZN(n5695)
         );
  INV_X1 U6843 ( .A(n5695), .ZN(n5696) );
  OAI21_X1 U6844 ( .B1(n6047), .B2(n6171), .A(n5696), .ZN(U2806) );
  AOI21_X1 U6845 ( .B1(n5699), .B2(n5697), .A(n5798), .ZN(n5909) );
  INV_X1 U6846 ( .A(n5909), .ZN(n5835) );
  OAI21_X1 U6847 ( .B1(n5716), .B2(n5700), .A(n5802), .ZN(n5701) );
  INV_X1 U6848 ( .A(n5701), .ZN(n6086) );
  AOI21_X1 U6849 ( .B1(n6264), .B2(EBX_REG_17__SCAN_IN), .A(n3952), .ZN(n5702)
         );
  OAI21_X1 U6850 ( .B1(n5907), .B2(n6258), .A(n5702), .ZN(n5709) );
  INV_X1 U6851 ( .A(n6246), .ZN(n5740) );
  NOR2_X1 U6852 ( .A1(n5740), .A2(n5703), .ZN(n5720) );
  INV_X1 U6853 ( .A(n5720), .ZN(n5704) );
  NOR2_X1 U6854 ( .A1(n5704), .A2(n6662), .ZN(n6018) );
  NOR2_X1 U6855 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6018), .ZN(n5707) );
  INV_X1 U6856 ( .A(n5705), .ZN(n5706) );
  OAI21_X1 U6857 ( .B1(n6236), .B2(n5706), .A(n6235), .ZN(n6137) );
  OAI22_X1 U6858 ( .A1(n5707), .A2(n6137), .B1(n3720), .B2(n6253), .ZN(n5708)
         );
  AOI211_X1 U6859 ( .C1(n6086), .C2(n6155), .A(n5709), .B(n5708), .ZN(n5710)
         );
  OAI21_X1 U6860 ( .B1(n5835), .B2(n6171), .A(n5710), .ZN(U2810) );
  INV_X1 U6861 ( .A(n5728), .ZN(n5712) );
  NAND2_X1 U6862 ( .A1(n5712), .A2(n5711), .ZN(n5713) );
  AND2_X1 U6863 ( .A1(n5697), .A2(n5713), .ZN(n6272) );
  INV_X1 U6864 ( .A(n6272), .ZN(n5807) );
  NOR2_X1 U6865 ( .A1(n5733), .A2(n5714), .ZN(n5715) );
  OR2_X1 U6866 ( .A1(n5716), .A2(n5715), .ZN(n6095) );
  INV_X1 U6867 ( .A(n6095), .ZN(n5726) );
  INV_X1 U6868 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5809) );
  OAI22_X1 U6869 ( .A1(n5913), .A2(n6258), .B1(n6180), .B2(n5809), .ZN(n5725)
         );
  OAI21_X1 U6871 ( .B1(n5740), .B2(n5717), .A(n5754), .ZN(n6149) );
  INV_X1 U6872 ( .A(n5718), .ZN(n5739) );
  NAND2_X1 U6873 ( .A1(n6246), .A2(n5739), .ZN(n6157) );
  NOR3_X1 U6874 ( .A1(n6157), .A2(REIP_REG_15__SCAN_IN), .A3(n5719), .ZN(n5734) );
  OAI33_X1 U6875 ( .A1(1'b0), .A2(n5720), .A3(REIP_REG_16__SCAN_IN), .B1(n6662), .B2(n6149), .B3(n5734), .ZN(n5722) );
  OAI211_X1 U6876 ( .C1(n6253), .C2(n5723), .A(n5722), .B(n6434), .ZN(n5724)
         );
  AOI211_X1 U6877 ( .C1(n5726), .C2(n6155), .A(n5725), .B(n5724), .ZN(n5727)
         );
  OAI21_X1 U6878 ( .B1(n5807), .B2(n6171), .A(n5727), .ZN(U2811) );
  AOI21_X1 U6879 ( .B1(n5729), .B2(n5459), .A(n5728), .ZN(n5922) );
  INV_X1 U6880 ( .A(n5922), .ZN(n5837) );
  AND2_X1 U6881 ( .A1(n5731), .A2(n5730), .ZN(n5732) );
  NOR2_X1 U6882 ( .A1(n5733), .A2(n5732), .ZN(n6103) );
  AOI211_X1 U6883 ( .C1(n6239), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n3952), 
        .B(n5734), .ZN(n5736) );
  AOI22_X1 U6884 ( .A1(n6149), .A2(REIP_REG_15__SCAN_IN), .B1(
        EBX_REG_15__SCAN_IN), .B2(n6264), .ZN(n5735) );
  OAI211_X1 U6885 ( .C1(n5920), .C2(n6258), .A(n5736), .B(n5735), .ZN(n5737)
         );
  AOI21_X1 U6886 ( .B1(n6103), .B2(n6155), .A(n5737), .ZN(n5738) );
  OAI21_X1 U6887 ( .B1(n5837), .B2(n6171), .A(n5738), .ZN(U2812) );
  NOR2_X1 U6888 ( .A1(n5740), .A2(n5739), .ZN(n5744) );
  OR2_X1 U6889 ( .A1(n5744), .A2(n6236), .ZN(n6174) );
  INV_X1 U6890 ( .A(n6174), .ZN(n5743) );
  INV_X1 U6891 ( .A(REIP_REG_11__SCAN_IN), .ZN(n5742) );
  OAI22_X1 U6892 ( .A1(n5743), .A2(n5742), .B1(n5741), .B2(n6258), .ZN(n5749)
         );
  AOI22_X1 U6893 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n6239), .B1(n5745), 
        .B2(n5744), .ZN(n5746) );
  OAI211_X1 U6894 ( .C1(n6180), .C2(n5747), .A(n5746), .B(n6434), .ZN(n5748)
         );
  AOI211_X1 U6895 ( .C1(n6363), .C2(n6155), .A(n5749), .B(n5748), .ZN(n5750)
         );
  OAI21_X1 U6896 ( .B1(n6171), .B2(n5751), .A(n5750), .ZN(U2816) );
  INV_X1 U6897 ( .A(n6255), .ZN(n6233) );
  NAND2_X1 U6898 ( .A1(n6196), .A2(n4546), .ZN(n5753) );
  NAND2_X1 U6899 ( .A1(n6239), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5752)
         );
  OAI211_X1 U6900 ( .C1(n5755), .C2(n5754), .A(n5753), .B(n5752), .ZN(n5756)
         );
  NOR2_X1 U6901 ( .A1(n5757), .A2(n5756), .ZN(n5759) );
  NAND2_X1 U6902 ( .A1(n6264), .A2(EBX_REG_1__SCAN_IN), .ZN(n5758) );
  OAI211_X1 U6903 ( .C1(n6417), .C2(n6257), .A(n5759), .B(n5758), .ZN(n5762)
         );
  NOR2_X1 U6904 ( .A1(n5760), .A2(n6260), .ZN(n5761) );
  AOI211_X1 U6905 ( .C1(n6233), .C2(n5763), .A(n5762), .B(n5761), .ZN(n5764)
         );
  INV_X1 U6906 ( .A(n5764), .ZN(U2826) );
  OAI222_X1 U6907 ( .A1(n5796), .A2(n5823), .B1(n5814), .B2(n6871), .C1(n5765), 
        .C2(n5808), .ZN(U2829) );
  AOI22_X1 U6908 ( .A1(n5929), .A2(n5811), .B1(n5805), .B2(EBX_REG_28__SCAN_IN), .ZN(n5766) );
  OAI21_X1 U6909 ( .B1(n5826), .B2(n5796), .A(n5766), .ZN(U2831) );
  INV_X1 U6910 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5767) );
  OAI222_X1 U6911 ( .A1(n5796), .A2(n5853), .B1(n5814), .B2(n5767), .C1(n5940), 
        .C2(n5808), .ZN(U2832) );
  OAI22_X1 U6912 ( .A1(n5952), .A2(n5808), .B1(n5768), .B2(n5814), .ZN(n5769)
         );
  INV_X1 U6913 ( .A(n5769), .ZN(n5770) );
  OAI21_X1 U6914 ( .B1(n6037), .B2(n5796), .A(n5770), .ZN(U2833) );
  INV_X1 U6915 ( .A(n5957), .ZN(n5771) );
  OAI222_X1 U6916 ( .A1(n5796), .A2(n5772), .B1(n5814), .B2(n5646), .C1(n5771), 
        .C2(n5808), .ZN(U2835) );
  OAI22_X1 U6917 ( .A1(n5964), .A2(n5808), .B1(n5773), .B2(n5814), .ZN(n5774)
         );
  INV_X1 U6918 ( .A(n5774), .ZN(n5775) );
  OAI21_X1 U6919 ( .B1(n5829), .B2(n5796), .A(n5775), .ZN(U2836) );
  OAI222_X1 U6920 ( .A1(n5776), .A2(n5814), .B1(n5796), .B2(n5883), .C1(n5808), 
        .C2(n5975), .ZN(U2837) );
  INV_X1 U6921 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5777) );
  OAI222_X1 U6922 ( .A1(n5777), .A2(n5814), .B1(n5808), .B2(n5982), .C1(n6047), 
        .C2(n5796), .ZN(U2838) );
  AND2_X1 U6923 ( .A1(n5785), .A2(n5778), .ZN(n5779) );
  OR2_X1 U6924 ( .A1(n5779), .A2(n5667), .ZN(n6017) );
  MUX2_X1 U6925 ( .A(n5781), .B(n5780), .S(n5789), .Z(n5783) );
  XNOR2_X1 U6926 ( .A(n5783), .B(n5782), .ZN(n6022) );
  OAI222_X1 U6927 ( .A1(n5796), .A2(n6017), .B1(n5808), .B2(n6022), .C1(n5784), 
        .C2(n5814), .ZN(U2839) );
  OAI21_X1 U6928 ( .B1(n5786), .B2(n3160), .A(n5785), .ZN(n6031) );
  NAND2_X1 U6929 ( .A1(n5788), .A2(n5787), .ZN(n5801) );
  INV_X1 U6930 ( .A(n5801), .ZN(n5791) );
  OR2_X1 U6931 ( .A1(n5789), .A2(n5791), .ZN(n5793) );
  OAI21_X1 U6932 ( .B1(n5802), .B2(n5791), .A(n5790), .ZN(n5792) );
  NAND2_X1 U6933 ( .A1(n5793), .A2(n5792), .ZN(n6030) );
  OAI22_X1 U6934 ( .A1(n6030), .A2(n5808), .B1(n6957), .B2(n5814), .ZN(n5794)
         );
  INV_X1 U6935 ( .A(n5794), .ZN(n5795) );
  OAI21_X1 U6936 ( .B1(n6031), .B2(n5796), .A(n5795), .ZN(U2840) );
  OR2_X1 U6937 ( .A1(n5798), .A2(n5797), .ZN(n5800) );
  AND2_X1 U6938 ( .A1(n5800), .A2(n5799), .ZN(n6268) );
  INV_X1 U6939 ( .A(n6268), .ZN(n5804) );
  XNOR2_X1 U6940 ( .A(n5802), .B(n5801), .ZN(n6140) );
  AOI22_X1 U6941 ( .A1(n6140), .A2(n5811), .B1(EBX_REG_18__SCAN_IN), .B2(n5805), .ZN(n5803) );
  OAI21_X1 U6942 ( .B1(n5804), .B2(n5796), .A(n5803), .ZN(U2841) );
  AOI22_X1 U6943 ( .A1(n6086), .A2(n5811), .B1(n5805), .B2(EBX_REG_17__SCAN_IN), .ZN(n5806) );
  OAI21_X1 U6944 ( .B1(n5835), .B2(n5796), .A(n5806), .ZN(U2842) );
  OAI222_X1 U6945 ( .A1(n5809), .A2(n5814), .B1(n5808), .B2(n6095), .C1(n5807), 
        .C2(n5796), .ZN(U2843) );
  INV_X1 U6946 ( .A(EBX_REG_15__SCAN_IN), .ZN(n7035) );
  NAND2_X1 U6947 ( .A1(n5922), .A2(n5810), .ZN(n5813) );
  NAND2_X1 U6948 ( .A1(n6103), .A2(n5811), .ZN(n5812) );
  OAI211_X1 U6949 ( .C1(n7035), .C2(n5814), .A(n5813), .B(n5812), .ZN(U2844)
         );
  AND2_X1 U6950 ( .A1(n5816), .A2(n5815), .ZN(n5817) );
  NAND2_X1 U6951 ( .A1(n5818), .A2(n5817), .ZN(n5820) );
  AOI22_X1 U6952 ( .A1(n6271), .A2(DATAI_31_), .B1(n6743), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5819) );
  NAND2_X1 U6953 ( .A1(n5820), .A2(n5819), .ZN(U2860) );
  AOI22_X1 U6954 ( .A1(n6271), .A2(DATAI_30_), .B1(n6743), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5822) );
  NAND2_X1 U6955 ( .A1(n6273), .A2(DATAI_14_), .ZN(n5821) );
  OAI211_X1 U6956 ( .C1(n5823), .C2(n5834), .A(n5822), .B(n5821), .ZN(U2861)
         );
  AOI22_X1 U6957 ( .A1(n6271), .A2(DATAI_28_), .B1(n6743), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5825) );
  NAND2_X1 U6958 ( .A1(n6273), .A2(DATAI_12_), .ZN(n5824) );
  OAI211_X1 U6959 ( .C1(n5826), .C2(n5834), .A(n5825), .B(n5824), .ZN(U2863)
         );
  AOI22_X1 U6960 ( .A1(n6271), .A2(DATAI_23_), .B1(n6743), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5828) );
  NAND2_X1 U6961 ( .A1(n6273), .A2(DATAI_7_), .ZN(n5827) );
  OAI211_X1 U6962 ( .C1(n5829), .C2(n5834), .A(n5828), .B(n5827), .ZN(U2868)
         );
  AOI22_X1 U6963 ( .A1(n6273), .A2(DATAI_3_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n6743), .ZN(n5831) );
  NAND2_X1 U6964 ( .A1(n6271), .A2(DATAI_19_), .ZN(n5830) );
  OAI211_X1 U6965 ( .C1(n6031), .C2(n5834), .A(n5831), .B(n5830), .ZN(U2872)
         );
  AOI22_X1 U6966 ( .A1(n6271), .A2(DATAI_17_), .B1(n6743), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U6967 ( .A1(n6273), .A2(DATAI_1_), .ZN(n5832) );
  OAI211_X1 U6968 ( .C1(n5835), .C2(n5834), .A(n5833), .B(n5832), .ZN(U2874)
         );
  AOI22_X1 U6969 ( .A1(n6742), .A2(DATAI_15_), .B1(n6743), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5836) );
  OAI21_X1 U6970 ( .B1(n5837), .B2(n5834), .A(n5836), .ZN(U2876) );
  NAND3_X1 U6971 ( .A1(n4442), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5880), .ZN(n5842) );
  INV_X1 U6972 ( .A(n5838), .ZN(n5840) );
  NAND2_X1 U6973 ( .A1(n6073), .A2(n5841), .ZN(n5948) );
  NOR2_X1 U6974 ( .A1(n5880), .A2(n5948), .ZN(n5839) );
  NAND2_X1 U6975 ( .A1(n5840), .A2(n5839), .ZN(n5849) );
  AOI22_X1 U6976 ( .A1(n5842), .A2(n5849), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5841), .ZN(n5843) );
  XNOR2_X1 U6977 ( .A(n5843), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5938)
         );
  NAND2_X1 U6978 ( .A1(n3952), .A2(REIP_REG_28__SCAN_IN), .ZN(n5934) );
  NAND2_X1 U6979 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5844)
         );
  OAI211_X1 U6980 ( .C1(n6352), .C2(n5845), .A(n5934), .B(n5844), .ZN(n5846)
         );
  AOI21_X1 U6981 ( .B1(n5847), .B2(n6347), .A(n5846), .ZN(n5848) );
  OAI21_X1 U6982 ( .B1(n6355), .B2(n5938), .A(n5848), .ZN(U2958) );
  NAND2_X1 U6983 ( .A1(n5850), .A2(n5849), .ZN(n5851) );
  XNOR2_X1 U6984 ( .A(n5851), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5946)
         );
  NAND2_X1 U6985 ( .A1(n3952), .A2(REIP_REG_27__SCAN_IN), .ZN(n5939) );
  OAI21_X1 U6986 ( .B1(n6342), .B2(n5852), .A(n5939), .ZN(n5855) );
  NOR2_X1 U6987 ( .A1(n5853), .A2(n6361), .ZN(n5854) );
  OAI21_X1 U6988 ( .B1(n5946), .B2(n6355), .A(n5857), .ZN(U2959) );
  NOR2_X1 U6989 ( .A1(n5880), .A2(n6897), .ZN(n5859) );
  OR2_X1 U6990 ( .A1(n5897), .A2(n5859), .ZN(n5861) );
  NAND2_X1 U6991 ( .A1(n5880), .A2(n6897), .ZN(n5860) );
  INV_X1 U6992 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n7011) );
  NAND2_X1 U6993 ( .A1(n5880), .A2(n7011), .ZN(n5863) );
  NOR2_X1 U6994 ( .A1(n5989), .A2(n7011), .ZN(n5862) );
  XNOR2_X1 U6995 ( .A(n5880), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5890)
         );
  INV_X1 U6996 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5971) );
  NAND3_X1 U6997 ( .A1(n5865), .A2(n5864), .A3(n5971), .ZN(n5872) );
  NAND3_X1 U6998 ( .A1(n5989), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5866) );
  INV_X1 U6999 ( .A(n5865), .ZN(n5888) );
  OAI21_X1 U7000 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5864), .A(n5888), 
        .ZN(n5882) );
  AOI22_X1 U7001 ( .A1(n5872), .A2(n5866), .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5882), .ZN(n5867) );
  XNOR2_X1 U7002 ( .A(n5867), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5961)
         );
  NOR2_X1 U7003 ( .A1(n6434), .A2(n6677), .ZN(n5956) );
  AOI21_X1 U7004 ( .B1(n6358), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5956), 
        .ZN(n5868) );
  OAI21_X1 U7005 ( .B1(n5869), .B2(n6352), .A(n5868), .ZN(n5870) );
  AOI21_X1 U7006 ( .B1(n6041), .B2(n6347), .A(n5870), .ZN(n5871) );
  OAI21_X1 U7007 ( .B1(n5961), .B2(n6355), .A(n5871), .ZN(U2962) );
  XNOR2_X1 U7008 ( .A(n5989), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5896)
         );
  NAND2_X1 U7009 ( .A1(n5897), .A2(n5896), .ZN(n5999) );
  OAI21_X1 U7010 ( .B1(n5873), .B2(n5999), .A(n5872), .ZN(n5874) );
  XNOR2_X1 U7011 ( .A(n5874), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5970)
         );
  NAND2_X1 U7012 ( .A1(n3952), .A2(REIP_REG_23__SCAN_IN), .ZN(n5963) );
  NAND2_X1 U7013 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5875)
         );
  OAI211_X1 U7014 ( .C1(n6352), .C2(n5876), .A(n5963), .B(n5875), .ZN(n5877)
         );
  AOI21_X1 U7015 ( .B1(n5878), .B2(n6347), .A(n5877), .ZN(n5879) );
  OAI21_X1 U7016 ( .B1(n5970), .B2(n6355), .A(n5879), .ZN(U2963) );
  XNOR2_X1 U7017 ( .A(n5880), .B(n5971), .ZN(n5881) );
  XNOR2_X1 U7018 ( .A(n5882), .B(n5881), .ZN(n5978) );
  INV_X1 U7019 ( .A(n5883), .ZN(n6044) );
  NAND2_X1 U7020 ( .A1(n3952), .A2(REIP_REG_22__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U7021 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5884)
         );
  OAI211_X1 U7022 ( .C1(n6352), .C2(n5885), .A(n5973), .B(n5884), .ZN(n5886)
         );
  AOI21_X1 U7023 ( .B1(n6044), .B2(n6347), .A(n5886), .ZN(n5887) );
  OAI21_X1 U7024 ( .B1(n5978), .B2(n6355), .A(n5887), .ZN(U2964) );
  OAI21_X1 U7025 ( .B1(n5890), .B2(n5889), .A(n5888), .ZN(n5980) );
  NAND2_X1 U7026 ( .A1(n5980), .A2(n4310), .ZN(n5895) );
  NAND2_X1 U7027 ( .A1(n3952), .A2(REIP_REG_21__SCAN_IN), .ZN(n5981) );
  OAI21_X1 U7028 ( .B1(n6342), .B2(n5891), .A(n5981), .ZN(n5892) );
  AOI21_X1 U7029 ( .B1(n6336), .B2(n5893), .A(n5892), .ZN(n5894) );
  OAI211_X1 U7030 ( .C1(n6361), .C2(n6047), .A(n5895), .B(n5894), .ZN(U2965)
         );
  OR2_X1 U7031 ( .A1(n5897), .A2(n5896), .ZN(n6000) );
  NAND3_X1 U7032 ( .A1(n6000), .A2(n5999), .A3(n4310), .ZN(n5901) );
  NAND2_X1 U7033 ( .A1(n3952), .A2(REIP_REG_19__SCAN_IN), .ZN(n6004) );
  OAI21_X1 U7034 ( .B1(n6342), .B2(n5898), .A(n6004), .ZN(n5899) );
  AOI21_X1 U7035 ( .B1(n6336), .B2(n6028), .A(n5899), .ZN(n5900) );
  OAI211_X1 U7036 ( .C1(n6361), .C2(n6031), .A(n5901), .B(n5900), .ZN(U2967)
         );
  NOR2_X1 U7037 ( .A1(n6061), .A2(n6100), .ZN(n5904) );
  NOR2_X1 U7038 ( .A1(n5916), .A2(n5989), .ZN(n6064) );
  OAI22_X1 U7039 ( .A1(n5904), .A2(n6064), .B1(n5989), .B2(n6100), .ZN(n5905)
         );
  XOR2_X1 U7040 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .B(n5905), .Z(n6083) );
  AOI22_X1 U7041 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .B1(n3952), 
        .B2(REIP_REG_17__SCAN_IN), .ZN(n5906) );
  OAI21_X1 U7042 ( .B1(n5907), .B2(n6352), .A(n5906), .ZN(n5908) );
  AOI21_X1 U7043 ( .B1(n5909), .B2(n6347), .A(n5908), .ZN(n5910) );
  OAI21_X1 U7044 ( .B1(n6083), .B2(n6355), .A(n5910), .ZN(U2969) );
  XNOR2_X1 U7045 ( .A(n5864), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5911)
         );
  XNOR2_X1 U7046 ( .A(n6061), .B(n5911), .ZN(n6096) );
  AOI22_X1 U7047 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n3952), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5912) );
  OAI21_X1 U7048 ( .B1(n5913), .B2(n6352), .A(n5912), .ZN(n5914) );
  AOI21_X1 U7049 ( .B1(n6272), .B2(n6347), .A(n5914), .ZN(n5915) );
  OAI21_X1 U7050 ( .B1(n6096), .B2(n6355), .A(n5915), .ZN(U2970) );
  OAI21_X1 U7051 ( .B1(n5918), .B2(n5917), .A(n5916), .ZN(n6104) );
  INV_X1 U7052 ( .A(n6104), .ZN(n5924) );
  AOI22_X1 U7053 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n3952), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5919) );
  OAI21_X1 U7054 ( .B1(n5920), .B2(n6352), .A(n5919), .ZN(n5921) );
  AOI21_X1 U7055 ( .B1(n5922), .B2(n6347), .A(n5921), .ZN(n5923) );
  OAI21_X1 U7056 ( .B1(n5924), .B2(n6355), .A(n5923), .ZN(U2971) );
  OAI22_X1 U7057 ( .A1(n6342), .A2(n6835), .B1(n6434), .B2(n6659), .ZN(n5926)
         );
  NOR2_X1 U7058 ( .A1(n6147), .A2(n6361), .ZN(n5925) );
  AOI211_X1 U7059 ( .C1(n6336), .C2(n6148), .A(n5926), .B(n5925), .ZN(n5927)
         );
  OAI21_X1 U7060 ( .B1(n5928), .B2(n6355), .A(n5927), .ZN(U2972) );
  INV_X1 U7061 ( .A(n5929), .ZN(n5935) );
  INV_X1 U7062 ( .A(n5941), .ZN(n5932) );
  NAND3_X1 U7063 ( .A1(n5932), .A2(n5931), .A3(n5930), .ZN(n5933) );
  OAI211_X1 U7064 ( .C1(n5935), .C2(n6424), .A(n5934), .B(n5933), .ZN(n5936)
         );
  AOI21_X1 U7065 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n5944), .A(n5936), 
        .ZN(n5937) );
  OAI21_X1 U7066 ( .B1(n5938), .B2(n6425), .A(n5937), .ZN(U2990) );
  OAI21_X1 U7067 ( .B1(n5940), .B2(n6424), .A(n5939), .ZN(n5943) );
  NOR2_X1 U7068 ( .A1(n5941), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5942)
         );
  AOI211_X1 U7069 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5944), .A(n5943), .B(n5942), .ZN(n5945) );
  OAI21_X1 U7070 ( .B1(n5946), .B2(n6425), .A(n5945), .ZN(U2991) );
  INV_X1 U7071 ( .A(n5947), .ZN(n5949) );
  NAND3_X1 U7072 ( .A1(n6074), .A2(n5949), .A3(n5948), .ZN(n5951) );
  OAI211_X1 U7073 ( .C1(n6424), .C2(n5952), .A(n5951), .B(n5950), .ZN(n5953)
         );
  AOI21_X1 U7074 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n6072), .A(n5953), 
        .ZN(n5954) );
  OAI21_X1 U7075 ( .B1(n5955), .B2(n6425), .A(n5954), .ZN(U2992) );
  AOI21_X1 U7076 ( .B1(n5957), .B2(n6390), .A(n5956), .ZN(n5960) );
  INV_X1 U7077 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n7031) );
  NOR2_X1 U7078 ( .A1(n5965), .A2(n7031), .ZN(n5958) );
  OAI21_X1 U7079 ( .B1(n5958), .B2(INSTADDRPOINTER_REG_24__SCAN_IN), .A(n6072), 
        .ZN(n5959) );
  OAI211_X1 U7080 ( .C1(n5961), .C2(n6425), .A(n5960), .B(n5959), .ZN(U2994)
         );
  INV_X1 U7081 ( .A(n5962), .ZN(n5968) );
  OAI21_X1 U7082 ( .B1(n5964), .B2(n6424), .A(n5963), .ZN(n5967) );
  NOR2_X1 U7083 ( .A1(n5965), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5966)
         );
  AOI211_X1 U7084 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5968), .A(n5967), .B(n5966), .ZN(n5969) );
  OAI21_X1 U7085 ( .B1(n5970), .B2(n6425), .A(n5969), .ZN(U2995) );
  XNOR2_X1 U7086 ( .A(n5971), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5972)
         );
  NAND2_X1 U7087 ( .A1(n5984), .A2(n5972), .ZN(n5974) );
  OAI211_X1 U7088 ( .C1(n6424), .C2(n5975), .A(n5974), .B(n5973), .ZN(n5976)
         );
  AOI21_X1 U7089 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5979), .A(n5976), 
        .ZN(n5977) );
  OAI21_X1 U7090 ( .B1(n5978), .B2(n6425), .A(n5977), .ZN(U2996) );
  INV_X1 U7091 ( .A(n5979), .ZN(n5988) );
  NAND2_X1 U7092 ( .A1(n5980), .A2(n6420), .ZN(n5986) );
  OAI21_X1 U7093 ( .B1(n5982), .B2(n6424), .A(n5981), .ZN(n5983) );
  AOI21_X1 U7094 ( .B1(n5984), .B2(n5987), .A(n5983), .ZN(n5985) );
  OAI211_X1 U7095 ( .C1(n5988), .C2(n5987), .A(n5986), .B(n5985), .ZN(U2997)
         );
  XNOR2_X1 U7096 ( .A(n5989), .B(n7011), .ZN(n5990) );
  XNOR2_X1 U7097 ( .A(n5991), .B(n5990), .ZN(n6055) );
  INV_X1 U7098 ( .A(n6055), .ZN(n5998) );
  NOR2_X1 U7099 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5992), .ZN(n6085)
         );
  NOR2_X1 U7100 ( .A1(n6085), .A2(n6087), .ZN(n6082) );
  OAI21_X1 U7101 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n6414), .A(n6082), 
        .ZN(n6006) );
  AOI21_X1 U7102 ( .B1(n7011), .B2(n6897), .A(n6001), .ZN(n5994) );
  AOI22_X1 U7103 ( .A1(n3952), .A2(REIP_REG_20__SCAN_IN), .B1(n5994), .B2(
        n5993), .ZN(n5995) );
  OAI21_X1 U7104 ( .B1(n6022), .B2(n6424), .A(n5995), .ZN(n5996) );
  AOI21_X1 U7105 ( .B1(n6006), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5996), 
        .ZN(n5997) );
  OAI21_X1 U7106 ( .B1(n5998), .B2(n6425), .A(n5997), .ZN(U2998) );
  NAND3_X1 U7107 ( .A1(n6000), .A2(n5999), .A3(n6420), .ZN(n6008) );
  INV_X1 U7108 ( .A(n6001), .ZN(n6002) );
  NAND2_X1 U7109 ( .A1(n6897), .A2(n6002), .ZN(n6003) );
  OAI211_X1 U7110 ( .C1(n6030), .C2(n6424), .A(n6004), .B(n6003), .ZN(n6005)
         );
  AOI21_X1 U7111 ( .B1(n6006), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n6005), 
        .ZN(n6007) );
  NAND2_X1 U7112 ( .A1(n6008), .A2(n6007), .ZN(U2999) );
  OAI211_X1 U7113 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n4640), .A(n6505), .B(
        n6442), .ZN(n6009) );
  OAI21_X1 U7114 ( .B1(n6013), .B2(n6010), .A(n6009), .ZN(n6011) );
  MUX2_X1 U7115 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n6011), .S(n6435), 
        .Z(U3464) );
  XNOR2_X1 U7116 ( .A(n6012), .B(n6505), .ZN(n6015) );
  OAI22_X1 U7117 ( .A1(n6015), .A2(n6729), .B1(n6014), .B2(n6013), .ZN(n6016)
         );
  MUX2_X1 U7118 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n6016), .S(n6435), 
        .Z(U3463) );
  INV_X1 U7119 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n6888) );
  NOR2_X1 U7120 ( .A1(n6888), .A2(n6301), .ZN(U2892) );
  AOI22_X1 U7121 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6264), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6239), .ZN(n6025) );
  INV_X1 U7122 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6668) );
  INV_X1 U7123 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6666) );
  NOR2_X1 U7124 ( .A1(n6668), .A2(n6666), .ZN(n6019) );
  AOI21_X1 U7125 ( .B1(n6027), .B2(n6019), .A(REIP_REG_20__SCAN_IN), .ZN(n6021) );
  OAI22_X1 U7126 ( .A1(n6022), .A2(n6257), .B1(n6021), .B2(n6020), .ZN(n6023)
         );
  AOI21_X1 U7127 ( .B1(n6054), .B2(n6220), .A(n6023), .ZN(n6024) );
  OAI211_X1 U7128 ( .C1(n6058), .C2(n6258), .A(n6025), .B(n6024), .ZN(U2807)
         );
  NAND2_X1 U7129 ( .A1(n6027), .A2(n6666), .ZN(n6142) );
  NOR2_X1 U7130 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6666), .ZN(n6026) );
  AOI22_X1 U7131 ( .A1(n6028), .A2(n6196), .B1(n6027), .B2(n6026), .ZN(n6029)
         );
  OAI211_X1 U7132 ( .C1(n6253), .C2(n5898), .A(n6029), .B(n6434), .ZN(n6033)
         );
  OAI22_X1 U7133 ( .A1(n6031), .A2(n6171), .B1(n6257), .B2(n6030), .ZN(n6032)
         );
  AOI211_X1 U7134 ( .C1(EBX_REG_19__SCAN_IN), .C2(n6264), .A(n6033), .B(n6032), 
        .ZN(n6034) );
  OAI221_X1 U7135 ( .B1(n6668), .B2(n6137), .C1(n6668), .C2(n6142), .A(n6034), 
        .ZN(U2808) );
  INV_X1 U7136 ( .A(n6271), .ZN(n6036) );
  OAI22_X1 U7137 ( .A1(n6037), .A2(n5834), .B1(n6036), .B2(n6035), .ZN(n6038)
         );
  INV_X1 U7138 ( .A(n6038), .ZN(n6040) );
  AOI22_X1 U7139 ( .A1(n6273), .A2(DATAI_10_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6743), .ZN(n6039) );
  NAND2_X1 U7140 ( .A1(n6040), .A2(n6039), .ZN(U2865) );
  AOI22_X1 U7141 ( .A1(n6041), .A2(n6744), .B1(n6271), .B2(DATAI_24_), .ZN(
        n6043) );
  AOI22_X1 U7142 ( .A1(n6273), .A2(DATAI_8_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6743), .ZN(n6042) );
  NAND2_X1 U7143 ( .A1(n6043), .A2(n6042), .ZN(U2867) );
  AOI22_X1 U7144 ( .A1(n6044), .A2(n6744), .B1(n6271), .B2(DATAI_22_), .ZN(
        n6046) );
  AOI22_X1 U7145 ( .A1(n6273), .A2(DATAI_6_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n6743), .ZN(n6045) );
  NAND2_X1 U7146 ( .A1(n6046), .A2(n6045), .ZN(U2869) );
  OR2_X1 U7147 ( .A1(n6047), .A2(n5834), .ZN(n6049) );
  NAND2_X1 U7148 ( .A1(n6271), .A2(DATAI_21_), .ZN(n6048) );
  AND2_X1 U7149 ( .A1(n6049), .A2(n6048), .ZN(n6051) );
  AOI22_X1 U7150 ( .A1(n6273), .A2(DATAI_5_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n6743), .ZN(n6050) );
  NAND2_X1 U7151 ( .A1(n6051), .A2(n6050), .ZN(U2870) );
  AOI22_X1 U7152 ( .A1(n6054), .A2(n6744), .B1(n6271), .B2(DATAI_20_), .ZN(
        n6053) );
  AOI22_X1 U7153 ( .A1(n6273), .A2(DATAI_4_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n6743), .ZN(n6052) );
  NAND2_X1 U7154 ( .A1(n6053), .A2(n6052), .ZN(U2871) );
  AOI22_X1 U7155 ( .A1(n3952), .A2(REIP_REG_20__SCAN_IN), .B1(n6358), .B2(
        PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6057) );
  AOI22_X1 U7156 ( .A1(n6055), .A2(n4310), .B1(n6347), .B2(n6054), .ZN(n6056)
         );
  OAI211_X1 U7157 ( .C1(n6352), .C2(n6058), .A(n6057), .B(n6056), .ZN(U2966)
         );
  AOI22_X1 U7158 ( .A1(n3952), .A2(REIP_REG_18__SCAN_IN), .B1(n6358), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6067) );
  NOR2_X1 U7159 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6063) );
  INV_X1 U7160 ( .A(n6059), .ZN(n6060) );
  NOR3_X1 U7161 ( .A1(n6061), .A2(n5864), .A3(n6060), .ZN(n6062) );
  AOI21_X1 U7162 ( .B1(n6064), .B2(n6063), .A(n6062), .ZN(n6065) );
  XNOR2_X1 U7163 ( .A(n6065), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6078)
         );
  AOI22_X1 U7164 ( .A1(n6078), .A2(n4310), .B1(n6347), .B2(n6268), .ZN(n6066)
         );
  OAI211_X1 U7165 ( .C1(n6352), .C2(n6138), .A(n6067), .B(n6066), .ZN(U2968)
         );
  INV_X1 U7166 ( .A(n6068), .ZN(n6069) );
  AOI22_X1 U7167 ( .A1(n6070), .A2(n6420), .B1(n6390), .B2(n6069), .ZN(n6076)
         );
  NOR2_X1 U7168 ( .A1(n6434), .A2(n6846), .ZN(n6071) );
  AOI221_X1 U7169 ( .B1(n6074), .B2(n6073), .C1(n6072), .C2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A(n6071), .ZN(n6075) );
  NAND2_X1 U7170 ( .A1(n6076), .A2(n6075), .ZN(U2993) );
  INV_X1 U7171 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6081) );
  AOI22_X1 U7172 ( .A1(REIP_REG_18__SCAN_IN), .A2(n3952), .B1(n6077), .B2(
        n6081), .ZN(n6080) );
  AOI22_X1 U7173 ( .A1(n6078), .A2(n6420), .B1(n6390), .B2(n6140), .ZN(n6079)
         );
  OAI211_X1 U7174 ( .C1(n6082), .C2(n6081), .A(n6080), .B(n6079), .ZN(U3000)
         );
  NOR2_X1 U7175 ( .A1(n6083), .A2(n6425), .ZN(n6084) );
  AOI211_X1 U7176 ( .C1(n3952), .C2(REIP_REG_17__SCAN_IN), .A(n6085), .B(n6084), .ZN(n6089) );
  AOI22_X1 U7177 ( .A1(n6087), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .B1(n6390), .B2(n6086), .ZN(n6088) );
  NAND2_X1 U7178 ( .A1(n6089), .A2(n6088), .ZN(U3001) );
  INV_X1 U7179 ( .A(n6092), .ZN(n6091) );
  AOI21_X1 U7180 ( .B1(n6091), .B2(n6090), .A(n6367), .ZN(n6101) );
  NAND3_X1 U7181 ( .A1(n6092), .A2(n7010), .A3(n6366), .ZN(n6105) );
  NOR3_X1 U7182 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n6094), .A3(n6093), 
        .ZN(n6098) );
  OAI22_X1 U7183 ( .A1(n6096), .A2(n6425), .B1(n6424), .B2(n6095), .ZN(n6097)
         );
  AOI211_X1 U7184 ( .C1(REIP_REG_16__SCAN_IN), .C2(n3952), .A(n6098), .B(n6097), .ZN(n6099) );
  OAI221_X1 U7185 ( .B1(n6100), .B2(n6101), .C1(n6100), .C2(n6105), .A(n6099), 
        .ZN(U3002) );
  INV_X1 U7186 ( .A(REIP_REG_15__SCAN_IN), .ZN(n7002) );
  INV_X1 U7187 ( .A(n6101), .ZN(n6102) );
  AOI222_X1 U7188 ( .A1(n6104), .A2(n6420), .B1(n6390), .B2(n6103), .C1(n6102), 
        .C2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6106) );
  OAI211_X1 U7189 ( .C1(n7002), .C2(n6434), .A(n6106), .B(n6105), .ZN(U3003)
         );
  INV_X1 U7190 ( .A(n6107), .ZN(n6111) );
  INV_X1 U7191 ( .A(n6108), .ZN(n6110) );
  NAND4_X1 U7192 ( .A1(n6111), .A2(n6110), .A3(n6109), .A4(n6234), .ZN(n6112)
         );
  OAI21_X1 U7193 ( .B1(n6713), .B2(n6113), .A(n6112), .ZN(U3455) );
  AOI21_X1 U7194 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6975), .A(n6628), .ZN(n6119) );
  INV_X1 U7195 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6114) );
  NOR2_X2 U7196 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6974), .ZN(n6741) );
  AOI21_X1 U7197 ( .B1(n6119), .B2(n6114), .A(n6741), .ZN(U2789) );
  INV_X1 U7198 ( .A(n6115), .ZN(n6116) );
  OAI21_X1 U7199 ( .B1(n6116), .B2(n6612), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6117) );
  OAI21_X1 U7200 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6611), .A(n6117), .ZN(
        U2790) );
  NOR2_X1 U7201 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n6120) );
  OAI21_X1 U7202 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6120), .A(n6727), .ZN(n6118)
         );
  OAI21_X1 U7203 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6727), .A(n6118), .ZN(
        U2791) );
  NOR2_X2 U7204 ( .A1(n6741), .A2(n6119), .ZN(n6697) );
  OAI21_X1 U7205 ( .B1(n6120), .B2(BS16_N), .A(n6697), .ZN(n6696) );
  OAI21_X1 U7206 ( .B1(n6697), .B2(n6121), .A(n6696), .ZN(U2792) );
  OAI21_X1 U7207 ( .B1(n6123), .B2(n6122), .A(n6355), .ZN(U2793) );
  INV_X1 U7208 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6959) );
  INV_X1 U7209 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6920) );
  INV_X1 U7210 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6917) );
  INV_X1 U7211 ( .A(DATAWIDTH_REG_31__SCAN_IN), .ZN(n6803) );
  NAND4_X1 U7212 ( .A1(n6959), .A2(n6920), .A3(n6917), .A4(n6803), .ZN(n6124)
         );
  AOI211_X1 U7213 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_13__SCAN_IN), .B(n6124), 
        .ZN(n6133) );
  NOR4_X1 U7214 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n6132) );
  NOR4_X1 U7215 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6131) );
  NOR4_X1 U7216 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6125) );
  INV_X1 U7217 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n6863) );
  NAND2_X1 U7218 ( .A1(n6125), .A2(n6863), .ZN(n7030) );
  NOR4_X1 U7219 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_4__SCAN_IN), .A4(
        DATAWIDTH_REG_5__SCAN_IN), .ZN(n6128) );
  NOR4_X1 U7220 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n6127) );
  NOR4_X1 U7221 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_10__SCAN_IN), .ZN(n6126) );
  NAND3_X1 U7222 ( .A1(n6128), .A2(n6127), .A3(n6126), .ZN(n6129) );
  NOR2_X1 U7223 ( .A1(n7030), .A2(n6129), .ZN(n6130) );
  NAND4_X1 U7224 ( .A1(n6133), .A2(n6132), .A3(n6131), .A4(n6130), .ZN(n6723)
         );
  NOR2_X1 U7225 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6723), .ZN(n6725) );
  INV_X1 U7226 ( .A(n6723), .ZN(n6720) );
  NOR2_X1 U7227 ( .A1(n6720), .A2(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6134) );
  INV_X1 U7228 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6717) );
  INV_X1 U7229 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6718) );
  NAND4_X1 U7230 ( .A1(n6720), .A2(n6724), .A3(n6717), .A4(n6718), .ZN(n6135)
         );
  OAI21_X1 U7231 ( .B1(n6725), .B2(n6134), .A(n6135), .ZN(U2794) );
  AOI22_X1 U7232 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(n6723), .B1(n6725), 
        .B2(n6717), .ZN(n6136) );
  NAND2_X1 U7233 ( .A1(n6136), .A2(n6135), .ZN(U2795) );
  OAI22_X1 U7234 ( .A1(n6138), .A2(n6258), .B1(n6666), .B2(n6137), .ZN(n6139)
         );
  AOI211_X1 U7235 ( .C1(n6239), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n3952), 
        .B(n6139), .ZN(n6144) );
  AOI22_X1 U7236 ( .A1(n6268), .A2(n6220), .B1(n6155), .B2(n6140), .ZN(n6143)
         );
  NAND2_X1 U7237 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6264), .ZN(n6141) );
  NAND4_X1 U7238 ( .A1(n6144), .A2(n6143), .A3(n6142), .A4(n6141), .ZN(U2809)
         );
  AOI22_X1 U7239 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6264), .B1(
        PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n6239), .ZN(n6153) );
  INV_X1 U7240 ( .A(n6145), .ZN(n6146) );
  AOI21_X1 U7241 ( .B1(n6146), .B2(n6155), .A(n3952), .ZN(n6152) );
  INV_X1 U7242 ( .A(n6147), .ZN(n6745) );
  AOI22_X1 U7243 ( .A1(n6745), .A2(n6220), .B1(n6196), .B2(n6148), .ZN(n6151)
         );
  NOR2_X1 U7244 ( .A1(n6157), .A2(n6808), .ZN(n6154) );
  OAI221_X1 U7245 ( .B1(REIP_REG_14__SCAN_IN), .B2(REIP_REG_13__SCAN_IN), .C1(
        REIP_REG_14__SCAN_IN), .C2(n6154), .A(n6149), .ZN(n6150) );
  NAND4_X1 U7246 ( .A1(n6153), .A2(n6152), .A3(n6151), .A4(n6150), .ZN(U2813)
         );
  AOI22_X1 U7247 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6264), .B1(n6154), .B2(n6657), .ZN(n6164) );
  AOI22_X1 U7248 ( .A1(n6156), .A2(n6155), .B1(PHYADDRPOINTER_REG_13__SCAN_IN), 
        .B2(n6239), .ZN(n6163) );
  NOR2_X1 U7249 ( .A1(n6157), .A2(REIP_REG_12__SCAN_IN), .ZN(n6168) );
  AOI221_X1 U7250 ( .B1(n6168), .B2(REIP_REG_13__SCAN_IN), .C1(n6174), .C2(
        REIP_REG_13__SCAN_IN), .A(n3952), .ZN(n6162) );
  OAI22_X1 U7251 ( .A1(n6159), .A2(n6171), .B1(n6158), .B2(n6258), .ZN(n6160)
         );
  INV_X1 U7252 ( .A(n6160), .ZN(n6161) );
  NAND4_X1 U7253 ( .A1(n6164), .A2(n6163), .A3(n6162), .A4(n6161), .ZN(U2814)
         );
  OAI22_X1 U7254 ( .A1(n6166), .A2(n6257), .B1(n6180), .B2(n6165), .ZN(n6167)
         );
  INV_X1 U7255 ( .A(n6167), .ZN(n6178) );
  AOI211_X1 U7256 ( .C1(n6239), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n3952), 
        .B(n6168), .ZN(n6177) );
  INV_X1 U7257 ( .A(n6169), .ZN(n6170) );
  OAI22_X1 U7258 ( .A1(n6172), .A2(n6171), .B1(n6170), .B2(n6258), .ZN(n6173)
         );
  INV_X1 U7259 ( .A(n6173), .ZN(n6176) );
  NAND2_X1 U7260 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6174), .ZN(n6175) );
  NAND4_X1 U7261 ( .A1(n6178), .A2(n6177), .A3(n6176), .A4(n6175), .ZN(U2815)
         );
  OAI22_X1 U7262 ( .A1(n6181), .A2(n6257), .B1(n6180), .B2(n6179), .ZN(n6182)
         );
  INV_X1 U7263 ( .A(n6182), .ZN(n6191) );
  AOI21_X1 U7264 ( .B1(n6200), .B2(n6183), .A(n6653), .ZN(n6186) );
  INV_X1 U7265 ( .A(n6206), .ZN(n6192) );
  NOR3_X1 U7266 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6184), .A3(n6192), .ZN(n6185) );
  AOI211_X1 U7267 ( .C1(n6239), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6186), 
        .B(n6185), .ZN(n6190) );
  AOI22_X1 U7268 ( .A1(n6188), .A2(n6220), .B1(n6196), .B2(n6187), .ZN(n6189)
         );
  NAND4_X1 U7269 ( .A1(n6191), .A2(n6190), .A3(n6189), .A4(n6434), .ZN(U2817)
         );
  NOR2_X1 U7270 ( .A1(n6645), .A2(n6192), .ZN(n6202) );
  AOI21_X1 U7271 ( .B1(REIP_REG_7__SCAN_IN), .B2(n6202), .A(
        REIP_REG_8__SCAN_IN), .ZN(n6201) );
  OAI22_X1 U7272 ( .A1(n6193), .A2(n6257), .B1(n6977), .B2(n6253), .ZN(n6194)
         );
  AOI211_X1 U7273 ( .C1(EBX_REG_8__SCAN_IN), .C2(n6264), .A(n3952), .B(n6194), 
        .ZN(n6199) );
  AOI22_X1 U7274 ( .A1(n6197), .A2(n6220), .B1(n6196), .B2(n6195), .ZN(n6198)
         );
  OAI211_X1 U7275 ( .C1(n6201), .C2(n6200), .A(n6199), .B(n6198), .ZN(U2819)
         );
  AOI22_X1 U7276 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6264), .B1(n6202), .B2(n6647), 
        .ZN(n6213) );
  INV_X1 U7277 ( .A(n6203), .ZN(n6211) );
  OR2_X1 U7278 ( .A1(n6205), .A2(n6204), .ZN(n6223) );
  NAND2_X1 U7279 ( .A1(n6206), .A2(n6645), .ZN(n6216) );
  AOI21_X1 U7280 ( .B1(n6223), .B2(n6216), .A(n6647), .ZN(n6207) );
  AOI211_X1 U7281 ( .C1(n6239), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3952), 
        .B(n6207), .ZN(n6208) );
  OAI21_X1 U7282 ( .B1(n6257), .B2(n6209), .A(n6208), .ZN(n6210) );
  AOI21_X1 U7283 ( .B1(n6211), .B2(n6220), .A(n6210), .ZN(n6212) );
  OAI211_X1 U7284 ( .C1(n6214), .C2(n6258), .A(n6213), .B(n6212), .ZN(U2820)
         );
  OAI22_X1 U7285 ( .A1(n6223), .A2(n6645), .B1(n6257), .B2(n6215), .ZN(n6219)
         );
  AOI22_X1 U7286 ( .A1(EBX_REG_6__SCAN_IN), .A2(n6264), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6239), .ZN(n6217) );
  NAND3_X1 U7287 ( .A1(n6217), .A2(n6434), .A3(n6216), .ZN(n6218) );
  AOI211_X1 U7288 ( .C1(n6338), .C2(n6220), .A(n6219), .B(n6218), .ZN(n6221)
         );
  OAI21_X1 U7289 ( .B1(n6335), .B2(n6258), .A(n6221), .ZN(U2821) );
  AOI21_X1 U7290 ( .B1(n6246), .B2(n6222), .A(REIP_REG_5__SCAN_IN), .ZN(n6224)
         );
  NOR2_X1 U7291 ( .A1(n6224), .A2(n6223), .ZN(n6230) );
  NOR2_X1 U7292 ( .A1(n6225), .A2(n6257), .ZN(n6226) );
  AOI211_X1 U7293 ( .C1(n6239), .C2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3952), 
        .B(n6226), .ZN(n6227) );
  OAI21_X1 U7294 ( .B1(n6228), .B2(n6260), .A(n6227), .ZN(n6229) );
  AOI211_X1 U7295 ( .C1(EBX_REG_5__SCAN_IN), .C2(n6264), .A(n6230), .B(n6229), 
        .ZN(n6231) );
  OAI21_X1 U7296 ( .B1(n6232), .B2(n6258), .A(n6231), .ZN(U2822) );
  AOI22_X1 U7297 ( .A1(n6234), .A2(n6233), .B1(EBX_REG_4__SCAN_IN), .B2(n6264), 
        .ZN(n6250) );
  OAI21_X1 U7298 ( .B1(n6236), .B2(n6244), .A(n6235), .ZN(n6267) );
  OAI22_X1 U7299 ( .A1(n6267), .A2(n6641), .B1(n6257), .B2(n6237), .ZN(n6238)
         );
  AOI211_X1 U7300 ( .C1(n6239), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3952), 
        .B(n6238), .ZN(n6249) );
  INV_X1 U7301 ( .A(n6240), .ZN(n6241) );
  OAI22_X1 U7302 ( .A1(n6242), .A2(n6260), .B1(n6241), .B2(n6258), .ZN(n6243)
         );
  INV_X1 U7303 ( .A(n6243), .ZN(n6248) );
  INV_X1 U7304 ( .A(n6244), .ZN(n6245) );
  NAND3_X1 U7305 ( .A1(n6246), .A2(n6641), .A3(n6245), .ZN(n6247) );
  NAND4_X1 U7306 ( .A1(n6250), .A2(n6249), .A3(n6248), .A4(n6247), .ZN(U2823)
         );
  INV_X1 U7307 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6761) );
  NAND2_X1 U7308 ( .A1(n6251), .A2(REIP_REG_2__SCAN_IN), .ZN(n6266) );
  INV_X1 U7309 ( .A(n6391), .ZN(n6256) );
  INV_X1 U7310 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6252) );
  OAI222_X1 U7311 ( .A1(n6257), .A2(n6256), .B1(n6255), .B2(n6254), .C1(n6253), 
        .C2(n6252), .ZN(n6263) );
  OAI22_X1 U7312 ( .A1(n6261), .A2(n6260), .B1(n6259), .B2(n6258), .ZN(n6262)
         );
  AOI211_X1 U7313 ( .C1(EBX_REG_3__SCAN_IN), .C2(n6264), .A(n6263), .B(n6262), 
        .ZN(n6265) );
  OAI221_X1 U7314 ( .B1(n6267), .B2(n6761), .C1(n6267), .C2(n6266), .A(n6265), 
        .ZN(U2824) );
  AOI22_X1 U7315 ( .A1(n6268), .A2(n6744), .B1(n6271), .B2(DATAI_18_), .ZN(
        n6270) );
  AOI22_X1 U7316 ( .A1(n6273), .A2(DATAI_2_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n6743), .ZN(n6269) );
  NAND2_X1 U7317 ( .A1(n6270), .A2(n6269), .ZN(U2873) );
  AOI22_X1 U7318 ( .A1(n6272), .A2(n6744), .B1(n6271), .B2(DATAI_16_), .ZN(
        n6275) );
  AOI22_X1 U7319 ( .A1(n6273), .A2(DATAI_0_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n6743), .ZN(n6274) );
  NAND2_X1 U7320 ( .A1(n6275), .A2(n6274), .ZN(U2875) );
  INV_X1 U7321 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n6874) );
  INV_X1 U7322 ( .A(n6276), .ZN(n6280) );
  AOI22_X1 U7323 ( .A1(n6280), .A2(EAX_REG_29__SCAN_IN), .B1(n6305), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n6277) );
  OAI21_X1 U7324 ( .B1(n6874), .B2(n6301), .A(n6277), .ZN(U2894) );
  AOI22_X1 U7325 ( .A1(n6304), .A2(DATAO_REG_27__SCAN_IN), .B1(n6280), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6278) );
  OAI21_X1 U7326 ( .B1(n4487), .B2(n6730), .A(n6278), .ZN(U2896) );
  INV_X1 U7327 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n6750) );
  AOI22_X1 U7328 ( .A1(n6280), .A2(EAX_REG_20__SCAN_IN), .B1(n6305), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n6279) );
  OAI21_X1 U7329 ( .B1(n6750), .B2(n6301), .A(n6279), .ZN(U2903) );
  INV_X1 U7330 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n6841) );
  AOI22_X1 U7331 ( .A1(n6280), .A2(EAX_REG_18__SCAN_IN), .B1(n6305), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n6281) );
  OAI21_X1 U7332 ( .B1(n6841), .B2(n6301), .A(n6281), .ZN(U2905) );
  INV_X1 U7333 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n6946) );
  AOI22_X1 U7334 ( .A1(EAX_REG_15__SCAN_IN), .A2(n6298), .B1(n6304), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6282) );
  OAI21_X1 U7335 ( .B1(n6946), .B2(n6730), .A(n6282), .ZN(U2908) );
  INV_X1 U7336 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6883) );
  AOI22_X1 U7337 ( .A1(n6305), .A2(LWORD_REG_14__SCAN_IN), .B1(n6304), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6283) );
  OAI21_X1 U7338 ( .B1(n6883), .B2(n6307), .A(n6283), .ZN(U2909) );
  AOI22_X1 U7339 ( .A1(n6305), .A2(LWORD_REG_13__SCAN_IN), .B1(n6304), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6284) );
  OAI21_X1 U7340 ( .B1(n5482), .B2(n6307), .A(n6284), .ZN(U2910) );
  INV_X1 U7341 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n6776) );
  AOI22_X1 U7342 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6298), .B1(n6305), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n6285) );
  OAI21_X1 U7343 ( .B1(n6776), .B2(n6301), .A(n6285), .ZN(U2911) );
  AOI22_X1 U7344 ( .A1(n6305), .A2(LWORD_REG_11__SCAN_IN), .B1(n6304), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6286) );
  OAI21_X1 U7345 ( .B1(n6287), .B2(n6307), .A(n6286), .ZN(U2912) );
  INV_X1 U7346 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6289) );
  AOI22_X1 U7347 ( .A1(n6305), .A2(LWORD_REG_10__SCAN_IN), .B1(n6304), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6288) );
  OAI21_X1 U7348 ( .B1(n6289), .B2(n6307), .A(n6288), .ZN(U2913) );
  INV_X1 U7349 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6291) );
  AOI22_X1 U7350 ( .A1(n6305), .A2(LWORD_REG_9__SCAN_IN), .B1(n6304), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6290) );
  OAI21_X1 U7351 ( .B1(n6291), .B2(n6307), .A(n6290), .ZN(U2914) );
  INV_X1 U7352 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6293) );
  AOI22_X1 U7353 ( .A1(n6305), .A2(LWORD_REG_8__SCAN_IN), .B1(n6304), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6292) );
  OAI21_X1 U7354 ( .B1(n6293), .B2(n6307), .A(n6292), .ZN(U2915) );
  INV_X1 U7355 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n6792) );
  OAI222_X1 U7356 ( .A1(n4480), .A2(n6730), .B1(n6307), .B2(n3569), .C1(n6792), 
        .C2(n6301), .ZN(U2916) );
  AOI22_X1 U7357 ( .A1(n6305), .A2(LWORD_REG_6__SCAN_IN), .B1(n6304), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6294) );
  OAI21_X1 U7358 ( .B1(n6295), .B2(n6307), .A(n6294), .ZN(U2917) );
  INV_X1 U7359 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n6297) );
  INV_X1 U7360 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n6912) );
  OAI222_X1 U7361 ( .A1(n6297), .A2(n6730), .B1(n6307), .B2(n6296), .C1(n6912), 
        .C2(n6301), .ZN(U2918) );
  AOI22_X1 U7362 ( .A1(EAX_REG_4__SCAN_IN), .A2(n6298), .B1(n6304), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6299) );
  OAI21_X1 U7363 ( .B1(n4518), .B2(n6730), .A(n6299), .ZN(U2919) );
  INV_X1 U7364 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n6818) );
  OAI222_X1 U7365 ( .A1(n6301), .A2(n6818), .B1(n6307), .B2(n6300), .C1(n4489), 
        .C2(n6730), .ZN(U2920) );
  AOI22_X1 U7366 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n6305), .B1(n6304), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6302) );
  OAI21_X1 U7367 ( .B1(n6953), .B2(n6307), .A(n6302), .ZN(U2921) );
  AOI22_X1 U7368 ( .A1(n6305), .A2(LWORD_REG_1__SCAN_IN), .B1(n6304), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6303) );
  OAI21_X1 U7369 ( .B1(n4510), .B2(n6307), .A(n6303), .ZN(U2922) );
  AOI22_X1 U7370 ( .A1(n6305), .A2(LWORD_REG_0__SCAN_IN), .B1(n6304), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6306) );
  OAI21_X1 U7371 ( .B1(n6308), .B2(n6307), .A(n6306), .ZN(U2923) );
  AOI22_X1 U7372 ( .A1(EAX_REG_24__SCAN_IN), .A2(n6330), .B1(n6327), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n6309) );
  NAND2_X1 U7373 ( .A1(n6331), .A2(DATAI_8_), .ZN(n6318) );
  NAND2_X1 U7374 ( .A1(n6309), .A2(n6318), .ZN(U2932) );
  AOI22_X1 U7375 ( .A1(EAX_REG_25__SCAN_IN), .A2(n6330), .B1(n6327), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n6310) );
  NAND2_X1 U7376 ( .A1(n6331), .A2(DATAI_9_), .ZN(n6320) );
  NAND2_X1 U7377 ( .A1(n6310), .A2(n6320), .ZN(U2933) );
  NAND2_X1 U7378 ( .A1(n6331), .A2(DATAI_10_), .ZN(n6322) );
  INV_X1 U7379 ( .A(n6322), .ZN(n6311) );
  AOI21_X1 U7380 ( .B1(n6327), .B2(UWORD_REG_10__SCAN_IN), .A(n6311), .ZN(
        n6312) );
  OAI21_X1 U7381 ( .B1(n6313), .B2(n6329), .A(n6312), .ZN(U2934) );
  AOI22_X1 U7382 ( .A1(EAX_REG_28__SCAN_IN), .A2(n6330), .B1(n6327), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n6314) );
  NAND2_X1 U7383 ( .A1(n6331), .A2(DATAI_12_), .ZN(n6324) );
  NAND2_X1 U7384 ( .A1(n6314), .A2(n6324), .ZN(U2936) );
  INV_X1 U7385 ( .A(DATAI_14_), .ZN(n6315) );
  NOR2_X1 U7386 ( .A1(n6316), .A2(n6315), .ZN(n6326) );
  AOI21_X1 U7387 ( .B1(n6327), .B2(UWORD_REG_14__SCAN_IN), .A(n6326), .ZN(
        n6317) );
  OAI21_X1 U7388 ( .B1(n6849), .B2(n6329), .A(n6317), .ZN(U2938) );
  AOI22_X1 U7389 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6330), .B1(n6327), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U7390 ( .A1(n6319), .A2(n6318), .ZN(U2947) );
  AOI22_X1 U7391 ( .A1(EAX_REG_9__SCAN_IN), .A2(n6330), .B1(n6327), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n6321) );
  NAND2_X1 U7392 ( .A1(n6321), .A2(n6320), .ZN(U2948) );
  AOI22_X1 U7393 ( .A1(EAX_REG_10__SCAN_IN), .A2(n6330), .B1(n6327), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n6323) );
  NAND2_X1 U7394 ( .A1(n6323), .A2(n6322), .ZN(U2949) );
  AOI22_X1 U7395 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6330), .B1(n6327), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U7396 ( .A1(n6325), .A2(n6324), .ZN(U2951) );
  AOI21_X1 U7397 ( .B1(n6327), .B2(LWORD_REG_14__SCAN_IN), .A(n6326), .ZN(
        n6328) );
  OAI21_X1 U7398 ( .B1(n6883), .B2(n6329), .A(n6328), .ZN(U2953) );
  AOI22_X1 U7399 ( .A1(n6331), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6330), .ZN(n6332) );
  OAI21_X1 U7400 ( .B1(n6946), .B2(n6333), .A(n6332), .ZN(U2954) );
  INV_X1 U7401 ( .A(n6334), .ZN(n6339) );
  INV_X1 U7402 ( .A(n6335), .ZN(n6337) );
  AOI222_X1 U7403 ( .A1(n4310), .A2(n6339), .B1(n6338), .B2(n6347), .C1(n6337), 
        .C2(n6336), .ZN(n6341) );
  OAI211_X1 U7404 ( .C1(n6890), .C2(n6342), .A(n6341), .B(n6340), .ZN(U2980)
         );
  AOI22_X1 U7405 ( .A1(n3952), .A2(REIP_REG_2__SCAN_IN), .B1(n6358), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6350) );
  XNOR2_X1 U7406 ( .A(n6343), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6345)
         );
  XNOR2_X1 U7407 ( .A(n6345), .B(n6344), .ZN(n6408) );
  INV_X1 U7408 ( .A(n6346), .ZN(n6348) );
  AOI22_X1 U7409 ( .A1(n6408), .A2(n4310), .B1(n6348), .B2(n6347), .ZN(n6349)
         );
  OAI211_X1 U7410 ( .C1(n6352), .C2(n6351), .A(n6350), .B(n6349), .ZN(U2984)
         );
  OAI21_X1 U7411 ( .B1(n6354), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n6353), 
        .ZN(n6426) );
  OAI22_X1 U7412 ( .A1(n6426), .A2(n6355), .B1(n6434), .B2(n6724), .ZN(n6356)
         );
  INV_X1 U7413 ( .A(n6356), .ZN(n6360) );
  OAI21_X1 U7414 ( .B1(n6358), .B2(n6357), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n6359) );
  OAI211_X1 U7415 ( .C1(n6362), .C2(n6361), .A(n6360), .B(n6359), .ZN(U2986)
         );
  AOI22_X1 U7416 ( .A1(n6364), .A2(n6420), .B1(n6390), .B2(n6363), .ZN(n6369)
         );
  AOI22_X1 U7417 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6367), .B1(n6366), .B2(n6365), .ZN(n6368) );
  OAI211_X1 U7418 ( .C1(n5742), .C2(n6434), .A(n6369), .B(n6368), .ZN(U3007)
         );
  INV_X1 U7419 ( .A(n6370), .ZN(n6378) );
  AOI21_X1 U7420 ( .B1(n6372), .B2(n6390), .A(n6371), .ZN(n6376) );
  AOI22_X1 U7421 ( .A1(n6374), .A2(n6377), .B1(n6373), .B2(n6420), .ZN(n6375)
         );
  OAI211_X1 U7422 ( .C1(n6378), .C2(n6377), .A(n6376), .B(n6375), .ZN(U3009)
         );
  AOI21_X1 U7423 ( .B1(n6380), .B2(n6390), .A(n6379), .ZN(n6383) );
  NAND2_X1 U7424 ( .A1(n6381), .A2(n6420), .ZN(n6382) );
  OAI211_X1 U7425 ( .C1(n6384), .C2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6383), 
        .B(n6382), .ZN(n6385) );
  INV_X1 U7426 ( .A(n6385), .ZN(n6386) );
  OAI21_X1 U7427 ( .B1(n6388), .B2(n6387), .A(n6386), .ZN(U3011) );
  INV_X1 U7428 ( .A(n6389), .ZN(n6398) );
  NAND2_X1 U7429 ( .A1(n6391), .A2(n6390), .ZN(n6393) );
  OAI211_X1 U7430 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n6394), .A(n6393), 
        .B(n6392), .ZN(n6395) );
  AOI21_X1 U7431 ( .B1(n6396), .B2(n6420), .A(n6395), .ZN(n6397) );
  OAI21_X1 U7432 ( .B1(n6398), .B2(n7003), .A(n6397), .ZN(U3015) );
  INV_X1 U7433 ( .A(n6399), .ZN(n6400) );
  NAND2_X1 U7434 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6400), .ZN(n6411)
         );
  OAI21_X1 U7435 ( .B1(n6402), .B2(n6416), .A(n6401), .ZN(n6404) );
  AOI22_X1 U7436 ( .A1(n6413), .A2(n6404), .B1(n3952), .B2(REIP_REG_2__SCAN_IN), .ZN(n6405) );
  OAI21_X1 U7437 ( .B1(n6424), .B2(n6406), .A(n6405), .ZN(n6407) );
  AOI21_X1 U7438 ( .B1(n6408), .B2(n6420), .A(n6407), .ZN(n6409) );
  OAI221_X1 U7439 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6411), .C1(n3973), .C2(n6410), .A(n6409), .ZN(U3016) );
  AOI21_X1 U7440 ( .B1(n6413), .B2(n6416), .A(n6412), .ZN(n6428) );
  AOI211_X1 U7441 ( .C1(n6416), .C2(n6415), .A(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .B(n6414), .ZN(n6419) );
  OAI22_X1 U7442 ( .A1(n6424), .A2(n6417), .B1(n5755), .B2(n6434), .ZN(n6418)
         );
  AOI211_X1 U7443 ( .C1(n6421), .C2(n6420), .A(n6419), .B(n6418), .ZN(n6422)
         );
  OAI21_X1 U7444 ( .B1(n6428), .B2(n6900), .A(n6422), .ZN(U3017) );
  OAI22_X1 U7445 ( .A1(n6426), .A2(n6425), .B1(n6424), .B2(n6423), .ZN(n6427)
         );
  INV_X1 U7446 ( .A(n6427), .ZN(n6433) );
  INV_X1 U7447 ( .A(n6428), .ZN(n6430) );
  OAI22_X1 U7448 ( .A1(n6431), .A2(n6430), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6429), .ZN(n6432) );
  OAI211_X1 U7449 ( .C1(n6724), .C2(n6434), .A(n6433), .B(n6432), .ZN(U3018)
         );
  NOR2_X1 U7450 ( .A1(n6590), .A2(n6435), .ZN(U3019) );
  NAND3_X1 U7451 ( .A1(n6437), .A2(n6436), .A3(n7014), .ZN(n6438) );
  OAI21_X1 U7452 ( .B1(n6440), .B2(n6439), .A(n6438), .ZN(n6476) );
  NOR2_X1 U7453 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6441), .ZN(n6475)
         );
  AOI22_X1 U7454 ( .A1(n6514), .A2(n6476), .B1(n6504), .B2(n6475), .ZN(n6453)
         );
  NAND3_X1 U7455 ( .A1(n6501), .A2(n6450), .A3(n6442), .ZN(n6445) );
  AOI21_X1 U7456 ( .B1(n6445), .B2(n6444), .A(n6443), .ZN(n6448) );
  OAI211_X1 U7457 ( .C1(n6475), .C2(n6702), .A(n6446), .B(n7014), .ZN(n6447)
         );
  AOI22_X1 U7458 ( .A1(n6479), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6451), 
        .B2(n6477), .ZN(n6452) );
  OAI211_X1 U7459 ( .C1(n6454), .C2(n6501), .A(n6453), .B(n6452), .ZN(U3068)
         );
  AOI22_X1 U7460 ( .A1(n6520), .A2(n6476), .B1(n6519), .B2(n6475), .ZN(n6457)
         );
  AOI22_X1 U7461 ( .A1(n6479), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6455), 
        .B2(n6477), .ZN(n6456) );
  OAI211_X1 U7462 ( .C1(n6458), .C2(n6501), .A(n6457), .B(n6456), .ZN(U3069)
         );
  AOI22_X1 U7463 ( .A1(n6526), .A2(n6476), .B1(n6525), .B2(n6475), .ZN(n6461)
         );
  AOI22_X1 U7464 ( .A1(n6479), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6459), 
        .B2(n6477), .ZN(n6460) );
  OAI211_X1 U7465 ( .C1(n6462), .C2(n6501), .A(n6461), .B(n6460), .ZN(U3070)
         );
  AOI22_X1 U7466 ( .A1(n6532), .A2(n6476), .B1(n6531), .B2(n6475), .ZN(n6465)
         );
  AOI22_X1 U7467 ( .A1(n6479), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6463), 
        .B2(n6477), .ZN(n6464) );
  OAI211_X1 U7468 ( .C1(n6466), .C2(n6501), .A(n6465), .B(n6464), .ZN(U3071)
         );
  AOI22_X1 U7469 ( .A1(n6538), .A2(n6476), .B1(n6537), .B2(n6475), .ZN(n6468)
         );
  AOI22_X1 U7470 ( .A1(n6479), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6536), 
        .B2(n6477), .ZN(n6467) );
  OAI211_X1 U7471 ( .C1(n6541), .C2(n6501), .A(n6468), .B(n6467), .ZN(U3072)
         );
  AOI22_X1 U7472 ( .A1(n6544), .A2(n6476), .B1(n6543), .B2(n6475), .ZN(n6471)
         );
  AOI22_X1 U7473 ( .A1(n6479), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6469), 
        .B2(n6477), .ZN(n6470) );
  OAI211_X1 U7474 ( .C1(n6472), .C2(n6501), .A(n6471), .B(n6470), .ZN(U3073)
         );
  AOI22_X1 U7475 ( .A1(n6551), .A2(n6476), .B1(n6550), .B2(n6475), .ZN(n6474)
         );
  AOI22_X1 U7476 ( .A1(n6479), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6548), 
        .B2(n6477), .ZN(n6473) );
  OAI211_X1 U7477 ( .C1(n6555), .C2(n6501), .A(n6474), .B(n6473), .ZN(U3074)
         );
  AOI22_X1 U7478 ( .A1(n6561), .A2(n6476), .B1(n6559), .B2(n6475), .ZN(n6481)
         );
  AOI22_X1 U7479 ( .A1(n6479), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6478), 
        .B2(n6477), .ZN(n6480) );
  OAI211_X1 U7480 ( .C1(n6482), .C2(n6501), .A(n6481), .B(n6480), .ZN(U3075)
         );
  AOI22_X1 U7481 ( .A1(n6504), .A2(n6496), .B1(n6503), .B2(n6495), .ZN(n6484)
         );
  AOI22_X1 U7482 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6498), .B1(n6514), 
        .B2(n6497), .ZN(n6483) );
  OAI211_X1 U7483 ( .C1(n6517), .C2(n6501), .A(n6484), .B(n6483), .ZN(U3076)
         );
  AOI22_X1 U7484 ( .A1(n6519), .A2(n6496), .B1(n6518), .B2(n6495), .ZN(n6486)
         );
  AOI22_X1 U7485 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6498), .B1(n6520), 
        .B2(n6497), .ZN(n6485) );
  OAI211_X1 U7486 ( .C1(n6523), .C2(n6501), .A(n6486), .B(n6485), .ZN(U3077)
         );
  AOI22_X1 U7487 ( .A1(n6531), .A2(n6496), .B1(n6530), .B2(n6495), .ZN(n6488)
         );
  AOI22_X1 U7488 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6498), .B1(n6532), 
        .B2(n6497), .ZN(n6487) );
  OAI211_X1 U7489 ( .C1(n6535), .C2(n6501), .A(n6488), .B(n6487), .ZN(U3079)
         );
  AOI22_X1 U7490 ( .A1(n6543), .A2(n6496), .B1(n6542), .B2(n6495), .ZN(n6490)
         );
  AOI22_X1 U7491 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6498), .B1(n6544), 
        .B2(n6497), .ZN(n6489) );
  OAI211_X1 U7492 ( .C1(n6547), .C2(n6501), .A(n6490), .B(n6489), .ZN(U3081)
         );
  AOI22_X1 U7493 ( .A1(n6550), .A2(n6496), .B1(n6491), .B2(n6495), .ZN(n6493)
         );
  AOI22_X1 U7494 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6498), .B1(n6551), 
        .B2(n6497), .ZN(n6492) );
  OAI211_X1 U7495 ( .C1(n6494), .C2(n6501), .A(n6493), .B(n6492), .ZN(U3082)
         );
  AOI22_X1 U7496 ( .A1(n6559), .A2(n6496), .B1(n6556), .B2(n6495), .ZN(n6500)
         );
  AOI22_X1 U7497 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6498), .B1(n6561), 
        .B2(n6497), .ZN(n6499) );
  OAI211_X1 U7498 ( .C1(n6566), .C2(n6501), .A(n6500), .B(n6499), .ZN(U3083)
         );
  NOR2_X1 U7499 ( .A1(n6502), .A2(n7014), .ZN(n6558) );
  AOI22_X1 U7500 ( .A1(n6504), .A2(n6558), .B1(n6557), .B2(n6503), .ZN(n6516)
         );
  OAI21_X1 U7501 ( .B1(n6506), .B2(n6505), .A(n6442), .ZN(n6513) );
  AOI21_X1 U7502 ( .B1(n6507), .B2(n6575), .A(n6558), .ZN(n6512) );
  INV_X1 U7503 ( .A(n6512), .ZN(n6510) );
  AOI21_X1 U7504 ( .B1(n6729), .B2(n6511), .A(n6508), .ZN(n6509) );
  OAI21_X1 U7505 ( .B1(n6513), .B2(n6510), .A(n6509), .ZN(n6562) );
  OAI22_X1 U7506 ( .A1(n6513), .A2(n6512), .B1(n6511), .B2(n6935), .ZN(n6560)
         );
  AOI22_X1 U7507 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6562), .B1(n6514), 
        .B2(n6560), .ZN(n6515) );
  OAI211_X1 U7508 ( .C1(n6517), .C2(n6565), .A(n6516), .B(n6515), .ZN(U3108)
         );
  AOI22_X1 U7509 ( .A1(n6519), .A2(n6558), .B1(n6557), .B2(n6518), .ZN(n6522)
         );
  AOI22_X1 U7510 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6562), .B1(n6520), 
        .B2(n6560), .ZN(n6521) );
  OAI211_X1 U7511 ( .C1(n6523), .C2(n6565), .A(n6522), .B(n6521), .ZN(U3109)
         );
  AOI22_X1 U7512 ( .A1(n6525), .A2(n6558), .B1(n6557), .B2(n6524), .ZN(n6528)
         );
  AOI22_X1 U7513 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6562), .B1(n6526), 
        .B2(n6560), .ZN(n6527) );
  OAI211_X1 U7514 ( .C1(n6529), .C2(n6565), .A(n6528), .B(n6527), .ZN(U3110)
         );
  AOI22_X1 U7515 ( .A1(n6531), .A2(n6558), .B1(n6557), .B2(n6530), .ZN(n6534)
         );
  AOI22_X1 U7516 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6562), .B1(n6532), 
        .B2(n6560), .ZN(n6533) );
  OAI211_X1 U7517 ( .C1(n6535), .C2(n6565), .A(n6534), .B(n6533), .ZN(U3111)
         );
  AOI22_X1 U7518 ( .A1(n6537), .A2(n6558), .B1(n6549), .B2(n6536), .ZN(n6540)
         );
  AOI22_X1 U7519 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6562), .B1(n6538), 
        .B2(n6560), .ZN(n6539) );
  OAI211_X1 U7520 ( .C1(n6541), .C2(n6554), .A(n6540), .B(n6539), .ZN(U3112)
         );
  AOI22_X1 U7521 ( .A1(n6543), .A2(n6558), .B1(n6557), .B2(n6542), .ZN(n6546)
         );
  AOI22_X1 U7522 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6562), .B1(n6544), 
        .B2(n6560), .ZN(n6545) );
  OAI211_X1 U7523 ( .C1(n6547), .C2(n6565), .A(n6546), .B(n6545), .ZN(U3113)
         );
  AOI22_X1 U7524 ( .A1(n6550), .A2(n6558), .B1(n6549), .B2(n6548), .ZN(n6553)
         );
  AOI22_X1 U7525 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6562), .B1(n6551), 
        .B2(n6560), .ZN(n6552) );
  OAI211_X1 U7526 ( .C1(n6555), .C2(n6554), .A(n6553), .B(n6552), .ZN(U3114)
         );
  AOI22_X1 U7527 ( .A1(n6559), .A2(n6558), .B1(n6557), .B2(n6556), .ZN(n6564)
         );
  AOI22_X1 U7528 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6562), .B1(n6561), 
        .B2(n6560), .ZN(n6563) );
  OAI211_X1 U7529 ( .C1(n6566), .C2(n6565), .A(n6564), .B(n6563), .ZN(U3115)
         );
  OAI21_X1 U7530 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6567), 
        .ZN(n6568) );
  NAND4_X1 U7531 ( .A1(n6571), .A2(n6570), .A3(n6569), .A4(n6568), .ZN(n6572)
         );
  NOR2_X1 U7532 ( .A1(n6573), .A2(n6572), .ZN(n6594) );
  NAND2_X1 U7533 ( .A1(n6592), .A2(n7014), .ZN(n6589) );
  AOI22_X1 U7534 ( .A1(n6575), .A2(n6574), .B1(n3704), .B2(n3921), .ZN(n6710)
         );
  NAND2_X1 U7535 ( .A1(n6576), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6716) );
  NAND3_X1 U7536 ( .A1(n6710), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6716), .ZN(n6578) );
  OAI21_X1 U7537 ( .B1(n6579), .B2(n6578), .A(n6577), .ZN(n6581) );
  NAND2_X1 U7538 ( .A1(n6579), .A2(n6578), .ZN(n6580) );
  OAI21_X1 U7539 ( .B1(n6582), .B2(n6581), .A(n6580), .ZN(n6587) );
  NAND2_X1 U7540 ( .A1(n6586), .A2(n6587), .ZN(n6583) );
  NAND2_X1 U7541 ( .A1(n6584), .A2(n6583), .ZN(n6585) );
  OAI21_X1 U7542 ( .B1(n6587), .B2(n6586), .A(n6585), .ZN(n6588) );
  NAND2_X1 U7543 ( .A1(n6589), .A2(n6588), .ZN(n6591) );
  OAI211_X1 U7544 ( .C1(n6592), .C2(n7014), .A(n6591), .B(n6590), .ZN(n6593)
         );
  NAND2_X1 U7545 ( .A1(n6594), .A2(n6593), .ZN(n6605) );
  OAI22_X1 U7546 ( .A1(n6605), .A2(n6612), .B1(n6630), .B2(n6730), .ZN(n6600)
         );
  INV_X1 U7547 ( .A(n6595), .ZN(n6598) );
  NOR3_X1 U7548 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .A3(n6596), .ZN(
        n6597) );
  NAND2_X1 U7549 ( .A1(n6598), .A2(n6597), .ZN(n6599) );
  AOI21_X1 U7550 ( .B1(READY_N), .B2(n6935), .A(n6698), .ZN(n6610) );
  NOR2_X1 U7551 ( .A1(n6702), .A2(n6616), .ZN(n6602) );
  AOI211_X1 U7552 ( .C1(n6602), .C2(n6601), .A(STATE2_REG_0__SCAN_IN), .B(
        n6698), .ZN(n6603) );
  AOI211_X1 U7553 ( .C1(n6606), .C2(n6605), .A(n6604), .B(n6603), .ZN(n6607)
         );
  OAI221_X1 U7554 ( .B1(n6609), .B2(n6610), .C1(n6609), .C2(n6608), .A(n6607), 
        .ZN(U3148) );
  NOR3_X1 U7555 ( .A1(n6619), .A2(n6610), .A3(n6709), .ZN(n6614) );
  AOI221_X1 U7556 ( .B1(READY_N), .B2(n6612), .C1(n6611), .C2(n6612), .A(n6698), .ZN(n6613) );
  OR3_X1 U7557 ( .A1(n6615), .A2(n6614), .A3(n6613), .ZN(U3149) );
  OAI211_X1 U7558 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6630), .A(n6699), .B(
        n6616), .ZN(n6618) );
  OAI21_X1 U7559 ( .B1(n6619), .B2(n6618), .A(n6617), .ZN(U3150) );
  NOR2_X1 U7560 ( .A1(n6697), .A2(n6803), .ZN(U3151) );
  INV_X1 U7561 ( .A(n6697), .ZN(n6695) );
  AND2_X1 U7562 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6695), .ZN(U3152) );
  AND2_X1 U7563 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6695), .ZN(U3153) );
  AND2_X1 U7564 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6695), .ZN(U3154) );
  INV_X1 U7565 ( .A(DATAWIDTH_REG_27__SCAN_IN), .ZN(n6861) );
  NOR2_X1 U7566 ( .A1(n6697), .A2(n6861), .ZN(U3155) );
  AND2_X1 U7567 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6695), .ZN(U3156) );
  AND2_X1 U7568 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6695), .ZN(U3157) );
  AND2_X1 U7569 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6695), .ZN(U3158) );
  AND2_X1 U7570 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6695), .ZN(U3159) );
  INV_X1 U7571 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6898) );
  NOR2_X1 U7572 ( .A1(n6697), .A2(n6898), .ZN(U3160) );
  NOR2_X1 U7573 ( .A1(n6697), .A2(n6920), .ZN(U3161) );
  AND2_X1 U7574 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6695), .ZN(U3162) );
  INV_X1 U7575 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n6833) );
  NOR2_X1 U7576 ( .A1(n6697), .A2(n6833), .ZN(U3163) );
  INV_X1 U7577 ( .A(DATAWIDTH_REG_18__SCAN_IN), .ZN(n6932) );
  NOR2_X1 U7578 ( .A1(n6697), .A2(n6932), .ZN(U3164) );
  AND2_X1 U7579 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6695), .ZN(U3165) );
  NOR2_X1 U7580 ( .A1(n6697), .A2(n6959), .ZN(U3166) );
  AND2_X1 U7581 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6695), .ZN(U3167) );
  AND2_X1 U7582 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6695), .ZN(U3168) );
  AND2_X1 U7583 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6695), .ZN(U3169) );
  INV_X1 U7584 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6777) );
  NOR2_X1 U7585 ( .A1(n6697), .A2(n6777), .ZN(U3170) );
  AND2_X1 U7586 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6695), .ZN(U3171) );
  AND2_X1 U7587 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6695), .ZN(U3172) );
  NOR2_X1 U7588 ( .A1(n6697), .A2(n6917), .ZN(U3173) );
  INV_X1 U7589 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6944) );
  NOR2_X1 U7590 ( .A1(n6697), .A2(n6944), .ZN(U3174) );
  INV_X1 U7591 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6929) );
  NOR2_X1 U7592 ( .A1(n6697), .A2(n6929), .ZN(U3175) );
  NOR2_X1 U7593 ( .A1(n6697), .A2(n6863), .ZN(U3176) );
  AND2_X1 U7594 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6695), .ZN(U3177) );
  AND2_X1 U7595 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6695), .ZN(U3178) );
  AND2_X1 U7596 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6695), .ZN(U3179) );
  INV_X1 U7597 ( .A(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6927) );
  NOR2_X1 U7598 ( .A1(n6697), .A2(n6927), .ZN(U3180) );
  NAND2_X1 U7599 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6624) );
  AND2_X1 U7600 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6623) );
  NAND2_X1 U7601 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .ZN(
        n6621) );
  NOR2_X1 U7602 ( .A1(n6630), .A2(n6974), .ZN(n6629) );
  AOI21_X1 U7603 ( .B1(NA_N), .B2(n6974), .A(n6975), .ZN(n6620) );
  NOR2_X1 U7604 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6620), .ZN(n6636) );
  AOI221_X1 U7605 ( .B1(n6623), .B2(n6621), .C1(n6629), .C2(n6621), .A(n6636), 
        .ZN(n6622) );
  OAI221_X1 U7606 ( .B1(n6741), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n6741), 
        .C2(n6624), .A(n6622), .ZN(U3181) );
  NAND2_X1 U7607 ( .A1(STATE_REG_0__SCAN_IN), .A2(REQUESTPENDING_REG_SCAN_IN), 
        .ZN(n6625) );
  AOI21_X1 U7608 ( .B1(n6625), .B2(n6624), .A(n6623), .ZN(n6626) );
  OR3_X1 U7609 ( .A1(n6627), .A2(n6629), .A3(n6626), .ZN(U3182) );
  AOI221_X1 U7610 ( .B1(HOLD), .B2(STATE_REG_2__SCAN_IN), .C1(n6629), .C2(
        STATE_REG_2__SCAN_IN), .A(n6628), .ZN(n6635) );
  NOR2_X1 U7611 ( .A1(NA_N), .A2(n6630), .ZN(n6632) );
  INV_X1 U7612 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6631) );
  OAI211_X1 U7613 ( .C1(n6632), .C2(n6974), .A(HOLD), .B(n6631), .ZN(n6634) );
  NAND4_X1 U7614 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .A3(
        REQUESTPENDING_REG_SCAN_IN), .A4(n6632), .ZN(n6633) );
  OAI221_X1 U7615 ( .B1(n6636), .B2(n6635), .C1(n6636), .C2(n6634), .A(n6633), 
        .ZN(U3183) );
  NAND2_X1 U7616 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6741), .ZN(n6681) );
  AOI22_X1 U7617 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6727), .ZN(n6637) );
  OAI21_X1 U7618 ( .B1(n5755), .B2(n6681), .A(n6637), .ZN(U3184) );
  INV_X1 U7619 ( .A(n6681), .ZN(n6687) );
  AOI22_X1 U7620 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6727), .ZN(n6638) );
  OAI21_X1 U7621 ( .B1(n5325), .B2(n6685), .A(n6638), .ZN(U3185) );
  AOI22_X1 U7622 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6727), .ZN(n6639) );
  OAI21_X1 U7623 ( .B1(n6761), .B2(n6685), .A(n6639), .ZN(U3186) );
  AOI22_X1 U7624 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6727), .ZN(n6640) );
  OAI21_X1 U7625 ( .B1(n6641), .B2(n6685), .A(n6640), .ZN(U3187) );
  INV_X1 U7626 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6643) );
  AOI22_X1 U7627 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6727), .ZN(n6642) );
  OAI21_X1 U7628 ( .B1(n6643), .B2(n6685), .A(n6642), .ZN(U3188) );
  AOI22_X1 U7629 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6727), .ZN(n6644) );
  OAI21_X1 U7630 ( .B1(n6645), .B2(n6685), .A(n6644), .ZN(U3189) );
  AOI22_X1 U7631 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6727), .ZN(n6646) );
  OAI21_X1 U7632 ( .B1(n6647), .B2(n6685), .A(n6646), .ZN(U3190) );
  AOI22_X1 U7633 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6727), .ZN(n6648) );
  OAI21_X1 U7634 ( .B1(n6649), .B2(n6685), .A(n6648), .ZN(U3191) );
  AOI22_X1 U7635 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6727), .ZN(n6650) );
  OAI21_X1 U7636 ( .B1(n6651), .B2(n6685), .A(n6650), .ZN(U3192) );
  AOI22_X1 U7637 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6727), .ZN(n6652) );
  OAI21_X1 U7638 ( .B1(n6653), .B2(n6685), .A(n6652), .ZN(U3193) );
  AOI22_X1 U7639 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6727), .ZN(n6654) );
  OAI21_X1 U7640 ( .B1(n5742), .B2(n6685), .A(n6654), .ZN(U3194) );
  AOI22_X1 U7641 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6727), .ZN(n6655) );
  OAI21_X1 U7642 ( .B1(n6808), .B2(n6685), .A(n6655), .ZN(U3195) );
  AOI22_X1 U7643 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6683), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6727), .ZN(n6656) );
  OAI21_X1 U7644 ( .B1(n6657), .B2(n6685), .A(n6656), .ZN(U3196) );
  AOI22_X1 U7645 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6683), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6727), .ZN(n6658) );
  OAI21_X1 U7646 ( .B1(n6659), .B2(n6681), .A(n6658), .ZN(U3197) );
  AOI22_X1 U7647 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6683), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6727), .ZN(n6660) );
  OAI21_X1 U7648 ( .B1(n7002), .B2(n6681), .A(n6660), .ZN(U3198) );
  AOI22_X1 U7649 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6683), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6727), .ZN(n6661) );
  OAI21_X1 U7650 ( .B1(n6662), .B2(n6681), .A(n6661), .ZN(U3199) );
  AOI22_X1 U7651 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6683), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6727), .ZN(n6663) );
  OAI21_X1 U7652 ( .B1(n6664), .B2(n6681), .A(n6663), .ZN(U3200) );
  AOI22_X1 U7653 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6683), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6727), .ZN(n6665) );
  OAI21_X1 U7654 ( .B1(n6666), .B2(n6681), .A(n6665), .ZN(U3201) );
  AOI22_X1 U7655 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6727), .ZN(n6667) );
  OAI21_X1 U7656 ( .B1(n6668), .B2(n6681), .A(n6667), .ZN(U3202) );
  AOI22_X1 U7657 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6687), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6727), .ZN(n6669) );
  OAI21_X1 U7658 ( .B1(n6670), .B2(n6689), .A(n6669), .ZN(U3203) );
  AOI22_X1 U7659 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6687), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6727), .ZN(n6671) );
  OAI21_X1 U7660 ( .B1(n6955), .B2(n6689), .A(n6671), .ZN(U3204) );
  AOI22_X1 U7661 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6687), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6727), .ZN(n6672) );
  OAI21_X1 U7662 ( .B1(n6674), .B2(n6689), .A(n6672), .ZN(U3205) );
  AOI22_X1 U7663 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6727), .ZN(n6673) );
  OAI21_X1 U7664 ( .B1(n6674), .B2(n6681), .A(n6673), .ZN(U3206) );
  AOI22_X1 U7665 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6727), .ZN(n6676) );
  OAI21_X1 U7666 ( .B1(n6677), .B2(n6681), .A(n6676), .ZN(U3207) );
  AOI22_X1 U7667 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6683), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6727), .ZN(n6678) );
  OAI21_X1 U7668 ( .B1(n6846), .B2(n6681), .A(n6678), .ZN(U3208) );
  INV_X1 U7669 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6832) );
  OAI222_X1 U7670 ( .A1(n6685), .A2(n6679), .B1(n6832), .B2(n6741), .C1(n6680), 
        .C2(n6689), .ZN(U3209) );
  INV_X1 U7671 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6873) );
  INV_X1 U7672 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6682) );
  OAI222_X1 U7673 ( .A1(n6681), .A2(n6680), .B1(n6873), .B2(n6741), .C1(n6682), 
        .C2(n6689), .ZN(U3210) );
  INV_X1 U7674 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6760) );
  OAI222_X1 U7675 ( .A1(n6685), .A2(n6682), .B1(n6760), .B2(n6741), .C1(n6686), 
        .C2(n6689), .ZN(U3211) );
  AOI22_X1 U7676 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6683), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6727), .ZN(n6684) );
  OAI21_X1 U7677 ( .B1(n6686), .B2(n6685), .A(n6684), .ZN(U3212) );
  INV_X1 U7678 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6690) );
  AOI22_X1 U7679 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6687), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6727), .ZN(n6688) );
  OAI21_X1 U7680 ( .B1(n6690), .B2(n6689), .A(n6688), .ZN(U3213) );
  INV_X1 U7681 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6691) );
  INV_X1 U7682 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n6886) );
  AOI22_X1 U7683 ( .A1(n6741), .A2(n6691), .B1(n6886), .B2(n6727), .ZN(U3445)
         );
  INV_X1 U7684 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6692) );
  INV_X1 U7685 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n6789) );
  AOI22_X1 U7686 ( .A1(n6741), .A2(n6692), .B1(n6789), .B2(n6727), .ZN(U3446)
         );
  INV_X1 U7687 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6693) );
  INV_X1 U7688 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n6848) );
  AOI22_X1 U7689 ( .A1(n6741), .A2(n6693), .B1(n6848), .B2(n6727), .ZN(U3447)
         );
  MUX2_X1 U7690 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6741), .Z(U3448) );
  INV_X1 U7691 ( .A(n6696), .ZN(n6694) );
  AOI21_X1 U7692 ( .B1(n6718), .B2(n6695), .A(n6694), .ZN(U3451) );
  OAI21_X1 U7693 ( .B1(n6697), .B2(n6717), .A(n6696), .ZN(U3452) );
  INV_X1 U7694 ( .A(n6698), .ZN(n6701) );
  OAI211_X1 U7695 ( .C1(n6702), .C2(n6701), .A(n6700), .B(n6699), .ZN(U3453)
         );
  INV_X1 U7696 ( .A(n6703), .ZN(n6706) );
  OAI22_X1 U7697 ( .A1(n6706), .A2(n6715), .B1(n6705), .B2(n6704), .ZN(n6708)
         );
  MUX2_X1 U7698 ( .A(n6708), .B(n6988), .S(n6707), .Z(U3456) );
  OAI22_X1 U7699 ( .A1(n6710), .A2(n6715), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6709), .ZN(n6712) );
  OAI22_X1 U7700 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6713), .B1(n6712), .B2(n6711), .ZN(n6714) );
  OAI21_X1 U7701 ( .B1(n6716), .B2(n6715), .A(n6714), .ZN(U3461) );
  OAI211_X1 U7702 ( .C1(n6718), .C2(n6724), .A(n6717), .B(n6725), .ZN(n6722)
         );
  OAI21_X1 U7703 ( .B1(n6724), .B2(n5755), .A(n6720), .ZN(n6719) );
  OAI21_X1 U7704 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(n6720), .A(n6719), .ZN(
        n6721) );
  NAND2_X1 U7705 ( .A1(n6722), .A2(n6721), .ZN(U3468) );
  INV_X1 U7706 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6859) );
  AOI22_X1 U7707 ( .A1(n6725), .A2(n6724), .B1(n6859), .B2(n6723), .ZN(U3469)
         );
  NAND2_X1 U7708 ( .A1(n6727), .A2(W_R_N_REG_SCAN_IN), .ZN(n6726) );
  OAI21_X1 U7709 ( .B1(n6727), .B2(READREQUEST_REG_SCAN_IN), .A(n6726), .ZN(
        U3470) );
  OAI211_X1 U7710 ( .C1(READY_N), .C2(n6730), .A(n6729), .B(n6728), .ZN(n6731)
         );
  NOR2_X1 U7711 ( .A1(n6732), .A2(n6731), .ZN(n6740) );
  INV_X1 U7712 ( .A(n6733), .ZN(n6734) );
  OAI211_X1 U7713 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6735), .A(n6734), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6737) );
  AOI21_X1 U7714 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6737), .A(n6736), .ZN(
        n6739) );
  NAND2_X1 U7715 ( .A1(n6740), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6738) );
  OAI21_X1 U7716 ( .B1(n6740), .B2(n6739), .A(n6738), .ZN(U3472) );
  MUX2_X1 U7717 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6741), .Z(U3473) );
  AOI222_X1 U7718 ( .A1(n6745), .A2(n6744), .B1(EAX_REG_14__SCAN_IN), .B2(
        n6743), .C1(DATAI_14_), .C2(n6742), .ZN(n6973) );
  INV_X1 U7719 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n6990) );
  AOI22_X1 U7720 ( .A1(n7031), .A2(keyinput10), .B1(n6990), .B2(keyinput55), 
        .ZN(n6746) );
  OAI221_X1 U7721 ( .B1(n7031), .B2(keyinput10), .C1(n6990), .C2(keyinput55), 
        .A(n6746), .ZN(n6755) );
  INV_X1 U7722 ( .A(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n7022) );
  AOI22_X1 U7723 ( .A1(n7022), .A2(keyinput3), .B1(keyinput5), .B2(n7014), 
        .ZN(n6747) );
  OAI221_X1 U7724 ( .B1(n7022), .B2(keyinput3), .C1(n7014), .C2(keyinput5), 
        .A(n6747), .ZN(n6754) );
  AOI22_X1 U7725 ( .A1(n6750), .A2(keyinput116), .B1(n6749), .B2(keyinput115), 
        .ZN(n6748) );
  OAI221_X1 U7726 ( .B1(n6750), .B2(keyinput116), .C1(n6749), .C2(keyinput115), 
        .A(n6748), .ZN(n6753) );
  AOI22_X1 U7727 ( .A1(n7009), .A2(keyinput106), .B1(keyinput59), .B2(n7003), 
        .ZN(n6751) );
  OAI221_X1 U7728 ( .B1(n7009), .B2(keyinput106), .C1(n7003), .C2(keyinput59), 
        .A(n6751), .ZN(n6752) );
  NOR4_X1 U7729 ( .A1(n6755), .A2(n6754), .A3(n6753), .A4(n6752), .ZN(n6800)
         );
  AOI22_X1 U7730 ( .A1(n6758), .A2(keyinput84), .B1(keyinput127), .B2(n6757), 
        .ZN(n6756) );
  OAI221_X1 U7731 ( .B1(n6758), .B2(keyinput84), .C1(n6757), .C2(keyinput127), 
        .A(n6756), .ZN(n6770) );
  AOI22_X1 U7732 ( .A1(n6761), .A2(keyinput107), .B1(keyinput118), .B2(n6760), 
        .ZN(n6759) );
  OAI221_X1 U7733 ( .B1(n6761), .B2(keyinput107), .C1(n6760), .C2(keyinput118), 
        .A(n6759), .ZN(n6769) );
  INV_X1 U7734 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n6764) );
  INV_X1 U7735 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n6763) );
  AOI22_X1 U7736 ( .A1(n6764), .A2(keyinput16), .B1(keyinput13), .B2(n6763), 
        .ZN(n6762) );
  OAI221_X1 U7737 ( .B1(n6764), .B2(keyinput16), .C1(n6763), .C2(keyinput13), 
        .A(n6762), .ZN(n6768) );
  INV_X1 U7738 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n6766) );
  AOI22_X1 U7739 ( .A1(n6766), .A2(keyinput40), .B1(keyinput19), .B2(n4968), 
        .ZN(n6765) );
  OAI221_X1 U7740 ( .B1(n6766), .B2(keyinput40), .C1(n4968), .C2(keyinput19), 
        .A(n6765), .ZN(n6767) );
  NOR4_X1 U7741 ( .A1(n6770), .A2(n6769), .A3(n6768), .A4(n6767), .ZN(n6799)
         );
  INV_X1 U7742 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n6772) );
  AOI22_X1 U7743 ( .A1(n6975), .A2(keyinput96), .B1(n6772), .B2(keyinput12), 
        .ZN(n6771) );
  OAI221_X1 U7744 ( .B1(n6975), .B2(keyinput96), .C1(n6772), .C2(keyinput12), 
        .A(n6771), .ZN(n6783) );
  AOI22_X1 U7745 ( .A1(n4679), .A2(keyinput49), .B1(n6774), .B2(keyinput114), 
        .ZN(n6773) );
  OAI221_X1 U7746 ( .B1(n4679), .B2(keyinput49), .C1(n6774), .C2(keyinput114), 
        .A(n6773), .ZN(n6782) );
  AOI22_X1 U7747 ( .A1(n6777), .A2(keyinput45), .B1(n6776), .B2(keyinput39), 
        .ZN(n6775) );
  OAI221_X1 U7748 ( .B1(n6777), .B2(keyinput45), .C1(n6776), .C2(keyinput39), 
        .A(n6775), .ZN(n6781) );
  XOR2_X1 U7749 ( .A(n5261), .B(keyinput14), .Z(n6779) );
  XNOR2_X1 U7750 ( .A(n6988), .B(keyinput124), .ZN(n6778) );
  NAND2_X1 U7751 ( .A1(n6779), .A2(n6778), .ZN(n6780) );
  NOR4_X1 U7752 ( .A1(n6783), .A2(n6782), .A3(n6781), .A4(n6780), .ZN(n6798)
         );
  INV_X1 U7753 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n6786) );
  INV_X1 U7754 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n6785) );
  AOI22_X1 U7755 ( .A1(n6786), .A2(keyinput41), .B1(n6785), .B2(keyinput38), 
        .ZN(n6784) );
  OAI221_X1 U7756 ( .B1(n6786), .B2(keyinput41), .C1(n6785), .C2(keyinput38), 
        .A(n6784), .ZN(n6796) );
  AOI22_X1 U7757 ( .A1(n4983), .A2(keyinput126), .B1(keyinput79), .B2(n4518), 
        .ZN(n6787) );
  OAI221_X1 U7758 ( .B1(n4983), .B2(keyinput126), .C1(n4518), .C2(keyinput79), 
        .A(n6787), .ZN(n6795) );
  INV_X1 U7759 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n6790) );
  AOI22_X1 U7760 ( .A1(n6790), .A2(keyinput50), .B1(keyinput76), .B2(n6789), 
        .ZN(n6788) );
  OAI221_X1 U7761 ( .B1(n6790), .B2(keyinput50), .C1(n6789), .C2(keyinput76), 
        .A(n6788), .ZN(n6794) );
  AOI22_X1 U7762 ( .A1(n4491), .A2(keyinput18), .B1(n6792), .B2(keyinput57), 
        .ZN(n6791) );
  OAI221_X1 U7763 ( .B1(n4491), .B2(keyinput18), .C1(n6792), .C2(keyinput57), 
        .A(n6791), .ZN(n6793) );
  NOR4_X1 U7764 ( .A1(n6796), .A2(n6795), .A3(n6794), .A4(n6793), .ZN(n6797)
         );
  NAND4_X1 U7765 ( .A1(n6800), .A2(n6799), .A3(n6798), .A4(n6797), .ZN(n6971)
         );
  INV_X1 U7766 ( .A(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n6983) );
  AOI22_X1 U7767 ( .A1(n7012), .A2(keyinput42), .B1(n6983), .B2(keyinput121), 
        .ZN(n6801) );
  OAI221_X1 U7768 ( .B1(n7012), .B2(keyinput42), .C1(n6983), .C2(keyinput121), 
        .A(n6801), .ZN(n6812) );
  INV_X1 U7769 ( .A(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n6804) );
  AOI22_X1 U7770 ( .A1(n6804), .A2(keyinput36), .B1(keyinput82), .B2(n6803), 
        .ZN(n6802) );
  OAI221_X1 U7771 ( .B1(n6804), .B2(keyinput36), .C1(n6803), .C2(keyinput82), 
        .A(n6802), .ZN(n6811) );
  INV_X1 U7772 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n6806) );
  AOI22_X1 U7773 ( .A1(n3419), .A2(keyinput111), .B1(keyinput7), .B2(n6806), 
        .ZN(n6805) );
  OAI221_X1 U7774 ( .B1(n3419), .B2(keyinput111), .C1(n6806), .C2(keyinput7), 
        .A(n6805), .ZN(n6810) );
  AOI22_X1 U7775 ( .A1(n7035), .A2(keyinput54), .B1(keyinput35), .B2(n6808), 
        .ZN(n6807) );
  OAI221_X1 U7776 ( .B1(n7035), .B2(keyinput54), .C1(n6808), .C2(keyinput35), 
        .A(n6807), .ZN(n6809) );
  NOR4_X1 U7777 ( .A1(n6812), .A2(n6811), .A3(n6810), .A4(n6809), .ZN(n6857)
         );
  INV_X1 U7778 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n6815) );
  AOI22_X1 U7779 ( .A1(n6815), .A2(keyinput64), .B1(keyinput6), .B2(n6814), 
        .ZN(n6813) );
  OAI221_X1 U7780 ( .B1(n6815), .B2(keyinput64), .C1(n6814), .C2(keyinput6), 
        .A(n6813), .ZN(n6827) );
  AOI22_X1 U7781 ( .A1(n6818), .A2(keyinput94), .B1(n6817), .B2(keyinput99), 
        .ZN(n6816) );
  OAI221_X1 U7782 ( .B1(n6818), .B2(keyinput94), .C1(n6817), .C2(keyinput99), 
        .A(n6816), .ZN(n6826) );
  INV_X1 U7783 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n6820) );
  INV_X1 U7784 ( .A(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n7008) );
  AOI22_X1 U7785 ( .A1(n6820), .A2(keyinput43), .B1(n7008), .B2(keyinput23), 
        .ZN(n6819) );
  OAI221_X1 U7786 ( .B1(n6820), .B2(keyinput43), .C1(n7008), .C2(keyinput23), 
        .A(n6819), .ZN(n6825) );
  AOI22_X1 U7787 ( .A1(n6823), .A2(keyinput17), .B1(n6822), .B2(keyinput97), 
        .ZN(n6821) );
  OAI221_X1 U7788 ( .B1(n6823), .B2(keyinput17), .C1(n6822), .C2(keyinput97), 
        .A(n6821), .ZN(n6824) );
  NOR4_X1 U7789 ( .A1(n6827), .A2(n6826), .A3(n6825), .A4(n6824), .ZN(n6856)
         );
  INV_X1 U7790 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n6829) );
  AOI22_X1 U7791 ( .A1(n6829), .A2(keyinput119), .B1(keyinput113), .B2(n7010), 
        .ZN(n6828) );
  OAI221_X1 U7792 ( .B1(n6829), .B2(keyinput119), .C1(n7010), .C2(keyinput113), 
        .A(n6828), .ZN(n6839) );
  AOI22_X1 U7793 ( .A1(n7002), .A2(keyinput63), .B1(keyinput123), .B2(n4521), 
        .ZN(n6830) );
  OAI221_X1 U7794 ( .B1(n7002), .B2(keyinput63), .C1(n4521), .C2(keyinput123), 
        .A(n6830), .ZN(n6838) );
  AOI22_X1 U7795 ( .A1(n6833), .A2(keyinput4), .B1(keyinput11), .B2(n6832), 
        .ZN(n6831) );
  OAI221_X1 U7796 ( .B1(n6833), .B2(keyinput4), .C1(n6832), .C2(keyinput11), 
        .A(n6831), .ZN(n6837) );
  INV_X1 U7797 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n6984) );
  NOR4_X1 U7798 ( .A1(n6839), .A2(n6838), .A3(n6837), .A4(n6836), .ZN(n6855)
         );
  INV_X1 U7799 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6842) );
  AOI22_X1 U7800 ( .A1(n6842), .A2(keyinput71), .B1(keyinput33), .B2(n6841), 
        .ZN(n6840) );
  OAI221_X1 U7801 ( .B1(n6842), .B2(keyinput71), .C1(n6841), .C2(keyinput33), 
        .A(n6840), .ZN(n6853) );
  AOI22_X1 U7802 ( .A1(n6844), .A2(keyinput80), .B1(n7011), .B2(keyinput25), 
        .ZN(n6843) );
  OAI221_X1 U7803 ( .B1(n6844), .B2(keyinput80), .C1(n7011), .C2(keyinput25), 
        .A(n6843), .ZN(n6852) );
  AOI22_X1 U7804 ( .A1(n6846), .A2(keyinput98), .B1(n6986), .B2(keyinput58), 
        .ZN(n6845) );
  OAI221_X1 U7805 ( .B1(n6846), .B2(keyinput98), .C1(n6986), .C2(keyinput58), 
        .A(n6845), .ZN(n6851) );
  AOI22_X1 U7806 ( .A1(n6849), .A2(keyinput31), .B1(keyinput24), .B2(n6848), 
        .ZN(n6847) );
  OAI221_X1 U7807 ( .B1(n6849), .B2(keyinput31), .C1(n6848), .C2(keyinput24), 
        .A(n6847), .ZN(n6850) );
  NOR4_X1 U7808 ( .A1(n6853), .A2(n6852), .A3(n6851), .A4(n6850), .ZN(n6854)
         );
  NAND4_X1 U7809 ( .A1(n6857), .A2(n6856), .A3(n6855), .A4(n6854), .ZN(n6970)
         );
  AOI22_X1 U7810 ( .A1(n4691), .A2(keyinput27), .B1(keyinput26), .B2(n6859), 
        .ZN(n6858) );
  OAI221_X1 U7811 ( .B1(n4691), .B2(keyinput27), .C1(n6859), .C2(keyinput26), 
        .A(n6858), .ZN(n6869) );
  AOI22_X1 U7812 ( .A1(n6861), .A2(keyinput91), .B1(n4673), .B2(keyinput100), 
        .ZN(n6860) );
  OAI221_X1 U7813 ( .B1(n6861), .B2(keyinput91), .C1(n4673), .C2(keyinput100), 
        .A(n6860), .ZN(n6868) );
  INV_X1 U7814 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6864) );
  AOI22_X1 U7815 ( .A1(n6864), .A2(keyinput89), .B1(keyinput74), .B2(n6863), 
        .ZN(n6862) );
  OAI221_X1 U7816 ( .B1(n6864), .B2(keyinput89), .C1(n6863), .C2(keyinput74), 
        .A(n6862), .ZN(n6867) );
  AOI22_X1 U7817 ( .A1(n3569), .A2(keyinput75), .B1(n6974), .B2(keyinput112), 
        .ZN(n6865) );
  OAI221_X1 U7818 ( .B1(n3569), .B2(keyinput75), .C1(n6974), .C2(keyinput112), 
        .A(n6865), .ZN(n6866) );
  NOR4_X1 U7819 ( .A1(n6869), .A2(n6868), .A3(n6867), .A4(n6866), .ZN(n6910)
         );
  INV_X1 U7820 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n7024) );
  AOI22_X1 U7821 ( .A1(n7024), .A2(keyinput28), .B1(keyinput78), .B2(n6871), 
        .ZN(n6870) );
  OAI221_X1 U7822 ( .B1(n7024), .B2(keyinput28), .C1(n6871), .C2(keyinput78), 
        .A(n6870), .ZN(n6881) );
  AOI22_X1 U7823 ( .A1(n6874), .A2(keyinput105), .B1(keyinput103), .B2(n6873), 
        .ZN(n6872) );
  OAI221_X1 U7824 ( .B1(n6874), .B2(keyinput105), .C1(n6873), .C2(keyinput103), 
        .A(n6872), .ZN(n6880) );
  AOI22_X1 U7825 ( .A1(n7013), .A2(keyinput1), .B1(n6981), .B2(keyinput37), 
        .ZN(n6875) );
  OAI221_X1 U7826 ( .B1(n7013), .B2(keyinput1), .C1(n6981), .C2(keyinput37), 
        .A(n6875), .ZN(n6879) );
  INV_X1 U7827 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n7021) );
  INV_X1 U7828 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n6877) );
  AOI22_X1 U7829 ( .A1(n7021), .A2(keyinput66), .B1(keyinput87), .B2(n6877), 
        .ZN(n6876) );
  OAI221_X1 U7830 ( .B1(n7021), .B2(keyinput66), .C1(n6877), .C2(keyinput87), 
        .A(n6876), .ZN(n6878) );
  NOR4_X1 U7831 ( .A1(n6881), .A2(n6880), .A3(n6879), .A4(n6878), .ZN(n6909)
         );
  INV_X1 U7832 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n6884) );
  AOI22_X1 U7833 ( .A1(n6884), .A2(keyinput117), .B1(keyinput15), .B2(n6883), 
        .ZN(n6882) );
  OAI221_X1 U7834 ( .B1(n6884), .B2(keyinput117), .C1(n6883), .C2(keyinput15), 
        .A(n6882), .ZN(n6894) );
  AOI22_X1 U7835 ( .A1(n6886), .A2(keyinput90), .B1(n4685), .B2(keyinput44), 
        .ZN(n6885) );
  OAI221_X1 U7836 ( .B1(n6886), .B2(keyinput90), .C1(n4685), .C2(keyinput44), 
        .A(n6885), .ZN(n6893) );
  AOI22_X1 U7837 ( .A1(n6888), .A2(keyinput67), .B1(n5325), .B2(keyinput69), 
        .ZN(n6887) );
  OAI221_X1 U7838 ( .B1(n6888), .B2(keyinput67), .C1(n5325), .C2(keyinput69), 
        .A(n6887), .ZN(n6892) );
  INV_X1 U7839 ( .A(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n6979) );
  AOI22_X1 U7840 ( .A1(n6890), .A2(keyinput62), .B1(n6979), .B2(keyinput85), 
        .ZN(n6889) );
  OAI221_X1 U7841 ( .B1(n6890), .B2(keyinput62), .C1(n6979), .C2(keyinput85), 
        .A(n6889), .ZN(n6891) );
  NOR4_X1 U7842 ( .A1(n6894), .A2(n6893), .A3(n6892), .A4(n6891), .ZN(n6908)
         );
  AOI22_X1 U7843 ( .A1(n7023), .A2(keyinput8), .B1(keyinput70), .B2(n4453), 
        .ZN(n6895) );
  OAI221_X1 U7844 ( .B1(n7023), .B2(keyinput8), .C1(n4453), .C2(keyinput70), 
        .A(n6895), .ZN(n6906) );
  AOI22_X1 U7845 ( .A1(n6898), .A2(keyinput60), .B1(n6897), .B2(keyinput104), 
        .ZN(n6896) );
  OAI221_X1 U7846 ( .B1(n6898), .B2(keyinput60), .C1(n6897), .C2(keyinput104), 
        .A(n6896), .ZN(n6905) );
  AOI22_X1 U7847 ( .A1(n6901), .A2(keyinput52), .B1(n6900), .B2(keyinput56), 
        .ZN(n6899) );
  OAI221_X1 U7848 ( .B1(n6901), .B2(keyinput52), .C1(n6900), .C2(keyinput56), 
        .A(n6899), .ZN(n6904) );
  AOI22_X1 U7849 ( .A1(n5755), .A2(keyinput46), .B1(keyinput95), .B2(n4489), 
        .ZN(n6902) );
  OAI221_X1 U7850 ( .B1(n5755), .B2(keyinput46), .C1(n4489), .C2(keyinput95), 
        .A(n6902), .ZN(n6903) );
  NOR4_X1 U7851 ( .A1(n6906), .A2(n6905), .A3(n6904), .A4(n6903), .ZN(n6907)
         );
  NAND4_X1 U7852 ( .A1(n6910), .A2(n6909), .A3(n6908), .A4(n6907), .ZN(n6969)
         );
  AOI22_X1 U7853 ( .A1(n6913), .A2(keyinput51), .B1(keyinput92), .B2(n6912), 
        .ZN(n6911) );
  OAI221_X1 U7854 ( .B1(n6913), .B2(keyinput51), .C1(n6912), .C2(keyinput92), 
        .A(n6911), .ZN(n6924) );
  INV_X1 U7855 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n6982) );
  INV_X1 U7856 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n6915) );
  AOI22_X1 U7857 ( .A1(n6982), .A2(keyinput73), .B1(n6915), .B2(keyinput109), 
        .ZN(n6914) );
  OAI221_X1 U7858 ( .B1(n6982), .B2(keyinput73), .C1(n6915), .C2(keyinput109), 
        .A(n6914), .ZN(n6923) );
  AOI22_X1 U7859 ( .A1(n6918), .A2(keyinput81), .B1(keyinput0), .B2(n6917), 
        .ZN(n6916) );
  OAI221_X1 U7860 ( .B1(n6918), .B2(keyinput81), .C1(n6917), .C2(keyinput0), 
        .A(n6916), .ZN(n6922) );
  INV_X1 U7861 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n7019) );
  AOI22_X1 U7862 ( .A1(n7019), .A2(keyinput9), .B1(keyinput122), .B2(n6920), 
        .ZN(n6919) );
  OAI221_X1 U7863 ( .B1(n7019), .B2(keyinput9), .C1(n6920), .C2(keyinput122), 
        .A(n6919), .ZN(n6921) );
  NOR4_X1 U7864 ( .A1(n6924), .A2(n6923), .A3(n6922), .A4(n6921), .ZN(n6967)
         );
  INV_X1 U7865 ( .A(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n6926) );
  AOI22_X1 U7866 ( .A1(n6927), .A2(keyinput20), .B1(n6926), .B2(keyinput110), 
        .ZN(n6925) );
  OAI221_X1 U7867 ( .B1(n6927), .B2(keyinput20), .C1(n6926), .C2(keyinput110), 
        .A(n6925), .ZN(n6939) );
  INV_X1 U7868 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n6930) );
  AOI22_X1 U7869 ( .A1(n6930), .A2(keyinput72), .B1(keyinput83), .B2(n6929), 
        .ZN(n6928) );
  OAI221_X1 U7870 ( .B1(n6930), .B2(keyinput72), .C1(n6929), .C2(keyinput83), 
        .A(n6928), .ZN(n6938) );
  INV_X1 U7871 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n6978) );
  AOI22_X1 U7872 ( .A1(n6978), .A2(keyinput34), .B1(keyinput29), .B2(n6932), 
        .ZN(n6931) );
  OAI221_X1 U7873 ( .B1(n6978), .B2(keyinput34), .C1(n6932), .C2(keyinput29), 
        .A(n6931), .ZN(n6937) );
  INV_X1 U7874 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n6934) );
  AOI22_X1 U7875 ( .A1(n6935), .A2(keyinput101), .B1(keyinput68), .B2(n6934), 
        .ZN(n6933) );
  OAI221_X1 U7876 ( .B1(n6935), .B2(keyinput101), .C1(n6934), .C2(keyinput68), 
        .A(n6933), .ZN(n6936) );
  NOR4_X1 U7877 ( .A1(n6939), .A2(n6938), .A3(n6937), .A4(n6936), .ZN(n6966)
         );
  INV_X1 U7878 ( .A(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n6941) );
  AOI22_X1 U7879 ( .A1(n6941), .A2(keyinput21), .B1(n6980), .B2(keyinput120), 
        .ZN(n6940) );
  OAI221_X1 U7880 ( .B1(n6941), .B2(keyinput21), .C1(n6980), .C2(keyinput120), 
        .A(n6940), .ZN(n6951) );
  AOI22_X1 U7881 ( .A1(n6944), .A2(keyinput22), .B1(n6943), .B2(keyinput77), 
        .ZN(n6942) );
  OAI221_X1 U7882 ( .B1(n6944), .B2(keyinput22), .C1(n6943), .C2(keyinput77), 
        .A(n6942), .ZN(n6950) );
  AOI22_X1 U7883 ( .A1(n6946), .A2(keyinput61), .B1(n4807), .B2(keyinput102), 
        .ZN(n6945) );
  OAI221_X1 U7884 ( .B1(n6946), .B2(keyinput61), .C1(n4807), .C2(keyinput102), 
        .A(n6945), .ZN(n6949) );
  INV_X1 U7885 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n7020) );
  AOI22_X1 U7886 ( .A1(n5619), .A2(keyinput86), .B1(n7020), .B2(keyinput30), 
        .ZN(n6947) );
  OAI221_X1 U7887 ( .B1(n5619), .B2(keyinput86), .C1(n7020), .C2(keyinput30), 
        .A(n6947), .ZN(n6948) );
  NOR4_X1 U7888 ( .A1(n6951), .A2(n6950), .A3(n6949), .A4(n6948), .ZN(n6965)
         );
  AOI22_X1 U7889 ( .A1(n6953), .A2(keyinput32), .B1(n6977), .B2(keyinput2), 
        .ZN(n6952) );
  OAI221_X1 U7890 ( .B1(n6953), .B2(keyinput32), .C1(n6977), .C2(keyinput2), 
        .A(n6952), .ZN(n6963) );
  INV_X1 U7891 ( .A(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n6985) );
  AOI22_X1 U7892 ( .A1(n6985), .A2(keyinput47), .B1(keyinput53), .B2(n6955), 
        .ZN(n6954) );
  OAI221_X1 U7893 ( .B1(n6985), .B2(keyinput47), .C1(n6955), .C2(keyinput53), 
        .A(n6954), .ZN(n6962) );
  AOI22_X1 U7894 ( .A1(n4487), .A2(keyinput125), .B1(n6957), .B2(keyinput88), 
        .ZN(n6956) );
  OAI221_X1 U7895 ( .B1(n4487), .B2(keyinput125), .C1(n6957), .C2(keyinput88), 
        .A(n6956), .ZN(n6961) );
  INV_X1 U7896 ( .A(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n7025) );
  AOI22_X1 U7897 ( .A1(n6959), .A2(keyinput65), .B1(n7025), .B2(keyinput48), 
        .ZN(n6958) );
  OAI221_X1 U7898 ( .B1(n6959), .B2(keyinput65), .C1(n7025), .C2(keyinput48), 
        .A(n6958), .ZN(n6960) );
  NOR4_X1 U7899 ( .A1(n6963), .A2(n6962), .A3(n6961), .A4(n6960), .ZN(n6964)
         );
  NAND4_X1 U7900 ( .A1(n6967), .A2(n6966), .A3(n6965), .A4(n6964), .ZN(n6968)
         );
  NOR4_X1 U7901 ( .A1(n6971), .A2(n6970), .A3(n6969), .A4(n6968), .ZN(n6972)
         );
  XNOR2_X1 U7902 ( .A(n6973), .B(n6972), .ZN(n7049) );
  NOR4_X1 U7903 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n6976) );
  NAND4_X1 U7904 ( .A1(n6976), .A2(n6975), .A3(n6974), .A4(n5619), .ZN(n6997)
         );
  NAND4_X1 U7905 ( .A1(n6980), .A2(n6979), .A3(n6978), .A4(n6977), .ZN(n6996)
         );
  NAND4_X1 U7906 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .A3(PHYADDRPOINTER_REG_2__SCAN_IN), 
        .A4(n6981), .ZN(n6995) );
  NOR4_X1 U7907 ( .A1(INSTQUEUE_REG_2__7__SCAN_IN), .A2(
        INSTQUEUE_REG_15__7__SCAN_IN), .A3(n6983), .A4(n6982), .ZN(n6993) );
  NOR4_X1 U7908 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(
        INSTQUEUE_REG_8__7__SCAN_IN), .A3(n6985), .A4(n6984), .ZN(n6992) );
  NOR4_X1 U7909 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(
        INSTQUEUE_REG_12__7__SCAN_IN), .A3(EAX_REG_14__SCAN_IN), .A4(n6986), 
        .ZN(n6987) );
  NAND2_X1 U7910 ( .A1(n6988), .A2(n6987), .ZN(n6989) );
  NOR4_X1 U7911 ( .A1(n6990), .A2(n6989), .A3(INSTQUEUE_REG_15__6__SCAN_IN), 
        .A4(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6991) );
  NAND3_X1 U7912 ( .A1(n6993), .A2(n6992), .A3(n6991), .ZN(n6994) );
  NOR4_X1 U7913 ( .A1(n6997), .A2(n6996), .A3(n6995), .A4(n6994), .ZN(n7047)
         );
  NAND4_X1 U7914 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        BE_N_REG_3__SCAN_IN), .A3(UWORD_REG_11__SCAN_IN), .A4(
        LWORD_REG_3__SCAN_IN), .ZN(n7001) );
  NAND4_X1 U7915 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_27__SCAN_IN), .A4(
        BYTEENABLE_REG_0__SCAN_IN), .ZN(n7000) );
  NAND4_X1 U7916 ( .A1(EBX_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_13__SCAN_IN), .A3(REIP_REG_3__SCAN_IN), .A4(
        DATAI_16_), .ZN(n6999) );
  NAND4_X1 U7917 ( .A1(DATAI_18_), .A2(DATAO_REG_7__SCAN_IN), .A3(
        DATAO_REG_21__SCAN_IN), .A4(UWORD_REG_5__SCAN_IN), .ZN(n6998) );
  NOR4_X1 U7918 ( .A1(n7001), .A2(n7000), .A3(n6999), .A4(n6998), .ZN(n7046)
         );
  NAND4_X1 U7919 ( .A1(EBX_REG_19__SCAN_IN), .A2(DATAI_30_), .A3(DATAI_27_), 
        .A4(DATAI_21_), .ZN(n7007) );
  NAND4_X1 U7920 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .A3(
        DATAI_31_), .A4(MEMORYFETCH_REG_SCAN_IN), .ZN(n7006) );
  NAND4_X1 U7921 ( .A1(DATAO_REG_29__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), 
        .A3(DATAWIDTH_REG_31__SCAN_IN), .A4(DATAWIDTH_REG_22__SCAN_IN), .ZN(
        n7005) );
  NAND4_X1 U7922 ( .A1(DATAO_REG_12__SCAN_IN), .A2(DATAO_REG_26__SCAN_IN), 
        .A3(n7003), .A4(n7002), .ZN(n7004) );
  NOR4_X1 U7923 ( .A1(n7007), .A2(n7006), .A3(n7005), .A4(n7004), .ZN(n7045)
         );
  NOR4_X1 U7924 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(
        INSTQUEUE_REG_0__0__SCAN_IN), .A3(INSTQUEUE_REG_9__1__SCAN_IN), .A4(
        n7008), .ZN(n7018) );
  NOR4_X1 U7925 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(
        INSTQUEUE_REG_11__1__SCAN_IN), .A3(n7009), .A4(n4968), .ZN(n7017) );
  NOR4_X1 U7926 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n7012), .A3(n7011), 
        .A4(n7010), .ZN(n7016) );
  NOR4_X1 U7927 ( .A1(EAX_REG_7__SCAN_IN), .A2(EAX_REG_2__SCAN_IN), .A3(n7014), 
        .A4(n7013), .ZN(n7015) );
  NAND4_X1 U7928 ( .A1(n7018), .A2(n7017), .A3(n7016), .A4(n7015), .ZN(n7043)
         );
  NOR4_X1 U7929 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n7021), .A3(n7020), 
        .A4(n7019), .ZN(n7029) );
  NOR4_X1 U7930 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(
        INSTQUEUE_REG_5__5__SCAN_IN), .A3(INSTQUEUE_REG_13__5__SCAN_IN), .A4(
        n7022), .ZN(n7028) );
  NOR4_X1 U7931 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(
        INSTQUEUE_REG_4__2__SCAN_IN), .A3(INSTQUEUE_REG_10__2__SCAN_IN), .A4(
        n7023), .ZN(n7027) );
  NOR4_X1 U7932 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(
        INSTQUEUE_REG_3__3__SCAN_IN), .A3(n7025), .A4(n7024), .ZN(n7026) );
  NAND4_X1 U7933 ( .A1(n7029), .A2(n7028), .A3(n7027), .A4(n7026), .ZN(n7042)
         );
  NOR4_X1 U7934 ( .A1(EAX_REG_22__SCAN_IN), .A2(DATAI_25_), .A3(DATAI_24_), 
        .A4(DATAI_4_), .ZN(n7034) );
  NOR4_X1 U7935 ( .A1(EBX_REG_8__SCAN_IN), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .A3(REIP_REG_1__SCAN_IN), .A4(REIP_REG_12__SCAN_IN), .ZN(n7033) );
  NOR4_X1 U7936 ( .A1(EAX_REG_30__SCAN_IN), .A2(DATAI_13_), .A3(DATAI_11_), 
        .A4(n7030), .ZN(n7032) );
  NAND4_X1 U7937 ( .A1(n7034), .A2(n7033), .A3(n7032), .A4(n7031), .ZN(n7041)
         );
  NOR4_X1 U7938 ( .A1(DATAO_REG_20__SCAN_IN), .A2(ADDRESS_REG_26__SCAN_IN), 
        .A3(ADDRESS_REG_25__SCAN_IN), .A4(DATAO_REG_3__SCAN_IN), .ZN(n7039) );
  NOR4_X1 U7939 ( .A1(DATAO_REG_31__SCAN_IN), .A2(LWORD_REG_15__SCAN_IN), .A3(
        DATAO_REG_18__SCAN_IN), .A4(n7035), .ZN(n7038) );
  NOR4_X1 U7940 ( .A1(REIP_REG_2__SCAN_IN), .A2(LWORD_REG_4__SCAN_IN), .A3(
        LWORD_REG_2__SCAN_IN), .A4(DATAO_REG_5__SCAN_IN), .ZN(n7037) );
  NOR4_X1 U7941 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        ADDRESS_REG_27__SCAN_IN), .A3(BE_N_REG_1__SCAN_IN), .A4(
        BE_N_REG_2__SCAN_IN), .ZN(n7036) );
  NAND4_X1 U7942 ( .A1(n7039), .A2(n7038), .A3(n7037), .A4(n7036), .ZN(n7040)
         );
  NOR4_X1 U7943 ( .A1(n7043), .A2(n7042), .A3(n7041), .A4(n7040), .ZN(n7044)
         );
  NAND4_X1 U7944 ( .A1(n7047), .A2(n7046), .A3(n7045), .A4(n7044), .ZN(n7048)
         );
  XNOR2_X1 U7945 ( .A(n7049), .B(n7048), .ZN(U2877) );
  AND2_X1 U3594 ( .A1(n4627), .A2(n5551), .ZN(n3352) );
  OR2_X1 U4168 ( .A1(n3197), .A2(n3196), .ZN(n4564) );
  CLKBUF_X1 U3584 ( .A(n4161), .Z(n4146) );
  CLKBUF_X1 U3604 ( .A(n3480), .Z(n4141) );
  AOI21_X1 U3609 ( .B1(n5763), .B2(n6609), .A(n3383), .ZN(n3440) );
  AND4_X1 U3625 ( .A1(n3268), .A2(n3267), .A3(n3266), .A4(n3265), .ZN(n3269)
         );
  CLKBUF_X1 U3647 ( .A(n3467), .Z(n4631) );
  CLKBUF_X1 U3667 ( .A(n5858), .Z(n5897) );
  CLKBUF_X1 U4070 ( .A(n3449), .Z(n5297) );
  CLKBUF_X1 U4234 ( .A(n3960), .Z(n4357) );
endmodule

