

module b14_C_AntiSAT_k_128_4 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795;

  INV_X1 U2293 ( .A(n2710), .ZN(n2880) );
  NOR2_X1 U2294 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2267)
         );
  INV_X1 U2295 ( .A(n2710), .ZN(n2731) );
  INV_X2 U2296 ( .A(n2874), .ZN(n2893) );
  INV_X1 U2297 ( .A(n2579), .ZN(n2456) );
  MUX2_X1 U2298 ( .A(n2279), .B(n2278), .S(n2255), .Z(n2051) );
  NAND2_X1 U2299 ( .A1(n2288), .A2(n2971), .ZN(n2535) );
  AND2_X1 U2300 ( .A1(n4366), .A2(n4365), .ZN(n4368) );
  NAND2_X2 U2301 ( .A1(n2639), .A2(n3786), .ZN(n3097) );
  XNOR2_X2 U2302 ( .A(n2566), .B(n2565), .ZN(n2639) );
  OAI21_X1 U2303 ( .B1(n3555), .B2(n2182), .A(n2180), .ZN(n2818) );
  OAI22_X1 U2304 ( .A1(n4668), .A2(n4664), .B1(REG2_REG_13__SCAN_IN), .B2(
        n4759), .ZN(n4053) );
  NAND2_X1 U2305 ( .A1(n4656), .A2(REG2_REG_12__SCAN_IN), .ZN(n4655) );
  XNOR2_X1 U2306 ( .A(n4051), .B(n2151), .ZN(n4656) );
  NAND2_X1 U2307 ( .A1(n4645), .A2(n4050), .ZN(n4051) );
  INV_X1 U2308 ( .A(n4110), .ZN(n2052) );
  XNOR2_X1 U2309 ( .A(n4048), .B(n2150), .ZN(n4634) );
  AND2_X1 U2310 ( .A1(n3258), .A2(n2087), .ZN(n4366) );
  INV_X2 U2311 ( .A(n3364), .ZN(n3626) );
  NAND2_X2 U2312 ( .A1(n3097), .A2(n2913), .ZN(n2874) );
  NAND3_X1 U2313 ( .A1(n4607), .A2(n2968), .A3(n4608), .ZN(n2937) );
  AND2_X2 U2314 ( .A1(n2287), .A2(n2289), .ZN(n2303) );
  INV_X1 U2315 ( .A(n2487), .ZN(n2489) );
  OR2_X1 U2316 ( .A1(n2476), .A2(n2075), .ZN(n2487) );
  AND2_X1 U2317 ( .A1(n2245), .A2(n2267), .ZN(n2139) );
  AND2_X1 U2318 ( .A1(n2323), .A2(n2265), .ZN(n2053) );
  NOR2_X1 U2319 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2297)
         );
  INV_X1 U2320 ( .A(IR_REG_5__SCAN_IN), .ZN(n2247) );
  AOI21_X2 U2321 ( .B1(n3382), .B2(n2871), .A(n2870), .ZN(n3506) );
  NAND2_X4 U2322 ( .A1(n2639), .A2(n2203), .ZN(n2710) );
  XNOR2_X1 U2323 ( .A(n2713), .B(n2874), .ZN(n2718) );
  NOR2_X1 U2324 ( .A1(n2204), .A2(n2921), .ZN(n2203) );
  INV_X1 U2325 ( .A(n2113), .ZN(n2112) );
  INV_X1 U2326 ( .A(n3657), .ZN(n2253) );
  INV_X1 U2327 ( .A(n2971), .ZN(n2289) );
  INV_X1 U2328 ( .A(n3741), .ZN(n2118) );
  INV_X1 U2329 ( .A(n4494), .ZN(n2587) );
  AND2_X1 U2330 ( .A1(n2275), .A2(n2274), .ZN(n2149) );
  NOR2_X1 U2331 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2275)
         );
  INV_X1 U2332 ( .A(IR_REG_22__SCAN_IN), .ZN(n2274) );
  INV_X1 U2333 ( .A(n2813), .ZN(n2816) );
  NOR2_X1 U2334 ( .A1(n3042), .A2(n3043), .ZN(n3041) );
  NAND2_X1 U2335 ( .A1(n4643), .A2(n4644), .ZN(n4642) );
  XNOR2_X1 U2336 ( .A(n4072), .B(n4054), .ZN(n4038) );
  NOR2_X1 U2337 ( .A1(n2163), .A2(n4709), .ZN(n4708) );
  INV_X1 U2338 ( .A(n2214), .ZN(n2213) );
  AOI22_X1 U2339 ( .A1(n4145), .A2(n2540), .B1(n4399), .B2(n4147), .ZN(n4126)
         );
  NAND2_X1 U2340 ( .A1(n4198), .A2(n2514), .ZN(n2137) );
  OAI21_X1 U2341 ( .B1(n4286), .B2(n2099), .A(n2097), .ZN(n4253) );
  INV_X1 U2342 ( .A(n2100), .ZN(n2099) );
  AOI21_X1 U2343 ( .B1(n2100), .B2(n2102), .A(n2098), .ZN(n2097) );
  INV_X1 U2344 ( .A(n4505), .ZN(n4529) );
  OR2_X1 U2345 ( .A1(n3088), .A2(n4609), .ZN(n3113) );
  AND2_X1 U2346 ( .A1(n2259), .A2(n2258), .ZN(n2257) );
  INV_X1 U2347 ( .A(IR_REG_21__SCAN_IN), .ZN(n2258) );
  AND2_X1 U2348 ( .A1(n3348), .A2(n2189), .ZN(n2188) );
  NOR2_X1 U2349 ( .A1(n2169), .A2(n3543), .ZN(n2168) );
  INV_X1 U2350 ( .A(n2170), .ZN(n2169) );
  INV_X1 U2351 ( .A(n3541), .ZN(n2171) );
  INV_X1 U2352 ( .A(n2937), .ZN(n2204) );
  OR2_X1 U2353 ( .A1(n2176), .A2(n2173), .ZN(n2172) );
  INV_X1 U2354 ( .A(n2179), .ZN(n2173) );
  AND2_X1 U2355 ( .A1(n3419), .A2(n2177), .ZN(n2176) );
  NAND2_X1 U2356 ( .A1(n3586), .A2(n3587), .ZN(n2177) );
  AND2_X1 U2357 ( .A1(n2092), .A2(n2091), .ZN(n2996) );
  NAND2_X1 U2358 ( .A1(n3004), .A2(REG1_REG_5__SCAN_IN), .ZN(n2091) );
  INV_X1 U2359 ( .A(n3660), .ZN(n2250) );
  INV_X1 U2360 ( .A(n2514), .ZN(n2133) );
  OR2_X1 U2361 ( .A1(n2390), .A2(n2389), .ZN(n2403) );
  NOR2_X1 U2362 ( .A1(n2403), .A2(n3578), .ZN(n2409) );
  INV_X1 U2363 ( .A(n2123), .ZN(n2121) );
  AND2_X1 U2364 ( .A1(n3692), .A2(n3691), .ZN(n2227) );
  NAND2_X1 U2365 ( .A1(n2125), .A2(n2124), .ZN(n2123) );
  NAND2_X1 U2366 ( .A1(n2347), .A2(n2126), .ZN(n2122) );
  NOR2_X1 U2367 ( .A1(n2355), .A2(n2127), .ZN(n2126) );
  INV_X1 U2368 ( .A(n2346), .ZN(n2127) );
  AND2_X1 U2369 ( .A1(n2269), .A2(n2268), .ZN(n2260) );
  NOR2_X1 U2370 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2269)
         );
  OR2_X1 U2371 ( .A1(n3599), .A2(n3598), .ZN(n2189) );
  NAND3_X1 U2372 ( .A1(n3484), .A2(n2725), .A3(n2191), .ZN(n2190) );
  NAND2_X1 U2373 ( .A1(n3599), .A2(n3598), .ZN(n2191) );
  AOI21_X1 U2374 ( .B1(n3983), .B2(n2731), .A(n2675), .ZN(n2680) );
  OR2_X1 U2375 ( .A1(n2533), .A2(n2532), .ZN(n2542) );
  XNOR2_X1 U2376 ( .A(n2671), .B(n2874), .ZN(n2684) );
  OAI22_X1 U2377 ( .A1(n3499), .A2(n2826), .B1(n2825), .B2(n3496), .ZN(n3590)
         );
  NOR2_X1 U2378 ( .A1(n3041), .A2(n2068), .ZN(n2993) );
  OR2_X1 U2379 ( .A1(n3030), .A2(n3029), .ZN(n2092) );
  XNOR2_X1 U2380 ( .A(n2996), .B(n3017), .ZN(n3014) );
  AOI21_X1 U2381 ( .B1(n3004), .B2(REG2_REG_5__SCAN_IN), .A(n3031), .ZN(n3005)
         );
  OAI21_X1 U2382 ( .B1(n3015), .B2(n2058), .A(n2093), .ZN(n4027) );
  INV_X1 U2383 ( .A(n2094), .ZN(n2093) );
  OAI21_X1 U2384 ( .B1(n2207), .B2(n2058), .A(n2205), .ZN(n2094) );
  NAND2_X1 U2385 ( .A1(n3058), .A2(REG1_REG_7__SCAN_IN), .ZN(n2205) );
  OAI22_X1 U2386 ( .A1(n4046), .A2(n4721), .B1(n4045), .B2(n4044), .ZN(n4625)
         );
  NAND2_X1 U2387 ( .A1(n4625), .A2(n4626), .ZN(n4624) );
  NAND2_X1 U2388 ( .A1(n4642), .A2(n4034), .ZN(n4035) );
  NAND2_X1 U2389 ( .A1(n4672), .A2(n4037), .ZN(n4072) );
  NAND2_X1 U2390 ( .A1(n4038), .A2(REG1_REG_14__SCAN_IN), .ZN(n4073) );
  NOR2_X1 U2391 ( .A1(n4678), .A2(n2156), .ZN(n4065) );
  AND2_X1 U2392 ( .A1(n4071), .A2(REG2_REG_15__SCAN_IN), .ZN(n2156) );
  NOR2_X1 U2393 ( .A1(n2214), .A2(n2212), .ZN(n2211) );
  INV_X1 U2394 ( .A(n4702), .ZN(n2212) );
  NAND2_X1 U2395 ( .A1(n2108), .A2(n2107), .ZN(n2649) );
  AOI21_X1 U2396 ( .B1(n2110), .B2(n2112), .A(n2076), .ZN(n2107) );
  NAND2_X1 U2397 ( .A1(n4126), .A2(n2110), .ZN(n2108) );
  AND2_X1 U2398 ( .A1(n2118), .A2(n2549), .ZN(n2114) );
  NAND2_X1 U2399 ( .A1(n2071), .A2(n2118), .ZN(n2113) );
  NAND2_X1 U2400 ( .A1(n4140), .A2(n3675), .ZN(n2217) );
  AOI22_X1 U2401 ( .A1(n4156), .A2(n2531), .B1(n3780), .B2(n4188), .ZN(n4145)
         );
  NOR2_X1 U2402 ( .A1(n4176), .A2(n2136), .ZN(n2135) );
  INV_X1 U2403 ( .A(n2515), .ZN(n2136) );
  AND2_X1 U2404 ( .A1(n4161), .A2(n2601), .ZN(n4176) );
  OAI211_X1 U2405 ( .C1(n4231), .C2(n4214), .A(n3750), .B(n4215), .ZN(n2509)
         );
  NAND2_X1 U2406 ( .A1(n2103), .A2(n2061), .ZN(n2100) );
  NAND3_X1 U2407 ( .A1(n2455), .A2(n2454), .A3(n2453), .ZN(n4286) );
  OR2_X1 U2408 ( .A1(n3268), .A2(n2443), .ZN(n2455) );
  NAND2_X1 U2409 ( .A1(n2106), .A2(n2105), .ZN(n4288) );
  INV_X1 U2410 ( .A(n4286), .ZN(n2106) );
  AOI21_X1 U2411 ( .B1(n2239), .B2(n2241), .A(n2083), .ZN(n2237) );
  NAND2_X1 U2412 ( .A1(n2238), .A2(n3709), .ZN(n4331) );
  NAND2_X1 U2413 ( .A1(n3267), .A2(n2242), .ZN(n2238) );
  OAI21_X1 U2414 ( .B1(n3267), .B2(n2241), .A(n2239), .ZN(n4332) );
  NAND2_X1 U2415 ( .A1(n3267), .A2(n3707), .ZN(n3292) );
  NAND2_X1 U2416 ( .A1(n3701), .A2(n3775), .ZN(n2225) );
  NAND2_X1 U2417 ( .A1(n2227), .A2(n3775), .ZN(n2226) );
  OR2_X1 U2418 ( .A1(n2375), .A2(n3961), .ZN(n2390) );
  AND2_X1 U2419 ( .A1(n3692), .A2(n4513), .ZN(n3777) );
  NOR2_X1 U2420 ( .A1(n2584), .A2(n2229), .ZN(n2233) );
  OAI21_X1 U2421 ( .B1(n3689), .B2(n2232), .A(n2082), .ZN(n2231) );
  NAND2_X1 U2422 ( .A1(n3686), .A2(n3698), .ZN(n2229) );
  NOR2_X1 U2423 ( .A1(n2584), .A2(n2228), .ZN(n2234) );
  INV_X1 U2424 ( .A(n3686), .ZN(n2228) );
  INV_X1 U2425 ( .A(n3521), .ZN(n3211) );
  AND2_X1 U2426 ( .A1(n3687), .A2(n3689), .ZN(n3765) );
  INV_X1 U2427 ( .A(n4130), .ZN(n4399) );
  AND2_X1 U2428 ( .A1(n2639), .A2(n3082), .ZN(n4258) );
  AND2_X1 U2429 ( .A1(n3672), .A2(n2607), .ZN(n4505) );
  MUX2_X1 U2430 ( .A(n4615), .B(DATAI_2_), .S(n2310), .Z(n3151) );
  AND3_X1 U2431 ( .A1(n2636), .A2(n2635), .A3(n2899), .ZN(n2644) );
  NAND2_X1 U2432 ( .A1(n2618), .A2(n4607), .ZN(n2973) );
  AND2_X1 U2433 ( .A1(n2937), .A2(n4750), .ZN(n3090) );
  AND2_X1 U2434 ( .A1(n2072), .A2(n2149), .ZN(n2138) );
  INV_X1 U2435 ( .A(IR_REG_25__SCAN_IN), .ZN(n2256) );
  INV_X1 U2436 ( .A(IR_REG_28__SCAN_IN), .ZN(n2575) );
  AND2_X1 U2437 ( .A1(n2569), .A2(n2274), .ZN(n2613) );
  INV_X1 U2438 ( .A(IR_REG_23__SCAN_IN), .ZN(n2620) );
  AND2_X1 U2439 ( .A1(n2273), .A2(n2260), .ZN(n2259) );
  AND4_X1 U2440 ( .A1(n2474), .A2(n2272), .A3(n2271), .A4(n2270), .ZN(n2273)
         );
  NOR2_X1 U2441 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2272)
         );
  NOR2_X1 U2442 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2271)
         );
  INV_X1 U2443 ( .A(IR_REG_20__SCAN_IN), .ZN(n2565) );
  NAND2_X1 U2444 ( .A1(n2564), .A2(IR_REG_31__SCAN_IN), .ZN(n2566) );
  NAND2_X1 U2445 ( .A1(n2501), .A2(n2500), .ZN(n2564) );
  NAND2_X1 U2446 ( .A1(n2489), .A2(n2488), .ZN(n2499) );
  XNOR2_X1 U2447 ( .A(n2477), .B(IR_REG_17__SCAN_IN), .ZN(n4080) );
  XNOR2_X1 U2448 ( .A(n2324), .B(IR_REG_3__SCAN_IN), .ZN(n3001) );
  NAND2_X1 U2449 ( .A1(n2194), .A2(n2192), .ZN(n2935) );
  NOR2_X1 U2450 ( .A1(n2193), .A2(n3359), .ZN(n2192) );
  INV_X1 U2451 ( .A(n2195), .ZN(n2193) );
  INV_X1 U2452 ( .A(n3517), .ZN(n3624) );
  NAND4_X1 U2453 ( .A1(n2338), .A2(n2337), .A3(n2336), .A4(n2335), .ZN(n3603)
         );
  NAND4_X1 U2454 ( .A1(n2322), .A2(n2321), .A3(n2320), .A4(n2319), .ZN(n3806)
         );
  XNOR2_X1 U2455 ( .A(n4035), .B(n2151), .ZN(n4661) );
  NAND2_X1 U2456 ( .A1(n4661), .A2(REG1_REG_12__SCAN_IN), .ZN(n4660) );
  NAND2_X1 U2457 ( .A1(n4673), .A2(n4674), .ZN(n4672) );
  XNOR2_X1 U2458 ( .A(n4065), .B(n4076), .ZN(n4690) );
  NAND2_X1 U2459 ( .A1(n4690), .A2(n4688), .ZN(n4689) );
  NOR2_X1 U2460 ( .A1(n4694), .A2(n4078), .ZN(n4703) );
  INV_X1 U2461 ( .A(n2095), .ZN(n4704) );
  OR2_X1 U2462 ( .A1(n4703), .A2(n4702), .ZN(n2095) );
  OAI21_X1 U2463 ( .B1(n4708), .B2(n2161), .A(n2160), .ZN(n2159) );
  AOI21_X1 U2464 ( .B1(n4711), .B2(ADDR_REG_18__SCAN_IN), .A(n4710), .ZN(n2160) );
  INV_X1 U2465 ( .A(n2162), .ZN(n2161) );
  AOI21_X1 U2466 ( .B1(n2163), .B2(n4709), .A(n4707), .ZN(n2162) );
  OR2_X1 U2467 ( .A1(n4704), .A2(n2214), .ZN(n4712) );
  AND2_X1 U2468 ( .A1(n3987), .A2(n3986), .ZN(n4713) );
  NAND2_X1 U2469 ( .A1(n2248), .A2(n2251), .ZN(n2651) );
  INV_X1 U2470 ( .A(n4611), .ZN(n4087) );
  OR2_X1 U2471 ( .A1(n3337), .A2(n4605), .ZN(n2641) );
  AND2_X2 U2472 ( .A1(n2644), .A2(n3095), .ZN(n4789) );
  NOR2_X1 U2473 ( .A1(n2285), .A2(IR_REG_29__SCAN_IN), .ZN(n2981) );
  AND2_X1 U2474 ( .A1(n2803), .A2(n2186), .ZN(n2185) );
  NAND2_X1 U2475 ( .A1(n2808), .A2(n3622), .ZN(n2186) );
  NAND2_X1 U2476 ( .A1(n2840), .A2(n2839), .ZN(n2179) );
  INV_X1 U2477 ( .A(IR_REG_10__SCAN_IN), .ZN(n2268) );
  AND2_X1 U2478 ( .A1(n2247), .A2(n2266), .ZN(n2245) );
  INV_X1 U2479 ( .A(IR_REG_6__SCAN_IN), .ZN(n2266) );
  AND2_X1 U2480 ( .A1(n2181), .A2(n2183), .ZN(n2180) );
  AND2_X1 U2481 ( .A1(n3474), .A2(n2184), .ZN(n2183) );
  NAND2_X1 U2482 ( .A1(n2185), .A2(n2796), .ZN(n2181) );
  OR2_X1 U2483 ( .A1(n2808), .A2(n3622), .ZN(n2184) );
  INV_X1 U2484 ( .A(n2185), .ZN(n2182) );
  INV_X1 U2485 ( .A(n2814), .ZN(n2815) );
  OR2_X1 U2486 ( .A1(n2525), .A2(n3385), .ZN(n2533) );
  AND2_X1 U2487 ( .A1(n2179), .A2(n3587), .ZN(n2170) );
  NAND2_X1 U2488 ( .A1(n2190), .A2(n2188), .ZN(n2740) );
  INV_X1 U2489 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2426) );
  OR2_X1 U2490 ( .A1(n2419), .A2(n3557), .ZN(n2427) );
  INV_X1 U2491 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2389) );
  AOI21_X1 U2492 ( .B1(n3058), .B2(REG2_REG_7__SCAN_IN), .A(n3053), .ZN(n4045)
         );
  INV_X1 U2493 ( .A(n2111), .ZN(n2110) );
  OAI21_X1 U2494 ( .B1(n2112), .B2(n2114), .A(n2117), .ZN(n2111) );
  NAND2_X1 U2495 ( .A1(n2052), .A2(n4098), .ZN(n2117) );
  NAND2_X1 U2496 ( .A1(n4270), .A2(n2081), .ZN(n4158) );
  NAND2_X1 U2497 ( .A1(n2466), .A2(n2280), .ZN(n2481) );
  NOR2_X1 U2498 ( .A1(n2591), .A2(n2243), .ZN(n2242) );
  INV_X1 U2499 ( .A(n3707), .ZN(n2243) );
  AOI21_X1 U2500 ( .B1(n3709), .B2(n2240), .A(n4334), .ZN(n2239) );
  INV_X1 U2501 ( .A(n2242), .ZN(n2240) );
  INV_X1 U2502 ( .A(n3694), .ZN(n2221) );
  AND3_X1 U2503 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2348) );
  AND2_X1 U2504 ( .A1(n2317), .A2(n3136), .ZN(n2129) );
  NAND2_X1 U2505 ( .A1(n2131), .A2(n2317), .ZN(n2130) );
  INV_X1 U2506 ( .A(n2311), .ZN(n2131) );
  NAND2_X1 U2507 ( .A1(n3068), .A2(n3078), .ZN(n3680) );
  AND2_X1 U2508 ( .A1(n2060), .A2(n4430), .ZN(n2146) );
  OR2_X1 U2509 ( .A1(n2449), .A2(n2448), .ZN(n4325) );
  OR2_X1 U2510 ( .A1(n2973), .A2(n2634), .ZN(n2899) );
  OR2_X1 U2511 ( .A1(n2973), .A2(D_REG_1__SCAN_IN), .ZN(n2900) );
  NOR2_X1 U2512 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2474)
         );
  NOR2_X1 U2513 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2270)
         );
  NAND3_X1 U2514 ( .A1(n3564), .A2(n3383), .A3(n3381), .ZN(n3382) );
  OR2_X1 U2515 ( .A1(n3396), .A2(n3394), .ZN(n3399) );
  AOI21_X1 U2516 ( .B1(n2077), .B2(n2197), .A(n2196), .ZN(n2195) );
  NOR2_X1 U2517 ( .A1(n2199), .A2(n2198), .ZN(n2197) );
  INV_X1 U2518 ( .A(n3610), .ZN(n2196) );
  INV_X1 U2519 ( .A(n3464), .ZN(n2199) );
  NAND2_X1 U2520 ( .A1(n2167), .A2(n2166), .ZN(n3443) );
  NAND2_X1 U2521 ( .A1(n2056), .A2(n2178), .ZN(n2166) );
  MUX2_X1 U2522 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2051), .Z(n2677) );
  NAND2_X1 U2523 ( .A1(n2174), .A2(n2172), .ZN(n3540) );
  NAND2_X1 U2524 ( .A1(n3590), .A2(n2170), .ZN(n2174) );
  OAI21_X2 U2525 ( .B1(n3454), .B2(n3450), .A(n3451), .ZN(n3555) );
  AOI21_X1 U2526 ( .B1(n2690), .B2(n2891), .A(n2689), .ZN(n2693) );
  AOI21_X1 U2527 ( .B1(n3507), .B2(n3509), .A(n3506), .ZN(n3466) );
  AND3_X1 U2528 ( .A1(n3094), .A2(n2901), .A3(n2900), .ZN(n2920) );
  AOI21_X1 U2529 ( .B1(n2187), .B2(n2803), .A(n2809), .ZN(n3620) );
  OR3_X1 U2530 ( .A1(n2710), .A2(n2936), .A3(n2913), .ZN(n2917) );
  OR2_X1 U2531 ( .A1(n2557), .A2(n2282), .ZN(n3361) );
  OR2_X1 U2532 ( .A1(n2552), .A2(n2551), .ZN(n3615) );
  INV_X1 U2533 ( .A(n4750), .ZN(n2936) );
  AND2_X1 U2534 ( .A1(n4010), .A2(n4009), .ZN(n4007) );
  XNOR2_X1 U2535 ( .A(n2216), .B(n3001), .ZN(n3042) );
  AOI22_X1 U2536 ( .A1(n3013), .A2(REG2_REG_6__SCAN_IN), .B1(n4613), .B2(n3006), .ZN(n3055) );
  OR2_X1 U2537 ( .A1(n2996), .A2(n3017), .ZN(n2207) );
  NAND2_X1 U2538 ( .A1(n4624), .A2(n4047), .ZN(n4048) );
  NAND2_X1 U2539 ( .A1(n4638), .A2(n4033), .ZN(n4643) );
  INV_X1 U2540 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3557) );
  AND2_X1 U2541 ( .A1(n4053), .A2(n4054), .ZN(n2155) );
  NOR2_X1 U2542 ( .A1(n2155), .A2(n4056), .ZN(n2154) );
  NAND2_X1 U2543 ( .A1(n4698), .A2(n2164), .ZN(n2163) );
  OR2_X1 U2544 ( .A1(n4080), .A2(REG2_REG_17__SCAN_IN), .ZN(n2164) );
  NAND2_X1 U2545 ( .A1(n4715), .A2(n2090), .ZN(n2214) );
  OAI21_X1 U2546 ( .B1(n2251), .B2(n2250), .A(n3651), .ZN(n2249) );
  NAND2_X1 U2547 ( .A1(n4108), .A2(n2055), .ZN(n2248) );
  AOI21_X1 U2548 ( .B1(n2055), .B2(n3648), .A(n2252), .ZN(n2251) );
  OAI21_X1 U2549 ( .B1(n4198), .B2(n2134), .A(n2132), .ZN(n4156) );
  AOI21_X1 U2550 ( .B1(n2135), .B2(n2133), .A(n2078), .ZN(n2132) );
  INV_X1 U2551 ( .A(n2135), .ZN(n2134) );
  AND2_X1 U2552 ( .A1(n2503), .A2(REG3_REG_20__SCAN_IN), .ZN(n2516) );
  AND2_X1 U2553 ( .A1(n3764), .A2(n4159), .ZN(n4199) );
  NOR2_X1 U2554 ( .A1(n2493), .A2(n2492), .ZN(n2503) );
  NAND2_X1 U2555 ( .A1(n4253), .A2(n2491), .ZN(n4231) );
  AND2_X1 U2556 ( .A1(n4270), .A2(n3755), .ZN(n4234) );
  INV_X1 U2557 ( .A(n4262), .ZN(n4259) );
  AND2_X1 U2558 ( .A1(n3291), .A2(n3707), .ZN(n3763) );
  NAND2_X1 U2559 ( .A1(n2588), .A2(n3700), .ZN(n3267) );
  OAI21_X1 U2560 ( .B1(n2586), .B2(n2222), .A(n2220), .ZN(n3256) );
  INV_X1 U2561 ( .A(n2223), .ZN(n2222) );
  AOI21_X1 U2562 ( .B1(n2226), .B2(n2223), .A(n2221), .ZN(n2220) );
  AND2_X1 U2563 ( .A1(n2225), .A2(n2224), .ZN(n2223) );
  NOR2_X1 U2564 ( .A1(n2383), .A2(n2121), .ZN(n2120) );
  NAND2_X1 U2565 ( .A1(n2586), .A2(n2227), .ZN(n4514) );
  NAND2_X1 U2566 ( .A1(n2122), .A2(n2123), .ZN(n3244) );
  NAND2_X1 U2567 ( .A1(n2586), .A2(n3691), .ZN(n3231) );
  INV_X1 U2568 ( .A(n3765), .ZN(n2327) );
  AND2_X1 U2569 ( .A1(n2899), .A2(n2974), .ZN(n3094) );
  NAND2_X1 U2570 ( .A1(n3138), .A2(n2311), .ZN(n3155) );
  INV_X1 U2571 ( .A(n2583), .ZN(n3762) );
  NAND2_X1 U2572 ( .A1(n2582), .A2(n3103), .ZN(n3137) );
  NAND2_X1 U2573 ( .A1(n3680), .A2(n3677), .ZN(n2582) );
  INV_X1 U2574 ( .A(n3078), .ZN(n3111) );
  AND2_X1 U2575 ( .A1(n3676), .A2(n3678), .ZN(n3778) );
  NOR2_X1 U2576 ( .A1(n4377), .A2(n4380), .ZN(n4376) );
  INV_X1 U2577 ( .A(n3669), .ZN(n4380) );
  NAND2_X1 U2578 ( .A1(n2143), .A2(n4128), .ZN(n2141) );
  NOR2_X1 U2579 ( .A1(n4383), .A2(n3338), .ZN(n2143) );
  OR2_X1 U2580 ( .A1(n2662), .A2(n3649), .ZN(n4377) );
  AND2_X1 U2581 ( .A1(n4114), .A2(n4098), .ZN(n4096) );
  NOR3_X1 U2582 ( .A1(n4146), .A2(n3614), .A3(n4395), .ZN(n4114) );
  NAND2_X1 U2583 ( .A1(n2051), .A2(DATAI_24_), .ZN(n4147) );
  AND2_X1 U2584 ( .A1(n4181), .A2(n4168), .ZN(n4170) );
  AND2_X1 U2585 ( .A1(n4200), .A2(n4191), .ZN(n4181) );
  AND2_X1 U2586 ( .A1(n4275), .A2(n2145), .ZN(n4200) );
  AND2_X1 U2587 ( .A1(n2146), .A2(n4202), .ZN(n2145) );
  NAND2_X1 U2588 ( .A1(n4275), .A2(n2146), .ZN(n4218) );
  NAND2_X1 U2589 ( .A1(n4275), .A2(n2060), .ZN(n4245) );
  NAND2_X1 U2590 ( .A1(n4275), .A2(n4259), .ZN(n4257) );
  AND2_X1 U2591 ( .A1(n4291), .A2(n4277), .ZN(n4275) );
  NOR2_X1 U2592 ( .A1(n4313), .A2(n4289), .ZN(n4291) );
  OR2_X1 U2593 ( .A1(n4337), .A2(n4458), .ZN(n4313) );
  INV_X1 U2594 ( .A(n4316), .ZN(n4462) );
  INV_X1 U2595 ( .A(n4466), .ZN(n4338) );
  NAND2_X1 U2596 ( .A1(n3258), .A2(n2062), .ZN(n3298) );
  NAND2_X1 U2597 ( .A1(n3258), .A2(n3305), .ZN(n3270) );
  INV_X1 U2598 ( .A(n3404), .ZN(n3305) );
  NOR2_X1 U2599 ( .A1(n4508), .A2(n3533), .ZN(n3258) );
  OR2_X1 U2600 ( .A1(n3228), .A2(n4517), .ZN(n4508) );
  INV_X1 U2601 ( .A(n4518), .ZN(n4500) );
  AND2_X1 U2602 ( .A1(n2089), .A2(n3212), .ZN(n3186) );
  NAND2_X1 U2603 ( .A1(n3212), .A2(n3211), .ZN(n3210) );
  AND2_X1 U2604 ( .A1(n4610), .A2(n3082), .ZN(n4518) );
  INV_X1 U2605 ( .A(n4519), .ZN(n4484) );
  AND2_X1 U2606 ( .A1(n3163), .A2(n2699), .ZN(n3212) );
  NOR2_X1 U2607 ( .A1(n3150), .A2(n3151), .ZN(n3163) );
  AND2_X1 U2608 ( .A1(n2283), .A2(IR_REG_31__SCAN_IN), .ZN(n2657) );
  AND2_X1 U2609 ( .A1(n2149), .A2(n2148), .ZN(n2147) );
  NOR2_X1 U2610 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .ZN(n2148)
         );
  NAND2_X1 U2611 ( .A1(n2201), .A2(IR_REG_31__SCAN_IN), .ZN(n2501) );
  NOR2_X1 U2612 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2202)
         );
  INV_X1 U2613 ( .A(IR_REG_19__SCAN_IN), .ZN(n2500) );
  NAND2_X1 U2614 ( .A1(n2434), .A2(n2433), .ZN(n2476) );
  INV_X1 U2615 ( .A(IR_REG_13__SCAN_IN), .ZN(n2433) );
  AND2_X1 U2616 ( .A1(n2396), .A2(n2260), .ZN(n2434) );
  NAND2_X1 U2617 ( .A1(n2053), .A2(n2247), .ZN(n2244) );
  NAND2_X1 U2618 ( .A1(n2246), .A2(n2053), .ZN(n2339) );
  INV_X1 U2619 ( .A(IR_REG_3__SCAN_IN), .ZN(n2323) );
  NAND2_X1 U2620 ( .A1(n2316), .A2(IR_REG_31__SCAN_IN), .ZN(n2324) );
  NAND2_X1 U2621 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2208)
         );
  AND2_X1 U2622 ( .A1(n2190), .A2(n2189), .ZN(n3349) );
  NAND2_X1 U2623 ( .A1(n2175), .A2(n3587), .ZN(n3420) );
  OR2_X1 U2624 ( .A1(n3590), .A2(n3586), .ZN(n2175) );
  INV_X1 U2625 ( .A(n4509), .ZN(n4517) );
  MUX2_X1 U2626 ( .A(n2997), .B(DATAI_1_), .S(n2310), .Z(n3078) );
  INV_X1 U2627 ( .A(n2723), .ZN(n3486) );
  INV_X1 U2628 ( .A(n2677), .ZN(n3112) );
  NAND4_X1 U2629 ( .A1(n2530), .A2(n2529), .A3(n2528), .A4(n2527), .ZN(n4188)
         );
  NAND4_X1 U2630 ( .A1(n2508), .A2(n2507), .A3(n2506), .A4(n2505), .ZN(n4242)
         );
  NAND4_X1 U2631 ( .A1(n2414), .A2(n2413), .A3(n2412), .A4(n2411), .ZN(n4496)
         );
  NAND2_X1 U2632 ( .A1(n2303), .A2(REG0_REG_12__SCAN_IN), .ZN(n2413) );
  NAND4_X1 U2633 ( .A1(n2408), .A2(n2407), .A3(n2406), .A4(n2405), .ZN(n3803)
         );
  NAND2_X1 U2634 ( .A1(n2303), .A2(REG0_REG_11__SCAN_IN), .ZN(n2407) );
  NAND4_X1 U2635 ( .A1(n2395), .A2(n2394), .A3(n2393), .A4(n2392), .ZN(n4494)
         );
  NAND4_X1 U2636 ( .A1(n2380), .A2(n2379), .A3(n2378), .A4(n2377), .ZN(n3434)
         );
  NAND4_X1 U2637 ( .A1(n2315), .A2(n2314), .A3(n2313), .A4(n2312), .ZN(n3981)
         );
  NAND4_X1 U2638 ( .A1(n2309), .A2(n2308), .A3(n2307), .A4(n2306), .ZN(n3983)
         );
  AOI22_X1 U2639 ( .A1(n4015), .A2(REG2_REG_4__SCAN_IN), .B1(n4614), .B2(n3003), .ZN(n3033) );
  NOR2_X1 U2640 ( .A1(n3033), .A2(n3032), .ZN(n3031) );
  NOR2_X1 U2641 ( .A1(n4016), .A2(n2066), .ZN(n3030) );
  INV_X1 U2642 ( .A(n2092), .ZN(n3028) );
  OR2_X1 U2643 ( .A1(n3014), .A2(n2995), .ZN(n3015) );
  NAND2_X1 U2644 ( .A1(n3015), .A2(n2207), .ZN(n3050) );
  XNOR2_X1 U2645 ( .A(n4027), .B(n4044), .ZN(n4029) );
  XNOR2_X1 U2646 ( .A(n4032), .B(n2150), .ZN(n4639) );
  NAND2_X1 U2647 ( .A1(n4639), .A2(REG1_REG_10__SCAN_IN), .ZN(n4638) );
  NAND2_X1 U2648 ( .A1(n4660), .A2(n4036), .ZN(n4673) );
  NAND2_X1 U2649 ( .A1(n4655), .A2(n4052), .ZN(n4668) );
  AND2_X1 U2650 ( .A1(n2154), .A2(n2153), .ZN(n4062) );
  NAND2_X1 U2651 ( .A1(n2153), .A2(n2152), .ZN(n4055) );
  INV_X1 U2652 ( .A(n2155), .ZN(n2152) );
  NAND2_X1 U2653 ( .A1(n4073), .A2(n4074), .ZN(n4684) );
  NAND2_X1 U2654 ( .A1(n4684), .A2(n4685), .ZN(n4683) );
  NOR2_X1 U2655 ( .A1(n2154), .A2(n4063), .ZN(n4680) );
  NAND2_X1 U2656 ( .A1(n4689), .A2(n4066), .ZN(n4697) );
  NOR2_X1 U2657 ( .A1(n2211), .A2(n2215), .ZN(n2210) );
  INV_X1 U2658 ( .A(n4666), .ZN(n4707) );
  AOI22_X1 U2659 ( .A1(n2649), .A2(n3743), .B1(n3338), .B2(n3802), .ZN(n2650)
         );
  NAND2_X1 U2660 ( .A1(n2254), .A2(n3657), .ZN(n4092) );
  AND3_X1 U2661 ( .A1(n2563), .A2(n2562), .A3(n2561), .ZN(n4386) );
  NAND2_X1 U2662 ( .A1(n2109), .A2(n2113), .ZN(n4094) );
  AND2_X1 U2663 ( .A1(n2115), .A2(n2119), .ZN(n4106) );
  NAND2_X1 U2664 ( .A1(n4126), .A2(n2549), .ZN(n2115) );
  NAND2_X1 U2665 ( .A1(n2217), .A2(n3747), .ZN(n4123) );
  NAND2_X1 U2666 ( .A1(n2137), .A2(n2135), .ZN(n4179) );
  NAND2_X1 U2667 ( .A1(n2137), .A2(n2515), .ZN(n4177) );
  NAND2_X1 U2668 ( .A1(n2096), .A2(n2100), .ZN(n4254) );
  NAND2_X1 U2669 ( .A1(n4286), .A2(n2101), .ZN(n2096) );
  NAND2_X1 U2670 ( .A1(n4288), .A2(n2465), .ZN(n4273) );
  AND2_X1 U2671 ( .A1(n4722), .A2(n4518), .ZN(n4340) );
  OAI21_X1 U2672 ( .B1(n2219), .B2(n2226), .A(n2225), .ZN(n3241) );
  INV_X1 U2673 ( .A(n2586), .ZN(n2219) );
  NAND2_X1 U2674 ( .A1(n2347), .A2(n2346), .ZN(n3169) );
  NAND2_X1 U2675 ( .A1(n2230), .A2(n3689), .ZN(n3180) );
  NAND2_X1 U2676 ( .A1(n2235), .A2(n2234), .ZN(n2230) );
  AND2_X1 U2677 ( .A1(n4722), .A2(n3171), .ZN(n4312) );
  NAND2_X1 U2678 ( .A1(n2235), .A2(n3686), .ZN(n3204) );
  NAND2_X1 U2679 ( .A1(n4722), .A2(n3128), .ZN(n4371) );
  OR2_X1 U2680 ( .A1(n2922), .A2(n3113), .ZN(n4719) );
  INV_X1 U2681 ( .A(n4719), .ZN(n4736) );
  INV_X2 U2682 ( .A(n4722), .ZN(n4744) );
  OR2_X1 U2683 ( .A1(n3337), .A2(n4533), .ZN(n2647) );
  OAI21_X1 U2684 ( .B1(n2140), .B2(n3656), .A(n4377), .ZN(n3331) );
  OR2_X1 U2685 ( .A1(n2981), .A2(n2982), .ZN(n2284) );
  XNOR2_X1 U2686 ( .A(n2286), .B(IR_REG_29__SCAN_IN), .ZN(n2971) );
  XNOR2_X1 U2687 ( .A(n2576), .B(n2575), .ZN(n4617) );
  AND3_X1 U2688 ( .A1(n2257), .A2(n2396), .A3(n2138), .ZN(n2574) );
  XNOR2_X1 U2689 ( .A(n2617), .B(IR_REG_26__SCAN_IN), .ZN(n4607) );
  NAND2_X1 U2690 ( .A1(n2614), .A2(IR_REG_31__SCAN_IN), .ZN(n2615) );
  AND2_X1 U2691 ( .A1(n2941), .A2(STATE_REG_SCAN_IN), .ZN(n4750) );
  XNOR2_X1 U2692 ( .A(n2572), .B(IR_REG_22__SCAN_IN), .ZN(n4609) );
  NAND2_X1 U2693 ( .A1(n2396), .A2(n2259), .ZN(n2567) );
  AND2_X1 U2694 ( .A1(n2564), .A2(n2502), .ZN(n4611) );
  OR2_X1 U2695 ( .A1(n2501), .A2(n2500), .ZN(n2502) );
  NOR2_X1 U2696 ( .A1(n2297), .A2(n2982), .ZN(n2158) );
  NAND2_X1 U2697 ( .A1(n2935), .A2(n2263), .ZN(n2932) );
  INV_X1 U2698 ( .A(n2159), .ZN(n4717) );
  AND2_X1 U2699 ( .A1(n2095), .A2(n2090), .ZN(n4714) );
  AOI21_X1 U2700 ( .B1(n2645), .B2(n4789), .A(n2642), .ZN(n2643) );
  NAND2_X1 U2701 ( .A1(n2641), .A2(n2261), .ZN(n2642) );
  NAND2_X1 U2702 ( .A1(n3555), .A2(n2797), .ZN(n2187) );
  OAI21_X1 U2703 ( .B1(n2105), .B2(n2104), .A(n2479), .ZN(n2103) );
  NOR2_X1 U2704 ( .A1(n3428), .A2(n2769), .ZN(n2054) );
  INV_X1 U2705 ( .A(n3805), .ZN(n2125) );
  NOR2_X1 U2706 ( .A1(n4095), .A2(n2253), .ZN(n2055) );
  NAND2_X1 U2707 ( .A1(n2187), .A2(n2088), .ZN(n3472) );
  INV_X1 U2708 ( .A(n2165), .ZN(n2316) );
  NAND3_X1 U2709 ( .A1(n2302), .A2(n2300), .A3(n2301), .ZN(n2673) );
  INV_X1 U2710 ( .A(IR_REG_17__SCAN_IN), .ZN(n2488) );
  NAND2_X1 U2711 ( .A1(n2172), .A2(n2171), .ZN(n2056) );
  NOR2_X1 U2712 ( .A1(n2769), .A2(n3398), .ZN(n2057) );
  OR2_X1 U2713 ( .A1(n4007), .A2(n2070), .ZN(n2216) );
  INV_X1 U2714 ( .A(n3709), .ZN(n2241) );
  INV_X1 U2715 ( .A(n2796), .ZN(n2797) );
  AND2_X1 U2716 ( .A1(n2206), .A2(n4793), .ZN(n2058) );
  AND3_X1 U2717 ( .A1(n2246), .A2(n2053), .A3(n2245), .ZN(n2059) );
  AND2_X1 U2718 ( .A1(n4259), .A2(n4246), .ZN(n2060) );
  NAND2_X1 U2719 ( .A1(n4296), .A2(n4446), .ZN(n2061) );
  AND2_X1 U2720 ( .A1(n3305), .A2(n4499), .ZN(n2062) );
  INV_X1 U2721 ( .A(n3698), .ZN(n2232) );
  INV_X1 U2722 ( .A(n4260), .ZN(n2098) );
  AND2_X1 U2723 ( .A1(n3638), .A2(n3755), .ZN(n2063) );
  INV_X1 U2724 ( .A(n4098), .ZN(n4383) );
  INV_X1 U2725 ( .A(n2674), .ZN(n2895) );
  INV_X1 U2726 ( .A(n2690), .ZN(n3074) );
  NAND4_X1 U2727 ( .A1(n2296), .A2(n2295), .A3(n2294), .A4(n2293), .ZN(n2690)
         );
  NOR2_X1 U2728 ( .A1(n2244), .A2(n2316), .ZN(n2341) );
  OR2_X1 U2729 ( .A1(n2610), .A2(IR_REG_25__SCAN_IN), .ZN(n2064) );
  INV_X1 U2730 ( .A(n2714), .ZN(n3489) );
  NOR3_X1 U2731 ( .A1(n4146), .A2(n2141), .A3(n3614), .ZN(n2140) );
  AND2_X1 U2732 ( .A1(n4396), .A2(n3614), .ZN(n2065) );
  INV_X1 U2733 ( .A(n2717), .ZN(n2200) );
  AND2_X1 U2734 ( .A1(n2994), .A2(n4614), .ZN(n2066) );
  XNOR2_X1 U2735 ( .A(n2284), .B(IR_REG_30__SCAN_IN), .ZN(n2288) );
  INV_X1 U2736 ( .A(IR_REG_2__SCAN_IN), .ZN(n2157) );
  NOR2_X1 U2737 ( .A1(n3518), .A2(n2723), .ZN(n2067) );
  AND2_X1 U2738 ( .A1(n2216), .A2(n3001), .ZN(n2068) );
  AND2_X1 U2739 ( .A1(n2571), .A2(n2570), .ZN(n3786) );
  NOR2_X1 U2740 ( .A1(n2388), .A2(n2387), .ZN(n2069) );
  AND2_X1 U2741 ( .A1(n4615), .A2(REG1_REG_2__SCAN_IN), .ZN(n2070) );
  OR2_X1 U2742 ( .A1(n2116), .A2(n2065), .ZN(n2071) );
  AND3_X1 U2743 ( .A1(n2276), .A2(n2256), .A3(n2255), .ZN(n2072) );
  AND2_X1 U2744 ( .A1(n2055), .A2(n3660), .ZN(n2073) );
  AND2_X1 U2745 ( .A1(n2130), .A2(n2318), .ZN(n2074) );
  OR2_X1 U2746 ( .A1(n2475), .A2(IR_REG_16__SCAN_IN), .ZN(n2075) );
  INV_X1 U2747 ( .A(n2330), .ZN(n2579) );
  AND2_X1 U2748 ( .A1(n2288), .A2(n2289), .ZN(n2330) );
  AND2_X1 U2749 ( .A1(n2396), .A2(n2268), .ZN(n2399) );
  INV_X1 U2750 ( .A(n3604), .ZN(n2124) );
  AOI21_X1 U2751 ( .B1(n4295), .B2(n4294), .A(n3639), .ZN(n4270) );
  INV_X1 U2752 ( .A(IR_REG_27__SCAN_IN), .ZN(n2255) );
  AND2_X1 U2753 ( .A1(n4110), .A2(n4383), .ZN(n2076) );
  INV_X1 U2754 ( .A(n3463), .ZN(n2198) );
  OR2_X1 U2755 ( .A1(n2886), .A2(n2885), .ZN(n2077) );
  AND2_X1 U2756 ( .A1(n4423), .A2(n2524), .ZN(n2078) );
  AND2_X1 U2757 ( .A1(n4270), .A2(n2063), .ZN(n2079) );
  INV_X1 U2758 ( .A(n3658), .ZN(n2252) );
  AND2_X1 U2759 ( .A1(n2297), .A2(n2157), .ZN(n2165) );
  INV_X1 U2760 ( .A(n2316), .ZN(n2246) );
  NAND2_X1 U2761 ( .A1(n4242), .A2(n4430), .ZN(n2080) );
  NOR2_X1 U2762 ( .A1(n4146), .A2(n4395), .ZN(n2142) );
  INV_X1 U2763 ( .A(n2102), .ZN(n2101) );
  NAND2_X1 U2764 ( .A1(n2465), .A2(n2061), .ZN(n2102) );
  INV_X1 U2765 ( .A(n3675), .ZN(n2218) );
  AND2_X1 U2766 ( .A1(n2063), .A2(n2080), .ZN(n2081) );
  NAND2_X1 U2767 ( .A1(n3603), .A2(n2714), .ZN(n2082) );
  AND2_X1 U2768 ( .A1(n2365), .A2(n2372), .ZN(n3058) );
  INV_X1 U2769 ( .A(n3058), .ZN(n2206) );
  OR2_X1 U2770 ( .A1(n4310), .A2(n2592), .ZN(n2083) );
  INV_X1 U2771 ( .A(n2465), .ZN(n2104) );
  INV_X1 U2772 ( .A(n3696), .ZN(n2224) );
  NAND2_X1 U2773 ( .A1(n3434), .A2(n3533), .ZN(n2084) );
  AND2_X1 U2774 ( .A1(n2077), .A2(n3463), .ZN(n2085) );
  INV_X1 U2775 ( .A(n2119), .ZN(n2116) );
  NAND2_X1 U2776 ( .A1(n4405), .A2(n4395), .ZN(n2119) );
  AND2_X1 U2777 ( .A1(n2604), .A2(n3747), .ZN(n2086) );
  AND2_X1 U2778 ( .A1(n2062), .A2(n4479), .ZN(n2087) );
  INV_X1 U2779 ( .A(IR_REG_31__SCAN_IN), .ZN(n2982) );
  NAND2_X1 U2780 ( .A1(n3156), .A2(n3761), .ZN(n2235) );
  XNOR2_X1 U2781 ( .A(n2718), .B(n2200), .ZN(n2723) );
  INV_X1 U2782 ( .A(n4116), .ZN(n3614) );
  NAND2_X1 U2783 ( .A1(n2310), .A2(DATAI_26_), .ZN(n4116) );
  AOI21_X1 U2784 ( .B1(n2122), .B2(n2120), .A(n2069), .ZN(n3257) );
  AOI21_X1 U2785 ( .B1(n2235), .B2(n2233), .A(n2231), .ZN(n3168) );
  NAND2_X1 U2786 ( .A1(n3484), .A2(n2725), .ZN(n3597) );
  AND2_X1 U2787 ( .A1(n3715), .A2(n3717), .ZN(n4294) );
  INV_X1 U2788 ( .A(n4294), .ZN(n2105) );
  NAND2_X1 U2789 ( .A1(n2051), .A2(DATAI_21_), .ZN(n4202) );
  AND2_X1 U2790 ( .A1(n2803), .A2(n2809), .ZN(n2088) );
  NAND2_X1 U2791 ( .A1(n2051), .A2(DATAI_20_), .ZN(n4430) );
  AND2_X1 U2792 ( .A1(n3211), .A2(n2714), .ZN(n2089) );
  NAND2_X1 U2793 ( .A1(n2310), .A2(DATAI_25_), .ZN(n4128) );
  AND2_X2 U2794 ( .A1(n2644), .A2(n2901), .ZN(n4795) );
  NAND4_X1 U2795 ( .A1(n3212), .A2(n3211), .A3(n2714), .A4(n2124), .ZN(n3230)
         );
  INV_X1 U2796 ( .A(n3230), .ZN(n2144) );
  NAND2_X1 U2797 ( .A1(n2310), .A2(DATAI_28_), .ZN(n2896) );
  NOR2_X1 U2798 ( .A1(n4753), .A2(n4081), .ZN(n2215) );
  INV_X1 U2799 ( .A(n4654), .ZN(n2151) );
  INV_X1 U2800 ( .A(n4632), .ZN(n2150) );
  OR2_X1 U2801 ( .A1(n4080), .A2(REG1_REG_17__SCAN_IN), .ZN(n2090) );
  NAND2_X1 U2802 ( .A1(n4126), .A2(n2114), .ZN(n2109) );
  NAND2_X1 U2803 ( .A1(n2673), .A2(n2731), .ZN(n2670) );
  NAND2_X1 U2804 ( .A1(n2074), .A2(n2128), .ZN(n3201) );
  NAND3_X1 U2805 ( .A1(n2583), .A2(n3137), .A3(n2129), .ZN(n2128) );
  NAND3_X1 U2806 ( .A1(n2583), .A2(n3137), .A3(n3136), .ZN(n3138) );
  AND2_X1 U2807 ( .A1(n2257), .A2(n2396), .ZN(n2569) );
  NAND4_X1 U2808 ( .A1(n2257), .A2(n2396), .A3(n2138), .A4(n2575), .ZN(n2285)
         );
  NAND3_X1 U2809 ( .A1(n2257), .A2(n2396), .A3(n2149), .ZN(n2610) );
  NOR2_X2 U2810 ( .A1(n2381), .A2(IR_REG_9__SCAN_IN), .ZN(n2396) );
  NAND3_X1 U2811 ( .A1(n2165), .A2(n2139), .A3(n2053), .ZN(n2381) );
  INV_X1 U2812 ( .A(n2140), .ZN(n2662) );
  INV_X1 U2813 ( .A(n2142), .ZN(n4127) );
  NAND2_X1 U2814 ( .A1(n2144), .A2(n3233), .ZN(n3228) );
  NAND2_X1 U2815 ( .A1(n2569), .A2(n2147), .ZN(n2283) );
  INV_X1 U2816 ( .A(n4063), .ZN(n2153) );
  MUX2_X1 U2817 ( .A(REG2_REG_2__SCAN_IN), .B(n4001), .S(n4615), .Z(n2999) );
  XNOR2_X2 U2818 ( .A(n2158), .B(n2157), .ZN(n4615) );
  NOR2_X1 U2819 ( .A1(n4053), .A2(n4054), .ZN(n4063) );
  NOR2_X1 U2820 ( .A1(n4680), .A2(n4679), .ZN(n4678) );
  NAND2_X1 U2821 ( .A1(n4699), .A2(n4697), .ZN(n4698) );
  NOR2_X1 U2822 ( .A1(n3055), .A2(n3054), .ZN(n3053) );
  NAND2_X1 U2823 ( .A1(n3590), .A2(n2168), .ZN(n2167) );
  INV_X1 U2824 ( .A(n3543), .ZN(n2178) );
  NAND2_X1 U2825 ( .A1(n3466), .A2(n2085), .ZN(n2194) );
  NAND2_X1 U2826 ( .A1(n2194), .A2(n2195), .ZN(n3360) );
  OAI21_X1 U2827 ( .B1(n3466), .B2(n3464), .A(n3463), .ZN(n3612) );
  NAND2_X1 U2828 ( .A1(n2489), .A2(n2202), .ZN(n2201) );
  XNOR2_X2 U2829 ( .A(n2208), .B(IR_REG_1__SCAN_IN), .ZN(n2997) );
  NAND2_X1 U2830 ( .A1(n2209), .A2(n2210), .ZN(n4084) );
  NAND2_X1 U2831 ( .A1(n4703), .A2(n2213), .ZN(n2209) );
  NAND2_X1 U2832 ( .A1(n2217), .A2(n2086), .ZN(n2605) );
  NAND2_X1 U2833 ( .A1(n3267), .A2(n2239), .ZN(n2236) );
  NAND2_X1 U2834 ( .A1(n2236), .A2(n2237), .ZN(n2593) );
  AOI21_X1 U2835 ( .B1(n4108), .B2(n2073), .A(n2249), .ZN(n2652) );
  OR2_X1 U2836 ( .A1(n4108), .A2(n3648), .ZN(n2254) );
  NAND2_X1 U2837 ( .A1(n4158), .A2(n3641), .ZN(n2603) );
  AND2_X1 U2838 ( .A1(n2299), .A2(n2298), .ZN(n2302) );
  INV_X1 U2839 ( .A(n2288), .ZN(n2287) );
  INV_X1 U2840 ( .A(n3414), .ZN(n2699) );
  NAND2_X1 U2841 ( .A1(n4368), .A2(n4338), .ZN(n4337) );
  NAND2_X1 U2842 ( .A1(n4170), .A2(n4147), .ZN(n4146) );
  NAND2_X1 U2843 ( .A1(n3681), .A2(n3684), .ZN(n2583) );
  OR2_X1 U2844 ( .A1(n3331), .A2(n4533), .ZN(n2667) );
  OR2_X1 U2845 ( .A1(n3331), .A2(n4605), .ZN(n2663) );
  OAI21_X1 U2846 ( .B1(n3676), .B2(n2582), .A(n3680), .ZN(n3142) );
  XNOR2_X1 U2847 ( .A(n2650), .B(n3779), .ZN(n3329) );
  MUX2_X2 U2848 ( .A(n2279), .B(n2278), .S(n2255), .Z(n2310) );
  OR2_X1 U2849 ( .A1(n4789), .A2(n2640), .ZN(n2261) );
  AND2_X1 U2850 ( .A1(n2659), .A2(n2658), .ZN(n2262) );
  INV_X1 U2851 ( .A(n4423), .ZN(n4207) );
  NAND2_X1 U2852 ( .A1(n2051), .A2(DATAI_22_), .ZN(n4191) );
  AND3_X1 U2853 ( .A1(n2931), .A2(n2930), .A3(n3624), .ZN(n2263) );
  AND2_X1 U2854 ( .A1(n2647), .A2(n2646), .ZN(n2264) );
  AND2_X1 U2855 ( .A1(n2923), .A2(n4719), .ZN(n3122) );
  NAND2_X2 U2856 ( .A1(n3096), .A2(n4719), .ZN(n4722) );
  OAI21_X1 U2857 ( .B1(n3369), .B2(n3552), .A(n3372), .ZN(n2796) );
  INV_X1 U2858 ( .A(IR_REG_4__SCAN_IN), .ZN(n2265) );
  INV_X1 U2859 ( .A(n2808), .ZN(n2809) );
  INV_X1 U2860 ( .A(n2657), .ZN(n2277) );
  INV_X1 U2861 ( .A(n2891), .ZN(n2892) );
  OR2_X1 U2862 ( .A1(n2535), .A2(n3129), .ZN(n2301) );
  AND2_X1 U2863 ( .A1(n3746), .A2(n4139), .ZN(n3675) );
  INV_X1 U2864 ( .A(n4191), .ZN(n2524) );
  INV_X1 U2865 ( .A(REG0_REG_28__SCAN_IN), .ZN(n2640) );
  INV_X1 U2866 ( .A(IR_REG_26__SCAN_IN), .ZN(n2276) );
  NAND2_X1 U2867 ( .A1(n2816), .A2(n2815), .ZN(n2817) );
  AOI21_X1 U2868 ( .B1(n2770), .B2(n2054), .A(n2057), .ZN(n3573) );
  NOR2_X1 U2869 ( .A1(n2427), .A2(n2426), .ZN(n2436) );
  OR2_X1 U2870 ( .A1(n2481), .A2(n2480), .ZN(n2493) );
  AND2_X1 U2871 ( .A1(n2436), .A2(REG3_REG_15__SCAN_IN), .ZN(n2466) );
  INV_X1 U2872 ( .A(n3656), .ZN(n3649) );
  INV_X1 U2873 ( .A(n4522), .ZN(n4495) );
  AND2_X1 U2874 ( .A1(n4609), .A2(n3786), .ZN(n2939) );
  INV_X1 U2875 ( .A(REG3_REG_7__SCAN_IN), .ZN(n3051) );
  NOR2_X1 U2876 ( .A1(n2542), .A2(n2541), .ZN(n2550) );
  AND2_X1 U2877 ( .A1(n2846), .A2(n2845), .ZN(n3543) );
  AND2_X1 U2878 ( .A1(n2552), .A2(REG3_REG_27__SCAN_IN), .ZN(n2557) );
  AND2_X1 U2879 ( .A1(n2550), .A2(REG3_REG_26__SCAN_IN), .ZN(n2552) );
  INV_X1 U2880 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3961) );
  INV_X1 U2881 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3578) );
  AND2_X1 U2882 ( .A1(n3775), .A2(n3774), .ZN(n4515) );
  AND2_X1 U2883 ( .A1(n3686), .A2(n3683), .ZN(n3761) );
  OR2_X1 U2884 ( .A1(n2973), .A2(D_REG_0__SCAN_IN), .ZN(n2638) );
  NAND2_X1 U2885 ( .A1(n2310), .A2(DATAI_23_), .ZN(n4168) );
  INV_X1 U2886 ( .A(n3558), .ZN(n4365) );
  AND2_X1 U2887 ( .A1(n2580), .A2(n2921), .ZN(n3082) );
  OR2_X1 U2888 ( .A1(n3090), .A2(n2942), .ZN(n2951) );
  INV_X1 U2889 ( .A(n4168), .ZN(n3780) );
  INV_X1 U2890 ( .A(n4202), .ZN(n4422) );
  INV_X1 U2891 ( .A(n4128), .ZN(n4395) );
  INV_X1 U2892 ( .A(n4430), .ZN(n3546) );
  AND2_X1 U2893 ( .A1(n2905), .A2(n3090), .ZN(n2906) );
  NAND2_X2 U2894 ( .A1(n2915), .A2(n3066), .ZN(n3630) );
  AND2_X1 U2895 ( .A1(n2943), .A2(n2951), .ZN(n3987) );
  AND2_X1 U2896 ( .A1(n3987), .A2(n3794), .ZN(n4666) );
  INV_X1 U2897 ( .A(n4371), .ZN(n4738) );
  AND2_X1 U2898 ( .A1(n2638), .A2(n2637), .ZN(n2901) );
  NAND2_X1 U2899 ( .A1(n2310), .A2(DATAI_27_), .ZN(n4098) );
  NAND2_X1 U2900 ( .A1(n4524), .A2(n3113), .ZN(n4492) );
  INV_X1 U2901 ( .A(n2901), .ZN(n3095) );
  XNOR2_X1 U2902 ( .A(n2621), .B(n2620), .ZN(n2941) );
  AND2_X1 U2903 ( .A1(n2401), .A2(n2400), .ZN(n4632) );
  AND2_X1 U2904 ( .A1(n2952), .A2(n2951), .ZN(n4711) );
  NAND2_X1 U2905 ( .A1(n2920), .A2(n2906), .ZN(n3517) );
  INV_X1 U2906 ( .A(n4386), .ZN(n3802) );
  NAND4_X1 U2907 ( .A1(n2548), .A2(n2547), .A3(n2546), .A4(n2545), .ZN(n4405)
         );
  OR2_X2 U2908 ( .A1(n2937), .A2(n2936), .ZN(n3982) );
  INV_X1 U2909 ( .A(n4713), .ZN(n3060) );
  NAND2_X1 U2910 ( .A1(n3987), .A2(n4617), .ZN(n4718) );
  INV_X1 U2911 ( .A(n4312), .ZN(n4375) );
  NAND2_X1 U2912 ( .A1(n4795), .A2(n4258), .ZN(n4533) );
  INV_X1 U2913 ( .A(n4795), .ZN(n4792) );
  NAND2_X1 U2914 ( .A1(n4789), .A2(n4258), .ZN(n4605) );
  INV_X1 U2915 ( .A(n4789), .ZN(n4787) );
  NAND2_X1 U2916 ( .A1(n2973), .A2(n3090), .ZN(n4749) );
  XNOR2_X1 U2917 ( .A(n2615), .B(IR_REG_24__SCAN_IN), .ZN(n4608) );
  INV_X1 U2918 ( .A(n4080), .ZN(n4754) );
  INV_X1 U2919 ( .A(n3017), .ZN(n4613) );
  INV_X1 U2920 ( .A(n3982), .ZN(U4043) );
  INV_X1 U2921 ( .A(n2643), .ZN(U3514) );
  NAND2_X1 U2922 ( .A1(n2657), .A2(IR_REG_28__SCAN_IN), .ZN(n2279) );
  NAND2_X1 U2923 ( .A1(n2277), .A2(n2575), .ZN(n2278) );
  NAND2_X1 U2924 ( .A1(n2348), .A2(REG3_REG_6__SCAN_IN), .ZN(n2356) );
  NOR2_X1 U2925 ( .A1(n2356), .A2(n3051), .ZN(n2366) );
  NAND2_X1 U2926 ( .A1(n2366), .A2(REG3_REG_8__SCAN_IN), .ZN(n2375) );
  NAND2_X1 U2927 ( .A1(n2409), .A2(REG3_REG_12__SCAN_IN), .ZN(n2419) );
  AND2_X1 U2928 ( .A1(REG3_REG_16__SCAN_IN), .A2(REG3_REG_17__SCAN_IN), .ZN(
        n2280) );
  INV_X1 U2929 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2480) );
  INV_X1 U2930 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2492) );
  AND2_X1 U2931 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2281) );
  NAND2_X1 U2932 ( .A1(n2516), .A2(n2281), .ZN(n2525) );
  INV_X1 U2933 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3385) );
  INV_X1 U2934 ( .A(REG3_REG_24__SCAN_IN), .ZN(n2532) );
  INV_X1 U2935 ( .A(REG3_REG_25__SCAN_IN), .ZN(n2541) );
  NOR2_X1 U2936 ( .A1(n2552), .A2(REG3_REG_27__SCAN_IN), .ZN(n2282) );
  NAND2_X1 U2937 ( .A1(n2285), .A2(IR_REG_31__SCAN_IN), .ZN(n2286) );
  AND2_X2 U2938 ( .A1(n2287), .A2(n2971), .ZN(n2304) );
  AOI22_X1 U2939 ( .A1(n2304), .A2(REG1_REG_27__SCAN_IN), .B1(n2303), .B2(
        REG0_REG_27__SCAN_IN), .ZN(n2291) );
  NAND2_X1 U2940 ( .A1(n2330), .A2(REG2_REG_27__SCAN_IN), .ZN(n2290) );
  OAI211_X2 U2941 ( .C1(n3361), .C2(n2535), .A(n2291), .B(n2290), .ZN(n4110)
         );
  NAND2_X1 U2942 ( .A1(n2303), .A2(REG0_REG_2__SCAN_IN), .ZN(n2296) );
  NAND2_X1 U2943 ( .A1(n2330), .A2(REG2_REG_2__SCAN_IN), .ZN(n2295) );
  NAND2_X1 U2944 ( .A1(n2304), .A2(REG1_REG_2__SCAN_IN), .ZN(n2294) );
  INV_X1 U2945 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2292) );
  OR2_X1 U2946 ( .A1(n2535), .A2(n2292), .ZN(n2293) );
  NAND2_X1 U2947 ( .A1(n3074), .A2(n3151), .ZN(n3681) );
  INV_X1 U2948 ( .A(n3151), .ZN(n3121) );
  NAND2_X1 U2949 ( .A1(n2690), .A2(n3121), .ZN(n3684) );
  NAND2_X1 U2950 ( .A1(n2303), .A2(REG0_REG_1__SCAN_IN), .ZN(n2299) );
  NAND2_X1 U2951 ( .A1(n2304), .A2(REG1_REG_1__SCAN_IN), .ZN(n2298) );
  INV_X1 U2952 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3129) );
  NAND2_X1 U2953 ( .A1(n2330), .A2(REG2_REG_1__SCAN_IN), .ZN(n2300) );
  INV_X1 U2954 ( .A(n2673), .ZN(n3068) );
  NAND2_X1 U2955 ( .A1(n2673), .A2(n3111), .ZN(n3677) );
  NAND2_X1 U2956 ( .A1(n2303), .A2(REG0_REG_0__SCAN_IN), .ZN(n2309) );
  NAND2_X1 U2957 ( .A1(n2330), .A2(REG2_REG_0__SCAN_IN), .ZN(n2308) );
  NAND2_X1 U2958 ( .A1(n2304), .A2(REG1_REG_0__SCAN_IN), .ZN(n2307) );
  INV_X1 U2959 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2305) );
  OR2_X1 U2960 ( .A1(n2535), .A2(n2305), .ZN(n2306) );
  AND2_X1 U2961 ( .A1(n3983), .A2(n2677), .ZN(n3103) );
  NAND2_X1 U2962 ( .A1(n2673), .A2(n3078), .ZN(n3136) );
  NAND2_X1 U2963 ( .A1(n3074), .A2(n3121), .ZN(n2311) );
  NAND2_X1 U2964 ( .A1(n2303), .A2(REG0_REG_3__SCAN_IN), .ZN(n2315) );
  NAND2_X1 U2965 ( .A1(n2456), .A2(REG2_REG_3__SCAN_IN), .ZN(n2314) );
  NAND2_X1 U2966 ( .A1(n2304), .A2(REG1_REG_3__SCAN_IN), .ZN(n2313) );
  OR2_X1 U2967 ( .A1(n2535), .A2(REG3_REG_3__SCAN_IN), .ZN(n2312) );
  MUX2_X1 U2968 ( .A(n3001), .B(DATAI_3_), .S(n2310), .Z(n3414) );
  NAND2_X1 U2969 ( .A1(n3981), .A2(n3414), .ZN(n2317) );
  INV_X1 U2970 ( .A(n3981), .ZN(n3144) );
  NAND2_X1 U2971 ( .A1(n3144), .A2(n2699), .ZN(n2318) );
  INV_X1 U2972 ( .A(n3201), .ZN(n2328) );
  NAND2_X1 U2973 ( .A1(n2304), .A2(REG1_REG_4__SCAN_IN), .ZN(n2322) );
  NAND2_X1 U2974 ( .A1(n2303), .A2(REG0_REG_4__SCAN_IN), .ZN(n2321) );
  NAND2_X1 U2975 ( .A1(n2456), .A2(REG2_REG_4__SCAN_IN), .ZN(n2320) );
  XNOR2_X1 U2976 ( .A(REG3_REG_4__SCAN_IN), .B(REG3_REG_3__SCAN_IN), .ZN(n3522) );
  OR2_X1 U2977 ( .A1(n2535), .A2(n3522), .ZN(n2319) );
  INV_X1 U2978 ( .A(n3806), .ZN(n3183) );
  NAND2_X1 U2979 ( .A1(n2324), .A2(n2323), .ZN(n2325) );
  NAND2_X1 U2980 ( .A1(n2325), .A2(IR_REG_31__SCAN_IN), .ZN(n2326) );
  XNOR2_X1 U2981 ( .A(n2326), .B(IR_REG_4__SCAN_IN), .ZN(n4614) );
  MUX2_X1 U2982 ( .A(n4614), .B(DATAI_4_), .S(n2051), .Z(n3521) );
  NAND2_X1 U2983 ( .A1(n3183), .A2(n3521), .ZN(n3687) );
  NAND2_X1 U2984 ( .A1(n3806), .A2(n3211), .ZN(n3689) );
  NAND2_X1 U2985 ( .A1(n2328), .A2(n2327), .ZN(n3203) );
  NAND2_X1 U2986 ( .A1(n3806), .A2(n3521), .ZN(n2329) );
  NAND2_X1 U2987 ( .A1(n3203), .A2(n2329), .ZN(n3179) );
  NAND2_X1 U2988 ( .A1(n2304), .A2(REG1_REG_5__SCAN_IN), .ZN(n2338) );
  NAND2_X1 U2989 ( .A1(n2303), .A2(REG0_REG_5__SCAN_IN), .ZN(n2337) );
  NAND2_X1 U2990 ( .A1(n2330), .A2(REG2_REG_5__SCAN_IN), .ZN(n2336) );
  INV_X1 U2991 ( .A(n2348), .ZN(n2334) );
  INV_X1 U2992 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2332) );
  NAND2_X1 U2993 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2331) );
  NAND2_X1 U2994 ( .A1(n2332), .A2(n2331), .ZN(n2333) );
  NAND2_X1 U2995 ( .A1(n2334), .A2(n2333), .ZN(n3490) );
  OR2_X1 U2996 ( .A1(n2535), .A2(n3490), .ZN(n2335) );
  INV_X1 U2997 ( .A(n3603), .ZN(n2585) );
  NAND2_X1 U2998 ( .A1(n2339), .A2(IR_REG_31__SCAN_IN), .ZN(n2340) );
  MUX2_X1 U2999 ( .A(IR_REG_31__SCAN_IN), .B(n2340), .S(IR_REG_5__SCAN_IN), 
        .Z(n2343) );
  INV_X1 U3000 ( .A(n2341), .ZN(n2342) );
  NAND2_X1 U3001 ( .A1(n2343), .A2(n2342), .ZN(n3035) );
  INV_X1 U3002 ( .A(DATAI_5_), .ZN(n2344) );
  MUX2_X1 U3003 ( .A(n3035), .B(n2344), .S(n2310), .Z(n2714) );
  NAND2_X1 U3004 ( .A1(n2585), .A2(n2714), .ZN(n2345) );
  NAND2_X1 U3005 ( .A1(n3179), .A2(n2345), .ZN(n2347) );
  NAND2_X1 U3006 ( .A1(n3603), .A2(n3489), .ZN(n2346) );
  NAND2_X1 U3007 ( .A1(n2304), .A2(REG1_REG_6__SCAN_IN), .ZN(n2352) );
  NAND2_X1 U3008 ( .A1(n2303), .A2(REG0_REG_6__SCAN_IN), .ZN(n2351) );
  NAND2_X1 U3009 ( .A1(n2456), .A2(REG2_REG_6__SCAN_IN), .ZN(n2350) );
  OAI21_X1 U3010 ( .B1(n2348), .B2(REG3_REG_6__SCAN_IN), .A(n2356), .ZN(n3173)
         );
  OR2_X1 U3011 ( .A1(n2535), .A2(n3173), .ZN(n2349) );
  NAND4_X1 U3012 ( .A1(n2352), .A2(n2351), .A3(n2350), .A4(n2349), .ZN(n3805)
         );
  NOR2_X1 U3013 ( .A1(n2341), .A2(n2982), .ZN(n2353) );
  MUX2_X1 U3014 ( .A(n2982), .B(n2353), .S(IR_REG_6__SCAN_IN), .Z(n2354) );
  OR2_X1 U3015 ( .A1(n2354), .A2(n2059), .ZN(n3017) );
  MUX2_X1 U3016 ( .A(n4613), .B(DATAI_6_), .S(n2310), .Z(n3604) );
  AND2_X1 U3017 ( .A1(n3805), .A2(n3604), .ZN(n2355) );
  NAND2_X1 U3018 ( .A1(n2304), .A2(REG1_REG_7__SCAN_IN), .ZN(n2361) );
  NAND2_X1 U3019 ( .A1(n2303), .A2(REG0_REG_7__SCAN_IN), .ZN(n2360) );
  NAND2_X1 U3020 ( .A1(n2456), .A2(REG2_REG_7__SCAN_IN), .ZN(n2359) );
  AND2_X1 U3021 ( .A1(n2356), .A2(n3051), .ZN(n2357) );
  OR2_X1 U3022 ( .A1(n2357), .A2(n2366), .ZN(n3353) );
  OR2_X1 U3023 ( .A1(n2535), .A2(n3353), .ZN(n2358) );
  NAND4_X1 U3024 ( .A1(n2361), .A2(n2360), .A3(n2359), .A4(n2358), .ZN(n4520)
         );
  INV_X1 U3025 ( .A(n4520), .ZN(n3216) );
  NOR2_X1 U3026 ( .A1(n2059), .A2(n2982), .ZN(n2362) );
  NAND2_X1 U3027 ( .A1(n2362), .A2(IR_REG_7__SCAN_IN), .ZN(n2365) );
  INV_X1 U3028 ( .A(n2362), .ZN(n2364) );
  INV_X1 U3029 ( .A(IR_REG_7__SCAN_IN), .ZN(n2363) );
  NAND2_X1 U3030 ( .A1(n2364), .A2(n2363), .ZN(n2372) );
  MUX2_X1 U3031 ( .A(n3058), .B(DATAI_7_), .S(n2051), .Z(n3352) );
  NAND2_X1 U3032 ( .A1(n3216), .A2(n3352), .ZN(n3692) );
  INV_X1 U3033 ( .A(n3352), .ZN(n3233) );
  NAND2_X1 U3034 ( .A1(n4520), .A2(n3233), .ZN(n4513) );
  NAND2_X1 U3035 ( .A1(n2304), .A2(REG1_REG_8__SCAN_IN), .ZN(n2371) );
  NAND2_X1 U3036 ( .A1(n2303), .A2(REG0_REG_8__SCAN_IN), .ZN(n2370) );
  NAND2_X1 U3037 ( .A1(n2456), .A2(REG2_REG_8__SCAN_IN), .ZN(n2369) );
  OR2_X1 U3038 ( .A1(n2366), .A2(REG3_REG_8__SCAN_IN), .ZN(n2367) );
  NAND2_X1 U3039 ( .A1(n2375), .A2(n2367), .ZN(n4720) );
  OR2_X1 U3040 ( .A1(n2535), .A2(n4720), .ZN(n2368) );
  NAND4_X1 U3041 ( .A1(n2371), .A2(n2370), .A3(n2369), .A4(n2368), .ZN(n3804)
         );
  INV_X1 U3042 ( .A(n3804), .ZN(n3282) );
  NAND2_X1 U3043 ( .A1(n2372), .A2(IR_REG_31__SCAN_IN), .ZN(n2374) );
  INV_X1 U3044 ( .A(IR_REG_8__SCAN_IN), .ZN(n2373) );
  XNOR2_X1 U3045 ( .A(n2374), .B(n2373), .ZN(n4044) );
  INV_X1 U3046 ( .A(DATAI_8_), .ZN(n2963) );
  MUX2_X1 U3047 ( .A(n4044), .B(n2963), .S(n2051), .Z(n4509) );
  AND2_X1 U3048 ( .A1(n3282), .A2(n4509), .ZN(n2386) );
  OR2_X1 U3049 ( .A1(n3777), .A2(n2386), .ZN(n3243) );
  NAND2_X1 U3050 ( .A1(n2304), .A2(REG1_REG_9__SCAN_IN), .ZN(n2380) );
  NAND2_X1 U3051 ( .A1(n2303), .A2(REG0_REG_9__SCAN_IN), .ZN(n2379) );
  NAND2_X1 U3052 ( .A1(n2456), .A2(REG2_REG_9__SCAN_IN), .ZN(n2378) );
  NAND2_X1 U3053 ( .A1(n2375), .A2(n3961), .ZN(n2376) );
  NAND2_X1 U3054 ( .A1(n2390), .A2(n2376), .ZN(n3534) );
  OR2_X1 U3055 ( .A1(n2535), .A2(n3534), .ZN(n2377) );
  INV_X1 U3056 ( .A(n3434), .ZN(n4523) );
  NAND2_X1 U3057 ( .A1(n2381), .A2(IR_REG_31__SCAN_IN), .ZN(n2382) );
  XNOR2_X1 U3058 ( .A(n2382), .B(IR_REG_9__SCAN_IN), .ZN(n4043) );
  MUX2_X1 U3059 ( .A(n4043), .B(DATAI_9_), .S(n2310), .Z(n3533) );
  INV_X1 U3060 ( .A(n3533), .ZN(n3278) );
  AND2_X1 U3061 ( .A1(n4523), .A2(n3278), .ZN(n2388) );
  OR2_X1 U3062 ( .A1(n3243), .A2(n2388), .ZN(n2383) );
  NAND2_X1 U3063 ( .A1(n4520), .A2(n3352), .ZN(n4511) );
  NAND2_X1 U3064 ( .A1(n3804), .A2(n4517), .ZN(n2384) );
  AND2_X1 U3065 ( .A1(n4511), .A2(n2384), .ZN(n2385) );
  OR2_X1 U3066 ( .A1(n2386), .A2(n2385), .ZN(n3245) );
  AND2_X1 U3067 ( .A1(n2084), .A2(n3245), .ZN(n2387) );
  NAND2_X1 U3068 ( .A1(n2304), .A2(REG1_REG_10__SCAN_IN), .ZN(n2395) );
  NAND2_X1 U3069 ( .A1(n2303), .A2(REG0_REG_10__SCAN_IN), .ZN(n2394) );
  NAND2_X1 U3070 ( .A1(n2456), .A2(REG2_REG_10__SCAN_IN), .ZN(n2393) );
  NAND2_X1 U3071 ( .A1(n2390), .A2(n2389), .ZN(n2391) );
  NAND2_X1 U3072 ( .A1(n2403), .A2(n2391), .ZN(n3259) );
  OR2_X1 U3073 ( .A1(n2535), .A2(n3259), .ZN(n2392) );
  INV_X1 U3074 ( .A(n2396), .ZN(n2397) );
  NAND2_X1 U3075 ( .A1(n2397), .A2(IR_REG_31__SCAN_IN), .ZN(n2398) );
  MUX2_X1 U3076 ( .A(IR_REG_31__SCAN_IN), .B(n2398), .S(IR_REG_10__SCAN_IN), 
        .Z(n2401) );
  INV_X1 U3077 ( .A(n2399), .ZN(n2400) );
  MUX2_X1 U3078 ( .A(n4632), .B(DATAI_10_), .S(n2310), .Z(n3404) );
  NOR2_X1 U3079 ( .A1(n4494), .A2(n3404), .ZN(n2402) );
  OAI22_X1 U3080 ( .A1(n3257), .A2(n2402), .B1(n2587), .B2(n3305), .ZN(n3268)
         );
  NAND2_X1 U3081 ( .A1(n2304), .A2(REG1_REG_11__SCAN_IN), .ZN(n2408) );
  NAND2_X1 U3082 ( .A1(n2456), .A2(REG2_REG_11__SCAN_IN), .ZN(n2406) );
  AND2_X1 U3083 ( .A1(n2403), .A2(n3578), .ZN(n2404) );
  OR2_X1 U3084 ( .A1(n2404), .A2(n2409), .ZN(n3580) );
  OR2_X1 U3085 ( .A1(n2535), .A2(n3580), .ZN(n2405) );
  INV_X1 U3086 ( .A(n3803), .ZN(n4485) );
  OR2_X1 U3087 ( .A1(n2399), .A2(n2982), .ZN(n2416) );
  XNOR2_X1 U3088 ( .A(n2416), .B(IR_REG_11__SCAN_IN), .ZN(n4762) );
  MUX2_X1 U3089 ( .A(n4762), .B(DATAI_11_), .S(n2051), .Z(n3579) );
  NAND2_X1 U3090 ( .A1(n4485), .A2(n3579), .ZN(n3291) );
  INV_X1 U3091 ( .A(n3579), .ZN(n4499) );
  NAND2_X1 U3092 ( .A1(n3803), .A2(n4499), .ZN(n3707) );
  NAND2_X1 U3093 ( .A1(n2304), .A2(REG1_REG_12__SCAN_IN), .ZN(n2414) );
  NAND2_X1 U3094 ( .A1(n2456), .A2(REG2_REG_12__SCAN_IN), .ZN(n2412) );
  OR2_X1 U3095 ( .A1(n2409), .A2(REG3_REG_12__SCAN_IN), .ZN(n2410) );
  NAND2_X1 U3096 ( .A1(n2419), .A2(n2410), .ZN(n3299) );
  OR2_X1 U3097 ( .A1(n2535), .A2(n3299), .ZN(n2411) );
  INV_X1 U3098 ( .A(IR_REG_11__SCAN_IN), .ZN(n2415) );
  NAND2_X1 U3099 ( .A1(n2416), .A2(n2415), .ZN(n2417) );
  NAND2_X1 U3100 ( .A1(n2417), .A2(IR_REG_31__SCAN_IN), .ZN(n2418) );
  XNOR2_X1 U3101 ( .A(n2418), .B(IR_REG_12__SCAN_IN), .ZN(n4654) );
  MUX2_X1 U3102 ( .A(n4654), .B(DATAI_12_), .S(n2310), .Z(n3457) );
  AND2_X1 U3103 ( .A1(n4496), .A2(n3457), .ZN(n2446) );
  OR2_X1 U3104 ( .A1(n3763), .A2(n2446), .ZN(n4352) );
  NAND2_X1 U3105 ( .A1(n2304), .A2(REG1_REG_13__SCAN_IN), .ZN(n2424) );
  NAND2_X1 U3106 ( .A1(n2303), .A2(REG0_REG_13__SCAN_IN), .ZN(n2423) );
  NAND2_X1 U3107 ( .A1(n2456), .A2(REG2_REG_13__SCAN_IN), .ZN(n2422) );
  NAND2_X1 U3108 ( .A1(n2419), .A2(n3557), .ZN(n2420) );
  NAND2_X1 U3109 ( .A1(n2427), .A2(n2420), .ZN(n3559) );
  OR2_X1 U3110 ( .A1(n2535), .A2(n3559), .ZN(n2421) );
  NAND4_X1 U3111 ( .A1(n2424), .A2(n2423), .A3(n2422), .A4(n2421), .ZN(n4481)
         );
  OR2_X1 U3112 ( .A1(n2434), .A2(n2982), .ZN(n2425) );
  XNOR2_X1 U3113 ( .A(n2425), .B(IR_REG_13__SCAN_IN), .ZN(n4759) );
  MUX2_X1 U3114 ( .A(n4759), .B(DATAI_13_), .S(n2051), .Z(n3558) );
  AND2_X1 U3115 ( .A1(n4481), .A2(n3558), .ZN(n2449) );
  OR2_X1 U3116 ( .A1(n4352), .A2(n2449), .ZN(n4324) );
  NAND2_X1 U3117 ( .A1(n2304), .A2(REG1_REG_14__SCAN_IN), .ZN(n2432) );
  NAND2_X1 U3118 ( .A1(n2303), .A2(REG0_REG_14__SCAN_IN), .ZN(n2431) );
  NAND2_X1 U3119 ( .A1(n2456), .A2(REG2_REG_14__SCAN_IN), .ZN(n2430) );
  AND2_X1 U3120 ( .A1(n2427), .A2(n2426), .ZN(n2428) );
  OR2_X1 U3121 ( .A1(n2428), .A2(n2436), .ZN(n3376) );
  OR2_X1 U3122 ( .A1(n2535), .A2(n3376), .ZN(n2429) );
  NAND4_X1 U3123 ( .A1(n2432), .A2(n2431), .A3(n2430), .A4(n2429), .ZN(n4316)
         );
  NAND2_X1 U3124 ( .A1(n2476), .A2(IR_REG_31__SCAN_IN), .ZN(n2435) );
  XNOR2_X1 U3125 ( .A(n2435), .B(IR_REG_14__SCAN_IN), .ZN(n4612) );
  MUX2_X1 U3126 ( .A(n4612), .B(DATAI_14_), .S(n2310), .Z(n4466) );
  NAND2_X1 U3127 ( .A1(n4462), .A2(n4466), .ZN(n4304) );
  NAND2_X1 U3128 ( .A1(n4316), .A2(n4338), .ZN(n3635) );
  NAND2_X1 U3129 ( .A1(n4304), .A2(n3635), .ZN(n4334) );
  INV_X1 U3130 ( .A(n4334), .ZN(n2450) );
  OR2_X1 U3131 ( .A1(n4324), .A2(n2450), .ZN(n4308) );
  NAND2_X1 U3132 ( .A1(n2304), .A2(REG1_REG_15__SCAN_IN), .ZN(n2441) );
  NAND2_X1 U3133 ( .A1(n2303), .A2(REG0_REG_15__SCAN_IN), .ZN(n2440) );
  NAND2_X1 U3134 ( .A1(n2456), .A2(REG2_REG_15__SCAN_IN), .ZN(n2439) );
  NOR2_X1 U3135 ( .A1(n2436), .A2(REG3_REG_15__SCAN_IN), .ZN(n2437) );
  OR2_X1 U3136 ( .A1(n2466), .A2(n2437), .ZN(n3629) );
  OR2_X1 U3137 ( .A1(n2535), .A2(n3629), .ZN(n2438) );
  NAND4_X1 U3138 ( .A1(n2441), .A2(n2440), .A3(n2439), .A4(n2438), .ZN(n4467)
         );
  OR2_X1 U3139 ( .A1(n2476), .A2(IR_REG_14__SCAN_IN), .ZN(n2442) );
  NAND2_X1 U3140 ( .A1(n2442), .A2(IR_REG_31__SCAN_IN), .ZN(n2462) );
  XNOR2_X1 U3141 ( .A(n2462), .B(IR_REG_15__SCAN_IN), .ZN(n4071) );
  MUX2_X1 U3142 ( .A(n4071), .B(DATAI_15_), .S(n2051), .Z(n4458) );
  AND2_X1 U3143 ( .A1(n4467), .A2(n4458), .ZN(n2452) );
  OR2_X1 U3144 ( .A1(n4308), .A2(n2452), .ZN(n2443) );
  INV_X1 U3145 ( .A(n4467), .ZN(n4345) );
  INV_X1 U3146 ( .A(n4458), .ZN(n4314) );
  NAND2_X1 U3147 ( .A1(n4345), .A2(n4314), .ZN(n2454) );
  NAND2_X1 U31480 ( .A1(n4462), .A2(n4338), .ZN(n2451) );
  OR2_X1 U31490 ( .A1(n4481), .A2(n3558), .ZN(n2447) );
  NAND2_X1 U3150 ( .A1(n4485), .A2(n4499), .ZN(n3295) );
  INV_X1 U3151 ( .A(n4496), .ZN(n2589) );
  INV_X1 U3152 ( .A(n3457), .ZN(n4479) );
  NAND2_X1 U3153 ( .A1(n2589), .A2(n4479), .ZN(n2444) );
  AND2_X1 U3154 ( .A1(n3295), .A2(n2444), .ZN(n2445) );
  OR2_X1 U3155 ( .A1(n2446), .A2(n2445), .ZN(n4353) );
  AND2_X1 U3156 ( .A1(n2447), .A2(n4353), .ZN(n2448) );
  OR2_X1 U3157 ( .A1(n2450), .A2(n4325), .ZN(n4327) );
  AND2_X1 U3158 ( .A1(n2451), .A2(n4327), .ZN(n4309) );
  OR2_X1 U3159 ( .A1(n2452), .A2(n4309), .ZN(n2453) );
  NAND2_X1 U3160 ( .A1(n2304), .A2(REG1_REG_16__SCAN_IN), .ZN(n2460) );
  NAND2_X1 U3161 ( .A1(n2303), .A2(REG0_REG_16__SCAN_IN), .ZN(n2459) );
  NAND2_X1 U3162 ( .A1(n2456), .A2(REG2_REG_16__SCAN_IN), .ZN(n2458) );
  XNOR2_X1 U3163 ( .A(n2466), .B(REG3_REG_16__SCAN_IN), .ZN(n4292) );
  OR2_X1 U3164 ( .A1(n2535), .A2(n4292), .ZN(n2457) );
  NAND4_X1 U3165 ( .A1(n2460), .A2(n2459), .A3(n2458), .A4(n2457), .ZN(n4459)
         );
  INV_X1 U3166 ( .A(n4459), .ZN(n4450) );
  INV_X1 U3167 ( .A(IR_REG_15__SCAN_IN), .ZN(n2461) );
  NAND2_X1 U3168 ( .A1(n2462), .A2(n2461), .ZN(n2463) );
  NAND2_X1 U3169 ( .A1(n2463), .A2(IR_REG_31__SCAN_IN), .ZN(n2464) );
  XNOR2_X1 U3170 ( .A(n2464), .B(IR_REG_16__SCAN_IN), .ZN(n4076) );
  MUX2_X1 U3171 ( .A(n4076), .B(DATAI_16_), .S(n2310), .Z(n4289) );
  NAND2_X1 U3172 ( .A1(n4450), .A2(n4289), .ZN(n3715) );
  INV_X1 U3173 ( .A(n4289), .ZN(n4299) );
  NAND2_X1 U3174 ( .A1(n4459), .A2(n4299), .ZN(n3717) );
  NAND2_X1 U3175 ( .A1(n4459), .A2(n4289), .ZN(n2465) );
  NAND2_X1 U3176 ( .A1(n2304), .A2(REG1_REG_17__SCAN_IN), .ZN(n2473) );
  NAND2_X1 U3177 ( .A1(n2303), .A2(REG0_REG_17__SCAN_IN), .ZN(n2472) );
  NAND2_X1 U3178 ( .A1(n2456), .A2(REG2_REG_17__SCAN_IN), .ZN(n2471) );
  NAND2_X1 U3179 ( .A1(n2466), .A2(REG3_REG_16__SCAN_IN), .ZN(n2468) );
  INV_X1 U3180 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2467) );
  NAND2_X1 U3181 ( .A1(n2468), .A2(n2467), .ZN(n2469) );
  NAND2_X1 U3182 ( .A1(n2469), .A2(n2481), .ZN(n3501) );
  OR2_X1 U3183 ( .A1(n2535), .A2(n3501), .ZN(n2470) );
  NAND4_X1 U3184 ( .A1(n2473), .A2(n2472), .A3(n2471), .A4(n2470), .ZN(n4296)
         );
  INV_X1 U3185 ( .A(n4296), .ZN(n4264) );
  INV_X1 U3186 ( .A(n2474), .ZN(n2475) );
  NAND2_X1 U3187 ( .A1(n2487), .A2(IR_REG_31__SCAN_IN), .ZN(n2477) );
  INV_X1 U3188 ( .A(DATAI_17_), .ZN(n2478) );
  MUX2_X1 U3189 ( .A(n4754), .B(n2478), .S(n2310), .Z(n4277) );
  NAND2_X1 U3190 ( .A1(n4264), .A2(n4277), .ZN(n2479) );
  INV_X1 U3191 ( .A(n4277), .ZN(n4446) );
  NAND2_X1 U3192 ( .A1(n2304), .A2(REG1_REG_18__SCAN_IN), .ZN(n2486) );
  NAND2_X1 U3193 ( .A1(n2303), .A2(REG0_REG_18__SCAN_IN), .ZN(n2485) );
  NAND2_X1 U3194 ( .A1(n2456), .A2(REG2_REG_18__SCAN_IN), .ZN(n2484) );
  NAND2_X1 U3195 ( .A1(n2481), .A2(n2480), .ZN(n2482) );
  NAND2_X1 U3196 ( .A1(n2493), .A2(n2482), .ZN(n3592) );
  OR2_X1 U3197 ( .A1(n2535), .A2(n3592), .ZN(n2483) );
  NAND4_X1 U3198 ( .A1(n2486), .A2(n2485), .A3(n2484), .A4(n2483), .ZN(n4447)
         );
  INV_X1 U3199 ( .A(n4447), .ZN(n4281) );
  NAND2_X1 U3200 ( .A1(n2499), .A2(IR_REG_31__SCAN_IN), .ZN(n2490) );
  XNOR2_X1 U3201 ( .A(n2490), .B(IR_REG_18__SCAN_IN), .ZN(n4069) );
  MUX2_X1 U3202 ( .A(n4069), .B(DATAI_18_), .S(n2051), .Z(n4262) );
  NAND2_X1 U3203 ( .A1(n4281), .A2(n4262), .ZN(n4237) );
  NAND2_X1 U3204 ( .A1(n4447), .A2(n4259), .ZN(n4235) );
  NAND2_X1 U3205 ( .A1(n4237), .A2(n4235), .ZN(n4260) );
  NAND2_X1 U3206 ( .A1(n4281), .A2(n4259), .ZN(n2491) );
  NAND2_X1 U3207 ( .A1(n2304), .A2(REG1_REG_19__SCAN_IN), .ZN(n2498) );
  NAND2_X1 U3208 ( .A1(n2303), .A2(REG0_REG_19__SCAN_IN), .ZN(n2497) );
  NAND2_X1 U3209 ( .A1(n2456), .A2(REG2_REG_19__SCAN_IN), .ZN(n2496) );
  AND2_X1 U32100 ( .A1(n2493), .A2(n2492), .ZN(n2494) );
  OR2_X1 U32110 ( .A1(n2494), .A2(n2503), .ZN(n4248) );
  OR2_X1 U32120 ( .A1(n2535), .A2(n4248), .ZN(n2495) );
  NAND4_X1 U32130 ( .A1(n2498), .A2(n2497), .A3(n2496), .A4(n2495), .ZN(n4433)
         );
  MUX2_X1 U32140 ( .A(n4611), .B(DATAI_19_), .S(n2310), .Z(n3422) );
  NOR2_X1 U32150 ( .A1(n4433), .A2(n3422), .ZN(n4214) );
  NAND2_X1 U32160 ( .A1(n2304), .A2(REG1_REG_20__SCAN_IN), .ZN(n2508) );
  NAND2_X1 U32170 ( .A1(n2303), .A2(REG0_REG_20__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U32180 ( .A1(n2456), .A2(REG2_REG_20__SCAN_IN), .ZN(n2506) );
  NOR2_X1 U32190 ( .A1(n2503), .A2(REG3_REG_20__SCAN_IN), .ZN(n2504) );
  OR2_X1 U32200 ( .A1(n2516), .A2(n2504), .ZN(n3547) );
  OR2_X1 U32210 ( .A1(n2535), .A2(n3547), .ZN(n2505) );
  NAND2_X1 U32220 ( .A1(n4242), .A2(n3546), .ZN(n3750) );
  NAND2_X1 U32230 ( .A1(n4433), .A2(n3422), .ZN(n4215) );
  INV_X1 U32240 ( .A(n4242), .ZN(n4426) );
  NAND2_X1 U32250 ( .A1(n4426), .A2(n4430), .ZN(n3751) );
  NAND2_X1 U32260 ( .A1(n2509), .A2(n3751), .ZN(n4198) );
  NAND2_X1 U32270 ( .A1(n2304), .A2(REG1_REG_21__SCAN_IN), .ZN(n2513) );
  NAND2_X1 U32280 ( .A1(n2303), .A2(REG0_REG_21__SCAN_IN), .ZN(n2512) );
  NAND2_X1 U32290 ( .A1(n2456), .A2(REG2_REG_21__SCAN_IN), .ZN(n2511) );
  XNOR2_X1 U32300 ( .A(n2516), .B(REG3_REG_21__SCAN_IN), .ZN(n3445) );
  OR2_X1 U32310 ( .A1(n2535), .A2(n3445), .ZN(n2510) );
  NAND4_X1 U32320 ( .A1(n2513), .A2(n2512), .A3(n2511), .A4(n2510), .ZN(n4220)
         );
  NAND2_X1 U32330 ( .A1(n4220), .A2(n4422), .ZN(n2514) );
  INV_X1 U32340 ( .A(n4220), .ZN(n4431) );
  NAND2_X1 U32350 ( .A1(n4431), .A2(n4202), .ZN(n2515) );
  NAND2_X1 U32360 ( .A1(n2304), .A2(REG1_REG_22__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U32370 ( .A1(n2303), .A2(REG0_REG_22__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U32380 ( .A1(n2456), .A2(REG2_REG_22__SCAN_IN), .ZN(n2521) );
  NAND2_X1 U32390 ( .A1(n2516), .A2(REG3_REG_21__SCAN_IN), .ZN(n2518) );
  INV_X1 U32400 ( .A(REG3_REG_22__SCAN_IN), .ZN(n2517) );
  NAND2_X1 U32410 ( .A1(n2518), .A2(n2517), .ZN(n2519) );
  NAND2_X1 U32420 ( .A1(n2519), .A2(n2525), .ZN(n4182) );
  OR2_X1 U32430 ( .A1(n2535), .A2(n4182), .ZN(n2520) );
  NAND4_X1 U32440 ( .A1(n2523), .A2(n2522), .A3(n2521), .A4(n2520), .ZN(n4423)
         );
  NAND2_X1 U32450 ( .A1(n4207), .A2(n2524), .ZN(n4161) );
  NAND2_X1 U32460 ( .A1(n4423), .A2(n4191), .ZN(n2601) );
  NAND2_X1 U32470 ( .A1(n2303), .A2(REG0_REG_23__SCAN_IN), .ZN(n2530) );
  NAND2_X1 U32480 ( .A1(n2330), .A2(REG2_REG_23__SCAN_IN), .ZN(n2529) );
  NAND2_X1 U32490 ( .A1(n2304), .A2(REG1_REG_23__SCAN_IN), .ZN(n2528) );
  NAND2_X1 U32500 ( .A1(n2525), .A2(n3385), .ZN(n2526) );
  NAND2_X1 U32510 ( .A1(n2533), .A2(n2526), .ZN(n3387) );
  OR2_X1 U32520 ( .A1(n2535), .A2(n3387), .ZN(n2527) );
  INV_X1 U32530 ( .A(n4188), .ZN(n4408) );
  NAND2_X1 U32540 ( .A1(n4408), .A2(n4168), .ZN(n2531) );
  NAND2_X1 U32550 ( .A1(n2304), .A2(REG1_REG_24__SCAN_IN), .ZN(n2539) );
  NAND2_X1 U32560 ( .A1(n2303), .A2(REG0_REG_24__SCAN_IN), .ZN(n2538) );
  NAND2_X1 U32570 ( .A1(n2330), .A2(REG2_REG_24__SCAN_IN), .ZN(n2537) );
  NAND2_X1 U32580 ( .A1(n2533), .A2(n2532), .ZN(n2534) );
  NAND2_X1 U32590 ( .A1(n2542), .A2(n2534), .ZN(n3512) );
  OR2_X1 U32600 ( .A1(n2535), .A2(n3512), .ZN(n2536) );
  NAND4_X1 U32610 ( .A1(n2539), .A2(n2538), .A3(n2537), .A4(n2536), .ZN(n4130)
         );
  INV_X1 U32620 ( .A(n4147), .ZN(n4404) );
  NAND2_X1 U32630 ( .A1(n4130), .A2(n4404), .ZN(n2540) );
  INV_X1 U32640 ( .A(n2535), .ZN(n2544) );
  AND2_X1 U32650 ( .A1(n2542), .A2(n2541), .ZN(n2543) );
  NOR2_X1 U32660 ( .A1(n2550), .A2(n2543), .ZN(n4131) );
  NAND2_X1 U32670 ( .A1(n2544), .A2(n4131), .ZN(n2548) );
  NAND2_X1 U32680 ( .A1(n2304), .A2(REG1_REG_25__SCAN_IN), .ZN(n2547) );
  NAND2_X1 U32690 ( .A1(n2303), .A2(REG0_REG_25__SCAN_IN), .ZN(n2546) );
  NAND2_X1 U32700 ( .A1(n2456), .A2(REG2_REG_25__SCAN_IN), .ZN(n2545) );
  INV_X1 U32710 ( .A(n4405), .ZN(n4151) );
  NAND2_X1 U32720 ( .A1(n4151), .A2(n4128), .ZN(n2549) );
  NOR2_X1 U32730 ( .A1(n2550), .A2(REG3_REG_26__SCAN_IN), .ZN(n2551) );
  NAND2_X1 U32740 ( .A1(n2304), .A2(REG1_REG_26__SCAN_IN), .ZN(n2554) );
  NAND2_X1 U32750 ( .A1(n2303), .A2(REG0_REG_26__SCAN_IN), .ZN(n2553) );
  AND2_X1 U32760 ( .A1(n2554), .A2(n2553), .ZN(n2556) );
  NAND2_X1 U32770 ( .A1(n2330), .A2(REG2_REG_26__SCAN_IN), .ZN(n2555) );
  OAI211_X2 U32780 ( .C1(n3615), .C2(n2535), .A(n2556), .B(n2555), .ZN(n4396)
         );
  NOR2_X1 U32790 ( .A1(n4396), .A2(n3614), .ZN(n3741) );
  NAND2_X1 U32800 ( .A1(n2557), .A2(REG3_REG_28__SCAN_IN), .ZN(n3330) );
  INV_X1 U32810 ( .A(n2557), .ZN(n2559) );
  INV_X1 U32820 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2558) );
  NAND2_X1 U32830 ( .A1(n2559), .A2(n2558), .ZN(n2560) );
  NAND2_X1 U32840 ( .A1(n3330), .A2(n2560), .ZN(n2908) );
  OR2_X1 U32850 ( .A1(n2908), .A2(n2535), .ZN(n2563) );
  AOI22_X1 U32860 ( .A1(n2304), .A2(REG1_REG_28__SCAN_IN), .B1(n2303), .B2(
        REG0_REG_28__SCAN_IN), .ZN(n2562) );
  NAND2_X1 U32870 ( .A1(n2330), .A2(REG2_REG_28__SCAN_IN), .ZN(n2561) );
  NAND2_X1 U32880 ( .A1(n3802), .A2(n2896), .ZN(n3660) );
  INV_X1 U32890 ( .A(n2896), .ZN(n3338) );
  NAND2_X1 U32900 ( .A1(n4386), .A2(n3338), .ZN(n3651) );
  NAND2_X1 U32910 ( .A1(n3660), .A2(n3651), .ZN(n3743) );
  XNOR2_X1 U32920 ( .A(n2649), .B(n3743), .ZN(n3347) );
  NAND2_X1 U32930 ( .A1(n2567), .A2(IR_REG_31__SCAN_IN), .ZN(n2568) );
  MUX2_X1 U32940 ( .A(IR_REG_31__SCAN_IN), .B(n2568), .S(IR_REG_21__SCAN_IN), 
        .Z(n2571) );
  INV_X1 U32950 ( .A(n2569), .ZN(n2570) );
  NAND2_X1 U32960 ( .A1(n2570), .A2(IR_REG_31__SCAN_IN), .ZN(n2572) );
  XNOR2_X1 U32970 ( .A(n3097), .B(n4609), .ZN(n2573) );
  NAND2_X1 U32980 ( .A1(n2573), .A2(n4087), .ZN(n4524) );
  NAND2_X1 U32990 ( .A1(n2639), .A2(n4611), .ZN(n3088) );
  INV_X1 U33000 ( .A(n4492), .ZN(n4781) );
  OR2_X1 U33010 ( .A1(n2574), .A2(n2982), .ZN(n2576) );
  INV_X1 U33020 ( .A(n2939), .ZN(n2902) );
  NOR2_X2 U33030 ( .A1(n4617), .A2(n2902), .ZN(n4519) );
  INV_X1 U33040 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3336) );
  OR2_X1 U33050 ( .A1(n3330), .A2(n2535), .ZN(n2578) );
  AOI22_X1 U33060 ( .A1(REG1_REG_29__SCAN_IN), .A2(n2304), .B1(n2303), .B2(
        REG0_REG_29__SCAN_IN), .ZN(n2577) );
  OAI211_X1 U33070 ( .C1(n2579), .C2(n3336), .A(n2578), .B(n2577), .ZN(n3801)
         );
  INV_X1 U33080 ( .A(n3801), .ZN(n3650) );
  NAND2_X1 U33090 ( .A1(n4617), .A2(n2939), .ZN(n4522) );
  INV_X1 U33100 ( .A(n2639), .ZN(n4610) );
  INV_X1 U33110 ( .A(n4609), .ZN(n2580) );
  INV_X1 U33120 ( .A(n3786), .ZN(n2921) );
  OAI22_X1 U33130 ( .A1(n3650), .A2(n4522), .B1(n4500), .B2(n2896), .ZN(n2581)
         );
  AOI21_X1 U33140 ( .B1(n4519), .B2(n4110), .A(n2581), .ZN(n2609) );
  INV_X1 U33150 ( .A(n3983), .ZN(n3076) );
  NAND2_X1 U33160 ( .A1(n3076), .A2(n2677), .ZN(n3676) );
  NAND2_X1 U33170 ( .A1(n3142), .A2(n3762), .ZN(n3141) );
  NAND2_X1 U33180 ( .A1(n3141), .A2(n3681), .ZN(n3156) );
  NAND2_X1 U33190 ( .A1(n3144), .A2(n3414), .ZN(n3686) );
  NAND2_X1 U33200 ( .A1(n3981), .A2(n2699), .ZN(n3683) );
  INV_X1 U33210 ( .A(n3687), .ZN(n2584) );
  NAND2_X1 U33220 ( .A1(n2585), .A2(n3489), .ZN(n3698) );
  NAND2_X1 U33230 ( .A1(n3805), .A2(n2124), .ZN(n3699) );
  NAND2_X1 U33240 ( .A1(n3168), .A2(n3699), .ZN(n2586) );
  NAND2_X1 U33250 ( .A1(n2125), .A2(n3604), .ZN(n3691) );
  NAND2_X1 U33260 ( .A1(n3804), .A2(n4509), .ZN(n3774) );
  NAND2_X1 U33270 ( .A1(n3282), .A2(n4517), .ZN(n3775) );
  AND2_X1 U33280 ( .A1(n3434), .A2(n3278), .ZN(n3696) );
  NAND2_X1 U33290 ( .A1(n4523), .A2(n3533), .ZN(n3694) );
  NAND2_X1 U33300 ( .A1(n4494), .A2(n3305), .ZN(n3706) );
  NAND2_X1 U33310 ( .A1(n3256), .A2(n3706), .ZN(n2588) );
  NAND2_X1 U33320 ( .A1(n2587), .A2(n3404), .ZN(n3700) );
  NAND2_X1 U33330 ( .A1(n4496), .A2(n4479), .ZN(n4357) );
  NAND2_X1 U33340 ( .A1(n4481), .A2(n4365), .ZN(n3752) );
  NAND2_X1 U33350 ( .A1(n4357), .A2(n3752), .ZN(n2591) );
  NAND2_X1 U33360 ( .A1(n2589), .A2(n3457), .ZN(n4356) );
  NAND2_X1 U33370 ( .A1(n3291), .A2(n4356), .ZN(n2590) );
  INV_X1 U33380 ( .A(n2591), .ZN(n3708) );
  NOR2_X1 U33390 ( .A1(n4481), .A2(n4365), .ZN(n3753) );
  AOI21_X1 U33400 ( .B1(n2590), .B2(n3708), .A(n3753), .ZN(n3709) );
  NAND2_X1 U33410 ( .A1(n4345), .A2(n4458), .ZN(n3637) );
  NAND2_X1 U33420 ( .A1(n4467), .A2(n4314), .ZN(n3636) );
  NAND2_X1 U33430 ( .A1(n3637), .A2(n3636), .ZN(n4310) );
  INV_X1 U33440 ( .A(n4304), .ZN(n2592) );
  NAND2_X1 U33450 ( .A1(n2593), .A2(n3636), .ZN(n4295) );
  INV_X1 U33460 ( .A(n3717), .ZN(n3639) );
  NAND2_X1 U33470 ( .A1(n4296), .A2(n4277), .ZN(n3755) );
  INV_X1 U33480 ( .A(n3422), .ZN(n4246) );
  NAND2_X1 U33490 ( .A1(n4433), .A2(n4246), .ZN(n2594) );
  AND2_X1 U33500 ( .A1(n4235), .A2(n2594), .ZN(n3638) );
  NAND2_X1 U33510 ( .A1(n4264), .A2(n4446), .ZN(n4232) );
  NAND2_X1 U33520 ( .A1(n4237), .A2(n4232), .ZN(n2595) );
  NAND2_X1 U3353 ( .A1(n2595), .A2(n3638), .ZN(n2597) );
  INV_X1 U33540 ( .A(n4433), .ZN(n2833) );
  NAND2_X1 U3355 ( .A1(n2833), .A2(n3422), .ZN(n2596) );
  NAND2_X1 U3356 ( .A1(n2597), .A2(n2596), .ZN(n4212) );
  NOR2_X1 U3357 ( .A1(n4242), .A2(n4430), .ZN(n2598) );
  OR2_X1 U3358 ( .A1(n4212), .A2(n2598), .ZN(n2599) );
  NAND2_X1 U3359 ( .A1(n2599), .A2(n2080), .ZN(n4157) );
  NAND2_X1 U3360 ( .A1(n4431), .A2(n4422), .ZN(n4159) );
  AND2_X1 U3361 ( .A1(n4161), .A2(n4159), .ZN(n3723) );
  AND2_X1 U3362 ( .A1(n4157), .A2(n3723), .ZN(n3641) );
  NAND2_X1 U3363 ( .A1(n4188), .A2(n4168), .ZN(n2600) );
  AND2_X1 U3364 ( .A1(n2601), .A2(n2600), .ZN(n3727) );
  AND2_X1 U3365 ( .A1(n4220), .A2(n4202), .ZN(n3721) );
  NAND2_X1 U3366 ( .A1(n4161), .A2(n3721), .ZN(n2602) );
  AND2_X1 U3367 ( .A1(n3727), .A2(n2602), .ZN(n3642) );
  NAND2_X1 U3368 ( .A1(n2603), .A2(n3642), .ZN(n4140) );
  NAND2_X1 U3369 ( .A1(n4399), .A2(n4404), .ZN(n3746) );
  NAND2_X1 U3370 ( .A1(n4408), .A2(n3780), .ZN(n4139) );
  AND2_X1 U3371 ( .A1(n4130), .A2(n4147), .ZN(n3646) );
  INV_X1 U3372 ( .A(n3646), .ZN(n3747) );
  AND2_X1 U3373 ( .A1(n4405), .A2(n4128), .ZN(n3744) );
  INV_X1 U3374 ( .A(n3744), .ZN(n2604) );
  OR2_X1 U3375 ( .A1(n4405), .A2(n4128), .ZN(n3647) );
  NAND2_X1 U3376 ( .A1(n2605), .A2(n3647), .ZN(n4108) );
  NOR2_X1 U3377 ( .A1(n4396), .A2(n4116), .ZN(n3648) );
  NAND2_X1 U3378 ( .A1(n4396), .A2(n4116), .ZN(n3657) );
  XNOR2_X1 U3379 ( .A(n4110), .B(n4098), .ZN(n4095) );
  OR2_X1 U3380 ( .A1(n4110), .A2(n4098), .ZN(n3658) );
  INV_X1 U3381 ( .A(n3743), .ZN(n2606) );
  XNOR2_X1 U3382 ( .A(n2651), .B(n2606), .ZN(n2608) );
  NAND2_X1 U3383 ( .A1(n4610), .A2(n3786), .ZN(n3672) );
  NAND2_X1 U3384 ( .A1(n4611), .A2(n4609), .ZN(n2607) );
  NAND2_X1 U3385 ( .A1(n2608), .A2(n4529), .ZN(n3342) );
  OAI211_X1 U3386 ( .C1(n3347), .C2(n4781), .A(n2609), .B(n3342), .ZN(n2645)
         );
  NAND2_X1 U3387 ( .A1(n2610), .A2(IR_REG_31__SCAN_IN), .ZN(n2611) );
  MUX2_X1 U3388 ( .A(IR_REG_31__SCAN_IN), .B(n2611), .S(IR_REG_25__SCAN_IN), 
        .Z(n2612) );
  NAND2_X1 U3389 ( .A1(n2612), .A2(n2064), .ZN(n2619) );
  NAND2_X1 U3390 ( .A1(n2619), .A2(B_REG_SCAN_IN), .ZN(n2616) );
  OR2_X1 U3391 ( .A1(n2613), .A2(n2982), .ZN(n2621) );
  NAND2_X1 U3392 ( .A1(n2621), .A2(n2620), .ZN(n2614) );
  MUX2_X1 U3393 ( .A(n2616), .B(B_REG_SCAN_IN), .S(n4608), .Z(n2618) );
  NAND2_X1 U3394 ( .A1(n2064), .A2(IR_REG_31__SCAN_IN), .ZN(n2617) );
  INV_X1 U3395 ( .A(n4607), .ZN(n2978) );
  NAND2_X1 U3396 ( .A1(n2978), .A2(n2619), .ZN(n2974) );
  NAND2_X1 U3397 ( .A1(n2900), .A2(n2974), .ZN(n2636) );
  INV_X1 U3398 ( .A(n2619), .ZN(n2968) );
  NAND2_X1 U3399 ( .A1(n2639), .A2(n4087), .ZN(n2622) );
  NAND2_X1 U3400 ( .A1(n2622), .A2(n2939), .ZN(n3093) );
  OAI211_X1 U3401 ( .C1(n3113), .C2(n3786), .A(n3090), .B(n3093), .ZN(n2623)
         );
  INV_X1 U3402 ( .A(n2623), .ZN(n2635) );
  NOR4_X1 U3403 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_17__SCAN_IN), .A4(D_REG_18__SCAN_IN), .ZN(n2627) );
  NOR4_X1 U3404 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2626) );
  NOR4_X1 U3405 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2625) );
  NOR4_X1 U3406 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_22__SCAN_IN), .ZN(n2624) );
  NAND4_X1 U3407 ( .A1(n2627), .A2(n2626), .A3(n2625), .A4(n2624), .ZN(n2633)
         );
  NOR2_X1 U3408 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_9__SCAN_IN), .ZN(n2631) );
  NOR4_X1 U3409 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2630) );
  NOR4_X1 U3410 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2629) );
  NOR4_X1 U3411 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2628) );
  NAND4_X1 U3412 ( .A1(n2631), .A2(n2630), .A3(n2629), .A4(n2628), .ZN(n2632)
         );
  NOR2_X1 U3413 ( .A1(n2633), .A2(n2632), .ZN(n2634) );
  INV_X1 U3414 ( .A(n4608), .ZN(n2977) );
  NAND2_X1 U3415 ( .A1(n2978), .A2(n2977), .ZN(n2637) );
  NAND2_X1 U3416 ( .A1(n3111), .A2(n3112), .ZN(n3150) );
  OAI21_X1 U3417 ( .B1(n4096), .B2(n2896), .A(n2662), .ZN(n3337) );
  NAND2_X1 U3418 ( .A1(n2645), .A2(n4795), .ZN(n2648) );
  NAND2_X1 U3419 ( .A1(n4792), .A2(REG1_REG_28__SCAN_IN), .ZN(n2646) );
  NAND2_X1 U3420 ( .A1(n2648), .A2(n2264), .ZN(U3546) );
  INV_X1 U3421 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2661) );
  NAND2_X1 U3422 ( .A1(n2051), .A2(DATAI_29_), .ZN(n3656) );
  XNOR2_X1 U3423 ( .A(n3801), .B(n3656), .ZN(n3779) );
  INV_X1 U3424 ( .A(n3651), .ZN(n3659) );
  INV_X1 U3425 ( .A(n2652), .ZN(n2653) );
  XNOR2_X1 U3426 ( .A(n2653), .B(n3779), .ZN(n2660) );
  NAND2_X1 U3427 ( .A1(n3802), .A2(n4519), .ZN(n2659) );
  NAND2_X1 U3428 ( .A1(n2304), .A2(REG1_REG_30__SCAN_IN), .ZN(n2656) );
  NAND2_X1 U3429 ( .A1(n2330), .A2(REG2_REG_30__SCAN_IN), .ZN(n2655) );
  NAND2_X1 U3430 ( .A1(n2303), .A2(REG0_REG_30__SCAN_IN), .ZN(n2654) );
  NAND3_X1 U3431 ( .A1(n2656), .A2(n2655), .A3(n2654), .ZN(n3800) );
  XNOR2_X1 U3432 ( .A(n2657), .B(n2255), .ZN(n4606) );
  AOI21_X1 U3433 ( .B1(B_REG_SCAN_IN), .B2(n4606), .A(n4522), .ZN(n3320) );
  AOI22_X1 U3434 ( .A1(n3800), .A2(n3320), .B1(n3649), .B2(n4518), .ZN(n2658)
         );
  OAI21_X1 U3435 ( .B1(n2660), .B2(n4505), .A(n2262), .ZN(n3333) );
  AOI21_X1 U3436 ( .B1(n3329), .B2(n4492), .A(n3333), .ZN(n2665) );
  MUX2_X1 U3437 ( .A(n2661), .B(n2665), .S(n4789), .Z(n2664) );
  NAND2_X1 U3438 ( .A1(n2664), .A2(n2663), .ZN(U3515) );
  INV_X1 U3439 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2666) );
  MUX2_X1 U3440 ( .A(n2666), .B(n2665), .S(n4795), .Z(n2668) );
  NAND2_X1 U3441 ( .A1(n2668), .A2(n2667), .ZN(U3547) );
  AND2_X2 U3442 ( .A1(n3097), .A2(n2937), .ZN(n2674) );
  NAND2_X1 U3443 ( .A1(n3078), .A2(n2674), .ZN(n2669) );
  NAND2_X1 U3444 ( .A1(n2670), .A2(n2669), .ZN(n2671) );
  NAND2_X1 U3445 ( .A1(n4087), .A2(n4609), .ZN(n2913) );
  INV_X1 U3446 ( .A(n4258), .ZN(n3229) );
  AND2_X4 U3447 ( .A1(n2674), .A2(n3229), .ZN(n2891) );
  NOR2_X1 U3448 ( .A1(n3111), .A2(n2710), .ZN(n2672) );
  AOI21_X1 U3449 ( .B1(n2673), .B2(n2891), .A(n2672), .ZN(n2682) );
  XNOR2_X1 U3450 ( .A(n2684), .B(n2682), .ZN(n3073) );
  NOR2_X1 U3451 ( .A1(n3112), .A2(n2895), .ZN(n2675) );
  INV_X1 U3452 ( .A(REG1_REG_0__SCAN_IN), .ZN(n3985) );
  OR2_X1 U3453 ( .A1(n2937), .A2(n3985), .ZN(n2676) );
  NAND2_X1 U3454 ( .A1(n2680), .A2(n2676), .ZN(n3064) );
  NAND2_X1 U3455 ( .A1(n3983), .A2(n2891), .ZN(n2679) );
  AOI22_X1 U3456 ( .A1(n2677), .A2(n2731), .B1(IR_REG_0__SCAN_IN), .B2(n2204), 
        .ZN(n2678) );
  NAND2_X1 U3457 ( .A1(n2679), .A2(n2678), .ZN(n3063) );
  NAND2_X1 U34580 ( .A1(n3064), .A2(n3063), .ZN(n3062) );
  NAND2_X1 U34590 ( .A1(n2680), .A2(n2893), .ZN(n2681) );
  NAND2_X1 U3460 ( .A1(n3062), .A2(n2681), .ZN(n3072) );
  NAND2_X1 U3461 ( .A1(n3073), .A2(n3072), .ZN(n3071) );
  INV_X1 U3462 ( .A(n2682), .ZN(n2683) );
  NAND2_X1 U3463 ( .A1(n2684), .A2(n2683), .ZN(n2685) );
  NAND2_X1 U3464 ( .A1(n3071), .A2(n2685), .ZN(n3118) );
  INV_X1 U3465 ( .A(n3118), .ZN(n2692) );
  NAND2_X1 U3466 ( .A1(n2690), .A2(n2731), .ZN(n2687) );
  NAND2_X1 U34670 ( .A1(n3151), .A2(n2674), .ZN(n2686) );
  NAND2_X1 U3468 ( .A1(n2687), .A2(n2686), .ZN(n2688) );
  XNOR2_X1 U34690 ( .A(n2688), .B(n2893), .ZN(n2694) );
  NOR2_X1 U3470 ( .A1(n3121), .A2(n2710), .ZN(n2689) );
  XNOR2_X1 U34710 ( .A(n2694), .B(n2693), .ZN(n3119) );
  INV_X1 U3472 ( .A(n3119), .ZN(n2691) );
  NAND2_X1 U34730 ( .A1(n2692), .A2(n2691), .ZN(n3116) );
  NAND2_X1 U3474 ( .A1(n2694), .A2(n2693), .ZN(n2695) );
  NAND2_X1 U34750 ( .A1(n3116), .A2(n2695), .ZN(n3411) );
  NAND2_X1 U3476 ( .A1(n3981), .A2(n2880), .ZN(n2697) );
  NAND2_X1 U34770 ( .A1(n3414), .A2(n2674), .ZN(n2696) );
  NAND2_X1 U3478 ( .A1(n2697), .A2(n2696), .ZN(n2698) );
  XNOR2_X1 U34790 ( .A(n2698), .B(n2874), .ZN(n2701) );
  NOR2_X1 U3480 ( .A1(n2699), .A2(n2710), .ZN(n2700) );
  AOI21_X1 U34810 ( .B1(n3981), .B2(n2891), .A(n2700), .ZN(n2702) );
  XNOR2_X1 U3482 ( .A(n2701), .B(n2702), .ZN(n3410) );
  NAND2_X1 U34830 ( .A1(n3411), .A2(n3410), .ZN(n2705) );
  INV_X1 U3484 ( .A(n2701), .ZN(n2703) );
  NAND2_X1 U34850 ( .A1(n2703), .A2(n2702), .ZN(n2704) );
  NAND2_X1 U3486 ( .A1(n2705), .A2(n2704), .ZN(n3481) );
  INV_X1 U34870 ( .A(n3481), .ZN(n2716) );
  NAND2_X1 U3488 ( .A1(n3806), .A2(n2880), .ZN(n2707) );
  NAND2_X1 U34890 ( .A1(n3521), .A2(n2674), .ZN(n2706) );
  NAND2_X1 U3490 ( .A1(n2707), .A2(n2706), .ZN(n2708) );
  XNOR2_X1 U34910 ( .A(n2708), .B(n2893), .ZN(n2719) );
  NOR2_X1 U3492 ( .A1(n3211), .A2(n2710), .ZN(n2709) );
  AOI21_X1 U34930 ( .B1(n3806), .B2(n2891), .A(n2709), .ZN(n2720) );
  XNOR2_X1 U3494 ( .A(n2719), .B(n2720), .ZN(n3518) );
  NAND2_X1 U34950 ( .A1(n3603), .A2(n2880), .ZN(n2712) );
  NAND2_X1 U3496 ( .A1(n3489), .A2(n2674), .ZN(n2711) );
  NAND2_X1 U34970 ( .A1(n2712), .A2(n2711), .ZN(n2713) );
  NOR2_X1 U3498 ( .A1(n2714), .A2(n2710), .ZN(n2715) );
  AOI21_X1 U34990 ( .B1(n3603), .B2(n2891), .A(n2715), .ZN(n2717) );
  NAND2_X1 U3500 ( .A1(n2716), .A2(n2067), .ZN(n3484) );
  NAND2_X1 U35010 ( .A1(n2718), .A2(n2200), .ZN(n2724) );
  INV_X1 U3502 ( .A(n2719), .ZN(n2722) );
  INV_X1 U35030 ( .A(n2720), .ZN(n2721) );
  NAND2_X1 U3504 ( .A1(n2722), .A2(n2721), .ZN(n3482) );
  OR2_X1 U35050 ( .A1(n2723), .A2(n3482), .ZN(n3483) );
  AND2_X1 U35060 ( .A1(n2724), .A2(n3483), .ZN(n2725) );
  NAND2_X1 U35070 ( .A1(n3805), .A2(n2891), .ZN(n2727) );
  NAND2_X1 U35080 ( .A1(n3604), .A2(n2880), .ZN(n2726) );
  NAND2_X1 U35090 ( .A1(n2727), .A2(n2726), .ZN(n3598) );
  NAND2_X1 U35100 ( .A1(n3805), .A2(n2880), .ZN(n2729) );
  NAND2_X1 U35110 ( .A1(n3604), .A2(n2674), .ZN(n2728) );
  NAND2_X1 U35120 ( .A1(n2729), .A2(n2728), .ZN(n2730) );
  XNOR2_X1 U35130 ( .A(n2730), .B(n2874), .ZN(n3599) );
  NAND2_X1 U35140 ( .A1(n4520), .A2(n2880), .ZN(n2733) );
  NAND2_X1 U35150 ( .A1(n3352), .A2(n2674), .ZN(n2732) );
  NAND2_X1 U35160 ( .A1(n2733), .A2(n2732), .ZN(n2734) );
  XNOR2_X1 U35170 ( .A(n2734), .B(n2874), .ZN(n2738) );
  NOR2_X1 U35180 ( .A1(n3233), .A2(n2710), .ZN(n2735) );
  AOI21_X1 U35190 ( .B1(n4520), .B2(n2891), .A(n2735), .ZN(n2736) );
  XNOR2_X1 U35200 ( .A(n2738), .B(n2736), .ZN(n3348) );
  INV_X1 U35210 ( .A(n2736), .ZN(n2737) );
  NAND2_X1 U35220 ( .A1(n2738), .A2(n2737), .ZN(n2739) );
  NAND2_X1 U35230 ( .A1(n2740), .A2(n2739), .ZN(n3392) );
  INV_X1 U35240 ( .A(n3392), .ZN(n2770) );
  NAND2_X1 U35250 ( .A1(n3804), .A2(n2731), .ZN(n2742) );
  NAND2_X1 U35260 ( .A1(n4517), .A2(n2674), .ZN(n2741) );
  NAND2_X1 U35270 ( .A1(n2742), .A2(n2741), .ZN(n2743) );
  XNOR2_X1 U35280 ( .A(n2743), .B(n2874), .ZN(n2763) );
  NAND2_X1 U35290 ( .A1(n3804), .A2(n2891), .ZN(n2745) );
  NAND2_X1 U35300 ( .A1(n4517), .A2(n2731), .ZN(n2744) );
  NAND2_X1 U35310 ( .A1(n2745), .A2(n2744), .ZN(n2764) );
  AND2_X1 U35320 ( .A1(n2763), .A2(n2764), .ZN(n3428) );
  NAND2_X1 U35330 ( .A1(n4494), .A2(n2880), .ZN(n2747) );
  NAND2_X1 U35340 ( .A1(n3404), .A2(n2674), .ZN(n2746) );
  NAND2_X1 U35350 ( .A1(n2747), .A2(n2746), .ZN(n2748) );
  XNOR2_X1 U35360 ( .A(n2748), .B(n2893), .ZN(n2753) );
  INV_X1 U35370 ( .A(n2753), .ZN(n2751) );
  NOR2_X1 U35380 ( .A1(n3305), .A2(n2710), .ZN(n2749) );
  AOI21_X1 U35390 ( .B1(n4494), .B2(n2891), .A(n2749), .ZN(n2752) );
  INV_X1 U35400 ( .A(n2752), .ZN(n2750) );
  NAND2_X1 U35410 ( .A1(n2751), .A2(n2750), .ZN(n2762) );
  XNOR2_X1 U35420 ( .A(n2753), .B(n2752), .ZN(n3396) );
  NAND2_X1 U35430 ( .A1(n3434), .A2(n2880), .ZN(n2755) );
  NAND2_X1 U35440 ( .A1(n3533), .A2(n2674), .ZN(n2754) );
  NAND2_X1 U35450 ( .A1(n2755), .A2(n2754), .ZN(n2756) );
  XNOR2_X1 U35460 ( .A(n2756), .B(n2874), .ZN(n2760) );
  INV_X1 U35470 ( .A(n2760), .ZN(n2758) );
  NOR2_X1 U35480 ( .A1(n3278), .A2(n2710), .ZN(n2757) );
  AOI21_X1 U35490 ( .B1(n3434), .B2(n2891), .A(n2757), .ZN(n2759) );
  NAND2_X1 U35500 ( .A1(n2758), .A2(n2759), .ZN(n2767) );
  INV_X1 U35510 ( .A(n2767), .ZN(n2761) );
  XNOR2_X1 U35520 ( .A(n2760), .B(n2759), .ZN(n3530) );
  OR2_X1 U35530 ( .A1(n2761), .A2(n3530), .ZN(n3394) );
  NAND2_X1 U35540 ( .A1(n2762), .A2(n3399), .ZN(n2769) );
  INV_X1 U35550 ( .A(n2763), .ZN(n2766) );
  INV_X1 U35560 ( .A(n2764), .ZN(n2765) );
  NAND2_X1 U35570 ( .A1(n2766), .A2(n2765), .ZN(n3528) );
  AND2_X1 U35580 ( .A1(n2767), .A2(n3528), .ZN(n3393) );
  INV_X1 U35590 ( .A(n3396), .ZN(n2768) );
  AND2_X1 U35600 ( .A1(n3393), .A2(n2768), .ZN(n3398) );
  NAND2_X1 U35610 ( .A1(n3803), .A2(n2891), .ZN(n2772) );
  NAND2_X1 U35620 ( .A1(n3579), .A2(n2880), .ZN(n2771) );
  NAND2_X1 U35630 ( .A1(n2772), .A2(n2771), .ZN(n3574) );
  NAND2_X1 U35640 ( .A1(n3803), .A2(n2731), .ZN(n2774) );
  NAND2_X1 U35650 ( .A1(n3579), .A2(n2674), .ZN(n2773) );
  NAND2_X1 U35660 ( .A1(n2774), .A2(n2773), .ZN(n2775) );
  XNOR2_X1 U35670 ( .A(n2775), .B(n2874), .ZN(n3575) );
  OAI21_X1 U35680 ( .B1(n3573), .B2(n3574), .A(n3575), .ZN(n2777) );
  NAND2_X1 U35690 ( .A1(n3573), .A2(n3574), .ZN(n2776) );
  NAND2_X1 U35700 ( .A1(n2777), .A2(n2776), .ZN(n3454) );
  NAND2_X1 U35710 ( .A1(n4496), .A2(n2880), .ZN(n2779) );
  NAND2_X1 U35720 ( .A1(n3457), .A2(n2674), .ZN(n2778) );
  NAND2_X1 U35730 ( .A1(n2779), .A2(n2778), .ZN(n2780) );
  XNOR2_X1 U35740 ( .A(n2780), .B(n2874), .ZN(n2783) );
  NAND2_X1 U35750 ( .A1(n4496), .A2(n2891), .ZN(n2782) );
  NAND2_X1 U35760 ( .A1(n3457), .A2(n2880), .ZN(n2781) );
  NAND2_X1 U35770 ( .A1(n2782), .A2(n2781), .ZN(n2784) );
  AND2_X1 U35780 ( .A1(n2783), .A2(n2784), .ZN(n3450) );
  INV_X1 U35790 ( .A(n2783), .ZN(n2786) );
  INV_X1 U35800 ( .A(n2784), .ZN(n2785) );
  NAND2_X1 U35810 ( .A1(n2786), .A2(n2785), .ZN(n3451) );
  NAND2_X1 U3582 ( .A1(n4481), .A2(n2731), .ZN(n2788) );
  NAND2_X1 U3583 ( .A1(n3558), .A2(n2674), .ZN(n2787) );
  NAND2_X1 U3584 ( .A1(n2788), .A2(n2787), .ZN(n2789) );
  XNOR2_X1 U3585 ( .A(n2789), .B(n2893), .ZN(n3369) );
  NOR2_X1 U3586 ( .A1(n4365), .A2(n2710), .ZN(n2790) );
  AOI21_X1 U3587 ( .B1(n4481), .B2(n2891), .A(n2790), .ZN(n3552) );
  NAND2_X1 U3588 ( .A1(n4316), .A2(n2880), .ZN(n2792) );
  NAND2_X1 U3589 ( .A1(n4466), .A2(n2674), .ZN(n2791) );
  NAND2_X1 U3590 ( .A1(n2792), .A2(n2791), .ZN(n2793) );
  XNOR2_X1 U3591 ( .A(n2793), .B(n2874), .ZN(n2798) );
  NAND2_X1 U3592 ( .A1(n4316), .A2(n2891), .ZN(n2795) );
  NAND2_X1 U3593 ( .A1(n4466), .A2(n2880), .ZN(n2794) );
  NAND2_X1 U3594 ( .A1(n2795), .A2(n2794), .ZN(n2799) );
  NAND2_X1 U3595 ( .A1(n2798), .A2(n2799), .ZN(n3372) );
  NAND3_X1 U3596 ( .A1(n3372), .A2(n3552), .A3(n3369), .ZN(n2802) );
  INV_X1 U3597 ( .A(n2798), .ZN(n2801) );
  INV_X1 U3598 ( .A(n2799), .ZN(n2800) );
  NAND2_X1 U3599 ( .A1(n2801), .A2(n2800), .ZN(n3371) );
  AND2_X1 U3600 ( .A1(n2802), .A2(n3371), .ZN(n2803) );
  NAND2_X1 U3601 ( .A1(n4467), .A2(n2880), .ZN(n2805) );
  NAND2_X1 U3602 ( .A1(n4458), .A2(n2674), .ZN(n2804) );
  NAND2_X1 U3603 ( .A1(n2805), .A2(n2804), .ZN(n2806) );
  XNOR2_X1 U3604 ( .A(n2806), .B(n2893), .ZN(n2808) );
  NOR2_X1 U3605 ( .A1(n4314), .A2(n2710), .ZN(n2807) );
  AOI21_X1 U3606 ( .B1(n4467), .B2(n2891), .A(n2807), .ZN(n3622) );
  NAND2_X1 U3607 ( .A1(n4459), .A2(n2880), .ZN(n2811) );
  NAND2_X1 U3608 ( .A1(n4289), .A2(n2674), .ZN(n2810) );
  NAND2_X1 U3609 ( .A1(n2811), .A2(n2810), .ZN(n2812) );
  XNOR2_X1 U3610 ( .A(n2812), .B(n2874), .ZN(n2813) );
  OAI22_X1 U3611 ( .A1(n4450), .A2(n2892), .B1(n4299), .B2(n2710), .ZN(n2814)
         );
  XOR2_X1 U3612 ( .A(n2813), .B(n2814), .Z(n3474) );
  NAND2_X1 U3613 ( .A1(n2818), .A2(n2817), .ZN(n3499) );
  NAND2_X1 U3614 ( .A1(n4296), .A2(n2731), .ZN(n2820) );
  NAND2_X1 U3615 ( .A1(n4446), .A2(n2674), .ZN(n2819) );
  NAND2_X1 U3616 ( .A1(n2820), .A2(n2819), .ZN(n2821) );
  XNOR2_X1 U3617 ( .A(n2821), .B(n2874), .ZN(n3497) );
  NAND2_X1 U3618 ( .A1(n4296), .A2(n2891), .ZN(n2823) );
  NAND2_X1 U3619 ( .A1(n4446), .A2(n2731), .ZN(n2822) );
  NAND2_X1 U3620 ( .A1(n2823), .A2(n2822), .ZN(n2824) );
  NOR2_X1 U3621 ( .A1(n3497), .A2(n2824), .ZN(n2826) );
  INV_X1 U3622 ( .A(n3497), .ZN(n2825) );
  INV_X1 U3623 ( .A(n2824), .ZN(n3496) );
  NAND2_X1 U3624 ( .A1(n4447), .A2(n2731), .ZN(n2828) );
  NAND2_X1 U3625 ( .A1(n4262), .A2(n2674), .ZN(n2827) );
  NAND2_X1 U3626 ( .A1(n2828), .A2(n2827), .ZN(n2829) );
  XNOR2_X1 U3627 ( .A(n2829), .B(n2893), .ZN(n2832) );
  NOR2_X1 U3628 ( .A1(n4259), .A2(n2710), .ZN(n2830) );
  AOI21_X1 U3629 ( .B1(n4447), .B2(n2891), .A(n2830), .ZN(n2831) );
  NOR2_X1 U3630 ( .A1(n2832), .A2(n2831), .ZN(n3586) );
  NAND2_X1 U3631 ( .A1(n2832), .A2(n2831), .ZN(n3587) );
  OAI22_X1 U3632 ( .A1(n2833), .A2(n2892), .B1(n2710), .B2(n4246), .ZN(n2838)
         );
  NAND2_X1 U3633 ( .A1(n4433), .A2(n2880), .ZN(n2835) );
  NAND2_X1 U3634 ( .A1(n3422), .A2(n2674), .ZN(n2834) );
  NAND2_X1 U3635 ( .A1(n2835), .A2(n2834), .ZN(n2836) );
  XNOR2_X1 U3636 ( .A(n2836), .B(n2874), .ZN(n2837) );
  XOR2_X1 U3637 ( .A(n2838), .B(n2837), .Z(n3419) );
  INV_X1 U3638 ( .A(n2837), .ZN(n2840) );
  INV_X1 U3639 ( .A(n2838), .ZN(n2839) );
  NAND2_X1 U3640 ( .A1(n4242), .A2(n2880), .ZN(n2842) );
  NAND2_X1 U3641 ( .A1(n3546), .A2(n2674), .ZN(n2841) );
  NAND2_X1 U3642 ( .A1(n2842), .A2(n2841), .ZN(n2843) );
  XNOR2_X1 U3643 ( .A(n2843), .B(n2893), .ZN(n2846) );
  NOR2_X1 U3644 ( .A1(n4430), .A2(n2710), .ZN(n2844) );
  AOI21_X1 U3645 ( .B1(n4242), .B2(n2891), .A(n2844), .ZN(n2845) );
  NOR2_X1 U3646 ( .A1(n2846), .A2(n2845), .ZN(n3541) );
  NAND2_X1 U3647 ( .A1(n4220), .A2(n2880), .ZN(n2848) );
  NAND2_X1 U3648 ( .A1(n4422), .A2(n2674), .ZN(n2847) );
  NAND2_X1 U3649 ( .A1(n2848), .A2(n2847), .ZN(n2849) );
  XNOR2_X1 U3650 ( .A(n2849), .B(n2893), .ZN(n3441) );
  NOR2_X1 U3651 ( .A1(n4202), .A2(n2710), .ZN(n2850) );
  AOI21_X1 U3652 ( .B1(n4220), .B2(n2891), .A(n2850), .ZN(n3440) );
  NAND2_X1 U3653 ( .A1(n3441), .A2(n3440), .ZN(n2853) );
  INV_X1 U3654 ( .A(n3441), .ZN(n2852) );
  INV_X1 U3655 ( .A(n3440), .ZN(n2851) );
  AOI22_X1 U3656 ( .A1(n3443), .A2(n2853), .B1(n2852), .B2(n2851), .ZN(n3565)
         );
  OAI22_X1 U3657 ( .A1(n4207), .A2(n2892), .B1(n4191), .B2(n2710), .ZN(n2862)
         );
  NAND2_X1 U3658 ( .A1(n4423), .A2(n2880), .ZN(n2855) );
  NAND2_X1 U3659 ( .A1(n2524), .A2(n2674), .ZN(n2854) );
  NAND2_X1 U3660 ( .A1(n2855), .A2(n2854), .ZN(n2856) );
  XNOR2_X1 U3661 ( .A(n2856), .B(n2874), .ZN(n2861) );
  XOR2_X1 U3662 ( .A(n2862), .B(n2861), .Z(n3566) );
  NAND2_X1 U3663 ( .A1(n3565), .A2(n3566), .ZN(n3564) );
  NAND2_X1 U3664 ( .A1(n4188), .A2(n2880), .ZN(n2858) );
  NAND2_X1 U3665 ( .A1(n3780), .A2(n2674), .ZN(n2857) );
  NAND2_X1 U3666 ( .A1(n2858), .A2(n2857), .ZN(n2859) );
  XNOR2_X1 U3667 ( .A(n2859), .B(n2874), .ZN(n2868) );
  NOR2_X1 U3668 ( .A1(n4168), .A2(n2710), .ZN(n2860) );
  AOI21_X1 U3669 ( .B1(n4188), .B2(n2891), .A(n2860), .ZN(n2866) );
  XNOR2_X1 U3670 ( .A(n2868), .B(n2866), .ZN(n3383) );
  INV_X1 U3671 ( .A(n2861), .ZN(n2864) );
  INV_X1 U3672 ( .A(n2862), .ZN(n2863) );
  NAND2_X1 U3673 ( .A1(n2864), .A2(n2863), .ZN(n3381) );
  NOR2_X1 U3674 ( .A1(n4147), .A2(n2710), .ZN(n2865) );
  AOI21_X1 U3675 ( .B1(n4130), .B2(n2891), .A(n2865), .ZN(n2870) );
  INV_X1 U3676 ( .A(n2866), .ZN(n2867) );
  NAND2_X1 U3677 ( .A1(n2868), .A2(n2867), .ZN(n2871) );
  NAND3_X1 U3678 ( .A1(n3382), .A2(n2870), .A3(n2871), .ZN(n3507) );
  OAI22_X1 U3679 ( .A1(n4399), .A2(n2710), .B1(n2895), .B2(n4147), .ZN(n2869)
         );
  XNOR2_X1 U3680 ( .A(n2869), .B(n2874), .ZN(n3509) );
  NAND2_X1 U3681 ( .A1(n4405), .A2(n2880), .ZN(n2873) );
  NAND2_X1 U3682 ( .A1(n4395), .A2(n2674), .ZN(n2872) );
  NAND2_X1 U3683 ( .A1(n2873), .A2(n2872), .ZN(n2875) );
  XNOR2_X1 U3684 ( .A(n2875), .B(n2874), .ZN(n2879) );
  NAND2_X1 U3685 ( .A1(n4405), .A2(n2891), .ZN(n2877) );
  NAND2_X1 U3686 ( .A1(n4395), .A2(n2880), .ZN(n2876) );
  NAND2_X1 U3687 ( .A1(n2877), .A2(n2876), .ZN(n2878) );
  NOR2_X1 U3688 ( .A1(n2879), .A2(n2878), .ZN(n3464) );
  NAND2_X1 U3689 ( .A1(n2879), .A2(n2878), .ZN(n3463) );
  NAND2_X1 U3690 ( .A1(n4396), .A2(n2880), .ZN(n2882) );
  NAND2_X1 U3691 ( .A1(n3614), .A2(n2674), .ZN(n2881) );
  NAND2_X1 U3692 ( .A1(n2882), .A2(n2881), .ZN(n2883) );
  XNOR2_X1 U3693 ( .A(n2883), .B(n2893), .ZN(n2886) );
  NOR2_X1 U3694 ( .A1(n4116), .A2(n2710), .ZN(n2884) );
  AOI21_X1 U3695 ( .B1(n4396), .B2(n2891), .A(n2884), .ZN(n2885) );
  NAND2_X1 U3696 ( .A1(n2886), .A2(n2885), .ZN(n3610) );
  NAND2_X1 U3697 ( .A1(n4110), .A2(n2880), .ZN(n2888) );
  NAND2_X1 U3698 ( .A1(n4383), .A2(n2674), .ZN(n2887) );
  NAND2_X1 U3699 ( .A1(n2888), .A2(n2887), .ZN(n2889) );
  XNOR2_X1 U3700 ( .A(n2889), .B(n2893), .ZN(n2927) );
  NOR2_X1 U3701 ( .A1(n4098), .A2(n2710), .ZN(n2890) );
  AOI21_X1 U3702 ( .B1(n4110), .B2(n2891), .A(n2890), .ZN(n2926) );
  XNOR2_X1 U3703 ( .A(n2927), .B(n2926), .ZN(n3359) );
  OAI22_X1 U3704 ( .A1(n4386), .A2(n2892), .B1(n2896), .B2(n2710), .ZN(n2894)
         );
  XNOR2_X1 U3705 ( .A(n2894), .B(n2893), .ZN(n2898) );
  OAI22_X1 U3706 ( .A1(n4386), .A2(n2710), .B1(n2896), .B2(n2895), .ZN(n2897)
         );
  XNOR2_X1 U3707 ( .A(n2898), .B(n2897), .ZN(n2931) );
  INV_X1 U3708 ( .A(n2931), .ZN(n2907) );
  NAND2_X1 U3709 ( .A1(n4611), .A2(n3082), .ZN(n2903) );
  NAND2_X1 U3710 ( .A1(n2903), .A2(n2902), .ZN(n2904) );
  OR2_X1 U3711 ( .A1(n4518), .A2(n2904), .ZN(n2909) );
  INV_X1 U3712 ( .A(n2909), .ZN(n2905) );
  NAND2_X1 U3713 ( .A1(n2907), .A2(n3624), .ZN(n2934) );
  INV_X1 U3714 ( .A(n2908), .ZN(n3339) );
  INV_X1 U3715 ( .A(n2920), .ZN(n2914) );
  NAND2_X1 U3716 ( .A1(n2909), .A2(n4500), .ZN(n2910) );
  NAND2_X1 U3717 ( .A1(n2914), .A2(n2910), .ZN(n2911) );
  NAND2_X1 U3718 ( .A1(n2911), .A2(n3093), .ZN(n3065) );
  NAND2_X1 U3719 ( .A1(n2937), .A2(n2941), .ZN(n2912) );
  OAI21_X1 U3720 ( .B1(n3065), .B2(n2912), .A(STATE_REG_SCAN_IN), .ZN(n2915)
         );
  INV_X1 U3721 ( .A(n2917), .ZN(n3793) );
  NAND2_X1 U3722 ( .A1(n2914), .A2(n3793), .ZN(n3066) );
  INV_X1 U3723 ( .A(n4617), .ZN(n3984) );
  NOR2_X1 U3724 ( .A1(n3984), .A2(n2917), .ZN(n2916) );
  NAND2_X1 U3725 ( .A1(n2920), .A2(n2916), .ZN(n3364) );
  NOR2_X1 U3726 ( .A1(n2917), .A2(n4617), .ZN(n2918) );
  AND2_X2 U3727 ( .A1(n2920), .A2(n2918), .ZN(n3627) );
  AND2_X1 U3728 ( .A1(n3090), .A2(n4518), .ZN(n2919) );
  NAND2_X1 U3729 ( .A1(n2920), .A2(n2919), .ZN(n2923) );
  NAND2_X1 U3730 ( .A1(n3090), .A2(n2921), .ZN(n2922) );
  INV_X2 U3731 ( .A(n3122), .ZN(n3628) );
  AOI22_X1 U3732 ( .A1(n4110), .A2(n3627), .B1(n3338), .B2(n3628), .ZN(n2925)
         );
  INV_X2 U3733 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X1 U3734 ( .A1(U3149), .A2(REG3_REG_28__SCAN_IN), .ZN(n2924) );
  OAI211_X1 U3735 ( .C1(n3650), .C2(n3364), .A(n2925), .B(n2924), .ZN(n2929)
         );
  OR2_X1 U3736 ( .A1(n2927), .A2(n2926), .ZN(n2930) );
  NOR3_X1 U3737 ( .A1(n2931), .A2(n3517), .A3(n2930), .ZN(n2928) );
  AOI211_X1 U3738 ( .C1(n3339), .C2(n3630), .A(n2929), .B(n2928), .ZN(n2933)
         );
  OAI211_X1 U3739 ( .C1(n2935), .C2(n2934), .A(n2933), .B(n2932), .ZN(U3217)
         );
  INV_X1 U3740 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2938) );
  XNOR2_X1 U3741 ( .A(n2997), .B(n2938), .ZN(n2945) );
  AND2_X1 U3742 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n2944)
         );
  NAND2_X1 U3743 ( .A1(n2941), .A2(n2939), .ZN(n2940) );
  NAND2_X1 U3744 ( .A1(n2310), .A2(n2940), .ZN(n2952) );
  INV_X1 U3745 ( .A(n2952), .ZN(n2943) );
  OR2_X1 U3746 ( .A1(n2941), .A2(U3149), .ZN(n3797) );
  INV_X1 U3747 ( .A(n3797), .ZN(n2942) );
  INV_X1 U3748 ( .A(n4606), .ZN(n3986) );
  NAND2_X1 U3749 ( .A1(n2945), .A2(n2944), .ZN(n2992) );
  OAI211_X1 U3750 ( .C1(n2945), .C2(n2944), .A(n4713), .B(n2992), .ZN(n2950)
         );
  NAND2_X1 U3751 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3993) );
  INV_X1 U3752 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2946) );
  MUX2_X1 U3753 ( .A(REG2_REG_1__SCAN_IN), .B(n2946), .S(n2997), .Z(n2948) );
  NOR2_X1 U3754 ( .A1(n4617), .A2(n3986), .ZN(n3794) );
  AND2_X1 U3755 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2947)
         );
  NAND2_X1 U3756 ( .A1(n2948), .A2(n2947), .ZN(n4003) );
  OAI211_X1 U3757 ( .C1(n2947), .C2(n2948), .A(n4666), .B(n4003), .ZN(n2949)
         );
  NAND2_X1 U3758 ( .A1(n2950), .A2(n2949), .ZN(n2955) );
  AND2_X1 U3759 ( .A1(n4711), .A2(ADDR_REG_1__SCAN_IN), .ZN(n2954) );
  INV_X1 U3760 ( .A(n2997), .ZN(n2957) );
  OAI22_X1 U3761 ( .A1(n4718), .A2(n2957), .B1(STATE_REG_SCAN_IN), .B2(n3129), 
        .ZN(n2953) );
  OR3_X1 U3762 ( .A1(n2955), .A2(n2954), .A3(n2953), .ZN(U3241) );
  INV_X1 U3763 ( .A(DATAI_1_), .ZN(n2956) );
  MUX2_X1 U3764 ( .A(n2957), .B(n2956), .S(U3149), .Z(n2958) );
  INV_X1 U3765 ( .A(n2958), .ZN(U3351) );
  INV_X1 U3766 ( .A(DATAI_3_), .ZN(n2959) );
  INV_X1 U3767 ( .A(n3001), .ZN(n3048) );
  MUX2_X1 U3768 ( .A(n2959), .B(n3048), .S(STATE_REG_SCAN_IN), .Z(n2960) );
  INV_X1 U3769 ( .A(n2960), .ZN(U3349) );
  INV_X1 U3770 ( .A(DATAI_7_), .ZN(n2961) );
  MUX2_X1 U3771 ( .A(n2961), .B(n2206), .S(STATE_REG_SCAN_IN), .Z(n2962) );
  INV_X1 U3772 ( .A(n2962), .ZN(U3345) );
  MUX2_X1 U3773 ( .A(n4044), .B(n2963), .S(U3149), .Z(n2964) );
  INV_X1 U3774 ( .A(n2964), .ZN(U3344) );
  MUX2_X1 U3775 ( .A(n3035), .B(n2344), .S(U3149), .Z(n2965) );
  INV_X1 U3776 ( .A(n2965), .ZN(U3347) );
  INV_X1 U3777 ( .A(DATAI_21_), .ZN(n2967) );
  NAND2_X1 U3778 ( .A1(n3786), .A2(STATE_REG_SCAN_IN), .ZN(n2966) );
  OAI21_X1 U3779 ( .B1(STATE_REG_SCAN_IN), .B2(n2967), .A(n2966), .ZN(U3331)
         );
  INV_X1 U3780 ( .A(DATAI_25_), .ZN(n2970) );
  NAND2_X1 U3781 ( .A1(n2968), .A2(STATE_REG_SCAN_IN), .ZN(n2969) );
  OAI21_X1 U3782 ( .B1(STATE_REG_SCAN_IN), .B2(n2970), .A(n2969), .ZN(U3327)
         );
  INV_X1 U3783 ( .A(DATAI_29_), .ZN(n3928) );
  NAND2_X1 U3784 ( .A1(n2971), .A2(STATE_REG_SCAN_IN), .ZN(n2972) );
  OAI21_X1 U3785 ( .B1(STATE_REG_SCAN_IN), .B2(n3928), .A(n2972), .ZN(U3323)
         );
  INV_X1 U3786 ( .A(D_REG_1__SCAN_IN), .ZN(n2976) );
  INV_X1 U3787 ( .A(n2974), .ZN(n2975) );
  AOI22_X1 U3788 ( .A1(n4749), .A2(n2976), .B1(n2975), .B2(n4750), .ZN(U3459)
         );
  INV_X1 U3789 ( .A(D_REG_0__SCAN_IN), .ZN(n2980) );
  AND2_X1 U3790 ( .A1(n2977), .A2(n4750), .ZN(n2979) );
  AOI22_X1 U3791 ( .A1(n4749), .A2(n2980), .B1(n2979), .B2(n2978), .ZN(U3458)
         );
  INV_X1 U3792 ( .A(DATAI_31_), .ZN(n2985) );
  INV_X1 U3793 ( .A(n2981), .ZN(n2983) );
  OR4_X1 U3794 ( .A1(n2983), .A2(IR_REG_30__SCAN_IN), .A3(n2982), .A4(U3149), 
        .ZN(n2984) );
  OAI21_X1 U3795 ( .B1(STATE_REG_SCAN_IN), .B2(n2985), .A(n2984), .ZN(U3321)
         );
  INV_X1 U3796 ( .A(DATAI_30_), .ZN(n2987) );
  NAND2_X1 U3797 ( .A1(n2288), .A2(STATE_REG_SCAN_IN), .ZN(n2986) );
  OAI21_X1 U3798 ( .B1(STATE_REG_SCAN_IN), .B2(n2987), .A(n2986), .ZN(U3322)
         );
  NOR2_X1 U3799 ( .A1(n4711), .A2(U4043), .ZN(U3148) );
  INV_X1 U3800 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n3947) );
  NAND2_X1 U3801 ( .A1(n2673), .A2(U4043), .ZN(n2988) );
  OAI21_X1 U3802 ( .B1(U4043), .B2(n3947), .A(n2988), .ZN(U3551) );
  INV_X1 U3803 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n3952) );
  NAND2_X1 U3804 ( .A1(n3603), .A2(U4043), .ZN(n2989) );
  OAI21_X1 U3805 ( .B1(U4043), .B2(n3952), .A(n2989), .ZN(U3555) );
  INV_X1 U3806 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4793) );
  INV_X1 U3807 ( .A(n3035), .ZN(n3004) );
  INV_X1 U3808 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2990) );
  XNOR2_X1 U3809 ( .A(n4615), .B(n2990), .ZN(n4010) );
  NAND2_X1 U3810 ( .A1(n2997), .A2(REG1_REG_1__SCAN_IN), .ZN(n2991) );
  NAND2_X1 U3811 ( .A1(n2992), .A2(n2991), .ZN(n4009) );
  INV_X1 U3812 ( .A(REG1_REG_3__SCAN_IN), .ZN(n3043) );
  INV_X1 U3813 ( .A(n2993), .ZN(n2994) );
  XOR2_X1 U3814 ( .A(n4614), .B(n2993), .Z(n4017) );
  INV_X1 U3815 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4790) );
  NOR2_X1 U3816 ( .A1(n4017), .A2(n4790), .ZN(n4016) );
  XOR2_X1 U3817 ( .A(REG1_REG_5__SCAN_IN), .B(n3035), .Z(n3029) );
  INV_X1 U3818 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2995) );
  XNOR2_X1 U3819 ( .A(n4029), .B(REG1_REG_8__SCAN_IN), .ZN(n3012) );
  INV_X1 U3820 ( .A(REG2_REG_2__SCAN_IN), .ZN(n4001) );
  INV_X1 U3821 ( .A(n4615), .ZN(n3999) );
  NAND2_X1 U3822 ( .A1(n2997), .A2(REG2_REG_1__SCAN_IN), .ZN(n4002) );
  NAND2_X1 U3823 ( .A1(n4003), .A2(n4002), .ZN(n2998) );
  NAND2_X1 U3824 ( .A1(n2999), .A2(n2998), .ZN(n4006) );
  OAI21_X1 U3825 ( .B1(n4001), .B2(n3999), .A(n4006), .ZN(n3000) );
  XOR2_X1 U3826 ( .A(n3001), .B(n3000), .Z(n3040) );
  AOI22_X1 U3827 ( .A1(n3040), .A2(REG2_REG_3__SCAN_IN), .B1(n3001), .B2(n3000), .ZN(n3002) );
  XNOR2_X1 U3828 ( .A(n3002), .B(n4614), .ZN(n4015) );
  INV_X1 U3829 ( .A(n3002), .ZN(n3003) );
  INV_X1 U3830 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3191) );
  MUX2_X1 U3831 ( .A(REG2_REG_5__SCAN_IN), .B(n3191), .S(n3035), .Z(n3032) );
  XNOR2_X1 U3832 ( .A(n3005), .B(n4613), .ZN(n3013) );
  INV_X1 U3833 ( .A(n3005), .ZN(n3006) );
  INV_X1 U3834 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3812) );
  MUX2_X1 U3835 ( .A(n3812), .B(REG2_REG_7__SCAN_IN), .S(n3058), .Z(n3054) );
  XNOR2_X1 U3836 ( .A(n4045), .B(n4044), .ZN(n4046) );
  XNOR2_X1 U3837 ( .A(REG2_REG_8__SCAN_IN), .B(n4046), .ZN(n3007) );
  NAND2_X1 U3838 ( .A1(n4666), .A2(n3007), .ZN(n3008) );
  NAND2_X1 U3839 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3432) );
  NAND2_X1 U3840 ( .A1(n3008), .A2(n3432), .ZN(n3010) );
  NOR2_X1 U3841 ( .A1(n4718), .A2(n4044), .ZN(n3009) );
  AOI211_X1 U3842 ( .C1(n4711), .C2(ADDR_REG_8__SCAN_IN), .A(n3010), .B(n3009), 
        .ZN(n3011) );
  OAI21_X1 U3843 ( .B1(n3012), .B2(n3060), .A(n3011), .ZN(U3248) );
  XNOR2_X1 U3844 ( .A(n3013), .B(REG2_REG_6__SCAN_IN), .ZN(n3021) );
  INV_X1 U3845 ( .A(n3014), .ZN(n3016) );
  OAI211_X1 U3846 ( .C1(n3016), .C2(REG1_REG_6__SCAN_IN), .A(n4713), .B(n3015), 
        .ZN(n3020) );
  AND2_X1 U3847 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3602) );
  NOR2_X1 U3848 ( .A1(n4718), .A2(n3017), .ZN(n3018) );
  AOI211_X1 U3849 ( .C1(n4711), .C2(ADDR_REG_6__SCAN_IN), .A(n3602), .B(n3018), 
        .ZN(n3019) );
  OAI211_X1 U3850 ( .C1(n3021), .C2(n4707), .A(n3020), .B(n3019), .ZN(U3246)
         );
  INV_X1 U3851 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n3023) );
  NAND2_X1 U3852 ( .A1(n4447), .A2(U4043), .ZN(n3022) );
  OAI21_X1 U3853 ( .B1(U4043), .B2(n3023), .A(n3022), .ZN(U3568) );
  INV_X1 U3854 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n3946) );
  NAND2_X1 U3855 ( .A1(n3434), .A2(U4043), .ZN(n3024) );
  OAI21_X1 U3856 ( .B1(U4043), .B2(n3946), .A(n3024), .ZN(U3559) );
  INV_X1 U3857 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n3949) );
  NAND2_X1 U3858 ( .A1(n4459), .A2(U4043), .ZN(n3025) );
  OAI21_X1 U3859 ( .B1(U4043), .B2(n3949), .A(n3025), .ZN(U3566) );
  INV_X1 U3860 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n3027) );
  NAND2_X1 U3861 ( .A1(n4520), .A2(U4043), .ZN(n3026) );
  OAI21_X1 U3862 ( .B1(U4043), .B2(n3027), .A(n3026), .ZN(U3557) );
  AOI211_X1 U3863 ( .C1(n3030), .C2(n3029), .A(n3060), .B(n3028), .ZN(n3038)
         );
  AOI211_X1 U3864 ( .C1(n3033), .C2(n3032), .A(n3031), .B(n4707), .ZN(n3037)
         );
  AND2_X1 U3865 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3488) );
  AOI21_X1 U3866 ( .B1(n4711), .B2(ADDR_REG_5__SCAN_IN), .A(n3488), .ZN(n3034)
         );
  OAI21_X1 U3867 ( .B1(n4718), .B2(n3035), .A(n3034), .ZN(n3036) );
  OR3_X1 U3868 ( .A1(n3038), .A2(n3037), .A3(n3036), .ZN(U3245) );
  INV_X1 U3869 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n3950) );
  NAND2_X1 U3870 ( .A1(n4130), .A2(U4043), .ZN(n3039) );
  OAI21_X1 U3871 ( .B1(U4043), .B2(n3950), .A(n3039), .ZN(U3574) );
  XOR2_X1 U3872 ( .A(REG2_REG_3__SCAN_IN), .B(n3040), .Z(n3045) );
  AOI211_X1 U3873 ( .C1(n3043), .C2(n3042), .A(n3041), .B(n3060), .ZN(n3044)
         );
  AOI21_X1 U3874 ( .B1(n4666), .B2(n3045), .A(n3044), .ZN(n3047) );
  INV_X1 U3875 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4730) );
  NOR2_X1 U3876 ( .A1(STATE_REG_SCAN_IN), .A2(n4730), .ZN(n3413) );
  AOI21_X1 U3877 ( .B1(n4711), .B2(ADDR_REG_3__SCAN_IN), .A(n3413), .ZN(n3046)
         );
  OAI211_X1 U3878 ( .C1(n3048), .C2(n4718), .A(n3047), .B(n3046), .ZN(U3243)
         );
  MUX2_X1 U3879 ( .A(REG1_REG_7__SCAN_IN), .B(n4793), .S(n3058), .Z(n3049) );
  XNOR2_X1 U3880 ( .A(n3050), .B(n3049), .ZN(n3061) );
  INV_X1 U3881 ( .A(n4718), .ZN(n4020) );
  NOR2_X1 U3882 ( .A1(STATE_REG_SCAN_IN), .A2(n3051), .ZN(n3351) );
  AOI21_X1 U3883 ( .B1(n4711), .B2(ADDR_REG_7__SCAN_IN), .A(n3351), .ZN(n3052)
         );
  INV_X1 U3884 ( .A(n3052), .ZN(n3057) );
  AOI211_X1 U3885 ( .C1(n3055), .C2(n3054), .A(n4707), .B(n3053), .ZN(n3056)
         );
  AOI211_X1 U3886 ( .C1(n4020), .C2(n3058), .A(n3057), .B(n3056), .ZN(n3059)
         );
  OAI21_X1 U3887 ( .B1(n3061), .B2(n3060), .A(n3059), .ZN(U3247) );
  OAI21_X1 U3888 ( .B1(n3064), .B2(n3063), .A(n3062), .ZN(n3995) );
  INV_X1 U3889 ( .A(n3065), .ZN(n3067) );
  NAND3_X1 U3890 ( .A1(n3067), .A2(n3090), .A3(n3066), .ZN(n3124) );
  OAI22_X1 U3891 ( .A1(n3122), .A2(n3112), .B1(n3068), .B2(n3364), .ZN(n3069)
         );
  AOI21_X1 U3892 ( .B1(REG3_REG_0__SCAN_IN), .B2(n3124), .A(n3069), .ZN(n3070)
         );
  OAI21_X1 U3893 ( .B1(n3995), .B2(n3517), .A(n3070), .ZN(U3229) );
  INV_X1 U3894 ( .A(n3124), .ZN(n3081) );
  OAI211_X1 U3895 ( .C1(n3073), .C2(n3072), .A(n3071), .B(n3624), .ZN(n3080)
         );
  INV_X1 U3896 ( .A(n3627), .ZN(n3075) );
  OAI22_X1 U3897 ( .A1(n3076), .A2(n3075), .B1(n3074), .B2(n3364), .ZN(n3077)
         );
  AOI21_X1 U3898 ( .B1(n3078), .B2(n3628), .A(n3077), .ZN(n3079) );
  OAI211_X1 U3899 ( .C1(n3081), .C2(n3129), .A(n3080), .B(n3079), .ZN(U3219)
         );
  INV_X1 U3900 ( .A(n3113), .ZN(n4778) );
  NAND2_X1 U3901 ( .A1(n3983), .A2(n3112), .ZN(n3678) );
  INV_X1 U3902 ( .A(n3778), .ZN(n3099) );
  INV_X1 U3903 ( .A(n3082), .ZN(n3083) );
  NOR2_X1 U3904 ( .A1(n3112), .A2(n3083), .ZN(n3089) );
  INV_X1 U3905 ( .A(n4524), .ZN(n3084) );
  NOR2_X1 U3906 ( .A1(n3084), .A2(n4529), .ZN(n3085) );
  OAI22_X1 U3907 ( .A1(n3778), .A2(n3085), .B1(n3068), .B2(n4522), .ZN(n3087)
         );
  AOI211_X1 U3908 ( .C1(n4778), .C2(n3099), .A(n3089), .B(n3087), .ZN(n4771)
         );
  NAND2_X1 U3909 ( .A1(n4792), .A2(REG1_REG_0__SCAN_IN), .ZN(n3086) );
  OAI21_X1 U3910 ( .B1(n4771), .B2(n4792), .A(n3086), .ZN(U3518) );
  AOI21_X1 U3911 ( .B1(n3089), .B2(n3088), .A(n3087), .ZN(n3102) );
  NAND2_X1 U3912 ( .A1(n3090), .A2(D_REG_1__SCAN_IN), .ZN(n3091) );
  NAND2_X1 U3913 ( .A1(n4749), .A2(n3091), .ZN(n3092) );
  NAND4_X1 U3914 ( .A1(n3095), .A2(n3094), .A3(n3093), .A4(n3092), .ZN(n3096)
         );
  AOI22_X1 U3915 ( .A1(n4744), .A2(REG2_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(n4736), .ZN(n3101) );
  OR2_X1 U3916 ( .A1(n3097), .A2(n4087), .ZN(n3170) );
  INV_X1 U3917 ( .A(n3170), .ZN(n3098) );
  NAND2_X1 U3918 ( .A1(n4722), .A2(n3098), .ZN(n4350) );
  INV_X1 U3919 ( .A(n4350), .ZN(n4739) );
  NAND2_X1 U3920 ( .A1(n3099), .A2(n4739), .ZN(n3100) );
  OAI211_X1 U3921 ( .C1(n3102), .C2(n4744), .A(n3101), .B(n3100), .ZN(U3290)
         );
  OR2_X1 U3922 ( .A1(n2582), .A2(n3103), .ZN(n3104) );
  NAND2_X1 U3923 ( .A1(n3137), .A2(n3104), .ZN(n3127) );
  NAND2_X1 U3924 ( .A1(n3983), .A2(n4519), .ZN(n3106) );
  NAND2_X1 U3925 ( .A1(n2690), .A2(n4495), .ZN(n3105) );
  OAI211_X1 U3926 ( .C1(n4500), .C2(n3111), .A(n3106), .B(n3105), .ZN(n3107)
         );
  INV_X1 U3927 ( .A(n3107), .ZN(n3110) );
  XNOR2_X1 U3928 ( .A(n2582), .B(n3676), .ZN(n3108) );
  NAND2_X1 U3929 ( .A1(n3108), .A2(n4529), .ZN(n3109) );
  OAI211_X1 U3930 ( .C1(n3127), .C2(n4524), .A(n3110), .B(n3109), .ZN(n3131)
         );
  OAI21_X1 U3931 ( .B1(n3112), .B2(n3111), .A(n3150), .ZN(n3130) );
  OAI22_X1 U3932 ( .A1(n3127), .A2(n3113), .B1(n3229), .B2(n3130), .ZN(n3114)
         );
  NOR2_X1 U3933 ( .A1(n3131), .A2(n3114), .ZN(n4773) );
  NAND2_X1 U3934 ( .A1(n4792), .A2(REG1_REG_1__SCAN_IN), .ZN(n3115) );
  OAI21_X1 U3935 ( .B1(n4773), .B2(n4792), .A(n3115), .ZN(U3519) );
  INV_X1 U3936 ( .A(n3116), .ZN(n3117) );
  AOI21_X1 U3937 ( .B1(n3119), .B2(n3118), .A(n3117), .ZN(n3126) );
  AOI22_X1 U3938 ( .A1(n3626), .A2(n3981), .B1(n3627), .B2(n2673), .ZN(n3120)
         );
  OAI21_X1 U3939 ( .B1(n3122), .B2(n3121), .A(n3120), .ZN(n3123) );
  AOI21_X1 U3940 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3124), .A(n3123), .ZN(n3125)
         );
  OAI21_X1 U3941 ( .B1(n3126), .B2(n3517), .A(n3125), .ZN(U3234) );
  INV_X1 U3942 ( .A(n3127), .ZN(n3134) );
  AND2_X1 U3943 ( .A1(n4258), .A2(n4087), .ZN(n3128) );
  OAI22_X1 U3944 ( .A1(n4371), .A2(n3130), .B1(n3129), .B2(n4719), .ZN(n3133)
         );
  MUX2_X1 U3945 ( .A(n3131), .B(REG2_REG_1__SCAN_IN), .S(n4744), .Z(n3132) );
  AOI211_X1 U3946 ( .C1(n3134), .C2(n4739), .A(n3133), .B(n3132), .ZN(n3135)
         );
  INV_X1 U3947 ( .A(n3135), .ZN(U3289) );
  NAND2_X1 U3948 ( .A1(n3137), .A2(n3136), .ZN(n3140) );
  INV_X1 U3949 ( .A(n3138), .ZN(n3139) );
  AOI21_X1 U3950 ( .B1(n3762), .B2(n3140), .A(n3139), .ZN(n3145) );
  INV_X1 U3951 ( .A(n3145), .ZN(n4740) );
  OAI21_X1 U3952 ( .B1(n3762), .B2(n3142), .A(n3141), .ZN(n3148) );
  AOI22_X1 U3953 ( .A1(n2673), .A2(n4519), .B1(n3151), .B2(n4518), .ZN(n3143)
         );
  OAI21_X1 U3954 ( .B1(n3144), .B2(n4522), .A(n3143), .ZN(n3147) );
  NOR2_X1 U3955 ( .A1(n3145), .A2(n4524), .ZN(n3146) );
  AOI211_X1 U3956 ( .C1(n4529), .C2(n3148), .A(n3147), .B(n3146), .ZN(n4743)
         );
  INV_X1 U3957 ( .A(n4743), .ZN(n3149) );
  AOI21_X1 U3958 ( .B1(n4778), .B2(n4740), .A(n3149), .ZN(n3154) );
  AOI21_X1 U3959 ( .B1(n3151), .B2(n3150), .A(n3163), .ZN(n4737) );
  INV_X1 U3960 ( .A(n4533), .ZN(n4490) );
  AOI22_X1 U3961 ( .A1(n4737), .A2(n4490), .B1(REG1_REG_2__SCAN_IN), .B2(n4792), .ZN(n3152) );
  OAI21_X1 U3962 ( .B1(n3154), .B2(n4792), .A(n3152), .ZN(U3520) );
  INV_X1 U3963 ( .A(n4605), .ZN(n4595) );
  AOI22_X1 U3964 ( .A1(n4737), .A2(n4595), .B1(REG0_REG_2__SCAN_IN), .B2(n4787), .ZN(n3153) );
  OAI21_X1 U3965 ( .B1(n3154), .B2(n4787), .A(n3153), .ZN(U3471) );
  XNOR2_X1 U3966 ( .A(n3155), .B(n3761), .ZN(n3158) );
  INV_X1 U3967 ( .A(n3158), .ZN(n4732) );
  XNOR2_X1 U3968 ( .A(n3156), .B(n3761), .ZN(n3161) );
  AOI22_X1 U3969 ( .A1(n2690), .A2(n4519), .B1(n4518), .B2(n3414), .ZN(n3157)
         );
  OAI21_X1 U3970 ( .B1(n3183), .B2(n4522), .A(n3157), .ZN(n3160) );
  NOR2_X1 U3971 ( .A1(n3158), .A2(n4524), .ZN(n3159) );
  AOI211_X1 U3972 ( .C1(n3161), .C2(n4529), .A(n3160), .B(n3159), .ZN(n4735)
         );
  INV_X1 U3973 ( .A(n4735), .ZN(n3162) );
  AOI21_X1 U3974 ( .B1(n4778), .B2(n4732), .A(n3162), .ZN(n3167) );
  INV_X1 U3975 ( .A(n3163), .ZN(n3164) );
  AOI21_X1 U3976 ( .B1(n3414), .B2(n3164), .A(n3212), .ZN(n4731) );
  AOI22_X1 U3977 ( .A1(n4731), .A2(n4490), .B1(REG1_REG_3__SCAN_IN), .B2(n4792), .ZN(n3165) );
  OAI21_X1 U3978 ( .B1(n3167), .B2(n4792), .A(n3165), .ZN(U3521) );
  AOI22_X1 U3979 ( .A1(n4731), .A2(n4595), .B1(REG0_REG_3__SCAN_IN), .B2(n4787), .ZN(n3166) );
  OAI21_X1 U3980 ( .B1(n3167), .B2(n4787), .A(n3166), .ZN(U3473) );
  NAND2_X1 U3981 ( .A1(n3691), .A2(n3699), .ZN(n3766) );
  XNOR2_X1 U3982 ( .A(n3168), .B(n3766), .ZN(n3219) );
  NAND2_X1 U3983 ( .A1(n4722), .A2(n4529), .ZN(n4230) );
  XOR2_X1 U3984 ( .A(n3766), .B(n3169), .Z(n3221) );
  NAND2_X1 U3985 ( .A1(n4524), .A2(n3170), .ZN(n3171) );
  NAND2_X1 U3986 ( .A1(n3221), .A2(n4312), .ZN(n3178) );
  INV_X1 U3987 ( .A(n3186), .ZN(n3172) );
  AOI21_X1 U3988 ( .B1(n3604), .B2(n3172), .A(n2144), .ZN(n3225) );
  INV_X1 U3989 ( .A(n4340), .ZN(n4225) );
  NAND2_X1 U3990 ( .A1(n4722), .A2(n4495), .ZN(n4344) );
  INV_X1 U3991 ( .A(n4344), .ZN(n4221) );
  AND2_X1 U3992 ( .A1(n4722), .A2(n4519), .ZN(n4339) );
  AOI22_X1 U3993 ( .A1(n4221), .A2(n4520), .B1(n4339), .B2(n3603), .ZN(n3175)
         );
  INV_X1 U3994 ( .A(n3173), .ZN(n3605) );
  AOI22_X1 U3995 ( .A1(n4744), .A2(REG2_REG_6__SCAN_IN), .B1(n3605), .B2(n4736), .ZN(n3174) );
  OAI211_X1 U3996 ( .C1(n2124), .C2(n4225), .A(n3175), .B(n3174), .ZN(n3176)
         );
  AOI21_X1 U3997 ( .B1(n3225), .B2(n4738), .A(n3176), .ZN(n3177) );
  OAI211_X1 U3998 ( .C1(n3219), .C2(n4230), .A(n3178), .B(n3177), .ZN(U3284)
         );
  NAND2_X1 U3999 ( .A1(n2082), .A2(n3698), .ZN(n3760) );
  XOR2_X1 U4000 ( .A(n3179), .B(n3760), .Z(n3199) );
  XNOR2_X1 U4001 ( .A(n3180), .B(n3760), .ZN(n3181) );
  NAND2_X1 U4002 ( .A1(n3181), .A2(n4529), .ZN(n3196) );
  AOI22_X1 U4003 ( .A1(n3805), .A2(n4495), .B1(n4518), .B2(n3489), .ZN(n3182)
         );
  OAI211_X1 U4004 ( .C1(n3183), .C2(n4484), .A(n3196), .B(n3182), .ZN(n3184)
         );
  AOI21_X1 U4005 ( .B1(n3199), .B2(n4492), .A(n3184), .ZN(n3189) );
  AND2_X1 U4006 ( .A1(n3210), .A2(n3489), .ZN(n3185) );
  NOR2_X1 U4007 ( .A1(n3186), .A2(n3185), .ZN(n3190) );
  AOI22_X1 U4008 ( .A1(n3190), .A2(n4490), .B1(REG1_REG_5__SCAN_IN), .B2(n4792), .ZN(n3187) );
  OAI21_X1 U4009 ( .B1(n3189), .B2(n4792), .A(n3187), .ZN(U3523) );
  AOI22_X1 U4010 ( .A1(n3190), .A2(n4595), .B1(REG0_REG_5__SCAN_IN), .B2(n4787), .ZN(n3188) );
  OAI21_X1 U4011 ( .B1(n3189), .B2(n4787), .A(n3188), .ZN(U3477) );
  NAND2_X1 U4012 ( .A1(n3190), .A2(n4738), .ZN(n3195) );
  OAI22_X1 U4013 ( .A1(n4722), .A2(n3191), .B1(n3490), .B2(n4719), .ZN(n3192)
         );
  AOI21_X1 U4014 ( .B1(n4221), .B2(n3805), .A(n3192), .ZN(n3194) );
  AOI22_X1 U4015 ( .A1(n4340), .A2(n3489), .B1(n4339), .B2(n3806), .ZN(n3193)
         );
  NAND3_X1 U4016 ( .A1(n3195), .A2(n3194), .A3(n3193), .ZN(n3198) );
  NOR2_X1 U4017 ( .A1(n3196), .A2(n4744), .ZN(n3197) );
  AOI211_X1 U4018 ( .C1(n3199), .C2(n4312), .A(n3198), .B(n3197), .ZN(n3200)
         );
  INV_X1 U4019 ( .A(n3200), .ZN(U3285) );
  NAND2_X1 U4020 ( .A1(n3201), .A2(n3765), .ZN(n3202) );
  NAND2_X1 U4021 ( .A1(n3203), .A2(n3202), .ZN(n4774) );
  XOR2_X1 U4022 ( .A(n3204), .B(n3765), .Z(n3209) );
  NAND2_X1 U4023 ( .A1(n3981), .A2(n4519), .ZN(n3205) );
  OAI21_X1 U4024 ( .B1(n4500), .B2(n3211), .A(n3205), .ZN(n3207) );
  NOR2_X1 U4025 ( .A1(n4774), .A2(n4524), .ZN(n3206) );
  AOI211_X1 U4026 ( .C1(n4495), .C2(n3603), .A(n3207), .B(n3206), .ZN(n3208)
         );
  OAI21_X1 U4027 ( .B1(n4505), .B2(n3209), .A(n3208), .ZN(n4776) );
  OAI211_X1 U4028 ( .C1(n3212), .C2(n3211), .A(n4258), .B(n3210), .ZN(n4775)
         );
  OAI22_X1 U4029 ( .A1(n4775), .A2(n4611), .B1(n4719), .B2(n3522), .ZN(n3213)
         );
  OAI21_X1 U4030 ( .B1(n4776), .B2(n3213), .A(n4722), .ZN(n3215) );
  NAND2_X1 U4031 ( .A1(n4744), .A2(REG2_REG_4__SCAN_IN), .ZN(n3214) );
  OAI211_X1 U4032 ( .C1(n4774), .C2(n4350), .A(n3215), .B(n3214), .ZN(U3286)
         );
  OAI22_X1 U4033 ( .A1(n3216), .A2(n4522), .B1(n4500), .B2(n2124), .ZN(n3217)
         );
  AOI21_X1 U4034 ( .B1(n4519), .B2(n3603), .A(n3217), .ZN(n3218) );
  OAI21_X1 U4035 ( .B1(n3219), .B2(n4505), .A(n3218), .ZN(n3220) );
  AOI21_X1 U4036 ( .B1(n3221), .B2(n4492), .A(n3220), .ZN(n3227) );
  AOI22_X1 U4037 ( .A1(n3225), .A2(n4490), .B1(n4792), .B2(REG1_REG_6__SCAN_IN), .ZN(n3222) );
  OAI21_X1 U4038 ( .B1(n3227), .B2(n4792), .A(n3222), .ZN(U3524) );
  INV_X1 U4039 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3223) );
  NOR2_X1 U4040 ( .A1(n4789), .A2(n3223), .ZN(n3224) );
  AOI21_X1 U4041 ( .B1(n3225), .B2(n4595), .A(n3224), .ZN(n3226) );
  OAI21_X1 U4042 ( .B1(n3227), .B2(n4787), .A(n3226), .ZN(U3479) );
  INV_X1 U40430 ( .A(n3228), .ZN(n4510) );
  AOI211_X1 U4044 ( .C1(n3352), .C2(n3230), .A(n3229), .B(n4510), .ZN(n4784)
         );
  XNOR2_X1 U4045 ( .A(n3231), .B(n3777), .ZN(n3232) );
  NAND2_X1 U4046 ( .A1(n3232), .A2(n4529), .ZN(n3236) );
  NOR2_X1 U4047 ( .A1(n3233), .A2(n4500), .ZN(n3234) );
  AOI21_X1 U4048 ( .B1(n3804), .B2(n4495), .A(n3234), .ZN(n3235) );
  OAI211_X1 U4049 ( .C1(n2125), .C2(n4484), .A(n3236), .B(n3235), .ZN(n4783)
         );
  AOI21_X1 U4050 ( .B1(n4784), .B2(n4087), .A(n4783), .ZN(n3240) );
  AND2_X1 U4051 ( .A1(n3244), .A2(n3777), .ZN(n4782) );
  NOR2_X1 U4052 ( .A1(n4782), .A2(n4375), .ZN(n3238) );
  OR2_X1 U4053 ( .A1(n3244), .A2(n3777), .ZN(n4785) );
  OAI22_X1 U4054 ( .A1(n4722), .A2(n3812), .B1(n3353), .B2(n4719), .ZN(n3237)
         );
  AOI21_X1 U4055 ( .B1(n3238), .B2(n4785), .A(n3237), .ZN(n3239) );
  OAI21_X1 U4056 ( .B1(n3240), .B2(n4744), .A(n3239), .ZN(U3283) );
  NAND2_X1 U4057 ( .A1(n2224), .A2(n3694), .ZN(n3767) );
  XNOR2_X1 U4058 ( .A(n3241), .B(n3767), .ZN(n3242) );
  NAND2_X1 U4059 ( .A1(n3242), .A2(n4529), .ZN(n3281) );
  OR2_X1 U4060 ( .A1(n3244), .A2(n3243), .ZN(n3246) );
  NAND2_X1 U4061 ( .A1(n3246), .A2(n3245), .ZN(n3247) );
  XOR2_X1 U4062 ( .A(n3767), .B(n3247), .Z(n3284) );
  NAND2_X1 U4063 ( .A1(n3284), .A2(n4312), .ZN(n3255) );
  INV_X1 U4064 ( .A(n4508), .ZN(n3249) );
  INV_X1 U4065 ( .A(n3258), .ZN(n3248) );
  OAI21_X1 U4066 ( .B1(n3249), .B2(n3278), .A(n3248), .ZN(n3290) );
  INV_X1 U4067 ( .A(n3290), .ZN(n3253) );
  INV_X1 U4068 ( .A(REG2_REG_9__SCAN_IN), .ZN(n4042) );
  OAI22_X1 U4069 ( .A1(n3534), .A2(n4719), .B1(n4042), .B2(n4722), .ZN(n3252)
         );
  AOI22_X1 U4070 ( .A1(n4221), .A2(n4494), .B1(n4339), .B2(n3804), .ZN(n3250)
         );
  OAI21_X1 U4071 ( .B1(n3278), .B2(n4225), .A(n3250), .ZN(n3251) );
  AOI211_X1 U4072 ( .C1(n3253), .C2(n4738), .A(n3252), .B(n3251), .ZN(n3254)
         );
  OAI211_X1 U4073 ( .C1(n4744), .C2(n3281), .A(n3255), .B(n3254), .ZN(U3281)
         );
  NAND2_X1 U4074 ( .A1(n3700), .A2(n3706), .ZN(n3758) );
  XNOR2_X1 U4075 ( .A(n3256), .B(n3758), .ZN(n3308) );
  XNOR2_X1 U4076 ( .A(n3257), .B(n3758), .ZN(n3310) );
  NAND2_X1 U4077 ( .A1(n3310), .A2(n4312), .ZN(n3265) );
  OAI21_X1 U4078 ( .B1(n3258), .B2(n3305), .A(n3270), .ZN(n3316) );
  INV_X1 U4079 ( .A(n3316), .ZN(n3263) );
  AOI22_X1 U4080 ( .A1(n4221), .A2(n3803), .B1(n4339), .B2(n3434), .ZN(n3261)
         );
  INV_X1 U4081 ( .A(n3259), .ZN(n3405) );
  AOI22_X1 U4082 ( .A1(n4744), .A2(REG2_REG_10__SCAN_IN), .B1(n3405), .B2(
        n4736), .ZN(n3260) );
  OAI211_X1 U4083 ( .C1(n3305), .C2(n4225), .A(n3261), .B(n3260), .ZN(n3262)
         );
  AOI21_X1 U4084 ( .B1(n3263), .B2(n4738), .A(n3262), .ZN(n3264) );
  OAI211_X1 U4085 ( .C1(n3308), .C2(n4230), .A(n3265), .B(n3264), .ZN(U3280)
         );
  INV_X1 U4086 ( .A(n3763), .ZN(n3266) );
  XNOR2_X1 U4087 ( .A(n3267), .B(n3266), .ZN(n4504) );
  OR2_X1 U4088 ( .A1(n3268), .A2(n3763), .ZN(n3296) );
  NAND2_X1 U4089 ( .A1(n3268), .A2(n3763), .ZN(n3269) );
  NAND2_X1 U4090 ( .A1(n3296), .A2(n3269), .ZN(n4493) );
  NAND2_X1 U4091 ( .A1(n3270), .A2(n3579), .ZN(n3271) );
  NAND2_X1 U4092 ( .A1(n3298), .A2(n3271), .ZN(n4601) );
  INV_X1 U4093 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3272) );
  OAI22_X1 U4094 ( .A1(n4722), .A2(n3272), .B1(n3580), .B2(n4719), .ZN(n3273)
         );
  AOI21_X1 U4095 ( .B1(n3579), .B2(n4340), .A(n3273), .ZN(n3275) );
  AOI22_X1 U4096 ( .A1(n4221), .A2(n4496), .B1(n4339), .B2(n4494), .ZN(n3274)
         );
  OAI211_X1 U4097 ( .C1(n4601), .C2(n4371), .A(n3275), .B(n3274), .ZN(n3276)
         );
  AOI21_X1 U4098 ( .B1(n4493), .B2(n4312), .A(n3276), .ZN(n3277) );
  OAI21_X1 U4099 ( .B1(n4230), .B2(n4504), .A(n3277), .ZN(U3279) );
  INV_X1 U4100 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3285) );
  NOR2_X1 U4101 ( .A1(n3278), .A2(n4500), .ZN(n3279) );
  AOI21_X1 U4102 ( .B1(n4494), .B2(n4495), .A(n3279), .ZN(n3280) );
  OAI211_X1 U4103 ( .C1(n3282), .C2(n4484), .A(n3281), .B(n3280), .ZN(n3283)
         );
  AOI21_X1 U4104 ( .B1(n3284), .B2(n4492), .A(n3283), .ZN(n3287) );
  MUX2_X1 U4105 ( .A(n3285), .B(n3287), .S(n4789), .Z(n3286) );
  OAI21_X1 U4106 ( .B1(n3290), .B2(n4605), .A(n3286), .ZN(U3485) );
  INV_X1 U4107 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3288) );
  MUX2_X1 U4108 ( .A(n3288), .B(n3287), .S(n4795), .Z(n3289) );
  OAI21_X1 U4109 ( .B1(n4533), .B2(n3290), .A(n3289), .ZN(U3527) );
  NAND2_X1 U4110 ( .A1(n3292), .A2(n3291), .ZN(n4359) );
  NAND2_X1 U4111 ( .A1(n4356), .A2(n4357), .ZN(n3759) );
  INV_X1 U4112 ( .A(n3759), .ZN(n3293) );
  XNOR2_X1 U4113 ( .A(n4359), .B(n3293), .ZN(n3294) );
  NAND2_X1 U4114 ( .A1(n3294), .A2(n4529), .ZN(n4483) );
  NAND2_X1 U4115 ( .A1(n3296), .A2(n3295), .ZN(n3297) );
  XNOR2_X1 U4116 ( .A(n3297), .B(n3759), .ZN(n4478) );
  NAND2_X1 U4117 ( .A1(n4478), .A2(n4312), .ZN(n3304) );
  AOI21_X1 U4118 ( .B1(n3457), .B2(n3298), .A(n4366), .ZN(n4596) );
  INV_X1 U4119 ( .A(n4481), .ZN(n4469) );
  AOI22_X1 U4120 ( .A1(n4340), .A2(n3457), .B1(n4339), .B2(n3803), .ZN(n3301)
         );
  INV_X1 U4121 ( .A(n3299), .ZN(n3458) );
  AOI22_X1 U4122 ( .A1(n4744), .A2(REG2_REG_12__SCAN_IN), .B1(n3458), .B2(
        n4736), .ZN(n3300) );
  OAI211_X1 U4123 ( .C1(n4469), .C2(n4344), .A(n3301), .B(n3300), .ZN(n3302)
         );
  AOI21_X1 U4124 ( .B1(n4596), .B2(n4738), .A(n3302), .ZN(n3303) );
  OAI211_X1 U4125 ( .C1(n4744), .C2(n4483), .A(n3304), .B(n3303), .ZN(U3278)
         );
  INV_X1 U4126 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3311) );
  OAI22_X1 U4127 ( .A1(n4485), .A2(n4522), .B1(n4500), .B2(n3305), .ZN(n3306)
         );
  AOI21_X1 U4128 ( .B1(n4519), .B2(n3434), .A(n3306), .ZN(n3307) );
  OAI21_X1 U4129 ( .B1(n3308), .B2(n4505), .A(n3307), .ZN(n3309) );
  AOI21_X1 U4130 ( .B1(n4492), .B2(n3310), .A(n3309), .ZN(n3313) );
  MUX2_X1 U4131 ( .A(n3311), .B(n3313), .S(n4795), .Z(n3312) );
  OAI21_X1 U4132 ( .B1(n3316), .B2(n4533), .A(n3312), .ZN(U3528) );
  INV_X1 U4133 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3314) );
  MUX2_X1 U4134 ( .A(n3314), .B(n3313), .S(n4789), .Z(n3315) );
  OAI21_X1 U4135 ( .B1(n3316), .B2(n4605), .A(n3315), .ZN(U3487) );
  NAND2_X1 U4136 ( .A1(n2051), .A2(DATAI_30_), .ZN(n3669) );
  NAND2_X1 U4137 ( .A1(n2051), .A2(DATAI_31_), .ZN(n3735) );
  XNOR2_X1 U4138 ( .A(n4376), .B(n3735), .ZN(n3328) );
  NAND2_X1 U4139 ( .A1(n2304), .A2(REG1_REG_31__SCAN_IN), .ZN(n3319) );
  NAND2_X1 U4140 ( .A1(n2330), .A2(REG2_REG_31__SCAN_IN), .ZN(n3318) );
  NAND2_X1 U4141 ( .A1(n2303), .A2(REG0_REG_31__SCAN_IN), .ZN(n3317) );
  NAND3_X1 U4142 ( .A1(n3319), .A2(n3318), .A3(n3317), .ZN(n3799) );
  NAND2_X1 U4143 ( .A1(n3799), .A2(n3320), .ZN(n4378) );
  OAI21_X1 U4144 ( .B1(n3735), .B2(n4500), .A(n4378), .ZN(n3325) );
  NAND2_X1 U4145 ( .A1(n3325), .A2(n4722), .ZN(n3322) );
  NAND2_X1 U4146 ( .A1(n4744), .A2(REG2_REG_31__SCAN_IN), .ZN(n3321) );
  OAI211_X1 U4147 ( .C1(n3328), .C2(n4371), .A(n3322), .B(n3321), .ZN(U3260)
         );
  NAND2_X1 U4148 ( .A1(n3325), .A2(n4795), .ZN(n3324) );
  NAND2_X1 U4149 ( .A1(n4792), .A2(REG1_REG_31__SCAN_IN), .ZN(n3323) );
  OAI211_X1 U4150 ( .C1(n3328), .C2(n4533), .A(n3324), .B(n3323), .ZN(U3549)
         );
  NAND2_X1 U4151 ( .A1(n3325), .A2(n4789), .ZN(n3327) );
  NAND2_X1 U4152 ( .A1(n4787), .A2(REG0_REG_31__SCAN_IN), .ZN(n3326) );
  OAI211_X1 U4153 ( .C1(n3328), .C2(n4605), .A(n3327), .B(n3326), .ZN(U3517)
         );
  NAND2_X1 U4154 ( .A1(n3329), .A2(n4312), .ZN(n3335) );
  OAI22_X1 U4155 ( .A1(n3331), .A2(n4371), .B1(n3330), .B2(n4719), .ZN(n3332)
         );
  OAI21_X1 U4156 ( .B1(n3333), .B2(n3332), .A(n4722), .ZN(n3334) );
  OAI211_X1 U4157 ( .C1(n4722), .C2(n3336), .A(n3335), .B(n3334), .ZN(U3354)
         );
  INV_X1 U4158 ( .A(n3337), .ZN(n3345) );
  AOI22_X1 U4159 ( .A1(n4110), .A2(n4339), .B1(n3338), .B2(n4340), .ZN(n3341)
         );
  AOI22_X1 U4160 ( .A1(n3339), .A2(n4736), .B1(n4744), .B2(
        REG2_REG_28__SCAN_IN), .ZN(n3340) );
  OAI211_X1 U4161 ( .C1(n3650), .C2(n4344), .A(n3341), .B(n3340), .ZN(n3344)
         );
  NOR2_X1 U4162 ( .A1(n3342), .A2(n4744), .ZN(n3343) );
  AOI211_X1 U4163 ( .C1(n4738), .C2(n3345), .A(n3344), .B(n3343), .ZN(n3346)
         );
  OAI21_X1 U4164 ( .B1(n3347), .B2(n4375), .A(n3346), .ZN(U3262) );
  XOR2_X1 U4165 ( .A(n3349), .B(n3348), .Z(n3350) );
  NAND2_X1 U4166 ( .A1(n3350), .A2(n3624), .ZN(n3358) );
  AOI21_X1 U4167 ( .B1(n3627), .B2(n3805), .A(n3351), .ZN(n3357) );
  AOI22_X1 U4168 ( .A1(n3626), .A2(n3804), .B1(n3628), .B2(n3352), .ZN(n3356)
         );
  INV_X1 U4169 ( .A(n3353), .ZN(n3354) );
  NAND2_X1 U4170 ( .A1(n3630), .A2(n3354), .ZN(n3355) );
  NAND4_X1 U4171 ( .A1(n3358), .A2(n3357), .A3(n3356), .A4(n3355), .ZN(U3210)
         );
  XNOR2_X1 U4172 ( .A(n3360), .B(n3359), .ZN(n3367) );
  INV_X1 U4173 ( .A(n3361), .ZN(n4099) );
  AOI22_X1 U4174 ( .A1(n4396), .A2(n3627), .B1(n3628), .B2(n4383), .ZN(n3363)
         );
  NAND2_X1 U4175 ( .A1(U3149), .A2(REG3_REG_27__SCAN_IN), .ZN(n3362) );
  OAI211_X1 U4176 ( .C1(n4386), .C2(n3364), .A(n3363), .B(n3362), .ZN(n3365)
         );
  AOI21_X1 U4177 ( .B1(n4099), .B2(n3630), .A(n3365), .ZN(n3366) );
  OAI21_X1 U4178 ( .B1(n3367), .B2(n3517), .A(n3366), .ZN(U3211) );
  INV_X1 U4179 ( .A(n3555), .ZN(n3368) );
  INV_X1 U4180 ( .A(n3369), .ZN(n3553) );
  NOR2_X1 U4181 ( .A1(n3368), .A2(n3553), .ZN(n3370) );
  OAI22_X1 U4182 ( .A1(n3370), .A2(n3552), .B1(n3369), .B2(n3555), .ZN(n3374)
         );
  NAND2_X1 U4183 ( .A1(n3372), .A2(n3371), .ZN(n3373) );
  XNOR2_X1 U4184 ( .A(n3374), .B(n3373), .ZN(n3375) );
  NAND2_X1 U4185 ( .A1(n3375), .A2(n3624), .ZN(n3380) );
  AND2_X1 U4186 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4039) );
  AOI21_X1 U4187 ( .B1(n3627), .B2(n4481), .A(n4039), .ZN(n3379) );
  AOI22_X1 U4188 ( .A1(n3626), .A2(n4467), .B1(n3628), .B2(n4466), .ZN(n3378)
         );
  INV_X1 U4189 ( .A(n3376), .ZN(n4341) );
  NAND2_X1 U4190 ( .A1(n3630), .A2(n4341), .ZN(n3377) );
  NAND4_X1 U4191 ( .A1(n3380), .A2(n3379), .A3(n3378), .A4(n3377), .ZN(U3212)
         );
  AND2_X1 U4192 ( .A1(n3564), .A2(n3381), .ZN(n3384) );
  OAI211_X1 U4193 ( .C1(n3384), .C2(n3383), .A(n3624), .B(n3382), .ZN(n3391)
         );
  NOR2_X1 U4194 ( .A1(n3385), .A2(STATE_REG_SCAN_IN), .ZN(n3386) );
  AOI21_X1 U4195 ( .B1(n3626), .B2(n4130), .A(n3386), .ZN(n3390) );
  AOI22_X1 U4196 ( .A1(n3780), .A2(n3628), .B1(n3627), .B2(n4423), .ZN(n3389)
         );
  INV_X1 U4197 ( .A(n3387), .ZN(n4171) );
  NAND2_X1 U4198 ( .A1(n3630), .A2(n4171), .ZN(n3388) );
  NAND4_X1 U4199 ( .A1(n3391), .A2(n3390), .A3(n3389), .A4(n3388), .ZN(U3213)
         );
  OR2_X1 U4200 ( .A1(n3392), .A2(n3428), .ZN(n3529) );
  NAND2_X1 U4201 ( .A1(n3529), .A2(n3393), .ZN(n3395) );
  AND2_X1 U4202 ( .A1(n3395), .A2(n3394), .ZN(n3397) );
  AOI21_X1 U4203 ( .B1(n3397), .B2(n3396), .A(n3517), .ZN(n3402) );
  NAND2_X1 U4204 ( .A1(n3529), .A2(n3398), .ZN(n3400) );
  AND2_X1 U4205 ( .A1(n3400), .A2(n3399), .ZN(n3401) );
  NAND2_X1 U4206 ( .A1(n3402), .A2(n3401), .ZN(n3409) );
  NAND2_X1 U4207 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4635) );
  INV_X1 U4208 ( .A(n4635), .ZN(n3403) );
  AOI21_X1 U4209 ( .B1(n3627), .B2(n3434), .A(n3403), .ZN(n3408) );
  AOI22_X1 U4210 ( .A1(n3626), .A2(n3803), .B1(n3628), .B2(n3404), .ZN(n3407)
         );
  NAND2_X1 U4211 ( .A1(n3630), .A2(n3405), .ZN(n3406) );
  NAND4_X1 U4212 ( .A1(n3409), .A2(n3408), .A3(n3407), .A4(n3406), .ZN(U3214)
         );
  XNOR2_X1 U4213 ( .A(n3411), .B(n3410), .ZN(n3412) );
  NAND2_X1 U4214 ( .A1(n3412), .A2(n3624), .ZN(n3418) );
  AOI21_X1 U4215 ( .B1(n3627), .B2(n2690), .A(n3413), .ZN(n3417) );
  AOI22_X1 U4216 ( .A1(n3626), .A2(n3806), .B1(n3628), .B2(n3414), .ZN(n3416)
         );
  NAND2_X1 U4217 ( .A1(n3630), .A2(n4730), .ZN(n3415) );
  NAND4_X1 U4218 ( .A1(n3418), .A2(n3417), .A3(n3416), .A4(n3415), .ZN(U3215)
         );
  XNOR2_X1 U4219 ( .A(n3420), .B(n3419), .ZN(n3421) );
  NAND2_X1 U4220 ( .A1(n3421), .A2(n3624), .ZN(n3427) );
  AND2_X1 U4221 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4085) );
  AOI21_X1 U4222 ( .B1(n3626), .B2(n4242), .A(n4085), .ZN(n3426) );
  AOI22_X1 U4223 ( .A1(n3422), .A2(n3628), .B1(n3627), .B2(n4447), .ZN(n3425)
         );
  INV_X1 U4224 ( .A(n4248), .ZN(n3423) );
  NAND2_X1 U4225 ( .A1(n3630), .A2(n3423), .ZN(n3424) );
  NAND4_X1 U4226 ( .A1(n3427), .A2(n3426), .A3(n3425), .A4(n3424), .ZN(U3216)
         );
  INV_X1 U4227 ( .A(n3428), .ZN(n3429) );
  NAND2_X1 U4228 ( .A1(n3429), .A2(n3528), .ZN(n3430) );
  XNOR2_X1 U4229 ( .A(n3392), .B(n3430), .ZN(n3431) );
  NAND2_X1 U4230 ( .A1(n3431), .A2(n3624), .ZN(n3439) );
  INV_X1 U4231 ( .A(n3432), .ZN(n3433) );
  AOI21_X1 U4232 ( .B1(n3627), .B2(n4520), .A(n3433), .ZN(n3438) );
  AOI22_X1 U4233 ( .A1(n3626), .A2(n3434), .B1(n3628), .B2(n4517), .ZN(n3437)
         );
  INV_X1 U4234 ( .A(n4720), .ZN(n3435) );
  NAND2_X1 U4235 ( .A1(n3630), .A2(n3435), .ZN(n3436) );
  NAND4_X1 U4236 ( .A1(n3439), .A2(n3438), .A3(n3437), .A4(n3436), .ZN(U3218)
         );
  XNOR2_X1 U4237 ( .A(n3441), .B(n3440), .ZN(n3442) );
  XNOR2_X1 U4238 ( .A(n3443), .B(n3442), .ZN(n3444) );
  NAND2_X1 U4239 ( .A1(n3444), .A2(n3624), .ZN(n3449) );
  AOI22_X1 U4240 ( .A1(n3626), .A2(n4423), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3448) );
  AOI22_X1 U4241 ( .A1(n4422), .A2(n3628), .B1(n3627), .B2(n4242), .ZN(n3447)
         );
  INV_X1 U4242 ( .A(n3445), .ZN(n4204) );
  NAND2_X1 U4243 ( .A1(n3630), .A2(n4204), .ZN(n3446) );
  NAND4_X1 U4244 ( .A1(n3449), .A2(n3448), .A3(n3447), .A4(n3446), .ZN(U3220)
         );
  INV_X1 U4245 ( .A(n3450), .ZN(n3452) );
  NAND2_X1 U4246 ( .A1(n3452), .A2(n3451), .ZN(n3453) );
  XNOR2_X1 U4247 ( .A(n3454), .B(n3453), .ZN(n3455) );
  NAND2_X1 U4248 ( .A1(n3455), .A2(n3624), .ZN(n3462) );
  NAND2_X1 U4249 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4657) );
  INV_X1 U4250 ( .A(n4657), .ZN(n3456) );
  AOI21_X1 U4251 ( .B1(n3627), .B2(n3803), .A(n3456), .ZN(n3461) );
  AOI22_X1 U4252 ( .A1(n3626), .A2(n4481), .B1(n3628), .B2(n3457), .ZN(n3460)
         );
  NAND2_X1 U4253 ( .A1(n3630), .A2(n3458), .ZN(n3459) );
  NAND4_X1 U4254 ( .A1(n3462), .A2(n3461), .A3(n3460), .A4(n3459), .ZN(U3221)
         );
  NOR2_X1 U4255 ( .A1(n3464), .A2(n2198), .ZN(n3465) );
  XNOR2_X1 U4256 ( .A(n3466), .B(n3465), .ZN(n3467) );
  NAND2_X1 U4257 ( .A1(n3467), .A2(n3624), .ZN(n3471) );
  AOI22_X1 U4258 ( .A1(n4396), .A2(n3626), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3470) );
  AOI22_X1 U4259 ( .A1(n4395), .A2(n3628), .B1(n3627), .B2(n4130), .ZN(n3469)
         );
  NAND2_X1 U4260 ( .A1(n3630), .A2(n4131), .ZN(n3468) );
  NAND4_X1 U4261 ( .A1(n3471), .A2(n3470), .A3(n3469), .A4(n3468), .ZN(U3222)
         );
  AOI21_X1 U4262 ( .B1(n3622), .B2(n3472), .A(n3620), .ZN(n3473) );
  XOR2_X1 U4263 ( .A(n3474), .B(n3473), .Z(n3475) );
  NAND2_X1 U4264 ( .A1(n3475), .A2(n3624), .ZN(n3480) );
  AND2_X1 U4265 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4692) );
  AOI21_X1 U4266 ( .B1(n3626), .B2(n4296), .A(n4692), .ZN(n3479) );
  AOI22_X1 U4267 ( .A1(n4289), .A2(n3628), .B1(n3627), .B2(n4467), .ZN(n3478)
         );
  INV_X1 U4268 ( .A(n4292), .ZN(n3476) );
  NAND2_X1 U4269 ( .A1(n3630), .A2(n3476), .ZN(n3477) );
  NAND4_X1 U4270 ( .A1(n3480), .A2(n3479), .A3(n3478), .A4(n3477), .ZN(U3223)
         );
  OR2_X1 U4271 ( .A1(n3481), .A2(n3518), .ZN(n3519) );
  NAND2_X1 U4272 ( .A1(n3519), .A2(n3482), .ZN(n3487) );
  AND2_X1 U4273 ( .A1(n3484), .A2(n3483), .ZN(n3485) );
  OAI211_X1 U4274 ( .C1(n3487), .C2(n3486), .A(n3485), .B(n3624), .ZN(n3495)
         );
  AOI21_X1 U4275 ( .B1(n3627), .B2(n3806), .A(n3488), .ZN(n3494) );
  AOI22_X1 U4276 ( .A1(n3626), .A2(n3805), .B1(n3628), .B2(n3489), .ZN(n3493)
         );
  INV_X1 U4277 ( .A(n3490), .ZN(n3491) );
  NAND2_X1 U4278 ( .A1(n3630), .A2(n3491), .ZN(n3492) );
  NAND4_X1 U4279 ( .A1(n3495), .A2(n3494), .A3(n3493), .A4(n3492), .ZN(U3224)
         );
  XNOR2_X1 U4280 ( .A(n3497), .B(n3496), .ZN(n3498) );
  XNOR2_X1 U4281 ( .A(n3499), .B(n3498), .ZN(n3500) );
  NAND2_X1 U4282 ( .A1(n3500), .A2(n3624), .ZN(n3505) );
  AND2_X1 U4283 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4701) );
  AOI21_X1 U4284 ( .B1(n3626), .B2(n4447), .A(n4701), .ZN(n3504) );
  AOI22_X1 U4285 ( .A1(n4446), .A2(n3628), .B1(n3627), .B2(n4459), .ZN(n3503)
         );
  INV_X1 U4286 ( .A(n3501), .ZN(n4278) );
  NAND2_X1 U4287 ( .A1(n3630), .A2(n4278), .ZN(n3502) );
  NAND4_X1 U4288 ( .A1(n3505), .A2(n3504), .A3(n3503), .A4(n3502), .ZN(U3225)
         );
  INV_X1 U4289 ( .A(n3506), .ZN(n3508) );
  NAND2_X1 U4290 ( .A1(n3508), .A2(n3507), .ZN(n3510) );
  XNOR2_X1 U4291 ( .A(n3510), .B(n3509), .ZN(n3511) );
  NAND2_X1 U4292 ( .A1(n3511), .A2(n3624), .ZN(n3516) );
  AOI22_X1 U4293 ( .A1(n3626), .A2(n4405), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3515) );
  AOI22_X1 U4294 ( .A1(n4404), .A2(n3628), .B1(n3627), .B2(n4188), .ZN(n3514)
         );
  INV_X1 U4295 ( .A(n3512), .ZN(n4148) );
  NAND2_X1 U4296 ( .A1(n3630), .A2(n4148), .ZN(n3513) );
  NAND4_X1 U4297 ( .A1(n3516), .A2(n3515), .A3(n3514), .A4(n3513), .ZN(U3226)
         );
  AOI21_X1 U4298 ( .B1(n3481), .B2(n3518), .A(n3517), .ZN(n3520) );
  NAND2_X1 U4299 ( .A1(n3520), .A2(n3519), .ZN(n3527) );
  AND2_X1 U4300 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n4014) );
  AOI21_X1 U4301 ( .B1(n3627), .B2(n3981), .A(n4014), .ZN(n3526) );
  AOI22_X1 U4302 ( .A1(n3626), .A2(n3603), .B1(n3628), .B2(n3521), .ZN(n3525)
         );
  INV_X1 U4303 ( .A(n3522), .ZN(n3523) );
  NAND2_X1 U4304 ( .A1(n3630), .A2(n3523), .ZN(n3524) );
  NAND4_X1 U4305 ( .A1(n3527), .A2(n3526), .A3(n3525), .A4(n3524), .ZN(U3227)
         );
  NAND2_X1 U4306 ( .A1(n3529), .A2(n3528), .ZN(n3531) );
  XNOR2_X1 U4307 ( .A(n3531), .B(n3530), .ZN(n3532) );
  NAND2_X1 U4308 ( .A1(n3532), .A2(n3624), .ZN(n3539) );
  NOR2_X1 U4309 ( .A1(STATE_REG_SCAN_IN), .A2(n3961), .ZN(n4630) );
  AOI21_X1 U4310 ( .B1(n3626), .B2(n4494), .A(n4630), .ZN(n3538) );
  AOI22_X1 U4311 ( .A1(n3533), .A2(n3628), .B1(n3627), .B2(n3804), .ZN(n3537)
         );
  INV_X1 U4312 ( .A(n3534), .ZN(n3535) );
  NAND2_X1 U4313 ( .A1(n3630), .A2(n3535), .ZN(n3536) );
  NAND4_X1 U4314 ( .A1(n3539), .A2(n3538), .A3(n3537), .A4(n3536), .ZN(U3228)
         );
  OR2_X1 U4315 ( .A1(n3540), .A2(n3541), .ZN(n3544) );
  OAI21_X1 U4316 ( .B1(n3543), .B2(n3541), .A(n3540), .ZN(n3542) );
  OAI21_X1 U4317 ( .B1(n3544), .B2(n3543), .A(n3542), .ZN(n3545) );
  NAND2_X1 U4318 ( .A1(n3545), .A2(n3624), .ZN(n3551) );
  AOI22_X1 U4319 ( .A1(n3626), .A2(n4220), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n3550) );
  AOI22_X1 U4320 ( .A1(n3546), .A2(n3628), .B1(n3627), .B2(n4433), .ZN(n3549)
         );
  INV_X1 U4321 ( .A(n3547), .ZN(n4222) );
  NAND2_X1 U4322 ( .A1(n3630), .A2(n4222), .ZN(n3548) );
  NAND4_X1 U4323 ( .A1(n3551), .A2(n3550), .A3(n3549), .A4(n3548), .ZN(U3230)
         );
  XNOR2_X1 U4324 ( .A(n3553), .B(n3552), .ZN(n3554) );
  XNOR2_X1 U4325 ( .A(n3555), .B(n3554), .ZN(n3556) );
  NAND2_X1 U4326 ( .A1(n3556), .A2(n3624), .ZN(n3563) );
  NOR2_X1 U4327 ( .A1(STATE_REG_SCAN_IN), .A2(n3557), .ZN(n4670) );
  AOI21_X1 U4328 ( .B1(n3626), .B2(n4316), .A(n4670), .ZN(n3562) );
  AOI22_X1 U4329 ( .A1(n3558), .A2(n3628), .B1(n3627), .B2(n4496), .ZN(n3561)
         );
  INV_X1 U4330 ( .A(n3559), .ZN(n4369) );
  NAND2_X1 U4331 ( .A1(n3630), .A2(n4369), .ZN(n3560) );
  NAND4_X1 U4332 ( .A1(n3563), .A2(n3562), .A3(n3561), .A4(n3560), .ZN(U3231)
         );
  OAI21_X1 U4333 ( .B1(n3566), .B2(n3565), .A(n3564), .ZN(n3567) );
  NAND2_X1 U4334 ( .A1(n3567), .A2(n3624), .ZN(n3572) );
  AOI22_X1 U4335 ( .A1(n3626), .A2(n4188), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n3571) );
  AOI22_X1 U4336 ( .A1(n2524), .A2(n3628), .B1(n3627), .B2(n4220), .ZN(n3570)
         );
  INV_X1 U4337 ( .A(n4182), .ZN(n3568) );
  NAND2_X1 U4338 ( .A1(n3630), .A2(n3568), .ZN(n3569) );
  NAND4_X1 U4339 ( .A1(n3572), .A2(n3571), .A3(n3570), .A4(n3569), .ZN(U3232)
         );
  XNOR2_X1 U4340 ( .A(n3575), .B(n3574), .ZN(n3576) );
  XNOR2_X1 U4341 ( .A(n3573), .B(n3576), .ZN(n3577) );
  NAND2_X1 U4342 ( .A1(n3577), .A2(n3624), .ZN(n3585) );
  NOR2_X1 U4343 ( .A1(STATE_REG_SCAN_IN), .A2(n3578), .ZN(n4652) );
  AOI21_X1 U4344 ( .B1(n3626), .B2(n4496), .A(n4652), .ZN(n3584) );
  AOI22_X1 U4345 ( .A1(n3579), .A2(n3628), .B1(n3627), .B2(n4494), .ZN(n3583)
         );
  INV_X1 U4346 ( .A(n3580), .ZN(n3581) );
  NAND2_X1 U4347 ( .A1(n3630), .A2(n3581), .ZN(n3582) );
  NAND4_X1 U4348 ( .A1(n3585), .A2(n3584), .A3(n3583), .A4(n3582), .ZN(U3233)
         );
  INV_X1 U4349 ( .A(n3586), .ZN(n3588) );
  NAND2_X1 U4350 ( .A1(n3588), .A2(n3587), .ZN(n3589) );
  XNOR2_X1 U4351 ( .A(n3590), .B(n3589), .ZN(n3591) );
  NAND2_X1 U4352 ( .A1(n3591), .A2(n3624), .ZN(n3596) );
  AND2_X1 U4353 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4710) );
  AOI21_X1 U4354 ( .B1(n3626), .B2(n4433), .A(n4710), .ZN(n3595) );
  AOI22_X1 U4355 ( .A1(n4262), .A2(n3628), .B1(n3627), .B2(n4296), .ZN(n3594)
         );
  INV_X1 U4356 ( .A(n3592), .ZN(n4256) );
  NAND2_X1 U4357 ( .A1(n3630), .A2(n4256), .ZN(n3593) );
  NAND4_X1 U4358 ( .A1(n3596), .A2(n3595), .A3(n3594), .A4(n3593), .ZN(U3235)
         );
  XNOR2_X1 U4359 ( .A(n3599), .B(n3598), .ZN(n3600) );
  XNOR2_X1 U4360 ( .A(n3597), .B(n3600), .ZN(n3601) );
  NAND2_X1 U4361 ( .A1(n3601), .A2(n3624), .ZN(n3609) );
  AOI21_X1 U4362 ( .B1(n3626), .B2(n4520), .A(n3602), .ZN(n3608) );
  AOI22_X1 U4363 ( .A1(n3604), .A2(n3628), .B1(n3627), .B2(n3603), .ZN(n3607)
         );
  NAND2_X1 U4364 ( .A1(n3630), .A2(n3605), .ZN(n3606) );
  NAND4_X1 U4365 ( .A1(n3609), .A2(n3608), .A3(n3607), .A4(n3606), .ZN(U3236)
         );
  NAND2_X1 U4366 ( .A1(n2077), .A2(n3610), .ZN(n3611) );
  XNOR2_X1 U4367 ( .A(n3612), .B(n3611), .ZN(n3613) );
  NAND2_X1 U4368 ( .A1(n3613), .A2(n3624), .ZN(n3619) );
  AOI22_X1 U4369 ( .A1(n4110), .A2(n3626), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3618) );
  AOI22_X1 U4370 ( .A1(n3627), .A2(n4405), .B1(n3628), .B2(n3614), .ZN(n3617)
         );
  INV_X1 U4371 ( .A(n3615), .ZN(n4117) );
  NAND2_X1 U4372 ( .A1(n3630), .A2(n4117), .ZN(n3616) );
  NAND4_X1 U4373 ( .A1(n3619), .A2(n3618), .A3(n3617), .A4(n3616), .ZN(U3237)
         );
  INV_X1 U4374 ( .A(n3472), .ZN(n3621) );
  NOR2_X1 U4375 ( .A1(n3621), .A2(n3620), .ZN(n3623) );
  XNOR2_X1 U4376 ( .A(n3623), .B(n3622), .ZN(n3625) );
  NAND2_X1 U4377 ( .A1(n3625), .A2(n3624), .ZN(n3634) );
  AND2_X1 U4378 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4682) );
  AOI21_X1 U4379 ( .B1(n3626), .B2(n4459), .A(n4682), .ZN(n3633) );
  AOI22_X1 U4380 ( .A1(n4458), .A2(n3628), .B1(n3627), .B2(n4316), .ZN(n3632)
         );
  INV_X1 U4381 ( .A(n3629), .ZN(n4317) );
  NAND2_X1 U4382 ( .A1(n3630), .A2(n4317), .ZN(n3631) );
  NAND4_X1 U4383 ( .A1(n3634), .A2(n3633), .A3(n3632), .A4(n3631), .ZN(U3238)
         );
  NAND2_X1 U4384 ( .A1(n4304), .A2(n3637), .ZN(n3711) );
  NAND2_X1 U4385 ( .A1(n3636), .A2(n3635), .ZN(n3697) );
  NAND2_X1 U4386 ( .A1(n3697), .A2(n3637), .ZN(n3710) );
  OAI21_X1 U4387 ( .B1(n4331), .B2(n3711), .A(n3710), .ZN(n3640) );
  NAND3_X1 U4388 ( .A1(n3638), .A2(n2080), .A3(n3755), .ZN(n3719) );
  AOI211_X1 U4389 ( .C1(n3640), .C2(n3715), .A(n3639), .B(n3719), .ZN(n3644)
         );
  INV_X1 U4390 ( .A(n3641), .ZN(n3643) );
  OAI21_X1 U4391 ( .B1(n3644), .B2(n3643), .A(n3642), .ZN(n3645) );
  NAND2_X1 U4392 ( .A1(n3645), .A2(n3675), .ZN(n3655) );
  NOR2_X1 U4393 ( .A1(n3744), .A2(n3646), .ZN(n3725) );
  INV_X1 U4394 ( .A(n3647), .ZN(n3745) );
  NOR2_X1 U4395 ( .A1(n3648), .A2(n3745), .ZN(n3731) );
  NAND2_X1 U4396 ( .A1(n3650), .A2(n3649), .ZN(n3662) );
  NAND4_X1 U4397 ( .A1(n3731), .A2(n3662), .A3(n3651), .A4(n3658), .ZN(n3654)
         );
  NAND2_X1 U4398 ( .A1(n3799), .A2(n3735), .ZN(n3738) );
  OR2_X1 U4399 ( .A1(n3800), .A2(n3669), .ZN(n3652) );
  AND2_X1 U4400 ( .A1(n3738), .A2(n3652), .ZN(n3776) );
  INV_X1 U4401 ( .A(n3776), .ZN(n3653) );
  AOI211_X1 U4402 ( .C1(n3655), .C2(n3725), .A(n3654), .B(n3653), .ZN(n3668)
         );
  INV_X1 U4403 ( .A(n4095), .ZN(n3666) );
  NAND2_X1 U4404 ( .A1(n3801), .A2(n3656), .ZN(n3661) );
  NAND3_X1 U4405 ( .A1(n3661), .A2(n3660), .A3(n3657), .ZN(n3728) );
  INV_X1 U4406 ( .A(n3728), .ZN(n3665) );
  NOR2_X1 U4407 ( .A1(n3659), .A2(n2252), .ZN(n3664) );
  NAND2_X1 U4408 ( .A1(n3661), .A2(n3660), .ZN(n3663) );
  OAI211_X1 U4409 ( .C1(n3664), .C2(n3663), .A(n3776), .B(n3662), .ZN(n3732)
         );
  AOI21_X1 U4410 ( .B1(n3666), .B2(n3665), .A(n3732), .ZN(n3667) );
  OAI22_X1 U4411 ( .A1(n3668), .A2(n3667), .B1(n3799), .B2(n3669), .ZN(n3674)
         );
  AND2_X1 U4412 ( .A1(n3800), .A2(n3669), .ZN(n3734) );
  INV_X1 U4413 ( .A(n3799), .ZN(n3671) );
  INV_X1 U4414 ( .A(n3735), .ZN(n3670) );
  OAI21_X1 U4415 ( .B1(n3734), .B2(n3671), .A(n3670), .ZN(n3673) );
  AOI21_X1 U4416 ( .B1(n3674), .B2(n3673), .A(n3672), .ZN(n3791) );
  INV_X1 U4417 ( .A(n3676), .ZN(n3679) );
  OAI211_X1 U4418 ( .C1(n3679), .C2(n3786), .A(n3678), .B(n3677), .ZN(n3682)
         );
  NAND3_X1 U4419 ( .A1(n3682), .A2(n3681), .A3(n3680), .ZN(n3685) );
  NAND3_X1 U4420 ( .A1(n3685), .A2(n3684), .A3(n3683), .ZN(n3688) );
  NAND3_X1 U4421 ( .A1(n3688), .A2(n3687), .A3(n3686), .ZN(n3690) );
  NAND4_X1 U4422 ( .A1(n3690), .A2(n3689), .A3(n3699), .A4(n2082), .ZN(n3693)
         );
  AND3_X1 U4423 ( .A1(n3693), .A2(n3692), .A3(n3691), .ZN(n3695) );
  NAND2_X1 U4424 ( .A1(n4513), .A2(n3774), .ZN(n3701) );
  OAI211_X1 U4425 ( .C1(n3695), .C2(n3701), .A(n3694), .B(n3775), .ZN(n3705)
         );
  NOR2_X1 U4426 ( .A1(n3697), .A2(n3696), .ZN(n3704) );
  NAND3_X1 U4427 ( .A1(n2232), .A2(n2224), .A3(n3699), .ZN(n3702) );
  OAI21_X1 U4428 ( .B1(n3702), .B2(n3701), .A(n3700), .ZN(n3703) );
  AOI22_X1 U4429 ( .A1(n3705), .A2(n3704), .B1(n3710), .B2(n3703), .ZN(n3714)
         );
  NAND3_X1 U4430 ( .A1(n3708), .A2(n3707), .A3(n3706), .ZN(n3713) );
  OAI21_X1 U4431 ( .B1(n2241), .B2(n3711), .A(n3710), .ZN(n3712) );
  OAI21_X1 U4432 ( .B1(n3714), .B2(n3713), .A(n3712), .ZN(n3718) );
  INV_X1 U4433 ( .A(n3715), .ZN(n3716) );
  AOI21_X1 U4434 ( .B1(n3718), .B2(n3717), .A(n3716), .ZN(n3720) );
  OAI21_X1 U4435 ( .B1(n3720), .B2(n3719), .A(n4157), .ZN(n3722) );
  INV_X1 U4436 ( .A(n3721), .ZN(n3764) );
  NAND2_X1 U4437 ( .A1(n3722), .A2(n3764), .ZN(n3724) );
  NAND2_X1 U4438 ( .A1(n3724), .A2(n3723), .ZN(n3726) );
  OAI221_X1 U4439 ( .B1(n2218), .B2(n3727), .C1(n2218), .C2(n3726), .A(n3725), 
        .ZN(n3730) );
  NOR2_X1 U4440 ( .A1(n2052), .A2(n4383), .ZN(n3729) );
  AOI211_X1 U4441 ( .C1(n3731), .C2(n3730), .A(n3729), .B(n3728), .ZN(n3733)
         );
  OR2_X1 U4442 ( .A1(n3733), .A2(n3732), .ZN(n3740) );
  INV_X1 U4443 ( .A(n3734), .ZN(n3737) );
  OR2_X1 U4444 ( .A1(n3799), .A2(n3735), .ZN(n3736) );
  NAND2_X1 U4445 ( .A1(n3737), .A2(n3736), .ZN(n3742) );
  NAND2_X1 U4446 ( .A1(n3742), .A2(n3738), .ZN(n3739) );
  NAND2_X1 U4447 ( .A1(n3740), .A2(n3739), .ZN(n3789) );
  NOR2_X1 U4448 ( .A1(n3741), .A2(n2065), .ZN(n4107) );
  OR3_X1 U4449 ( .A1(n3743), .A2(n4107), .A3(n3742), .ZN(n3748) );
  NOR2_X1 U4450 ( .A1(n3745), .A2(n3744), .ZN(n4125) );
  INV_X1 U4451 ( .A(n4125), .ZN(n4122) );
  NAND2_X1 U4452 ( .A1(n3747), .A2(n3746), .ZN(n4144) );
  NOR4_X1 U4453 ( .A1(n3748), .A2(n4122), .A3(n4095), .A4(n4144), .ZN(n3773)
         );
  INV_X1 U4454 ( .A(n4215), .ZN(n3749) );
  OR2_X1 U4455 ( .A1(n3749), .A2(n4214), .ZN(n4238) );
  INV_X1 U4456 ( .A(n4238), .ZN(n3757) );
  NAND2_X1 U4457 ( .A1(n3751), .A2(n3750), .ZN(n4216) );
  INV_X1 U4458 ( .A(n4216), .ZN(n3756) );
  INV_X1 U4459 ( .A(n3752), .ZN(n3754) );
  OR2_X1 U4460 ( .A1(n3754), .A2(n3753), .ZN(n4361) );
  NAND2_X1 U4461 ( .A1(n4232), .A2(n3755), .ZN(n4274) );
  NOR4_X1 U4462 ( .A1(n3757), .A2(n3756), .A3(n4361), .A4(n4274), .ZN(n3772)
         );
  NOR4_X1 U4463 ( .A1(n2582), .A2(n3760), .A3(n3759), .A4(n3758), .ZN(n3771)
         );
  NAND4_X1 U4464 ( .A1(n2098), .A2(n3763), .A3(n3762), .A4(n3761), .ZN(n3769)
         );
  NAND2_X1 U4465 ( .A1(n4199), .A2(n3765), .ZN(n3768) );
  NOR4_X1 U4466 ( .A1(n3769), .A2(n3768), .A3(n3767), .A4(n3766), .ZN(n3770)
         );
  NAND4_X1 U4467 ( .A1(n3773), .A2(n3772), .A3(n3771), .A4(n3770), .ZN(n3785)
         );
  INV_X1 U4468 ( .A(n4310), .ZN(n4305) );
  NAND4_X1 U4469 ( .A1(n2450), .A2(n4305), .A3(n4294), .A4(n4515), .ZN(n3784)
         );
  NAND4_X1 U4470 ( .A1(n4176), .A2(n3778), .A3(n3777), .A4(n3776), .ZN(n3783)
         );
  INV_X1 U4471 ( .A(n3779), .ZN(n3781) );
  XNOR2_X1 U4472 ( .A(n4188), .B(n3780), .ZN(n4162) );
  NAND2_X1 U4473 ( .A1(n3781), .A2(n4162), .ZN(n3782) );
  NOR4_X1 U4474 ( .A1(n3785), .A2(n3784), .A3(n3783), .A4(n3782), .ZN(n3787)
         );
  NOR2_X1 U4475 ( .A1(n3787), .A2(n3786), .ZN(n3788) );
  MUX2_X1 U4476 ( .A(n3789), .B(n3788), .S(n4610), .Z(n3790) );
  NOR2_X1 U4477 ( .A1(n3791), .A2(n3790), .ZN(n3792) );
  XNOR2_X1 U4478 ( .A(n3792), .B(n4611), .ZN(n3798) );
  NAND2_X1 U4479 ( .A1(n3794), .A2(n3793), .ZN(n3795) );
  OAI211_X1 U4480 ( .C1(n4609), .C2(n3797), .A(n3795), .B(B_REG_SCAN_IN), .ZN(
        n3796) );
  OAI21_X1 U4481 ( .B1(n3798), .B2(n3797), .A(n3796), .ZN(U3239) );
  MUX2_X1 U4482 ( .A(n3799), .B(DATAO_REG_31__SCAN_IN), .S(n3982), .Z(U3581)
         );
  MUX2_X1 U4483 ( .A(n3800), .B(DATAO_REG_30__SCAN_IN), .S(n3982), .Z(U3580)
         );
  MUX2_X1 U4484 ( .A(n3801), .B(DATAO_REG_29__SCAN_IN), .S(n3982), .Z(U3579)
         );
  MUX2_X1 U4485 ( .A(DATAO_REG_28__SCAN_IN), .B(n3802), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4486 ( .A(n4110), .B(DATAO_REG_27__SCAN_IN), .S(n3982), .Z(U3577)
         );
  MUX2_X1 U4487 ( .A(n4396), .B(DATAO_REG_26__SCAN_IN), .S(n3982), .Z(U3576)
         );
  MUX2_X1 U4488 ( .A(n4405), .B(DATAO_REG_25__SCAN_IN), .S(n3982), .Z(U3575)
         );
  MUX2_X1 U4489 ( .A(n4188), .B(DATAO_REG_23__SCAN_IN), .S(n3982), .Z(U3573)
         );
  MUX2_X1 U4490 ( .A(n4423), .B(DATAO_REG_22__SCAN_IN), .S(n3982), .Z(U3572)
         );
  MUX2_X1 U4491 ( .A(n4220), .B(DATAO_REG_21__SCAN_IN), .S(n3982), .Z(U3571)
         );
  MUX2_X1 U4492 ( .A(n4242), .B(DATAO_REG_20__SCAN_IN), .S(n3982), .Z(U3570)
         );
  MUX2_X1 U4493 ( .A(n4433), .B(DATAO_REG_19__SCAN_IN), .S(n3982), .Z(U3569)
         );
  MUX2_X1 U4494 ( .A(n4296), .B(DATAO_REG_17__SCAN_IN), .S(n3982), .Z(U3567)
         );
  MUX2_X1 U4495 ( .A(n4467), .B(DATAO_REG_15__SCAN_IN), .S(n3982), .Z(U3565)
         );
  MUX2_X1 U4496 ( .A(n4316), .B(DATAO_REG_14__SCAN_IN), .S(n3982), .Z(U3564)
         );
  MUX2_X1 U4497 ( .A(n4481), .B(DATAO_REG_13__SCAN_IN), .S(n3982), .Z(U3563)
         );
  MUX2_X1 U4498 ( .A(n4496), .B(DATAO_REG_12__SCAN_IN), .S(n3982), .Z(U3562)
         );
  MUX2_X1 U4499 ( .A(n3803), .B(DATAO_REG_11__SCAN_IN), .S(n3982), .Z(U3561)
         );
  MUX2_X1 U4500 ( .A(n4494), .B(DATAO_REG_10__SCAN_IN), .S(n3982), .Z(U3560)
         );
  MUX2_X1 U4501 ( .A(n3804), .B(DATAO_REG_8__SCAN_IN), .S(n3982), .Z(U3558) );
  MUX2_X1 U4502 ( .A(n3805), .B(DATAO_REG_6__SCAN_IN), .S(n3982), .Z(U3556) );
  MUX2_X1 U4503 ( .A(n3806), .B(DATAO_REG_4__SCAN_IN), .S(n3982), .Z(n3980) );
  INV_X1 U4504 ( .A(ADDR_REG_10__SCAN_IN), .ZN(n3926) );
  OAI22_X1 U4505 ( .A1(n4730), .A2(keyinput118), .B1(n3926), .B2(keyinput121), 
        .ZN(n3807) );
  AOI221_X1 U4506 ( .B1(n4730), .B2(keyinput118), .C1(keyinput121), .C2(n3926), 
        .A(n3807), .ZN(n3816) );
  INV_X1 U4507 ( .A(ADDR_REG_1__SCAN_IN), .ZN(n3809) );
  OAI22_X1 U4508 ( .A1(n3809), .A2(keyinput80), .B1(IR_REG_18__SCAN_IN), .B2(
        keyinput87), .ZN(n3808) );
  AOI221_X1 U4509 ( .B1(n3809), .B2(keyinput80), .C1(keyinput87), .C2(
        IR_REG_18__SCAN_IN), .A(n3808), .ZN(n3815) );
  INV_X1 U4510 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4025) );
  OAI22_X1 U4511 ( .A1(n4025), .A2(keyinput120), .B1(n3288), .B2(keyinput127), 
        .ZN(n3810) );
  AOI221_X1 U4512 ( .B1(n4025), .B2(keyinput120), .C1(keyinput127), .C2(n3288), 
        .A(n3810), .ZN(n3814) );
  INV_X1 U4513 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3925) );
  OAI22_X1 U4514 ( .A1(n3925), .A2(keyinput124), .B1(n3812), .B2(keyinput104), 
        .ZN(n3811) );
  AOI221_X1 U4515 ( .B1(n3925), .B2(keyinput124), .C1(keyinput104), .C2(n3812), 
        .A(n3811), .ZN(n3813) );
  NAND4_X1 U4516 ( .A1(n3816), .A2(n3815), .A3(n3814), .A4(n3813), .ZN(n3851)
         );
  OAI22_X1 U4517 ( .A1(IR_REG_23__SCAN_IN), .A2(keyinput116), .B1(keyinput70), 
        .B2(DATAO_REG_4__SCAN_IN), .ZN(n3817) );
  AOI221_X1 U4518 ( .B1(IR_REG_23__SCAN_IN), .B2(keyinput116), .C1(
        DATAO_REG_4__SCAN_IN), .C2(keyinput70), .A(n3817), .ZN(n3824) );
  OAI22_X1 U4519 ( .A1(REG0_REG_29__SCAN_IN), .A2(keyinput103), .B1(
        REG3_REG_6__SCAN_IN), .B2(keyinput119), .ZN(n3818) );
  AOI221_X1 U4520 ( .B1(REG0_REG_29__SCAN_IN), .B2(keyinput103), .C1(
        keyinput119), .C2(REG3_REG_6__SCAN_IN), .A(n3818), .ZN(n3823) );
  OAI22_X1 U4521 ( .A1(DATAO_REG_1__SCAN_IN), .A2(keyinput113), .B1(
        DATAO_REG_9__SCAN_IN), .B2(keyinput85), .ZN(n3819) );
  AOI221_X1 U4522 ( .B1(DATAO_REG_1__SCAN_IN), .B2(keyinput113), .C1(
        keyinput85), .C2(DATAO_REG_9__SCAN_IN), .A(n3819), .ZN(n3822) );
  OAI22_X1 U4523 ( .A1(DATAO_REG_24__SCAN_IN), .A2(keyinput123), .B1(
        DATAO_REG_16__SCAN_IN), .B2(keyinput84), .ZN(n3820) );
  AOI221_X1 U4524 ( .B1(DATAO_REG_24__SCAN_IN), .B2(keyinput123), .C1(
        keyinput84), .C2(DATAO_REG_16__SCAN_IN), .A(n3820), .ZN(n3821) );
  NAND4_X1 U4525 ( .A1(n3824), .A2(n3823), .A3(n3822), .A4(n3821), .ZN(n3850)
         );
  INV_X1 U4526 ( .A(DATAI_19_), .ZN(n3826) );
  AOI22_X1 U4527 ( .A1(n3826), .A2(keyinput66), .B1(keyinput93), .B2(n3952), 
        .ZN(n3825) );
  OAI221_X1 U4528 ( .B1(n3826), .B2(keyinput66), .C1(n3952), .C2(keyinput93), 
        .A(n3825), .ZN(n3837) );
  INV_X1 U4529 ( .A(ADDR_REG_18__SCAN_IN), .ZN(n3829) );
  INV_X1 U4530 ( .A(ADDR_REG_6__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4531 ( .A1(n3829), .A2(keyinput81), .B1(keyinput126), .B2(n3828), 
        .ZN(n3827) );
  OAI221_X1 U4532 ( .B1(n3829), .B2(keyinput81), .C1(n3828), .C2(keyinput126), 
        .A(n3827), .ZN(n3836) );
  INV_X1 U4533 ( .A(REG1_REG_31__SCAN_IN), .ZN(n3830) );
  XOR2_X1 U4534 ( .A(n3830), .B(keyinput105), .Z(n3834) );
  XNOR2_X1 U4535 ( .A(IR_REG_8__SCAN_IN), .B(keyinput92), .ZN(n3833) );
  XNOR2_X1 U4536 ( .A(IR_REG_12__SCAN_IN), .B(keyinput111), .ZN(n3832) );
  XNOR2_X1 U4537 ( .A(IR_REG_25__SCAN_IN), .B(keyinput65), .ZN(n3831) );
  NAND4_X1 U4538 ( .A1(n3834), .A2(n3833), .A3(n3832), .A4(n3831), .ZN(n3835)
         );
  OR3_X1 U4539 ( .A1(n3837), .A2(n3836), .A3(n3835), .ZN(n3849) );
  INV_X1 U4540 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3839) );
  INV_X1 U4541 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4788) );
  OAI22_X1 U4542 ( .A1(n3839), .A2(keyinput71), .B1(n4788), .B2(keyinput91), 
        .ZN(n3838) );
  AOI221_X1 U4543 ( .B1(n3839), .B2(keyinput71), .C1(keyinput91), .C2(n4788), 
        .A(n3838), .ZN(n3847) );
  INV_X1 U4544 ( .A(D_REG_25__SCAN_IN), .ZN(n4746) );
  INV_X1 U4545 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4542) );
  OAI22_X1 U4546 ( .A1(n4746), .A2(keyinput122), .B1(n4542), .B2(keyinput73), 
        .ZN(n3840) );
  AOI221_X1 U4547 ( .B1(n4746), .B2(keyinput122), .C1(keyinput73), .C2(n4542), 
        .A(n3840), .ZN(n3846) );
  XNOR2_X1 U4548 ( .A(IR_REG_11__SCAN_IN), .B(keyinput86), .ZN(n3844) );
  XNOR2_X1 U4549 ( .A(REG1_REG_12__SCAN_IN), .B(keyinput109), .ZN(n3843) );
  XNOR2_X1 U4550 ( .A(IR_REG_28__SCAN_IN), .B(keyinput75), .ZN(n3842) );
  XNOR2_X1 U4551 ( .A(keyinput107), .B(REG1_REG_29__SCAN_IN), .ZN(n3841) );
  AND4_X1 U4552 ( .A1(n3844), .A2(n3843), .A3(n3842), .A4(n3841), .ZN(n3845)
         );
  NAND3_X1 U4553 ( .A1(n3847), .A2(n3846), .A3(n3845), .ZN(n3848) );
  NOR4_X1 U4554 ( .A1(n3851), .A2(n3850), .A3(n3849), .A4(n3848), .ZN(n3978)
         );
  OAI22_X1 U4555 ( .A1(REG0_REG_27__SCAN_IN), .A2(keyinput96), .B1(
        REG3_REG_1__SCAN_IN), .B2(keyinput94), .ZN(n3852) );
  AOI221_X1 U4556 ( .B1(REG0_REG_27__SCAN_IN), .B2(keyinput96), .C1(keyinput94), .C2(REG3_REG_1__SCAN_IN), .A(n3852), .ZN(n3859) );
  OAI22_X1 U4557 ( .A1(DATAI_29_), .A2(keyinput67), .B1(keyinput72), .B2(
        REG1_REG_20__SCAN_IN), .ZN(n3853) );
  AOI221_X1 U4558 ( .B1(DATAI_29_), .B2(keyinput67), .C1(REG1_REG_20__SCAN_IN), 
        .C2(keyinput72), .A(n3853), .ZN(n3858) );
  OAI22_X1 U4559 ( .A1(REG3_REG_5__SCAN_IN), .A2(keyinput74), .B1(keyinput77), 
        .B2(ADDR_REG_5__SCAN_IN), .ZN(n3854) );
  AOI221_X1 U4560 ( .B1(REG3_REG_5__SCAN_IN), .B2(keyinput74), .C1(
        ADDR_REG_5__SCAN_IN), .C2(keyinput77), .A(n3854), .ZN(n3857) );
  OAI22_X1 U4561 ( .A1(IR_REG_0__SCAN_IN), .A2(keyinput83), .B1(keyinput112), 
        .B2(REG3_REG_11__SCAN_IN), .ZN(n3855) );
  AOI221_X1 U4562 ( .B1(IR_REG_0__SCAN_IN), .B2(keyinput83), .C1(
        REG3_REG_11__SCAN_IN), .C2(keyinput112), .A(n3855), .ZN(n3856) );
  NAND4_X1 U4563 ( .A1(n3859), .A2(n3858), .A3(n3857), .A4(n3856), .ZN(n3887)
         );
  OAI22_X1 U4564 ( .A1(DATAI_1_), .A2(keyinput69), .B1(DATAI_24_), .B2(
        keyinput88), .ZN(n3860) );
  AOI221_X1 U4565 ( .B1(DATAI_1_), .B2(keyinput69), .C1(keyinput88), .C2(
        DATAI_24_), .A(n3860), .ZN(n3867) );
  OAI22_X1 U4566 ( .A1(REG2_REG_25__SCAN_IN), .A2(keyinput106), .B1(
        REG2_REG_17__SCAN_IN), .B2(keyinput95), .ZN(n3861) );
  AOI221_X1 U4567 ( .B1(REG2_REG_25__SCAN_IN), .B2(keyinput106), .C1(
        keyinput95), .C2(REG2_REG_17__SCAN_IN), .A(n3861), .ZN(n3866) );
  OAI22_X1 U4568 ( .A1(REG3_REG_22__SCAN_IN), .A2(keyinput99), .B1(
        REG2_REG_26__SCAN_IN), .B2(keyinput98), .ZN(n3862) );
  AOI221_X1 U4569 ( .B1(REG3_REG_22__SCAN_IN), .B2(keyinput99), .C1(keyinput98), .C2(REG2_REG_26__SCAN_IN), .A(n3862), .ZN(n3865) );
  OAI22_X1 U4570 ( .A1(DATAI_20_), .A2(keyinput115), .B1(keyinput90), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n3863) );
  AOI221_X1 U4571 ( .B1(DATAI_20_), .B2(keyinput115), .C1(DATAO_REG_7__SCAN_IN), .C2(keyinput90), .A(n3863), .ZN(n3864) );
  NAND4_X1 U4572 ( .A1(n3867), .A2(n3866), .A3(n3865), .A4(n3864), .ZN(n3886)
         );
  OAI22_X1 U4573 ( .A1(D_REG_31__SCAN_IN), .A2(keyinput64), .B1(keyinput76), 
        .B2(REG3_REG_9__SCAN_IN), .ZN(n3868) );
  AOI221_X1 U4574 ( .B1(D_REG_31__SCAN_IN), .B2(keyinput64), .C1(
        REG3_REG_9__SCAN_IN), .C2(keyinput76), .A(n3868), .ZN(n3875) );
  OAI22_X1 U4575 ( .A1(REG1_REG_10__SCAN_IN), .A2(keyinput89), .B1(keyinput79), 
        .B2(REG1_REG_8__SCAN_IN), .ZN(n3869) );
  AOI221_X1 U4576 ( .B1(REG1_REG_10__SCAN_IN), .B2(keyinput89), .C1(
        REG1_REG_8__SCAN_IN), .C2(keyinput79), .A(n3869), .ZN(n3874) );
  OAI22_X1 U4577 ( .A1(REG1_REG_21__SCAN_IN), .A2(keyinput114), .B1(
        keyinput108), .B2(DATAO_REG_18__SCAN_IN), .ZN(n3870) );
  AOI221_X1 U4578 ( .B1(REG1_REG_21__SCAN_IN), .B2(keyinput114), .C1(
        DATAO_REG_18__SCAN_IN), .C2(keyinput108), .A(n3870), .ZN(n3873) );
  OAI22_X1 U4579 ( .A1(D_REG_3__SCAN_IN), .A2(keyinput110), .B1(
        REG1_REG_16__SCAN_IN), .B2(keyinput97), .ZN(n3871) );
  AOI221_X1 U4580 ( .B1(D_REG_3__SCAN_IN), .B2(keyinput110), .C1(keyinput97), 
        .C2(REG1_REG_16__SCAN_IN), .A(n3871), .ZN(n3872) );
  NAND4_X1 U4581 ( .A1(n3875), .A2(n3874), .A3(n3873), .A4(n3872), .ZN(n3885)
         );
  OAI22_X1 U4582 ( .A1(D_REG_27__SCAN_IN), .A2(keyinput78), .B1(keyinput125), 
        .B2(REG1_REG_1__SCAN_IN), .ZN(n3876) );
  AOI221_X1 U4583 ( .B1(D_REG_27__SCAN_IN), .B2(keyinput78), .C1(
        REG1_REG_1__SCAN_IN), .C2(keyinput125), .A(n3876), .ZN(n3883) );
  OAI22_X1 U4584 ( .A1(REG1_REG_11__SCAN_IN), .A2(keyinput68), .B1(keyinput101), .B2(ADDR_REG_11__SCAN_IN), .ZN(n3877) );
  AOI221_X1 U4585 ( .B1(REG1_REG_11__SCAN_IN), .B2(keyinput68), .C1(
        ADDR_REG_11__SCAN_IN), .C2(keyinput101), .A(n3877), .ZN(n3882) );
  OAI22_X1 U4586 ( .A1(IR_REG_31__SCAN_IN), .A2(keyinput117), .B1(
        REG0_REG_12__SCAN_IN), .B2(keyinput82), .ZN(n3878) );
  AOI221_X1 U4587 ( .B1(IR_REG_31__SCAN_IN), .B2(keyinput117), .C1(keyinput82), 
        .C2(REG0_REG_12__SCAN_IN), .A(n3878), .ZN(n3881) );
  OAI22_X1 U4588 ( .A1(D_REG_9__SCAN_IN), .A2(keyinput102), .B1(keyinput100), 
        .B2(D_REG_14__SCAN_IN), .ZN(n3879) );
  AOI221_X1 U4589 ( .B1(D_REG_9__SCAN_IN), .B2(keyinput102), .C1(
        D_REG_14__SCAN_IN), .C2(keyinput100), .A(n3879), .ZN(n3880) );
  NAND4_X1 U4590 ( .A1(n3883), .A2(n3882), .A3(n3881), .A4(n3880), .ZN(n3884)
         );
  NOR4_X1 U4591 ( .A1(n3887), .A2(n3886), .A3(n3885), .A4(n3884), .ZN(n3977)
         );
  AOI22_X1 U4592 ( .A1(REG2_REG_26__SCAN_IN), .A2(keyinput34), .B1(
        REG3_REG_3__SCAN_IN), .B2(keyinput54), .ZN(n3888) );
  OAI221_X1 U4593 ( .B1(REG2_REG_26__SCAN_IN), .B2(keyinput34), .C1(
        REG3_REG_3__SCAN_IN), .C2(keyinput54), .A(n3888), .ZN(n3895) );
  AOI22_X1 U4594 ( .A1(DATAO_REG_7__SCAN_IN), .A2(keyinput26), .B1(
        REG2_REG_25__SCAN_IN), .B2(keyinput42), .ZN(n3889) );
  OAI221_X1 U4595 ( .B1(DATAO_REG_7__SCAN_IN), .B2(keyinput26), .C1(
        REG2_REG_25__SCAN_IN), .C2(keyinput42), .A(n3889), .ZN(n3894) );
  AOI22_X1 U4596 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput30), .B1(
        REG3_REG_5__SCAN_IN), .B2(keyinput10), .ZN(n3890) );
  OAI221_X1 U4597 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput30), .C1(
        REG3_REG_5__SCAN_IN), .C2(keyinput10), .A(n3890), .ZN(n3893) );
  AOI22_X1 U4598 ( .A1(D_REG_9__SCAN_IN), .A2(keyinput38), .B1(
        D_REG_27__SCAN_IN), .B2(keyinput14), .ZN(n3891) );
  OAI221_X1 U4599 ( .B1(D_REG_9__SCAN_IN), .B2(keyinput38), .C1(
        D_REG_27__SCAN_IN), .C2(keyinput14), .A(n3891), .ZN(n3892) );
  NOR4_X1 U4600 ( .A1(n3895), .A2(n3894), .A3(n3893), .A4(n3892), .ZN(n3923)
         );
  AOI22_X1 U4601 ( .A1(REG0_REG_12__SCAN_IN), .A2(keyinput18), .B1(
        IR_REG_11__SCAN_IN), .B2(keyinput22), .ZN(n3896) );
  OAI221_X1 U4602 ( .B1(REG0_REG_12__SCAN_IN), .B2(keyinput18), .C1(
        IR_REG_11__SCAN_IN), .C2(keyinput22), .A(n3896), .ZN(n3903) );
  AOI22_X1 U4603 ( .A1(ADDR_REG_6__SCAN_IN), .A2(keyinput62), .B1(DATAI_1_), 
        .B2(keyinput5), .ZN(n3897) );
  OAI221_X1 U4604 ( .B1(ADDR_REG_6__SCAN_IN), .B2(keyinput62), .C1(DATAI_1_), 
        .C2(keyinput5), .A(n3897), .ZN(n3902) );
  AOI22_X1 U4605 ( .A1(DATAI_24_), .A2(keyinput24), .B1(DATAI_20_), .B2(
        keyinput51), .ZN(n3898) );
  OAI221_X1 U4606 ( .B1(DATAI_24_), .B2(keyinput24), .C1(DATAI_20_), .C2(
        keyinput51), .A(n3898), .ZN(n3901) );
  AOI22_X1 U4607 ( .A1(REG1_REG_20__SCAN_IN), .A2(keyinput8), .B1(
        REG3_REG_22__SCAN_IN), .B2(keyinput35), .ZN(n3899) );
  OAI221_X1 U4608 ( .B1(REG1_REG_20__SCAN_IN), .B2(keyinput8), .C1(
        REG3_REG_22__SCAN_IN), .C2(keyinput35), .A(n3899), .ZN(n3900) );
  NOR4_X1 U4609 ( .A1(n3903), .A2(n3902), .A3(n3901), .A4(n3900), .ZN(n3922)
         );
  AOI22_X1 U4610 ( .A1(REG0_REG_27__SCAN_IN), .A2(keyinput32), .B1(
        REG3_REG_11__SCAN_IN), .B2(keyinput48), .ZN(n3904) );
  OAI221_X1 U4611 ( .B1(REG0_REG_27__SCAN_IN), .B2(keyinput32), .C1(
        REG3_REG_11__SCAN_IN), .C2(keyinput48), .A(n3904), .ZN(n3911) );
  AOI22_X1 U4612 ( .A1(ADDR_REG_1__SCAN_IN), .A2(keyinput16), .B1(
        IR_REG_0__SCAN_IN), .B2(keyinput19), .ZN(n3905) );
  OAI221_X1 U4613 ( .B1(ADDR_REG_1__SCAN_IN), .B2(keyinput16), .C1(
        IR_REG_0__SCAN_IN), .C2(keyinput19), .A(n3905), .ZN(n3910) );
  AOI22_X1 U4614 ( .A1(ADDR_REG_5__SCAN_IN), .A2(keyinput13), .B1(
        ADDR_REG_11__SCAN_IN), .B2(keyinput37), .ZN(n3906) );
  OAI221_X1 U4615 ( .B1(ADDR_REG_5__SCAN_IN), .B2(keyinput13), .C1(
        ADDR_REG_11__SCAN_IN), .C2(keyinput37), .A(n3906), .ZN(n3909) );
  AOI22_X1 U4616 ( .A1(REG2_REG_7__SCAN_IN), .A2(keyinput40), .B1(
        REG1_REG_13__SCAN_IN), .B2(keyinput56), .ZN(n3907) );
  OAI221_X1 U4617 ( .B1(REG2_REG_7__SCAN_IN), .B2(keyinput40), .C1(
        REG1_REG_13__SCAN_IN), .C2(keyinput56), .A(n3907), .ZN(n3908) );
  NOR4_X1 U4618 ( .A1(n3911), .A2(n3910), .A3(n3909), .A4(n3908), .ZN(n3921)
         );
  AOI22_X1 U4619 ( .A1(REG1_REG_9__SCAN_IN), .A2(keyinput63), .B1(
        REG1_REG_11__SCAN_IN), .B2(keyinput4), .ZN(n3912) );
  OAI221_X1 U4620 ( .B1(REG1_REG_9__SCAN_IN), .B2(keyinput63), .C1(
        REG1_REG_11__SCAN_IN), .C2(keyinput4), .A(n3912), .ZN(n3919) );
  AOI22_X1 U4621 ( .A1(REG1_REG_8__SCAN_IN), .A2(keyinput15), .B1(
        D_REG_14__SCAN_IN), .B2(keyinput36), .ZN(n3913) );
  OAI221_X1 U4622 ( .B1(REG1_REG_8__SCAN_IN), .B2(keyinput15), .C1(
        D_REG_14__SCAN_IN), .C2(keyinput36), .A(n3913), .ZN(n3918) );
  AOI22_X1 U4623 ( .A1(REG1_REG_10__SCAN_IN), .A2(keyinput25), .B1(
        REG1_REG_12__SCAN_IN), .B2(keyinput45), .ZN(n3914) );
  OAI221_X1 U4624 ( .B1(REG1_REG_10__SCAN_IN), .B2(keyinput25), .C1(
        REG1_REG_12__SCAN_IN), .C2(keyinput45), .A(n3914), .ZN(n3917) );
  AOI22_X1 U4625 ( .A1(REG0_REG_7__SCAN_IN), .A2(keyinput27), .B1(
        REG0_REG_13__SCAN_IN), .B2(keyinput7), .ZN(n3915) );
  OAI221_X1 U4626 ( .B1(REG0_REG_7__SCAN_IN), .B2(keyinput27), .C1(
        REG0_REG_13__SCAN_IN), .C2(keyinput7), .A(n3915), .ZN(n3916) );
  NOR4_X1 U4627 ( .A1(n3919), .A2(n3918), .A3(n3917), .A4(n3916), .ZN(n3920)
         );
  NAND4_X1 U4628 ( .A1(n3923), .A2(n3922), .A3(n3921), .A4(n3920), .ZN(n3976)
         );
  AOI22_X1 U4629 ( .A1(n3926), .A2(keyinput57), .B1(n3925), .B2(keyinput60), 
        .ZN(n3924) );
  OAI221_X1 U4630 ( .B1(n3926), .B2(keyinput57), .C1(n3925), .C2(keyinput60), 
        .A(n3924), .ZN(n3936) );
  INV_X1 U4631 ( .A(REG2_REG_17__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4632 ( .A1(n3929), .A2(keyinput31), .B1(n3928), .B2(keyinput3), 
        .ZN(n3927) );
  OAI221_X1 U4633 ( .B1(n3929), .B2(keyinput31), .C1(n3928), .C2(keyinput3), 
        .A(n3927), .ZN(n3935) );
  AOI22_X1 U4634 ( .A1(ADDR_REG_18__SCAN_IN), .A2(keyinput17), .B1(
        IR_REG_25__SCAN_IN), .B2(keyinput1), .ZN(n3930) );
  OAI221_X1 U4635 ( .B1(ADDR_REG_18__SCAN_IN), .B2(keyinput17), .C1(
        IR_REG_25__SCAN_IN), .C2(keyinput1), .A(n3930), .ZN(n3934) );
  XNOR2_X1 U4636 ( .A(REG1_REG_1__SCAN_IN), .B(keyinput61), .ZN(n3932) );
  XNOR2_X1 U4637 ( .A(IR_REG_31__SCAN_IN), .B(keyinput53), .ZN(n3931) );
  NAND2_X1 U4638 ( .A1(n3932), .A2(n3931), .ZN(n3933) );
  NOR4_X1 U4639 ( .A1(n3936), .A2(n3935), .A3(n3934), .A4(n3933), .ZN(n3974)
         );
  AOI22_X1 U4640 ( .A1(REG3_REG_6__SCAN_IN), .A2(keyinput55), .B1(
        IR_REG_28__SCAN_IN), .B2(keyinput11), .ZN(n3937) );
  OAI221_X1 U4641 ( .B1(REG3_REG_6__SCAN_IN), .B2(keyinput55), .C1(
        IR_REG_28__SCAN_IN), .C2(keyinput11), .A(n3937), .ZN(n3944) );
  AOI22_X1 U4642 ( .A1(DATAO_REG_18__SCAN_IN), .A2(keyinput44), .B1(
        REG1_REG_29__SCAN_IN), .B2(keyinput43), .ZN(n3938) );
  OAI221_X1 U4643 ( .B1(DATAO_REG_18__SCAN_IN), .B2(keyinput44), .C1(
        REG1_REG_29__SCAN_IN), .C2(keyinput43), .A(n3938), .ZN(n3943) );
  AOI22_X1 U4644 ( .A1(REG1_REG_31__SCAN_IN), .A2(keyinput41), .B1(
        IR_REG_8__SCAN_IN), .B2(keyinput28), .ZN(n3939) );
  OAI221_X1 U4645 ( .B1(REG1_REG_31__SCAN_IN), .B2(keyinput41), .C1(
        IR_REG_8__SCAN_IN), .C2(keyinput28), .A(n3939), .ZN(n3942) );
  AOI22_X1 U4646 ( .A1(IR_REG_12__SCAN_IN), .A2(keyinput47), .B1(
        IR_REG_23__SCAN_IN), .B2(keyinput52), .ZN(n3940) );
  OAI221_X1 U4647 ( .B1(IR_REG_12__SCAN_IN), .B2(keyinput47), .C1(
        IR_REG_23__SCAN_IN), .C2(keyinput52), .A(n3940), .ZN(n3941) );
  NOR4_X1 U4648 ( .A1(n3944), .A2(n3943), .A3(n3942), .A4(n3941), .ZN(n3973)
         );
  AOI22_X1 U4649 ( .A1(n3947), .A2(keyinput49), .B1(keyinput21), .B2(n3946), 
        .ZN(n3945) );
  OAI221_X1 U4650 ( .B1(n3947), .B2(keyinput49), .C1(n3946), .C2(keyinput21), 
        .A(n3945), .ZN(n3958) );
  AOI22_X1 U4651 ( .A1(n3950), .A2(keyinput59), .B1(keyinput20), .B2(n3949), 
        .ZN(n3948) );
  OAI221_X1 U4652 ( .B1(n3950), .B2(keyinput59), .C1(n3949), .C2(keyinput20), 
        .A(n3948), .ZN(n3957) );
  AOI22_X1 U4653 ( .A1(n3952), .A2(keyinput29), .B1(n4542), .B2(keyinput9), 
        .ZN(n3951) );
  OAI221_X1 U4654 ( .B1(n3952), .B2(keyinput29), .C1(n4542), .C2(keyinput9), 
        .A(n3951), .ZN(n3956) );
  XNOR2_X1 U4655 ( .A(IR_REG_18__SCAN_IN), .B(keyinput23), .ZN(n3954) );
  XNOR2_X1 U4656 ( .A(keyinput2), .B(DATAI_19_), .ZN(n3953) );
  NAND2_X1 U4657 ( .A1(n3954), .A2(n3953), .ZN(n3955) );
  NOR4_X1 U4658 ( .A1(n3958), .A2(n3957), .A3(n3956), .A4(n3955), .ZN(n3972)
         );
  INV_X1 U4659 ( .A(D_REG_31__SCAN_IN), .ZN(n4745) );
  INV_X1 U4660 ( .A(D_REG_3__SCAN_IN), .ZN(n4747) );
  AOI22_X1 U4661 ( .A1(n4745), .A2(keyinput0), .B1(keyinput46), .B2(n4747), 
        .ZN(n3959) );
  OAI221_X1 U4662 ( .B1(n4745), .B2(keyinput0), .C1(n4747), .C2(keyinput46), 
        .A(n3959), .ZN(n3970) );
  AOI22_X1 U4663 ( .A1(n3961), .A2(keyinput12), .B1(n4746), .B2(keyinput58), 
        .ZN(n3960) );
  OAI221_X1 U4664 ( .B1(n3961), .B2(keyinput12), .C1(n4746), .C2(keyinput58), 
        .A(n3960), .ZN(n3969) );
  INV_X1 U4665 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4666 ( .A1(n2661), .A2(keyinput39), .B1(keyinput6), .B2(n3963), 
        .ZN(n3962) );
  OAI221_X1 U4667 ( .B1(n2661), .B2(keyinput39), .C1(n3963), .C2(keyinput6), 
        .A(n3962), .ZN(n3968) );
  INV_X1 U4668 ( .A(REG1_REG_16__SCAN_IN), .ZN(n3966) );
  INV_X1 U4669 ( .A(REG1_REG_21__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U4670 ( .A1(n3966), .A2(keyinput33), .B1(n3965), .B2(keyinput50), 
        .ZN(n3964) );
  OAI221_X1 U4671 ( .B1(n3966), .B2(keyinput33), .C1(n3965), .C2(keyinput50), 
        .A(n3964), .ZN(n3967) );
  NOR4_X1 U4672 ( .A1(n3970), .A2(n3969), .A3(n3968), .A4(n3967), .ZN(n3971)
         );
  NAND4_X1 U4673 ( .A1(n3974), .A2(n3973), .A3(n3972), .A4(n3971), .ZN(n3975)
         );
  AOI211_X1 U4674 ( .C1(n3978), .C2(n3977), .A(n3976), .B(n3975), .ZN(n3979)
         );
  XOR2_X1 U4675 ( .A(n3980), .B(n3979), .Z(U3554) );
  MUX2_X1 U4676 ( .A(n3981), .B(DATAO_REG_3__SCAN_IN), .S(n3982), .Z(U3553) );
  MUX2_X1 U4677 ( .A(n2690), .B(DATAO_REG_2__SCAN_IN), .S(n3982), .Z(U3552) );
  MUX2_X1 U4678 ( .A(n3983), .B(DATAO_REG_0__SCAN_IN), .S(n3982), .Z(U3550) );
  INV_X1 U4679 ( .A(IR_REG_0__SCAN_IN), .ZN(n4769) );
  NAND3_X1 U4680 ( .A1(n4713), .A2(n3985), .A3(IR_REG_0__SCAN_IN), .ZN(n3992)
         );
  AOI22_X1 U4681 ( .A1(n4711), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n3991) );
  OAI21_X1 U4682 ( .B1(REG2_REG_0__SCAN_IN), .B2(n3986), .A(n3984), .ZN(n3989)
         );
  AOI21_X1 U4683 ( .B1(n3986), .B2(n3985), .A(IR_REG_0__SCAN_IN), .ZN(n3988)
         );
  NAND2_X1 U4684 ( .A1(n3989), .A2(n4769), .ZN(n3996) );
  OAI211_X1 U4685 ( .C1(n3989), .C2(n3988), .A(n3996), .B(n3987), .ZN(n3990)
         );
  NAND3_X1 U4686 ( .A1(n3992), .A2(n3991), .A3(n3990), .ZN(U3240) );
  AOI21_X1 U4687 ( .B1(n4606), .B2(n3993), .A(n4617), .ZN(n3994) );
  OAI21_X1 U4688 ( .B1(n3995), .B2(n4606), .A(n3994), .ZN(n3997) );
  NAND3_X1 U4689 ( .A1(n3997), .A2(U4043), .A3(n3996), .ZN(n4024) );
  AOI22_X1 U4690 ( .A1(n4711), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3998) );
  OAI21_X1 U4691 ( .B1(n4718), .B2(n3999), .A(n3998), .ZN(n4000) );
  INV_X1 U4692 ( .A(n4000), .ZN(n4013) );
  MUX2_X1 U4693 ( .A(n4001), .B(REG2_REG_2__SCAN_IN), .S(n4615), .Z(n4004) );
  NAND3_X1 U4694 ( .A1(n4004), .A2(n4003), .A3(n4002), .ZN(n4005) );
  NAND3_X1 U4695 ( .A1(n4666), .A2(n4006), .A3(n4005), .ZN(n4012) );
  INV_X1 U4696 ( .A(n4007), .ZN(n4008) );
  OAI211_X1 U4697 ( .C1(n4010), .C2(n4009), .A(n4713), .B(n4008), .ZN(n4011)
         );
  NAND4_X1 U4698 ( .A1(n4024), .A2(n4013), .A3(n4012), .A4(n4011), .ZN(U3242)
         );
  AOI21_X1 U4699 ( .B1(n4711), .B2(ADDR_REG_4__SCAN_IN), .A(n4014), .ZN(n4023)
         );
  XOR2_X1 U4700 ( .A(REG2_REG_4__SCAN_IN), .B(n4015), .Z(n4019) );
  AOI21_X1 U4701 ( .B1(n4790), .B2(n4017), .A(n4016), .ZN(n4018) );
  AOI22_X1 U4702 ( .A1(n4666), .A2(n4019), .B1(n4713), .B2(n4018), .ZN(n4022)
         );
  NAND2_X1 U4703 ( .A1(n4020), .A2(n4614), .ZN(n4021) );
  NAND4_X1 U4704 ( .A1(n4024), .A2(n4023), .A3(n4022), .A4(n4021), .ZN(U3244)
         );
  INV_X1 U4705 ( .A(n4612), .ZN(n4054) );
  NAND2_X1 U4706 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4759), .ZN(n4037) );
  INV_X1 U4707 ( .A(n4759), .ZN(n4677) );
  AOI22_X1 U4708 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4759), .B1(n4677), .B2(
        n4025), .ZN(n4674) );
  NAND2_X1 U4709 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4762), .ZN(n4034) );
  INV_X1 U4710 ( .A(n4762), .ZN(n4650) );
  INV_X1 U4711 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U4712 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4762), .B1(n4650), .B2(
        n4026), .ZN(n4644) );
  NAND2_X1 U4713 ( .A1(n4043), .A2(REG1_REG_9__SCAN_IN), .ZN(n4031) );
  INV_X1 U4714 ( .A(n4043), .ZN(n4766) );
  AOI22_X1 U4715 ( .A1(n4043), .A2(REG1_REG_9__SCAN_IN), .B1(n3288), .B2(n4766), .ZN(n4623) );
  INV_X1 U4716 ( .A(n4044), .ZN(n4028) );
  AOI22_X1 U4717 ( .A1(n4029), .A2(REG1_REG_8__SCAN_IN), .B1(n4028), .B2(n4027), .ZN(n4030) );
  INV_X1 U4718 ( .A(n4030), .ZN(n4622) );
  NAND2_X1 U4719 ( .A1(n4623), .A2(n4622), .ZN(n4621) );
  NAND2_X1 U4720 ( .A1(n4031), .A2(n4621), .ZN(n4032) );
  NAND2_X1 U4721 ( .A1(n4632), .A2(n4032), .ZN(n4033) );
  NAND2_X1 U4722 ( .A1(n4654), .A2(n4035), .ZN(n4036) );
  OAI211_X1 U4723 ( .C1(n4038), .C2(REG1_REG_14__SCAN_IN), .A(n4713), .B(n4073), .ZN(n4041) );
  AOI21_X1 U4724 ( .B1(n4711), .B2(ADDR_REG_14__SCAN_IN), .A(n4039), .ZN(n4040) );
  OAI211_X1 U4725 ( .C1(n4718), .C2(n4054), .A(n4041), .B(n4040), .ZN(n4058)
         );
  INV_X1 U4726 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4056) );
  NAND2_X1 U4727 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4762), .ZN(n4050) );
  AOI22_X1 U4728 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4762), .B1(n4650), .B2(
        n3272), .ZN(n4647) );
  NAND2_X1 U4729 ( .A1(n4043), .A2(REG2_REG_9__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U4730 ( .A1(n4043), .A2(REG2_REG_9__SCAN_IN), .B1(n4042), .B2(n4766), .ZN(n4626) );
  INV_X1 U4731 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4721) );
  NAND2_X1 U4732 ( .A1(n4632), .A2(n4048), .ZN(n4049) );
  NAND2_X1 U4733 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4634), .ZN(n4633) );
  NAND2_X1 U4734 ( .A1(n4049), .A2(n4633), .ZN(n4646) );
  NAND2_X1 U4735 ( .A1(n4647), .A2(n4646), .ZN(n4645) );
  NAND2_X1 U4736 ( .A1(n4654), .A2(n4051), .ZN(n4052) );
  INV_X1 U4737 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4665) );
  NOR2_X1 U4738 ( .A1(n4665), .A2(n4677), .ZN(n4664) );
  AOI211_X1 U4739 ( .C1(n4056), .C2(n4055), .A(n4062), .B(n4707), .ZN(n4057)
         );
  OR2_X1 U4740 ( .A1(n4058), .A2(n4057), .ZN(U3254) );
  INV_X1 U4741 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4059) );
  MUX2_X1 U4742 ( .A(REG2_REG_19__SCAN_IN), .B(n4059), .S(n4611), .Z(n4068) );
  INV_X1 U4743 ( .A(n4069), .ZN(n4753) );
  INV_X1 U4744 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U4745 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4753), .B1(n4069), .B2(
        n4060), .ZN(n4709) );
  NOR2_X1 U4746 ( .A1(n4080), .A2(REG2_REG_17__SCAN_IN), .ZN(n4061) );
  AOI21_X1 U4747 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4080), .A(n4061), .ZN(n4699) );
  NAND2_X1 U4748 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4071), .ZN(n4064) );
  OAI21_X1 U4749 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4071), .A(n4064), .ZN(n4679) );
  INV_X1 U4750 ( .A(n4076), .ZN(n4756) );
  NAND2_X1 U4751 ( .A1(n4065), .A2(n4756), .ZN(n4066) );
  INV_X1 U4752 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4688) );
  AOI21_X1 U4753 ( .B1(n4069), .B2(REG2_REG_18__SCAN_IN), .A(n4708), .ZN(n4067) );
  XOR2_X1 U4754 ( .A(n4068), .B(n4067), .Z(n4091) );
  INV_X1 U4755 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4081) );
  AOI22_X1 U4756 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4069), .B1(n4753), .B2(
        n4081), .ZN(n4715) );
  NAND2_X1 U4757 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4071), .ZN(n4075) );
  INV_X1 U4758 ( .A(n4071), .ZN(n4758) );
  INV_X1 U4759 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4070) );
  AOI22_X1 U4760 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4071), .B1(n4758), .B2(
        n4070), .ZN(n4685) );
  NAND2_X1 U4761 ( .A1(n4072), .A2(n4612), .ZN(n4074) );
  NAND2_X1 U4762 ( .A1(n4075), .A2(n4683), .ZN(n4077) );
  NOR2_X1 U4763 ( .A1(n4076), .A2(n4077), .ZN(n4078) );
  XNOR2_X1 U4764 ( .A(n4077), .B(n4076), .ZN(n4693) );
  NOR2_X1 U4765 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4693), .ZN(n4694) );
  INV_X1 U4766 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4079) );
  AOI22_X1 U4767 ( .A1(n4080), .A2(n4079), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4754), .ZN(n4702) );
  INV_X1 U4768 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4082) );
  MUX2_X1 U4769 ( .A(n4082), .B(REG1_REG_19__SCAN_IN), .S(n4611), .Z(n4083) );
  XNOR2_X1 U4770 ( .A(n4084), .B(n4083), .ZN(n4089) );
  AOI21_X1 U4771 ( .B1(n4711), .B2(ADDR_REG_19__SCAN_IN), .A(n4085), .ZN(n4086) );
  OAI21_X1 U4772 ( .B1(n4718), .B2(n4087), .A(n4086), .ZN(n4088) );
  AOI21_X1 U4773 ( .B1(n4089), .B2(n4713), .A(n4088), .ZN(n4090) );
  OAI21_X1 U4774 ( .B1(n4091), .B2(n4707), .A(n4090), .ZN(U3259) );
  XNOR2_X1 U4775 ( .A(n4092), .B(n4095), .ZN(n4093) );
  NAND2_X1 U4776 ( .A1(n4093), .A2(n4529), .ZN(n4385) );
  XOR2_X1 U4777 ( .A(n4095), .B(n4094), .Z(n4388) );
  NAND2_X1 U4778 ( .A1(n4388), .A2(n4312), .ZN(n4105) );
  INV_X1 U4779 ( .A(n4096), .ZN(n4097) );
  OAI21_X1 U4780 ( .B1(n4114), .B2(n4098), .A(n4097), .ZN(n4540) );
  INV_X1 U4781 ( .A(n4540), .ZN(n4103) );
  AOI22_X1 U4782 ( .A1(n4099), .A2(n4736), .B1(n4744), .B2(
        REG2_REG_27__SCAN_IN), .ZN(n4101) );
  AOI22_X1 U4783 ( .A1(n4339), .A2(n4396), .B1(n4340), .B2(n4383), .ZN(n4100)
         );
  OAI211_X1 U4784 ( .C1(n4386), .C2(n4344), .A(n4101), .B(n4100), .ZN(n4102)
         );
  AOI21_X1 U4785 ( .B1(n4103), .B2(n4738), .A(n4102), .ZN(n4104) );
  OAI211_X1 U4786 ( .C1(n4744), .C2(n4385), .A(n4105), .B(n4104), .ZN(U3263)
         );
  XNOR2_X1 U4787 ( .A(n4106), .B(n4107), .ZN(n4392) );
  INV_X1 U4788 ( .A(n4392), .ZN(n4121) );
  XNOR2_X1 U4789 ( .A(n4108), .B(n4107), .ZN(n4113) );
  NOR2_X1 U4790 ( .A1(n4116), .A2(n4500), .ZN(n4109) );
  AOI21_X1 U4791 ( .B1(n4110), .B2(n4495), .A(n4109), .ZN(n4112) );
  NAND2_X1 U4792 ( .A1(n4405), .A2(n4519), .ZN(n4111) );
  OAI211_X1 U4793 ( .C1(n4113), .C2(n4505), .A(n4112), .B(n4111), .ZN(n4391)
         );
  INV_X1 U4794 ( .A(n4114), .ZN(n4115) );
  OAI21_X1 U4795 ( .B1(n2142), .B2(n4116), .A(n4115), .ZN(n4544) );
  AOI22_X1 U4796 ( .A1(n4744), .A2(REG2_REG_26__SCAN_IN), .B1(n4117), .B2(
        n4736), .ZN(n4118) );
  OAI21_X1 U4797 ( .B1(n4544), .B2(n4371), .A(n4118), .ZN(n4119) );
  AOI21_X1 U4798 ( .B1(n4391), .B2(n4722), .A(n4119), .ZN(n4120) );
  OAI21_X1 U4799 ( .B1(n4121), .B2(n4375), .A(n4120), .ZN(U3264) );
  XNOR2_X1 U4800 ( .A(n4123), .B(n4122), .ZN(n4124) );
  NAND2_X1 U4801 ( .A1(n4124), .A2(n4529), .ZN(n4398) );
  XNOR2_X1 U4802 ( .A(n4126), .B(n4125), .ZN(n4401) );
  NAND2_X1 U4803 ( .A1(n4401), .A2(n4312), .ZN(n4138) );
  INV_X1 U4804 ( .A(n4146), .ZN(n4129) );
  OAI21_X1 U4805 ( .B1(n4129), .B2(n4128), .A(n4127), .ZN(n4548) );
  INV_X1 U4806 ( .A(n4548), .ZN(n4136) );
  INV_X1 U4807 ( .A(n4396), .ZN(n4134) );
  AOI22_X1 U4808 ( .A1(n4395), .A2(n4340), .B1(n4339), .B2(n4130), .ZN(n4133)
         );
  AOI22_X1 U4809 ( .A1(n4744), .A2(REG2_REG_25__SCAN_IN), .B1(n4131), .B2(
        n4736), .ZN(n4132) );
  OAI211_X1 U4810 ( .C1(n4134), .C2(n4344), .A(n4133), .B(n4132), .ZN(n4135)
         );
  AOI21_X1 U4811 ( .B1(n4136), .B2(n4738), .A(n4135), .ZN(n4137) );
  OAI211_X1 U4812 ( .C1(n4744), .C2(n4398), .A(n4138), .B(n4137), .ZN(U3265)
         );
  NAND2_X1 U4813 ( .A1(n4140), .A2(n4139), .ZN(n4142) );
  INV_X1 U4814 ( .A(n4144), .ZN(n4141) );
  XNOR2_X1 U4815 ( .A(n4142), .B(n4141), .ZN(n4143) );
  NAND2_X1 U4816 ( .A1(n4143), .A2(n4529), .ZN(n4407) );
  XNOR2_X1 U4817 ( .A(n4145), .B(n4144), .ZN(n4410) );
  NAND2_X1 U4818 ( .A1(n4410), .A2(n4312), .ZN(n4155) );
  OAI21_X1 U4819 ( .B1(n4170), .B2(n4147), .A(n4146), .ZN(n4552) );
  INV_X1 U4820 ( .A(n4552), .ZN(n4153) );
  AOI22_X1 U4821 ( .A1(n4404), .A2(n4340), .B1(n4339), .B2(n4188), .ZN(n4150)
         );
  AOI22_X1 U4822 ( .A1(n4744), .A2(REG2_REG_24__SCAN_IN), .B1(n4148), .B2(
        n4736), .ZN(n4149) );
  OAI211_X1 U4823 ( .C1(n4151), .C2(n4344), .A(n4150), .B(n4149), .ZN(n4152)
         );
  AOI21_X1 U4824 ( .B1(n4153), .B2(n4738), .A(n4152), .ZN(n4154) );
  OAI211_X1 U4825 ( .C1(n4744), .C2(n4407), .A(n4155), .B(n4154), .ZN(U3266)
         );
  XNOR2_X1 U4826 ( .A(n4156), .B(n4162), .ZN(n4414) );
  INV_X1 U4827 ( .A(n4414), .ZN(n4175) );
  NAND2_X1 U4828 ( .A1(n4158), .A2(n4157), .ZN(n4196) );
  INV_X1 U4829 ( .A(n4159), .ZN(n4160) );
  AOI21_X1 U4830 ( .B1(n4196), .B2(n4199), .A(n4160), .ZN(n4187) );
  INV_X1 U4831 ( .A(n4176), .ZN(n4186) );
  OAI21_X1 U4832 ( .B1(n4187), .B2(n4186), .A(n4161), .ZN(n4164) );
  INV_X1 U4833 ( .A(n4162), .ZN(n4163) );
  XNOR2_X1 U4834 ( .A(n4164), .B(n4163), .ZN(n4167) );
  OAI22_X1 U4835 ( .A1(n4399), .A2(n4522), .B1(n4500), .B2(n4168), .ZN(n4165)
         );
  AOI21_X1 U4836 ( .B1(n4519), .B2(n4423), .A(n4165), .ZN(n4166) );
  OAI21_X1 U4837 ( .B1(n4167), .B2(n4505), .A(n4166), .ZN(n4413) );
  NOR2_X1 U4838 ( .A1(n4181), .A2(n4168), .ZN(n4169) );
  OR2_X1 U4839 ( .A1(n4170), .A2(n4169), .ZN(n4556) );
  AOI22_X1 U4840 ( .A1(n4744), .A2(REG2_REG_23__SCAN_IN), .B1(n4171), .B2(
        n4736), .ZN(n4172) );
  OAI21_X1 U4841 ( .B1(n4556), .B2(n4371), .A(n4172), .ZN(n4173) );
  AOI21_X1 U4842 ( .B1(n4413), .B2(n4722), .A(n4173), .ZN(n4174) );
  OAI21_X1 U4843 ( .B1(n4175), .B2(n4375), .A(n4174), .ZN(U3267) );
  NAND2_X1 U4844 ( .A1(n4177), .A2(n4176), .ZN(n4178) );
  NAND2_X1 U4845 ( .A1(n4179), .A2(n4178), .ZN(n4417) );
  NOR2_X1 U4846 ( .A1(n4200), .A2(n4191), .ZN(n4180) );
  OR2_X1 U4847 ( .A1(n4181), .A2(n4180), .ZN(n4560) );
  INV_X1 U4848 ( .A(n4560), .ZN(n4185) );
  INV_X1 U4849 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4183) );
  OAI22_X1 U4850 ( .A1(n4722), .A2(n4183), .B1(n4182), .B2(n4719), .ZN(n4184)
         );
  AOI21_X1 U4851 ( .B1(n4185), .B2(n4738), .A(n4184), .ZN(n4195) );
  XNOR2_X1 U4852 ( .A(n4187), .B(n4186), .ZN(n4193) );
  NAND2_X1 U4853 ( .A1(n4220), .A2(n4519), .ZN(n4190) );
  NAND2_X1 U4854 ( .A1(n4188), .A2(n4495), .ZN(n4189) );
  OAI211_X1 U4855 ( .C1(n4500), .C2(n4191), .A(n4190), .B(n4189), .ZN(n4192)
         );
  AOI21_X1 U4856 ( .B1(n4193), .B2(n4529), .A(n4192), .ZN(n4418) );
  OR2_X1 U4857 ( .A1(n4418), .A2(n4744), .ZN(n4194) );
  OAI211_X1 U4858 ( .C1(n4417), .C2(n4375), .A(n4195), .B(n4194), .ZN(U3268)
         );
  XNOR2_X1 U4859 ( .A(n4196), .B(n4199), .ZN(n4197) );
  NAND2_X1 U4860 ( .A1(n4197), .A2(n4529), .ZN(n4425) );
  XOR2_X1 U4861 ( .A(n4199), .B(n4198), .Z(n4428) );
  NAND2_X1 U4862 ( .A1(n4428), .A2(n4312), .ZN(n4211) );
  INV_X1 U4863 ( .A(n4218), .ZN(n4203) );
  INV_X1 U4864 ( .A(n4200), .ZN(n4201) );
  OAI21_X1 U4865 ( .B1(n4203), .B2(n4202), .A(n4201), .ZN(n4564) );
  INV_X1 U4866 ( .A(n4564), .ZN(n4209) );
  AOI22_X1 U4867 ( .A1(n4340), .A2(n4422), .B1(n4339), .B2(n4242), .ZN(n4206)
         );
  AOI22_X1 U4868 ( .A1(n4744), .A2(REG2_REG_21__SCAN_IN), .B1(n4204), .B2(
        n4736), .ZN(n4205) );
  OAI211_X1 U4869 ( .C1(n4207), .C2(n4344), .A(n4206), .B(n4205), .ZN(n4208)
         );
  AOI21_X1 U4870 ( .B1(n4209), .B2(n4738), .A(n4208), .ZN(n4210) );
  OAI211_X1 U4871 ( .C1(n4744), .C2(n4425), .A(n4211), .B(n4210), .ZN(U3269)
         );
  NOR2_X1 U4872 ( .A1(n2079), .A2(n4212), .ZN(n4213) );
  XNOR2_X1 U4873 ( .A(n4213), .B(n4216), .ZN(n4435) );
  AOI21_X1 U4874 ( .B1(n4231), .B2(n4215), .A(n4214), .ZN(n4217) );
  XNOR2_X1 U4875 ( .A(n4217), .B(n4216), .ZN(n4437) );
  NAND2_X1 U4876 ( .A1(n4437), .A2(n4312), .ZN(n4229) );
  INV_X1 U4877 ( .A(n4245), .ZN(n4219) );
  OAI21_X1 U4878 ( .B1(n4219), .B2(n4430), .A(n4218), .ZN(n4568) );
  INV_X1 U4879 ( .A(n4568), .ZN(n4227) );
  AOI22_X1 U4880 ( .A1(n4221), .A2(n4220), .B1(n4339), .B2(n4433), .ZN(n4224)
         );
  AOI22_X1 U4881 ( .A1(n4744), .A2(REG2_REG_20__SCAN_IN), .B1(n4222), .B2(
        n4736), .ZN(n4223) );
  OAI211_X1 U4882 ( .C1(n4430), .C2(n4225), .A(n4224), .B(n4223), .ZN(n4226)
         );
  AOI21_X1 U4883 ( .B1(n4227), .B2(n4738), .A(n4226), .ZN(n4228) );
  OAI211_X1 U4884 ( .C1(n4435), .C2(n4230), .A(n4229), .B(n4228), .ZN(U3270)
         );
  XOR2_X1 U4885 ( .A(n4238), .B(n4231), .Z(n4441) );
  INV_X1 U4886 ( .A(n4441), .ZN(n4252) );
  INV_X1 U4887 ( .A(n4232), .ZN(n4233) );
  NOR2_X1 U4888 ( .A1(n4234), .A2(n4233), .ZN(n4261) );
  INV_X1 U4889 ( .A(n4235), .ZN(n4236) );
  AOI21_X1 U4890 ( .B1(n4261), .B2(n4237), .A(n4236), .ZN(n4239) );
  XNOR2_X1 U4891 ( .A(n4239), .B(n4238), .ZN(n4240) );
  NAND2_X1 U4892 ( .A1(n4240), .A2(n4529), .ZN(n4244) );
  NOR2_X1 U4893 ( .A1(n4246), .A2(n4500), .ZN(n4241) );
  AOI21_X1 U4894 ( .B1(n4242), .B2(n4495), .A(n4241), .ZN(n4243) );
  OAI211_X1 U4895 ( .C1(n4281), .C2(n4484), .A(n4244), .B(n4243), .ZN(n4440)
         );
  INV_X1 U4896 ( .A(n4257), .ZN(n4247) );
  OAI21_X1 U4897 ( .B1(n4247), .B2(n4246), .A(n4245), .ZN(n4572) );
  NOR2_X1 U4898 ( .A1(n4572), .A2(n4371), .ZN(n4250) );
  OAI22_X1 U4899 ( .A1(n4722), .A2(n4059), .B1(n4248), .B2(n4719), .ZN(n4249)
         );
  AOI211_X1 U4900 ( .C1(n4440), .C2(n4722), .A(n4250), .B(n4249), .ZN(n4251)
         );
  OAI21_X1 U4901 ( .B1(n4252), .B2(n4375), .A(n4251), .ZN(U3271) );
  OAI21_X1 U4902 ( .B1(n4254), .B2(n4260), .A(n4253), .ZN(n4255) );
  INV_X1 U4903 ( .A(n4255), .ZN(n4445) );
  AOI22_X1 U4904 ( .A1(n4744), .A2(REG2_REG_18__SCAN_IN), .B1(n4256), .B2(
        n4736), .ZN(n4269) );
  OAI211_X1 U4905 ( .C1(n4275), .C2(n4259), .A(n4258), .B(n4257), .ZN(n4443)
         );
  XNOR2_X1 U4906 ( .A(n4261), .B(n4260), .ZN(n4266) );
  AOI22_X1 U4907 ( .A1(n4433), .A2(n4495), .B1(n4518), .B2(n4262), .ZN(n4263)
         );
  OAI21_X1 U4908 ( .B1(n4264), .B2(n4484), .A(n4263), .ZN(n4265) );
  AOI21_X1 U4909 ( .B1(n4266), .B2(n4529), .A(n4265), .ZN(n4444) );
  OAI21_X1 U4910 ( .B1(n4611), .B2(n4443), .A(n4444), .ZN(n4267) );
  NAND2_X1 U4911 ( .A1(n4267), .A2(n4722), .ZN(n4268) );
  OAI211_X1 U4912 ( .C1(n4445), .C2(n4375), .A(n4269), .B(n4268), .ZN(U3272)
         );
  INV_X1 U4913 ( .A(n4274), .ZN(n4271) );
  XNOR2_X1 U4914 ( .A(n4270), .B(n4271), .ZN(n4272) );
  NAND2_X1 U4915 ( .A1(n4272), .A2(n4529), .ZN(n4449) );
  XOR2_X1 U4916 ( .A(n4274), .B(n4273), .Z(n4452) );
  NAND2_X1 U4917 ( .A1(n4452), .A2(n4312), .ZN(n4285) );
  INV_X1 U4918 ( .A(n4275), .ZN(n4276) );
  OAI21_X1 U4919 ( .B1(n4291), .B2(n4277), .A(n4276), .ZN(n4577) );
  INV_X1 U4920 ( .A(n4577), .ZN(n4283) );
  AOI22_X1 U4921 ( .A1(n4340), .A2(n4446), .B1(n4339), .B2(n4459), .ZN(n4280)
         );
  AOI22_X1 U4922 ( .A1(n4744), .A2(REG2_REG_17__SCAN_IN), .B1(n4278), .B2(
        n4736), .ZN(n4279) );
  OAI211_X1 U4923 ( .C1(n4281), .C2(n4344), .A(n4280), .B(n4279), .ZN(n4282)
         );
  AOI21_X1 U4924 ( .B1(n4283), .B2(n4738), .A(n4282), .ZN(n4284) );
  OAI211_X1 U4925 ( .C1(n4744), .C2(n4449), .A(n4285), .B(n4284), .ZN(U3273)
         );
  NAND2_X1 U4926 ( .A1(n4286), .A2(n4294), .ZN(n4287) );
  NAND2_X1 U4927 ( .A1(n4288), .A2(n4287), .ZN(n4455) );
  AND2_X1 U4928 ( .A1(n4313), .A2(n4289), .ZN(n4290) );
  NOR2_X1 U4929 ( .A1(n4291), .A2(n4290), .ZN(n4580) );
  OAI22_X1 U4930 ( .A1(n4722), .A2(n4688), .B1(n4292), .B2(n4719), .ZN(n4293)
         );
  AOI21_X1 U4931 ( .B1(n4580), .B2(n4738), .A(n4293), .ZN(n4303) );
  XNOR2_X1 U4932 ( .A(n4295), .B(n2105), .ZN(n4301) );
  NAND2_X1 U4933 ( .A1(n4467), .A2(n4519), .ZN(n4298) );
  NAND2_X1 U4934 ( .A1(n4296), .A2(n4495), .ZN(n4297) );
  OAI211_X1 U4935 ( .C1(n4500), .C2(n4299), .A(n4298), .B(n4297), .ZN(n4300)
         );
  AOI21_X1 U4936 ( .B1(n4301), .B2(n4529), .A(n4300), .ZN(n4454) );
  OR2_X1 U4937 ( .A1(n4454), .A2(n4744), .ZN(n4302) );
  OAI211_X1 U4938 ( .C1(n4455), .C2(n4375), .A(n4303), .B(n4302), .ZN(U3274)
         );
  NAND2_X1 U4939 ( .A1(n4332), .A2(n4304), .ZN(n4306) );
  XNOR2_X1 U4940 ( .A(n4306), .B(n4305), .ZN(n4307) );
  NAND2_X1 U4941 ( .A1(n4307), .A2(n4529), .ZN(n4461) );
  OR2_X1 U4942 ( .A1(n3268), .A2(n4308), .ZN(n4328) );
  NAND2_X1 U4943 ( .A1(n4328), .A2(n4309), .ZN(n4311) );
  XNOR2_X1 U4944 ( .A(n4311), .B(n4310), .ZN(n4464) );
  NAND2_X1 U4945 ( .A1(n4464), .A2(n4312), .ZN(n4323) );
  INV_X1 U4946 ( .A(n4337), .ZN(n4315) );
  OAI21_X1 U4947 ( .B1(n4315), .B2(n4314), .A(n4313), .ZN(n4585) );
  INV_X1 U4948 ( .A(n4585), .ZN(n4321) );
  AOI22_X1 U4949 ( .A1(n4340), .A2(n4458), .B1(n4339), .B2(n4316), .ZN(n4319)
         );
  AOI22_X1 U4950 ( .A1(n4744), .A2(REG2_REG_15__SCAN_IN), .B1(n4317), .B2(
        n4736), .ZN(n4318) );
  OAI211_X1 U4951 ( .C1(n4450), .C2(n4344), .A(n4319), .B(n4318), .ZN(n4320)
         );
  AOI21_X1 U4952 ( .B1(n4321), .B2(n4738), .A(n4320), .ZN(n4322) );
  OAI211_X1 U4953 ( .C1(n4744), .C2(n4461), .A(n4323), .B(n4322), .ZN(U3275)
         );
  OR2_X1 U4954 ( .A1(n3268), .A2(n4324), .ZN(n4326) );
  NAND2_X1 U4955 ( .A1(n4326), .A2(n4325), .ZN(n4330) );
  AND2_X1 U4956 ( .A1(n4328), .A2(n4327), .ZN(n4329) );
  OAI21_X1 U4957 ( .B1(n4330), .B2(n4334), .A(n4329), .ZN(n4472) );
  INV_X1 U4958 ( .A(n4472), .ZN(n4351) );
  INV_X1 U4959 ( .A(n4331), .ZN(n4335) );
  INV_X1 U4960 ( .A(n4332), .ZN(n4333) );
  AOI21_X1 U4961 ( .B1(n4335), .B2(n4334), .A(n4333), .ZN(n4336) );
  OAI22_X1 U4962 ( .A1(n4351), .A2(n4524), .B1(n4505), .B2(n4336), .ZN(n4470)
         );
  NAND2_X1 U4963 ( .A1(n4470), .A2(n4722), .ZN(n4349) );
  OAI21_X1 U4964 ( .B1(n4368), .B2(n4338), .A(n4337), .ZN(n4589) );
  INV_X1 U4965 ( .A(n4589), .ZN(n4347) );
  AOI22_X1 U4966 ( .A1(n4466), .A2(n4340), .B1(n4339), .B2(n4481), .ZN(n4343)
         );
  AOI22_X1 U4967 ( .A1(n4744), .A2(REG2_REG_14__SCAN_IN), .B1(n4341), .B2(
        n4736), .ZN(n4342) );
  OAI211_X1 U4968 ( .C1(n4345), .C2(n4344), .A(n4343), .B(n4342), .ZN(n4346)
         );
  AOI21_X1 U4969 ( .B1(n4347), .B2(n4738), .A(n4346), .ZN(n4348) );
  OAI211_X1 U4970 ( .C1(n4351), .C2(n4350), .A(n4349), .B(n4348), .ZN(U3276)
         );
  OR2_X1 U4971 ( .A1(n3268), .A2(n4352), .ZN(n4354) );
  NAND2_X1 U4972 ( .A1(n4354), .A2(n4353), .ZN(n4355) );
  XNOR2_X1 U4973 ( .A(n4355), .B(n4361), .ZN(n4476) );
  INV_X1 U4974 ( .A(n4476), .ZN(n4374) );
  INV_X1 U4975 ( .A(n4356), .ZN(n4358) );
  OAI21_X1 U4976 ( .B1(n4359), .B2(n4358), .A(n4357), .ZN(n4360) );
  XOR2_X1 U4977 ( .A(n4361), .B(n4360), .Z(n4364) );
  OAI22_X1 U4978 ( .A1(n4462), .A2(n4522), .B1(n4500), .B2(n4365), .ZN(n4362)
         );
  AOI21_X1 U4979 ( .B1(n4519), .B2(n4496), .A(n4362), .ZN(n4363) );
  OAI21_X1 U4980 ( .B1(n4364), .B2(n4505), .A(n4363), .ZN(n4475) );
  NOR2_X1 U4981 ( .A1(n4366), .A2(n4365), .ZN(n4367) );
  OR2_X1 U4982 ( .A1(n4368), .A2(n4367), .ZN(n4592) );
  AOI22_X1 U4983 ( .A1(n4744), .A2(REG2_REG_13__SCAN_IN), .B1(n4369), .B2(
        n4736), .ZN(n4370) );
  OAI21_X1 U4984 ( .B1(n4592), .B2(n4371), .A(n4370), .ZN(n4372) );
  AOI21_X1 U4985 ( .B1(n4475), .B2(n4722), .A(n4372), .ZN(n4373) );
  OAI21_X1 U4986 ( .B1(n4375), .B2(n4374), .A(n4373), .ZN(U3277) );
  AOI21_X1 U4987 ( .B1(n4380), .B2(n4377), .A(n4376), .ZN(n4618) );
  INV_X1 U4988 ( .A(n4618), .ZN(n4536) );
  INV_X1 U4989 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4381) );
  INV_X1 U4990 ( .A(n4378), .ZN(n4379) );
  AOI21_X1 U4991 ( .B1(n4380), .B2(n4518), .A(n4379), .ZN(n4620) );
  MUX2_X1 U4992 ( .A(n4381), .B(n4620), .S(n4795), .Z(n4382) );
  OAI21_X1 U4993 ( .B1(n4536), .B2(n4533), .A(n4382), .ZN(U3548) );
  INV_X1 U4994 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4389) );
  AOI22_X1 U4995 ( .A1(n4396), .A2(n4519), .B1(n4383), .B2(n4518), .ZN(n4384)
         );
  OAI211_X1 U4996 ( .C1(n4386), .C2(n4522), .A(n4385), .B(n4384), .ZN(n4387)
         );
  AOI21_X1 U4997 ( .B1(n4388), .B2(n4492), .A(n4387), .ZN(n4537) );
  MUX2_X1 U4998 ( .A(n4389), .B(n4537), .S(n4795), .Z(n4390) );
  OAI21_X1 U4999 ( .B1(n4533), .B2(n4540), .A(n4390), .ZN(U3545) );
  INV_X1 U5000 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4393) );
  AOI21_X1 U5001 ( .B1(n4392), .B2(n4492), .A(n4391), .ZN(n4541) );
  MUX2_X1 U5002 ( .A(n4393), .B(n4541), .S(n4795), .Z(n4394) );
  OAI21_X1 U5003 ( .B1(n4533), .B2(n4544), .A(n4394), .ZN(U3544) );
  INV_X1 U5004 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4402) );
  AOI22_X1 U5005 ( .A1(n4396), .A2(n4495), .B1(n4518), .B2(n4395), .ZN(n4397)
         );
  OAI211_X1 U5006 ( .C1(n4399), .C2(n4484), .A(n4398), .B(n4397), .ZN(n4400)
         );
  AOI21_X1 U5007 ( .B1(n4401), .B2(n4492), .A(n4400), .ZN(n4545) );
  MUX2_X1 U5008 ( .A(n4402), .B(n4545), .S(n4795), .Z(n4403) );
  OAI21_X1 U5009 ( .B1(n4533), .B2(n4548), .A(n4403), .ZN(U3543) );
  INV_X1 U5010 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4411) );
  AOI22_X1 U5011 ( .A1(n4405), .A2(n4495), .B1(n4518), .B2(n4404), .ZN(n4406)
         );
  OAI211_X1 U5012 ( .C1(n4408), .C2(n4484), .A(n4407), .B(n4406), .ZN(n4409)
         );
  AOI21_X1 U5013 ( .B1(n4410), .B2(n4492), .A(n4409), .ZN(n4549) );
  MUX2_X1 U5014 ( .A(n4411), .B(n4549), .S(n4795), .Z(n4412) );
  OAI21_X1 U5015 ( .B1(n4533), .B2(n4552), .A(n4412), .ZN(U3542) );
  INV_X1 U5016 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4415) );
  AOI21_X1 U5017 ( .B1(n4414), .B2(n4492), .A(n4413), .ZN(n4553) );
  MUX2_X1 U5018 ( .A(n4415), .B(n4553), .S(n4795), .Z(n4416) );
  OAI21_X1 U5019 ( .B1(n4533), .B2(n4556), .A(n4416), .ZN(U3541) );
  OR2_X1 U5020 ( .A1(n4417), .A2(n4781), .ZN(n4419) );
  NAND2_X1 U5021 ( .A1(n4419), .A2(n4418), .ZN(n4557) );
  MUX2_X1 U5022 ( .A(REG1_REG_22__SCAN_IN), .B(n4557), .S(n4795), .Z(n4420) );
  INV_X1 U5023 ( .A(n4420), .ZN(n4421) );
  OAI21_X1 U5024 ( .B1(n4533), .B2(n4560), .A(n4421), .ZN(U3540) );
  AOI22_X1 U5025 ( .A1(n4423), .A2(n4495), .B1(n4518), .B2(n4422), .ZN(n4424)
         );
  OAI211_X1 U5026 ( .C1(n4426), .C2(n4484), .A(n4425), .B(n4424), .ZN(n4427)
         );
  AOI21_X1 U5027 ( .B1(n4428), .B2(n4492), .A(n4427), .ZN(n4561) );
  MUX2_X1 U5028 ( .A(n3965), .B(n4561), .S(n4795), .Z(n4429) );
  OAI21_X1 U5029 ( .B1(n4533), .B2(n4564), .A(n4429), .ZN(U3539) );
  INV_X1 U5030 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4438) );
  OAI22_X1 U5031 ( .A1(n4431), .A2(n4522), .B1(n4430), .B2(n4500), .ZN(n4432)
         );
  AOI21_X1 U5032 ( .B1(n4519), .B2(n4433), .A(n4432), .ZN(n4434) );
  OAI21_X1 U5033 ( .B1(n4435), .B2(n4505), .A(n4434), .ZN(n4436) );
  AOI21_X1 U5034 ( .B1(n4437), .B2(n4492), .A(n4436), .ZN(n4565) );
  MUX2_X1 U5035 ( .A(n4438), .B(n4565), .S(n4795), .Z(n4439) );
  OAI21_X1 U5036 ( .B1(n4533), .B2(n4568), .A(n4439), .ZN(U3538) );
  AOI21_X1 U5037 ( .B1(n4441), .B2(n4492), .A(n4440), .ZN(n4569) );
  MUX2_X1 U5038 ( .A(n4082), .B(n4569), .S(n4795), .Z(n4442) );
  OAI21_X1 U5039 ( .B1(n4533), .B2(n4572), .A(n4442), .ZN(U3537) );
  OAI211_X1 U5040 ( .C1(n4445), .C2(n4781), .A(n4444), .B(n4443), .ZN(n4573)
         );
  MUX2_X1 U5041 ( .A(REG1_REG_18__SCAN_IN), .B(n4573), .S(n4795), .Z(U3536) );
  AOI22_X1 U5042 ( .A1(n4447), .A2(n4495), .B1(n4518), .B2(n4446), .ZN(n4448)
         );
  OAI211_X1 U5043 ( .C1(n4450), .C2(n4484), .A(n4449), .B(n4448), .ZN(n4451)
         );
  AOI21_X1 U5044 ( .B1(n4452), .B2(n4492), .A(n4451), .ZN(n4575) );
  MUX2_X1 U5045 ( .A(n4575), .B(n4079), .S(n4792), .Z(n4453) );
  OAI21_X1 U5046 ( .B1(n4533), .B2(n4577), .A(n4453), .ZN(U3535) );
  OAI21_X1 U5047 ( .B1(n4455), .B2(n4781), .A(n4454), .ZN(n4578) );
  MUX2_X1 U5048 ( .A(REG1_REG_16__SCAN_IN), .B(n4578), .S(n4795), .Z(n4456) );
  AOI21_X1 U5049 ( .B1(n4490), .B2(n4580), .A(n4456), .ZN(n4457) );
  INV_X1 U5050 ( .A(n4457), .ZN(U3534) );
  AOI22_X1 U5051 ( .A1(n4459), .A2(n4495), .B1(n4518), .B2(n4458), .ZN(n4460)
         );
  OAI211_X1 U5052 ( .C1(n4462), .C2(n4484), .A(n4461), .B(n4460), .ZN(n4463)
         );
  AOI21_X1 U5053 ( .B1(n4464), .B2(n4492), .A(n4463), .ZN(n4583) );
  MUX2_X1 U5054 ( .A(n4583), .B(n4070), .S(n4792), .Z(n4465) );
  OAI21_X1 U5055 ( .B1(n4533), .B2(n4585), .A(n4465), .ZN(U3533) );
  INV_X1 U5056 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4473) );
  AOI22_X1 U5057 ( .A1(n4467), .A2(n4495), .B1(n4466), .B2(n4518), .ZN(n4468)
         );
  OAI21_X1 U5058 ( .B1(n4469), .B2(n4484), .A(n4468), .ZN(n4471) );
  AOI211_X1 U5059 ( .C1(n4778), .C2(n4472), .A(n4471), .B(n4470), .ZN(n4586)
         );
  MUX2_X1 U5060 ( .A(n4473), .B(n4586), .S(n4795), .Z(n4474) );
  OAI21_X1 U5061 ( .B1(n4533), .B2(n4589), .A(n4474), .ZN(U3532) );
  AOI21_X1 U5062 ( .B1(n4492), .B2(n4476), .A(n4475), .ZN(n4590) );
  MUX2_X1 U5063 ( .A(n4025), .B(n4590), .S(n4795), .Z(n4477) );
  OAI21_X1 U5064 ( .B1(n4533), .B2(n4592), .A(n4477), .ZN(U3531) );
  NAND2_X1 U5065 ( .A1(n4478), .A2(n4492), .ZN(n4488) );
  NOR2_X1 U5066 ( .A1(n4479), .A2(n4500), .ZN(n4480) );
  AOI21_X1 U5067 ( .B1(n4481), .B2(n4495), .A(n4480), .ZN(n4482) );
  OAI211_X1 U5068 ( .C1(n4485), .C2(n4484), .A(n4483), .B(n4482), .ZN(n4486)
         );
  INV_X1 U5069 ( .A(n4486), .ZN(n4487) );
  NAND2_X1 U5070 ( .A1(n4488), .A2(n4487), .ZN(n4593) );
  MUX2_X1 U5071 ( .A(REG1_REG_12__SCAN_IN), .B(n4593), .S(n4795), .Z(n4489) );
  AOI21_X1 U5072 ( .B1(n4490), .B2(n4596), .A(n4489), .ZN(n4491) );
  INV_X1 U5073 ( .A(n4491), .ZN(U3530) );
  NAND2_X1 U5074 ( .A1(n4493), .A2(n4492), .ZN(n4503) );
  NAND2_X1 U5075 ( .A1(n4494), .A2(n4519), .ZN(n4498) );
  NAND2_X1 U5076 ( .A1(n4496), .A2(n4495), .ZN(n4497) );
  OAI211_X1 U5077 ( .C1(n4500), .C2(n4499), .A(n4498), .B(n4497), .ZN(n4501)
         );
  INV_X1 U5078 ( .A(n4501), .ZN(n4502) );
  OAI211_X1 U5079 ( .C1(n4505), .C2(n4504), .A(n4503), .B(n4502), .ZN(n4598)
         );
  MUX2_X1 U5080 ( .A(REG1_REG_11__SCAN_IN), .B(n4598), .S(n4795), .Z(n4506) );
  INV_X1 U5081 ( .A(n4506), .ZN(n4507) );
  OAI21_X1 U5082 ( .B1(n4533), .B2(n4601), .A(n4507), .ZN(U3529) );
  OAI21_X1 U5083 ( .B1(n4510), .B2(n4509), .A(n4508), .ZN(n4724) );
  INV_X1 U5084 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4531) );
  NAND2_X1 U5085 ( .A1(n4785), .A2(n4511), .ZN(n4512) );
  XOR2_X1 U5086 ( .A(n4515), .B(n4512), .Z(n4525) );
  INV_X1 U5087 ( .A(n4525), .ZN(n4726) );
  NAND2_X1 U5088 ( .A1(n4514), .A2(n4513), .ZN(n4516) );
  XOR2_X1 U5089 ( .A(n4516), .B(n4515), .Z(n4528) );
  AOI22_X1 U5090 ( .A1(n4520), .A2(n4519), .B1(n4518), .B2(n4517), .ZN(n4521)
         );
  OAI21_X1 U5091 ( .B1(n4523), .B2(n4522), .A(n4521), .ZN(n4527) );
  NOR2_X1 U5092 ( .A1(n4525), .A2(n4524), .ZN(n4526) );
  AOI211_X1 U5093 ( .C1(n4529), .C2(n4528), .A(n4527), .B(n4526), .ZN(n4729)
         );
  INV_X1 U5094 ( .A(n4729), .ZN(n4530) );
  AOI21_X1 U5095 ( .B1(n4778), .B2(n4726), .A(n4530), .ZN(n4602) );
  MUX2_X1 U5096 ( .A(n4531), .B(n4602), .S(n4795), .Z(n4532) );
  OAI21_X1 U5097 ( .B1(n4724), .B2(n4533), .A(n4532), .ZN(U3526) );
  INV_X1 U5098 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4534) );
  MUX2_X1 U5099 ( .A(n4534), .B(n4620), .S(n4789), .Z(n4535) );
  OAI21_X1 U5100 ( .B1(n4536), .B2(n4605), .A(n4535), .ZN(U3516) );
  INV_X1 U5101 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4538) );
  MUX2_X1 U5102 ( .A(n4538), .B(n4537), .S(n4789), .Z(n4539) );
  OAI21_X1 U5103 ( .B1(n4540), .B2(n4605), .A(n4539), .ZN(U3513) );
  MUX2_X1 U5104 ( .A(n4542), .B(n4541), .S(n4789), .Z(n4543) );
  OAI21_X1 U5105 ( .B1(n4544), .B2(n4605), .A(n4543), .ZN(U3512) );
  INV_X1 U5106 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4546) );
  MUX2_X1 U5107 ( .A(n4546), .B(n4545), .S(n4789), .Z(n4547) );
  OAI21_X1 U5108 ( .B1(n4548), .B2(n4605), .A(n4547), .ZN(U3511) );
  INV_X1 U5109 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4550) );
  MUX2_X1 U5110 ( .A(n4550), .B(n4549), .S(n4789), .Z(n4551) );
  OAI21_X1 U5111 ( .B1(n4552), .B2(n4605), .A(n4551), .ZN(U3510) );
  INV_X1 U5112 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4554) );
  MUX2_X1 U5113 ( .A(n4554), .B(n4553), .S(n4789), .Z(n4555) );
  OAI21_X1 U5114 ( .B1(n4556), .B2(n4605), .A(n4555), .ZN(U3509) );
  MUX2_X1 U5115 ( .A(REG0_REG_22__SCAN_IN), .B(n4557), .S(n4789), .Z(n4558) );
  INV_X1 U5116 ( .A(n4558), .ZN(n4559) );
  OAI21_X1 U5117 ( .B1(n4560), .B2(n4605), .A(n4559), .ZN(U3508) );
  INV_X1 U5118 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4562) );
  MUX2_X1 U5119 ( .A(n4562), .B(n4561), .S(n4789), .Z(n4563) );
  OAI21_X1 U5120 ( .B1(n4564), .B2(n4605), .A(n4563), .ZN(U3507) );
  INV_X1 U5121 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4566) );
  MUX2_X1 U5122 ( .A(n4566), .B(n4565), .S(n4789), .Z(n4567) );
  OAI21_X1 U5123 ( .B1(n4568), .B2(n4605), .A(n4567), .ZN(U3506) );
  INV_X1 U5124 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4570) );
  MUX2_X1 U5125 ( .A(n4570), .B(n4569), .S(n4789), .Z(n4571) );
  OAI21_X1 U5126 ( .B1(n4572), .B2(n4605), .A(n4571), .ZN(U3505) );
  MUX2_X1 U5127 ( .A(REG0_REG_18__SCAN_IN), .B(n4573), .S(n4789), .Z(U3503) );
  INV_X1 U5128 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4574) );
  MUX2_X1 U5129 ( .A(n4575), .B(n4574), .S(n4787), .Z(n4576) );
  OAI21_X1 U5130 ( .B1(n4577), .B2(n4605), .A(n4576), .ZN(U3501) );
  MUX2_X1 U5131 ( .A(REG0_REG_16__SCAN_IN), .B(n4578), .S(n4789), .Z(n4579) );
  AOI21_X1 U5132 ( .B1(n4580), .B2(n4595), .A(n4579), .ZN(n4581) );
  INV_X1 U5133 ( .A(n4581), .ZN(U3499) );
  INV_X1 U5134 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4582) );
  MUX2_X1 U5135 ( .A(n4583), .B(n4582), .S(n4787), .Z(n4584) );
  OAI21_X1 U5136 ( .B1(n4585), .B2(n4605), .A(n4584), .ZN(U3497) );
  INV_X1 U5137 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4587) );
  MUX2_X1 U5138 ( .A(n4587), .B(n4586), .S(n4789), .Z(n4588) );
  OAI21_X1 U5139 ( .B1(n4589), .B2(n4605), .A(n4588), .ZN(U3495) );
  MUX2_X1 U5140 ( .A(n3839), .B(n4590), .S(n4789), .Z(n4591) );
  OAI21_X1 U5141 ( .B1(n4592), .B2(n4605), .A(n4591), .ZN(U3493) );
  MUX2_X1 U5142 ( .A(REG0_REG_12__SCAN_IN), .B(n4593), .S(n4789), .Z(n4594) );
  AOI21_X1 U5143 ( .B1(n4596), .B2(n4595), .A(n4594), .ZN(n4597) );
  INV_X1 U5144 ( .A(n4597), .ZN(U3491) );
  MUX2_X1 U5145 ( .A(n4598), .B(REG0_REG_11__SCAN_IN), .S(n4787), .Z(n4599) );
  INV_X1 U5146 ( .A(n4599), .ZN(n4600) );
  OAI21_X1 U5147 ( .B1(n4601), .B2(n4605), .A(n4600), .ZN(U3489) );
  INV_X1 U5148 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4603) );
  MUX2_X1 U5149 ( .A(n4603), .B(n4602), .S(n4789), .Z(n4604) );
  OAI21_X1 U5150 ( .B1(n4724), .B2(n4605), .A(n4604), .ZN(U3483) );
  MUX2_X1 U5151 ( .A(n4606), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U5152 ( .A(n4607), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5153 ( .A(n4608), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U5154 ( .A(n4609), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U5155 ( .A(DATAI_20_), .B(n4610), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5156 ( .A(n4611), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5157 ( .A(DATAI_14_), .B(n4612), .S(STATE_REG_SCAN_IN), .Z(U3338)
         );
  MUX2_X1 U5158 ( .A(n4613), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5159 ( .A(DATAI_4_), .B(n4614), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5160 ( .A(n4615), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  INV_X1 U5161 ( .A(DATAI_28_), .ZN(n4616) );
  AOI22_X1 U5162 ( .A1(STATE_REG_SCAN_IN), .A2(n4617), .B1(n4616), .B2(U3149), 
        .ZN(U3324) );
  AOI22_X1 U5163 ( .A1(n4618), .A2(n4738), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4744), .ZN(n4619) );
  OAI21_X1 U5164 ( .B1(n4744), .B2(n4620), .A(n4619), .ZN(U3261) );
  OAI211_X1 U5165 ( .C1(n4623), .C2(n4622), .A(n4713), .B(n4621), .ZN(n4628)
         );
  OAI211_X1 U5166 ( .C1(n4626), .C2(n4625), .A(n4666), .B(n4624), .ZN(n4627)
         );
  OAI211_X1 U5167 ( .C1(n4718), .C2(n4766), .A(n4628), .B(n4627), .ZN(n4629)
         );
  AOI211_X1 U5168 ( .C1(n4711), .C2(ADDR_REG_9__SCAN_IN), .A(n4630), .B(n4629), 
        .ZN(n4631) );
  INV_X1 U5169 ( .A(n4631), .ZN(U3249) );
  OAI211_X1 U5170 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4634), .A(n4666), .B(n4633), .ZN(n4636) );
  NAND2_X1 U5171 ( .A1(n4636), .A2(n4635), .ZN(n4637) );
  AOI21_X1 U5172 ( .B1(n4711), .B2(ADDR_REG_10__SCAN_IN), .A(n4637), .ZN(n4641) );
  OAI211_X1 U5173 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4639), .A(n4713), .B(n4638), .ZN(n4640) );
  OAI211_X1 U5174 ( .C1(n4718), .C2(n2150), .A(n4641), .B(n4640), .ZN(U3250)
         );
  OAI211_X1 U5175 ( .C1(n4644), .C2(n4643), .A(n4713), .B(n4642), .ZN(n4649)
         );
  OAI211_X1 U5176 ( .C1(n4647), .C2(n4646), .A(n4666), .B(n4645), .ZN(n4648)
         );
  OAI211_X1 U5177 ( .C1(n4718), .C2(n4650), .A(n4649), .B(n4648), .ZN(n4651)
         );
  AOI211_X1 U5178 ( .C1(n4711), .C2(ADDR_REG_11__SCAN_IN), .A(n4652), .B(n4651), .ZN(n4653) );
  INV_X1 U5179 ( .A(n4653), .ZN(U3251) );
  OAI211_X1 U5180 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4656), .A(n4666), .B(n4655), .ZN(n4658) );
  NAND2_X1 U5181 ( .A1(n4658), .A2(n4657), .ZN(n4659) );
  AOI21_X1 U5182 ( .B1(n4711), .B2(ADDR_REG_12__SCAN_IN), .A(n4659), .ZN(n4663) );
  OAI211_X1 U5183 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4661), .A(n4713), .B(n4660), .ZN(n4662) );
  OAI211_X1 U5184 ( .C1(n4718), .C2(n2151), .A(n4663), .B(n4662), .ZN(U3252)
         );
  AOI21_X1 U5185 ( .B1(n4665), .B2(n4677), .A(n4664), .ZN(n4669) );
  OAI21_X1 U5186 ( .B1(n4669), .B2(n4668), .A(n4666), .ZN(n4667) );
  AOI21_X1 U5187 ( .B1(n4669), .B2(n4668), .A(n4667), .ZN(n4671) );
  AOI211_X1 U5188 ( .C1(n4711), .C2(ADDR_REG_13__SCAN_IN), .A(n4671), .B(n4670), .ZN(n4676) );
  OAI211_X1 U5189 ( .C1(n4674), .C2(n4673), .A(n4713), .B(n4672), .ZN(n4675)
         );
  OAI211_X1 U5190 ( .C1(n4718), .C2(n4677), .A(n4676), .B(n4675), .ZN(U3253)
         );
  AOI211_X1 U5191 ( .C1(n4680), .C2(n4679), .A(n4678), .B(n4707), .ZN(n4681)
         );
  AOI211_X1 U5192 ( .C1(n4711), .C2(ADDR_REG_15__SCAN_IN), .A(n4682), .B(n4681), .ZN(n4687) );
  OAI211_X1 U5193 ( .C1(n4685), .C2(n4684), .A(n4713), .B(n4683), .ZN(n4686)
         );
  OAI211_X1 U5194 ( .C1(n4718), .C2(n4758), .A(n4687), .B(n4686), .ZN(U3255)
         );
  AOI221_X1 U5195 ( .B1(n4690), .B2(n4689), .C1(n4688), .C2(n4689), .A(n4707), 
        .ZN(n4691) );
  AOI211_X1 U5196 ( .C1(n4711), .C2(ADDR_REG_16__SCAN_IN), .A(n4692), .B(n4691), .ZN(n4696) );
  OAI221_X1 U5197 ( .B1(n4694), .B2(REG1_REG_16__SCAN_IN), .C1(n4694), .C2(
        n4693), .A(n4713), .ZN(n4695) );
  OAI211_X1 U5198 ( .C1(n4718), .C2(n4756), .A(n4696), .B(n4695), .ZN(U3256)
         );
  AOI221_X1 U5199 ( .B1(n4699), .B2(n4698), .C1(n4697), .C2(n4698), .A(n4707), 
        .ZN(n4700) );
  AOI211_X1 U5200 ( .C1(n4711), .C2(ADDR_REG_17__SCAN_IN), .A(n4701), .B(n4700), .ZN(n4706) );
  OAI221_X1 U5201 ( .B1(n4704), .B2(n4703), .C1(n4704), .C2(n4702), .A(n4713), 
        .ZN(n4705) );
  OAI211_X1 U5202 ( .C1(n4718), .C2(n4754), .A(n4706), .B(n4705), .ZN(U3257)
         );
  OAI211_X1 U5203 ( .C1(n4715), .C2(n4714), .A(n4713), .B(n4712), .ZN(n4716)
         );
  OAI211_X1 U5204 ( .C1(n4718), .C2(n4753), .A(n4717), .B(n4716), .ZN(U3258)
         );
  OAI22_X1 U5205 ( .A1(n4722), .A2(n4721), .B1(n4720), .B2(n4719), .ZN(n4723)
         );
  INV_X1 U5206 ( .A(n4723), .ZN(n4728) );
  INV_X1 U5207 ( .A(n4724), .ZN(n4725) );
  AOI22_X1 U5208 ( .A1(n4726), .A2(n4739), .B1(n4738), .B2(n4725), .ZN(n4727)
         );
  OAI211_X1 U5209 ( .C1(n4744), .C2(n4729), .A(n4728), .B(n4727), .ZN(U3282)
         );
  AOI22_X1 U5210 ( .A1(n4744), .A2(REG2_REG_3__SCAN_IN), .B1(n4736), .B2(n4730), .ZN(n4734) );
  AOI22_X1 U5211 ( .A1(n4732), .A2(n4739), .B1(n4738), .B2(n4731), .ZN(n4733)
         );
  OAI211_X1 U5212 ( .C1(n4744), .C2(n4735), .A(n4734), .B(n4733), .ZN(U3287)
         );
  AOI22_X1 U5213 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4744), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4736), .ZN(n4742) );
  AOI22_X1 U5214 ( .A1(n4740), .A2(n4739), .B1(n4738), .B2(n4737), .ZN(n4741)
         );
  OAI211_X1 U5215 ( .C1(n4744), .C2(n4743), .A(n4742), .B(n4741), .ZN(U3288)
         );
  INV_X1 U5216 ( .A(n4749), .ZN(n4748) );
  NOR2_X1 U5217 ( .A1(n4748), .A2(n4745), .ZN(U3291) );
  AND2_X1 U5218 ( .A1(D_REG_30__SCAN_IN), .A2(n4749), .ZN(U3292) );
  AND2_X1 U5219 ( .A1(D_REG_29__SCAN_IN), .A2(n4749), .ZN(U3293) );
  AND2_X1 U5220 ( .A1(D_REG_28__SCAN_IN), .A2(n4749), .ZN(U3294) );
  AND2_X1 U5221 ( .A1(n4749), .A2(D_REG_27__SCAN_IN), .ZN(U3295) );
  AND2_X1 U5222 ( .A1(D_REG_26__SCAN_IN), .A2(n4749), .ZN(U3296) );
  NOR2_X1 U5223 ( .A1(n4748), .A2(n4746), .ZN(U3297) );
  AND2_X1 U5224 ( .A1(D_REG_24__SCAN_IN), .A2(n4749), .ZN(U3298) );
  AND2_X1 U5225 ( .A1(D_REG_23__SCAN_IN), .A2(n4749), .ZN(U3299) );
  AND2_X1 U5226 ( .A1(D_REG_22__SCAN_IN), .A2(n4749), .ZN(U3300) );
  AND2_X1 U5227 ( .A1(D_REG_21__SCAN_IN), .A2(n4749), .ZN(U3301) );
  AND2_X1 U5228 ( .A1(D_REG_20__SCAN_IN), .A2(n4749), .ZN(U3302) );
  AND2_X1 U5229 ( .A1(D_REG_19__SCAN_IN), .A2(n4749), .ZN(U3303) );
  AND2_X1 U5230 ( .A1(D_REG_18__SCAN_IN), .A2(n4749), .ZN(U3304) );
  AND2_X1 U5231 ( .A1(D_REG_17__SCAN_IN), .A2(n4749), .ZN(U3305) );
  AND2_X1 U5232 ( .A1(D_REG_16__SCAN_IN), .A2(n4749), .ZN(U3306) );
  AND2_X1 U5233 ( .A1(D_REG_15__SCAN_IN), .A2(n4749), .ZN(U3307) );
  AND2_X1 U5234 ( .A1(n4749), .A2(D_REG_14__SCAN_IN), .ZN(U3308) );
  AND2_X1 U5235 ( .A1(D_REG_13__SCAN_IN), .A2(n4749), .ZN(U3309) );
  AND2_X1 U5236 ( .A1(D_REG_12__SCAN_IN), .A2(n4749), .ZN(U3310) );
  AND2_X1 U5237 ( .A1(D_REG_11__SCAN_IN), .A2(n4749), .ZN(U3311) );
  AND2_X1 U5238 ( .A1(D_REG_10__SCAN_IN), .A2(n4749), .ZN(U3312) );
  AND2_X1 U5239 ( .A1(n4749), .A2(D_REG_9__SCAN_IN), .ZN(U3313) );
  AND2_X1 U5240 ( .A1(D_REG_8__SCAN_IN), .A2(n4749), .ZN(U3314) );
  AND2_X1 U5241 ( .A1(D_REG_7__SCAN_IN), .A2(n4749), .ZN(U3315) );
  AND2_X1 U5242 ( .A1(D_REG_6__SCAN_IN), .A2(n4749), .ZN(U3316) );
  AND2_X1 U5243 ( .A1(D_REG_5__SCAN_IN), .A2(n4749), .ZN(U3317) );
  AND2_X1 U5244 ( .A1(D_REG_4__SCAN_IN), .A2(n4749), .ZN(U3318) );
  NOR2_X1 U5245 ( .A1(n4748), .A2(n4747), .ZN(U3319) );
  AND2_X1 U5246 ( .A1(D_REG_2__SCAN_IN), .A2(n4749), .ZN(U3320) );
  INV_X1 U5247 ( .A(DATAI_23_), .ZN(n4751) );
  AOI21_X1 U5248 ( .B1(U3149), .B2(n4751), .A(n4750), .ZN(U3329) );
  INV_X1 U5249 ( .A(DATAI_18_), .ZN(n4752) );
  AOI22_X1 U5250 ( .A1(STATE_REG_SCAN_IN), .A2(n4753), .B1(n4752), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5251 ( .A1(STATE_REG_SCAN_IN), .A2(n4754), .B1(n2478), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5252 ( .A(DATAI_16_), .ZN(n4755) );
  AOI22_X1 U5253 ( .A1(STATE_REG_SCAN_IN), .A2(n4756), .B1(n4755), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5254 ( .A(DATAI_15_), .ZN(n4757) );
  AOI22_X1 U5255 ( .A1(STATE_REG_SCAN_IN), .A2(n4758), .B1(n4757), .B2(U3149), 
        .ZN(U3337) );
  OAI22_X1 U5256 ( .A1(U3149), .A2(n4759), .B1(DATAI_13_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4760) );
  INV_X1 U5257 ( .A(n4760), .ZN(U3339) );
  INV_X1 U5258 ( .A(DATAI_12_), .ZN(n4761) );
  AOI22_X1 U5259 ( .A1(STATE_REG_SCAN_IN), .A2(n2151), .B1(n4761), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U5260 ( .A1(U3149), .A2(n4762), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4763) );
  INV_X1 U5261 ( .A(n4763), .ZN(U3341) );
  INV_X1 U5262 ( .A(DATAI_10_), .ZN(n4764) );
  AOI22_X1 U5263 ( .A1(STATE_REG_SCAN_IN), .A2(n2150), .B1(n4764), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5264 ( .A(DATAI_9_), .ZN(n4765) );
  AOI22_X1 U5265 ( .A1(STATE_REG_SCAN_IN), .A2(n4766), .B1(n4765), .B2(U3149), 
        .ZN(U3343) );
  INV_X1 U5266 ( .A(DATAI_0_), .ZN(n4768) );
  AOI22_X1 U5267 ( .A1(STATE_REG_SCAN_IN), .A2(n4769), .B1(n4768), .B2(U3149), 
        .ZN(U3352) );
  INV_X1 U5268 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4770) );
  AOI22_X1 U5269 ( .A1(n4789), .A2(n4771), .B1(n4770), .B2(n4787), .ZN(U3467)
         );
  INV_X1 U5270 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4772) );
  AOI22_X1 U5271 ( .A1(n4789), .A2(n4773), .B1(n4772), .B2(n4787), .ZN(U3469)
         );
  INV_X1 U5272 ( .A(n4774), .ZN(n4779) );
  INV_X1 U5273 ( .A(n4775), .ZN(n4777) );
  AOI211_X1 U5274 ( .C1(n4779), .C2(n4778), .A(n4777), .B(n4776), .ZN(n4791)
         );
  INV_X1 U5275 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4780) );
  AOI22_X1 U5276 ( .A1(n4789), .A2(n4791), .B1(n4780), .B2(n4787), .ZN(U3475)
         );
  NOR2_X1 U5277 ( .A1(n4782), .A2(n4781), .ZN(n4786) );
  AOI211_X1 U5278 ( .C1(n4786), .C2(n4785), .A(n4784), .B(n4783), .ZN(n4794)
         );
  AOI22_X1 U5279 ( .A1(n4789), .A2(n4794), .B1(n4788), .B2(n4787), .ZN(U3481)
         );
  AOI22_X1 U5280 ( .A1(n4795), .A2(n4791), .B1(n4790), .B2(n4792), .ZN(U3522)
         );
  AOI22_X1 U5281 ( .A1(n4795), .A2(n4794), .B1(n4793), .B2(n4792), .ZN(U3525)
         );
endmodule

