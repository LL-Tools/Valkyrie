

module b15_C_gen_AntiSAT_k_128_10 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, 
        U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, 
        U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, 
        U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, 
        U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, 
        U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, 
        U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, 
        U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, 
        U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, 
        U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, 
        U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, 
        U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, 
        U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, 
        U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, 
        U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, 
        U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, 
        U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, 
        U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, 
        U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, 
        U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, 
        U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, 
        U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, 
        U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, 
        U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, 
        U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, 
        U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, 
        U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, 
        U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, 
        U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, 
        U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, 
        U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, 
        U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, 
        U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, 
        U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, 
        U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, 
        U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, 
        U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, 
        U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, 
        U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, 
        U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, 
        U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, 
        U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, 
        U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, 
        U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, 
        U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, 
        U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1,
         keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6,
         keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11,
         keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16,
         keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21,
         keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26,
         keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31,
         keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36,
         keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41,
         keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46,
         keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51,
         keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56,
         keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61,
         keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791;

  XNOR2_X1 U3431 ( .A(n4112), .B(n4111), .ZN(n5528) );
  XNOR2_X1 U3432 ( .A(n5366), .B(n5365), .ZN(n5374) );
  INV_X1 U3433 ( .A(n2984), .ZN(n5440) );
  INV_X2 U3434 ( .A(n6175), .ZN(n6162) );
  NAND2_X1 U3435 ( .A1(n3533), .A2(n3078), .ZN(n3535) );
  BUF_X1 U3436 ( .A(n4401), .Z(n3021) );
  CLKBUF_X2 U3437 ( .A(n4504), .Z(n3029) );
  INV_X1 U3438 ( .A(n5097), .ZN(n3419) );
  CLKBUF_X2 U3439 ( .A(n2990), .Z(n2991) );
  NAND2_X1 U3440 ( .A1(n3325), .A2(n3324), .ZN(n3326) );
  CLKBUF_X2 U3441 ( .A(n3335), .Z(n4084) );
  NAND2_X1 U3442 ( .A1(n3240), .A2(n3239), .ZN(n4124) );
  CLKBUF_X2 U3443 ( .A(n3333), .Z(n3334) );
  CLKBUF_X2 U3444 ( .A(n3269), .Z(n4091) );
  CLKBUF_X2 U34450 ( .A(n3026), .Z(n3022) );
  CLKBUF_X2 U34460 ( .A(n3185), .Z(n3027) );
  CLKBUF_X2 U34470 ( .A(n3328), .Z(n4062) );
  CLKBUF_X1 U3449 ( .A(n3211), .Z(n4529) );
  INV_X1 U3450 ( .A(n4268), .ZN(n4525) );
  NAND4_X2 U34510 ( .A1(n3209), .A2(n3208), .A3(n3207), .A4(n3206), .ZN(n4145)
         );
  AND2_X1 U34520 ( .A1(n3137), .A2(n3136), .ZN(n3211) );
  AND4_X1 U34530 ( .A1(n3115), .A2(n3114), .A3(n3113), .A4(n3112), .ZN(n3116)
         );
  AND2_X2 U3454 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4471) );
  AND2_X2 U34550 ( .A1(n3359), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4391) );
  INV_X1 U34560 ( .A(n5782), .ZN(n2983) );
  XNOR2_X1 U3457 ( .A(n3292), .B(n3291), .ZN(n4370) );
  CLKBUF_X1 U34590 ( .A(n4722), .Z(n2985) );
  CLKBUF_X1 U34600 ( .A(n5250), .Z(n2986) );
  CLKBUF_X1 U34610 ( .A(n5195), .Z(n2987) );
  XNOR2_X1 U34630 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3580) );
  XNOR2_X1 U34640 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3560) );
  AND2_X2 U34650 ( .A1(n4375), .A2(n3100), .ZN(n3201) );
  AND2_X1 U3466 ( .A1(n3099), .A2(n4471), .ZN(n3335) );
  INV_X1 U34680 ( .A(n4251), .ZN(n5471) );
  AND2_X1 U34690 ( .A1(n4418), .A2(n4419), .ZN(n4416) );
  NAND2_X1 U34700 ( .A1(n4525), .A2(n2993), .ZN(n3545) );
  INV_X1 U34710 ( .A(n6022), .ZN(n5993) );
  AND2_X2 U34720 ( .A1(n4391), .A2(n3099), .ZN(n3185) );
  AND4_X1 U34730 ( .A1(n3168), .A2(n3167), .A3(n3166), .A4(n3165), .ZN(n2989)
         );
  XNOR2_X1 U34740 ( .A(n3439), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4439)
         );
  AND2_X1 U3475 ( .A1(n4445), .A2(n3426), .ZN(n6157) );
  AND2_X1 U3478 ( .A1(n4754), .A2(n3715), .ZN(n4906) );
  CLKBUF_X2 U3479 ( .A(n6088), .Z(n6152) );
  AND2_X1 U3480 ( .A1(n4574), .A2(n3041), .ZN(n4494) );
  AND2_X1 U3481 ( .A1(n3284), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3569) );
  CLKBUF_X2 U3482 ( .A(n3370), .Z(n3307) );
  BUF_X2 U3483 ( .A(n3196), .Z(n3721) );
  CLKBUF_X1 U3485 ( .A(n3293), .Z(n2990) );
  BUF_X2 U3486 ( .A(n3174), .Z(n4067) );
  NOR2_X1 U3487 ( .A1(n5372), .A2(n5371), .ZN(n5373) );
  AOI22_X1 U3488 ( .A1(n5752), .A2(n5572), .B1(n5621), .B2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5611) );
  AND2_X1 U3489 ( .A1(n5481), .A2(n5480), .ZN(n5838) );
  AND2_X1 U3490 ( .A1(n5562), .A2(n5478), .ZN(n5841) );
  CLKBUF_X1 U3491 ( .A(n5413), .Z(n5414) );
  NAND2_X1 U3492 ( .A1(n5637), .A2(n5638), .ZN(n5620) );
  NAND2_X1 U3493 ( .A1(n3506), .A2(n3002), .ZN(n2999) );
  BUF_X1 U3494 ( .A(n5214), .Z(n2998) );
  NAND2_X1 U3495 ( .A1(n3497), .A2(n3496), .ZN(n5195) );
  NAND3_X1 U3496 ( .A1(n3733), .A2(n3035), .A3(n4906), .ZN(n3769) );
  NAND2_X1 U3497 ( .A1(n3667), .A2(n3094), .ZN(n4754) );
  XNOR2_X1 U3498 ( .A(n3514), .B(n4182), .ZN(n4961) );
  NAND2_X1 U3499 ( .A1(n5621), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3522) );
  INV_X2 U3500 ( .A(n5621), .ZN(n2992) );
  NAND2_X1 U3501 ( .A1(n3518), .A2(n3513), .ZN(n3514) );
  XNOR2_X1 U3502 ( .A(n3507), .B(n3500), .ZN(n3662) );
  NAND2_X2 U3503 ( .A1(n3507), .A2(n3509), .ZN(n3518) );
  OAI21_X1 U3504 ( .B1(n3646), .B2(n3788), .A(n3652), .ZN(n4560) );
  OAI21_X1 U3505 ( .B1(n3646), .B2(n3467), .A(n3466), .ZN(n3469) );
  NAND2_X1 U3506 ( .A1(n3460), .A2(n3459), .ZN(n3488) );
  OR2_X1 U3507 ( .A1(n3460), .A2(n3459), .ZN(n3461) );
  XNOR2_X1 U3508 ( .A(n3446), .B(n3444), .ZN(n3637) );
  NAND2_X1 U3509 ( .A1(n3380), .A2(n4503), .ZN(n3446) );
  XNOR2_X1 U3510 ( .A(n3425), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4447)
         );
  OR2_X2 U3511 ( .A1(n6156), .A2(n6170), .ZN(n6166) );
  NOR2_X1 U3512 ( .A1(n4555), .A2(n5527), .ZN(n6443) );
  XNOR2_X1 U3513 ( .A(n3288), .B(n3287), .ZN(n3428) );
  CLKBUF_X1 U3514 ( .A(n4382), .Z(n6277) );
  NAND2_X1 U3515 ( .A1(n3305), .A2(n3304), .ZN(n3407) );
  NAND2_X2 U3516 ( .A1(n6071), .A2(n6473), .ZN(n5914) );
  NAND2_X1 U3517 ( .A1(n3283), .A2(n3282), .ZN(n3288) );
  AND2_X1 U3518 ( .A1(n3805), .A2(n3064), .ZN(n3063) );
  NAND2_X1 U3519 ( .A1(n3267), .A2(n3266), .ZN(n3357) );
  NAND2_X1 U3520 ( .A1(n3322), .A2(n3323), .ZN(n3327) );
  NAND2_X1 U3521 ( .A1(n3226), .A2(n3225), .ZN(n3322) );
  AND2_X1 U3522 ( .A1(n3257), .A2(n3256), .ZN(n3258) );
  NOR2_X1 U3523 ( .A1(n3224), .A2(n3223), .ZN(n3225) );
  NAND2_X1 U3524 ( .A1(n3172), .A2(n3171), .ZN(n3243) );
  AND2_X1 U3525 ( .A1(n3415), .A2(n3345), .ZN(n3346) );
  OR2_X1 U3526 ( .A1(n3342), .A2(n3343), .ZN(n3415) );
  OR2_X1 U3527 ( .A1(n4251), .A2(n3610), .ZN(n4371) );
  NOR2_X1 U3528 ( .A1(n4150), .A2(n6490), .ZN(n3508) );
  INV_X1 U3529 ( .A(n3211), .ZN(n4150) );
  AND2_X1 U3530 ( .A1(n3546), .A2(n4268), .ZN(n3550) );
  OR2_X1 U3531 ( .A1(n3303), .A2(n3302), .ZN(n3409) );
  OR2_X1 U3532 ( .A1(n3341), .A2(n3340), .ZN(n3421) );
  AND2_X1 U3533 ( .A1(n4554), .A2(n3219), .ZN(n3616) );
  NAND2_X1 U3534 ( .A1(n3219), .A2(n3611), .ZN(n4271) );
  NAND2_X2 U3535 ( .A1(n3032), .A2(n2989), .ZN(n3420) );
  INV_X1 U3536 ( .A(n3170), .ZN(n3160) );
  INV_X1 U3537 ( .A(n4145), .ZN(n2993) );
  AND4_X2 U3538 ( .A1(n3157), .A2(n3156), .A3(n3155), .A4(n3154), .ZN(n4537)
         );
  AND4_X1 U3539 ( .A1(n3131), .A2(n3130), .A3(n3129), .A4(n3128), .ZN(n3137)
         );
  AND4_X1 U3540 ( .A1(n3190), .A2(n3189), .A3(n3188), .A4(n3187), .ZN(n3209)
         );
  AND4_X1 U3541 ( .A1(n3195), .A2(n3194), .A3(n3193), .A4(n3192), .ZN(n3208)
         );
  NAND2_X2 U3542 ( .A1(n3117), .A2(n3116), .ZN(n3611) );
  OR2_X2 U3543 ( .A1(n3107), .A2(n3106), .ZN(n3219) );
  AND4_X1 U3544 ( .A1(n3145), .A2(n3144), .A3(n3143), .A4(n3142), .ZN(n3156)
         );
  AND4_X1 U3545 ( .A1(n3111), .A2(n3110), .A3(n3109), .A4(n3108), .ZN(n3117)
         );
  AND4_X1 U3546 ( .A1(n3164), .A2(n3163), .A3(n3162), .A4(n3161), .ZN(n3032)
         );
  AND4_X1 U3547 ( .A1(n3153), .A2(n3152), .A3(n3151), .A4(n3150), .ZN(n3154)
         );
  AND4_X1 U3548 ( .A1(n3149), .A2(n3148), .A3(n3147), .A4(n3146), .ZN(n3155)
         );
  AND4_X1 U3549 ( .A1(n3141), .A2(n3140), .A3(n3139), .A4(n3138), .ZN(n3157)
         );
  INV_X2 U3550 ( .A(n4388), .ZN(n4090) );
  AND4_X1 U3551 ( .A1(n3178), .A2(n3177), .A3(n3176), .A4(n3175), .ZN(n3183)
         );
  AND4_X1 U3552 ( .A1(n3121), .A2(n3120), .A3(n3119), .A4(n3118), .ZN(n3127)
         );
  AND4_X1 U3553 ( .A1(n3205), .A2(n3204), .A3(n3203), .A4(n3202), .ZN(n3206)
         );
  AND4_X1 U3554 ( .A1(n3135), .A2(n3134), .A3(n3133), .A4(n3132), .ZN(n3136)
         );
  BUF_X2 U3555 ( .A(n3186), .Z(n4085) );
  BUF_X2 U3556 ( .A(n3191), .Z(n4092) );
  AND2_X2 U3557 ( .A1(n4385), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4392)
         );
  CLKBUF_X1 U3558 ( .A(n6157), .Z(n2994) );
  AND2_X2 U3559 ( .A1(n2999), .A2(n3000), .ZN(n2995) );
  OR2_X1 U3560 ( .A1(n3001), .A2(n3005), .ZN(n3000) );
  NAND2_X1 U3561 ( .A1(n2999), .A2(n3000), .ZN(n5165) );
  INV_X2 U3562 ( .A(n5577), .ZN(n5604) );
  NAND2_X2 U3563 ( .A1(n3486), .A2(n3485), .ZN(n3507) );
  NAND2_X1 U3564 ( .A1(n3772), .A2(n3771), .ZN(n2996) );
  AND2_X2 U3565 ( .A1(n2996), .A2(n2997), .ZN(n5266) );
  AND2_X1 U3566 ( .A1(n3063), .A2(n5185), .ZN(n2997) );
  INV_X1 U3567 ( .A(n3003), .ZN(n3001) );
  AND2_X1 U3568 ( .A1(n3505), .A2(n3003), .ZN(n3002) );
  OR2_X1 U3569 ( .A1(n3004), .A2(n3076), .ZN(n3003) );
  INV_X1 U3570 ( .A(n3516), .ZN(n3004) );
  AND2_X1 U3571 ( .A1(n4961), .A2(n3516), .ZN(n3005) );
  INV_X1 U3572 ( .A(n5343), .ZN(n3006) );
  CLKBUF_X1 U3573 ( .A(n4446), .Z(n3007) );
  NAND2_X1 U3574 ( .A1(n3413), .A2(n3412), .ZN(n4446) );
  NOR2_X2 U3575 ( .A1(n5478), .A2(n5479), .ZN(n5315) );
  NAND2_X1 U3576 ( .A1(n3524), .A2(n3011), .ZN(n3008) );
  AND2_X2 U3577 ( .A1(n3008), .A2(n3009), .ZN(n5618) );
  OR2_X1 U3578 ( .A1(n3010), .A2(n5638), .ZN(n3009) );
  INV_X1 U3579 ( .A(n3074), .ZN(n3010) );
  AND2_X1 U3580 ( .A1(n3523), .A2(n3074), .ZN(n3011) );
  CLKBUF_X1 U3581 ( .A(n4445), .Z(n3012) );
  CLKBUF_X1 U3582 ( .A(n5296), .Z(n3013) );
  AND2_X2 U3583 ( .A1(n3535), .A2(n3534), .ZN(n3014) );
  AND2_X4 U3584 ( .A1(n4392), .A2(n4375), .ZN(n3333) );
  AND2_X1 U3585 ( .A1(n3099), .A2(n4392), .ZN(n3015) );
  AND2_X4 U3586 ( .A1(n4392), .A2(n3101), .ZN(n3328) );
  AND2_X2 U3587 ( .A1(n3100), .A2(n4374), .ZN(n3191) );
  AND2_X1 U3588 ( .A1(n4374), .A2(n4471), .ZN(n3309) );
  AND2_X2 U3589 ( .A1(n4375), .A2(n4471), .ZN(n3174) );
  AND2_X2 U3590 ( .A1(n4391), .A2(n4375), .ZN(n3269) );
  AND2_X1 U3591 ( .A1(n3099), .A2(n4471), .ZN(n3018) );
  AND2_X1 U3592 ( .A1(n4391), .A2(n3101), .ZN(n3268) );
  AND2_X1 U3593 ( .A1(n3101), .A2(n4471), .ZN(n3019) );
  AND2_X1 U3594 ( .A1(n4537), .A2(n3420), .ZN(n4269) );
  NAND2_X1 U3595 ( .A1(n3398), .A2(n3397), .ZN(n3441) );
  NAND2_X1 U3596 ( .A1(n3404), .A2(n3403), .ZN(n3439) );
  AOI21_X2 U3597 ( .B1(n5611), .B2(n5612), .A(n5574), .ZN(n5606) );
  NOR2_X2 U3598 ( .A1(n4461), .A2(n4462), .ZN(n4463) );
  NAND2_X1 U3599 ( .A1(n3351), .A2(n3414), .ZN(n3418) );
  NAND2_X2 U3600 ( .A1(n5585), .A2(n3528), .ZN(n5752) );
  NAND2_X2 U3601 ( .A1(n3127), .A2(n3126), .ZN(n3170) );
  XNOR2_X1 U3602 ( .A(n3428), .B(n3427), .ZN(n4502) );
  OAI21_X2 U3603 ( .B1(n4439), .B2(n4438), .A(n3440), .ZN(n4490) );
  AND2_X1 U3604 ( .A1(n4392), .A2(n4374), .ZN(n3020) );
  AND2_X2 U3605 ( .A1(n5453), .A2(n5454), .ZN(n5439) );
  NOR2_X2 U3606 ( .A1(n5465), .A2(n5512), .ZN(n5453) );
  INV_X2 U3607 ( .A(n3518), .ZN(n5621) );
  NAND2_X2 U3608 ( .A1(n3327), .A2(n3326), .ZN(n3617) );
  NAND2_X2 U3609 ( .A1(n5576), .A2(n5575), .ZN(n5577) );
  OR2_X2 U3611 ( .A1(n3218), .A2(n4533), .ZN(n3215) );
  XNOR2_X1 U3612 ( .A(n3356), .B(n3357), .ZN(n4401) );
  NOR2_X4 U3613 ( .A1(n5413), .A2(n5415), .ZN(n4308) );
  AND2_X4 U3614 ( .A1(n3099), .A2(n3100), .ZN(n3023) );
  AND2_X1 U3615 ( .A1(n3099), .A2(n3100), .ZN(n3274) );
  AND2_X1 U3616 ( .A1(n4374), .A2(n4471), .ZN(n3024) );
  AND2_X2 U3617 ( .A1(n4374), .A2(n4471), .ZN(n3025) );
  AND2_X1 U3618 ( .A1(n4392), .A2(n4374), .ZN(n3293) );
  AND2_X1 U3619 ( .A1(n4391), .A2(n3101), .ZN(n3026) );
  BUF_X1 U3620 ( .A(n4504), .Z(n3028) );
  XNOR2_X1 U3621 ( .A(n3408), .B(n3407), .ZN(n4504) );
  OR2_X1 U3622 ( .A1(n5407), .A2(n4369), .ZN(n4351) );
  NAND2_X1 U3623 ( .A1(n3508), .A2(n3499), .ZN(n3342) );
  OR2_X1 U3624 ( .A1(n3594), .A2(n3482), .ZN(n3483) );
  INV_X1 U3625 ( .A(n3444), .ZN(n3445) );
  OR2_X1 U3626 ( .A1(n3590), .A2(n6234), .ZN(n3592) );
  AOI21_X1 U3627 ( .B1(n3196), .B2(INSTQUEUE_REG_9__0__SCAN_IN), .A(n3200), 
        .ZN(n3207) );
  AND2_X1 U3628 ( .A1(n4525), .A2(n4145), .ZN(n3395) );
  AND2_X1 U3629 ( .A1(n5490), .A2(n4307), .ZN(n3061) );
  OR2_X2 U3630 ( .A1(n5683), .A2(n5682), .ZN(n3045) );
  NAND2_X1 U3631 ( .A1(n3259), .A2(n3258), .ZN(n3290) );
  NAND2_X1 U3632 ( .A1(n3254), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3259) );
  AOI22_X1 U3633 ( .A1(n3174), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3112) );
  INV_X1 U3634 ( .A(n4335), .ZN(n6580) );
  AND2_X1 U3635 ( .A1(n6585), .A2(n4318), .ZN(n5963) );
  NAND2_X1 U3636 ( .A1(n6071), .A2(n4424), .ZN(n6105) );
  NAND2_X1 U3637 ( .A1(n5484), .A2(n5318), .ZN(n5320) );
  OR2_X1 U3638 ( .A1(n3344), .A2(n6490), .ZN(n3345) );
  INV_X1 U3639 ( .A(n3394), .ZN(n3462) );
  INV_X1 U3640 ( .A(n3487), .ZN(n3485) );
  INV_X1 U3641 ( .A(n3488), .ZN(n3486) );
  NAND2_X1 U3642 ( .A1(n4150), .A2(n4145), .ZN(n3365) );
  OR2_X1 U3643 ( .A1(n3376), .A2(n3375), .ZN(n3400) );
  NAND2_X1 U3644 ( .A1(n3365), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3594) );
  BUF_X1 U3645 ( .A(n3611), .Z(n3612) );
  OR2_X1 U3646 ( .A1(n3698), .A2(n4947), .ZN(n3714) );
  INV_X1 U3647 ( .A(n3649), .ZN(n4105) );
  AND2_X1 U3648 ( .A1(n4227), .A2(n5472), .ZN(n4231) );
  NOR2_X1 U3649 ( .A1(n3050), .A2(n5287), .ZN(n3049) );
  INV_X1 U3650 ( .A(n5516), .ZN(n3050) );
  NAND2_X1 U3651 ( .A1(n3252), .A2(n3083), .ZN(n3289) );
  NAND2_X1 U3652 ( .A1(n3358), .A2(n3357), .ZN(n4478) );
  NAND2_X1 U3653 ( .A1(n3364), .A2(n3363), .ZN(n6282) );
  INV_X1 U3654 ( .A(n3029), .ZN(n4646) );
  NOR2_X1 U3655 ( .A1(n4373), .A2(n4278), .ZN(n5400) );
  NOR2_X1 U3656 ( .A1(n5965), .A2(n4325), .ZN(n5189) );
  INV_X1 U3657 ( .A(n5089), .ZN(n5347) );
  NAND2_X1 U3658 ( .A1(n5418), .A2(n3043), .ZN(n5683) );
  NOR2_X1 U3659 ( .A1(n4246), .A2(n5491), .ZN(n3043) );
  AOI21_X1 U3660 ( .B1(n4419), .B2(n3056), .A(n4109), .ZN(n3055) );
  INV_X1 U3661 ( .A(n4419), .ZN(n3058) );
  INV_X1 U3662 ( .A(n3615), .ZN(n3056) );
  NAND2_X1 U3663 ( .A1(n3038), .A2(n3245), .ZN(n4420) );
  NAND2_X1 U3664 ( .A1(n4058), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4117)
         );
  AND2_X1 U3665 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n4034), .ZN(n4035)
         );
  NAND2_X1 U3666 ( .A1(n4035), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4057)
         );
  AND2_X1 U3667 ( .A1(n3061), .A2(n5561), .ZN(n3060) );
  AND2_X1 U3668 ( .A1(n3835), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3836)
         );
  NAND2_X1 U3669 ( .A1(n3836), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3870)
         );
  NAND2_X1 U3670 ( .A1(n3059), .A2(n3615), .ZN(n4418) );
  NOR2_X1 U3671 ( .A1(n3080), .A2(n3079), .ZN(n3078) );
  INV_X1 U3672 ( .A(n3532), .ZN(n3079) );
  INV_X1 U3673 ( .A(n3033), .ZN(n3080) );
  AOI21_X1 U3674 ( .B1(n5241), .B2(n3071), .A(n3070), .ZN(n3069) );
  INV_X1 U3675 ( .A(n5242), .ZN(n3070) );
  AND2_X1 U3676 ( .A1(n4573), .A2(n3031), .ZN(n3041) );
  XNOR2_X1 U3677 ( .A(n4159), .B(n4563), .ZN(n4448) );
  OAI21_X1 U3678 ( .B1(n4351), .B2(n4143), .A(n4142), .ZN(n4285) );
  NAND2_X1 U3679 ( .A1(n3418), .A2(n3352), .ZN(n3406) );
  OAI211_X1 U3680 ( .C1(n3321), .C2(n3320), .A(n3319), .B(n3342), .ZN(n3405)
         );
  AND2_X1 U3681 ( .A1(n3029), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6368) );
  XNOR2_X1 U3682 ( .A(n4478), .B(n6282), .ZN(n4382) );
  INV_X1 U3683 ( .A(n4376), .ZN(n5334) );
  AND2_X1 U3684 ( .A1(n3604), .A2(n3603), .ZN(n5407) );
  NAND2_X1 U3685 ( .A1(n4507), .A2(n4647), .ZN(n6367) );
  NAND2_X1 U3686 ( .A1(n4646), .A2(n5097), .ZN(n4833) );
  INV_X1 U3687 ( .A(n4520), .ZN(n4837) );
  AND2_X1 U3688 ( .A1(n6493), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3605) );
  INV_X1 U3689 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6656) );
  NAND2_X1 U3690 ( .A1(n5388), .A2(n5387), .ZN(n5389) );
  NAND2_X1 U3691 ( .A1(n5383), .A2(REIP_REG_30__SCAN_IN), .ZN(n5388) );
  AND2_X1 U3692 ( .A1(n5386), .A2(n5385), .ZN(n5387) );
  AND3_X1 U3693 ( .A1(n5797), .A2(REIP_REG_28__SCAN_IN), .A3(
        REIP_REG_27__SCAN_IN), .ZN(n5392) );
  OR2_X1 U3694 ( .A1(n5963), .A2(n4319), .ZN(n5971) );
  OR2_X1 U3695 ( .A1(n5484), .A2(n5318), .ZN(n5319) );
  AND2_X1 U3696 ( .A1(n5526), .A2(n5376), .ZN(n6046) );
  INV_X1 U3697 ( .A(n5526), .ZN(n6045) );
  AND2_X1 U3698 ( .A1(n5526), .A2(n4427), .ZN(n5225) );
  INV_X1 U3699 ( .A(n6225), .ZN(n6210) );
  OR2_X1 U3700 ( .A1(n3281), .A2(n3280), .ZN(n3393) );
  AND2_X2 U3701 ( .A1(n3234), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3101)
         );
  OAI21_X1 U3702 ( .B1(n3611), .B2(n3211), .A(n4537), .ZN(n3158) );
  INV_X1 U3703 ( .A(n3542), .ZN(n3561) );
  NAND2_X1 U3704 ( .A1(n3392), .A2(n3391), .ZN(n3444) );
  NAND2_X1 U3705 ( .A1(n3458), .A2(n3457), .ZN(n3459) );
  OR2_X1 U3706 ( .A1(n3481), .A2(n3480), .ZN(n3491) );
  OR2_X1 U3707 ( .A1(n3456), .A2(n3455), .ZN(n3464) );
  NAND2_X1 U3708 ( .A1(n3214), .A2(n3219), .ZN(n3238) );
  INV_X1 U3709 ( .A(n3213), .ZN(n3214) );
  NAND2_X1 U3710 ( .A1(n3569), .A2(n3550), .ZN(n3600) );
  AOI22_X1 U3711 ( .A1(n3026), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3186), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3166) );
  AOI22_X1 U3712 ( .A1(n3328), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3185), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3125) );
  AOI22_X1 U3713 ( .A1(n3015), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3019), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3119) );
  AOI22_X1 U3714 ( .A1(n3020), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3186), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3120) );
  AOI22_X1 U3715 ( .A1(n3333), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3024), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3118) );
  AOI22_X1 U3716 ( .A1(n3328), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3268), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3111) );
  AOI22_X1 U3717 ( .A1(n3185), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3186), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3110) );
  AOI22_X1 U3718 ( .A1(n3020), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3109) );
  AOI22_X1 U3719 ( .A1(n3023), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3114) );
  AND2_X1 U3720 ( .A1(n4269), .A2(n3227), .ZN(n3239) );
  INV_X1 U3721 ( .A(n3238), .ZN(n3240) );
  NOR2_X1 U3722 ( .A1(n3213), .A2(n3616), .ZN(n3171) );
  AND2_X1 U3723 ( .A1(n3956), .A2(n3925), .ZN(n3065) );
  NAND2_X1 U3725 ( .A1(n3628), .A2(n3627), .ZN(n4455) );
  NAND2_X1 U3726 ( .A1(n3436), .A2(n3435), .ZN(n3437) );
  NOR2_X1 U3727 ( .A1(n3219), .A2(n6481), .ZN(n3623) );
  NAND2_X1 U3728 ( .A1(n3535), .A2(n3534), .ZN(n5360) );
  NAND2_X1 U3729 ( .A1(n2992), .A2(n5879), .ZN(n3534) );
  NAND2_X1 U3730 ( .A1(n5621), .A2(n3531), .ZN(n3532) );
  INV_X1 U3731 ( .A(n5605), .ZN(n5575) );
  NOR2_X1 U3732 ( .A1(n3075), .A2(n5629), .ZN(n3074) );
  INV_X1 U3733 ( .A(n3525), .ZN(n3075) );
  AND2_X1 U3734 ( .A1(n4998), .A2(n3036), .ZN(n4910) );
  INV_X1 U3735 ( .A(n4909), .ZN(n3046) );
  NOR2_X1 U3736 ( .A1(n3072), .A2(n3068), .ZN(n3067) );
  INV_X1 U3737 ( .A(n5241), .ZN(n3072) );
  INV_X1 U3738 ( .A(n3034), .ZN(n3068) );
  INV_X1 U3739 ( .A(n5166), .ZN(n3071) );
  INV_X1 U3740 ( .A(n4234), .ZN(n4254) );
  NAND2_X1 U3741 ( .A1(n4156), .A2(n3054), .ZN(n4159) );
  NAND2_X1 U3742 ( .A1(n4161), .A2(n4570), .ZN(n3054) );
  NAND2_X1 U3743 ( .A1(n6167), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3425)
         );
  INV_X1 U3744 ( .A(n3421), .ZN(n3343) );
  INV_X1 U3745 ( .A(n3510), .ZN(n3499) );
  OR3_X1 U3746 ( .A1(n4267), .A2(n4277), .A3(n4276), .ZN(n4373) );
  NAND2_X1 U3747 ( .A1(n3593), .A2(n3592), .ZN(n4138) );
  OAI21_X1 U3748 ( .B1(n4482), .B2(n4484), .A(n6483), .ZN(n4523) );
  NAND2_X1 U3749 ( .A1(n4382), .A2(n6490), .ZN(n3379) );
  NAND2_X1 U3750 ( .A1(n3241), .A2(n4145), .ZN(n5401) );
  AND2_X1 U3751 ( .A1(n3909), .A2(n3908), .ZN(n5441) );
  NOR2_X1 U3752 ( .A1(n5285), .A2(n4326), .ZN(n5821) );
  NOR2_X1 U3753 ( .A1(n3735), .A2(n3734), .ZN(n3753) );
  NAND2_X1 U3754 ( .A1(n5418), .A2(n4331), .ZN(n5492) );
  AND2_X1 U3755 ( .A1(n5430), .A2(n5416), .ZN(n5418) );
  NOR2_X1 U3756 ( .A1(n5504), .A2(n5431), .ZN(n5430) );
  AND2_X1 U3757 ( .A1(n5800), .A2(n4105), .ZN(n4014) );
  NOR2_X1 U3758 ( .A1(n4351), .A2(n4350), .ZN(n6049) );
  CLKBUF_X1 U3759 ( .A(n3395), .Z(n4335) );
  INV_X1 U3760 ( .A(n6480), .ZN(n6070) );
  AND2_X1 U3761 ( .A1(n4037), .A2(n4036), .ZN(n5561) );
  AND2_X1 U3762 ( .A1(n3997), .A2(n3996), .ZN(n4307) );
  NAND2_X1 U3763 ( .A1(n3993), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4033)
         );
  NOR2_X1 U3764 ( .A1(n3950), .A2(n5600), .ZN(n3951) );
  AND2_X1 U3765 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n3906), .ZN(n3907)
         );
  INV_X1 U3766 ( .A(n3905), .ZN(n3906) );
  NAND2_X1 U3767 ( .A1(n3907), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3950)
         );
  AND2_X1 U3768 ( .A1(n3889), .A2(n3888), .ZN(n5454) );
  NOR2_X1 U3769 ( .A1(n3870), .A2(n5624), .ZN(n3871) );
  NAND2_X1 U3770 ( .A1(n3871), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3905)
         );
  CLKBUF_X1 U3771 ( .A(n5465), .Z(n5466) );
  AND2_X1 U3772 ( .A1(n3838), .A2(n3837), .ZN(n5280) );
  NOR2_X1 U3773 ( .A1(n3807), .A2(n3806), .ZN(n3835) );
  INV_X1 U3774 ( .A(n5267), .ZN(n3064) );
  NAND2_X1 U3775 ( .A1(n3789), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3807)
         );
  NOR2_X1 U3776 ( .A1(n3784), .A2(n3783), .ZN(n3789) );
  NAND2_X1 U3777 ( .A1(n3753), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3784)
         );
  INV_X1 U3778 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3783) );
  INV_X1 U3779 ( .A(n3769), .ZN(n5012) );
  NAND2_X1 U3780 ( .A1(n3716), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3735)
         );
  INV_X1 U3781 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3734) );
  NOR2_X1 U3782 ( .A1(n3683), .A2(n3682), .ZN(n3716) );
  NAND2_X1 U3783 ( .A1(n3699), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3683)
         );
  NAND2_X1 U3784 ( .A1(n3663), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3668)
         );
  NAND2_X1 U3785 ( .A1(n3662), .A2(n3798), .ZN(n3667) );
  INV_X1 U3786 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3656) );
  NOR2_X1 U3787 ( .A1(n3653), .A2(n3656), .ZN(n3663) );
  NOR2_X1 U3788 ( .A1(n3642), .A2(n6000), .ZN(n3648) );
  NAND2_X1 U3789 ( .A1(n3648), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3653)
         );
  NOR2_X1 U3790 ( .A1(n3651), .A2(n3650), .ZN(n3652) );
  NOR2_X1 U3791 ( .A1(n5992), .A2(n3649), .ZN(n3650) );
  INV_X1 U3792 ( .A(n3647), .ZN(n3651) );
  INV_X1 U3793 ( .A(n3630), .ZN(n3631) );
  NAND2_X1 U3794 ( .A1(n3631), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3642)
         );
  NAND2_X1 U3795 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3630) );
  INV_X1 U3796 ( .A(n5482), .ZN(n3044) );
  AND2_X1 U3797 ( .A1(n4240), .A2(n4239), .ZN(n5501) );
  OR2_X1 U3798 ( .A1(n5502), .A2(n5501), .ZN(n5504) );
  NOR2_X1 U3799 ( .A1(n5286), .A2(n3048), .ZN(n5445) );
  NAND2_X1 U3800 ( .A1(n3085), .A2(n3049), .ZN(n3048) );
  AND2_X1 U3801 ( .A1(n4237), .A2(n4236), .ZN(n5444) );
  INV_X1 U3802 ( .A(n5471), .ZN(n4275) );
  INV_X1 U3803 ( .A(n3049), .ZN(n3047) );
  AND2_X1 U3804 ( .A1(n5866), .A2(n3527), .ZN(n3528) );
  NAND2_X1 U3805 ( .A1(n5268), .A2(n5269), .ZN(n5286) );
  NOR2_X1 U3806 ( .A1(n5286), .A2(n5287), .ZN(n5514) );
  NAND2_X1 U3807 ( .A1(n5216), .A2(n5188), .ZN(n5227) );
  NAND2_X1 U3808 ( .A1(n4910), .A2(n5015), .ZN(n5217) );
  NOR2_X2 U3809 ( .A1(n5217), .A2(n5218), .ZN(n5216) );
  NOR2_X1 U3810 ( .A1(n4968), .A2(n4953), .ZN(n4998) );
  NAND2_X1 U3811 ( .A1(n4998), .A2(n4999), .ZN(n4997) );
  NAND2_X1 U3812 ( .A1(n4960), .A2(n4961), .ZN(n3077) );
  NAND2_X1 U3813 ( .A1(n4756), .A2(n4967), .ZN(n4968) );
  XNOR2_X1 U3814 ( .A(n3504), .B(n6203), .ZN(n5196) );
  NAND2_X1 U3815 ( .A1(n3053), .A2(n3051), .ZN(n4757) );
  NOR2_X1 U3816 ( .A1(n4577), .A2(n3052), .ZN(n3051) );
  INV_X1 U3817 ( .A(n4576), .ZN(n3053) );
  INV_X1 U3818 ( .A(n4725), .ZN(n3052) );
  XNOR2_X1 U3819 ( .A(n3495), .B(n4176), .ZN(n4723) );
  NOR2_X1 U3820 ( .A1(n4576), .A2(n4577), .ZN(n4724) );
  NAND2_X1 U3821 ( .A1(n4494), .A2(n4495), .ZN(n4576) );
  INV_X1 U3822 ( .A(n5770), .ZN(n5740) );
  AND2_X1 U3823 ( .A1(n4158), .A2(n4157), .ZN(n4563) );
  INV_X1 U3824 ( .A(n4502), .ZN(n4507) );
  NAND2_X1 U3825 ( .A1(n3260), .A2(n3290), .ZN(n3356) );
  OR2_X1 U3826 ( .A1(n3360), .A2(n4385), .ZN(n3267) );
  NAND2_X1 U3827 ( .A1(n6490), .A2(n4523), .ZN(n4520) );
  OR2_X1 U3828 ( .A1(n3608), .A2(n3607), .ZN(n4376) );
  AND4_X1 U3829 ( .A1(n4533), .A2(n2993), .A3(n4537), .A4(n4150), .ZN(n3216)
         );
  AND3_X1 U3830 ( .A1(n4368), .A2(n4367), .A3(n4568), .ZN(n6459) );
  AND2_X1 U3831 ( .A1(n4696), .A2(n6328), .ZN(n4698) );
  AND2_X1 U3832 ( .A1(n5101), .A2(n6277), .ZN(n6371) );
  INV_X1 U3833 ( .A(n3420), .ZN(n4533) );
  INV_X1 U3834 ( .A(n3611), .ZN(n4554) );
  OR2_X1 U3835 ( .A1(n6367), .A2(n6271), .ZN(n5105) );
  NAND2_X1 U3836 ( .A1(n4524), .A2(n4523), .ZN(n4555) );
  OR2_X1 U3837 ( .A1(n4858), .A2(n4646), .ZN(n4581) );
  NAND2_X1 U3838 ( .A1(n6236), .A2(n4503), .ZN(n4858) );
  NOR2_X1 U3839 ( .A1(n4581), .A2(n3419), .ZN(n4859) );
  INV_X1 U3840 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6468) );
  NOR2_X1 U3841 ( .A1(n4147), .A2(n3610), .ZN(n6473) );
  AND2_X1 U3842 ( .A1(n6072), .A2(n4347), .ZN(n6585) );
  NAND2_X1 U3843 ( .A1(n5347), .A2(n4322), .ZN(n5965) );
  INV_X1 U3844 ( .A(n5971), .ZN(n5982) );
  INV_X1 U3845 ( .A(n5965), .ZN(n6005) );
  INV_X1 U3846 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6000) );
  INV_X1 U3847 ( .A(n5967), .ZN(n6002) );
  INV_X1 U3848 ( .A(n5524), .ZN(n5833) );
  INV_X1 U3849 ( .A(n5837), .ZN(n6043) );
  NAND2_X1 U3850 ( .A1(n4425), .A2(n6105), .ZN(n5526) );
  INV_X1 U3851 ( .A(n5225), .ZN(n5221) );
  INV_X1 U3852 ( .A(n6588), .ZN(n4431) );
  AND2_X1 U3854 ( .A1(n6490), .A2(n4484), .ZN(n6067) );
  XNOR2_X1 U3855 ( .A(n4119), .B(n4118), .ZN(n4323) );
  OR2_X1 U3856 ( .A1(n4117), .A2(n5367), .ZN(n4119) );
  OR2_X1 U3857 ( .A1(n3535), .A2(n3536), .ZN(n3537) );
  AND2_X1 U3858 ( .A1(n5715), .A2(n4301), .ZN(n5880) );
  NOR2_X1 U3859 ( .A1(n5727), .A2(n4300), .ZN(n5715) );
  CLKBUF_X1 U3860 ( .A(n5585), .Z(n5589) );
  OR2_X1 U3861 ( .A1(n5888), .A2(n4299), .ZN(n5727) );
  CLKBUF_X1 U3862 ( .A(n5294), .Z(n5295) );
  NAND2_X1 U3863 ( .A1(n2995), .A2(n3034), .ZN(n3073) );
  OAI21_X1 U3864 ( .B1(n4743), .B2(n5736), .A(n5896), .ZN(n6177) );
  NOR2_X1 U3865 ( .A1(n3039), .A2(n3031), .ZN(n3042) );
  NAND2_X1 U3866 ( .A1(n4285), .A2(n4152), .ZN(n6225) );
  AND2_X1 U3867 ( .A1(n4285), .A2(n4149), .ZN(n6227) );
  INV_X1 U3868 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6454) );
  XNOR2_X1 U3869 ( .A(n3406), .B(n3405), .ZN(n3408) );
  INV_X1 U3870 ( .A(n4507), .ZN(n6236) );
  CLKBUF_X1 U3871 ( .A(n3629), .Z(n4647) );
  NOR2_X1 U3872 ( .A1(n6573), .A2(n5407), .ZN(n5336) );
  NOR2_X1 U3873 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5340) );
  NOR2_X1 U3874 ( .A1(n4701), .A2(n3419), .ZN(n4797) );
  INV_X1 U3875 ( .A(n6243), .ZN(n6265) );
  OAI21_X1 U3876 ( .B1(n4617), .B2(n4616), .A(n4615), .ZN(n4639) );
  OAI21_X1 U3877 ( .B1(n4921), .B2(n4922), .A(n4920), .ZN(n6363) );
  INV_X1 U3878 ( .A(n6451), .ZN(n6421) );
  INV_X1 U3879 ( .A(n6407), .ZN(n6437) );
  INV_X1 U3880 ( .A(n6427), .ZN(n6445) );
  INV_X1 U3881 ( .A(n5029), .ZN(n5076) );
  AND2_X1 U3882 ( .A1(n3605), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6491) );
  INV_X1 U3883 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6493) );
  INV_X1 U3884 ( .A(READY_N), .ZN(n6728) );
  INV_X1 U3885 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6573) );
  AOI21_X1 U3886 ( .B1(n5390), .B2(n6020), .A(n5389), .ZN(n5394) );
  NOR2_X1 U3887 ( .A1(n5328), .A2(n5327), .ZN(n5329) );
  OAI21_X1 U3888 ( .B1(n5370), .B2(n6166), .A(n5369), .ZN(n5371) );
  AND2_X2 U3889 ( .A1(n3101), .A2(n3100), .ZN(n3186) );
  NAND2_X1 U3890 ( .A1(n3062), .A2(n3805), .ZN(n5224) );
  NAND2_X1 U3891 ( .A1(n2984), .A2(n3925), .ZN(n5426) );
  AND2_X1 U3892 ( .A1(n3533), .A2(n3532), .ZN(n3030) );
  NAND2_X1 U3893 ( .A1(n3461), .A2(n3488), .ZN(n3646) );
  AND2_X1 U3894 ( .A1(n4169), .A2(n4168), .ZN(n3031) );
  AND2_X1 U3895 ( .A1(n5471), .A2(n4565), .ZN(n4161) );
  AND2_X2 U3896 ( .A1(n4391), .A2(n4374), .ZN(n3275) );
  NAND2_X1 U3897 ( .A1(n4533), .A2(n4145), .ZN(n4211) );
  INV_X1 U3898 ( .A(n4145), .ZN(n4548) );
  NAND2_X1 U3899 ( .A1(n5620), .A2(n3525), .ZN(n5631) );
  NAND2_X1 U3900 ( .A1(n3014), .A2(n3091), .ZN(n5558) );
  INV_X1 U3901 ( .A(n4503), .ZN(n4506) );
  NAND2_X1 U3902 ( .A1(n3379), .A2(n3378), .ZN(n4503) );
  AND2_X1 U3903 ( .A1(n4308), .A2(n3061), .ZN(n5488) );
  AND2_X1 U3904 ( .A1(n2992), .A2(n5774), .ZN(n5629) );
  NAND2_X1 U3905 ( .A1(n4308), .A2(n3060), .ZN(n5478) );
  AND2_X1 U3906 ( .A1(n4308), .A2(n4307), .ZN(n4309) );
  AND2_X2 U3907 ( .A1(n3101), .A2(n4471), .ZN(n3370) );
  INV_X1 U3908 ( .A(n3219), .ZN(n5527) );
  INV_X1 U3909 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3251) );
  AND2_X1 U3910 ( .A1(n3222), .A2(n3221), .ZN(n3606) );
  NAND2_X1 U3911 ( .A1(n3066), .A2(n3069), .ZN(n5250) );
  NAND2_X1 U3912 ( .A1(n3073), .A2(n5166), .ZN(n5240) );
  NAND2_X1 U3913 ( .A1(n3077), .A2(n3515), .ZN(n5200) );
  OAI22_X1 U3914 ( .A1(n3233), .A2(n3212), .B1(n4548), .B2(n4537), .ZN(n4267)
         );
  NAND2_X1 U3915 ( .A1(n3772), .A2(n3771), .ZN(n5183) );
  XNOR2_X1 U3916 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(n2992), .ZN(n3033)
         );
  INV_X1 U3917 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6490) );
  INV_X1 U3918 ( .A(n5184), .ZN(n3062) );
  NOR2_X1 U3919 ( .A1(n5286), .A2(n3047), .ZN(n5456) );
  NAND2_X1 U3920 ( .A1(n3518), .A2(n3517), .ZN(n3034) );
  AND2_X1 U3921 ( .A1(n4908), .A2(n3752), .ZN(n3035) );
  AND2_X1 U3922 ( .A1(n4999), .A2(n3046), .ZN(n3036) );
  NAND2_X1 U3923 ( .A1(n2992), .A2(n5756), .ZN(n3037) );
  NAND2_X1 U3924 ( .A1(n3418), .A2(n3417), .ZN(n5097) );
  INV_X1 U3925 ( .A(n3754), .ZN(n4109) );
  NOR2_X1 U3926 ( .A1(n4757), .A2(n4758), .ZN(n4756) );
  XNOR2_X1 U3927 ( .A(n3469), .B(n3468), .ZN(n4739) );
  OAI211_X1 U3928 ( .C1(n3059), .C2(n3058), .A(n3057), .B(n3055), .ZN(n4454)
         );
  INV_X1 U3929 ( .A(n4124), .ZN(n3241) );
  INV_X1 U3930 ( .A(n5223), .ZN(n3805) );
  AND3_X1 U3931 ( .A1(n3227), .A2(n4533), .A3(n4537), .ZN(n3038) );
  AND2_X1 U3932 ( .A1(n4574), .A2(n4573), .ZN(n3039) );
  AND2_X1 U3933 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3040) );
  INV_X1 U3934 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3806) );
  NOR2_X1 U3935 ( .A1(n4494), .A2(n3042), .ZN(n6019) );
  INV_X1 U3936 ( .A(n3045), .ZN(n5685) );
  NOR2_X4 U3937 ( .A1(n3045), .A2(n3044), .ZN(n5484) );
  NAND2_X1 U3938 ( .A1(n5445), .A2(n5444), .ZN(n5502) );
  INV_X2 U3939 ( .A(n4565), .ZN(n5396) );
  NAND2_X1 U3940 ( .A1(n4502), .A2(n3798), .ZN(n3057) );
  NAND2_X1 U3941 ( .A1(n3057), .A2(n3754), .ZN(n3626) );
  NAND2_X1 U3942 ( .A1(n3028), .A2(n3798), .ZN(n3059) );
  NAND2_X1 U3943 ( .A1(n5266), .A2(n5280), .ZN(n5279) );
  NAND3_X1 U3944 ( .A1(n3733), .A2(n4906), .A3(n4908), .ZN(n4907) );
  NAND2_X1 U3945 ( .A1(n2984), .A2(n3065), .ZN(n5413) );
  NAND2_X1 U3946 ( .A1(n2995), .A2(n3067), .ZN(n3066) );
  AND2_X1 U3947 ( .A1(n3081), .A2(n3515), .ZN(n3076) );
  INV_X1 U3948 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3234) );
  INV_X1 U3950 ( .A(n3170), .ZN(n3227) );
  INV_X1 U3951 ( .A(n3327), .ZN(n3291) );
  OR2_X1 U3952 ( .A1(n3518), .A2(n6194), .ZN(n3081) );
  NOR2_X1 U3953 ( .A1(n6274), .A2(n4764), .ZN(n3082) );
  OR2_X1 U3954 ( .A1(n3255), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3083)
         );
  AND3_X1 U3955 ( .A1(n3696), .A2(n3695), .A3(n3694), .ZN(n3084) );
  AND2_X1 U3956 ( .A1(n4233), .A2(n4232), .ZN(n3085) );
  OR2_X1 U3957 ( .A1(n5476), .A2(n6009), .ZN(n3086) );
  NAND2_X1 U3958 ( .A1(n5320), .A2(n5319), .ZN(n5476) );
  AND4_X1 U3959 ( .A1(n3315), .A2(n3314), .A3(n3313), .A4(n3312), .ZN(n3087)
         );
  AND2_X1 U3960 ( .A1(n3311), .A2(n3310), .ZN(n3088) );
  NOR2_X1 U3961 ( .A1(n5513), .A2(n5453), .ZN(n3089) );
  AND4_X1 U3962 ( .A1(n3182), .A2(n3181), .A3(n3180), .A4(n3179), .ZN(n3090)
         );
  AND2_X1 U3963 ( .A1(n5836), .A2(n5527), .ZN(n5831) );
  NAND2_X1 U3964 ( .A1(n6481), .A2(n6656), .ZN(n3649) );
  AND2_X1 U3965 ( .A1(n2992), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3091)
         );
  OR2_X1 U3966 ( .A1(n4561), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3092)
         );
  INV_X1 U3967 ( .A(n3623), .ZN(n3973) );
  NOR2_X1 U3968 ( .A1(n6274), .A2(n4836), .ZN(n3093) );
  AND3_X1 U3969 ( .A1(n3666), .A2(n3665), .A3(n3664), .ZN(n3094) );
  INV_X1 U3970 ( .A(n5836), .ZN(n5499) );
  AND2_X2 U3971 ( .A1(n4569), .A2(n6491), .ZN(n5836) );
  AND2_X2 U3972 ( .A1(n5914), .A2(n4114), .ZN(n6156) );
  OR2_X1 U3973 ( .A1(n3548), .A2(n3559), .ZN(n3553) );
  NOR2_X1 U3974 ( .A1(n6490), .A2(n5343), .ZN(n3235) );
  OR2_X1 U3975 ( .A1(n3390), .A2(n3389), .ZN(n3394) );
  NAND2_X1 U3976 ( .A1(n3508), .A2(n3393), .ZN(n3282) );
  OR2_X1 U3977 ( .A1(n3594), .A2(n3462), .ZN(n3391) );
  INV_X1 U3978 ( .A(n5468), .ZN(n3854) );
  OR2_X1 U3979 ( .A1(n3594), .A2(n3489), .ZN(n3457) );
  INV_X1 U3980 ( .A(n3308), .ZN(n3318) );
  AOI22_X1 U3981 ( .A1(n3015), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3275), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3168) );
  INV_X1 U3982 ( .A(n3365), .ZN(n3284) );
  OR2_X1 U3983 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n3592), .ZN(n3584)
         );
  INV_X1 U3984 ( .A(n5506), .ZN(n3925) );
  INV_X1 U3985 ( .A(n4900), .ZN(n3660) );
  OR2_X1 U3986 ( .A1(n3318), .A2(n3317), .ZN(n3510) );
  INV_X1 U3987 ( .A(n3464), .ZN(n3489) );
  AND2_X1 U3988 ( .A1(n3585), .A2(n3584), .ZN(n4135) );
  INV_X1 U3989 ( .A(n5427), .ZN(n3956) );
  NOR2_X1 U3990 ( .A1(n4057), .A2(n4056), .ZN(n4058) );
  AND2_X1 U3991 ( .A1(n3484), .A2(n3483), .ZN(n3487) );
  AND3_X1 U3992 ( .A1(n3508), .A2(n3550), .A3(n3510), .ZN(n3509) );
  AND2_X1 U3993 ( .A1(n4565), .A2(n4251), .ZN(n4234) );
  NAND2_X1 U3994 ( .A1(n5334), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4078) );
  AND2_X1 U3995 ( .A1(n3951), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3992)
         );
  INV_X1 U3996 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3682) );
  OR2_X1 U3997 ( .A1(n3437), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6159)
         );
  OR2_X1 U3998 ( .A1(n3021), .A2(n5782), .ZN(n5100) );
  AOI21_X1 U3999 ( .B1(n5351), .B2(REIP_REG_31__SCAN_IN), .A(n5350), .ZN(n5352) );
  NAND2_X1 U4000 ( .A1(n5189), .A2(REIP_REG_14__SCAN_IN), .ZN(n5285) );
  INV_X1 U4001 ( .A(n3668), .ZN(n3699) );
  OR2_X1 U4002 ( .A1(n5963), .A2(n6573), .ZN(n6023) );
  OR2_X1 U4003 ( .A1(n5963), .A2(n6481), .ZN(n5089) );
  INV_X1 U4004 ( .A(n4110), .ZN(n4111) );
  AND2_X1 U4005 ( .A1(n3992), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3993)
         );
  INV_X1 U4006 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5624) );
  INV_X1 U4007 ( .A(n4754), .ZN(n4755) );
  INV_X1 U4008 ( .A(n6156), .ZN(n6171) );
  AND2_X1 U4009 ( .A1(n2992), .A2(n5573), .ZN(n5574) );
  INV_X1 U4010 ( .A(n6215), .ZN(n5900) );
  INV_X1 U4011 ( .A(n5336), .ZN(n6483) );
  INV_X1 U4012 ( .A(n6491), .ZN(n4369) );
  INV_X1 U4013 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4695) );
  INV_X1 U4014 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5106) );
  AOI21_X1 U4015 ( .B1(n6454), .B2(STATE2_REG_3__SCAN_IN), .A(n4520), .ZN(
        n6326) );
  OR2_X1 U4016 ( .A1(n4124), .A2(n6580), .ZN(n6480) );
  OR2_X1 U4017 ( .A1(n4344), .A2(n4369), .ZN(n4347) );
  INV_X1 U4018 ( .A(n5352), .ZN(n5353) );
  NAND2_X1 U4019 ( .A1(n3086), .A2(n5329), .ZN(n5330) );
  NAND2_X1 U4020 ( .A1(n5347), .A2(n4334), .ZN(n6009) );
  NOR2_X1 U4021 ( .A1(n6756), .A2(n5460), .ZN(n5442) );
  OR2_X1 U4022 ( .A1(n4323), .A2(n6493), .ZN(n4319) );
  INV_X1 U4023 ( .A(n6023), .ZN(n5978) );
  INV_X1 U4024 ( .A(n6009), .ZN(n6020) );
  XNOR2_X1 U4025 ( .A(n4266), .B(n4265), .ZN(n5344) );
  AND2_X1 U4026 ( .A1(n5526), .A2(n5375), .ZN(n6042) );
  NOR2_X1 U4027 ( .A1(n6049), .A2(n4431), .ZN(n6066) );
  OAI21_X1 U4028 ( .B1(n4335), .B2(n6728), .A(n6073), .ZN(n6088) );
  INV_X1 U4029 ( .A(n6105), .ZN(n6151) );
  INV_X1 U4030 ( .A(n6166), .ZN(n5642) );
  INV_X1 U4031 ( .A(n4351), .ZN(n6071) );
  INV_X1 U4032 ( .A(n5914), .ZN(n6173) );
  CLKBUF_X1 U4033 ( .A(n4490), .Z(n4491) );
  INV_X1 U4034 ( .A(n5739), .ZN(n6209) );
  OAI21_X1 U4035 ( .B1(n4802), .B2(n4803), .A(n4801), .ZN(n4825) );
  INV_X1 U4036 ( .A(n4721), .ZN(n4691) );
  OAI21_X1 U4037 ( .B1(n6249), .B2(n6248), .A(n6247), .ZN(n6267) );
  AND2_X1 U4038 ( .A1(n4760), .A2(n3419), .ZN(n6266) );
  NOR2_X1 U4039 ( .A1(n6272), .A2(n4857), .ZN(n6314) );
  INV_X1 U4040 ( .A(n6318), .ZN(n6345) );
  INV_X1 U4041 ( .A(n6366), .ZN(n6346) );
  OR2_X1 U4042 ( .A1(n3029), .A2(n5097), .ZN(n4857) );
  INV_X1 U4043 ( .A(n5105), .ZN(n6422) );
  INV_X1 U4044 ( .A(n6397), .ZN(n6431) );
  OAI211_X1 U4045 ( .C1(n6442), .C2(n6573), .A(n4839), .B(n4838), .ZN(n6448)
         );
  NOR2_X2 U4046 ( .A1(n4858), .A2(n4833), .ZN(n6446) );
  NOR2_X1 U4047 ( .A1(n4858), .A2(n4857), .ZN(n5029) );
  INV_X2 U4048 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6481) );
  INV_X1 U4049 ( .A(n6564), .ZN(n6559) );
  NAND2_X1 U4050 ( .A1(n6071), .A2(n4312), .ZN(n6072) );
  AND2_X1 U4051 ( .A1(n4126), .A2(STATE_REG_1__SCAN_IN), .ZN(n6789) );
  AOI21_X1 U4052 ( .B1(n5344), .B2(n6020), .A(n5353), .ZN(n5355) );
  INV_X1 U4053 ( .A(n6018), .ZN(n5954) );
  OR2_X1 U4054 ( .A1(n5963), .A2(n5397), .ZN(n5967) );
  OR2_X1 U4055 ( .A1(n5963), .A2(n4324), .ZN(n6022) );
  INV_X1 U4056 ( .A(n5344), .ZN(n5358) );
  NAND2_X1 U4057 ( .A1(n5836), .A2(n3219), .ZN(n5524) );
  OR2_X1 U4058 ( .A1(n4978), .A2(n4977), .ZN(n5177) );
  NAND2_X1 U4059 ( .A1(n5526), .A2(n4426), .ZN(n5837) );
  INV_X1 U4060 ( .A(n6049), .ZN(n6069) );
  OR2_X1 U4061 ( .A1(n4976), .A2(n4952), .ZN(n5206) );
  INV_X1 U4062 ( .A(n6227), .ZN(n5779) );
  INV_X1 U4063 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6234) );
  INV_X1 U4064 ( .A(n4797), .ZN(n4832) );
  NAND2_X1 U4065 ( .A1(n4650), .A2(n3419), .ZN(n4721) );
  AOI21_X1 U4066 ( .B1(n4655), .B2(n4654), .A(n4653), .ZN(n4694) );
  INV_X1 U4067 ( .A(n6266), .ZN(n4795) );
  OR2_X1 U4068 ( .A1(n6272), .A2(n6271), .ZN(n6318) );
  OR2_X1 U4069 ( .A1(n6272), .A2(n4914), .ZN(n6366) );
  OR2_X1 U4070 ( .A1(n6367), .A2(n4857), .ZN(n5140) );
  AOI22_X1 U4071 ( .A1(n5108), .A2(n6371), .B1(n6274), .B2(n5104), .ZN(n5143)
         );
  OR2_X1 U4072 ( .A1(n6367), .A2(n4914), .ZN(n6451) );
  INV_X1 U4073 ( .A(n4859), .ZN(n4899) );
  INV_X1 U4074 ( .A(n6568), .ZN(n6503) );
  INV_X1 U4075 ( .A(n6562), .ZN(n6561) );
  AND2_X4 U4076 ( .A1(n3251), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3099)
         );
  AND2_X2 U4077 ( .A1(n3099), .A2(n4392), .ZN(n3196) );
  AOI22_X1 U4078 ( .A1(n3196), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3098) );
  NOR2_X4 U4079 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3100) );
  INV_X1 U4080 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4081 ( .A1(n3023), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3268), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3097) );
  NOR2_X4 U4082 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4375) );
  AOI22_X1 U4083 ( .A1(n3333), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3096) );
  AND2_X4 U4084 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4374) );
  AOI22_X1 U4085 ( .A1(n3335), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3191), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3095) );
  NAND4_X1 U4086 ( .A1(n3098), .A2(n3097), .A3(n3096), .A4(n3095), .ZN(n3107)
         );
  AOI22_X1 U4087 ( .A1(n3275), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3201), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3105) );
  AOI22_X1 U4088 ( .A1(n3185), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3186), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3104) );
  AOI22_X1 U4089 ( .A1(n3328), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3020), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3103) );
  AOI22_X1 U4090 ( .A1(n3269), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3102) );
  NAND4_X1 U4091 ( .A1(n3105), .A2(n3104), .A3(n3103), .A4(n3102), .ZN(n3106)
         );
  AOI22_X1 U4092 ( .A1(n3335), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3191), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3108) );
  AOI22_X1 U4093 ( .A1(n3015), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3275), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3115) );
  AOI22_X1 U4094 ( .A1(n3370), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3201), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3113) );
  AOI22_X1 U4095 ( .A1(n3023), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3121) );
  AOI22_X1 U4096 ( .A1(n3018), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3191), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3124) );
  AOI22_X1 U4097 ( .A1(n3026), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3123) );
  AOI22_X1 U4098 ( .A1(n3275), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3201), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3122) );
  AND4_X2 U4099 ( .A1(n3125), .A2(n3124), .A3(n3123), .A4(n3122), .ZN(n3126)
         );
  AOI22_X1 U4100 ( .A1(n3185), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        INSTQUEUE_REG_2__4__SCAN_IN), .B2(n3186), .ZN(n3131) );
  AOI22_X1 U4101 ( .A1(n3328), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3268), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3130) );
  AOI22_X1 U4102 ( .A1(n3293), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3129) );
  AOI22_X1 U4103 ( .A1(n3335), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3191), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3128) );
  AOI22_X1 U4104 ( .A1(n3196), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3275), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3135) );
  AOI22_X1 U4105 ( .A1(n3023), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3134) );
  AOI22_X1 U4106 ( .A1(n3370), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3201), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3133) );
  AOI22_X1 U4107 ( .A1(n3174), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3132) );
  NAND2_X1 U4108 ( .A1(n3196), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3141) );
  NAND2_X1 U4109 ( .A1(n3370), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3140)
         );
  NAND2_X1 U4110 ( .A1(n3275), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3139) );
  NAND2_X1 U4111 ( .A1(n3201), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3138) );
  NAND2_X1 U4112 ( .A1(n3185), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3145) );
  NAND2_X1 U4113 ( .A1(n3186), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3144) );
  NAND2_X1 U4114 ( .A1(n3335), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3143)
         );
  NAND2_X1 U4115 ( .A1(n3191), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3142) );
  NAND2_X1 U4116 ( .A1(n3293), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3149)
         );
  NAND2_X1 U4117 ( .A1(n3328), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3148)
         );
  NAND2_X1 U4118 ( .A1(n3026), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3147) );
  NAND2_X1 U4119 ( .A1(n3269), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3146) );
  NAND2_X1 U4120 ( .A1(n3023), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3153) );
  NAND2_X1 U4121 ( .A1(n3333), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3152) );
  NAND2_X1 U4122 ( .A1(n3309), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3151)
         );
  NAND2_X1 U4123 ( .A1(n3174), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3150)
         );
  NAND2_X1 U4124 ( .A1(n3158), .A2(n3219), .ZN(n3159) );
  OAI21_X1 U4125 ( .B1(n4271), .B2(n3546), .A(n3159), .ZN(n3169) );
  NOR2_X2 U4126 ( .A1(n3160), .A2(n3611), .ZN(n3218) );
  AOI22_X1 U4127 ( .A1(n3023), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3164) );
  AOI22_X1 U4128 ( .A1(n3328), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3185), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3163) );
  AOI22_X1 U4129 ( .A1(n3020), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3162) );
  AOI22_X1 U4130 ( .A1(n3174), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3161) );
  AOI22_X1 U4131 ( .A1(n3018), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3191), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3167) );
  AOI22_X1 U4132 ( .A1(n3370), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3201), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3165) );
  AND2_X2 U4133 ( .A1(n3169), .A2(n3215), .ZN(n3172) );
  NAND2_X1 U4134 ( .A1(n3227), .A2(n3611), .ZN(n3220) );
  NAND2_X1 U4135 ( .A1(n3220), .A2(n3211), .ZN(n3213) );
  NAND2_X1 U4136 ( .A1(n3172), .A2(n4537), .ZN(n3173) );
  NAND2_X1 U4137 ( .A1(n3243), .A2(n3173), .ZN(n3184) );
  AOI22_X1 U4138 ( .A1(n3023), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3178) );
  AOI22_X1 U4139 ( .A1(n3196), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3275), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3177) );
  AOI22_X1 U4140 ( .A1(n3370), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3201), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3176) );
  AOI22_X1 U4141 ( .A1(n3174), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3175) );
  AOI22_X1 U4142 ( .A1(n3293), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3182) );
  AOI22_X1 U4143 ( .A1(n3335), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3191), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3181) );
  AOI22_X1 U4144 ( .A1(n3328), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3268), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3180) );
  AOI22_X1 U4145 ( .A1(n3185), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3186), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3179) );
  NAND2_X2 U4146 ( .A1(n3183), .A2(n3090), .ZN(n4268) );
  NAND2_X1 U4147 ( .A1(n3184), .A2(n4525), .ZN(n3210) );
  NAND2_X1 U4148 ( .A1(n3333), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3190) );
  NAND2_X1 U4149 ( .A1(n3185), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3189) );
  NAND2_X1 U4150 ( .A1(n3186), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3188) );
  NAND2_X1 U4151 ( .A1(n3269), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3187) );
  NAND2_X1 U4152 ( .A1(n3328), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3195)
         );
  NAND2_X1 U4153 ( .A1(n3268), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3194) );
  NAND2_X1 U4154 ( .A1(n3335), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3193)
         );
  NAND2_X1 U4155 ( .A1(n3191), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3192) );
  NAND2_X1 U4156 ( .A1(n3275), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3199) );
  NAND2_X1 U4157 ( .A1(n3370), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3198)
         );
  NAND2_X1 U4158 ( .A1(n3309), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3197)
         );
  NAND3_X1 U4159 ( .A1(n3199), .A2(n3198), .A3(n3197), .ZN(n3200) );
  NAND2_X1 U4160 ( .A1(n3293), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3205)
         );
  NAND2_X1 U4161 ( .A1(n3023), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3204) );
  NAND2_X1 U4162 ( .A1(n3174), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3203)
         );
  NAND2_X1 U4163 ( .A1(n3201), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3202) );
  NAND2_X1 U4164 ( .A1(n3210), .A2(n4548), .ZN(n3233) );
  AND2_X1 U4165 ( .A1(n3550), .A2(n4529), .ZN(n3212) );
  INV_X1 U4166 ( .A(n4267), .ZN(n3226) );
  OAI21_X1 U4167 ( .B1(n3238), .B2(n3215), .A(n3395), .ZN(n3217) );
  AND2_X1 U4168 ( .A1(n5340), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6492) );
  NAND2_X2 U4169 ( .A1(n3420), .A2(n4268), .ZN(n4251) );
  NAND2_X1 U4170 ( .A1(n3211), .A2(n3546), .ZN(n3610) );
  NAND2_X1 U4171 ( .A1(n3216), .A2(n3616), .ZN(n4403) );
  NAND4_X1 U4172 ( .A1(n3217), .A2(n6492), .A3(n4371), .A4(n4403), .ZN(n3224)
         );
  NAND2_X1 U4173 ( .A1(n3218), .A2(n4529), .ZN(n3222) );
  AND2_X1 U4174 ( .A1(n3220), .A2(n3219), .ZN(n3221) );
  OAI211_X1 U4175 ( .C1(n4529), .C2(n3218), .A(n3606), .B(n3420), .ZN(n3230)
         );
  AND2_X1 U4176 ( .A1(n3230), .A2(n4268), .ZN(n3223) );
  NAND2_X1 U4177 ( .A1(n3238), .A2(n3395), .ZN(n3229) );
  XNOR2_X1 U4178 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .ZN(
        n4125) );
  NAND2_X1 U4179 ( .A1(n4525), .A2(n4125), .ZN(n3242) );
  INV_X1 U4180 ( .A(n4537), .ZN(n4272) );
  AOI21_X1 U4181 ( .B1(n3227), .B2(n3242), .A(n4272), .ZN(n3228) );
  NAND3_X1 U4182 ( .A1(n4371), .A2(n3229), .A3(n3228), .ZN(n3231) );
  NOR2_X1 U4183 ( .A1(n3231), .A2(n3230), .ZN(n3232) );
  NAND2_X1 U4184 ( .A1(n3233), .A2(n3232), .ZN(n3253) );
  NAND2_X1 U4185 ( .A1(n3253), .A2(n3235), .ZN(n3237) );
  NAND2_X1 U4186 ( .A1(n5340), .A2(n6490), .ZN(n6587) );
  MUX2_X1 U4187 ( .A(n6587), .B(n3605), .S(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .Z(n3236) );
  NAND2_X1 U4188 ( .A1(n3237), .A2(n3236), .ZN(n3323) );
  INV_X1 U4189 ( .A(n3242), .ZN(n3247) );
  INV_X1 U4190 ( .A(n3243), .ZN(n3244) );
  INV_X1 U4191 ( .A(n3545), .ZN(n3245) );
  NAND2_X1 U4192 ( .A1(n3244), .A2(n3245), .ZN(n4144) );
  INV_X1 U4193 ( .A(n4420), .ZN(n3246) );
  INV_X1 U4194 ( .A(n4271), .ZN(n5375) );
  NAND2_X1 U4195 ( .A1(n3246), .A2(n5375), .ZN(n4151) );
  OAI211_X1 U4196 ( .C1(n5401), .C2(n3247), .A(n4144), .B(n4151), .ZN(n3248)
         );
  NAND2_X1 U4197 ( .A1(n3248), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3257) );
  INV_X1 U4198 ( .A(n3257), .ZN(n3252) );
  INV_X1 U4199 ( .A(n6587), .ZN(n3265) );
  XNOR2_X1 U4200 ( .A(n5106), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6274)
         );
  NAND2_X1 U4201 ( .A1(n3265), .A2(n6274), .ZN(n3250) );
  INV_X1 U4202 ( .A(n3605), .ZN(n3264) );
  NAND2_X1 U4203 ( .A1(n3264), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3249) );
  NAND2_X1 U4204 ( .A1(n3250), .A2(n3249), .ZN(n3255) );
  NAND2_X1 U4205 ( .A1(n3327), .A2(n3289), .ZN(n3260) );
  NAND2_X1 U4206 ( .A1(n3253), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3360) );
  INV_X1 U4207 ( .A(n3360), .ZN(n3254) );
  INV_X1 U4208 ( .A(n3255), .ZN(n3256) );
  INV_X1 U4209 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4385) );
  AND2_X1 U4210 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3261) );
  NAND2_X1 U4211 ( .A1(n3261), .A2(n4695), .ZN(n6372) );
  INV_X1 U4212 ( .A(n3261), .ZN(n3262) );
  NAND2_X1 U4213 ( .A1(n3262), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3263) );
  NAND2_X1 U4214 ( .A1(n6372), .A2(n3263), .ZN(n4656) );
  AOI22_X1 U4215 ( .A1(n3265), .A2(n4656), .B1(n3264), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3266) );
  NAND2_X1 U4216 ( .A1(n4401), .A2(n6490), .ZN(n3283) );
  AOI22_X1 U4217 ( .A1(n4062), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3273) );
  AOI22_X1 U4218 ( .A1(n3027), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3272) );
  AOI22_X1 U4219 ( .A1(n2990), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3271) );
  AOI22_X1 U4220 ( .A1(n4084), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3270) );
  NAND4_X1 U4221 ( .A1(n3273), .A2(n3272), .A3(n3271), .A4(n3270), .ZN(n3281)
         );
  AOI22_X1 U4222 ( .A1(n3023), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3334), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3279) );
  INV_X1 U4223 ( .A(n3275), .ZN(n4388) );
  AOI22_X1 U4224 ( .A1(n3196), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3278) );
  AOI22_X1 U4225 ( .A1(n3370), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3277) );
  AOI22_X1 U4226 ( .A1(n4067), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3276) );
  NAND4_X1 U4227 ( .A1(n3279), .A2(n3278), .A3(n3277), .A4(n3276), .ZN(n3280)
         );
  NAND2_X1 U4228 ( .A1(n3569), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3286) );
  NOR2_X1 U4229 ( .A1(n4145), .A2(n6490), .ZN(n3306) );
  NAND2_X1 U4230 ( .A1(n3306), .A2(n3393), .ZN(n3285) );
  NAND2_X1 U4231 ( .A1(n3286), .A2(n3285), .ZN(n3287) );
  INV_X1 U4232 ( .A(n3428), .ZN(n3355) );
  NAND2_X1 U4233 ( .A1(n3290), .A2(n3289), .ZN(n3292) );
  NAND2_X1 U4234 ( .A1(n4370), .A2(n6490), .ZN(n3305) );
  AOI22_X1 U4235 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n3022), .B1(n2990), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3297) );
  AOI22_X1 U4236 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n4084), .B1(n3027), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4237 ( .A1(n3019), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3295) );
  AOI22_X1 U4238 ( .A1(n3023), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3294) );
  NAND4_X1 U4239 ( .A1(n3297), .A2(n3296), .A3(n3295), .A4(n3294), .ZN(n3303)
         );
  AOI22_X1 U4240 ( .A1(n3196), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4241 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n4062), .B1(n4091), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U4242 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n3334), .B1(n3016), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4243 ( .A1(n3186), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3191), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3298) );
  NAND4_X1 U4244 ( .A1(n3301), .A2(n3300), .A3(n3299), .A4(n3298), .ZN(n3302)
         );
  NAND2_X1 U4245 ( .A1(n3508), .A2(n3409), .ZN(n3304) );
  INV_X1 U4246 ( .A(n3409), .ZN(n3321) );
  INV_X1 U4247 ( .A(n3306), .ZN(n3320) );
  NAND2_X1 U4248 ( .A1(n3569), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3319) );
  AOI22_X1 U4249 ( .A1(n3370), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4250 ( .A1(n4067), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4251 ( .A1(n3027), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3018), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U4252 ( .A1(n3186), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4253 ( .A1(n3023), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3334), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3315) );
  AOI22_X1 U4254 ( .A1(n2990), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4255 ( .A1(n3196), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4256 ( .A1(n4062), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3191), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3312) );
  NAND3_X1 U4257 ( .A1(n3316), .A2(n3088), .A3(n3087), .ZN(n3317) );
  INV_X1 U4258 ( .A(n3322), .ZN(n3325) );
  INV_X1 U4259 ( .A(n3323), .ZN(n3324) );
  AOI22_X1 U4260 ( .A1(n3196), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3019), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3332) );
  AOI22_X1 U4261 ( .A1(n3023), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3331) );
  AOI22_X1 U4262 ( .A1(n4062), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3330) );
  AOI22_X1 U4263 ( .A1(n3027), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3186), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3329) );
  NAND4_X1 U4264 ( .A1(n3332), .A2(n3331), .A3(n3330), .A4(n3329), .ZN(n3341)
         );
  AOI22_X1 U4265 ( .A1(n3334), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3339) );
  AOI22_X1 U4266 ( .A1(n4090), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3338) );
  AOI22_X1 U4267 ( .A1(n4084), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3191), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3337) );
  AOI22_X1 U4268 ( .A1(n4067), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3336) );
  NAND4_X1 U4269 ( .A1(n3339), .A2(n3338), .A3(n3337), .A4(n3336), .ZN(n3340)
         );
  NAND2_X1 U4270 ( .A1(n3343), .A2(n4529), .ZN(n3344) );
  OAI21_X2 U4271 ( .B1(n3617), .B2(STATE2_REG_0__SCAN_IN), .A(n3346), .ZN(
        n3351) );
  NAND2_X1 U4272 ( .A1(n3569), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3350) );
  NAND2_X1 U4273 ( .A1(n4548), .A2(n3421), .ZN(n3347) );
  OAI211_X1 U4274 ( .C1(n3499), .C2(n4150), .A(STATE2_REG_0__SCAN_IN), .B(
        n3347), .ZN(n3348) );
  INV_X1 U4275 ( .A(n3348), .ZN(n3349) );
  NAND2_X1 U4276 ( .A1(n3350), .A2(n3349), .ZN(n3414) );
  NAND2_X1 U4277 ( .A1(n3508), .A2(n3510), .ZN(n3352) );
  OAI21_X1 U4278 ( .B1(n3407), .B2(n3405), .A(n2988), .ZN(n3354) );
  NAND2_X1 U4279 ( .A1(n3407), .A2(n3405), .ZN(n3353) );
  NAND2_X1 U4280 ( .A1(n3354), .A2(n3353), .ZN(n3427) );
  INV_X1 U4281 ( .A(n3399), .ZN(n3380) );
  INV_X1 U4282 ( .A(n3356), .ZN(n3358) );
  OR2_X1 U4283 ( .A1(n3360), .A2(n3359), .ZN(n3364) );
  NOR3_X1 U4284 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4695), .A3(n5106), 
        .ZN(n6329) );
  NAND2_X1 U4285 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6329), .ZN(n6321) );
  NAND2_X1 U4286 ( .A1(n6468), .A2(n6321), .ZN(n3361) );
  NOR3_X1 U4287 ( .A1(n6468), .A2(n4695), .A3(n5106), .ZN(n4862) );
  NAND2_X1 U4288 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4862), .ZN(n4606) );
  NAND2_X1 U4289 ( .A1(n3361), .A2(n4606), .ZN(n4836) );
  OAI22_X1 U4290 ( .A1(n6587), .A2(n4836), .B1(n3605), .B2(n6468), .ZN(n3362)
         );
  INV_X1 U4291 ( .A(n3362), .ZN(n3363) );
  INV_X1 U4292 ( .A(n3594), .ZN(n3377) );
  AOI22_X1 U4293 ( .A1(n4062), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4294 ( .A1(n3027), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4295 ( .A1(n2991), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4296 ( .A1(n4084), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3366) );
  NAND4_X1 U4297 ( .A1(n3369), .A2(n3368), .A3(n3367), .A4(n3366), .ZN(n3376)
         );
  AOI22_X1 U4298 ( .A1(n3023), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3334), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4299 ( .A1(n3721), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4300 ( .A1(n3307), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3372) );
  AOI22_X1 U4301 ( .A1(n4067), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3371) );
  NAND4_X1 U4302 ( .A1(n3374), .A2(n3373), .A3(n3372), .A4(n3371), .ZN(n3375)
         );
  AOI22_X1 U4303 ( .A1(n3377), .A2(n3400), .B1(n3569), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3378) );
  NAND2_X1 U4304 ( .A1(n3569), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3392) );
  AOI22_X1 U4305 ( .A1(n4062), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3384) );
  AOI22_X1 U4306 ( .A1(n3027), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3383) );
  AOI22_X1 U4307 ( .A1(n2991), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4308 ( .A1(n4084), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3381) );
  NAND4_X1 U4309 ( .A1(n3384), .A2(n3383), .A3(n3382), .A4(n3381), .ZN(n3390)
         );
  AOI22_X1 U4310 ( .A1(n3023), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3334), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3388) );
  AOI22_X1 U4311 ( .A1(n3721), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3387) );
  AOI22_X1 U4312 ( .A1(n3307), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3386) );
  AOI22_X1 U4313 ( .A1(n4067), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3385) );
  NAND4_X1 U4314 ( .A1(n3388), .A2(n3387), .A3(n3386), .A4(n3385), .ZN(n3389)
         );
  NAND2_X1 U4315 ( .A1(n3637), .A2(n3550), .ZN(n3398) );
  NAND2_X1 U4316 ( .A1(n3421), .A2(n3409), .ZN(n3431) );
  INV_X1 U4317 ( .A(n3393), .ZN(n3430) );
  NAND2_X1 U4318 ( .A1(n3431), .A2(n3430), .ZN(n3429) );
  NAND2_X1 U4319 ( .A1(n3429), .A2(n3400), .ZN(n3463) );
  XNOR2_X1 U4320 ( .A(n3463), .B(n3394), .ZN(n3396) );
  NAND2_X1 U4321 ( .A1(n3396), .A2(n4335), .ZN(n3397) );
  INV_X1 U4322 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4170) );
  XNOR2_X1 U4323 ( .A(n3441), .B(n4170), .ZN(n4489) );
  NAND2_X1 U4324 ( .A1(n3629), .A2(n3550), .ZN(n3404) );
  INV_X1 U4325 ( .A(n3400), .ZN(n3401) );
  XNOR2_X1 U4326 ( .A(n3429), .B(n3401), .ZN(n3402) );
  NAND2_X1 U4327 ( .A1(n3402), .A2(n4335), .ZN(n3403) );
  NAND2_X1 U4328 ( .A1(n3029), .A2(n3550), .ZN(n3413) );
  OAI21_X1 U4329 ( .B1(n3409), .B2(n3421), .A(n3431), .ZN(n3410) );
  OAI211_X1 U4330 ( .C1(n3410), .C2(n6580), .A(n4269), .B(n3546), .ZN(n3411)
         );
  INV_X1 U4331 ( .A(n3411), .ZN(n3412) );
  INV_X1 U4332 ( .A(n3414), .ZN(n3416) );
  NAND2_X1 U4333 ( .A1(n3416), .A2(n3415), .ZN(n3417) );
  NAND2_X1 U4334 ( .A1(n3419), .A2(n3550), .ZN(n3424) );
  NAND2_X1 U4335 ( .A1(n4548), .A2(n3420), .ZN(n3432) );
  OAI21_X1 U4336 ( .B1(n6580), .B2(n3421), .A(n3432), .ZN(n3422) );
  INV_X1 U4337 ( .A(n3422), .ZN(n3423) );
  NAND2_X1 U4338 ( .A1(n3424), .A2(n3423), .ZN(n6167) );
  NAND2_X1 U4339 ( .A1(n4446), .A2(n4447), .ZN(n4445) );
  INV_X1 U4340 ( .A(n3425), .ZN(n6168) );
  NAND2_X1 U4341 ( .A1(n6168), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3426)
         );
  NAND2_X1 U4342 ( .A1(n4502), .A2(n3550), .ZN(n3436) );
  OAI21_X1 U4343 ( .B1(n3431), .B2(n3430), .A(n3429), .ZN(n3434) );
  INV_X1 U4344 ( .A(n3432), .ZN(n3433) );
  AOI21_X1 U4345 ( .B1(n3434), .B2(n4335), .A(n3433), .ZN(n3435) );
  NAND2_X1 U4346 ( .A1(n3437), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6158)
         );
  NAND2_X1 U4347 ( .A1(n6157), .A2(n6158), .ZN(n3438) );
  NAND2_X1 U4348 ( .A1(n3438), .A2(n6159), .ZN(n4438) );
  NAND2_X1 U4349 ( .A1(n3439), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3440)
         );
  NAND2_X1 U4350 ( .A1(n4489), .A2(n4490), .ZN(n3443) );
  NAND2_X1 U4351 ( .A1(n3441), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3442)
         );
  NAND2_X1 U4352 ( .A1(n3443), .A2(n3442), .ZN(n4740) );
  NOR2_X2 U4353 ( .A1(n3446), .A2(n3445), .ZN(n3460) );
  NAND2_X1 U4354 ( .A1(n3569), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3458) );
  AOI22_X1 U4355 ( .A1(n4062), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4356 ( .A1(n3027), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4357 ( .A1(n2991), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3448) );
  AOI22_X1 U4358 ( .A1(n4084), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3447) );
  NAND4_X1 U4359 ( .A1(n3450), .A2(n3449), .A3(n3448), .A4(n3447), .ZN(n3456)
         );
  AOI22_X1 U4360 ( .A1(n3023), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3334), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4361 ( .A1(n3721), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3453) );
  AOI22_X1 U4362 ( .A1(n3307), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3452) );
  AOI22_X1 U4363 ( .A1(n4067), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3451) );
  NAND4_X1 U4364 ( .A1(n3454), .A2(n3453), .A3(n3452), .A4(n3451), .ZN(n3455)
         );
  INV_X1 U4365 ( .A(n3550), .ZN(n3467) );
  OR2_X1 U4366 ( .A1(n3463), .A2(n3462), .ZN(n3490) );
  XNOR2_X1 U4367 ( .A(n3490), .B(n3464), .ZN(n3465) );
  NAND2_X1 U4368 ( .A1(n3465), .A2(n4335), .ZN(n3466) );
  INV_X1 U4369 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3468) );
  NAND2_X1 U4370 ( .A1(n4740), .A2(n4739), .ZN(n3471) );
  NAND2_X1 U4371 ( .A1(n3469), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3470)
         );
  NAND2_X1 U4372 ( .A1(n3471), .A2(n3470), .ZN(n4722) );
  NAND2_X1 U4373 ( .A1(n3569), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3484) );
  AOI22_X1 U4374 ( .A1(n3721), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3475) );
  AOI22_X1 U4375 ( .A1(n4062), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3474) );
  AOI22_X1 U4376 ( .A1(n3334), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3473) );
  AOI22_X1 U4377 ( .A1(n4067), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3472) );
  NAND4_X1 U4378 ( .A1(n3475), .A2(n3474), .A3(n3473), .A4(n3472), .ZN(n3481)
         );
  AOI22_X1 U4379 ( .A1(n3023), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3479) );
  AOI22_X1 U4380 ( .A1(n3022), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3478) );
  AOI22_X1 U4381 ( .A1(n3307), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3477) );
  AOI22_X1 U4382 ( .A1(n4084), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3476) );
  NAND4_X1 U4383 ( .A1(n3479), .A2(n3478), .A3(n3477), .A4(n3476), .ZN(n3480)
         );
  INV_X1 U4384 ( .A(n3491), .ZN(n3482) );
  NAND2_X1 U4385 ( .A1(n3488), .A2(n3487), .ZN(n3659) );
  NAND3_X1 U4386 ( .A1(n3507), .A2(n3659), .A3(n3550), .ZN(n3494) );
  NOR2_X1 U4387 ( .A1(n3490), .A2(n3489), .ZN(n3492) );
  NAND2_X1 U4388 ( .A1(n3492), .A2(n3491), .ZN(n3512) );
  OAI211_X1 U4389 ( .C1(n3492), .C2(n3491), .A(n3512), .B(n4335), .ZN(n3493)
         );
  NAND2_X1 U4390 ( .A1(n3494), .A2(n3493), .ZN(n3495) );
  INV_X1 U4391 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4176) );
  NAND2_X1 U4392 ( .A1(n4722), .A2(n4723), .ZN(n3497) );
  NAND2_X1 U4393 ( .A1(n3495), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3496)
         );
  NAND2_X1 U4394 ( .A1(n3569), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3498) );
  OAI21_X1 U4395 ( .B1(n3499), .B2(n3594), .A(n3498), .ZN(n3500) );
  NAND2_X1 U4396 ( .A1(n3662), .A2(n3550), .ZN(n3503) );
  XNOR2_X1 U4397 ( .A(n3512), .B(n3510), .ZN(n3501) );
  NAND2_X1 U4398 ( .A1(n3501), .A2(n4335), .ZN(n3502) );
  NAND2_X1 U4399 ( .A1(n3503), .A2(n3502), .ZN(n3504) );
  NAND2_X1 U4400 ( .A1(n5195), .A2(n5196), .ZN(n3506) );
  NAND2_X1 U4401 ( .A1(n3504), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3505)
         );
  NAND2_X1 U4402 ( .A1(n3506), .A2(n3505), .ZN(n4960) );
  NAND2_X1 U4403 ( .A1(n4335), .A2(n3510), .ZN(n3511) );
  OR2_X1 U4404 ( .A1(n3512), .A2(n3511), .ZN(n3513) );
  INV_X1 U4405 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4182) );
  NAND2_X1 U4406 ( .A1(n3514), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3515)
         );
  INV_X1 U4407 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U4408 ( .A1(n3518), .A2(n6194), .ZN(n3516) );
  INV_X1 U4409 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3517) );
  NAND2_X1 U4410 ( .A1(n5621), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5166) );
  INV_X1 U4411 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3519) );
  NAND2_X1 U4412 ( .A1(n3518), .A2(n3519), .ZN(n5241) );
  NAND2_X1 U4413 ( .A1(n5621), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5242) );
  INV_X1 U4414 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3520) );
  NOR2_X1 U4415 ( .A1(n2992), .A2(n3520), .ZN(n5253) );
  NAND2_X1 U4416 ( .A1(n2992), .A2(n3520), .ZN(n5251) );
  OAI21_X1 U4417 ( .B1(n5250), .B2(n5253), .A(n5251), .ZN(n5294) );
  XNOR2_X1 U4418 ( .A(n2992), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5297)
         );
  NAND2_X1 U4419 ( .A1(n5294), .A2(n5297), .ZN(n5296) );
  INV_X1 U4420 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4284) );
  NAND2_X1 U4421 ( .A1(n2992), .A2(n4284), .ZN(n3521) );
  NAND2_X1 U4422 ( .A1(n5296), .A2(n3521), .ZN(n5646) );
  NAND2_X1 U4423 ( .A1(n5646), .A2(n3522), .ZN(n3524) );
  INV_X1 U4424 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U4425 ( .A1(n2992), .A2(n5906), .ZN(n3523) );
  NAND2_X1 U4426 ( .A1(n3524), .A2(n3523), .ZN(n5637) );
  XNOR2_X1 U4427 ( .A(n2992), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5638)
         );
  INV_X1 U4428 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U4429 ( .A1(n2992), .A2(n5893), .ZN(n3525) );
  INV_X1 U4430 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5774) );
  INV_X1 U4431 ( .A(n5618), .ZN(n3526) );
  NAND2_X1 U4432 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U4433 ( .A1(n3526), .A2(n3037), .ZN(n5585) );
  NAND2_X1 U4434 ( .A1(n5621), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5866) );
  OAI21_X1 U4435 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5621), .ZN(n3527) );
  AND2_X1 U4436 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5720) );
  AND2_X1 U4437 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4301) );
  AND2_X1 U4438 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5586) );
  NAND3_X1 U4439 ( .A1(n5720), .A2(n4301), .A3(n5586), .ZN(n3529) );
  NAND2_X1 U4440 ( .A1(n2992), .A2(n3529), .ZN(n3530) );
  NAND2_X1 U4441 ( .A1(n5752), .A2(n3530), .ZN(n3533) );
  NOR2_X1 U4442 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5719) );
  NOR2_X1 U4443 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5704) );
  NOR2_X1 U4444 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5741) );
  NAND3_X1 U4445 ( .A1(n5719), .A2(n5704), .A3(n5741), .ZN(n3531) );
  INV_X1 U4446 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5879) );
  NAND2_X1 U4447 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5676) );
  NOR2_X2 U4448 ( .A1(n5558), .A2(n5676), .ZN(n5541) );
  NAND2_X1 U4449 ( .A1(n5541), .A2(n3040), .ZN(n3538) );
  INV_X1 U4450 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5690) );
  INV_X1 U4451 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4255) );
  NAND2_X1 U4452 ( .A1(n5690), .A2(n4255), .ZN(n5677) );
  NOR3_X1 U4453 ( .A1(n2992), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n5677), 
        .ZN(n5359) );
  INV_X1 U4454 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5660) );
  INV_X1 U4455 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5669) );
  NAND3_X1 U4456 ( .A1(n5359), .A2(n5660), .A3(n5669), .ZN(n3536) );
  NAND2_X1 U4457 ( .A1(n3538), .A2(n3537), .ZN(n3539) );
  XNOR2_X1 U4458 ( .A(n3539), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4306)
         );
  OR2_X1 U4459 ( .A1(n3594), .A2(n4525), .ZN(n3540) );
  NAND2_X1 U4460 ( .A1(n3540), .A2(n3546), .ZN(n3554) );
  NAND2_X1 U4461 ( .A1(n6454), .A2(n3006), .ZN(n3542) );
  INV_X1 U4462 ( .A(n3560), .ZN(n3541) );
  XNOR2_X1 U4463 ( .A(n3561), .B(n3541), .ZN(n4136) );
  OAI21_X1 U4464 ( .B1(n3006), .B2(n6454), .A(n3542), .ZN(n3543) );
  NOR2_X1 U4465 ( .A1(n3594), .A2(n3543), .ZN(n3549) );
  INV_X1 U4466 ( .A(n3543), .ZN(n3544) );
  AOI21_X1 U4467 ( .B1(n3610), .B2(n3544), .A(n4548), .ZN(n3548) );
  NAND2_X1 U4468 ( .A1(n4525), .A2(n3546), .ZN(n3547) );
  NAND2_X1 U4469 ( .A1(n3545), .A2(n3547), .ZN(n3559) );
  OAI211_X1 U4470 ( .C1(n3554), .C2(n4136), .A(n3549), .B(n3553), .ZN(n3552)
         );
  NAND3_X1 U4471 ( .A1(n3554), .A2(STATE2_REG_0__SCAN_IN), .A3(n4136), .ZN(
        n3551) );
  NAND3_X1 U4472 ( .A1(n3552), .A2(n3600), .A3(n3551), .ZN(n3558) );
  INV_X1 U4473 ( .A(n3553), .ZN(n3556) );
  INV_X1 U4474 ( .A(n3554), .ZN(n3555) );
  NAND3_X1 U4475 ( .A1(n3556), .A2(n3555), .A3(n4136), .ZN(n3557) );
  NAND2_X1 U4476 ( .A1(n3558), .A2(n3557), .ZN(n3568) );
  INV_X1 U4477 ( .A(n3559), .ZN(n3570) );
  NAND2_X1 U4478 ( .A1(n3568), .A2(n3570), .ZN(n3567) );
  NAND2_X1 U4479 ( .A1(n3561), .A2(n3560), .ZN(n3563) );
  NAND2_X1 U4480 ( .A1(n5106), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3562) );
  NAND2_X1 U4481 ( .A1(n3563), .A2(n3562), .ZN(n3576) );
  MUX2_X1 U4482 ( .A(n4695), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n3575) );
  INV_X1 U4483 ( .A(n3575), .ZN(n3564) );
  XNOR2_X1 U4484 ( .A(n3576), .B(n3564), .ZN(n4134) );
  INV_X1 U4485 ( .A(n4134), .ZN(n3565) );
  NOR2_X1 U4486 ( .A1(n3594), .A2(n3565), .ZN(n3566) );
  NAND2_X1 U4487 ( .A1(n3567), .A2(n3566), .ZN(n3574) );
  INV_X1 U4488 ( .A(n3568), .ZN(n3572) );
  INV_X1 U4489 ( .A(n3569), .ZN(n3586) );
  OAI21_X1 U4490 ( .B1(n4134), .B2(n3586), .A(n3570), .ZN(n3571) );
  NAND2_X1 U4491 ( .A1(n3572), .A2(n3571), .ZN(n3573) );
  NAND2_X1 U4492 ( .A1(n3574), .A2(n3573), .ZN(n3589) );
  NAND2_X1 U4493 ( .A1(n3576), .A2(n3575), .ZN(n3578) );
  NAND2_X1 U4494 ( .A1(n4695), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3577) );
  NAND2_X1 U4495 ( .A1(n3578), .A2(n3577), .ZN(n3581) );
  INV_X1 U4496 ( .A(n3580), .ZN(n3579) );
  XNOR2_X1 U4497 ( .A(n3581), .B(n3579), .ZN(n3585) );
  NAND2_X1 U4498 ( .A1(n3581), .A2(n3580), .ZN(n3583) );
  NAND2_X1 U4499 ( .A1(n6468), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3582) );
  NAND2_X1 U4500 ( .A1(n3583), .A2(n3582), .ZN(n3590) );
  INV_X1 U4501 ( .A(n4135), .ZN(n3587) );
  NAND2_X1 U4502 ( .A1(n3587), .A2(n3586), .ZN(n3588) );
  NAND2_X1 U4503 ( .A1(n3589), .A2(n3588), .ZN(n3599) );
  NAND2_X1 U4504 ( .A1(n3590), .A2(n6234), .ZN(n3591) );
  INV_X1 U4505 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3640) );
  NAND2_X1 U4506 ( .A1(n3591), .A2(n3640), .ZN(n3593) );
  NOR2_X1 U4507 ( .A1(n3594), .A2(n4138), .ZN(n3595) );
  AOI21_X1 U4508 ( .B1(n6490), .B2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(n3595), 
        .ZN(n3596) );
  OAI21_X1 U4509 ( .B1(n3600), .B2(n4135), .A(n3596), .ZN(n3597) );
  INV_X1 U4510 ( .A(n3597), .ZN(n3598) );
  NAND2_X1 U4511 ( .A1(n3599), .A2(n3598), .ZN(n3604) );
  INV_X1 U4512 ( .A(n3600), .ZN(n3602) );
  INV_X1 U4513 ( .A(n4138), .ZN(n3601) );
  NAND2_X1 U4514 ( .A1(n3602), .A2(n3601), .ZN(n3603) );
  INV_X1 U4515 ( .A(n3218), .ZN(n3608) );
  NAND2_X1 U4516 ( .A1(n3219), .A2(n4150), .ZN(n3607) );
  NAND2_X1 U4517 ( .A1(n4376), .A2(n4548), .ZN(n3609) );
  NAND3_X1 U4518 ( .A1(n3606), .A2(n4269), .A3(n3609), .ZN(n4147) );
  NOR2_X2 U4519 ( .A1(n3612), .A2(n6481), .ZN(n3798) );
  AOI22_X1 U4520 ( .A1(n3623), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6481), .ZN(n3614) );
  AND2_X1 U4521 ( .A1(n5375), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3622) );
  NAND2_X1 U4522 ( .A1(n3622), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3613) );
  AND2_X1 U4523 ( .A1(n3614), .A2(n3613), .ZN(n3615) );
  AOI21_X1 U4524 ( .B1(n5097), .B2(n3616), .A(n6481), .ZN(n4458) );
  INV_X1 U4525 ( .A(n3798), .ZN(n3788) );
  AOI22_X1 U4526 ( .A1(n3623), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6481), .ZN(n3619) );
  NAND2_X1 U4527 ( .A1(n3622), .A2(n3006), .ZN(n3618) );
  AND2_X1 U4528 ( .A1(n3619), .A2(n3618), .ZN(n3620) );
  OAI21_X1 U4529 ( .B1(n3617), .B2(n3788), .A(n3620), .ZN(n4457) );
  NAND2_X1 U4530 ( .A1(n4458), .A2(n4457), .ZN(n4460) );
  OR2_X1 U4531 ( .A1(n4457), .A2(n3649), .ZN(n3621) );
  NAND2_X1 U4532 ( .A1(n4460), .A2(n3621), .ZN(n4419) );
  NAND2_X1 U4533 ( .A1(n6481), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3754) );
  INV_X1 U4534 ( .A(n3622), .ZN(n3641) );
  OAI21_X1 U4535 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3630), .ZN(n6165) );
  AOI22_X1 U4536 ( .A1(n4105), .A2(n6165), .B1(n4109), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3625) );
  INV_X2 U4537 ( .A(n3973), .ZN(n3902) );
  NAND2_X1 U4538 ( .A1(n3902), .A2(EAX_REG_2__SCAN_IN), .ZN(n3624) );
  OAI211_X1 U4539 ( .C1(n3641), .C2(n4385), .A(n3625), .B(n3624), .ZN(n4456)
         );
  NAND2_X1 U4540 ( .A1(n4454), .A2(n4456), .ZN(n3628) );
  NAND2_X1 U4541 ( .A1(n3626), .A2(n4416), .ZN(n3627) );
  NAND2_X1 U4542 ( .A1(n3629), .A2(n3798), .ZN(n3636) );
  OAI21_X1 U4543 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3631), .A(n3642), 
        .ZN(n6021) );
  AOI22_X1 U4544 ( .A1(n4105), .A2(n6021), .B1(n4109), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3633) );
  NAND2_X1 U4545 ( .A1(n3902), .A2(EAX_REG_3__SCAN_IN), .ZN(n3632) );
  OAI211_X1 U4546 ( .C1(n3641), .C2(n3359), .A(n3633), .B(n3632), .ZN(n3634)
         );
  INV_X1 U4547 ( .A(n3634), .ZN(n3635) );
  NAND2_X1 U4548 ( .A1(n3636), .A2(n3635), .ZN(n4466) );
  NAND2_X1 U4549 ( .A1(n4455), .A2(n4466), .ZN(n4461) );
  OAI21_X1 U4550 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n6656), .A(n6481), 
        .ZN(n3639) );
  NAND2_X1 U4551 ( .A1(n3902), .A2(EAX_REG_4__SCAN_IN), .ZN(n3638) );
  OAI211_X1 U4552 ( .C1(n3641), .C2(n3640), .A(n3639), .B(n3638), .ZN(n3644)
         );
  AOI21_X1 U4553 ( .B1(n3642), .B2(n6000), .A(n3648), .ZN(n5148) );
  NAND2_X1 U4554 ( .A1(n5148), .A2(n4105), .ZN(n3643) );
  AND2_X1 U4555 ( .A1(n3644), .A2(n3643), .ZN(n3645) );
  AOI21_X1 U4556 ( .B1(n3637), .B2(n3798), .A(n3645), .ZN(n4462) );
  AOI22_X1 U4557 ( .A1(n3902), .A2(EAX_REG_5__SCAN_IN), .B1(n4109), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3647) );
  OAI21_X1 U4558 ( .B1(n3648), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3653), 
        .ZN(n4987) );
  INV_X1 U4559 ( .A(n4987), .ZN(n5992) );
  NAND2_X1 U4560 ( .A1(n4463), .A2(n4560), .ZN(n4559) );
  INV_X1 U4561 ( .A(n4559), .ZN(n3661) );
  NAND2_X1 U4562 ( .A1(n3653), .A2(n3656), .ZN(n3655) );
  INV_X1 U4563 ( .A(n3663), .ZN(n3654) );
  NAND2_X1 U4564 ( .A1(n3655), .A2(n3654), .ZN(n5986) );
  INV_X1 U4565 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4904) );
  OAI22_X1 U4566 ( .A1(n3973), .A2(n4904), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3656), .ZN(n3657) );
  MUX2_X1 U4567 ( .A(n5986), .B(n3657), .S(n3649), .Z(n3658) );
  AOI21_X1 U4568 ( .B1(n3659), .B2(n3798), .A(n3658), .ZN(n4900) );
  NAND2_X1 U4569 ( .A1(n3661), .A2(n3660), .ZN(n4752) );
  INV_X1 U4570 ( .A(n4752), .ZN(n3733) );
  OAI21_X1 U4571 ( .B1(n3663), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3668), 
        .ZN(n5970) );
  NAND2_X1 U4572 ( .A1(n5970), .A2(n4105), .ZN(n3666) );
  NAND2_X1 U4573 ( .A1(n3902), .A2(EAX_REG_7__SCAN_IN), .ZN(n3665) );
  NAND2_X1 U4574 ( .A1(n4109), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3664)
         );
  XOR2_X1 U4575 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3716), .Z(n5180) );
  AOI22_X1 U4576 ( .A1(n3307), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4577 ( .A1(n4062), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4578 ( .A1(n2991), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4579 ( .A1(n4085), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3669) );
  NAND4_X1 U4580 ( .A1(n3672), .A2(n3671), .A3(n3670), .A4(n3669), .ZN(n3678)
         );
  AOI22_X1 U4581 ( .A1(n3023), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3334), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3676) );
  AOI22_X1 U4582 ( .A1(n3027), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4084), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3675) );
  AOI22_X1 U4583 ( .A1(n3721), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3674) );
  AOI22_X1 U4584 ( .A1(n4067), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3673) );
  NAND4_X1 U4585 ( .A1(n3676), .A2(n3675), .A3(n3674), .A4(n3673), .ZN(n3677)
         );
  OR2_X1 U4586 ( .A1(n3678), .A2(n3677), .ZN(n3679) );
  AOI22_X1 U4587 ( .A1(n3798), .A2(n3679), .B1(n4109), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3681) );
  NAND2_X1 U4588 ( .A1(n3902), .A2(EAX_REG_10__SCAN_IN), .ZN(n3680) );
  OAI211_X1 U4589 ( .C1(n5180), .C2(n3649), .A(n3681), .B(n3680), .ZN(n4975)
         );
  INV_X1 U4590 ( .A(n4975), .ZN(n3698) );
  XNOR2_X1 U4591 ( .A(n3683), .B(n3682), .ZN(n5202) );
  NAND2_X1 U4592 ( .A1(n5202), .A2(n4105), .ZN(n3697) );
  AOI22_X1 U4593 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n4062), .B1(n2991), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4594 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n3027), .B1(n4085), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4595 ( .A1(n4091), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4596 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n4084), .B1(n4092), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3684) );
  NAND4_X1 U4597 ( .A1(n3687), .A2(n3686), .A3(n3685), .A4(n3684), .ZN(n3693)
         );
  AOI22_X1 U4598 ( .A1(n3023), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4599 ( .A1(n3721), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4600 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(n3307), .B1(n3016), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4601 ( .A1(n3334), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3688) );
  NAND4_X1 U4602 ( .A1(n3691), .A2(n3690), .A3(n3689), .A4(n3688), .ZN(n3692)
         );
  OAI21_X1 U4603 ( .B1(n3693), .B2(n3692), .A(n3798), .ZN(n3696) );
  NAND2_X1 U4604 ( .A1(n3902), .A2(EAX_REG_9__SCAN_IN), .ZN(n3695) );
  NAND2_X1 U4605 ( .A1(n4109), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3694)
         );
  NAND2_X1 U4606 ( .A1(n3697), .A2(n3084), .ZN(n4951) );
  INV_X1 U4607 ( .A(n4951), .ZN(n4947) );
  XOR2_X1 U4608 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3699), .Z(n5956) );
  INV_X1 U4609 ( .A(n5956), .ZN(n5003) );
  AOI22_X1 U4610 ( .A1(n3022), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4611 ( .A1(n3027), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4084), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3702) );
  AOI22_X1 U4612 ( .A1(n3307), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3701) );
  AOI22_X1 U4613 ( .A1(n3274), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3700) );
  NAND4_X1 U4614 ( .A1(n3703), .A2(n3702), .A3(n3701), .A4(n3700), .ZN(n3709)
         );
  AOI22_X1 U4615 ( .A1(n3721), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3707) );
  AOI22_X1 U4616 ( .A1(n2991), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4617 ( .A1(n3334), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4618 ( .A1(n4062), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3704) );
  NAND4_X1 U4619 ( .A1(n3707), .A2(n3706), .A3(n3705), .A4(n3704), .ZN(n3708)
         );
  OAI21_X1 U4620 ( .B1(n3709), .B2(n3708), .A(n3798), .ZN(n3712) );
  NAND2_X1 U4621 ( .A1(n3902), .A2(EAX_REG_8__SCAN_IN), .ZN(n3711) );
  NAND2_X1 U4622 ( .A1(n4109), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3710)
         );
  NAND3_X1 U4623 ( .A1(n3712), .A2(n3711), .A3(n3710), .ZN(n3713) );
  AOI21_X1 U4624 ( .B1(n5003), .B2(n4105), .A(n3713), .ZN(n4994) );
  NOR2_X1 U4625 ( .A1(n3714), .A2(n4994), .ZN(n3715) );
  XNOR2_X1 U4626 ( .A(n3735), .B(n3734), .ZN(n5245) );
  NAND2_X1 U4627 ( .A1(n5245), .A2(n4105), .ZN(n3732) );
  AOI22_X1 U4628 ( .A1(n4062), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4629 ( .A1(n3307), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4630 ( .A1(n4091), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4631 ( .A1(n4084), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3717) );
  NAND4_X1 U4632 ( .A1(n3720), .A2(n3719), .A3(n3718), .A4(n3717), .ZN(n3727)
         );
  AOI22_X1 U4633 ( .A1(n3274), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3725) );
  AOI22_X1 U4634 ( .A1(n3022), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4635 ( .A1(n3721), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4636 ( .A1(n3334), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3722) );
  NAND4_X1 U4637 ( .A1(n3725), .A2(n3724), .A3(n3723), .A4(n3722), .ZN(n3726)
         );
  OAI21_X1 U4638 ( .B1(n3727), .B2(n3726), .A(n3798), .ZN(n3730) );
  NAND2_X1 U4639 ( .A1(n3902), .A2(EAX_REG_11__SCAN_IN), .ZN(n3729) );
  NAND2_X1 U4640 ( .A1(n4109), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3728)
         );
  AND3_X1 U4641 ( .A1(n3730), .A2(n3729), .A3(n3728), .ZN(n3731) );
  NAND2_X1 U4642 ( .A1(n3732), .A2(n3731), .ZN(n4908) );
  XOR2_X1 U4643 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3753), .Z(n5946) );
  INV_X1 U4644 ( .A(n5946), .ZN(n5256) );
  INV_X1 U4645 ( .A(EAX_REG_12__SCAN_IN), .ZN(n3737) );
  INV_X1 U4646 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3736) );
  OAI22_X1 U4647 ( .A1(n3973), .A2(n3737), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3736), .ZN(n3738) );
  NAND2_X1 U4648 ( .A1(n3738), .A2(n3649), .ZN(n3750) );
  AOI22_X1 U4649 ( .A1(n4062), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4650 ( .A1(n4085), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4084), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3741) );
  AOI22_X1 U4651 ( .A1(n3721), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4652 ( .A1(n4091), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3739) );
  NAND4_X1 U4653 ( .A1(n3742), .A2(n3741), .A3(n3740), .A4(n3739), .ZN(n3748)
         );
  AOI22_X1 U4654 ( .A1(n3274), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3746) );
  AOI22_X1 U4655 ( .A1(n3307), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3745) );
  AOI22_X1 U4656 ( .A1(n3334), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3744) );
  AOI22_X1 U4657 ( .A1(n3027), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3743) );
  NAND4_X1 U4658 ( .A1(n3746), .A2(n3745), .A3(n3744), .A4(n3743), .ZN(n3747)
         );
  OAI21_X1 U4659 ( .B1(n3748), .B2(n3747), .A(n3798), .ZN(n3749) );
  NAND2_X1 U4660 ( .A1(n3750), .A2(n3749), .ZN(n3751) );
  AOI21_X1 U4661 ( .B1(n5256), .B2(n4105), .A(n3751), .ZN(n5013) );
  INV_X1 U4662 ( .A(n5013), .ZN(n3752) );
  XNOR2_X1 U4663 ( .A(n3784), .B(n3783), .ZN(n5932) );
  NAND2_X1 U4664 ( .A1(n5932), .A2(n4105), .ZN(n3757) );
  NOR2_X1 U4665 ( .A1(n3754), .A2(n3783), .ZN(n3755) );
  AOI21_X1 U4666 ( .B1(n3902), .B2(EAX_REG_13__SCAN_IN), .A(n3755), .ZN(n3756)
         );
  NAND2_X1 U4667 ( .A1(n3757), .A2(n3756), .ZN(n3770) );
  AOI22_X1 U4668 ( .A1(n3721), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4669 ( .A1(n3274), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4670 ( .A1(n4062), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4084), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3759) );
  AOI22_X1 U4671 ( .A1(n4067), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3758) );
  NAND4_X1 U4672 ( .A1(n3761), .A2(n3760), .A3(n3759), .A4(n3758), .ZN(n3767)
         );
  AOI22_X1 U4673 ( .A1(n2991), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4674 ( .A1(n3334), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3764) );
  AOI22_X1 U4675 ( .A1(n4090), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4676 ( .A1(n3027), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3762) );
  NAND4_X1 U4677 ( .A1(n3765), .A2(n3764), .A3(n3763), .A4(n3762), .ZN(n3766)
         );
  OR2_X1 U4678 ( .A1(n3767), .A2(n3766), .ZN(n3768) );
  AND2_X1 U4679 ( .A1(n3798), .A2(n3768), .ZN(n5215) );
  NAND2_X1 U4680 ( .A1(n5214), .A2(n5215), .ZN(n3772) );
  NAND2_X1 U4681 ( .A1(n5012), .A2(n3770), .ZN(n3771) );
  AOI22_X1 U4682 ( .A1(n4062), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4683 ( .A1(n3027), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4084), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4684 ( .A1(n3721), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4685 ( .A1(n3334), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3773) );
  NAND4_X1 U4686 ( .A1(n3776), .A2(n3775), .A3(n3774), .A4(n3773), .ZN(n3782)
         );
  AOI22_X1 U4687 ( .A1(n2991), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4688 ( .A1(n3307), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4689 ( .A1(n3022), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4690 ( .A1(n3274), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3777) );
  NAND4_X1 U4691 ( .A1(n3780), .A2(n3779), .A3(n3778), .A4(n3777), .ZN(n3781)
         );
  NOR2_X1 U4692 ( .A1(n3782), .A2(n3781), .ZN(n3787) );
  XNOR2_X1 U4693 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3789), .ZN(n5650)
         );
  AOI22_X1 U4694 ( .A1(n4105), .A2(n5650), .B1(n4109), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3786) );
  NAND2_X1 U4695 ( .A1(n3902), .A2(EAX_REG_14__SCAN_IN), .ZN(n3785) );
  OAI211_X1 U4696 ( .C1(n3788), .C2(n3787), .A(n3786), .B(n3785), .ZN(n5185)
         );
  NAND2_X1 U4697 ( .A1(n5183), .A2(n5185), .ZN(n5184) );
  XOR2_X1 U4698 ( .A(n3806), .B(n3807), .Z(n5641) );
  INV_X1 U4699 ( .A(n5641), .ZN(n5230) );
  AOI22_X1 U4700 ( .A1(n4062), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4701 ( .A1(n3274), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4702 ( .A1(n4090), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4703 ( .A1(n4085), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3790) );
  NAND4_X1 U4704 ( .A1(n3793), .A2(n3792), .A3(n3791), .A4(n3790), .ZN(n3800)
         );
  AOI22_X1 U4705 ( .A1(n3721), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4706 ( .A1(n3334), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4707 ( .A1(n3027), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4084), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4708 ( .A1(n3016), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3794) );
  NAND4_X1 U4709 ( .A1(n3797), .A2(n3796), .A3(n3795), .A4(n3794), .ZN(n3799)
         );
  OAI21_X1 U4710 ( .B1(n3800), .B2(n3799), .A(n3798), .ZN(n3803) );
  NAND2_X1 U4711 ( .A1(n3902), .A2(EAX_REG_15__SCAN_IN), .ZN(n3802) );
  NAND2_X1 U4712 ( .A1(n4109), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3801)
         );
  NAND3_X1 U4713 ( .A1(n3803), .A2(n3802), .A3(n3801), .ZN(n3804) );
  AOI21_X1 U4714 ( .B1(n5230), .B2(n4105), .A(n3804), .ZN(n5223) );
  XNOR2_X1 U4715 ( .A(n3835), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5634)
         );
  AOI22_X1 U4716 ( .A1(n4062), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4717 ( .A1(n3027), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4084), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4718 ( .A1(n3274), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4719 ( .A1(n3307), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3808) );
  NAND4_X1 U4720 ( .A1(n3811), .A2(n3810), .A3(n3809), .A4(n3808), .ZN(n3817)
         );
  AOI22_X1 U4721 ( .A1(n3334), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4722 ( .A1(n3721), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4723 ( .A1(n3016), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4724 ( .A1(n3022), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3812) );
  NAND4_X1 U4725 ( .A1(n3815), .A2(n3814), .A3(n3813), .A4(n3812), .ZN(n3816)
         );
  NOR2_X1 U4726 ( .A1(n3817), .A2(n3816), .ZN(n3819) );
  AOI22_X1 U4727 ( .A1(n3902), .A2(EAX_REG_16__SCAN_IN), .B1(n4109), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3818) );
  OAI21_X1 U4728 ( .B1(n4078), .B2(n3819), .A(n3818), .ZN(n3820) );
  AOI21_X1 U4729 ( .B1(n5634), .B2(n4105), .A(n3820), .ZN(n5267) );
  AOI22_X1 U4730 ( .A1(n4062), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4731 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(n4084), .B1(n4085), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4732 ( .A1(n3307), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4733 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n4091), .B1(n4067), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3821) );
  NAND4_X1 U4734 ( .A1(n3824), .A2(n3823), .A3(n3822), .A4(n3821), .ZN(n3830)
         );
  AOI22_X1 U4735 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n2991), .B1(n3274), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4736 ( .A1(n3721), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4737 ( .A1(n3334), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4738 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(n3027), .B1(n4092), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3825) );
  NAND4_X1 U4739 ( .A1(n3828), .A2(n3827), .A3(n3826), .A4(n3825), .ZN(n3829)
         );
  NOR2_X1 U4740 ( .A1(n3830), .A2(n3829), .ZN(n3834) );
  NAND2_X1 U4741 ( .A1(n6481), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3831)
         );
  NAND2_X1 U4742 ( .A1(n3649), .A2(n3831), .ZN(n3832) );
  AOI21_X1 U4743 ( .B1(n3902), .B2(EAX_REG_17__SCAN_IN), .A(n3832), .ZN(n3833)
         );
  OAI21_X1 U4744 ( .B1(n4078), .B2(n3834), .A(n3833), .ZN(n3838) );
  OAI21_X1 U4745 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3836), .A(n3870), 
        .ZN(n5873) );
  OR2_X1 U4746 ( .A1(n3649), .A2(n5873), .ZN(n3837) );
  INV_X1 U4747 ( .A(n5279), .ZN(n3855) );
  AOI22_X1 U4748 ( .A1(n4062), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4749 ( .A1(n3027), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4750 ( .A1(n2991), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4751 ( .A1(n4084), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3839) );
  NAND4_X1 U4752 ( .A1(n3842), .A2(n3841), .A3(n3840), .A4(n3839), .ZN(n3848)
         );
  AOI22_X1 U4753 ( .A1(n3274), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3334), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4754 ( .A1(n3721), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4755 ( .A1(n3307), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4756 ( .A1(n4067), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3843) );
  NAND4_X1 U4757 ( .A1(n3846), .A2(n3845), .A3(n3844), .A4(n3843), .ZN(n3847)
         );
  NOR2_X1 U4758 ( .A1(n3848), .A2(n3847), .ZN(n3851) );
  AOI21_X1 U4759 ( .B1(n5624), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3849) );
  AOI21_X1 U4760 ( .B1(n3902), .B2(EAX_REG_18__SCAN_IN), .A(n3849), .ZN(n3850)
         );
  OAI21_X1 U4761 ( .B1(n4078), .B2(n3851), .A(n3850), .ZN(n3853) );
  XNOR2_X1 U4762 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3870), .ZN(n5626)
         );
  NAND2_X1 U4763 ( .A1(n4105), .A2(n5626), .ZN(n3852) );
  NAND2_X1 U4764 ( .A1(n3853), .A2(n3852), .ZN(n5468) );
  NAND2_X1 U4765 ( .A1(n3855), .A2(n3854), .ZN(n5465) );
  AOI22_X1 U4766 ( .A1(n4062), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4767 ( .A1(n4085), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4084), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4768 ( .A1(n3721), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4769 ( .A1(n4091), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3856) );
  NAND4_X1 U4770 ( .A1(n3859), .A2(n3858), .A3(n3857), .A4(n3856), .ZN(n3865)
         );
  AOI22_X1 U4771 ( .A1(n3274), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4772 ( .A1(n3307), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4773 ( .A1(n3027), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4774 ( .A1(n3334), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3860) );
  NAND4_X1 U4775 ( .A1(n3863), .A2(n3862), .A3(n3861), .A4(n3860), .ZN(n3864)
         );
  NOR2_X1 U4776 ( .A1(n3865), .A2(n3864), .ZN(n3869) );
  NAND2_X1 U4777 ( .A1(n6481), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3866)
         );
  NAND2_X1 U4778 ( .A1(n3649), .A2(n3866), .ZN(n3867) );
  AOI21_X1 U4779 ( .B1(n3902), .B2(EAX_REG_19__SCAN_IN), .A(n3867), .ZN(n3868)
         );
  OAI21_X1 U4780 ( .B1(n4078), .B2(n3869), .A(n3868), .ZN(n3873) );
  OAI21_X1 U4781 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n3871), .A(n3905), 
        .ZN(n5865) );
  OR2_X1 U4782 ( .A1(n3649), .A2(n5865), .ZN(n3872) );
  NAND2_X1 U4783 ( .A1(n3873), .A2(n3872), .ZN(n5512) );
  AOI22_X1 U4784 ( .A1(n4062), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4785 ( .A1(n4085), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4084), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4786 ( .A1(n3334), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4787 ( .A1(n3307), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3874) );
  NAND4_X1 U4788 ( .A1(n3877), .A2(n3876), .A3(n3875), .A4(n3874), .ZN(n3883)
         );
  AOI22_X1 U4789 ( .A1(n3274), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4790 ( .A1(n3721), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4791 ( .A1(n4067), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4792 ( .A1(n3027), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3878) );
  NAND4_X1 U4793 ( .A1(n3881), .A2(n3880), .A3(n3879), .A4(n3878), .ZN(n3882)
         );
  NOR2_X1 U4794 ( .A1(n3883), .A2(n3882), .ZN(n3887) );
  NAND2_X1 U4795 ( .A1(n6481), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3884)
         );
  NAND2_X1 U4796 ( .A1(n3649), .A2(n3884), .ZN(n3885) );
  AOI21_X1 U4797 ( .B1(n3902), .B2(EAX_REG_20__SCAN_IN), .A(n3885), .ZN(n3886)
         );
  OAI21_X1 U4798 ( .B1(n4078), .B2(n3887), .A(n3886), .ZN(n3889) );
  XNOR2_X1 U4799 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n3905), .ZN(n5616)
         );
  NAND2_X1 U4800 ( .A1(n5616), .A2(n4105), .ZN(n3888) );
  AOI22_X1 U4801 ( .A1(n2991), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4802 ( .A1(n4062), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4803 ( .A1(n3721), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4804 ( .A1(n3274), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3890) );
  NAND4_X1 U4805 ( .A1(n3893), .A2(n3892), .A3(n3891), .A4(n3890), .ZN(n3899)
         );
  AOI22_X1 U4806 ( .A1(n3307), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4807 ( .A1(n3027), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4808 ( .A1(n3334), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4809 ( .A1(n4084), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3894) );
  NAND4_X1 U4810 ( .A1(n3897), .A2(n3896), .A3(n3895), .A4(n3894), .ZN(n3898)
         );
  NOR2_X1 U4811 ( .A1(n3899), .A2(n3898), .ZN(n3904) );
  NAND2_X1 U4812 ( .A1(n6481), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3900)
         );
  NAND2_X1 U4813 ( .A1(n3649), .A2(n3900), .ZN(n3901) );
  AOI21_X1 U4814 ( .B1(n3902), .B2(EAX_REG_21__SCAN_IN), .A(n3901), .ZN(n3903)
         );
  OAI21_X1 U4815 ( .B1(n4078), .B2(n3904), .A(n3903), .ZN(n3909) );
  OAI21_X1 U4816 ( .B1(n3907), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n3950), 
        .ZN(n5608) );
  OR2_X1 U4817 ( .A1(n5608), .A2(n3649), .ZN(n3908) );
  AOI22_X1 U4818 ( .A1(n3334), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4819 ( .A1(n3022), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4820 ( .A1(n3721), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4821 ( .A1(n4084), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3910) );
  NAND4_X1 U4822 ( .A1(n3913), .A2(n3912), .A3(n3911), .A4(n3910), .ZN(n3919)
         );
  AOI22_X1 U4823 ( .A1(n3307), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4824 ( .A1(n4062), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4825 ( .A1(n3274), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4826 ( .A1(n3016), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3914) );
  NAND4_X1 U4827 ( .A1(n3917), .A2(n3916), .A3(n3915), .A4(n3914), .ZN(n3918)
         );
  NOR2_X1 U4828 ( .A1(n3919), .A2(n3918), .ZN(n3922) );
  INV_X1 U4829 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5600) );
  OAI21_X1 U4830 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5600), .A(n3649), .ZN(
        n3920) );
  AOI21_X1 U4831 ( .B1(n3902), .B2(EAX_REG_22__SCAN_IN), .A(n3920), .ZN(n3921)
         );
  OAI21_X1 U4832 ( .B1(n4078), .B2(n3922), .A(n3921), .ZN(n3924) );
  XNOR2_X1 U4833 ( .A(n3950), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5810)
         );
  NAND2_X1 U4834 ( .A1(n5810), .A2(n4105), .ZN(n3923) );
  NAND2_X1 U4835 ( .A1(n3924), .A2(n3923), .ZN(n5506) );
  AOI22_X1 U4836 ( .A1(n3721), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4837 ( .A1(n3016), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4838 ( .A1(n3027), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4839 ( .A1(n3334), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3926) );
  NAND4_X1 U4840 ( .A1(n3929), .A2(n3928), .A3(n3927), .A4(n3926), .ZN(n3935)
         );
  AOI22_X1 U4841 ( .A1(n3307), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3274), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4842 ( .A1(n4062), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4843 ( .A1(n4085), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4084), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4844 ( .A1(n2991), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3930) );
  NAND4_X1 U4845 ( .A1(n3933), .A2(n3932), .A3(n3931), .A4(n3930), .ZN(n3934)
         );
  NOR2_X1 U4846 ( .A1(n3935), .A2(n3934), .ZN(n3957) );
  AOI22_X1 U4847 ( .A1(n4062), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4848 ( .A1(n3274), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3938) );
  AOI22_X1 U4849 ( .A1(n4090), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4850 ( .A1(n4084), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3936) );
  NAND4_X1 U4851 ( .A1(n3939), .A2(n3938), .A3(n3937), .A4(n3936), .ZN(n3945)
         );
  AOI22_X1 U4852 ( .A1(n3721), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4853 ( .A1(n3334), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4854 ( .A1(n3022), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4855 ( .A1(n4067), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3940) );
  NAND4_X1 U4856 ( .A1(n3943), .A2(n3942), .A3(n3941), .A4(n3940), .ZN(n3944)
         );
  NOR2_X1 U4857 ( .A1(n3945), .A2(n3944), .ZN(n3958) );
  XNOR2_X1 U4858 ( .A(n3957), .B(n3958), .ZN(n3949) );
  NAND2_X1 U4859 ( .A1(n6481), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3946)
         );
  NAND2_X1 U4860 ( .A1(n3649), .A2(n3946), .ZN(n3947) );
  AOI21_X1 U4861 ( .B1(n3902), .B2(EAX_REG_23__SCAN_IN), .A(n3947), .ZN(n3948)
         );
  OAI21_X1 U4862 ( .B1(n4078), .B2(n3949), .A(n3948), .ZN(n3955) );
  NOR2_X1 U4863 ( .A1(n3951), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3952)
         );
  OR2_X1 U4864 ( .A1(n3992), .A2(n3952), .ZN(n5593) );
  INV_X1 U4865 ( .A(n5593), .ZN(n3953) );
  NAND2_X1 U4866 ( .A1(n3953), .A2(n4105), .ZN(n3954) );
  NAND2_X1 U4867 ( .A1(n3955), .A2(n3954), .ZN(n5427) );
  NOR2_X1 U4868 ( .A1(n3958), .A2(n3957), .ZN(n3987) );
  AOI22_X1 U4869 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n4062), .B1(n3022), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4870 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n3027), .B1(n4085), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4871 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n2991), .B1(n4091), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4872 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4084), .B1(n4092), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3959) );
  NAND4_X1 U4873 ( .A1(n3962), .A2(n3961), .A3(n3960), .A4(n3959), .ZN(n3968)
         );
  AOI22_X1 U4874 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n3334), .B1(n3274), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3966) );
  AOI22_X1 U4875 ( .A1(n3721), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U4876 ( .A1(n3307), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U4877 ( .A1(n4067), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3963) );
  NAND4_X1 U4878 ( .A1(n3966), .A2(n3965), .A3(n3964), .A4(n3963), .ZN(n3967)
         );
  OR2_X1 U4879 ( .A1(n3968), .A2(n3967), .ZN(n3986) );
  INV_X1 U4880 ( .A(n3986), .ZN(n3969) );
  XNOR2_X1 U4881 ( .A(n3987), .B(n3969), .ZN(n3975) );
  INV_X1 U4882 ( .A(n4078), .ZN(n4101) );
  INV_X1 U4883 ( .A(EAX_REG_24__SCAN_IN), .ZN(n3972) );
  NAND2_X1 U4884 ( .A1(n4109), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3971)
         );
  XNOR2_X1 U4885 ( .A(n3992), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5581)
         );
  NAND2_X1 U4886 ( .A1(n5581), .A2(n4105), .ZN(n3970) );
  OAI211_X1 U4887 ( .C1(n3973), .C2(n3972), .A(n3971), .B(n3970), .ZN(n3974)
         );
  AOI21_X1 U4888 ( .B1(n3975), .B2(n4101), .A(n3974), .ZN(n5415) );
  AOI22_X1 U4889 ( .A1(n3721), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4890 ( .A1(n4085), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4891 ( .A1(n4067), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4892 ( .A1(n4084), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3976) );
  NAND4_X1 U4893 ( .A1(n3979), .A2(n3978), .A3(n3977), .A4(n3976), .ZN(n3985)
         );
  AOI22_X1 U4894 ( .A1(n3274), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3334), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4895 ( .A1(n2991), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4896 ( .A1(n4062), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4897 ( .A1(n3307), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3980) );
  NAND4_X1 U4898 ( .A1(n3983), .A2(n3982), .A3(n3981), .A4(n3980), .ZN(n3984)
         );
  NOR2_X1 U4899 ( .A1(n3985), .A2(n3984), .ZN(n3999) );
  NAND2_X1 U4900 ( .A1(n3987), .A2(n3986), .ZN(n3998) );
  XNOR2_X1 U4901 ( .A(n3999), .B(n3998), .ZN(n3991) );
  NAND2_X1 U4902 ( .A1(n6481), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3988)
         );
  NAND2_X1 U4903 ( .A1(n3649), .A2(n3988), .ZN(n3989) );
  AOI21_X1 U4904 ( .B1(n3902), .B2(EAX_REG_25__SCAN_IN), .A(n3989), .ZN(n3990)
         );
  OAI21_X1 U4905 ( .B1(n3991), .B2(n4078), .A(n3990), .ZN(n3997) );
  OR2_X1 U4906 ( .A1(n3993), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3994)
         );
  NAND2_X1 U4907 ( .A1(n3994), .A2(n4033), .ZN(n5861) );
  INV_X1 U4908 ( .A(n5861), .ZN(n3995) );
  NAND2_X1 U4909 ( .A1(n3995), .A2(n4105), .ZN(n3996) );
  NOR2_X1 U4910 ( .A1(n3999), .A2(n3998), .ZN(n4028) );
  AOI22_X1 U4911 ( .A1(n4062), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U4912 ( .A1(n3027), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4913 ( .A1(n2991), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U4914 ( .A1(n4084), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4000) );
  NAND4_X1 U4915 ( .A1(n4003), .A2(n4002), .A3(n4001), .A4(n4000), .ZN(n4009)
         );
  AOI22_X1 U4916 ( .A1(n3274), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3334), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4917 ( .A1(n3721), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4918 ( .A1(n3307), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4005) );
  AOI22_X1 U4919 ( .A1(n4067), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4004) );
  NAND4_X1 U4920 ( .A1(n4007), .A2(n4006), .A3(n4005), .A4(n4004), .ZN(n4008)
         );
  OR2_X1 U4921 ( .A1(n4009), .A2(n4008), .ZN(n4027) );
  INV_X1 U4922 ( .A(n4027), .ZN(n4010) );
  XNOR2_X1 U4923 ( .A(n4028), .B(n4010), .ZN(n4011) );
  NAND2_X1 U4924 ( .A1(n4011), .A2(n4101), .ZN(n4016) );
  NAND2_X1 U4925 ( .A1(n6481), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4012)
         );
  NAND2_X1 U4926 ( .A1(n3649), .A2(n4012), .ZN(n4013) );
  AOI21_X1 U4927 ( .B1(n3902), .B2(EAX_REG_26__SCAN_IN), .A(n4013), .ZN(n4015)
         );
  XNOR2_X1 U4928 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .B(n4033), .ZN(n5800)
         );
  AOI21_X1 U4929 ( .B1(n4016), .B2(n4015), .A(n4014), .ZN(n5490) );
  AOI22_X1 U4930 ( .A1(n3274), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U4931 ( .A1(n3328), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U4932 ( .A1(n3307), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U4933 ( .A1(n3334), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4017) );
  NAND4_X1 U4934 ( .A1(n4020), .A2(n4019), .A3(n4018), .A4(n4017), .ZN(n4026)
         );
  AOI22_X1 U4935 ( .A1(n2991), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U4936 ( .A1(n3721), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U4937 ( .A1(n4091), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U4938 ( .A1(n4084), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4021) );
  NAND4_X1 U4939 ( .A1(n4024), .A2(n4023), .A3(n4022), .A4(n4021), .ZN(n4025)
         );
  NOR2_X1 U4940 ( .A1(n4026), .A2(n4025), .ZN(n4039) );
  NAND2_X1 U4941 ( .A1(n4028), .A2(n4027), .ZN(n4038) );
  XNOR2_X1 U4942 ( .A(n4039), .B(n4038), .ZN(n4032) );
  NAND2_X1 U4943 ( .A1(n6481), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4029)
         );
  NAND2_X1 U4944 ( .A1(n3649), .A2(n4029), .ZN(n4030) );
  AOI21_X1 U4945 ( .B1(n3902), .B2(EAX_REG_27__SCAN_IN), .A(n4030), .ZN(n4031)
         );
  OAI21_X1 U4946 ( .B1(n4032), .B2(n4078), .A(n4031), .ZN(n4037) );
  INV_X1 U4947 ( .A(n4033), .ZN(n4034) );
  OAI21_X1 U4948 ( .B1(n4035), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n4057), 
        .ZN(n5794) );
  OR2_X1 U4949 ( .A1(n5794), .A2(n3649), .ZN(n4036) );
  NOR2_X1 U4950 ( .A1(n4039), .A2(n4038), .ZN(n4075) );
  AOI22_X1 U4951 ( .A1(n3328), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U4952 ( .A1(n3027), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U4953 ( .A1(n2991), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U4954 ( .A1(n4084), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4040) );
  NAND4_X1 U4955 ( .A1(n4043), .A2(n4042), .A3(n4041), .A4(n4040), .ZN(n4049)
         );
  AOI22_X1 U4956 ( .A1(n3274), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3334), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U4957 ( .A1(n3721), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U4958 ( .A1(n3307), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U4959 ( .A1(n4067), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4044) );
  NAND4_X1 U4960 ( .A1(n4047), .A2(n4046), .A3(n4045), .A4(n4044), .ZN(n4048)
         );
  OR2_X1 U4961 ( .A1(n4049), .A2(n4048), .ZN(n4074) );
  XNOR2_X1 U4962 ( .A(n4075), .B(n4074), .ZN(n4053) );
  NAND2_X1 U4963 ( .A1(n6481), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4050)
         );
  NAND2_X1 U4964 ( .A1(n3649), .A2(n4050), .ZN(n4051) );
  AOI21_X1 U4965 ( .B1(n3902), .B2(EAX_REG_28__SCAN_IN), .A(n4051), .ZN(n4052)
         );
  OAI21_X1 U4966 ( .B1(n4053), .B2(n4078), .A(n4052), .ZN(n4055) );
  XNOR2_X1 U4967 ( .A(n4057), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5786)
         );
  NAND2_X1 U4968 ( .A1(n5786), .A2(n4105), .ZN(n4054) );
  NAND2_X1 U4969 ( .A1(n4055), .A2(n4054), .ZN(n5479) );
  INV_X1 U4970 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4056) );
  INV_X1 U4971 ( .A(n4058), .ZN(n4060) );
  INV_X1 U4972 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4059) );
  NAND2_X1 U4973 ( .A1(n4060), .A2(n4059), .ZN(n4061) );
  NAND2_X1 U4974 ( .A1(n4117), .A2(n4061), .ZN(n5546) );
  AOI22_X1 U4975 ( .A1(n3307), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3334), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U4976 ( .A1(n4062), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U4977 ( .A1(n3721), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U4978 ( .A1(n4085), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4063) );
  NAND4_X1 U4979 ( .A1(n4066), .A2(n4065), .A3(n4064), .A4(n4063), .ZN(n4073)
         );
  AOI22_X1 U4980 ( .A1(n3027), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4084), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U4981 ( .A1(n3022), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4070) );
  AOI22_X1 U4982 ( .A1(n3016), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U4983 ( .A1(n3274), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4068) );
  NAND4_X1 U4984 ( .A1(n4071), .A2(n4070), .A3(n4069), .A4(n4068), .ZN(n4072)
         );
  NOR2_X1 U4985 ( .A1(n4073), .A2(n4072), .ZN(n4083) );
  NAND2_X1 U4986 ( .A1(n4075), .A2(n4074), .ZN(n4082) );
  XNOR2_X1 U4987 ( .A(n4083), .B(n4082), .ZN(n4079) );
  AOI21_X1 U4988 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6481), .A(n4105), 
        .ZN(n4077) );
  NAND2_X1 U4989 ( .A1(n3902), .A2(EAX_REG_29__SCAN_IN), .ZN(n4076) );
  OAI211_X1 U4990 ( .C1(n4079), .C2(n4078), .A(n4077), .B(n4076), .ZN(n4080)
         );
  OAI21_X1 U4991 ( .B1(n3649), .B2(n5546), .A(n4080), .ZN(n5316) );
  INV_X1 U4992 ( .A(n5316), .ZN(n4081) );
  AND2_X2 U4993 ( .A1(n5315), .A2(n4081), .ZN(n5366) );
  NOR2_X1 U4994 ( .A1(n4083), .A2(n4082), .ZN(n4100) );
  AOI22_X1 U4995 ( .A1(n3274), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3334), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U4996 ( .A1(n2991), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3022), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4088) );
  AOI22_X1 U4997 ( .A1(n4085), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4084), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4087) );
  AOI22_X1 U4998 ( .A1(n3721), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4086) );
  NAND4_X1 U4999 ( .A1(n4089), .A2(n4088), .A3(n4087), .A4(n4086), .ZN(n4098)
         );
  AOI22_X1 U5000 ( .A1(n3307), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4096) );
  AOI22_X1 U5001 ( .A1(n3328), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4095) );
  AOI22_X1 U5002 ( .A1(n4067), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3025), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4094) );
  AOI22_X1 U5003 ( .A1(n3027), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4093) );
  NAND4_X1 U5004 ( .A1(n4096), .A2(n4095), .A3(n4094), .A4(n4093), .ZN(n4097)
         );
  NOR2_X1 U5005 ( .A1(n4098), .A2(n4097), .ZN(n4099) );
  XNOR2_X1 U5006 ( .A(n4100), .B(n4099), .ZN(n4102) );
  NAND2_X1 U5007 ( .A1(n4102), .A2(n4101), .ZN(n4108) );
  NAND2_X1 U5008 ( .A1(n6481), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4103)
         );
  NAND2_X1 U5009 ( .A1(n3649), .A2(n4103), .ZN(n4104) );
  AOI21_X1 U5010 ( .B1(n3902), .B2(EAX_REG_30__SCAN_IN), .A(n4104), .ZN(n4107)
         );
  XNOR2_X1 U5011 ( .A(n4117), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5384)
         );
  AND2_X1 U5012 ( .A1(n5384), .A2(n4105), .ZN(n4106) );
  AOI21_X1 U5013 ( .B1(n4108), .B2(n4107), .A(n4106), .ZN(n5365) );
  NAND2_X1 U5014 ( .A1(n5366), .A2(n5365), .ZN(n4112) );
  AOI22_X1 U5015 ( .A1(n3902), .A2(EAX_REG_31__SCAN_IN), .B1(n4109), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4110) );
  NAND3_X1 U5016 ( .A1(n6490), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6499) );
  NAND2_X2 U5017 ( .A1(n6481), .A2(n6573), .ZN(n6586) );
  OR2_X2 U5018 ( .A1(n6499), .A2(n6586), .ZN(n6175) );
  NAND2_X1 U5019 ( .A1(n5528), .A2(n6162), .ZN(n4123) );
  NAND2_X1 U5020 ( .A1(n6587), .A2(n6586), .ZN(n4113) );
  NAND2_X1 U5021 ( .A1(n4113), .A2(n6490), .ZN(n4114) );
  NAND2_X1 U5022 ( .A1(n6490), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4116) );
  NAND2_X1 U5023 ( .A1(n6656), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4115) );
  AND2_X1 U5024 ( .A1(n4116), .A2(n4115), .ZN(n6170) );
  INV_X1 U5025 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5367) );
  INV_X1 U5026 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4118) );
  NAND2_X1 U5027 ( .A1(n6490), .A2(n6481), .ZN(n4314) );
  INV_X1 U5028 ( .A(n4314), .ZN(n6501) );
  AND2_X2 U5029 ( .A1(n5340), .A2(n6501), .ZN(n6215) );
  AND2_X1 U5030 ( .A1(n6215), .A2(REIP_REG_31__SCAN_IN), .ZN(n4296) );
  AOI21_X1 U5031 ( .B1(n6156), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n4296), 
        .ZN(n4120) );
  OAI21_X1 U5032 ( .B1(n6166), .B2(n4323), .A(n4120), .ZN(n4121) );
  INV_X1 U5033 ( .A(n4121), .ZN(n4122) );
  OAI211_X1 U5034 ( .C1(n4306), .C2(n5914), .A(n4123), .B(n4122), .ZN(U2955)
         );
  INV_X1 U5035 ( .A(n4125), .ZN(n4127) );
  INV_X1 U5036 ( .A(STATE_REG_0__SCAN_IN), .ZN(n4126) );
  NAND2_X1 U5037 ( .A1(n4127), .A2(n4126), .ZN(n6509) );
  NAND2_X1 U5038 ( .A1(n4525), .A2(n6509), .ZN(n4321) );
  NAND2_X1 U5039 ( .A1(n4321), .A2(n6728), .ZN(n4128) );
  OAI211_X1 U5040 ( .C1(n4124), .C2(n4128), .A(n4145), .B(n4271), .ZN(n4129)
         );
  NAND2_X1 U5041 ( .A1(n4129), .A2(n4537), .ZN(n4143) );
  NAND2_X1 U5042 ( .A1(n5334), .A2(n4268), .ZN(n4278) );
  INV_X1 U5043 ( .A(n4278), .ZN(n4130) );
  NAND2_X1 U5044 ( .A1(n5407), .A2(n4130), .ZN(n4140) );
  NOR2_X1 U5045 ( .A1(n3243), .A2(n4145), .ZN(n5405) );
  OAI21_X1 U5046 ( .B1(n4548), .B2(n3218), .A(n6580), .ZN(n4131) );
  OAI21_X1 U5047 ( .B1(n3238), .B2(n3218), .A(n4131), .ZN(n4132) );
  INV_X1 U5048 ( .A(n4132), .ZN(n4277) );
  NOR2_X1 U5049 ( .A1(n4277), .A2(n4147), .ZN(n4133) );
  OR2_X1 U5050 ( .A1(n5405), .A2(n4133), .ZN(n4364) );
  INV_X1 U5051 ( .A(n6509), .ZN(n5410) );
  NAND3_X1 U5052 ( .A1(n4136), .A2(n4135), .A3(n4134), .ZN(n4137) );
  NAND2_X1 U5053 ( .A1(n4138), .A2(n4137), .ZN(n5404) );
  NOR2_X1 U5054 ( .A1(READY_N), .A2(n5404), .ZN(n4359) );
  OAI211_X1 U5055 ( .C1(n4525), .C2(n5410), .A(n4272), .B(n4359), .ZN(n4139)
         );
  NAND3_X1 U5056 ( .A1(n4140), .A2(n4364), .A3(n4139), .ZN(n4141) );
  NAND2_X1 U5057 ( .A1(n4141), .A2(n6491), .ZN(n4142) );
  AND2_X4 U5058 ( .A1(n4145), .A2(n4268), .ZN(n4565) );
  OR2_X1 U5059 ( .A1(n4124), .A2(n5396), .ZN(n4423) );
  OAI211_X1 U5060 ( .C1(n4529), .C2(n4151), .A(n4144), .B(n4423), .ZN(n4146)
         );
  INV_X1 U5061 ( .A(n4146), .ZN(n4148) );
  INV_X1 U5062 ( .A(n6473), .ZN(n5403) );
  OR2_X1 U5063 ( .A1(n4147), .A2(n3545), .ZN(n5402) );
  NAND3_X1 U5064 ( .A1(n4148), .A2(n5403), .A3(n5402), .ZN(n4149) );
  OAI21_X1 U5065 ( .B1(n4151), .B2(n4150), .A(n6480), .ZN(n4152) );
  INV_X1 U5066 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4570) );
  INV_X1 U5067 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4153) );
  NAND2_X1 U5068 ( .A1(n4211), .A2(n4153), .ZN(n4155) );
  NAND2_X1 U5069 ( .A1(n4565), .A2(n4570), .ZN(n4154) );
  NAND3_X1 U5070 ( .A1(n4155), .A2(n4251), .A3(n4154), .ZN(n4156) );
  NAND2_X1 U5071 ( .A1(n4211), .A2(EBX_REG_0__SCAN_IN), .ZN(n4158) );
  INV_X1 U5072 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5209) );
  NAND2_X1 U5073 ( .A1(n4251), .A2(n5209), .ZN(n4157) );
  OAI21_X1 U5074 ( .B1(n4448), .B2(n5396), .A(n4159), .ZN(n4160) );
  INV_X1 U5075 ( .A(n4160), .ZN(n4574) );
  INV_X1 U5076 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4575) );
  NAND2_X1 U5077 ( .A1(n4161), .A2(n4575), .ZN(n4164) );
  NAND2_X1 U5078 ( .A1(n4165), .A2(n5396), .ZN(n4217) );
  INV_X1 U5079 ( .A(n4211), .ZN(n4165) );
  OR2_X1 U5080 ( .A1(n4211), .A2(n4575), .ZN(n4163) );
  NAND2_X1 U5081 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n5396), .ZN(n4162)
         );
  NAND4_X1 U5082 ( .A1(n4164), .A2(n4217), .A3(n4163), .A4(n4162), .ZN(n4573)
         );
  INV_X1 U5083 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4735) );
  NAND2_X1 U5084 ( .A1(n4234), .A2(n4735), .ZN(n4169) );
  NAND2_X1 U5085 ( .A1(n4565), .A2(n4735), .ZN(n4167) );
  NAND2_X1 U5086 ( .A1(n4275), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4166)
         );
  NAND3_X1 U5087 ( .A1(n4167), .A2(n4211), .A3(n4166), .ZN(n4168) );
  INV_X1 U5088 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4732) );
  NAND2_X1 U5089 ( .A1(n4161), .A2(n4732), .ZN(n4174) );
  NAND2_X1 U5090 ( .A1(n4211), .A2(n4170), .ZN(n4172) );
  NAND2_X1 U5091 ( .A1(n4565), .A2(n4732), .ZN(n4171) );
  NAND3_X1 U5092 ( .A1(n4172), .A2(n4275), .A3(n4171), .ZN(n4173) );
  NAND2_X1 U5093 ( .A1(n4174), .A2(n4173), .ZN(n4495) );
  MUX2_X1 U5094 ( .A(n4254), .B(n4275), .S(EBX_REG_5__SCAN_IN), .Z(n4175) );
  NAND2_X1 U5095 ( .A1(n4211), .A2(n4275), .ZN(n4561) );
  NAND2_X1 U5096 ( .A1(n4175), .A2(n3092), .ZN(n4577) );
  INV_X1 U5097 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4901) );
  NAND2_X1 U5098 ( .A1(n4161), .A2(n4901), .ZN(n4180) );
  NAND2_X1 U5099 ( .A1(n4211), .A2(n4176), .ZN(n4178) );
  NAND2_X1 U5100 ( .A1(n4565), .A2(n4901), .ZN(n4177) );
  NAND3_X1 U5101 ( .A1(n4178), .A2(n4275), .A3(n4177), .ZN(n4179) );
  NAND2_X1 U5102 ( .A1(n4180), .A2(n4179), .ZN(n4725) );
  MUX2_X1 U5103 ( .A(n4254), .B(n4275), .S(EBX_REG_7__SCAN_IN), .Z(n4181) );
  OAI21_X1 U5104 ( .B1(n4561), .B2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n4181), 
        .ZN(n4758) );
  INV_X1 U5105 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U5106 ( .A1(n4161), .A2(n5953), .ZN(n4186) );
  NAND2_X1 U5107 ( .A1(n4211), .A2(n4182), .ZN(n4184) );
  NAND2_X1 U5108 ( .A1(n4565), .A2(n5953), .ZN(n4183) );
  NAND3_X1 U5109 ( .A1(n4184), .A2(n4275), .A3(n4183), .ZN(n4185) );
  NAND2_X1 U5110 ( .A1(n4186), .A2(n4185), .ZN(n4967) );
  INV_X1 U5111 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4956) );
  NAND2_X1 U5112 ( .A1(n4234), .A2(n4956), .ZN(n4190) );
  NAND2_X1 U5113 ( .A1(n4565), .A2(n4956), .ZN(n4188) );
  NAND2_X1 U5114 ( .A1(n4251), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4187)
         );
  NAND3_X1 U5115 ( .A1(n4188), .A2(n4211), .A3(n4187), .ZN(n4189) );
  NAND2_X1 U5116 ( .A1(n4190), .A2(n4189), .ZN(n4953) );
  INV_X1 U5117 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4191) );
  NAND2_X1 U5118 ( .A1(n4161), .A2(n4191), .ZN(n4194) );
  OR2_X1 U5119 ( .A1(n4211), .A2(n4191), .ZN(n4193) );
  NAND2_X1 U5120 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n5396), .ZN(n4192) );
  NAND4_X1 U5121 ( .A1(n4194), .A2(n4217), .A3(n4193), .A4(n4192), .ZN(n4999)
         );
  INV_X1 U5122 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5079) );
  NAND2_X1 U5123 ( .A1(n4234), .A2(n5079), .ZN(n4198) );
  NAND2_X1 U5124 ( .A1(n4565), .A2(n5079), .ZN(n4196) );
  NAND2_X1 U5125 ( .A1(n4251), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4195) );
  NAND3_X1 U5126 ( .A1(n4196), .A2(n4211), .A3(n4195), .ZN(n4197) );
  NAND2_X1 U5127 ( .A1(n4198), .A2(n4197), .ZN(n4909) );
  INV_X1 U5128 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5017) );
  NAND2_X1 U5129 ( .A1(n4161), .A2(n5017), .ZN(n4201) );
  OR2_X1 U5130 ( .A1(n4211), .A2(n5017), .ZN(n4200) );
  NAND2_X1 U5131 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n5396), .ZN(n4199) );
  NAND4_X1 U5132 ( .A1(n4201), .A2(n4217), .A3(n4200), .A4(n4199), .ZN(n5015)
         );
  INV_X1 U5133 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5930) );
  NAND2_X1 U5134 ( .A1(n4234), .A2(n5930), .ZN(n4205) );
  NAND2_X1 U5135 ( .A1(n4565), .A2(n5930), .ZN(n4203) );
  NAND2_X1 U5136 ( .A1(n4251), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4202) );
  NAND3_X1 U5137 ( .A1(n4203), .A2(n4211), .A3(n4202), .ZN(n4204) );
  NAND2_X1 U5138 ( .A1(n4205), .A2(n4204), .ZN(n5218) );
  INV_X1 U5139 ( .A(EBX_REG_14__SCAN_IN), .ZN(n4206) );
  NAND2_X1 U5140 ( .A1(n4161), .A2(n4206), .ZN(n4209) );
  OR2_X1 U5141 ( .A1(n4211), .A2(n4206), .ZN(n4208) );
  NAND2_X1 U5142 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5396), .ZN(n4207) );
  NAND4_X1 U5143 ( .A1(n4209), .A2(n4217), .A3(n4208), .A4(n4207), .ZN(n5188)
         );
  INV_X1 U5144 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5236) );
  NAND2_X1 U5145 ( .A1(n4234), .A2(n5236), .ZN(n4214) );
  NAND2_X1 U5146 ( .A1(n4565), .A2(n5236), .ZN(n4212) );
  NAND2_X1 U5147 ( .A1(n4275), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4210) );
  NAND3_X1 U5148 ( .A1(n4212), .A2(n4211), .A3(n4210), .ZN(n4213) );
  NAND2_X1 U5149 ( .A1(n4214), .A2(n4213), .ZN(n5229) );
  NOR2_X2 U5150 ( .A1(n5227), .A2(n5229), .ZN(n5268) );
  INV_X1 U5151 ( .A(EBX_REG_16__SCAN_IN), .ZN(n4215) );
  NAND2_X1 U5152 ( .A1(n4161), .A2(n4215), .ZN(n4219) );
  OR2_X1 U5153 ( .A1(n4211), .A2(n4215), .ZN(n4218) );
  NAND2_X1 U5154 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n5396), .ZN(n4216) );
  NAND4_X1 U5155 ( .A1(n4219), .A2(n4218), .A3(n4217), .A4(n4216), .ZN(n5269)
         );
  AOI21_X1 U5156 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n4275), .A(n4165), 
        .ZN(n4220) );
  OAI21_X1 U5157 ( .B1(EBX_REG_17__SCAN_IN), .B2(n5396), .A(n4220), .ZN(n4221)
         );
  OAI21_X1 U5158 ( .B1(EBX_REG_17__SCAN_IN), .B2(n4254), .A(n4221), .ZN(n5287)
         );
  INV_X1 U5159 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U5160 ( .A1(n4161), .A2(n5830), .ZN(n4225) );
  INV_X1 U5161 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U5162 ( .A1(n4211), .A2(n5753), .ZN(n4223) );
  NAND2_X1 U5163 ( .A1(n4565), .A2(n5830), .ZN(n4222) );
  NAND3_X1 U5164 ( .A1(n4223), .A2(n4251), .A3(n4222), .ZN(n4224) );
  NAND2_X1 U5165 ( .A1(n4225), .A2(n4224), .ZN(n5516) );
  OR2_X1 U5166 ( .A1(n4561), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4227)
         );
  INV_X1 U5167 ( .A(EBX_REG_18__SCAN_IN), .ZN(n4226) );
  NAND2_X1 U5168 ( .A1(n4565), .A2(n4226), .ZN(n5472) );
  OR2_X1 U5169 ( .A1(n4561), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4229)
         );
  INV_X1 U5170 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5511) );
  NAND2_X1 U5171 ( .A1(n4565), .A2(n5511), .ZN(n4228) );
  NAND2_X1 U5172 ( .A1(n4229), .A2(n4228), .ZN(n5457) );
  NOR2_X1 U5173 ( .A1(n4275), .A2(n5511), .ZN(n4230) );
  AOI21_X1 U5174 ( .B1(n4231), .B2(n5457), .A(n4230), .ZN(n4233) );
  INV_X1 U5175 ( .A(n4231), .ZN(n5473) );
  NAND2_X1 U5176 ( .A1(n5473), .A2(n4275), .ZN(n4232) );
  INV_X1 U5177 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5508) );
  NAND2_X1 U5178 ( .A1(n4234), .A2(n5508), .ZN(n4237) );
  NAND2_X1 U5179 ( .A1(n4275), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4235) );
  OAI211_X1 U5180 ( .C1(n5396), .C2(EBX_REG_21__SCAN_IN), .A(n4211), .B(n4235), 
        .ZN(n4236) );
  AOI22_X1 U5181 ( .A1(n4165), .A2(EBX_REG_22__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5396), .ZN(n4240) );
  INV_X1 U5182 ( .A(EBX_REG_22__SCAN_IN), .ZN(n4238) );
  NAND2_X1 U5183 ( .A1(n4161), .A2(n4238), .ZN(n4239) );
  NAND2_X1 U5184 ( .A1(n4251), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4241) );
  OAI211_X1 U5185 ( .C1(n5396), .C2(EBX_REG_23__SCAN_IN), .A(n4211), .B(n4241), 
        .ZN(n4242) );
  OAI21_X1 U5186 ( .B1(n4254), .B2(EBX_REG_23__SCAN_IN), .A(n4242), .ZN(n5431)
         );
  AOI22_X1 U5187 ( .A1(n4165), .A2(EBX_REG_24__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n5396), .ZN(n4244) );
  INV_X1 U5188 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U5189 ( .A1(n4161), .A2(n5422), .ZN(n4243) );
  NAND2_X1 U5190 ( .A1(n4244), .A2(n4243), .ZN(n5416) );
  MUX2_X1 U5191 ( .A(n4254), .B(n4275), .S(EBX_REG_25__SCAN_IN), .Z(n4245) );
  OAI21_X1 U5192 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n4561), .A(n4245), 
        .ZN(n4246) );
  INV_X1 U5193 ( .A(n4246), .ZN(n4331) );
  INV_X1 U5194 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5809) );
  NAND2_X1 U5195 ( .A1(n4161), .A2(n5809), .ZN(n4250) );
  INV_X1 U5196 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U5197 ( .A1(n4211), .A2(n5551), .ZN(n4248) );
  NAND2_X1 U5198 ( .A1(n4565), .A2(n5809), .ZN(n4247) );
  NAND3_X1 U5199 ( .A1(n4248), .A2(n4251), .A3(n4247), .ZN(n4249) );
  AND2_X1 U5200 ( .A1(n4250), .A2(n4249), .ZN(n5491) );
  NAND2_X1 U5201 ( .A1(n4251), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4252) );
  OAI211_X1 U5202 ( .C1(n5396), .C2(EBX_REG_27__SCAN_IN), .A(n4211), .B(n4252), 
        .ZN(n4253) );
  OAI21_X1 U5203 ( .B1(n4254), .B2(EBX_REG_27__SCAN_IN), .A(n4253), .ZN(n5682)
         );
  INV_X1 U5204 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5485) );
  NAND2_X1 U5205 ( .A1(n4161), .A2(n5485), .ZN(n4259) );
  NAND2_X1 U5206 ( .A1(n4211), .A2(n4255), .ZN(n4257) );
  NAND2_X1 U5207 ( .A1(n4565), .A2(n5485), .ZN(n4256) );
  NAND3_X1 U5208 ( .A1(n4257), .A2(n4275), .A3(n4256), .ZN(n4258) );
  NAND2_X1 U5209 ( .A1(n4259), .A2(n4258), .ZN(n5482) );
  OAI22_X1 U5210 ( .A1(n4561), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n5396), .ZN(n5379) );
  INV_X1 U5211 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5477) );
  NOR2_X1 U5212 ( .A1(n4275), .A2(n5477), .ZN(n4262) );
  AOI21_X1 U5213 ( .B1(n5379), .B2(n4275), .A(n4262), .ZN(n5318) );
  AND2_X1 U5214 ( .A1(n5396), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4260)
         );
  AOI21_X1 U5215 ( .B1(n4561), .B2(EBX_REG_30__SCAN_IN), .A(n4260), .ZN(n5380)
         );
  INV_X1 U5216 ( .A(n5484), .ZN(n4261) );
  NAND2_X1 U5217 ( .A1(n4261), .A2(n5471), .ZN(n4264) );
  INV_X1 U5218 ( .A(n4262), .ZN(n4263) );
  OAI211_X1 U5219 ( .C1(n5320), .C2(n5380), .A(n4264), .B(n4263), .ZN(n4266)
         );
  OAI22_X1 U5220 ( .A1(n4561), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n5396), .ZN(n4265) );
  AND2_X1 U5221 ( .A1(n5405), .A2(n4268), .ZN(n4402) );
  NAND2_X1 U5222 ( .A1(n4285), .A2(n4402), .ZN(n6231) );
  AND2_X1 U5223 ( .A1(n4548), .A2(n4268), .ZN(n5087) );
  AND2_X1 U5224 ( .A1(n5087), .A2(n4537), .ZN(n4362) );
  INV_X1 U5225 ( .A(n4269), .ZN(n4270) );
  OAI21_X1 U5226 ( .B1(n4362), .B2(n4561), .A(n4270), .ZN(n4274) );
  NAND2_X1 U5227 ( .A1(n4272), .A2(n4271), .ZN(n4273) );
  OAI211_X1 U5228 ( .C1(n3606), .C2(n4275), .A(n4274), .B(n4273), .ZN(n4276)
         );
  NAND2_X1 U5229 ( .A1(n4285), .A2(n5400), .ZN(n5739) );
  INV_X1 U5230 ( .A(n4373), .ZN(n4279) );
  OAI211_X1 U5231 ( .C1(n4371), .C2(n4145), .A(n4279), .B(n4403), .ZN(n4280)
         );
  NAND2_X1 U5232 ( .A1(n4285), .A2(n4280), .ZN(n5897) );
  NAND2_X1 U5233 ( .A1(n5739), .A2(n5897), .ZN(n5303) );
  INV_X1 U5234 ( .A(n5303), .ZN(n4281) );
  NAND2_X1 U5235 ( .A1(n6231), .A2(n4281), .ZN(n5770) );
  AND2_X1 U5236 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U5237 ( .A1(n6231), .A2(n5897), .ZN(n5735) );
  INV_X1 U5238 ( .A(n6231), .ZN(n4282) );
  NOR2_X1 U5239 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n4282), .ZN(n4449)
         );
  INV_X1 U5240 ( .A(n4449), .ZN(n4283) );
  NAND2_X1 U5241 ( .A1(n5735), .A2(n4283), .ZN(n4743) );
  INV_X1 U5242 ( .A(n4743), .ZN(n6217) );
  NOR2_X1 U5243 ( .A1(n6217), .A2(n6209), .ZN(n4292) );
  INV_X1 U5244 ( .A(n5720), .ZN(n4300) );
  INV_X1 U5245 ( .A(n5735), .ZN(n4963) );
  NAND2_X1 U5246 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5305) );
  NOR2_X1 U5247 ( .A1(n4284), .A2(n5305), .ZN(n5895) );
  NAND2_X1 U5248 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5895), .ZN(n5771) );
  NAND2_X1 U5249 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5772) );
  NOR2_X1 U5250 ( .A1(n5771), .A2(n5772), .ZN(n4298) );
  INV_X1 U5251 ( .A(n4298), .ZN(n5734) );
  INV_X1 U5252 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6203) );
  NOR2_X1 U5253 ( .A1(n6203), .A2(n4182), .ZN(n5171) );
  INV_X1 U5254 ( .A(n5171), .ZN(n5168) );
  NAND2_X1 U5255 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5169) );
  NOR2_X1 U5256 ( .A1(n5168), .A2(n5169), .ZN(n4287) );
  NAND4_X1 U5257 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4742) );
  NOR3_X1 U5258 ( .A1(n3468), .A2(n4176), .A3(n4742), .ZN(n4962) );
  NAND2_X1 U5259 ( .A1(n4287), .A2(n4962), .ZN(n5736) );
  INV_X1 U5260 ( .A(n5756), .ZN(n5744) );
  NAND2_X1 U5261 ( .A1(n5744), .A2(n5586), .ZN(n4299) );
  NOR3_X1 U5262 ( .A1(n5734), .A2(n5736), .A3(n4299), .ZN(n4291) );
  OR2_X1 U5263 ( .A1(n5897), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4286)
         );
  OR2_X1 U5264 ( .A1(n4285), .A2(n6215), .ZN(n6230) );
  NAND2_X1 U5265 ( .A1(n4286), .A2(n6230), .ZN(n5733) );
  INV_X1 U5266 ( .A(n5733), .ZN(n4290) );
  INV_X1 U5267 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U5268 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U5269 ( .A1(n6216), .A2(n6207), .ZN(n6206) );
  NAND3_X1 U5270 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n6206), .ZN(n4744) );
  NOR2_X1 U5271 ( .A1(n3468), .A2(n4744), .ZN(n4727) );
  AND2_X1 U5272 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4727), .ZN(n4971)
         );
  NAND2_X1 U5273 ( .A1(n4971), .A2(n4287), .ZN(n4297) );
  NOR2_X1 U5274 ( .A1(n4297), .A2(n5734), .ZN(n5738) );
  INV_X1 U5275 ( .A(n5738), .ZN(n4288) );
  OAI21_X1 U5276 ( .B1(n4299), .B2(n4288), .A(n6209), .ZN(n4289) );
  OAI211_X1 U5277 ( .C1(n4963), .C2(n4291), .A(n4290), .B(n4289), .ZN(n5730)
         );
  AOI21_X1 U5278 ( .B1(n4300), .B2(n5770), .A(n5730), .ZN(n5712) );
  OAI21_X1 U5279 ( .B1(n4301), .B2(n4292), .A(n5712), .ZN(n5878) );
  INV_X1 U5280 ( .A(n5878), .ZN(n4293) );
  OAI21_X1 U5281 ( .B1(n5696), .B2(n5740), .A(n4293), .ZN(n5681) );
  AOI21_X1 U5282 ( .B1(n5676), .B2(n5770), .A(n5681), .ZN(n5664) );
  OAI21_X1 U5283 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5740), .A(n5664), 
        .ZN(n5655) );
  AOI21_X1 U5284 ( .B1(n5660), .B2(n5770), .A(n5655), .ZN(n4294) );
  INV_X1 U5285 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4379) );
  NOR2_X1 U5286 ( .A1(n4294), .A2(n4379), .ZN(n4295) );
  AOI211_X1 U5287 ( .C1(n6210), .C2(n5344), .A(n4296), .B(n4295), .ZN(n4304)
         );
  INV_X1 U5288 ( .A(n4297), .ZN(n5260) );
  NAND2_X1 U5289 ( .A1(n6209), .A2(n5260), .ZN(n5896) );
  NAND2_X1 U5290 ( .A1(n6177), .A2(n4298), .ZN(n5888) );
  NAND2_X1 U5291 ( .A1(n5880), .A2(n5696), .ZN(n5668) );
  INV_X1 U5292 ( .A(n5676), .ZN(n5670) );
  NAND2_X1 U5293 ( .A1(n5670), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4302) );
  NOR2_X1 U5294 ( .A1(n5668), .A2(n4302), .ZN(n5661) );
  NAND3_X1 U5295 ( .A1(n5661), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n4379), .ZN(n4303) );
  AND2_X1 U5296 ( .A1(n4304), .A2(n4303), .ZN(n4305) );
  OAI21_X1 U5297 ( .B1(n4306), .B2(n5779), .A(n4305), .ZN(U2987) );
  INV_X1 U5298 ( .A(n4307), .ZN(n4311) );
  INV_X1 U5299 ( .A(n4308), .ZN(n4310) );
  AOI21_X1 U5300 ( .B1(n4311), .B2(n4310), .A(n4309), .ZN(n5858) );
  INV_X1 U5301 ( .A(n5858), .ZN(n5497) );
  INV_X1 U5302 ( .A(n5401), .ZN(n4312) );
  INV_X1 U5303 ( .A(n5404), .ZN(n4313) );
  NAND2_X1 U5304 ( .A1(n5405), .A2(n4313), .ZN(n4344) );
  NOR2_X1 U5305 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n4482) );
  INV_X1 U5306 ( .A(n4482), .ZN(n6583) );
  NOR3_X1 U5307 ( .A1(n6490), .A2(n6573), .A3(n6583), .ZN(n6486) );
  INV_X1 U5308 ( .A(n6486), .ZN(n4316) );
  NOR3_X1 U5309 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n4314), .A3(n6493), .ZN(
        n6495) );
  INV_X1 U5310 ( .A(n6495), .ZN(n4315) );
  NAND2_X1 U5311 ( .A1(n4316), .A2(n4315), .ZN(n4317) );
  NOR2_X1 U5312 ( .A1(n6215), .A2(n4317), .ZN(n4318) );
  NOR2_X1 U5313 ( .A1(n5497), .A2(n5971), .ZN(n4343) );
  INV_X1 U5314 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6687) );
  INV_X1 U5315 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6756) );
  NAND2_X1 U5316 ( .A1(n6728), .A2(n6656), .ZN(n4336) );
  INV_X1 U5317 ( .A(n4336), .ZN(n4320) );
  AND3_X1 U5318 ( .A1(n4321), .A2(n4145), .A3(n4320), .ZN(n4322) );
  INV_X1 U5319 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6538) );
  INV_X1 U5320 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6528) );
  INV_X1 U5321 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6525) );
  NAND3_X1 U5322 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6003) );
  NOR2_X1 U5323 ( .A1(n6525), .A2(n6003), .ZN(n5987) );
  NAND2_X1 U5324 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5987), .ZN(n5964) );
  NOR2_X1 U5325 ( .A1(n6528), .A2(n5964), .ZN(n5951) );
  NAND3_X1 U5326 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        n5951), .ZN(n5019) );
  NAND2_X1 U5327 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n5020) );
  NOR2_X1 U5328 ( .A1(n5019), .A2(n5020), .ZN(n5082) );
  NAND2_X1 U5329 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5082), .ZN(n5935) );
  NOR2_X1 U5330 ( .A1(n6538), .A2(n5935), .ZN(n5937) );
  NAND2_X1 U5331 ( .A1(REIP_REG_13__SCAN_IN), .A2(n5937), .ZN(n4325) );
  NAND3_X1 U5332 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n4326) );
  NAND3_X1 U5333 ( .A1(n5821), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n5460) );
  NAND4_X1 U5334 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5442), .ZN(n5317) );
  OR2_X1 U5335 ( .A1(n6687), .A2(n5317), .ZN(n5801) );
  NOR2_X1 U5336 ( .A1(n5801), .A2(REIP_REG_25__SCAN_IN), .ZN(n4342) );
  NAND2_X1 U5337 ( .A1(n4323), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4324) );
  NAND2_X1 U5338 ( .A1(n5978), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4330)
         );
  NAND3_X1 U5339 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4327) );
  INV_X1 U5340 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6540) );
  OR3_X1 U5341 ( .A1(n6540), .A2(n4325), .A3(n5963), .ZN(n5187) );
  NOR2_X1 U5342 ( .A1(n4326), .A2(n5187), .ZN(n5283) );
  NAND4_X1 U5343 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .A4(n5283), .ZN(n5443) );
  NOR2_X1 U5344 ( .A1(n4327), .A2(n5443), .ZN(n4328) );
  INV_X1 U5345 ( .A(n5963), .ZN(n5999) );
  NAND2_X1 U5346 ( .A1(n5965), .A2(n5999), .ZN(n5962) );
  INV_X1 U5347 ( .A(n5962), .ZN(n5282) );
  OR2_X1 U5348 ( .A1(n4328), .A2(n5282), .ZN(n5323) );
  INV_X1 U5349 ( .A(n5323), .ZN(n5436) );
  NOR2_X1 U5350 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5317), .ZN(n5423) );
  OAI21_X1 U5351 ( .B1(n5436), .B2(n5423), .A(REIP_REG_25__SCAN_IN), .ZN(n4329) );
  OAI211_X1 U5352 ( .C1(n6022), .C2(n5861), .A(n4330), .B(n4329), .ZN(n4341)
         );
  OR2_X1 U5353 ( .A1(n5418), .A2(n4331), .ZN(n4332) );
  NAND2_X1 U5354 ( .A1(n5492), .A2(n4332), .ZN(n5874) );
  NAND2_X1 U5355 ( .A1(n4336), .A2(EBX_REG_31__SCAN_IN), .ZN(n4333) );
  NOR2_X1 U5356 ( .A1(n5396), .A2(n4333), .ZN(n4334) );
  NAND3_X1 U5357 ( .A1(n6728), .A2(n6656), .A3(n5410), .ZN(n6479) );
  AND2_X1 U5358 ( .A1(n4335), .A2(n6479), .ZN(n5346) );
  INV_X1 U5359 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5357) );
  AND3_X1 U5360 ( .A1(n4145), .A2(n5357), .A3(n4336), .ZN(n4337) );
  NOR2_X1 U5361 ( .A1(n5346), .A2(n4337), .ZN(n4338) );
  NOR2_X4 U5362 ( .A1(n5089), .A2(n4338), .ZN(n6018) );
  NAND2_X1 U5363 ( .A1(n6018), .A2(EBX_REG_25__SCAN_IN), .ZN(n4339) );
  OAI21_X1 U5364 ( .B1(n5874), .B2(n6009), .A(n4339), .ZN(n4340) );
  OR4_X1 U5365 ( .A1(n4343), .A2(n4342), .A3(n4341), .A4(n4340), .ZN(U2802) );
  AOI22_X1 U5366 ( .A1(n5407), .A2(n3545), .B1(n5401), .B2(n4344), .ZN(n5412)
         );
  AND2_X1 U5367 ( .A1(n5412), .A2(n6491), .ZN(n4346) );
  INV_X1 U5368 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6713) );
  NAND3_X1 U5369 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4482), .A3(n6573), .ZN(
        n4345) );
  OAI21_X1 U5370 ( .B1(n4346), .B2(n6713), .A(n4345), .ZN(U2790) );
  INV_X1 U5371 ( .A(n4347), .ZN(n4349) );
  INV_X1 U5372 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n4348) );
  OR2_X1 U5373 ( .A1(n6586), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5397) );
  OAI211_X1 U5374 ( .C1(n4349), .C2(n4348), .A(n6072), .B(n5397), .ZN(U2788)
         );
  OAI21_X1 U5375 ( .B1(n4402), .B2(n6070), .A(n5410), .ZN(n4350) );
  NAND2_X1 U5376 ( .A1(n6049), .A2(n4145), .ZN(n4437) );
  NOR2_X1 U5377 ( .A1(n6493), .A2(n6481), .ZN(n4484) );
  INV_X1 U5378 ( .A(n6067), .ZN(n6588) );
  AOI22_X1 U5379 ( .A1(n4431), .A2(UWORD_REG_8__SCAN_IN), .B1(n6066), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4352) );
  OAI21_X1 U5380 ( .B1(n3972), .B2(n4437), .A(n4352), .ZN(U2899) );
  INV_X1 U5381 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6097) );
  AOI22_X1 U5382 ( .A1(n4431), .A2(UWORD_REG_10__SCAN_IN), .B1(n6066), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4353) );
  OAI21_X1 U5383 ( .B1(n6097), .B2(n4437), .A(n4353), .ZN(U2897) );
  INV_X1 U5384 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6099) );
  AOI22_X1 U5385 ( .A1(n4431), .A2(UWORD_REG_11__SCAN_IN), .B1(n6066), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4354) );
  OAI21_X1 U5386 ( .B1(n6099), .B2(n4437), .A(n4354), .ZN(U2896) );
  INV_X1 U5387 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6101) );
  AOI22_X1 U5388 ( .A1(n4431), .A2(UWORD_REG_12__SCAN_IN), .B1(n6066), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4355) );
  OAI21_X1 U5389 ( .B1(n6101), .B2(n4437), .A(n4355), .ZN(U2895) );
  INV_X1 U5390 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6103) );
  AOI22_X1 U5391 ( .A1(n4431), .A2(UWORD_REG_13__SCAN_IN), .B1(n6066), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4356) );
  OAI21_X1 U5392 ( .B1(n6103), .B2(n4437), .A(n4356), .ZN(U2894) );
  INV_X1 U5393 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6095) );
  AOI22_X1 U5394 ( .A1(n4431), .A2(UWORD_REG_9__SCAN_IN), .B1(n6066), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4357) );
  OAI21_X1 U5395 ( .B1(n6095), .B2(n4437), .A(n4357), .ZN(U2898) );
  INV_X1 U5396 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6107) );
  AOI22_X1 U5397 ( .A1(n4431), .A2(UWORD_REG_14__SCAN_IN), .B1(n6066), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4358) );
  OAI21_X1 U5398 ( .B1(n6107), .B2(n4437), .A(n4358), .ZN(U2893) );
  NAND2_X1 U5399 ( .A1(n6490), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6571) );
  INV_X1 U5400 ( .A(n6571), .ZN(n4524) );
  INV_X1 U5401 ( .A(n4359), .ZN(n4360) );
  OAI22_X1 U5402 ( .A1(n5407), .A2(n5402), .B1(n4144), .B2(n4360), .ZN(n4422)
         );
  INV_X1 U5403 ( .A(n4422), .ZN(n4368) );
  INV_X1 U5404 ( .A(n5407), .ZN(n5399) );
  OAI21_X1 U5405 ( .B1(n4402), .B2(n3241), .A(n5410), .ZN(n4361) );
  AOI21_X1 U5406 ( .B1(n4361), .B2(n4423), .A(READY_N), .ZN(n4366) );
  INV_X1 U5407 ( .A(n4362), .ZN(n4363) );
  NAND2_X1 U5408 ( .A1(n4364), .A2(n4363), .ZN(n4365) );
  AOI21_X1 U5409 ( .B1(n5399), .B2(n4366), .A(n4365), .ZN(n4367) );
  NAND2_X1 U5410 ( .A1(n5400), .A2(n5407), .ZN(n4568) );
  NAND2_X1 U5411 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4484), .ZN(n6570) );
  INV_X1 U5412 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6674) );
  OAI22_X1 U5413 ( .A1(n6459), .A2(n4369), .B1(n6570), .B2(n6674), .ZN(n5908)
         );
  NOR2_X1 U5414 ( .A1(n4524), .A2(n5908), .ZN(n5332) );
  INV_X1 U5415 ( .A(n4370), .ZN(n5782) );
  NAND4_X1 U5416 ( .A1(n4144), .A2(n4124), .A3(n4420), .A4(n4371), .ZN(n4372)
         );
  NOR2_X1 U5417 ( .A1(n4373), .A2(n4372), .ZN(n5333) );
  NOR3_X1 U5418 ( .A1(n4376), .A2(n4374), .A3(n4375), .ZN(n4377) );
  AOI21_X1 U5419 ( .B1(n4402), .B2(n3251), .A(n4377), .ZN(n4378) );
  OAI21_X1 U5420 ( .B1(n5782), .B2(n5333), .A(n4378), .ZN(n6457) );
  AOI22_X1 U5421 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4379), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4153), .ZN(n4400) );
  INV_X1 U5422 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6232) );
  NOR2_X1 U5423 ( .A1(n6493), .A2(n6232), .ZN(n4411) );
  INV_X1 U5424 ( .A(n4375), .ZN(n4477) );
  NOR2_X1 U5425 ( .A1(n4374), .A2(n6483), .ZN(n4413) );
  AOI222_X1 U5426 ( .A1(n6457), .A2(n5340), .B1(n4400), .B2(n4411), .C1(n4477), 
        .C2(n4413), .ZN(n4381) );
  NAND2_X1 U5427 ( .A1(n5332), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4380) );
  OAI21_X1 U5428 ( .B1(n5332), .B2(n4381), .A(n4380), .ZN(U3460) );
  INV_X1 U5429 ( .A(n6277), .ZN(n4917) );
  NAND2_X1 U5430 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4383) );
  INV_X1 U5431 ( .A(n4383), .ZN(n4384) );
  MUX2_X1 U5432 ( .A(n4384), .B(n4383), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4390) );
  INV_X1 U5433 ( .A(n4403), .ZN(n4389) );
  INV_X1 U5434 ( .A(n4374), .ZN(n4386) );
  OAI21_X1 U5435 ( .B1(n4386), .B2(n4385), .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .ZN(n4387) );
  NAND2_X1 U5436 ( .A1(n4388), .A2(n4387), .ZN(n4397) );
  AOI22_X1 U5437 ( .A1(n4402), .A2(n4390), .B1(n4389), .B2(n4397), .ZN(n4396)
         );
  MUX2_X1 U5438 ( .A(n4392), .B(n3359), .S(n4374), .Z(n4394) );
  INV_X1 U5439 ( .A(n5400), .ZN(n4393) );
  NAND2_X1 U5440 ( .A1(n4393), .A2(n5402), .ZN(n4407) );
  OAI21_X1 U5441 ( .B1(n4391), .B2(n4394), .A(n4407), .ZN(n4395) );
  OAI211_X1 U5442 ( .C1(n4917), .C2(n5333), .A(n4396), .B(n4395), .ZN(n4472)
         );
  AOI22_X1 U5443 ( .A1(n4472), .A2(n5340), .B1(n5336), .B2(n4397), .ZN(n4399)
         );
  NAND2_X1 U5444 ( .A1(n5332), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4398) );
  OAI21_X1 U5445 ( .B1(n5332), .B2(n4399), .A(n4398), .ZN(U3456) );
  INV_X1 U5446 ( .A(n4400), .ZN(n4412) );
  NOR2_X1 U5447 ( .A1(n6483), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4410)
         );
  INV_X1 U5448 ( .A(n3021), .ZN(n4409) );
  XNOR2_X1 U5449 ( .A(n4374), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4406)
         );
  INV_X1 U5450 ( .A(n4402), .ZN(n5339) );
  XNOR2_X1 U5451 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4404) );
  OAI22_X1 U5452 ( .A1(n5339), .A2(n4404), .B1(n4403), .B2(n4406), .ZN(n4405)
         );
  AOI21_X1 U5453 ( .B1(n4407), .B2(n4406), .A(n4405), .ZN(n4408) );
  OAI21_X1 U5454 ( .B1(n4409), .B2(n5333), .A(n4408), .ZN(n4473) );
  AOI222_X1 U5455 ( .A1(n4412), .A2(n4411), .B1(n4374), .B2(n4410), .C1(n4473), 
        .C2(n5340), .ZN(n4415) );
  OAI21_X1 U5456 ( .B1(n5332), .B2(n4413), .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .ZN(n4414) );
  OAI21_X1 U5457 ( .B1(n5332), .B2(n4415), .A(n4414), .ZN(U3459) );
  INV_X1 U5458 ( .A(n4416), .ZN(n4417) );
  OAI21_X1 U5459 ( .B1(n4419), .B2(n4418), .A(n4417), .ZN(n5096) );
  NAND3_X1 U5460 ( .A1(n5527), .A2(n4529), .A3(n3612), .ZN(n4564) );
  NOR2_X1 U5461 ( .A1(n4420), .A2(n4564), .ZN(n4421) );
  OAI21_X1 U5462 ( .B1(n4422), .B2(n4421), .A(n6491), .ZN(n4425) );
  NOR2_X1 U5463 ( .A1(n4423), .A2(READY_N), .ZN(n4424) );
  OR2_X1 U5464 ( .A1(n3218), .A2(n5527), .ZN(n4426) );
  INV_X1 U5465 ( .A(n4426), .ZN(n4427) );
  INV_X1 U5466 ( .A(DATAI_1_), .ZN(n6737) );
  INV_X1 U5467 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6113) );
  OAI222_X1 U5468 ( .A1(n5096), .A2(n5837), .B1(n5221), .B2(n6737), .C1(n5526), 
        .C2(n6113), .ZN(U2890) );
  INV_X1 U5469 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6086) );
  AOI22_X1 U5470 ( .A1(n4431), .A2(UWORD_REG_5__SCAN_IN), .B1(n6062), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4428) );
  OAI21_X1 U5471 ( .B1(n6086), .B2(n4437), .A(n4428), .ZN(U2902) );
  INV_X1 U5472 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6090) );
  AOI22_X1 U5473 ( .A1(n4431), .A2(UWORD_REG_6__SCAN_IN), .B1(n6062), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4429) );
  OAI21_X1 U5474 ( .B1(n6090), .B2(n4437), .A(n4429), .ZN(U2901) );
  INV_X1 U5475 ( .A(EAX_REG_20__SCAN_IN), .ZN(n6084) );
  AOI22_X1 U5476 ( .A1(n4431), .A2(UWORD_REG_4__SCAN_IN), .B1(n6062), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4430) );
  OAI21_X1 U5477 ( .B1(n6084), .B2(n4437), .A(n4430), .ZN(U2903) );
  INV_X1 U5478 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6092) );
  AOI22_X1 U5479 ( .A1(n4431), .A2(UWORD_REG_7__SCAN_IN), .B1(n6062), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4432) );
  OAI21_X1 U5480 ( .B1(n6092), .B2(n4437), .A(n4432), .ZN(U2900) );
  INV_X1 U5481 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6077) );
  AOI22_X1 U5482 ( .A1(n6067), .A2(UWORD_REG_1__SCAN_IN), .B1(n6062), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4433) );
  OAI21_X1 U5483 ( .B1(n6077), .B2(n4437), .A(n4433), .ZN(U2906) );
  INV_X1 U5484 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6079) );
  AOI22_X1 U5485 ( .A1(n6067), .A2(UWORD_REG_2__SCAN_IN), .B1(n6062), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4434) );
  OAI21_X1 U5486 ( .B1(n6079), .B2(n4437), .A(n4434), .ZN(U2905) );
  INV_X1 U5487 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6081) );
  AOI22_X1 U5488 ( .A1(n6067), .A2(UWORD_REG_3__SCAN_IN), .B1(n6062), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4435) );
  OAI21_X1 U5489 ( .B1(n6081), .B2(n4437), .A(n4435), .ZN(U2904) );
  INV_X1 U5490 ( .A(EAX_REG_16__SCAN_IN), .ZN(n6075) );
  AOI22_X1 U5491 ( .A1(n6067), .A2(UWORD_REG_0__SCAN_IN), .B1(n6062), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4436) );
  OAI21_X1 U5492 ( .B1(n6075), .B2(n4437), .A(n4436), .ZN(U2907) );
  XNOR2_X1 U5493 ( .A(n4438), .B(n4439), .ZN(n4945) );
  NAND2_X1 U5494 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4440) );
  AOI21_X1 U5495 ( .B1(n4440), .B2(n5735), .A(n5733), .ZN(n6212) );
  OAI21_X1 U5496 ( .B1(n5739), .B2(n6206), .A(n6212), .ZN(n4497) );
  OAI21_X1 U5497 ( .B1(n4743), .B2(n4440), .A(n5739), .ZN(n4970) );
  AND2_X1 U5498 ( .A1(n6206), .A2(n4970), .ZN(n4442) );
  INV_X1 U5499 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4441) );
  AOI22_X1 U5500 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4497), .B1(n4442), 
        .B2(n4441), .ZN(n4444) );
  AND2_X1 U5501 ( .A1(n6215), .A2(REIP_REG_3__SCAN_IN), .ZN(n4941) );
  AOI21_X1 U5502 ( .B1(n6210), .B2(n6019), .A(n4941), .ZN(n4443) );
  OAI211_X1 U5503 ( .C1(n4945), .C2(n5779), .A(n4444), .B(n4443), .ZN(U3015)
         );
  OAI21_X1 U5504 ( .B1(n4447), .B2(n3007), .A(n3012), .ZN(n4983) );
  NAND2_X1 U5505 ( .A1(n6232), .A2(n5303), .ZN(n6223) );
  AOI21_X1 U5506 ( .B1(n6230), .B2(n6223), .A(n4153), .ZN(n4452) );
  AND2_X1 U5507 ( .A1(n6215), .A2(REIP_REG_1__SCAN_IN), .ZN(n4979) );
  XNOR2_X1 U5508 ( .A(n4448), .B(n4565), .ZN(n5086) );
  NOR2_X1 U5509 ( .A1(n6225), .A2(n5086), .ZN(n4451) );
  NOR3_X1 U5510 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4449), .A3(n5740), 
        .ZN(n4450) );
  NOR4_X1 U5511 ( .A1(n4452), .A2(n4979), .A3(n4451), .A4(n4450), .ZN(n4453)
         );
  OAI21_X1 U5512 ( .B1(n5779), .B2(n4983), .A(n4453), .ZN(U3017) );
  INV_X1 U5513 ( .A(n4455), .ZN(n4468) );
  OAI21_X1 U5514 ( .B1(n4456), .B2(n4454), .A(n4468), .ZN(n5154) );
  INV_X1 U5515 ( .A(DATAI_2_), .ZN(n6721) );
  INV_X1 U5516 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6116) );
  OAI222_X1 U5517 ( .A1(n5154), .A2(n5837), .B1(n5221), .B2(n6721), .C1(n5526), 
        .C2(n6116), .ZN(U2889) );
  OR2_X1 U5518 ( .A1(n4458), .A2(n4457), .ZN(n4459) );
  NAND2_X1 U5519 ( .A1(n4460), .A2(n4459), .ZN(n6176) );
  INV_X1 U5520 ( .A(DATAI_0_), .ZN(n6628) );
  INV_X1 U5521 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6110) );
  OAI222_X1 U5522 ( .A1(n6176), .A2(n5837), .B1(n5221), .B2(n6628), .C1(n5526), 
        .C2(n6110), .ZN(U2891) );
  AND2_X1 U5523 ( .A1(n4461), .A2(n4462), .ZN(n4464) );
  OR2_X1 U5524 ( .A1(n4464), .A2(n4463), .ZN(n4731) );
  AOI22_X1 U5525 ( .A1(n5225), .A2(DATAI_4_), .B1(n6045), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n4465) );
  OAI21_X1 U5526 ( .B1(n4731), .B2(n5837), .A(n4465), .ZN(U2887) );
  INV_X1 U5527 ( .A(n4466), .ZN(n4467) );
  NAND2_X1 U5528 ( .A1(n4468), .A2(n4467), .ZN(n4469) );
  AND2_X1 U5529 ( .A1(n4461), .A2(n4469), .ZN(n6031) );
  INV_X1 U5530 ( .A(n6031), .ZN(n4470) );
  INV_X1 U5531 ( .A(DATAI_3_), .ZN(n6658) );
  INV_X1 U5532 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6119) );
  OAI222_X1 U5533 ( .A1(n4470), .A2(n5837), .B1(n5221), .B2(n6658), .C1(n5526), 
        .C2(n6119), .ZN(U2888) );
  NAND2_X1 U5534 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6674), .ZN(n4476) );
  INV_X1 U5535 ( .A(n4471), .ZN(n4475) );
  MUX2_X1 U5536 ( .A(n4472), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6459), 
        .Z(n6467) );
  MUX2_X1 U5537 ( .A(n4473), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(n6459), 
        .Z(n6463) );
  NAND3_X1 U5538 ( .A1(n6467), .A2(n6493), .A3(n6463), .ZN(n4474) );
  OAI21_X1 U5539 ( .B1(n4476), .B2(n4475), .A(n4474), .ZN(n6474) );
  NAND2_X1 U5540 ( .A1(n6474), .A2(n4477), .ZN(n4485) );
  MUX2_X1 U5541 ( .A(n6459), .B(n6674), .S(STATE2_REG_1__SCAN_IN), .Z(n4481)
         );
  INV_X1 U5542 ( .A(n6282), .ZN(n4834) );
  OR2_X1 U5543 ( .A1(n4478), .A2(n4834), .ZN(n4479) );
  XNOR2_X1 U5544 ( .A(n4479), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6006)
         );
  INV_X1 U5545 ( .A(n6006), .ZN(n4480) );
  NOR3_X1 U5546 ( .A1(n4480), .A2(STATE2_REG_1__SCAN_IN), .A3(n4144), .ZN(
        n5909) );
  AOI21_X1 U5547 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n4481), .A(n5909), 
        .ZN(n6476) );
  AND3_X1 U5548 ( .A1(n4485), .A2(n6674), .A3(n6476), .ZN(n4483) );
  OAI21_X1 U5549 ( .B1(n4483), .B2(n6570), .A(n4520), .ZN(n6233) );
  NAND3_X1 U5550 ( .A1(n4485), .A2(n6476), .A3(n4484), .ZN(n6489) );
  INV_X1 U5551 ( .A(n6489), .ZN(n4487) );
  NAND2_X1 U5552 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6573), .ZN(n4510) );
  INV_X1 U5553 ( .A(n4510), .ZN(n5783) );
  OAI22_X1 U5554 ( .A1(n5097), .A2(n6586), .B1(n3617), .B2(n5783), .ZN(n4486)
         );
  OAI21_X1 U5555 ( .B1(n4487), .B2(n4486), .A(n6233), .ZN(n4488) );
  OAI21_X1 U5556 ( .B1(n6233), .B2(n6454), .A(n4488), .ZN(U3465) );
  XNOR2_X1 U5557 ( .A(n4489), .B(n4491), .ZN(n5153) );
  OAI211_X1 U5558 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4970), .B(n6206), .ZN(n4493) );
  AND2_X1 U5559 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4492) );
  NOR2_X1 U5560 ( .A1(n4493), .A2(n4492), .ZN(n4500) );
  AND2_X1 U5561 ( .A1(n6215), .A2(REIP_REG_4__SCAN_IN), .ZN(n5149) );
  OR2_X1 U5562 ( .A1(n4495), .A2(n4494), .ZN(n4496) );
  NAND2_X1 U5563 ( .A1(n4496), .A2(n4576), .ZN(n6010) );
  NOR2_X1 U5564 ( .A1(n6225), .A2(n6010), .ZN(n4499) );
  AND2_X1 U5565 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n4497), .ZN(n4498)
         );
  NOR4_X1 U5566 ( .A1(n4500), .A2(n5149), .A3(n4499), .A4(n4498), .ZN(n4501)
         );
  OAI21_X1 U5567 ( .B1(n5779), .B2(n5153), .A(n4501), .ZN(U3014) );
  INV_X1 U5568 ( .A(n6233), .ZN(n4514) );
  INV_X1 U5569 ( .A(n4858), .ZN(n4505) );
  NOR2_X1 U5570 ( .A1(n3029), .A2(n6656), .ZN(n4612) );
  NAND2_X1 U5571 ( .A1(n4505), .A2(n4612), .ZN(n5034) );
  NAND2_X1 U5572 ( .A1(n6236), .A2(n4506), .ZN(n6272) );
  INV_X1 U5573 ( .A(n6272), .ZN(n4613) );
  NAND2_X1 U5574 ( .A1(n4613), .A2(n6368), .ZN(n6320) );
  NAND3_X1 U5575 ( .A1(n5034), .A2(n6320), .A3(n6367), .ZN(n6237) );
  INV_X1 U5576 ( .A(n6586), .ZN(n6328) );
  NOR2_X1 U5577 ( .A1(n6586), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6280) );
  AOI222_X1 U5578 ( .A1(n6237), .A2(n6328), .B1(n6277), .B2(n4510), .C1(n4647), 
        .C2(n6280), .ZN(n4509) );
  NAND2_X1 U5579 ( .A1(n4514), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4508) );
  OAI21_X1 U5580 ( .B1(n4514), .B2(n4509), .A(n4508), .ZN(U3462) );
  INV_X1 U5581 ( .A(n6368), .ZN(n6235) );
  XNOR2_X1 U5582 ( .A(n6235), .B(n6236), .ZN(n4511) );
  AOI22_X1 U5583 ( .A1(n4511), .A2(n6328), .B1(n4510), .B2(n3021), .ZN(n4513)
         );
  NAND2_X1 U5584 ( .A1(n4514), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4512) );
  OAI21_X1 U5585 ( .B1(n4514), .B2(n4513), .A(n4512), .ZN(U3463) );
  NOR2_X1 U5586 ( .A1(n6175), .A2(n6668), .ZN(n6389) );
  INV_X1 U5587 ( .A(n6389), .ZN(n6294) );
  INV_X1 U5588 ( .A(n4612), .ZN(n4515) );
  OAI21_X1 U5589 ( .B1(n6367), .B2(n4515), .A(n6328), .ZN(n4521) );
  OR2_X1 U5590 ( .A1(n3021), .A2(n4370), .ZN(n4916) );
  INV_X1 U5591 ( .A(n3617), .ZN(n6370) );
  NAND2_X1 U5592 ( .A1(n6277), .A2(n6370), .ZN(n5030) );
  OR2_X1 U5593 ( .A1(n4916), .A2(n5030), .ZN(n4517) );
  NAND3_X1 U5594 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4695), .A3(n5106), .ZN(n4918) );
  NOR2_X1 U5595 ( .A1(n6454), .A2(n4918), .ZN(n4556) );
  INV_X1 U5596 ( .A(n4556), .ZN(n4516) );
  AND2_X1 U5597 ( .A1(n4517), .A2(n4516), .ZN(n4522) );
  INV_X1 U5598 ( .A(n4522), .ZN(n4519) );
  INV_X1 U5599 ( .A(n6326), .ZN(n6379) );
  AOI21_X1 U5600 ( .B1(n6586), .B2(n4918), .A(n6379), .ZN(n4518) );
  OAI21_X1 U5601 ( .B1(n4521), .B2(n4519), .A(n4518), .ZN(n4553) );
  NAND2_X1 U5602 ( .A1(DATAI_1_), .A2(n4837), .ZN(n6393) );
  INV_X1 U5603 ( .A(n6393), .ZN(n6291) );
  OAI22_X1 U5604 ( .A1(n4522), .A2(n4521), .B1(n6481), .B2(n4918), .ZN(n4552)
         );
  AOI22_X1 U5605 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4553), .B1(n6291), 
        .B2(n4552), .ZN(n4527) );
  NOR2_X2 U5606 ( .A1(n6367), .A2(n4833), .ZN(n6362) );
  INV_X1 U5607 ( .A(DATAI_25_), .ZN(n6693) );
  NOR2_X2 U5608 ( .A1(n6175), .A2(n6693), .ZN(n6390) );
  NOR2_X1 U5609 ( .A1(n4555), .A2(n4525), .ZN(n6388) );
  AOI22_X1 U5610 ( .A1(n6362), .A2(n6390), .B1(n6388), .B2(n4556), .ZN(n4526)
         );
  OAI211_X1 U5611 ( .C1(n6294), .C2(n5140), .A(n4527), .B(n4526), .ZN(U3093)
         );
  INV_X1 U5612 ( .A(DATAI_20_), .ZN(n4528) );
  NOR2_X1 U5613 ( .A1(n6175), .A2(n4528), .ZN(n6438) );
  INV_X1 U5614 ( .A(n6438), .ZN(n6304) );
  NAND2_X1 U5615 ( .A1(DATAI_4_), .A2(n4837), .ZN(n6407) );
  AOI22_X1 U5616 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4553), .B1(n6437), 
        .B2(n4552), .ZN(n4531) );
  NAND2_X1 U5617 ( .A1(n6162), .A2(DATAI_28_), .ZN(n6441) );
  INV_X1 U5618 ( .A(n6441), .ZN(n6404) );
  NOR2_X1 U5619 ( .A1(n4555), .A2(n4529), .ZN(n6436) );
  AOI22_X1 U5620 ( .A1(n6362), .A2(n6404), .B1(n6436), .B2(n4556), .ZN(n4530)
         );
  OAI211_X1 U5621 ( .C1(n6304), .C2(n5140), .A(n4531), .B(n4530), .ZN(U3096)
         );
  INV_X1 U5622 ( .A(DATAI_19_), .ZN(n4532) );
  NOR2_X1 U5623 ( .A1(n6175), .A2(n4532), .ZN(n6400) );
  INV_X1 U5624 ( .A(n6400), .ZN(n6301) );
  NAND2_X1 U5625 ( .A1(DATAI_3_), .A2(n4837), .ZN(n6403) );
  INV_X1 U5626 ( .A(n6403), .ZN(n6298) );
  AOI22_X1 U5627 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4553), .B1(n6298), 
        .B2(n4552), .ZN(n4535) );
  INV_X1 U5628 ( .A(DATAI_27_), .ZN(n6730) );
  NOR2_X2 U5629 ( .A1(n6175), .A2(n6730), .ZN(n6399) );
  NOR2_X1 U5630 ( .A1(n4555), .A2(n4533), .ZN(n6398) );
  AOI22_X1 U5631 ( .A1(n6362), .A2(n6399), .B1(n6398), .B2(n4556), .ZN(n4534)
         );
  OAI211_X1 U5632 ( .C1(n6301), .C2(n5140), .A(n4535), .B(n4534), .ZN(U3095)
         );
  INV_X1 U5633 ( .A(DATAI_18_), .ZN(n4536) );
  NOR2_X1 U5634 ( .A1(n6175), .A2(n4536), .ZN(n6432) );
  INV_X1 U5635 ( .A(n6432), .ZN(n6297) );
  NAND2_X1 U5636 ( .A1(DATAI_2_), .A2(n4837), .ZN(n6397) );
  AOI22_X1 U5637 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4553), .B1(n6431), 
        .B2(n4552), .ZN(n4539) );
  NAND2_X1 U5638 ( .A1(n6162), .A2(DATAI_26_), .ZN(n6435) );
  INV_X1 U5639 ( .A(n6435), .ZN(n6394) );
  NOR2_X1 U5640 ( .A1(n4555), .A2(n4537), .ZN(n6430) );
  AOI22_X1 U5641 ( .A1(n6362), .A2(n6394), .B1(n6430), .B2(n4556), .ZN(n4538)
         );
  OAI211_X1 U5642 ( .C1(n6297), .C2(n5140), .A(n4539), .B(n4538), .ZN(U3094)
         );
  INV_X1 U5643 ( .A(DATAI_23_), .ZN(n4540) );
  NOR2_X1 U5644 ( .A1(n6175), .A2(n4540), .ZN(n6447) );
  INV_X1 U5645 ( .A(n6447), .ZN(n6319) );
  NAND2_X1 U5646 ( .A1(DATAI_7_), .A2(n4837), .ZN(n6427) );
  AOI22_X1 U5647 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4553), .B1(n6445), 
        .B2(n4552), .ZN(n4543) );
  INV_X1 U5648 ( .A(DATAI_31_), .ZN(n4541) );
  NOR2_X1 U5649 ( .A1(n6175), .A2(n4541), .ZN(n6423) );
  AOI22_X1 U5650 ( .A1(n6362), .A2(n6423), .B1(n6443), .B2(n4556), .ZN(n4542)
         );
  OAI211_X1 U5651 ( .C1(n6319), .C2(n5140), .A(n4543), .B(n4542), .ZN(U3099)
         );
  INV_X1 U5652 ( .A(DATAI_21_), .ZN(n4544) );
  NOR2_X1 U5653 ( .A1(n6175), .A2(n4544), .ZN(n6409) );
  INV_X1 U5654 ( .A(n6409), .ZN(n6308) );
  NAND2_X1 U5655 ( .A1(DATAI_5_), .A2(n4837), .ZN(n6413) );
  INV_X1 U5656 ( .A(n6413), .ZN(n6305) );
  AOI22_X1 U5657 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4553), .B1(n6305), 
        .B2(n4552), .ZN(n4546) );
  INV_X1 U5658 ( .A(DATAI_29_), .ZN(n6736) );
  NOR2_X2 U5659 ( .A1(n6175), .A2(n6736), .ZN(n6410) );
  NOR2_X1 U5660 ( .A1(n4555), .A2(n3160), .ZN(n6408) );
  AOI22_X1 U5661 ( .A1(n6362), .A2(n6410), .B1(n6408), .B2(n4556), .ZN(n4545)
         );
  OAI211_X1 U5662 ( .C1(n6308), .C2(n5140), .A(n4546), .B(n4545), .ZN(U3097)
         );
  INV_X1 U5663 ( .A(DATAI_16_), .ZN(n4547) );
  NOR2_X1 U5664 ( .A1(n6175), .A2(n4547), .ZN(n6376) );
  INV_X1 U5665 ( .A(n6376), .ZN(n6290) );
  NAND2_X1 U5666 ( .A1(DATAI_0_), .A2(n4837), .ZN(n6387) );
  INV_X1 U5667 ( .A(n6387), .ZN(n6279) );
  AOI22_X1 U5668 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4553), .B1(n6279), 
        .B2(n4552), .ZN(n4550) );
  INV_X1 U5669 ( .A(DATAI_24_), .ZN(n6695) );
  NOR2_X2 U5670 ( .A1(n6175), .A2(n6695), .ZN(n6384) );
  NOR2_X1 U5671 ( .A1(n4555), .A2(n4548), .ZN(n6375) );
  AOI22_X1 U5672 ( .A1(n6362), .A2(n6384), .B1(n6375), .B2(n4556), .ZN(n4549)
         );
  OAI211_X1 U5673 ( .C1(n6290), .C2(n5140), .A(n4550), .B(n4549), .ZN(U3092)
         );
  INV_X1 U5674 ( .A(DATAI_22_), .ZN(n4551) );
  NOR2_X1 U5675 ( .A1(n6175), .A2(n4551), .ZN(n6416) );
  INV_X1 U5676 ( .A(n6416), .ZN(n6311) );
  NAND2_X1 U5677 ( .A1(DATAI_6_), .A2(n4837), .ZN(n6419) );
  INV_X1 U5678 ( .A(n6419), .ZN(n6356) );
  AOI22_X1 U5679 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4553), .B1(n6356), 
        .B2(n4552), .ZN(n4558) );
  INV_X1 U5680 ( .A(DATAI_30_), .ZN(n6703) );
  NOR2_X1 U5681 ( .A1(n6175), .A2(n6703), .ZN(n6415) );
  NOR2_X1 U5682 ( .A1(n4555), .A2(n4554), .ZN(n6414) );
  AOI22_X1 U5683 ( .A1(n6362), .A2(n6415), .B1(n6414), .B2(n4556), .ZN(n4557)
         );
  OAI211_X1 U5684 ( .C1(n6311), .C2(n5140), .A(n4558), .B(n4557), .ZN(U3098)
         );
  OAI21_X1 U5685 ( .B1(n4463), .B2(n4560), .A(n4559), .ZN(n5991) );
  INV_X1 U5686 ( .A(DATAI_5_), .ZN(n6787) );
  INV_X1 U5687 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6125) );
  OAI222_X1 U5688 ( .A1(n5991), .A2(n5837), .B1(n5221), .B2(n6787), .C1(n5526), 
        .C2(n6125), .ZN(U2886) );
  NOR2_X1 U5689 ( .A1(n4561), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4562)
         );
  OR2_X1 U5690 ( .A1(n4563), .A2(n4562), .ZN(n6224) );
  INV_X1 U5691 ( .A(n4564), .ZN(n4566) );
  NAND3_X1 U5692 ( .A1(n3038), .A2(n4566), .A3(n4565), .ZN(n4567) );
  NAND2_X1 U5693 ( .A1(n4568), .A2(n4567), .ZN(n4569) );
  INV_X2 U5694 ( .A(n5831), .ZN(n5522) );
  OAI222_X1 U5695 ( .A1(n6224), .A2(n5522), .B1(n5836), .B2(n5209), .C1(n6176), 
        .C2(n5524), .ZN(U2859) );
  OAI22_X1 U5696 ( .A1(n5522), .A2(n5086), .B1(n5836), .B2(n4570), .ZN(n4571)
         );
  INV_X1 U5697 ( .A(n4571), .ZN(n4572) );
  OAI21_X1 U5698 ( .B1(n5096), .B2(n5524), .A(n4572), .ZN(U2858) );
  XNOR2_X1 U5699 ( .A(n4574), .B(n4573), .ZN(n6205) );
  OAI222_X1 U5700 ( .A1(n5524), .A2(n5154), .B1(n4575), .B2(n5836), .C1(n5522), 
        .C2(n6205), .ZN(U2857) );
  INV_X1 U5701 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4578) );
  AOI21_X1 U5702 ( .B1(n4577), .B2(n4576), .A(n4724), .ZN(n4748) );
  INV_X1 U5703 ( .A(n4748), .ZN(n5989) );
  OAI222_X1 U5704 ( .A1(n5991), .A2(n5524), .B1(n5836), .B2(n4578), .C1(n5989), 
        .C2(n5522), .ZN(U2854) );
  INV_X1 U5705 ( .A(n6390), .ZN(n5124) );
  NAND2_X1 U5706 ( .A1(n3029), .A2(n3419), .ZN(n4914) );
  NOR2_X2 U5707 ( .A1(n4858), .A2(n4914), .ZN(n4829) );
  NAND2_X1 U5708 ( .A1(n3021), .A2(n2983), .ZN(n6283) );
  OR2_X1 U5709 ( .A1(n5030), .A2(n6283), .ZN(n4579) );
  NAND2_X1 U5710 ( .A1(n4579), .A2(n4606), .ZN(n4582) );
  AOI22_X1 U5711 ( .A1(n4582), .A2(n6328), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4862), .ZN(n4607) );
  INV_X1 U5712 ( .A(n6388), .ZN(n4923) );
  OAI22_X1 U5713 ( .A1(n6393), .A2(n4607), .B1(n4606), .B2(n4923), .ZN(n4580)
         );
  AOI21_X1 U5714 ( .B1(n6389), .B2(n4829), .A(n4580), .ZN(n4587) );
  AND2_X1 U5715 ( .A1(n4581), .A2(n6162), .ZN(n4584) );
  INV_X1 U5716 ( .A(n4582), .ZN(n4583) );
  OAI21_X1 U5717 ( .B1(n4584), .B2(n6280), .A(n4583), .ZN(n4585) );
  OAI211_X1 U5718 ( .C1(n4862), .C2(n6328), .A(n4585), .B(n6326), .ZN(n4609)
         );
  NAND2_X1 U5719 ( .A1(n4609), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4586)
         );
  OAI211_X1 U5720 ( .C1(n4899), .C2(n5124), .A(n4587), .B(n4586), .ZN(U3141)
         );
  INV_X1 U5721 ( .A(n6430), .ZN(n4868) );
  OAI22_X1 U5722 ( .A1(n6397), .A2(n4607), .B1(n4606), .B2(n4868), .ZN(n4588)
         );
  AOI21_X1 U5723 ( .B1(n6432), .B2(n4829), .A(n4588), .ZN(n4590) );
  NAND2_X1 U5724 ( .A1(n4609), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4589)
         );
  OAI211_X1 U5725 ( .C1(n4899), .C2(n6435), .A(n4590), .B(n4589), .ZN(U3142)
         );
  INV_X1 U5726 ( .A(n6384), .ZN(n5116) );
  INV_X1 U5727 ( .A(n6375), .ZN(n4936) );
  OAI22_X1 U5728 ( .A1(n6387), .A2(n4607), .B1(n4606), .B2(n4936), .ZN(n4591)
         );
  AOI21_X1 U5729 ( .B1(n6376), .B2(n4829), .A(n4591), .ZN(n4593) );
  NAND2_X1 U5730 ( .A1(n4609), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4592)
         );
  OAI211_X1 U5731 ( .C1(n4899), .C2(n5116), .A(n4593), .B(n4592), .ZN(U3140)
         );
  INV_X1 U5732 ( .A(n6423), .ZN(n6452) );
  INV_X1 U5733 ( .A(n6443), .ZN(n4888) );
  OAI22_X1 U5734 ( .A1(n6427), .A2(n4607), .B1(n4606), .B2(n4888), .ZN(n4594)
         );
  AOI21_X1 U5735 ( .B1(n6447), .B2(n4829), .A(n4594), .ZN(n4596) );
  NAND2_X1 U5736 ( .A1(n4609), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4595)
         );
  OAI211_X1 U5737 ( .C1(n4899), .C2(n6452), .A(n4596), .B(n4595), .ZN(U3147)
         );
  INV_X1 U5738 ( .A(n6399), .ZN(n5131) );
  INV_X1 U5739 ( .A(n6398), .ZN(n4927) );
  OAI22_X1 U5740 ( .A1(n6403), .A2(n4607), .B1(n4606), .B2(n4927), .ZN(n4597)
         );
  AOI21_X1 U5741 ( .B1(n6400), .B2(n4829), .A(n4597), .ZN(n4599) );
  NAND2_X1 U5742 ( .A1(n4609), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4598)
         );
  OAI211_X1 U5743 ( .C1(n4899), .C2(n5131), .A(n4599), .B(n4598), .ZN(U3143)
         );
  INV_X1 U5744 ( .A(n6436), .ZN(n4894) );
  OAI22_X1 U5745 ( .A1(n6407), .A2(n4607), .B1(n4606), .B2(n4894), .ZN(n4600)
         );
  AOI21_X1 U5746 ( .B1(n6438), .B2(n4829), .A(n4600), .ZN(n4602) );
  NAND2_X1 U5747 ( .A1(n4609), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4601)
         );
  OAI211_X1 U5748 ( .C1(n4899), .C2(n6441), .A(n4602), .B(n4601), .ZN(U3144)
         );
  INV_X1 U5749 ( .A(n6410), .ZN(n5120) );
  INV_X1 U5750 ( .A(n6408), .ZN(n4931) );
  OAI22_X1 U5751 ( .A1(n6413), .A2(n4607), .B1(n4606), .B2(n4931), .ZN(n4603)
         );
  AOI21_X1 U5752 ( .B1(n6409), .B2(n4829), .A(n4603), .ZN(n4605) );
  NAND2_X1 U5753 ( .A1(n4609), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4604)
         );
  OAI211_X1 U5754 ( .C1(n4899), .C2(n5120), .A(n4605), .B(n4604), .ZN(U3145)
         );
  INV_X1 U5755 ( .A(n6415), .ZN(n6359) );
  INV_X1 U5756 ( .A(n6414), .ZN(n4875) );
  OAI22_X1 U5757 ( .A1(n6419), .A2(n4607), .B1(n4606), .B2(n4875), .ZN(n4608)
         );
  AOI21_X1 U5758 ( .B1(n6416), .B2(n4829), .A(n4608), .ZN(n4611) );
  NAND2_X1 U5759 ( .A1(n4609), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4610)
         );
  OAI211_X1 U5760 ( .C1(n4899), .C2(n6359), .A(n4611), .B(n4610), .ZN(U3146)
         );
  AOI21_X1 U5761 ( .B1(n4613), .B2(n4612), .A(n6586), .ZN(n4762) );
  NAND2_X1 U5762 ( .A1(n3021), .A2(n5782), .ZN(n5031) );
  OR2_X1 U5763 ( .A1(n5031), .A2(n6282), .ZN(n4761) );
  NAND2_X1 U5764 ( .A1(n5106), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5038) );
  OR2_X1 U5765 ( .A1(n5038), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4763)
         );
  OR2_X1 U5766 ( .A1(n6454), .A2(n4763), .ZN(n4640) );
  OAI21_X1 U5767 ( .B1(n4761), .B2(n3617), .A(n4640), .ZN(n4616) );
  INV_X1 U5768 ( .A(n4763), .ZN(n4614) );
  AOI22_X1 U5769 ( .A1(n4762), .A2(n4616), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4614), .ZN(n4645) );
  INV_X1 U5770 ( .A(n4762), .ZN(n4617) );
  AOI21_X1 U5771 ( .B1(n6586), .B2(n4763), .A(n6379), .ZN(n4615) );
  NAND2_X1 U5772 ( .A1(n4639), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4620) );
  NOR2_X2 U5773 ( .A1(n6272), .A2(n4833), .ZN(n4792) );
  INV_X1 U5774 ( .A(n6314), .ZN(n4641) );
  OAI22_X1 U5775 ( .A1(n4641), .A2(n6304), .B1(n4894), .B2(n4640), .ZN(n4618)
         );
  AOI21_X1 U5776 ( .B1(n6404), .B2(n4792), .A(n4618), .ZN(n4619) );
  OAI211_X1 U5777 ( .C1(n4645), .C2(n6407), .A(n4620), .B(n4619), .ZN(U3064)
         );
  NAND2_X1 U5778 ( .A1(n4639), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4623) );
  OAI22_X1 U5779 ( .A1(n4641), .A2(n6311), .B1(n4875), .B2(n4640), .ZN(n4621)
         );
  AOI21_X1 U5780 ( .B1(n6415), .B2(n4792), .A(n4621), .ZN(n4622) );
  OAI211_X1 U5781 ( .C1(n4645), .C2(n6419), .A(n4623), .B(n4622), .ZN(U3066)
         );
  NAND2_X1 U5782 ( .A1(n4639), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4626) );
  OAI22_X1 U5783 ( .A1(n4641), .A2(n6319), .B1(n4888), .B2(n4640), .ZN(n4624)
         );
  AOI21_X1 U5784 ( .B1(n6423), .B2(n4792), .A(n4624), .ZN(n4625) );
  OAI211_X1 U5785 ( .C1(n4645), .C2(n6427), .A(n4626), .B(n4625), .ZN(U3067)
         );
  NAND2_X1 U5786 ( .A1(n4639), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4629) );
  OAI22_X1 U5787 ( .A1(n4641), .A2(n6301), .B1(n4927), .B2(n4640), .ZN(n4627)
         );
  AOI21_X1 U5788 ( .B1(n6399), .B2(n4792), .A(n4627), .ZN(n4628) );
  OAI211_X1 U5789 ( .C1(n4645), .C2(n6403), .A(n4629), .B(n4628), .ZN(U3063)
         );
  NAND2_X1 U5790 ( .A1(n4639), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4632) );
  OAI22_X1 U5791 ( .A1(n4641), .A2(n6290), .B1(n4936), .B2(n4640), .ZN(n4630)
         );
  AOI21_X1 U5792 ( .B1(n6384), .B2(n4792), .A(n4630), .ZN(n4631) );
  OAI211_X1 U5793 ( .C1(n4645), .C2(n6387), .A(n4632), .B(n4631), .ZN(U3060)
         );
  NAND2_X1 U5794 ( .A1(n4639), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4635) );
  OAI22_X1 U5795 ( .A1(n4641), .A2(n6294), .B1(n4923), .B2(n4640), .ZN(n4633)
         );
  AOI21_X1 U5796 ( .B1(n6390), .B2(n4792), .A(n4633), .ZN(n4634) );
  OAI211_X1 U5797 ( .C1(n4645), .C2(n6393), .A(n4635), .B(n4634), .ZN(U3061)
         );
  NAND2_X1 U5798 ( .A1(n4639), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4638) );
  OAI22_X1 U5799 ( .A1(n4641), .A2(n6308), .B1(n4931), .B2(n4640), .ZN(n4636)
         );
  AOI21_X1 U5800 ( .B1(n6410), .B2(n4792), .A(n4636), .ZN(n4637) );
  OAI211_X1 U5801 ( .C1(n4645), .C2(n6413), .A(n4638), .B(n4637), .ZN(U3065)
         );
  NAND2_X1 U5802 ( .A1(n4639), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4644) );
  OAI22_X1 U5803 ( .A1(n4641), .A2(n6297), .B1(n4868), .B2(n4640), .ZN(n4642)
         );
  AOI21_X1 U5804 ( .B1(n6394), .B2(n4792), .A(n4642), .ZN(n4643) );
  OAI211_X1 U5805 ( .C1(n4645), .C2(n6397), .A(n4644), .B(n4643), .ZN(U3062)
         );
  NOR3_X1 U5806 ( .A1(n4647), .A2(n6236), .A3(n4646), .ZN(n4760) );
  NAND2_X1 U5807 ( .A1(n4760), .A2(n5097), .ZN(n6243) );
  INV_X1 U5808 ( .A(n4647), .ZN(n4649) );
  NOR2_X1 U5809 ( .A1(n3029), .A2(n6236), .ZN(n4648) );
  NAND2_X1 U5810 ( .A1(n4649), .A2(n4648), .ZN(n4701) );
  INV_X1 U5811 ( .A(n4701), .ZN(n4650) );
  AOI21_X1 U5812 ( .B1(n6243), .B2(n4721), .A(n6280), .ZN(n4651) );
  NOR2_X1 U5813 ( .A1(n6277), .A2(n5100), .ZN(n6239) );
  OAI21_X1 U5814 ( .B1(n4651), .B2(n6239), .A(n6573), .ZN(n4655) );
  NOR3_X1 U5815 ( .A1(n5106), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6242) );
  INV_X1 U5816 ( .A(n6242), .ZN(n6246) );
  NOR2_X1 U5817 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6246), .ZN(n4687)
         );
  INV_X1 U5818 ( .A(n4687), .ZN(n4654) );
  INV_X1 U5819 ( .A(n4656), .ZN(n4652) );
  NOR2_X1 U5820 ( .A1(n4652), .A2(n6481), .ZN(n6275) );
  OAI21_X1 U5821 ( .B1(n6274), .B2(n6481), .A(n4837), .ZN(n4861) );
  NOR2_X1 U5822 ( .A1(n6275), .A2(n4861), .ZN(n5111) );
  INV_X1 U5823 ( .A(n5111), .ZN(n4653) );
  INV_X1 U5824 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4662) );
  INV_X1 U5825 ( .A(n6239), .ZN(n4658) );
  NOR2_X1 U5826 ( .A1(n4656), .A2(n6481), .ZN(n5102) );
  NAND3_X1 U5827 ( .A1(n5102), .A2(n6274), .A3(n6468), .ZN(n4657) );
  OAI21_X1 U5828 ( .B1(n4658), .B2(n6586), .A(n4657), .ZN(n4688) );
  AOI22_X1 U5829 ( .A1(n6291), .A2(n4688), .B1(n6388), .B2(n4687), .ZN(n4659)
         );
  OAI21_X1 U5830 ( .B1(n6243), .B2(n6294), .A(n4659), .ZN(n4660) );
  AOI21_X1 U5831 ( .B1(n4691), .B2(n6390), .A(n4660), .ZN(n4661) );
  OAI21_X1 U5832 ( .B1(n4694), .B2(n4662), .A(n4661), .ZN(U3037) );
  INV_X1 U5833 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4666) );
  AOI22_X1 U5834 ( .A1(n6305), .A2(n4688), .B1(n6408), .B2(n4687), .ZN(n4663)
         );
  OAI21_X1 U5835 ( .B1(n6243), .B2(n6308), .A(n4663), .ZN(n4664) );
  AOI21_X1 U5836 ( .B1(n4691), .B2(n6410), .A(n4664), .ZN(n4665) );
  OAI21_X1 U5837 ( .B1(n4694), .B2(n4666), .A(n4665), .ZN(U3041) );
  INV_X1 U5838 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4670) );
  AOI22_X1 U5839 ( .A1(n6298), .A2(n4688), .B1(n6398), .B2(n4687), .ZN(n4667)
         );
  OAI21_X1 U5840 ( .B1(n6243), .B2(n6301), .A(n4667), .ZN(n4668) );
  AOI21_X1 U5841 ( .B1(n4691), .B2(n6399), .A(n4668), .ZN(n4669) );
  OAI21_X1 U5842 ( .B1(n4694), .B2(n4670), .A(n4669), .ZN(U3039) );
  INV_X1 U5843 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4674) );
  AOI22_X1 U5844 ( .A1(n6431), .A2(n4688), .B1(n6430), .B2(n4687), .ZN(n4671)
         );
  OAI21_X1 U5845 ( .B1(n6243), .B2(n6297), .A(n4671), .ZN(n4672) );
  AOI21_X1 U5846 ( .B1(n4691), .B2(n6394), .A(n4672), .ZN(n4673) );
  OAI21_X1 U5847 ( .B1(n4694), .B2(n4674), .A(n4673), .ZN(U3038) );
  INV_X1 U5848 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4678) );
  AOI22_X1 U5849 ( .A1(n6445), .A2(n4688), .B1(n6443), .B2(n4687), .ZN(n4675)
         );
  OAI21_X1 U5850 ( .B1(n6243), .B2(n6319), .A(n4675), .ZN(n4676) );
  AOI21_X1 U5851 ( .B1(n4691), .B2(n6423), .A(n4676), .ZN(n4677) );
  OAI21_X1 U5852 ( .B1(n4694), .B2(n4678), .A(n4677), .ZN(U3043) );
  INV_X1 U5853 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4682) );
  AOI22_X1 U5854 ( .A1(n6279), .A2(n4688), .B1(n6375), .B2(n4687), .ZN(n4679)
         );
  OAI21_X1 U5855 ( .B1(n6243), .B2(n6290), .A(n4679), .ZN(n4680) );
  AOI21_X1 U5856 ( .B1(n4691), .B2(n6384), .A(n4680), .ZN(n4681) );
  OAI21_X1 U5857 ( .B1(n4694), .B2(n4682), .A(n4681), .ZN(U3036) );
  INV_X1 U5858 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4686) );
  AOI22_X1 U5859 ( .A1(n6356), .A2(n4688), .B1(n6414), .B2(n4687), .ZN(n4683)
         );
  OAI21_X1 U5860 ( .B1(n6243), .B2(n6311), .A(n4683), .ZN(n4684) );
  AOI21_X1 U5861 ( .B1(n4691), .B2(n6415), .A(n4684), .ZN(n4685) );
  OAI21_X1 U5862 ( .B1(n4694), .B2(n4686), .A(n4685), .ZN(U3042) );
  INV_X1 U5863 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4693) );
  AOI22_X1 U5864 ( .A1(n6437), .A2(n4688), .B1(n6436), .B2(n4687), .ZN(n4689)
         );
  OAI21_X1 U5865 ( .B1(n6243), .B2(n6304), .A(n4689), .ZN(n4690) );
  AOI21_X1 U5866 ( .B1(n4691), .B2(n6404), .A(n4690), .ZN(n4692) );
  OAI21_X1 U5867 ( .B1(n4694), .B2(n4693), .A(n4692), .ZN(U3040) );
  NOR2_X1 U5868 ( .A1(n6277), .A2(n4916), .ZN(n4803) );
  NAND3_X1 U5869 ( .A1(n6468), .A2(n4695), .A3(n5106), .ZN(n4799) );
  NOR2_X1 U5870 ( .A1(n6454), .A2(n4799), .ZN(n4718) );
  AOI21_X1 U5871 ( .B1(n4803), .B2(n6370), .A(n4718), .ZN(n4700) );
  OR2_X1 U5872 ( .A1(n4701), .A2(n6656), .ZN(n4696) );
  AOI22_X1 U5873 ( .A1(n4700), .A2(n4698), .B1(n6586), .B2(n4799), .ZN(n4697)
         );
  NAND2_X1 U5874 ( .A1(n6326), .A2(n4697), .ZN(n4717) );
  INV_X1 U5875 ( .A(n4698), .ZN(n4699) );
  OAI22_X1 U5876 ( .A1(n4700), .A2(n4699), .B1(n6481), .B2(n4799), .ZN(n4716)
         );
  AOI22_X1 U5877 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4717), .B1(n6437), 
        .B2(n4716), .ZN(n4703) );
  AOI22_X1 U5878 ( .A1(n4797), .A2(n6404), .B1(n4718), .B2(n6436), .ZN(n4702)
         );
  OAI211_X1 U5879 ( .C1(n4721), .C2(n6304), .A(n4703), .B(n4702), .ZN(U3032)
         );
  AOI22_X1 U5880 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4717), .B1(n6298), 
        .B2(n4716), .ZN(n4705) );
  AOI22_X1 U5881 ( .A1(n4797), .A2(n6399), .B1(n4718), .B2(n6398), .ZN(n4704)
         );
  OAI211_X1 U5882 ( .C1(n4721), .C2(n6301), .A(n4705), .B(n4704), .ZN(U3031)
         );
  AOI22_X1 U5883 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4717), .B1(n6431), 
        .B2(n4716), .ZN(n4707) );
  AOI22_X1 U5884 ( .A1(n4797), .A2(n6394), .B1(n4718), .B2(n6430), .ZN(n4706)
         );
  OAI211_X1 U5885 ( .C1(n4721), .C2(n6297), .A(n4707), .B(n4706), .ZN(U3030)
         );
  AOI22_X1 U5886 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4717), .B1(n6445), 
        .B2(n4716), .ZN(n4709) );
  AOI22_X1 U5887 ( .A1(n4797), .A2(n6423), .B1(n4718), .B2(n6443), .ZN(n4708)
         );
  OAI211_X1 U5888 ( .C1(n4721), .C2(n6319), .A(n4709), .B(n4708), .ZN(U3035)
         );
  AOI22_X1 U5889 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4717), .B1(n6279), 
        .B2(n4716), .ZN(n4711) );
  AOI22_X1 U5890 ( .A1(n4797), .A2(n6384), .B1(n6375), .B2(n4718), .ZN(n4710)
         );
  OAI211_X1 U5891 ( .C1(n4721), .C2(n6290), .A(n4711), .B(n4710), .ZN(U3028)
         );
  AOI22_X1 U5892 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4717), .B1(n6305), 
        .B2(n4716), .ZN(n4713) );
  AOI22_X1 U5893 ( .A1(n4797), .A2(n6410), .B1(n4718), .B2(n6408), .ZN(n4712)
         );
  OAI211_X1 U5894 ( .C1(n4721), .C2(n6308), .A(n4713), .B(n4712), .ZN(U3033)
         );
  AOI22_X1 U5895 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4717), .B1(n6291), 
        .B2(n4716), .ZN(n4715) );
  AOI22_X1 U5896 ( .A1(n4797), .A2(n6390), .B1(n4718), .B2(n6388), .ZN(n4714)
         );
  OAI211_X1 U5897 ( .C1(n4721), .C2(n6294), .A(n4715), .B(n4714), .ZN(U3029)
         );
  AOI22_X1 U5898 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4717), .B1(n6356), 
        .B2(n4716), .ZN(n4720) );
  AOI22_X1 U5899 ( .A1(n4797), .A2(n6415), .B1(n4718), .B2(n6414), .ZN(n4719)
         );
  OAI211_X1 U5900 ( .C1(n4721), .C2(n6311), .A(n4720), .B(n4719), .ZN(U3034)
         );
  XNOR2_X1 U5901 ( .A(n2985), .B(n4723), .ZN(n5147) );
  OAI21_X1 U5902 ( .B1(n4727), .B2(n5740), .A(n6212), .ZN(n4745) );
  OR2_X1 U5903 ( .A1(n4725), .A2(n4724), .ZN(n4726) );
  NAND2_X1 U5904 ( .A1(n4726), .A2(n4757), .ZN(n5980) );
  OAI22_X1 U5905 ( .A1(n6225), .A2(n5980), .B1(n6528), .B2(n5900), .ZN(n4729)
         );
  AND3_X1 U5906 ( .A1(n4727), .A2(n4176), .A3(n4970), .ZN(n4728) );
  AOI211_X1 U5907 ( .C1(INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n4745), .A(n4729), 
        .B(n4728), .ZN(n4730) );
  OAI21_X1 U5908 ( .B1(n5147), .B2(n5779), .A(n4730), .ZN(U3012) );
  INV_X1 U5909 ( .A(n4731), .ZN(n6012) );
  OAI22_X1 U5910 ( .A1(n5522), .A2(n6010), .B1(n5836), .B2(n4732), .ZN(n4733)
         );
  AOI21_X1 U5911 ( .B1(n6012), .B2(n5833), .A(n4733), .ZN(n4734) );
  INV_X1 U5912 ( .A(n4734), .ZN(U2855) );
  INV_X1 U5913 ( .A(n6019), .ZN(n4736) );
  OAI22_X1 U5914 ( .A1(n5522), .A2(n4736), .B1(n5836), .B2(n4735), .ZN(n4737)
         );
  AOI21_X1 U5915 ( .B1(n6031), .B2(n5833), .A(n4737), .ZN(n4738) );
  INV_X1 U5916 ( .A(n4738), .ZN(U2856) );
  CLKBUF_X1 U5917 ( .A(n4740), .Z(n4741) );
  XOR2_X1 U5918 ( .A(n4739), .B(n4741), .Z(n4986) );
  INV_X1 U5919 ( .A(n4986), .ZN(n4751) );
  OAI22_X1 U5920 ( .A1(n5739), .A2(n4744), .B1(n4743), .B2(n4742), .ZN(n4746)
         );
  OAI21_X1 U5921 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4746), .A(n4745), 
        .ZN(n4750) );
  INV_X1 U5922 ( .A(REIP_REG_5__SCAN_IN), .ZN(n4747) );
  NOR2_X1 U5923 ( .A1(n5900), .A2(n4747), .ZN(n4989) );
  AOI21_X1 U5924 ( .B1(n6210), .B2(n4748), .A(n4989), .ZN(n4749) );
  OAI211_X1 U5925 ( .C1(n4751), .C2(n5779), .A(n4750), .B(n4749), .ZN(U3013)
         );
  INV_X1 U5926 ( .A(n4752), .ZN(n4949) );
  OR2_X1 U5927 ( .A1(n4752), .A2(n4755), .ZN(n4993) );
  OAI21_X1 U5928 ( .B1(n4949), .B2(n4754), .A(n4993), .ZN(n5972) );
  AOI21_X1 U5929 ( .B1(n4758), .B2(n4757), .A(n4756), .ZN(n6197) );
  AOI22_X1 U5930 ( .A1(n5831), .A2(n6197), .B1(EBX_REG_7__SCAN_IN), .B2(n5499), 
        .ZN(n4759) );
  OAI21_X1 U5931 ( .B1(n5972), .B2(n5524), .A(n4759), .ZN(U2852) );
  OAI211_X1 U5932 ( .C1(n4795), .C2(n6280), .A(n4762), .B(n4761), .ZN(n4766)
         );
  OR2_X1 U5933 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4763), .ZN(n4789)
         );
  INV_X1 U5934 ( .A(n4836), .ZN(n4764) );
  OAI21_X1 U5935 ( .B1(n3082), .B2(n6481), .A(n4837), .ZN(n4800) );
  AOI211_X1 U5936 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4789), .A(n5102), .B(
        n4800), .ZN(n4765) );
  NAND2_X1 U5937 ( .A1(n4766), .A2(n4765), .ZN(n4788) );
  NAND2_X1 U5938 ( .A1(n4788), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4769) );
  NOR2_X1 U5939 ( .A1(n5031), .A2(n6586), .ZN(n4840) );
  AOI22_X1 U5940 ( .A1(n4840), .A2(n4917), .B1(n6275), .B2(n3082), .ZN(n4790)
         );
  OAI22_X1 U5941 ( .A1(n6397), .A2(n4790), .B1(n4868), .B2(n4789), .ZN(n4767)
         );
  AOI21_X1 U5942 ( .B1(n6432), .B2(n4792), .A(n4767), .ZN(n4768) );
  OAI211_X1 U5943 ( .C1(n4795), .C2(n6435), .A(n4769), .B(n4768), .ZN(U3054)
         );
  NAND2_X1 U5944 ( .A1(n4788), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4772) );
  OAI22_X1 U5945 ( .A1(n6407), .A2(n4790), .B1(n4894), .B2(n4789), .ZN(n4770)
         );
  AOI21_X1 U5946 ( .B1(n6438), .B2(n4792), .A(n4770), .ZN(n4771) );
  OAI211_X1 U5947 ( .C1(n4795), .C2(n6441), .A(n4772), .B(n4771), .ZN(U3056)
         );
  NAND2_X1 U5948 ( .A1(n4788), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4775) );
  OAI22_X1 U5949 ( .A1(n6413), .A2(n4790), .B1(n4931), .B2(n4789), .ZN(n4773)
         );
  AOI21_X1 U5950 ( .B1(n6409), .B2(n4792), .A(n4773), .ZN(n4774) );
  OAI211_X1 U5951 ( .C1(n4795), .C2(n5120), .A(n4775), .B(n4774), .ZN(U3057)
         );
  NAND2_X1 U5952 ( .A1(n4788), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4778) );
  OAI22_X1 U5953 ( .A1(n6387), .A2(n4790), .B1(n4936), .B2(n4789), .ZN(n4776)
         );
  AOI21_X1 U5954 ( .B1(n6376), .B2(n4792), .A(n4776), .ZN(n4777) );
  OAI211_X1 U5955 ( .C1(n4795), .C2(n5116), .A(n4778), .B(n4777), .ZN(U3052)
         );
  NAND2_X1 U5956 ( .A1(n4788), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4781) );
  OAI22_X1 U5957 ( .A1(n6419), .A2(n4790), .B1(n4875), .B2(n4789), .ZN(n4779)
         );
  AOI21_X1 U5958 ( .B1(n6416), .B2(n4792), .A(n4779), .ZN(n4780) );
  OAI211_X1 U5959 ( .C1(n4795), .C2(n6359), .A(n4781), .B(n4780), .ZN(U3058)
         );
  NAND2_X1 U5960 ( .A1(n4788), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4784) );
  OAI22_X1 U5961 ( .A1(n6403), .A2(n4790), .B1(n4927), .B2(n4789), .ZN(n4782)
         );
  AOI21_X1 U5962 ( .B1(n6400), .B2(n4792), .A(n4782), .ZN(n4783) );
  OAI211_X1 U5963 ( .C1(n4795), .C2(n5131), .A(n4784), .B(n4783), .ZN(U3055)
         );
  NAND2_X1 U5964 ( .A1(n4788), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4787) );
  OAI22_X1 U5965 ( .A1(n6427), .A2(n4790), .B1(n4888), .B2(n4789), .ZN(n4785)
         );
  AOI21_X1 U5966 ( .B1(n6447), .B2(n4792), .A(n4785), .ZN(n4786) );
  OAI211_X1 U5967 ( .C1(n4795), .C2(n6452), .A(n4787), .B(n4786), .ZN(U3059)
         );
  NAND2_X1 U5968 ( .A1(n4788), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4794) );
  OAI22_X1 U5969 ( .A1(n6393), .A2(n4790), .B1(n4923), .B2(n4789), .ZN(n4791)
         );
  AOI21_X1 U5970 ( .B1(n6389), .B2(n4792), .A(n4791), .ZN(n4793) );
  OAI211_X1 U5971 ( .C1(n4795), .C2(n5124), .A(n4794), .B(n4793), .ZN(U3053)
         );
  INV_X1 U5972 ( .A(DATAI_7_), .ZN(n4796) );
  INV_X1 U5973 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6130) );
  OAI222_X1 U5974 ( .A1(n5972), .A2(n5837), .B1(n5221), .B2(n4796), .C1(n5526), 
        .C2(n6130), .ZN(U2884) );
  NOR3_X1 U5975 ( .A1(n4797), .A2(n4829), .A3(n6586), .ZN(n4798) );
  NOR2_X1 U5976 ( .A1(n4798), .A2(n6280), .ZN(n4802) );
  OR2_X1 U5977 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4799), .ZN(n4826)
         );
  AOI211_X1 U5978 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4826), .A(n6275), .B(
        n4800), .ZN(n4801) );
  NAND2_X1 U5979 ( .A1(n4825), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4806) );
  AOI22_X1 U5980 ( .A1(n4803), .A2(n6328), .B1(n5102), .B2(n3082), .ZN(n4827)
         );
  OAI22_X1 U5981 ( .A1(n6407), .A2(n4827), .B1(n4894), .B2(n4826), .ZN(n4804)
         );
  AOI21_X1 U5982 ( .B1(n6404), .B2(n4829), .A(n4804), .ZN(n4805) );
  OAI211_X1 U5983 ( .C1(n6304), .C2(n4832), .A(n4806), .B(n4805), .ZN(U3024)
         );
  NAND2_X1 U5984 ( .A1(n4825), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4809) );
  OAI22_X1 U5985 ( .A1(n6387), .A2(n4827), .B1(n4936), .B2(n4826), .ZN(n4807)
         );
  AOI21_X1 U5986 ( .B1(n6384), .B2(n4829), .A(n4807), .ZN(n4808) );
  OAI211_X1 U5987 ( .C1(n4832), .C2(n6290), .A(n4809), .B(n4808), .ZN(U3020)
         );
  NAND2_X1 U5988 ( .A1(n4825), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4812) );
  OAI22_X1 U5989 ( .A1(n6397), .A2(n4827), .B1(n4868), .B2(n4826), .ZN(n4810)
         );
  AOI21_X1 U5990 ( .B1(n6394), .B2(n4829), .A(n4810), .ZN(n4811) );
  OAI211_X1 U5991 ( .C1(n6297), .C2(n4832), .A(n4812), .B(n4811), .ZN(U3022)
         );
  NAND2_X1 U5992 ( .A1(n4825), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4815) );
  OAI22_X1 U5993 ( .A1(n6393), .A2(n4827), .B1(n4923), .B2(n4826), .ZN(n4813)
         );
  AOI21_X1 U5994 ( .B1(n6390), .B2(n4829), .A(n4813), .ZN(n4814) );
  OAI211_X1 U5995 ( .C1(n6294), .C2(n4832), .A(n4815), .B(n4814), .ZN(U3021)
         );
  NAND2_X1 U5996 ( .A1(n4825), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4818) );
  OAI22_X1 U5997 ( .A1(n6403), .A2(n4827), .B1(n4927), .B2(n4826), .ZN(n4816)
         );
  AOI21_X1 U5998 ( .B1(n6399), .B2(n4829), .A(n4816), .ZN(n4817) );
  OAI211_X1 U5999 ( .C1(n6301), .C2(n4832), .A(n4818), .B(n4817), .ZN(U3023)
         );
  NAND2_X1 U6000 ( .A1(n4825), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4821) );
  OAI22_X1 U6001 ( .A1(n6413), .A2(n4827), .B1(n4931), .B2(n4826), .ZN(n4819)
         );
  AOI21_X1 U6002 ( .B1(n6410), .B2(n4829), .A(n4819), .ZN(n4820) );
  OAI211_X1 U6003 ( .C1(n6308), .C2(n4832), .A(n4821), .B(n4820), .ZN(U3025)
         );
  NAND2_X1 U6004 ( .A1(n4825), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4824) );
  OAI22_X1 U6005 ( .A1(n6419), .A2(n4827), .B1(n4875), .B2(n4826), .ZN(n4822)
         );
  AOI21_X1 U6006 ( .B1(n6415), .B2(n4829), .A(n4822), .ZN(n4823) );
  OAI211_X1 U6007 ( .C1(n6311), .C2(n4832), .A(n4824), .B(n4823), .ZN(U3026)
         );
  NAND2_X1 U6008 ( .A1(n4825), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4831) );
  OAI22_X1 U6009 ( .A1(n6427), .A2(n4827), .B1(n4888), .B2(n4826), .ZN(n4828)
         );
  AOI21_X1 U6010 ( .B1(n6423), .B2(n4829), .A(n4828), .ZN(n4830) );
  OAI211_X1 U6011 ( .C1(n6319), .C2(n4832), .A(n4831), .B(n4830), .ZN(U3027)
         );
  OR2_X1 U6012 ( .A1(n6468), .A2(n5038), .ZN(n5037) );
  NOR2_X1 U6013 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5037), .ZN(n6442)
         );
  NOR3_X1 U6014 ( .A1(n6421), .A2(n6446), .A3(n6586), .ZN(n4835) );
  OAI22_X1 U6015 ( .A1(n4835), .A2(n6280), .B1(n4834), .B2(n5031), .ZN(n4839)
         );
  OAI21_X1 U6016 ( .B1(n3093), .B2(n6481), .A(n4837), .ZN(n4919) );
  NOR2_X1 U6017 ( .A1(n5102), .A2(n4919), .ZN(n4838) );
  NAND2_X1 U6018 ( .A1(n6448), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4843)
         );
  AOI22_X1 U6019 ( .A1(n4840), .A2(n6277), .B1(n3093), .B2(n6275), .ZN(n6429)
         );
  INV_X1 U6020 ( .A(n6442), .ZN(n4853) );
  OAI22_X1 U6021 ( .A1(n6419), .A2(n6429), .B1(n4875), .B2(n4853), .ZN(n4841)
         );
  AOI21_X1 U6022 ( .B1(n6416), .B2(n6446), .A(n4841), .ZN(n4842) );
  OAI211_X1 U6023 ( .C1(n6451), .C2(n6359), .A(n4843), .B(n4842), .ZN(U3122)
         );
  NAND2_X1 U6024 ( .A1(n6448), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4846)
         );
  OAI22_X1 U6025 ( .A1(n6403), .A2(n6429), .B1(n4927), .B2(n4853), .ZN(n4844)
         );
  AOI21_X1 U6026 ( .B1(n6400), .B2(n6446), .A(n4844), .ZN(n4845) );
  OAI211_X1 U6027 ( .C1(n6451), .C2(n5131), .A(n4846), .B(n4845), .ZN(U3119)
         );
  NAND2_X1 U6028 ( .A1(n6448), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4849)
         );
  OAI22_X1 U6029 ( .A1(n6393), .A2(n6429), .B1(n4923), .B2(n4853), .ZN(n4847)
         );
  AOI21_X1 U6030 ( .B1(n6389), .B2(n6446), .A(n4847), .ZN(n4848) );
  OAI211_X1 U6031 ( .C1(n6451), .C2(n5124), .A(n4849), .B(n4848), .ZN(U3117)
         );
  NAND2_X1 U6032 ( .A1(n6448), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4852)
         );
  OAI22_X1 U6033 ( .A1(n6387), .A2(n6429), .B1(n4936), .B2(n4853), .ZN(n4850)
         );
  AOI21_X1 U6034 ( .B1(n6376), .B2(n6446), .A(n4850), .ZN(n4851) );
  OAI211_X1 U6035 ( .C1(n6451), .C2(n5116), .A(n4852), .B(n4851), .ZN(U3116)
         );
  NAND2_X1 U6036 ( .A1(n6448), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4856)
         );
  OAI22_X1 U6037 ( .A1(n6413), .A2(n6429), .B1(n4931), .B2(n4853), .ZN(n4854)
         );
  AOI21_X1 U6038 ( .B1(n6409), .B2(n6446), .A(n4854), .ZN(n4855) );
  OAI211_X1 U6039 ( .C1(n6451), .C2(n5120), .A(n4856), .B(n4855), .ZN(U3121)
         );
  NOR3_X1 U6040 ( .A1(n4859), .A2(n5029), .A3(n6586), .ZN(n4860) );
  OAI21_X1 U6041 ( .B1(n4860), .B2(n6280), .A(n6283), .ZN(n4865) );
  NOR2_X1 U6042 ( .A1(n5102), .A2(n4861), .ZN(n6286) );
  INV_X1 U6043 ( .A(n4862), .ZN(n4863) );
  OR2_X1 U6044 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4863), .ZN(n4893)
         );
  AOI21_X1 U6045 ( .B1(n4893), .B2(STATE2_REG_3__SCAN_IN), .A(n6468), .ZN(
        n4864) );
  NAND3_X1 U6046 ( .A1(n4865), .A2(n6286), .A3(n4864), .ZN(n4892) );
  NAND2_X1 U6047 ( .A1(n4892), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4871)
         );
  NOR2_X1 U6048 ( .A1(n6283), .A2(n6586), .ZN(n6273) );
  INV_X1 U6049 ( .A(n6275), .ZN(n4866) );
  NOR2_X1 U6050 ( .A1(n4866), .A2(n6468), .ZN(n4867) );
  AOI22_X1 U6051 ( .A1(n6273), .A2(n6277), .B1(n6274), .B2(n4867), .ZN(n4895)
         );
  OAI22_X1 U6052 ( .A1(n6397), .A2(n4895), .B1(n4868), .B2(n4893), .ZN(n4869)
         );
  AOI21_X1 U6053 ( .B1(n6394), .B2(n5029), .A(n4869), .ZN(n4870) );
  OAI211_X1 U6054 ( .C1(n4899), .C2(n6297), .A(n4871), .B(n4870), .ZN(U3134)
         );
  NAND2_X1 U6055 ( .A1(n4892), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4874)
         );
  OAI22_X1 U6056 ( .A1(n6403), .A2(n4895), .B1(n4927), .B2(n4893), .ZN(n4872)
         );
  AOI21_X1 U6057 ( .B1(n6399), .B2(n5029), .A(n4872), .ZN(n4873) );
  OAI211_X1 U6058 ( .C1(n4899), .C2(n6301), .A(n4874), .B(n4873), .ZN(U3135)
         );
  NAND2_X1 U6059 ( .A1(n4892), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4878)
         );
  OAI22_X1 U6060 ( .A1(n6419), .A2(n4895), .B1(n4875), .B2(n4893), .ZN(n4876)
         );
  AOI21_X1 U6061 ( .B1(n6415), .B2(n5029), .A(n4876), .ZN(n4877) );
  OAI211_X1 U6062 ( .C1(n4899), .C2(n6311), .A(n4878), .B(n4877), .ZN(U3138)
         );
  NAND2_X1 U6063 ( .A1(n4892), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4881)
         );
  OAI22_X1 U6064 ( .A1(n6393), .A2(n4895), .B1(n4923), .B2(n4893), .ZN(n4879)
         );
  AOI21_X1 U6065 ( .B1(n6390), .B2(n5029), .A(n4879), .ZN(n4880) );
  OAI211_X1 U6066 ( .C1(n4899), .C2(n6294), .A(n4881), .B(n4880), .ZN(U3133)
         );
  NAND2_X1 U6067 ( .A1(n4892), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4884)
         );
  OAI22_X1 U6068 ( .A1(n6413), .A2(n4895), .B1(n4931), .B2(n4893), .ZN(n4882)
         );
  AOI21_X1 U6069 ( .B1(n6410), .B2(n5029), .A(n4882), .ZN(n4883) );
  OAI211_X1 U6070 ( .C1(n4899), .C2(n6308), .A(n4884), .B(n4883), .ZN(U3137)
         );
  NAND2_X1 U6071 ( .A1(n4892), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4887)
         );
  OAI22_X1 U6072 ( .A1(n6387), .A2(n4895), .B1(n4936), .B2(n4893), .ZN(n4885)
         );
  AOI21_X1 U6073 ( .B1(n6384), .B2(n5029), .A(n4885), .ZN(n4886) );
  OAI211_X1 U6074 ( .C1(n4899), .C2(n6290), .A(n4887), .B(n4886), .ZN(U3132)
         );
  NAND2_X1 U6075 ( .A1(n4892), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4891)
         );
  OAI22_X1 U6076 ( .A1(n6427), .A2(n4895), .B1(n4888), .B2(n4893), .ZN(n4889)
         );
  AOI21_X1 U6077 ( .B1(n6423), .B2(n5029), .A(n4889), .ZN(n4890) );
  OAI211_X1 U6078 ( .C1(n4899), .C2(n6319), .A(n4891), .B(n4890), .ZN(U3139)
         );
  NAND2_X1 U6079 ( .A1(n4892), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4898)
         );
  OAI22_X1 U6080 ( .A1(n6407), .A2(n4895), .B1(n4894), .B2(n4893), .ZN(n4896)
         );
  AOI21_X1 U6081 ( .B1(n6404), .B2(n5029), .A(n4896), .ZN(n4897) );
  OAI211_X1 U6082 ( .C1(n4899), .C2(n6304), .A(n4898), .B(n4897), .ZN(U3136)
         );
  AOI21_X1 U6083 ( .B1(n4900), .B2(n4559), .A(n4949), .ZN(n5983) );
  OAI22_X1 U6084 ( .A1(n5522), .A2(n5980), .B1(n5836), .B2(n4901), .ZN(n4902)
         );
  AOI21_X1 U6085 ( .B1(n5983), .B2(n5833), .A(n4902), .ZN(n4903) );
  INV_X1 U6086 ( .A(n4903), .ZN(U2853) );
  INV_X1 U6087 ( .A(n5983), .ZN(n4905) );
  INV_X1 U6088 ( .A(DATAI_6_), .ZN(n6087) );
  OAI222_X1 U6089 ( .A1(n4905), .A2(n5837), .B1(n5526), .B2(n4904), .C1(n5221), 
        .C2(n6087), .ZN(U2885) );
  AND2_X1 U6090 ( .A1(n4906), .A2(n4949), .ZN(n4978) );
  OAI21_X1 U6091 ( .B1(n4978), .B2(n4908), .A(n4907), .ZN(n5249) );
  NAND2_X1 U6092 ( .A1(n4909), .A2(n4997), .ZN(n4911) );
  INV_X1 U6093 ( .A(n4910), .ZN(n5014) );
  NAND2_X1 U6094 ( .A1(n4911), .A2(n5014), .ZN(n6178) );
  OAI22_X1 U6095 ( .A1(n5522), .A2(n6178), .B1(n5836), .B2(n5079), .ZN(n4912)
         );
  INV_X1 U6096 ( .A(n4912), .ZN(n4913) );
  OAI21_X1 U6097 ( .B1(n5249), .B2(n5524), .A(n4913), .ZN(U2848) );
  INV_X1 U6098 ( .A(n6362), .ZN(n4940) );
  NOR3_X1 U6099 ( .A1(n6362), .A2(n6346), .A3(n6586), .ZN(n4915) );
  NOR2_X1 U6100 ( .A1(n4915), .A2(n6280), .ZN(n4921) );
  NOR2_X1 U6101 ( .A1(n4917), .A2(n4916), .ZN(n4922) );
  NOR2_X1 U6102 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4918), .ZN(n6360)
         );
  INV_X1 U6103 ( .A(n6360), .ZN(n4935) );
  AOI211_X1 U6104 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4935), .A(n6275), .B(
        n4919), .ZN(n4920) );
  NAND2_X1 U6105 ( .A1(n6363), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4926) );
  AOI22_X1 U6106 ( .A1(n4922), .A2(n6328), .B1(n5102), .B2(n3093), .ZN(n6351)
         );
  OAI22_X1 U6107 ( .A1(n6393), .A2(n6351), .B1(n4923), .B2(n4935), .ZN(n4924)
         );
  AOI21_X1 U6108 ( .B1(n6390), .B2(n6346), .A(n4924), .ZN(n4925) );
  OAI211_X1 U6109 ( .C1(n4940), .C2(n6294), .A(n4926), .B(n4925), .ZN(U3085)
         );
  NAND2_X1 U6110 ( .A1(n6363), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4930) );
  OAI22_X1 U6111 ( .A1(n6403), .A2(n6351), .B1(n4927), .B2(n4935), .ZN(n4928)
         );
  AOI21_X1 U6112 ( .B1(n6399), .B2(n6346), .A(n4928), .ZN(n4929) );
  OAI211_X1 U6113 ( .C1(n4940), .C2(n6301), .A(n4930), .B(n4929), .ZN(U3087)
         );
  NAND2_X1 U6114 ( .A1(n6363), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4934) );
  OAI22_X1 U6115 ( .A1(n6413), .A2(n6351), .B1(n4931), .B2(n4935), .ZN(n4932)
         );
  AOI21_X1 U6116 ( .B1(n6410), .B2(n6346), .A(n4932), .ZN(n4933) );
  OAI211_X1 U6117 ( .C1(n4940), .C2(n6308), .A(n4934), .B(n4933), .ZN(U3089)
         );
  NAND2_X1 U6118 ( .A1(n6363), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4939) );
  OAI22_X1 U6119 ( .A1(n6387), .A2(n6351), .B1(n4936), .B2(n4935), .ZN(n4937)
         );
  AOI21_X1 U6120 ( .B1(n6384), .B2(n6346), .A(n4937), .ZN(n4938) );
  OAI211_X1 U6121 ( .C1(n4940), .C2(n6290), .A(n4939), .B(n4938), .ZN(U3084)
         );
  AOI21_X1 U6122 ( .B1(n6156), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4941), 
        .ZN(n4942) );
  OAI21_X1 U6123 ( .B1(n6166), .B2(n6021), .A(n4942), .ZN(n4943) );
  AOI21_X1 U6124 ( .B1(n6031), .B2(n6162), .A(n4943), .ZN(n4944) );
  OAI21_X1 U6125 ( .B1(n4945), .B2(n5914), .A(n4944), .ZN(U2983) );
  INV_X1 U6126 ( .A(n4994), .ZN(n4946) );
  NAND2_X1 U6127 ( .A1(n4754), .A2(n4946), .ZN(n4950) );
  NOR2_X1 U6128 ( .A1(n4950), .A2(n4947), .ZN(n4948) );
  AND2_X1 U6129 ( .A1(n4949), .A2(n4948), .ZN(n4976) );
  NOR2_X1 U6130 ( .A1(n4752), .A2(n4950), .ZN(n4992) );
  NOR2_X1 U6131 ( .A1(n4992), .A2(n4951), .ZN(n4952) );
  NAND2_X1 U6132 ( .A1(n4953), .A2(n4968), .ZN(n4955) );
  INV_X1 U6133 ( .A(n4998), .ZN(n4954) );
  NAND2_X1 U6134 ( .A1(n4955), .A2(n4954), .ZN(n6187) );
  OAI22_X1 U6135 ( .A1(n5522), .A2(n6187), .B1(n5836), .B2(n4956), .ZN(n4957)
         );
  INV_X1 U6136 ( .A(n4957), .ZN(n4958) );
  OAI21_X1 U6137 ( .B1(n5206), .B2(n5524), .A(n4958), .ZN(U2850) );
  INV_X1 U6138 ( .A(DATAI_11_), .ZN(n6631) );
  INV_X1 U6139 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6142) );
  OAI222_X1 U6140 ( .A1(n5249), .A2(n5837), .B1(n5221), .B2(n6631), .C1(n5526), 
        .C2(n6142), .ZN(U2880) );
  INV_X1 U6141 ( .A(DATAI_9_), .ZN(n4959) );
  INV_X1 U6142 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6136) );
  OAI222_X1 U6143 ( .A1(n5206), .A2(n5837), .B1(n5221), .B2(n4959), .C1(n5526), 
        .C2(n6136), .ZN(U2882) );
  XNOR2_X1 U6144 ( .A(n4960), .B(n4961), .ZN(n5006) );
  NOR2_X1 U6145 ( .A1(n4963), .A2(n4962), .ZN(n4966) );
  NOR2_X1 U6146 ( .A1(n5739), .A2(n4971), .ZN(n4964) );
  OR2_X1 U6147 ( .A1(n5733), .A2(n4964), .ZN(n4965) );
  OR2_X1 U6148 ( .A1(n4966), .A2(n4965), .ZN(n5170) );
  OR2_X1 U6149 ( .A1(n4967), .A2(n4756), .ZN(n4969) );
  NAND2_X1 U6150 ( .A1(n4969), .A2(n4968), .ZN(n5952) );
  NAND2_X1 U6151 ( .A1(n6215), .A2(REIP_REG_8__SCAN_IN), .ZN(n5002) );
  OAI21_X1 U6152 ( .B1(n6225), .B2(n5952), .A(n5002), .ZN(n4973) );
  NAND2_X1 U6153 ( .A1(n4971), .A2(n4970), .ZN(n6199) );
  AOI211_X1 U6154 ( .C1(n6203), .C2(n4182), .A(n5171), .B(n6199), .ZN(n4972)
         );
  AOI211_X1 U6155 ( .C1(INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n5170), .A(n4973), 
        .B(n4972), .ZN(n4974) );
  OAI21_X1 U6156 ( .B1(n5779), .B2(n5006), .A(n4974), .ZN(U3010) );
  NOR2_X1 U6157 ( .A1(n4976), .A2(n4975), .ZN(n4977) );
  INV_X1 U6158 ( .A(DATAI_10_), .ZN(n6640) );
  INV_X1 U6159 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6139) );
  OAI222_X1 U6160 ( .A1(n5177), .A2(n5837), .B1(n5221), .B2(n6640), .C1(n5526), 
        .C2(n6139), .ZN(U2881) );
  AOI21_X1 U6161 ( .B1(n6156), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4979), 
        .ZN(n4982) );
  INV_X1 U6162 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4980) );
  NAND2_X1 U6163 ( .A1(n5642), .A2(n4980), .ZN(n4981) );
  OAI211_X1 U6164 ( .C1(n4983), .C2(n5914), .A(n4982), .B(n4981), .ZN(n4984)
         );
  INV_X1 U6165 ( .A(n4984), .ZN(n4985) );
  OAI21_X1 U6166 ( .B1(n6175), .B2(n5096), .A(n4985), .ZN(U2985) );
  NAND2_X1 U6167 ( .A1(n4986), .A2(n6173), .ZN(n4991) );
  NOR2_X1 U6168 ( .A1(n6166), .A2(n4987), .ZN(n4988) );
  AOI211_X1 U6169 ( .C1(n6156), .C2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4989), 
        .B(n4988), .ZN(n4990) );
  OAI211_X1 U6170 ( .C1(n6175), .C2(n5991), .A(n4991), .B(n4990), .ZN(U2981)
         );
  AOI21_X1 U6171 ( .B1(n4994), .B2(n4993), .A(n4992), .ZN(n5957) );
  OAI22_X1 U6172 ( .A1(n5522), .A2(n5952), .B1(n5836), .B2(n5953), .ZN(n4995)
         );
  AOI21_X1 U6173 ( .B1(n5957), .B2(n5833), .A(n4995), .ZN(n4996) );
  INV_X1 U6174 ( .A(n4996), .ZN(U2851) );
  OAI21_X1 U6175 ( .B1(n4999), .B2(n4998), .A(n4997), .ZN(n5172) );
  OAI222_X1 U6176 ( .A1(n5172), .A2(n5522), .B1(n5836), .B2(n4191), .C1(n5177), 
        .C2(n5524), .ZN(U2849) );
  INV_X1 U6177 ( .A(n5957), .ZN(n5000) );
  INV_X1 U6178 ( .A(DATAI_8_), .ZN(n6661) );
  INV_X1 U6179 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6133) );
  OAI222_X1 U6180 ( .A1(n5000), .A2(n5837), .B1(n5221), .B2(n6661), .C1(n5526), 
        .C2(n6133), .ZN(U2883) );
  NAND2_X1 U6181 ( .A1(n6156), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5001)
         );
  OAI211_X1 U6182 ( .C1(n6166), .C2(n5003), .A(n5002), .B(n5001), .ZN(n5004)
         );
  AOI21_X1 U6183 ( .B1(n5957), .B2(n6162), .A(n5004), .ZN(n5005) );
  OAI21_X1 U6184 ( .B1(n5914), .B2(n5006), .A(n5005), .ZN(U2978) );
  INV_X1 U6185 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6533) );
  OAI21_X1 U6186 ( .B1(n5963), .B2(n5019), .A(n5962), .ZN(n5960) );
  AOI22_X1 U6187 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6018), .B1(
        PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n5978), .ZN(n5007) );
  OAI211_X1 U6188 ( .C1(n6533), .C2(n5960), .A(n5007), .B(n5967), .ZN(n5010)
         );
  NOR3_X1 U6189 ( .A1(n5965), .A2(n5019), .A3(REIP_REG_9__SCAN_IN), .ZN(n5009)
         );
  OAI22_X1 U6190 ( .A1(n6009), .A2(n6187), .B1(n5202), .B2(n6022), .ZN(n5008)
         );
  NOR3_X1 U6191 ( .A1(n5010), .A2(n5009), .A3(n5008), .ZN(n5011) );
  OAI21_X1 U6192 ( .B1(n5206), .B2(n5971), .A(n5011), .ZN(U2818) );
  AOI21_X1 U6193 ( .B1(n5013), .B2(n4907), .A(n5012), .ZN(n5947) );
  INV_X1 U6194 ( .A(n5947), .ZN(n5018) );
  INV_X1 U6195 ( .A(DATAI_12_), .ZN(n6625) );
  OAI222_X1 U6196 ( .A1(n5018), .A2(n5837), .B1(n5221), .B2(n6625), .C1(n5526), 
        .C2(n3737), .ZN(U2879) );
  XNOR2_X1 U6197 ( .A(n5015), .B(n5014), .ZN(n5942) );
  INV_X1 U6198 ( .A(n5942), .ZN(n5016) );
  OAI222_X1 U6199 ( .A1(n5018), .A2(n5524), .B1(n5017), .B2(n5836), .C1(n5522), 
        .C2(n5016), .ZN(U2847) );
  INV_X1 U6200 ( .A(n5172), .ZN(n5027) );
  INV_X1 U6201 ( .A(n5019), .ZN(n5021) );
  OAI211_X1 U6202 ( .C1(REIP_REG_10__SCAN_IN), .C2(REIP_REG_9__SCAN_IN), .A(
        n5021), .B(n5020), .ZN(n5023) );
  INV_X1 U6203 ( .A(n5180), .ZN(n5022) );
  OAI22_X1 U6204 ( .A1(n5965), .A2(n5023), .B1(n6022), .B2(n5022), .ZN(n5026)
         );
  INV_X1 U6205 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6535) );
  AOI22_X1 U6206 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6018), .B1(
        PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n5978), .ZN(n5024) );
  OAI211_X1 U6207 ( .C1(n6535), .C2(n5960), .A(n5024), .B(n5967), .ZN(n5025)
         );
  AOI211_X1 U6208 ( .C1(n5027), .C2(n6020), .A(n5026), .B(n5025), .ZN(n5028)
         );
  OAI21_X1 U6209 ( .B1(n5177), .B2(n5971), .A(n5028), .ZN(U2817) );
  INV_X1 U6210 ( .A(n5030), .ZN(n5033) );
  INV_X1 U6211 ( .A(n5031), .ZN(n5032) );
  NOR2_X1 U6212 ( .A1(n6454), .A2(n5037), .ZN(n5069) );
  AOI21_X1 U6213 ( .B1(n5033), .B2(n5032), .A(n5069), .ZN(n5040) );
  NAND2_X1 U6214 ( .A1(n5040), .A2(n5034), .ZN(n5035) );
  NOR2_X1 U6215 ( .A1(n6586), .A2(n5035), .ZN(n5036) );
  AOI211_X2 U6216 ( .C1(n6586), .C2(n5037), .A(n5036), .B(n6379), .ZN(n5073)
         );
  INV_X1 U6217 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n5042) );
  NAND2_X1 U6218 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5039) );
  OAI22_X1 U6219 ( .A1(n5040), .A2(n6586), .B1(n5039), .B2(n5038), .ZN(n5070)
         );
  AOI22_X1 U6220 ( .A1(n6356), .A2(n5070), .B1(n6414), .B2(n5069), .ZN(n5041)
         );
  OAI21_X1 U6221 ( .B1(n5073), .B2(n5042), .A(n5041), .ZN(n5043) );
  AOI21_X1 U6222 ( .B1(n6415), .B2(n6446), .A(n5043), .ZN(n5044) );
  OAI21_X1 U6223 ( .B1(n6311), .B2(n5076), .A(n5044), .ZN(U3130) );
  INV_X1 U6224 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n5046) );
  AOI22_X1 U6225 ( .A1(n6445), .A2(n5070), .B1(n6443), .B2(n5069), .ZN(n5045)
         );
  OAI21_X1 U6226 ( .B1(n5073), .B2(n5046), .A(n5045), .ZN(n5047) );
  AOI21_X1 U6227 ( .B1(n6423), .B2(n6446), .A(n5047), .ZN(n5048) );
  OAI21_X1 U6228 ( .B1(n6319), .B2(n5076), .A(n5048), .ZN(U3131) );
  INV_X1 U6229 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n5050) );
  AOI22_X1 U6230 ( .A1(n6431), .A2(n5070), .B1(n6430), .B2(n5069), .ZN(n5049)
         );
  OAI21_X1 U6231 ( .B1(n5073), .B2(n5050), .A(n5049), .ZN(n5051) );
  AOI21_X1 U6232 ( .B1(n6394), .B2(n6446), .A(n5051), .ZN(n5052) );
  OAI21_X1 U6233 ( .B1(n6297), .B2(n5076), .A(n5052), .ZN(U3126) );
  INV_X1 U6234 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n5054) );
  AOI22_X1 U6235 ( .A1(n6279), .A2(n5070), .B1(n6375), .B2(n5069), .ZN(n5053)
         );
  OAI21_X1 U6236 ( .B1(n5073), .B2(n5054), .A(n5053), .ZN(n5055) );
  AOI21_X1 U6237 ( .B1(n6384), .B2(n6446), .A(n5055), .ZN(n5056) );
  OAI21_X1 U6238 ( .B1(n6290), .B2(n5076), .A(n5056), .ZN(U3124) );
  INV_X1 U6239 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n5058) );
  AOI22_X1 U6240 ( .A1(n6291), .A2(n5070), .B1(n6388), .B2(n5069), .ZN(n5057)
         );
  OAI21_X1 U6241 ( .B1(n5073), .B2(n5058), .A(n5057), .ZN(n5059) );
  AOI21_X1 U6242 ( .B1(n6390), .B2(n6446), .A(n5059), .ZN(n5060) );
  OAI21_X1 U6243 ( .B1(n6294), .B2(n5076), .A(n5060), .ZN(U3125) );
  INV_X1 U6244 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n5062) );
  AOI22_X1 U6245 ( .A1(n6437), .A2(n5070), .B1(n6436), .B2(n5069), .ZN(n5061)
         );
  OAI21_X1 U6246 ( .B1(n5073), .B2(n5062), .A(n5061), .ZN(n5063) );
  AOI21_X1 U6247 ( .B1(n6404), .B2(n6446), .A(n5063), .ZN(n5064) );
  OAI21_X1 U6248 ( .B1(n6304), .B2(n5076), .A(n5064), .ZN(U3128) );
  INV_X1 U6249 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n5066) );
  AOI22_X1 U6250 ( .A1(n6305), .A2(n5070), .B1(n6408), .B2(n5069), .ZN(n5065)
         );
  OAI21_X1 U6251 ( .B1(n5073), .B2(n5066), .A(n5065), .ZN(n5067) );
  AOI21_X1 U6252 ( .B1(n6410), .B2(n6446), .A(n5067), .ZN(n5068) );
  OAI21_X1 U6253 ( .B1(n6308), .B2(n5076), .A(n5068), .ZN(U3129) );
  INV_X1 U6254 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n5072) );
  AOI22_X1 U6255 ( .A1(n6298), .A2(n5070), .B1(n6398), .B2(n5069), .ZN(n5071)
         );
  OAI21_X1 U6256 ( .B1(n5073), .B2(n5072), .A(n5071), .ZN(n5074) );
  AOI21_X1 U6257 ( .B1(n6399), .B2(n6446), .A(n5074), .ZN(n5075) );
  OAI21_X1 U6258 ( .B1(n6301), .B2(n5076), .A(n5075), .ZN(U3127) );
  INV_X1 U6259 ( .A(n5935), .ZN(n5077) );
  NOR2_X1 U6260 ( .A1(n5965), .A2(n5077), .ZN(n5083) );
  OAI22_X1 U6261 ( .A1(n6009), .A2(n6178), .B1(n5245), .B2(n6022), .ZN(n5081)
         );
  NOR2_X1 U6262 ( .A1(n5963), .A2(n5083), .ZN(n5943) );
  INV_X1 U6263 ( .A(n5943), .ZN(n5936) );
  AOI22_X1 U6264 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n5978), .B1(
        REIP_REG_11__SCAN_IN), .B2(n5936), .ZN(n5078) );
  OAI211_X1 U6265 ( .C1(n5954), .C2(n5079), .A(n5078), .B(n5967), .ZN(n5080)
         );
  AOI211_X1 U6266 ( .C1(n5083), .C2(n5082), .A(n5081), .B(n5080), .ZN(n5084)
         );
  OAI21_X1 U6267 ( .B1(n5249), .B2(n5971), .A(n5084), .ZN(U2816) );
  OAI21_X1 U6268 ( .B1(n5089), .B2(n3545), .A(n5971), .ZN(n6030) );
  INV_X1 U6269 ( .A(n6030), .ZN(n5213) );
  INV_X1 U6270 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5085) );
  NAND2_X1 U6271 ( .A1(n6005), .A2(n5085), .ZN(n5155) );
  INV_X1 U6272 ( .A(n5155), .ZN(n5094) );
  INV_X1 U6273 ( .A(n5086), .ZN(n5090) );
  INV_X1 U6274 ( .A(n5087), .ZN(n5088) );
  NOR2_X1 U6275 ( .A1(n5089), .A2(n5088), .ZN(n6026) );
  AOI22_X1 U6276 ( .A1(n6020), .A2(n5090), .B1(n6026), .B2(n2983), .ZN(n5092)
         );
  AOI22_X1 U6277 ( .A1(n5978), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n5963), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5091) );
  OAI211_X1 U6278 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6022), .A(n5092), 
        .B(n5091), .ZN(n5093) );
  AOI211_X1 U6279 ( .C1(n6018), .C2(EBX_REG_1__SCAN_IN), .A(n5094), .B(n5093), 
        .ZN(n5095) );
  OAI21_X1 U6280 ( .B1(n5213), .B2(n5096), .A(n5095), .ZN(U2826) );
  NAND2_X1 U6281 ( .A1(n3029), .A2(n5097), .ZN(n6271) );
  NAND3_X1 U6282 ( .A1(n5105), .A2(n5140), .A3(n6328), .ZN(n5099) );
  INV_X1 U6283 ( .A(n6280), .ZN(n5098) );
  NAND2_X1 U6284 ( .A1(n5099), .A2(n5098), .ZN(n5108) );
  INV_X1 U6285 ( .A(n5100), .ZN(n5101) );
  INV_X1 U6286 ( .A(n5102), .ZN(n5103) );
  NOR2_X1 U6287 ( .A1(n5103), .A2(n6468), .ZN(n5104) );
  NOR3_X1 U6288 ( .A1(n6468), .A2(n5106), .A3(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), 
        .ZN(n6378) );
  NAND2_X1 U6289 ( .A1(n6454), .A2(n6378), .ZN(n5109) );
  INV_X1 U6290 ( .A(n5109), .ZN(n5138) );
  INV_X1 U6291 ( .A(n6371), .ZN(n5107) );
  AOI22_X1 U6292 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n5109), .B1(n5108), .B2(
        n5107), .ZN(n5110) );
  OAI211_X1 U6293 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6481), .A(n5111), .B(n5110), .ZN(n5137) );
  AOI22_X1 U6294 ( .A1(n6443), .A2(n5138), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5137), .ZN(n5112) );
  OAI21_X1 U6295 ( .B1(n6452), .B2(n5140), .A(n5112), .ZN(n5113) );
  AOI21_X1 U6296 ( .B1(n6447), .B2(n6422), .A(n5113), .ZN(n5114) );
  OAI21_X1 U6297 ( .B1(n5143), .B2(n6427), .A(n5114), .ZN(U3107) );
  AOI22_X1 U6298 ( .A1(n6375), .A2(n5138), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5137), .ZN(n5115) );
  OAI21_X1 U6299 ( .B1(n5116), .B2(n5140), .A(n5115), .ZN(n5117) );
  AOI21_X1 U6300 ( .B1(n6376), .B2(n6422), .A(n5117), .ZN(n5118) );
  OAI21_X1 U6301 ( .B1(n5143), .B2(n6387), .A(n5118), .ZN(U3100) );
  AOI22_X1 U6302 ( .A1(n6408), .A2(n5138), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5137), .ZN(n5119) );
  OAI21_X1 U6303 ( .B1(n5120), .B2(n5140), .A(n5119), .ZN(n5121) );
  AOI21_X1 U6304 ( .B1(n6409), .B2(n6422), .A(n5121), .ZN(n5122) );
  OAI21_X1 U6305 ( .B1(n5143), .B2(n6413), .A(n5122), .ZN(U3105) );
  AOI22_X1 U6306 ( .A1(n6388), .A2(n5138), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5137), .ZN(n5123) );
  OAI21_X1 U6307 ( .B1(n5124), .B2(n5140), .A(n5123), .ZN(n5125) );
  AOI21_X1 U6308 ( .B1(n6389), .B2(n6422), .A(n5125), .ZN(n5126) );
  OAI21_X1 U6309 ( .B1(n5143), .B2(n6393), .A(n5126), .ZN(U3101) );
  AOI22_X1 U6310 ( .A1(n6414), .A2(n5138), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5137), .ZN(n5127) );
  OAI21_X1 U6311 ( .B1(n6359), .B2(n5140), .A(n5127), .ZN(n5128) );
  AOI21_X1 U6312 ( .B1(n6416), .B2(n6422), .A(n5128), .ZN(n5129) );
  OAI21_X1 U6313 ( .B1(n5143), .B2(n6419), .A(n5129), .ZN(U3106) );
  AOI22_X1 U6314 ( .A1(n6398), .A2(n5138), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5137), .ZN(n5130) );
  OAI21_X1 U6315 ( .B1(n5131), .B2(n5140), .A(n5130), .ZN(n5132) );
  AOI21_X1 U6316 ( .B1(n6400), .B2(n6422), .A(n5132), .ZN(n5133) );
  OAI21_X1 U6317 ( .B1(n5143), .B2(n6403), .A(n5133), .ZN(U3103) );
  AOI22_X1 U6318 ( .A1(n6436), .A2(n5138), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5137), .ZN(n5134) );
  OAI21_X1 U6319 ( .B1(n6441), .B2(n5140), .A(n5134), .ZN(n5135) );
  AOI21_X1 U6320 ( .B1(n6438), .B2(n6422), .A(n5135), .ZN(n5136) );
  OAI21_X1 U6321 ( .B1(n5143), .B2(n6407), .A(n5136), .ZN(U3104) );
  AOI22_X1 U6322 ( .A1(n6430), .A2(n5138), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5137), .ZN(n5139) );
  OAI21_X1 U6323 ( .B1(n6435), .B2(n5140), .A(n5139), .ZN(n5141) );
  AOI21_X1 U6324 ( .B1(n6432), .B2(n6422), .A(n5141), .ZN(n5142) );
  OAI21_X1 U6325 ( .B1(n5143), .B2(n6397), .A(n5142), .ZN(U3102) );
  AOI22_X1 U6326 ( .A1(n6156), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .B1(n6215), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n5144) );
  OAI21_X1 U6327 ( .B1(n6166), .B2(n5986), .A(n5144), .ZN(n5145) );
  AOI21_X1 U6328 ( .B1(n5983), .B2(n6162), .A(n5145), .ZN(n5146) );
  OAI21_X1 U6329 ( .B1(n5914), .B2(n5147), .A(n5146), .ZN(U2980) );
  INV_X1 U6330 ( .A(n5148), .ZN(n6015) );
  AOI21_X1 U6331 ( .B1(n6156), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5149), 
        .ZN(n5150) );
  OAI21_X1 U6332 ( .B1(n6166), .B2(n6015), .A(n5150), .ZN(n5151) );
  AOI21_X1 U6333 ( .B1(n6012), .B2(n6162), .A(n5151), .ZN(n5152) );
  OAI21_X1 U6334 ( .B1(n5914), .B2(n5153), .A(n5152), .ZN(U2982) );
  INV_X1 U6335 ( .A(n5154), .ZN(n6161) );
  NOR2_X1 U6336 ( .A1(n6009), .A2(n6205), .ZN(n5163) );
  NAND2_X1 U6337 ( .A1(n5155), .A2(n5999), .ZN(n6017) );
  NAND2_X1 U6338 ( .A1(n6017), .A2(REIP_REG_2__SCAN_IN), .ZN(n5161) );
  INV_X1 U6339 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5156) );
  OAI22_X1 U6340 ( .A1(n6165), .A2(n6022), .B1(n6023), .B2(n5156), .ZN(n5157)
         );
  INV_X1 U6341 ( .A(n5157), .ZN(n5160) );
  AOI22_X1 U6342 ( .A1(EBX_REG_2__SCAN_IN), .A2(n6018), .B1(n6026), .B2(n3021), 
        .ZN(n5159) );
  INV_X1 U6343 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6016) );
  NAND3_X1 U6344 ( .A1(n6005), .A2(REIP_REG_1__SCAN_IN), .A3(n6016), .ZN(n5158) );
  NAND4_X1 U6345 ( .A1(n5161), .A2(n5160), .A3(n5159), .A4(n5158), .ZN(n5162)
         );
  AOI211_X1 U6346 ( .C1(n6161), .C2(n6030), .A(n5163), .B(n5162), .ZN(n5164)
         );
  INV_X1 U6347 ( .A(n5164), .ZN(U2825) );
  NAND2_X1 U6348 ( .A1(n3034), .A2(n5166), .ZN(n5167) );
  XNOR2_X1 U6349 ( .A(n5165), .B(n5167), .ZN(n5182) );
  NOR2_X1 U6350 ( .A1(n5168), .A2(n6199), .ZN(n6190) );
  OAI211_X1 U6351 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6190), .B(n5169), .ZN(n5175) );
  INV_X1 U6352 ( .A(n5170), .ZN(n6204) );
  OAI21_X1 U6353 ( .B1(n5171), .B2(n5740), .A(n6204), .ZN(n6186) );
  OAI22_X1 U6354 ( .A1(n6225), .A2(n5172), .B1(n6535), .B2(n5900), .ZN(n5173)
         );
  AOI21_X1 U6355 ( .B1(n6186), .B2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n5173), 
        .ZN(n5174) );
  OAI211_X1 U6356 ( .C1(n5182), .C2(n5779), .A(n5175), .B(n5174), .ZN(U3008)
         );
  INV_X1 U6357 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5176) );
  OAI22_X1 U6358 ( .A1(n6171), .A2(n5176), .B1(n5900), .B2(n6535), .ZN(n5179)
         );
  NOR2_X1 U6359 ( .A1(n5177), .A2(n6175), .ZN(n5178) );
  AOI211_X1 U6360 ( .C1(n5642), .C2(n5180), .A(n5179), .B(n5178), .ZN(n5181)
         );
  OAI21_X1 U6361 ( .B1(n5914), .B2(n5182), .A(n5181), .ZN(U2976) );
  OAI21_X1 U6362 ( .B1(n5183), .B2(n5185), .A(n5184), .ZN(n5648) );
  AOI22_X1 U6363 ( .A1(n5225), .A2(DATAI_14_), .B1(n6045), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5186) );
  OAI21_X1 U6364 ( .B1(n5648), .B2(n5837), .A(n5186), .ZN(U2877) );
  AND2_X1 U6365 ( .A1(n5962), .A2(n5187), .ZN(n5271) );
  OAI21_X1 U6366 ( .B1(n5188), .B2(n5216), .A(n5227), .ZN(n5901) );
  OAI22_X1 U6367 ( .A1(n6009), .A2(n5901), .B1(n5650), .B2(n6022), .ZN(n5193)
         );
  INV_X1 U6368 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5191) );
  AOI22_X1 U6369 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6018), .B1(n5189), .B2(n6540), .ZN(n5190) );
  OAI211_X1 U6370 ( .C1(n6023), .C2(n5191), .A(n5190), .B(n5967), .ZN(n5192)
         );
  AOI211_X1 U6371 ( .C1(n5271), .C2(REIP_REG_14__SCAN_IN), .A(n5193), .B(n5192), .ZN(n5194) );
  OAI21_X1 U6372 ( .B1(n5648), .B2(n5971), .A(n5194), .ZN(U2813) );
  XOR2_X1 U6373 ( .A(n5196), .B(n2987), .Z(n6201) );
  NAND2_X1 U6374 ( .A1(n6201), .A2(n6173), .ZN(n5199) );
  INV_X1 U6375 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6530) );
  NOR2_X1 U6376 ( .A1(n5900), .A2(n6530), .ZN(n6196) );
  NOR2_X1 U6377 ( .A1(n6166), .A2(n5970), .ZN(n5197) );
  AOI211_X1 U6378 ( .C1(n6156), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6196), 
        .B(n5197), .ZN(n5198) );
  OAI211_X1 U6379 ( .C1(n6175), .C2(n5972), .A(n5199), .B(n5198), .ZN(U2979)
         );
  XNOR2_X1 U6380 ( .A(n2992), .B(n6194), .ZN(n5201) );
  XNOR2_X1 U6381 ( .A(n5200), .B(n5201), .ZN(n6191) );
  NAND2_X1 U6382 ( .A1(n6191), .A2(n6173), .ZN(n5205) );
  NOR2_X1 U6383 ( .A1(n5900), .A2(n6533), .ZN(n6188) );
  NOR2_X1 U6384 ( .A1(n6166), .A2(n5202), .ZN(n5203) );
  AOI211_X1 U6385 ( .C1(n6156), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6188), 
        .B(n5203), .ZN(n5204) );
  OAI211_X1 U6386 ( .C1(n6175), .C2(n5206), .A(n5205), .B(n5204), .ZN(U2977)
         );
  INV_X1 U6387 ( .A(n6026), .ZN(n5208) );
  OAI21_X1 U6388 ( .B1(n5978), .B2(n5993), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5207) );
  OAI21_X1 U6389 ( .B1(n5208), .B2(n3617), .A(n5207), .ZN(n5211) );
  OAI22_X1 U6390 ( .A1(n5954), .A2(n5209), .B1(n6009), .B2(n6224), .ZN(n5210)
         );
  AOI211_X1 U6391 ( .C1(REIP_REG_0__SCAN_IN), .C2(n5962), .A(n5211), .B(n5210), 
        .ZN(n5212) );
  OAI21_X1 U6392 ( .B1(n5213), .B2(n6176), .A(n5212), .ZN(U2827) );
  OAI222_X1 U6393 ( .A1(n5648), .A2(n5524), .B1(n5836), .B2(n4206), .C1(n5901), 
        .C2(n5522), .ZN(U2845) );
  XOR2_X1 U6394 ( .A(n5215), .B(n2998), .Z(n5934) );
  AOI21_X1 U6395 ( .B1(n5218), .B2(n5217), .A(n5216), .ZN(n5308) );
  INV_X1 U6396 ( .A(n5308), .ZN(n5929) );
  OAI22_X1 U6397 ( .A1(n5522), .A2(n5929), .B1(n5836), .B2(n5930), .ZN(n5219)
         );
  AOI21_X1 U6398 ( .B1(n5934), .B2(n5833), .A(n5219), .ZN(n5220) );
  INV_X1 U6399 ( .A(n5220), .ZN(U2846) );
  INV_X1 U6400 ( .A(n5934), .ZN(n5222) );
  INV_X1 U6401 ( .A(DATAI_13_), .ZN(n6720) );
  INV_X1 U6402 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6147) );
  OAI222_X1 U6403 ( .A1(n5837), .A2(n5222), .B1(n5221), .B2(n6720), .C1(n5526), 
        .C2(n6147), .ZN(U2878) );
  OAI21_X1 U6404 ( .B1(n3062), .B2(n3805), .A(n5224), .ZN(n5645) );
  AOI22_X1 U6405 ( .A1(n5225), .A2(DATAI_15_), .B1(n6045), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5226) );
  OAI21_X1 U6406 ( .B1(n5645), .B2(n5837), .A(n5226), .ZN(U2876) );
  INV_X1 U6407 ( .A(n5285), .ZN(n5234) );
  INV_X1 U6408 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5639) );
  INV_X1 U6409 ( .A(n5227), .ZN(n5228) );
  XNOR2_X1 U6410 ( .A(n5229), .B(n5228), .ZN(n5889) );
  INV_X1 U6411 ( .A(n5889), .ZN(n5237) );
  OAI22_X1 U6412 ( .A1(n6009), .A2(n5237), .B1(n6022), .B2(n5230), .ZN(n5233)
         );
  AOI22_X1 U6413 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n5978), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5271), .ZN(n5231) );
  OAI211_X1 U6414 ( .C1(n5954), .C2(n5236), .A(n5231), .B(n5967), .ZN(n5232)
         );
  AOI211_X1 U6415 ( .C1(n5234), .C2(n5639), .A(n5233), .B(n5232), .ZN(n5235)
         );
  OAI21_X1 U6416 ( .B1(n5645), .B2(n5971), .A(n5235), .ZN(U2812) );
  OAI22_X1 U6417 ( .A1(n5522), .A2(n5237), .B1(n5836), .B2(n5236), .ZN(n5238)
         );
  INV_X1 U6418 ( .A(n5238), .ZN(n5239) );
  OAI21_X1 U6419 ( .B1(n5645), .B2(n5524), .A(n5239), .ZN(U2844) );
  NAND2_X1 U6420 ( .A1(n5242), .A2(n5241), .ZN(n5243) );
  XNOR2_X1 U6421 ( .A(n5240), .B(n5243), .ZN(n6181) );
  NAND2_X1 U6422 ( .A1(n6181), .A2(n6173), .ZN(n5248) );
  INV_X1 U6423 ( .A(REIP_REG_11__SCAN_IN), .ZN(n5244) );
  NOR2_X1 U6424 ( .A1(n5900), .A2(n5244), .ZN(n6179) );
  NOR2_X1 U6425 ( .A1(n6166), .A2(n5245), .ZN(n5246) );
  AOI211_X1 U6426 ( .C1(n6156), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6179), 
        .B(n5246), .ZN(n5247) );
  OAI211_X1 U6427 ( .C1(n6175), .C2(n5249), .A(n5248), .B(n5247), .ZN(U2975)
         );
  INV_X1 U6428 ( .A(n5251), .ZN(n5252) );
  NOR2_X1 U6429 ( .A1(n5253), .A2(n5252), .ZN(n5254) );
  XNOR2_X1 U6430 ( .A(n2986), .B(n5254), .ZN(n5265) );
  NOR2_X1 U6431 ( .A1(n5900), .A2(n6538), .ZN(n5262) );
  AOI21_X1 U6432 ( .B1(n6156), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n5262), 
        .ZN(n5255) );
  OAI21_X1 U6433 ( .B1(n6166), .B2(n5256), .A(n5255), .ZN(n5257) );
  AOI21_X1 U6434 ( .B1(n5947), .B2(n6162), .A(n5257), .ZN(n5258) );
  OAI21_X1 U6435 ( .B1(n5265), .B2(n5914), .A(n5258), .ZN(U2974) );
  AOI21_X1 U6436 ( .B1(n5735), .B2(n5736), .A(n5733), .ZN(n5259) );
  OAI21_X1 U6437 ( .B1(n5260), .B2(n5739), .A(n5259), .ZN(n6182) );
  XOR2_X1 U6438 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .B(
        INSTADDRPOINTER_REG_11__SCAN_IN), .Z(n5261) );
  AOI22_X1 U6439 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6182), .B1(n6177), .B2(n5261), .ZN(n5264) );
  AOI21_X1 U6440 ( .B1(n6210), .B2(n5942), .A(n5262), .ZN(n5263) );
  OAI211_X1 U6441 ( .C1(n5265), .C2(n5779), .A(n5264), .B(n5263), .ZN(U3006)
         );
  AOI21_X1 U6442 ( .B1(n5267), .B2(n5224), .A(n5266), .ZN(n6044) );
  INV_X1 U6443 ( .A(n6044), .ZN(n5278) );
  OAI21_X1 U6444 ( .B1(n5269), .B2(n5268), .A(n5286), .ZN(n5277) );
  INV_X1 U6445 ( .A(n5277), .ZN(n5777) );
  AOI21_X1 U6446 ( .B1(n5978), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6002), 
        .ZN(n5270) );
  OAI21_X1 U6447 ( .B1(n5634), .B2(n6022), .A(n5270), .ZN(n5275) );
  NAND2_X1 U6448 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n5284) );
  OAI21_X1 U6449 ( .B1(REIP_REG_16__SCAN_IN), .B2(REIP_REG_15__SCAN_IN), .A(
        n5284), .ZN(n5273) );
  AOI22_X1 U6450 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6018), .B1(
        REIP_REG_16__SCAN_IN), .B2(n5271), .ZN(n5272) );
  OAI21_X1 U6451 ( .B1(n5285), .B2(n5273), .A(n5272), .ZN(n5274) );
  AOI211_X1 U6452 ( .C1(n5777), .C2(n6020), .A(n5275), .B(n5274), .ZN(n5276)
         );
  OAI21_X1 U6453 ( .B1(n5278), .B2(n5971), .A(n5276), .ZN(U2811) );
  OAI222_X1 U6454 ( .A1(n5278), .A2(n5524), .B1(n5836), .B2(n4215), .C1(n5277), 
        .C2(n5522), .ZN(U2843) );
  OR2_X1 U6455 ( .A1(n5266), .A2(n5280), .ZN(n5281) );
  AND2_X1 U6456 ( .A1(n5279), .A2(n5281), .ZN(n6039) );
  INV_X1 U6457 ( .A(n6039), .ZN(n5312) );
  NOR2_X1 U6458 ( .A1(n5283), .A2(n5282), .ZN(n5825) );
  INV_X1 U6459 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6544) );
  OAI21_X1 U6460 ( .B1(n5285), .B2(n5284), .A(n6544), .ZN(n5292) );
  AOI21_X1 U6461 ( .B1(n5287), .B2(n5286), .A(n5514), .ZN(n5884) );
  INV_X1 U6462 ( .A(n5884), .ZN(n5314) );
  NAND2_X1 U6463 ( .A1(n6018), .A2(EBX_REG_17__SCAN_IN), .ZN(n5288) );
  OAI211_X1 U6464 ( .C1(n5314), .C2(n6009), .A(n5288), .B(n5967), .ZN(n5291)
         );
  INV_X1 U6465 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5289) );
  OAI22_X1 U6466 ( .A1(n5289), .A2(n6023), .B1(n5873), .B2(n6022), .ZN(n5290)
         );
  AOI211_X1 U6467 ( .C1(n5825), .C2(n5292), .A(n5291), .B(n5290), .ZN(n5293)
         );
  OAI21_X1 U6468 ( .B1(n5312), .B2(n5971), .A(n5293), .ZN(U2810) );
  OAI21_X1 U6469 ( .B1(n5295), .B2(n5297), .A(n3013), .ZN(n5298) );
  INV_X1 U6470 ( .A(n5298), .ZN(n5311) );
  INV_X1 U6471 ( .A(REIP_REG_13__SCAN_IN), .ZN(n5299) );
  NOR2_X1 U6472 ( .A1(n5900), .A2(n5299), .ZN(n5307) );
  AOI21_X1 U6473 ( .B1(n6156), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5307), 
        .ZN(n5300) );
  OAI21_X1 U6474 ( .B1(n6166), .B2(n5932), .A(n5300), .ZN(n5301) );
  AOI21_X1 U6475 ( .B1(n5934), .B2(n6162), .A(n5301), .ZN(n5302) );
  OAI21_X1 U6476 ( .B1(n5311), .B2(n5914), .A(n5302), .ZN(U2973) );
  AOI21_X1 U6477 ( .B1(n5305), .B2(n5303), .A(n6182), .ZN(n5304) );
  OAI21_X1 U6478 ( .B1(n5895), .B2(n6231), .A(n5304), .ZN(n5898) );
  NOR2_X1 U6479 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5305), .ZN(n5306)
         );
  AOI22_X1 U6480 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5898), .B1(n5306), .B2(n6177), .ZN(n5310) );
  AOI21_X1 U6481 ( .B1(n6210), .B2(n5308), .A(n5307), .ZN(n5309) );
  OAI211_X1 U6482 ( .C1(n5311), .C2(n5779), .A(n5310), .B(n5309), .ZN(U3005)
         );
  INV_X1 U6483 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5313) );
  OAI222_X1 U6484 ( .A1(n5314), .A2(n5522), .B1(n5313), .B2(n5836), .C1(n5312), 
        .C2(n5524), .ZN(U2842) );
  INV_X1 U6485 ( .A(n5315), .ZN(n5481) );
  AOI21_X1 U6486 ( .B1(n5316), .B2(n5481), .A(n5366), .ZN(n5548) );
  INV_X1 U6487 ( .A(n5548), .ZN(n5533) );
  INV_X1 U6488 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6660) );
  INV_X1 U6489 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6690) );
  OR3_X1 U6490 ( .A1(n6687), .A2(n6660), .A3(n6690), .ZN(n5321) );
  NOR2_X1 U6491 ( .A1(n5317), .A2(n5321), .ZN(n5797) );
  INV_X1 U6492 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6733) );
  OAI22_X1 U6493 ( .A1(n4059), .A2(n6023), .B1(n6022), .B2(n5546), .ZN(n5328)
         );
  NAND2_X1 U6494 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5324) );
  NAND2_X1 U6495 ( .A1(n5962), .A2(n5321), .ZN(n5322) );
  NAND2_X1 U6496 ( .A1(n5323), .A2(n5322), .ZN(n5806) );
  AOI21_X1 U6497 ( .B1(n6005), .B2(n5324), .A(n5806), .ZN(n5345) );
  OR2_X1 U6498 ( .A1(n5345), .A2(n6733), .ZN(n5326) );
  NAND2_X1 U6499 ( .A1(n6018), .A2(EBX_REG_29__SCAN_IN), .ZN(n5325) );
  NAND2_X1 U6500 ( .A1(n5326), .A2(n5325), .ZN(n5327) );
  AOI21_X1 U6501 ( .B1(n5392), .B2(n6733), .A(n5330), .ZN(n5331) );
  OAI21_X1 U6502 ( .B1(n5533), .B2(n5971), .A(n5331), .ZN(U2798) );
  INV_X1 U6503 ( .A(n5332), .ZN(n5911) );
  INV_X1 U6504 ( .A(n5333), .ZN(n5335) );
  AOI22_X1 U6505 ( .A1(n6370), .A2(n5335), .B1(n5334), .B2(n5343), .ZN(n6453)
         );
  INV_X1 U6506 ( .A(n5340), .ZN(n5338) );
  AOI22_X1 U6507 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6232), .B1(n5343), .B2(
        n5336), .ZN(n5337) );
  OAI21_X1 U6508 ( .B1(n6453), .B2(n5338), .A(n5337), .ZN(n5341) );
  NOR2_X1 U6509 ( .A1(n5339), .A2(n5343), .ZN(n6455) );
  AOI22_X1 U6510 ( .A1(n5911), .A2(n5341), .B1(n5340), .B2(n6455), .ZN(n5342)
         );
  OAI21_X1 U6511 ( .B1(n5343), .B2(n5911), .A(n5342), .ZN(U3461) );
  INV_X1 U6512 ( .A(n5528), .ZN(n5356) );
  INV_X1 U6513 ( .A(n5345), .ZN(n5785) );
  AOI21_X1 U6514 ( .B1(n6005), .B2(n6733), .A(n5785), .ZN(n5382) );
  OAI21_X1 U6515 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5965), .A(n5382), .ZN(n5351) );
  NAND2_X1 U6516 ( .A1(n5978), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5349)
         );
  NAND3_X1 U6517 ( .A1(n5347), .A2(EBX_REG_31__SCAN_IN), .A3(n5346), .ZN(n5348) );
  NAND2_X1 U6518 ( .A1(n5349), .A2(n5348), .ZN(n5350) );
  INV_X1 U6519 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6691) );
  NAND4_X1 U6520 ( .A1(n5392), .A2(REIP_REG_30__SCAN_IN), .A3(
        REIP_REG_29__SCAN_IN), .A4(n6691), .ZN(n5354) );
  OAI211_X1 U6521 ( .C1(n5356), .C2(n5971), .A(n5355), .B(n5354), .ZN(U2796)
         );
  OAI22_X1 U6522 ( .A1(n5358), .A2(n5522), .B1(n5836), .B2(n5357), .ZN(U2828)
         );
  NAND2_X1 U6523 ( .A1(n5360), .A2(n5359), .ZN(n5542) );
  INV_X1 U6524 ( .A(n5542), .ZN(n5361) );
  NAND2_X1 U6525 ( .A1(n5361), .A2(n5669), .ZN(n5363) );
  NAND2_X1 U6526 ( .A1(n5541), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6527 ( .A1(n5363), .A2(n5362), .ZN(n5364) );
  XNOR2_X1 U6528 ( .A(n5364), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5663)
         );
  NOR2_X1 U6529 ( .A1(n5374), .A2(n6175), .ZN(n5372) );
  INV_X1 U6530 ( .A(n5384), .ZN(n5370) );
  NAND2_X1 U6531 ( .A1(n6215), .A2(REIP_REG_30__SCAN_IN), .ZN(n5656) );
  OAI21_X1 U6532 ( .B1(n6171), .B2(n5367), .A(n5656), .ZN(n5368) );
  INV_X1 U6533 ( .A(n5368), .ZN(n5369) );
  OAI21_X1 U6534 ( .B1(n5663), .B2(n5914), .A(n5373), .ZN(U2956) );
  AOI22_X1 U6535 ( .A1(n6042), .A2(DATAI_30_), .B1(n6045), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5378) );
  AND2_X1 U6536 ( .A1(n3227), .A2(n3219), .ZN(n5376) );
  NAND2_X1 U6537 ( .A1(n6046), .A2(DATAI_14_), .ZN(n5377) );
  OAI211_X1 U6538 ( .C1(n5374), .C2(n5837), .A(n5378), .B(n5377), .ZN(U2861)
         );
  MUX2_X1 U6539 ( .A(n4275), .B(n5379), .S(n5484), .Z(n5381) );
  XNOR2_X1 U6540 ( .A(n5381), .B(n5380), .ZN(n5658) );
  INV_X1 U6541 ( .A(n5658), .ZN(n5390) );
  INV_X1 U6542 ( .A(n5382), .ZN(n5383) );
  AOI22_X1 U6543 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n5978), .B1(n5993), 
        .B2(n5384), .ZN(n5386) );
  NAND2_X1 U6544 ( .A1(n6018), .A2(EBX_REG_30__SCAN_IN), .ZN(n5385) );
  INV_X1 U6545 ( .A(REIP_REG_30__SCAN_IN), .ZN(n5391) );
  NAND3_X1 U6546 ( .A1(n5392), .A2(REIP_REG_29__SCAN_IN), .A3(n5391), .ZN(
        n5393) );
  OAI211_X1 U6547 ( .C1(n5374), .C2(n5971), .A(n5394), .B(n5393), .ZN(U2797)
         );
  INV_X1 U6548 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5395) );
  OAI222_X1 U6549 ( .A1(n5524), .A2(n5374), .B1(n5395), .B2(n5836), .C1(n5522), 
        .C2(n5658), .ZN(U2829) );
  NAND2_X1 U6550 ( .A1(n5396), .A2(n3545), .ZN(n5411) );
  INV_X1 U6551 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6673) );
  NAND2_X1 U6552 ( .A1(n5397), .A2(n6673), .ZN(n5398) );
  MUX2_X1 U6553 ( .A(n5411), .B(n5398), .S(n6585), .Z(U3474) );
  NAND2_X1 U6554 ( .A1(n5400), .A2(n5399), .ZN(n5409) );
  NAND3_X1 U6555 ( .A1(n5403), .A2(n5402), .A3(n5401), .ZN(n5406) );
  AOI22_X1 U6556 ( .A1(n5407), .A2(n5406), .B1(n5405), .B2(n5404), .ZN(n5408)
         );
  NAND2_X1 U6557 ( .A1(n5409), .A2(n5408), .ZN(n6471) );
  NOR2_X1 U6558 ( .A1(n5411), .A2(n5410), .ZN(n6582) );
  OAI21_X1 U6559 ( .B1(READY_N), .B2(n6582), .A(n5412), .ZN(n6469) );
  AND2_X1 U6560 ( .A1(n6469), .A2(n6491), .ZN(n5915) );
  MUX2_X1 U6561 ( .A(MORE_REG_SCAN_IN), .B(n6471), .S(n5915), .Z(U3471) );
  AOI21_X1 U6562 ( .B1(n5415), .B2(n5414), .A(n4308), .ZN(n5583) );
  INV_X1 U6563 ( .A(n5583), .ZN(n5538) );
  NOR2_X1 U6564 ( .A1(n5430), .A2(n5416), .ZN(n5417) );
  OR2_X1 U6565 ( .A1(n5418), .A2(n5417), .ZN(n5498) );
  INV_X1 U6566 ( .A(n5498), .ZN(n5703) );
  INV_X1 U6567 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5419) );
  OAI22_X1 U6568 ( .A1(n5419), .A2(n6023), .B1(n6022), .B2(n5581), .ZN(n5420)
         );
  AOI21_X1 U6569 ( .B1(n6020), .B2(n5703), .A(n5420), .ZN(n5421) );
  OAI21_X1 U6570 ( .B1(n5422), .B2(n5954), .A(n5421), .ZN(n5424) );
  AOI211_X1 U6571 ( .C1(n5436), .C2(REIP_REG_24__SCAN_IN), .A(n5424), .B(n5423), .ZN(n5425) );
  OAI21_X1 U6572 ( .B1(n5538), .B2(n5971), .A(n5425), .ZN(U2803) );
  NAND2_X1 U6573 ( .A1(n5426), .A2(n5427), .ZN(n5428) );
  NAND2_X1 U6574 ( .A1(n5414), .A2(n5428), .ZN(n5591) );
  INV_X1 U6575 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6552) );
  NAND2_X1 U6576 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5442), .ZN(n5812) );
  INV_X1 U6577 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6718) );
  OAI21_X1 U6578 ( .B1(n6552), .B2(n5812), .A(n6718), .ZN(n5437) );
  INV_X1 U6579 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5429) );
  OAI22_X1 U6580 ( .A1(n5429), .A2(n6023), .B1(n5593), .B2(n6022), .ZN(n5435)
         );
  INV_X1 U6581 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5433) );
  AOI21_X1 U6582 ( .B1(n5431), .B2(n5504), .A(n5430), .ZN(n5709) );
  INV_X1 U6583 ( .A(n5709), .ZN(n5432) );
  OAI22_X1 U6584 ( .A1(n5954), .A2(n5433), .B1(n5432), .B2(n6009), .ZN(n5434)
         );
  AOI211_X1 U6585 ( .C1(n5437), .C2(n5436), .A(n5435), .B(n5434), .ZN(n5438)
         );
  OAI21_X1 U6586 ( .B1(n5591), .B2(n5971), .A(n5438), .ZN(U2804) );
  OAI21_X1 U6587 ( .B1(n5439), .B2(n5441), .A(n5440), .ZN(n5507) );
  INV_X1 U6588 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6734) );
  NAND2_X1 U6589 ( .A1(n5442), .A2(n6734), .ZN(n5818) );
  NAND2_X1 U6590 ( .A1(n5962), .A2(n5443), .ZN(n5819) );
  XNOR2_X1 U6591 ( .A(n5445), .B(n5444), .ZN(n5726) );
  INV_X1 U6592 ( .A(n5726), .ZN(n5448) );
  INV_X1 U6593 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5446) );
  OAI22_X1 U6594 ( .A1(n5446), .A2(n6023), .B1(n6022), .B2(n5608), .ZN(n5447)
         );
  AOI21_X1 U6595 ( .B1(n6020), .B2(n5448), .A(n5447), .ZN(n5450) );
  NAND2_X1 U6596 ( .A1(n6018), .A2(EBX_REG_21__SCAN_IN), .ZN(n5449) );
  OAI211_X1 U6597 ( .C1(n5819), .C2(n6734), .A(n5450), .B(n5449), .ZN(n5451)
         );
  INV_X1 U6598 ( .A(n5451), .ZN(n5452) );
  OAI211_X1 U6599 ( .C1(n5507), .C2(n5971), .A(n5818), .B(n5452), .ZN(U2806)
         );
  NOR2_X1 U6600 ( .A1(n5453), .A2(n5454), .ZN(n5455) );
  OR2_X1 U6601 ( .A1(n5439), .A2(n5455), .ZN(n5852) );
  MUX2_X1 U6602 ( .A(n4275), .B(n5473), .S(n5456), .Z(n5458) );
  XNOR2_X1 U6603 ( .A(n5458), .B(n5457), .ZN(n5748) );
  INV_X1 U6604 ( .A(n5748), .ZN(n5463) );
  INV_X1 U6605 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5613) );
  AOI22_X1 U6606 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6018), .B1(n5616), .B2(n5993), .ZN(n5459) );
  OAI21_X1 U6607 ( .B1(n6023), .B2(n5613), .A(n5459), .ZN(n5462) );
  AOI21_X1 U6608 ( .B1(n6756), .B2(n5460), .A(n5819), .ZN(n5461) );
  AOI211_X1 U6609 ( .C1(n5463), .C2(n6020), .A(n5462), .B(n5461), .ZN(n5464)
         );
  OAI21_X1 U6610 ( .B1(n5852), .B2(n5971), .A(n5464), .ZN(U2807) );
  INV_X1 U6611 ( .A(n5466), .ZN(n5467) );
  AOI21_X1 U6612 ( .B1(n5468), .B2(n5279), .A(n5467), .ZN(n6036) );
  INV_X1 U6613 ( .A(n6036), .ZN(n5525) );
  INV_X1 U6614 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6547) );
  AOI22_X1 U6615 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6018), .B1(n5821), .B2(n6547), .ZN(n5469) );
  OAI211_X1 U6616 ( .C1(n6023), .C2(n5624), .A(n5469), .B(n5967), .ZN(n5470)
         );
  AOI21_X1 U6617 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5825), .A(n5470), .ZN(n5475) );
  MUX2_X1 U6618 ( .A(n5473), .B(n5472), .S(n5471), .Z(n5519) );
  XNOR2_X1 U6619 ( .A(n5519), .B(n5514), .ZN(n5767) );
  AOI22_X1 U6620 ( .A1(n6020), .A2(n5767), .B1(n5993), .B2(n5626), .ZN(n5474)
         );
  OAI211_X1 U6621 ( .C1(n5525), .C2(n5971), .A(n5475), .B(n5474), .ZN(U2809)
         );
  OAI222_X1 U6622 ( .A1(n5524), .A2(n5533), .B1(n5477), .B2(n5836), .C1(n5476), 
        .C2(n5522), .ZN(U2830) );
  NAND2_X1 U6623 ( .A1(n5478), .A2(n5479), .ZN(n5480) );
  NOR2_X1 U6624 ( .A1(n5685), .A2(n5482), .ZN(n5483) );
  OR2_X1 U6625 ( .A1(n5484), .A2(n5483), .ZN(n5787) );
  OAI22_X1 U6626 ( .A1(n5787), .A2(n5522), .B1(n5485), .B2(n5836), .ZN(n5486)
         );
  AOI21_X1 U6627 ( .B1(n5838), .B2(n5833), .A(n5486), .ZN(n5487) );
  INV_X1 U6628 ( .A(n5487), .ZN(U2831) );
  INV_X1 U6629 ( .A(n5488), .ZN(n5489) );
  OAI21_X1 U6630 ( .B1(n5490), .B2(n4309), .A(n5489), .ZN(n5803) );
  INV_X1 U6631 ( .A(n5803), .ZN(n5570) );
  NAND2_X1 U6632 ( .A1(n5492), .A2(n5491), .ZN(n5493) );
  NAND2_X1 U6633 ( .A1(n5683), .A2(n5493), .ZN(n5802) );
  OAI22_X1 U6634 ( .A1(n5522), .A2(n5802), .B1(n5809), .B2(n5836), .ZN(n5494)
         );
  AOI21_X1 U6635 ( .B1(n5570), .B2(n5833), .A(n5494), .ZN(n5495) );
  INV_X1 U6636 ( .A(n5495), .ZN(U2833) );
  INV_X1 U6637 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5496) );
  OAI222_X1 U6638 ( .A1(n5497), .A2(n5524), .B1(n5496), .B2(n5836), .C1(n5874), 
        .C2(n5522), .ZN(U2834) );
  OAI222_X1 U6639 ( .A1(n5524), .A2(n5538), .B1(n5836), .B2(n5422), .C1(n5498), 
        .C2(n5522), .ZN(U2835) );
  AOI22_X1 U6640 ( .A1(n5831), .A2(n5709), .B1(EBX_REG_23__SCAN_IN), .B2(n5499), .ZN(n5500) );
  OAI21_X1 U6641 ( .B1(n5591), .B2(n5524), .A(n5500), .ZN(U2836) );
  NAND2_X1 U6642 ( .A1(n5502), .A2(n5501), .ZN(n5503) );
  NAND2_X1 U6643 ( .A1(n5504), .A2(n5503), .ZN(n5813) );
  INV_X1 U6644 ( .A(n5426), .ZN(n5505) );
  AOI21_X1 U6645 ( .B1(n5506), .B2(n5440), .A(n5505), .ZN(n5602) );
  INV_X1 U6646 ( .A(n5602), .ZN(n5814) );
  OAI222_X1 U6647 ( .A1(n5522), .A2(n5813), .B1(n5836), .B2(n4238), .C1(n5814), 
        .C2(n5524), .ZN(U2837) );
  INV_X1 U6648 ( .A(n5507), .ZN(n5849) );
  OAI22_X1 U6649 ( .A1(n5522), .A2(n5726), .B1(n5508), .B2(n5836), .ZN(n5509)
         );
  AOI21_X1 U6650 ( .B1(n5849), .B2(n5833), .A(n5509), .ZN(n5510) );
  INV_X1 U6651 ( .A(n5510), .ZN(U2838) );
  OAI222_X1 U6652 ( .A1(n5852), .A2(n5524), .B1(n5511), .B2(n5836), .C1(n5522), 
        .C2(n5748), .ZN(U2839) );
  AND2_X1 U6653 ( .A1(n5466), .A2(n5512), .ZN(n5513) );
  INV_X1 U6654 ( .A(n5456), .ZN(n5518) );
  INV_X1 U6655 ( .A(n5514), .ZN(n5515) );
  NOR2_X1 U6656 ( .A1(n5515), .A2(n5519), .ZN(n5517) );
  OAI22_X1 U6657 ( .A1(n5519), .A2(n5518), .B1(n5517), .B2(n5516), .ZN(n5826)
         );
  OAI22_X1 U6658 ( .A1(n5522), .A2(n5826), .B1(n5830), .B2(n5836), .ZN(n5520)
         );
  AOI21_X1 U6659 ( .B1(n3089), .B2(n5833), .A(n5520), .ZN(n5521) );
  INV_X1 U6660 ( .A(n5521), .ZN(U2840) );
  INV_X1 U6661 ( .A(n5767), .ZN(n5523) );
  OAI222_X1 U6662 ( .A1(n5525), .A2(n5524), .B1(n5836), .B2(n4226), .C1(n5523), 
        .C2(n5522), .ZN(U2841) );
  NAND3_X1 U6663 ( .A1(n5528), .A2(n5527), .A3(n5526), .ZN(n5530) );
  AOI22_X1 U6664 ( .A1(n6042), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6045), .ZN(n5529) );
  NAND2_X1 U6665 ( .A1(n5530), .A2(n5529), .ZN(U2860) );
  AOI22_X1 U6666 ( .A1(n6042), .A2(DATAI_29_), .B1(n6045), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U6667 ( .A1(n6046), .A2(DATAI_13_), .ZN(n5531) );
  OAI211_X1 U6668 ( .C1(n5533), .C2(n5837), .A(n5532), .B(n5531), .ZN(U2862)
         );
  AOI22_X1 U6669 ( .A1(n6046), .A2(DATAI_10_), .B1(n6045), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U6670 ( .A1(n6042), .A2(DATAI_26_), .ZN(n5534) );
  OAI211_X1 U6671 ( .C1(n5803), .C2(n5837), .A(n5535), .B(n5534), .ZN(U2865)
         );
  AOI22_X1 U6672 ( .A1(n6042), .A2(DATAI_24_), .B1(n6045), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U6673 ( .A1(n6046), .A2(DATAI_8_), .ZN(n5536) );
  OAI211_X1 U6674 ( .C1(n5538), .C2(n5837), .A(n5537), .B(n5536), .ZN(U2867)
         );
  AOI22_X1 U6675 ( .A1(n6046), .A2(DATAI_6_), .B1(n6045), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5540) );
  NAND2_X1 U6676 ( .A1(n6042), .A2(DATAI_22_), .ZN(n5539) );
  OAI211_X1 U6677 ( .C1(n5814), .C2(n5837), .A(n5540), .B(n5539), .ZN(U2869)
         );
  INV_X1 U6678 ( .A(n5541), .ZN(n5543) );
  NAND2_X1 U6679 ( .A1(n5543), .A2(n5542), .ZN(n5544) );
  XNOR2_X1 U6680 ( .A(n5544), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5673)
         );
  AND2_X1 U6681 ( .A1(n6215), .A2(REIP_REG_29__SCAN_IN), .ZN(n5666) );
  AOI21_X1 U6682 ( .B1(n6156), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5666), 
        .ZN(n5545) );
  OAI21_X1 U6683 ( .B1(n6166), .B2(n5546), .A(n5545), .ZN(n5547) );
  AOI21_X1 U6684 ( .B1(n5548), .B2(n6162), .A(n5547), .ZN(n5549) );
  OAI21_X1 U6685 ( .B1(n5673), .B2(n5914), .A(n5549), .ZN(U2957) );
  NAND3_X1 U6686 ( .A1(n3014), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n2992), .ZN(n5552) );
  NAND2_X1 U6687 ( .A1(n5879), .A2(n5551), .ZN(n5697) );
  NOR2_X1 U6688 ( .A1(n2992), .A2(n5697), .ZN(n5550) );
  NAND2_X1 U6689 ( .A1(n3030), .A2(n5550), .ZN(n5559) );
  AOI22_X1 U6690 ( .A1(n5552), .A2(n5559), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5551), .ZN(n5553) );
  XNOR2_X1 U6691 ( .A(n5553), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5680)
         );
  INV_X1 U6692 ( .A(n5786), .ZN(n5555) );
  AND2_X1 U6693 ( .A1(n6215), .A2(REIP_REG_28__SCAN_IN), .ZN(n5675) );
  AOI21_X1 U6694 ( .B1(n6156), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5675), 
        .ZN(n5554) );
  OAI21_X1 U6695 ( .B1(n6166), .B2(n5555), .A(n5554), .ZN(n5556) );
  AOI21_X1 U6696 ( .B1(n5838), .B2(n6162), .A(n5556), .ZN(n5557) );
  OAI21_X1 U6697 ( .B1(n5914), .B2(n5680), .A(n5557), .ZN(U2958) );
  NAND2_X1 U6698 ( .A1(n5558), .A2(n5559), .ZN(n5560) );
  XNOR2_X1 U6699 ( .A(n5560), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5693)
         );
  OR2_X1 U6700 ( .A1(n5488), .A2(n5561), .ZN(n5562) );
  AND2_X1 U6701 ( .A1(n6215), .A2(REIP_REG_27__SCAN_IN), .ZN(n5686) );
  AOI21_X1 U6702 ( .B1(n6156), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5686), 
        .ZN(n5563) );
  OAI21_X1 U6703 ( .B1(n6166), .B2(n5794), .A(n5563), .ZN(n5564) );
  AOI21_X1 U6704 ( .B1(n5841), .B2(n6162), .A(n5564), .ZN(n5565) );
  OAI21_X1 U6705 ( .B1(n5693), .B2(n5914), .A(n5565), .ZN(U2959) );
  XNOR2_X1 U6706 ( .A(n2992), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5566)
         );
  XNOR2_X1 U6707 ( .A(n3014), .B(n5566), .ZN(n5701) );
  INV_X1 U6708 ( .A(n5800), .ZN(n5568) );
  AND2_X1 U6709 ( .A1(n6215), .A2(REIP_REG_26__SCAN_IN), .ZN(n5695) );
  AOI21_X1 U6710 ( .B1(n6156), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5695), 
        .ZN(n5567) );
  OAI21_X1 U6711 ( .B1(n6166), .B2(n5568), .A(n5567), .ZN(n5569) );
  AOI21_X1 U6712 ( .B1(n5570), .B2(n6162), .A(n5569), .ZN(n5571) );
  OAI21_X1 U6713 ( .B1(n5914), .B2(n5701), .A(n5571), .ZN(U2960) );
  NAND2_X1 U6714 ( .A1(n2992), .A2(n5753), .ZN(n5572) );
  XNOR2_X1 U6715 ( .A(n2992), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5612)
         );
  INV_X1 U6716 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5573) );
  INV_X1 U6717 ( .A(n5606), .ZN(n5576) );
  XNOR2_X1 U6718 ( .A(n5621), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5605)
         );
  NOR2_X1 U6719 ( .A1(n2992), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5596)
         );
  NAND2_X1 U6720 ( .A1(n5604), .A2(n5596), .ZN(n5587) );
  NAND3_X1 U6721 ( .A1(n2992), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5578) );
  OAI21_X1 U6722 ( .B1(n5621), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5577), 
        .ZN(n5598) );
  OAI22_X2 U6723 ( .A1(n5587), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5578), .B2(n5598), .ZN(n5579) );
  XNOR2_X1 U6724 ( .A(n5579), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5708)
         );
  NOR2_X1 U6725 ( .A1(n5900), .A2(n6687), .ZN(n5702) );
  AOI21_X1 U6726 ( .B1(n6156), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5702), 
        .ZN(n5580) );
  OAI21_X1 U6727 ( .B1(n6166), .B2(n5581), .A(n5580), .ZN(n5582) );
  AOI21_X1 U6728 ( .B1(n5583), .B2(n6162), .A(n5582), .ZN(n5584) );
  OAI21_X1 U6729 ( .B1(n5708), .B2(n5914), .A(n5584), .ZN(U2962) );
  NAND3_X1 U6730 ( .A1(n2992), .A2(n5720), .A3(n5586), .ZN(n5588) );
  OAI21_X1 U6731 ( .B1(n5589), .B2(n5588), .A(n5587), .ZN(n5590) );
  XNOR2_X1 U6732 ( .A(n5590), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5717)
         );
  INV_X1 U6733 ( .A(n5591), .ZN(n5846) );
  NAND2_X1 U6734 ( .A1(n6215), .A2(REIP_REG_23__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U6735 ( .A1(n6156), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5592)
         );
  OAI211_X1 U6736 ( .C1(n6166), .C2(n5593), .A(n5711), .B(n5592), .ZN(n5594)
         );
  AOI21_X1 U6737 ( .B1(n5846), .B2(n6162), .A(n5594), .ZN(n5595) );
  OAI21_X1 U6738 ( .B1(n5717), .B2(n5914), .A(n5595), .ZN(U2963) );
  AOI21_X1 U6739 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n2992), .A(n5596), 
        .ZN(n5597) );
  XNOR2_X1 U6740 ( .A(n5598), .B(n5597), .ZN(n5724) );
  NAND2_X1 U6741 ( .A1(n5642), .A2(n5810), .ZN(n5599) );
  NAND2_X1 U6742 ( .A1(n6215), .A2(REIP_REG_22__SCAN_IN), .ZN(n5718) );
  OAI211_X1 U6743 ( .C1(n6171), .C2(n5600), .A(n5599), .B(n5718), .ZN(n5601)
         );
  AOI21_X1 U6744 ( .B1(n5602), .B2(n6162), .A(n5601), .ZN(n5603) );
  OAI21_X1 U6745 ( .B1(n5724), .B2(n5914), .A(n5603), .ZN(U2964) );
  AOI21_X1 U6746 ( .B1(n5606), .B2(n5605), .A(n5604), .ZN(n5732) );
  NAND2_X1 U6747 ( .A1(n6215), .A2(REIP_REG_21__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U6748 ( .A1(n6156), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5607)
         );
  OAI211_X1 U6749 ( .C1(n6166), .C2(n5608), .A(n5725), .B(n5607), .ZN(n5609)
         );
  AOI21_X1 U6750 ( .B1(n5849), .B2(n6162), .A(n5609), .ZN(n5610) );
  OAI21_X1 U6751 ( .B1(n5732), .B2(n5914), .A(n5610), .ZN(U2965) );
  XOR2_X1 U6752 ( .A(n5612), .B(n5611), .Z(n5751) );
  NAND2_X1 U6753 ( .A1(n6215), .A2(REIP_REG_20__SCAN_IN), .ZN(n5746) );
  OAI21_X1 U6754 ( .B1(n6171), .B2(n5613), .A(n5746), .ZN(n5615) );
  NOR2_X1 U6755 ( .A1(n5852), .A2(n6175), .ZN(n5614) );
  AOI211_X1 U6756 ( .C1(n5642), .C2(n5616), .A(n5615), .B(n5614), .ZN(n5617)
         );
  OAI21_X1 U6757 ( .B1(n5751), .B2(n5914), .A(n5617), .ZN(U2966) );
  BUF_X1 U6758 ( .A(n5618), .Z(n5619) );
  NAND2_X1 U6759 ( .A1(n2992), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5870) );
  INV_X1 U6760 ( .A(n5620), .ZN(n5622) );
  INV_X1 U6761 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5762) );
  NAND4_X1 U6762 ( .A1(n5622), .A2(n5621), .A3(n5774), .A4(n5762), .ZN(n5868)
         );
  OAI21_X1 U6763 ( .B1(n5619), .B2(n5870), .A(n5868), .ZN(n5623) );
  XNOR2_X1 U6764 ( .A(n5623), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5769)
         );
  OAI22_X1 U6765 ( .A1(n6171), .A2(n5624), .B1(n5900), .B2(n6547), .ZN(n5625)
         );
  AOI21_X1 U6766 ( .B1(n5642), .B2(n5626), .A(n5625), .ZN(n5628) );
  NAND2_X1 U6767 ( .A1(n6036), .A2(n6162), .ZN(n5627) );
  OAI211_X1 U6768 ( .C1(n5769), .C2(n5914), .A(n5628), .B(n5627), .ZN(U2968)
         );
  INV_X1 U6769 ( .A(n5866), .ZN(n5630) );
  NOR2_X1 U6770 ( .A1(n5630), .A2(n5629), .ZN(n5632) );
  XOR2_X1 U6771 ( .A(n5632), .B(n5631), .Z(n5780) );
  AND2_X1 U6772 ( .A1(n6215), .A2(REIP_REG_16__SCAN_IN), .ZN(n5776) );
  AOI21_X1 U6773 ( .B1(n6156), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5776), 
        .ZN(n5633) );
  OAI21_X1 U6774 ( .B1(n6166), .B2(n5634), .A(n5633), .ZN(n5635) );
  AOI21_X1 U6775 ( .B1(n6044), .B2(n6162), .A(n5635), .ZN(n5636) );
  OAI21_X1 U6776 ( .B1(n5780), .B2(n5914), .A(n5636), .ZN(U2970) );
  OAI21_X1 U6777 ( .B1(n5637), .B2(n5638), .A(n5620), .ZN(n5890) );
  NAND2_X1 U6778 ( .A1(n5890), .A2(n6173), .ZN(n5644) );
  OAI22_X1 U6779 ( .A1(n6171), .A2(n3806), .B1(n5900), .B2(n5639), .ZN(n5640)
         );
  AOI21_X1 U6780 ( .B1(n5642), .B2(n5641), .A(n5640), .ZN(n5643) );
  OAI211_X1 U6781 ( .C1(n6175), .C2(n5645), .A(n5644), .B(n5643), .ZN(U2971)
         );
  XNOR2_X1 U6782 ( .A(n2992), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5647)
         );
  XNOR2_X1 U6783 ( .A(n5646), .B(n5647), .ZN(n5903) );
  INV_X1 U6784 ( .A(n5903), .ZN(n5654) );
  INV_X1 U6785 ( .A(n5648), .ZN(n5652) );
  AOI22_X1 U6786 ( .A1(n6156), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6215), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5649) );
  OAI21_X1 U6787 ( .B1(n6166), .B2(n5650), .A(n5649), .ZN(n5651) );
  AOI21_X1 U6788 ( .B1(n5652), .B2(n6162), .A(n5651), .ZN(n5653) );
  OAI21_X1 U6789 ( .B1(n5654), .B2(n5914), .A(n5653), .ZN(U2972) );
  NAND2_X1 U6790 ( .A1(n5655), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5657) );
  OAI211_X1 U6791 ( .C1(n5658), .C2(n6225), .A(n5657), .B(n5656), .ZN(n5659)
         );
  AOI21_X1 U6792 ( .B1(n5661), .B2(n5660), .A(n5659), .ZN(n5662) );
  OAI21_X1 U6793 ( .B1(n5663), .B2(n5779), .A(n5662), .ZN(U2988) );
  INV_X1 U6794 ( .A(n5476), .ZN(n5667) );
  NOR2_X1 U6795 ( .A1(n5664), .A2(n5669), .ZN(n5665) );
  AOI211_X1 U6796 ( .C1(n6210), .C2(n5667), .A(n5666), .B(n5665), .ZN(n5672)
         );
  INV_X1 U6797 ( .A(n5668), .ZN(n5691) );
  NAND3_X1 U6798 ( .A1(n5691), .A2(n5670), .A3(n5669), .ZN(n5671) );
  OAI211_X1 U6799 ( .C1(n5673), .C2(n5779), .A(n5672), .B(n5671), .ZN(U2989)
         );
  NOR2_X1 U6800 ( .A1(n5787), .A2(n6225), .ZN(n5674) );
  AOI211_X1 U6801 ( .C1(n5681), .C2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n5675), .B(n5674), .ZN(n5679) );
  NAND3_X1 U6802 ( .A1(n5691), .A2(n5677), .A3(n5676), .ZN(n5678) );
  OAI211_X1 U6803 ( .C1(n5680), .C2(n5779), .A(n5679), .B(n5678), .ZN(U2990)
         );
  INV_X1 U6804 ( .A(n5681), .ZN(n5688) );
  AND2_X1 U6805 ( .A1(n5683), .A2(n5682), .ZN(n5684) );
  NOR2_X1 U6806 ( .A1(n5685), .A2(n5684), .ZN(n5832) );
  AOI21_X1 U6807 ( .B1(n5832), .B2(n6210), .A(n5686), .ZN(n5687) );
  OAI21_X1 U6808 ( .B1(n5688), .B2(n5690), .A(n5687), .ZN(n5689) );
  AOI21_X1 U6809 ( .B1(n5691), .B2(n5690), .A(n5689), .ZN(n5692) );
  OAI21_X1 U6810 ( .B1(n5693), .B2(n5779), .A(n5692), .ZN(U2991) );
  NOR2_X1 U6811 ( .A1(n5802), .A2(n6225), .ZN(n5694) );
  AOI211_X1 U6812 ( .C1(n5878), .C2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5695), .B(n5694), .ZN(n5700) );
  INV_X1 U6813 ( .A(n5696), .ZN(n5698) );
  NAND3_X1 U6814 ( .A1(n5880), .A2(n5698), .A3(n5697), .ZN(n5699) );
  OAI211_X1 U6815 ( .C1(n5701), .C2(n5779), .A(n5700), .B(n5699), .ZN(U2992)
         );
  AOI21_X1 U6816 ( .B1(n6210), .B2(n5703), .A(n5702), .ZN(n5707) );
  INV_X1 U6817 ( .A(n5704), .ZN(n5705) );
  OAI211_X1 U6818 ( .C1(n5715), .C2(INSTADDRPOINTER_REG_24__SCAN_IN), .A(n5878), .B(n5705), .ZN(n5706) );
  OAI211_X1 U6819 ( .C1(n5708), .C2(n5779), .A(n5707), .B(n5706), .ZN(U2994)
         );
  INV_X1 U6820 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5714) );
  NAND2_X1 U6821 ( .A1(n6210), .A2(n5709), .ZN(n5710) );
  OAI211_X1 U6822 ( .C1(n5712), .C2(n5714), .A(n5711), .B(n5710), .ZN(n5713)
         );
  AOI21_X1 U6823 ( .B1(n5715), .B2(n5714), .A(n5713), .ZN(n5716) );
  OAI21_X1 U6824 ( .B1(n5717), .B2(n5779), .A(n5716), .ZN(U2995) );
  OAI21_X1 U6825 ( .B1(n6225), .B2(n5813), .A(n5718), .ZN(n5722) );
  NOR3_X1 U6826 ( .A1(n5727), .A2(n5720), .A3(n5719), .ZN(n5721) );
  AOI211_X1 U6827 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5730), .A(n5722), .B(n5721), .ZN(n5723) );
  OAI21_X1 U6828 ( .B1(n5724), .B2(n5779), .A(n5723), .ZN(U2996) );
  OAI21_X1 U6829 ( .B1(n6225), .B2(n5726), .A(n5725), .ZN(n5729) );
  NOR2_X1 U6830 ( .A1(n5727), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5728)
         );
  AOI211_X1 U6831 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5730), .A(n5729), .B(n5728), .ZN(n5731) );
  OAI21_X1 U6832 ( .B1(n5732), .B2(n5779), .A(n5731), .ZN(U2997) );
  AOI221_X1 U6833 ( .B1(n5736), .B2(n5735), .C1(n5734), .C2(n5735), .A(n5733), 
        .ZN(n5737) );
  OAI221_X1 U6834 ( .B1(n5739), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .C1(
        n5739), .C2(n5738), .A(n5737), .ZN(n5883) );
  AOI21_X1 U6835 ( .B1(n6217), .B2(n5762), .A(n5883), .ZN(n5764) );
  OAI21_X1 U6836 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5740), .A(n5764), 
        .ZN(n5759) );
  INV_X1 U6837 ( .A(n5888), .ZN(n5745) );
  NAND2_X1 U6838 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5743) );
  INV_X1 U6839 ( .A(n5741), .ZN(n5742) );
  NAND4_X1 U6840 ( .A1(n5745), .A2(n5744), .A3(n5743), .A4(n5742), .ZN(n5747)
         );
  OAI211_X1 U6841 ( .C1(n6225), .C2(n5748), .A(n5747), .B(n5746), .ZN(n5749)
         );
  AOI21_X1 U6842 ( .B1(INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n5759), .A(n5749), 
        .ZN(n5750) );
  OAI21_X1 U6843 ( .B1(n5751), .B2(n5779), .A(n5750), .ZN(U2998) );
  XNOR2_X1 U6844 ( .A(n2992), .B(n5753), .ZN(n5754) );
  XNOR2_X1 U6845 ( .A(n5752), .B(n5754), .ZN(n5862) );
  INV_X1 U6846 ( .A(n5862), .ZN(n5761) );
  INV_X1 U6847 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5755) );
  OAI22_X1 U6848 ( .A1(n6225), .A2(n5826), .B1(n5900), .B2(n5755), .ZN(n5758)
         );
  NOR3_X1 U6849 ( .A1(n5888), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .A3(n5756), 
        .ZN(n5757) );
  AOI211_X1 U6850 ( .C1(n5759), .C2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5758), .B(n5757), .ZN(n5760) );
  OAI21_X1 U6851 ( .B1(n5761), .B2(n5779), .A(n5760), .ZN(U2999) );
  NOR3_X1 U6852 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5762), .A3(n5888), 
        .ZN(n5766) );
  INV_X1 U6853 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5763) );
  OAI22_X1 U6854 ( .A1(n5764), .A2(n5763), .B1(n5900), .B2(n6547), .ZN(n5765)
         );
  AOI211_X1 U6855 ( .C1(n6210), .C2(n5767), .A(n5766), .B(n5765), .ZN(n5768)
         );
  OAI21_X1 U6856 ( .B1(n5769), .B2(n5779), .A(n5768), .ZN(U3000) );
  AOI21_X1 U6857 ( .B1(n5771), .B2(n5770), .A(n6182), .ZN(n5892) );
  NAND3_X1 U6858 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5895), .A3(n6177), .ZN(n5894) );
  OAI21_X1 U6859 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5772), .ZN(n5773) );
  OAI22_X1 U6860 ( .A1(n5892), .A2(n5774), .B1(n5894), .B2(n5773), .ZN(n5775)
         );
  AOI211_X1 U6861 ( .C1(n6210), .C2(n5777), .A(n5776), .B(n5775), .ZN(n5778)
         );
  OAI21_X1 U6862 ( .B1(n5780), .B2(n5779), .A(n5778), .ZN(U3002) );
  OAI211_X1 U6863 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n3029), .A(n6235), .B(
        n6328), .ZN(n5781) );
  OAI21_X1 U6864 ( .B1(n5783), .B2(n5782), .A(n5781), .ZN(n5784) );
  MUX2_X1 U6865 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5784), .S(n6233), 
        .Z(U3464) );
  AND2_X1 U6866 ( .A1(n6062), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U6867 ( .A1(EBX_REG_28__SCAN_IN), .A2(n6018), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n5978), .ZN(n5792) );
  AOI22_X1 U6868 ( .A1(n5786), .A2(n5993), .B1(REIP_REG_28__SCAN_IN), .B2(
        n5785), .ZN(n5791) );
  NOR2_X1 U6869 ( .A1(n6009), .A2(n5787), .ZN(n5788) );
  AOI21_X1 U6870 ( .B1(n5838), .B2(n5982), .A(n5788), .ZN(n5790) );
  INV_X1 U6871 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6626) );
  NAND3_X1 U6872 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5797), .A3(n6626), .ZN(
        n5789) );
  NAND4_X1 U6873 ( .A1(n5792), .A2(n5791), .A3(n5790), .A4(n5789), .ZN(U2799)
         );
  INV_X1 U6874 ( .A(REIP_REG_27__SCAN_IN), .ZN(n5796) );
  AOI22_X1 U6875 ( .A1(EBX_REG_27__SCAN_IN), .A2(n6018), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n5978), .ZN(n5793) );
  OAI21_X1 U6876 ( .B1(n5794), .B2(n6022), .A(n5793), .ZN(n5795) );
  AOI221_X1 U6877 ( .B1(n5806), .B2(REIP_REG_27__SCAN_IN), .C1(n5797), .C2(
        n5796), .A(n5795), .ZN(n5799) );
  AOI22_X1 U6878 ( .A1(n5841), .A2(n5982), .B1(n5832), .B2(n6020), .ZN(n5798)
         );
  NAND2_X1 U6879 ( .A1(n5799), .A2(n5798), .ZN(U2800) );
  AOI22_X1 U6880 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n5978), .B1(n5800), 
        .B2(n5993), .ZN(n5808) );
  OAI21_X1 U6881 ( .B1(n6690), .B2(n5801), .A(n6660), .ZN(n5805) );
  OAI22_X1 U6882 ( .A1(n5803), .A2(n5971), .B1(n6009), .B2(n5802), .ZN(n5804)
         );
  AOI21_X1 U6883 ( .B1(n5806), .B2(n5805), .A(n5804), .ZN(n5807) );
  OAI211_X1 U6884 ( .C1(n5809), .C2(n5954), .A(n5808), .B(n5807), .ZN(U2801)
         );
  AOI22_X1 U6885 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n5978), .B1(n5810), 
        .B2(n5993), .ZN(n5811) );
  OAI21_X1 U6886 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5812), .A(n5811), .ZN(n5816) );
  OAI22_X1 U6887 ( .A1(n5814), .A2(n5971), .B1(n5813), .B2(n6009), .ZN(n5815)
         );
  AOI211_X1 U6888 ( .C1(EBX_REG_22__SCAN_IN), .C2(n6018), .A(n5816), .B(n5815), 
        .ZN(n5817) );
  OAI221_X1 U6889 ( .B1(n6552), .B2(n5819), .C1(n6552), .C2(n5818), .A(n5817), 
        .ZN(U2805) );
  INV_X1 U6890 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5823) );
  NAND2_X1 U6891 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5820) );
  OAI211_X1 U6892 ( .C1(REIP_REG_19__SCAN_IN), .C2(REIP_REG_18__SCAN_IN), .A(
        n5821), .B(n5820), .ZN(n5822) );
  OAI211_X1 U6893 ( .C1(n6023), .C2(n5823), .A(n5822), .B(n5967), .ZN(n5824)
         );
  AOI21_X1 U6894 ( .B1(REIP_REG_19__SCAN_IN), .B2(n5825), .A(n5824), .ZN(n5829) );
  OAI22_X1 U6895 ( .A1(n6009), .A2(n5826), .B1(n5865), .B2(n6022), .ZN(n5827)
         );
  AOI21_X1 U6896 ( .B1(n3089), .B2(n5982), .A(n5827), .ZN(n5828) );
  OAI211_X1 U6897 ( .C1(n5830), .C2(n5954), .A(n5829), .B(n5828), .ZN(U2808)
         );
  INV_X1 U6898 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5835) );
  AOI22_X1 U6899 ( .A1(n5841), .A2(n5833), .B1(n5832), .B2(n5831), .ZN(n5834)
         );
  OAI21_X1 U6900 ( .B1(n5836), .B2(n5835), .A(n5834), .ZN(U2832) );
  AOI22_X1 U6901 ( .A1(n5838), .A2(n6043), .B1(n6042), .B2(DATAI_28_), .ZN(
        n5840) );
  AOI22_X1 U6902 ( .A1(n6046), .A2(DATAI_12_), .B1(n6045), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U6903 ( .A1(n5840), .A2(n5839), .ZN(U2863) );
  AOI22_X1 U6904 ( .A1(n5841), .A2(n6043), .B1(n6042), .B2(DATAI_27_), .ZN(
        n5843) );
  AOI22_X1 U6905 ( .A1(n6046), .A2(DATAI_11_), .B1(n6045), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5842) );
  NAND2_X1 U6906 ( .A1(n5843), .A2(n5842), .ZN(U2864) );
  AOI22_X1 U6907 ( .A1(n5858), .A2(n6043), .B1(n6042), .B2(DATAI_25_), .ZN(
        n5845) );
  AOI22_X1 U6908 ( .A1(n6046), .A2(DATAI_9_), .B1(n6045), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5844) );
  NAND2_X1 U6909 ( .A1(n5845), .A2(n5844), .ZN(U2866) );
  AOI22_X1 U6910 ( .A1(n5846), .A2(n6043), .B1(n6042), .B2(DATAI_23_), .ZN(
        n5848) );
  AOI22_X1 U6911 ( .A1(n6046), .A2(DATAI_7_), .B1(n6045), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U6912 ( .A1(n5848), .A2(n5847), .ZN(U2868) );
  AOI22_X1 U6913 ( .A1(n5849), .A2(n6043), .B1(n6042), .B2(DATAI_21_), .ZN(
        n5851) );
  AOI22_X1 U6914 ( .A1(n6046), .A2(DATAI_5_), .B1(n6045), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U6915 ( .A1(n5851), .A2(n5850), .ZN(U2870) );
  INV_X1 U6916 ( .A(n5852), .ZN(n5853) );
  AOI22_X1 U6917 ( .A1(n5853), .A2(n6043), .B1(n6042), .B2(DATAI_20_), .ZN(
        n5855) );
  AOI22_X1 U6918 ( .A1(n6046), .A2(DATAI_4_), .B1(n6045), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U6919 ( .A1(n5855), .A2(n5854), .ZN(U2871) );
  AOI22_X1 U6920 ( .A1(n3089), .A2(n6043), .B1(n6042), .B2(DATAI_19_), .ZN(
        n5857) );
  AOI22_X1 U6921 ( .A1(n6046), .A2(DATAI_3_), .B1(n6045), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5856) );
  NAND2_X1 U6922 ( .A1(n5857), .A2(n5856), .ZN(U2872) );
  AOI22_X1 U6923 ( .A1(n6215), .A2(REIP_REG_25__SCAN_IN), .B1(n6156), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5860) );
  OAI21_X1 U6924 ( .B1(n3033), .B2(n3030), .A(n3535), .ZN(n5876) );
  AOI22_X1 U6925 ( .A1(n5858), .A2(n6162), .B1(n6173), .B2(n5876), .ZN(n5859)
         );
  OAI211_X1 U6926 ( .C1(n6166), .C2(n5861), .A(n5860), .B(n5859), .ZN(U2961)
         );
  AOI22_X1 U6927 ( .A1(n6215), .A2(REIP_REG_19__SCAN_IN), .B1(n6156), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5864) );
  AOI22_X1 U6928 ( .A1(n5862), .A2(n6173), .B1(n3089), .B2(n6162), .ZN(n5863)
         );
  OAI211_X1 U6929 ( .C1(n6166), .C2(n5865), .A(n5864), .B(n5863), .ZN(U2967)
         );
  AOI22_X1 U6930 ( .A1(n6215), .A2(REIP_REG_17__SCAN_IN), .B1(n6156), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5872) );
  NAND2_X1 U6931 ( .A1(n5619), .A2(n5866), .ZN(n5867) );
  OAI211_X1 U6932 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n2992), .A(n5867), .B(n5870), .ZN(n5869) );
  OAI211_X1 U6933 ( .C1(n3526), .C2(n5870), .A(n5869), .B(n5868), .ZN(n5885)
         );
  AOI22_X1 U6934 ( .A1(n5885), .A2(n6173), .B1(n6162), .B2(n6039), .ZN(n5871)
         );
  OAI211_X1 U6935 ( .C1(n6166), .C2(n5873), .A(n5872), .B(n5871), .ZN(U2969)
         );
  INV_X1 U6936 ( .A(n5874), .ZN(n5875) );
  AOI22_X1 U6937 ( .A1(n5876), .A2(n6227), .B1(n6210), .B2(n5875), .ZN(n5882)
         );
  NOR2_X1 U6938 ( .A1(n5900), .A2(n6690), .ZN(n5877) );
  AOI221_X1 U6939 ( .B1(n5880), .B2(n5879), .C1(n5878), .C2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5877), .ZN(n5881) );
  NAND2_X1 U6940 ( .A1(n5882), .A2(n5881), .ZN(U2993) );
  AOI22_X1 U6941 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5883), .B1(n6215), .B2(REIP_REG_17__SCAN_IN), .ZN(n5887) );
  AOI22_X1 U6942 ( .A1(n5885), .A2(n6227), .B1(n6210), .B2(n5884), .ZN(n5886)
         );
  OAI211_X1 U6943 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5888), .A(n5887), .B(n5886), .ZN(U3001) );
  AOI222_X1 U6944 ( .A1(n5890), .A2(n6227), .B1(REIP_REG_15__SCAN_IN), .B2(
        n6215), .C1(n5889), .C2(n6210), .ZN(n5891) );
  OAI221_X1 U6945 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n5894), .C1(
        n5893), .C2(n5892), .A(n5891), .ZN(U3003) );
  NAND2_X1 U6946 ( .A1(n5895), .A2(n6177), .ZN(n5907) );
  AOI21_X1 U6947 ( .B1(n5897), .B2(n5896), .A(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5899) );
  NOR2_X1 U6948 ( .A1(n5899), .A2(n5898), .ZN(n5905) );
  OAI22_X1 U6949 ( .A1(n6225), .A2(n5901), .B1(n6540), .B2(n5900), .ZN(n5902)
         );
  AOI21_X1 U6950 ( .B1(n5903), .B2(n6227), .A(n5902), .ZN(n5904) );
  OAI221_X1 U6951 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n5907), .C1(
        n5906), .C2(n5905), .A(n5904), .ZN(U3004) );
  NAND3_X1 U6952 ( .A1(n5909), .A2(n6573), .A3(n5908), .ZN(n5910) );
  OAI21_X1 U6953 ( .B1(n5911), .B2(n3640), .A(n5910), .ZN(U3455) );
  INV_X1 U6954 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6716) );
  INV_X1 U6955 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6519) );
  INV_X2 U6956 ( .A(n6789), .ZN(n6788) );
  OAI221_X1 U6957 ( .B1(n6519), .B2(n4126), .C1(STATE_REG_1__SCAN_IN), .C2(
        n4126), .A(n6788), .ZN(n6502) );
  INV_X1 U6958 ( .A(n6502), .ZN(n6568) );
  OAI21_X1 U6959 ( .B1(n6716), .B2(n4126), .A(n6503), .ZN(U2789) );
  INV_X1 U6960 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6704) );
  NOR2_X1 U6961 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5913) );
  NOR2_X1 U6962 ( .A1(n6789), .A2(n5913), .ZN(n5912) );
  AOI22_X1 U6963 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n6789), .B1(n6704), .B2(
        n5912), .ZN(U2791) );
  OAI21_X1 U6964 ( .B1(BS16_N), .B2(n5913), .A(n6568), .ZN(n6566) );
  OAI21_X1 U6965 ( .B1(n6568), .B2(n6656), .A(n6566), .ZN(U2792) );
  OAI21_X1 U6966 ( .B1(n5915), .B2(n6674), .A(n5914), .ZN(U2793) );
  NOR4_X1 U6967 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n5919) );
  NOR4_X1 U6968 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n5918) );
  NOR4_X1 U6969 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5917) );
  NOR4_X1 U6970 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5916) );
  NAND4_X1 U6971 ( .A1(n5919), .A2(n5918), .A3(n5917), .A4(n5916), .ZN(n5925)
         );
  NOR4_X1 U6972 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n5923) );
  AOI211_X1 U6973 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_2__SCAN_IN), .B(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n5922) );
  NOR4_X1 U6974 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n5921) );
  NOR4_X1 U6975 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n5920) );
  NAND4_X1 U6976 ( .A1(n5923), .A2(n5922), .A3(n5921), .A4(n5920), .ZN(n5924)
         );
  NOR2_X1 U6977 ( .A1(n5925), .A2(n5924), .ZN(n6578) );
  INV_X1 U6978 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6706) );
  NOR3_X1 U6979 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5927) );
  OAI21_X1 U6980 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5927), .A(n6578), .ZN(n5926)
         );
  OAI21_X1 U6981 ( .B1(n6578), .B2(n6706), .A(n5926), .ZN(U2794) );
  INV_X1 U6982 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6567) );
  AOI21_X1 U6983 ( .B1(n5085), .B2(n6567), .A(n5927), .ZN(n5928) );
  INV_X1 U6984 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6670) );
  INV_X1 U6985 ( .A(n6578), .ZN(n6575) );
  AOI22_X1 U6986 ( .A1(n6578), .A2(n5928), .B1(n6670), .B2(n6575), .ZN(U2795)
         );
  OAI22_X1 U6987 ( .A1(n5954), .A2(n5930), .B1(n6009), .B2(n5929), .ZN(n5931)
         );
  AOI211_X1 U6988 ( .C1(n5978), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6002), 
        .B(n5931), .ZN(n5941) );
  INV_X1 U6989 ( .A(n5932), .ZN(n5933) );
  AOI22_X1 U6990 ( .A1(n5934), .A2(n5982), .B1(n5993), .B2(n5933), .ZN(n5940)
         );
  NOR3_X1 U6991 ( .A1(n5965), .A2(REIP_REG_12__SCAN_IN), .A3(n5935), .ZN(n5945) );
  OAI21_X1 U6992 ( .B1(n5945), .B2(n5936), .A(REIP_REG_13__SCAN_IN), .ZN(n5939) );
  NAND3_X1 U6993 ( .A1(n6005), .A2(n5299), .A3(n5937), .ZN(n5938) );
  NAND4_X1 U6994 ( .A1(n5941), .A2(n5940), .A3(n5939), .A4(n5938), .ZN(U2814)
         );
  AOI22_X1 U6995 ( .A1(n6020), .A2(n5942), .B1(PHYADDRPOINTER_REG_12__SCAN_IN), 
        .B2(n5978), .ZN(n5950) );
  NOR2_X1 U6996 ( .A1(n5943), .A2(n6538), .ZN(n5944) );
  AOI211_X1 U6997 ( .C1(n6018), .C2(EBX_REG_12__SCAN_IN), .A(n5945), .B(n5944), 
        .ZN(n5949) );
  AOI22_X1 U6998 ( .A1(n5947), .A2(n5982), .B1(n5946), .B2(n5993), .ZN(n5948)
         );
  NAND4_X1 U6999 ( .A1(n5950), .A2(n5949), .A3(n5948), .A4(n5967), .ZN(U2815)
         );
  AND2_X1 U7000 ( .A1(n6005), .A2(n5951), .ZN(n5966) );
  AOI21_X1 U7001 ( .B1(REIP_REG_7__SCAN_IN), .B2(n5966), .A(
        REIP_REG_8__SCAN_IN), .ZN(n5961) );
  OAI22_X1 U7002 ( .A1(n5954), .A2(n5953), .B1(n6009), .B2(n5952), .ZN(n5955)
         );
  AOI211_X1 U7003 ( .C1(n5978), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6002), 
        .B(n5955), .ZN(n5959) );
  AOI22_X1 U7004 ( .A1(n5957), .A2(n5982), .B1(n5993), .B2(n5956), .ZN(n5958)
         );
  OAI211_X1 U7005 ( .C1(n5961), .C2(n5960), .A(n5959), .B(n5958), .ZN(U2819)
         );
  OAI21_X1 U7006 ( .B1(n5963), .B2(n5964), .A(n5962), .ZN(n5997) );
  OR3_X1 U7007 ( .A1(n5965), .A2(REIP_REG_6__SCAN_IN), .A3(n5964), .ZN(n5976)
         );
  INV_X1 U7008 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5969) );
  AOI22_X1 U7009 ( .A1(n5966), .A2(n6530), .B1(n6020), .B2(n6197), .ZN(n5968)
         );
  OAI211_X1 U7010 ( .C1(n6023), .C2(n5969), .A(n5968), .B(n5967), .ZN(n5974)
         );
  OAI22_X1 U7011 ( .A1(n5972), .A2(n5971), .B1(n5970), .B2(n6022), .ZN(n5973)
         );
  AOI211_X1 U7012 ( .C1(EBX_REG_7__SCAN_IN), .C2(n6018), .A(n5974), .B(n5973), 
        .ZN(n5975) );
  OAI221_X1 U7013 ( .B1(n6530), .B2(n5997), .C1(n6530), .C2(n5976), .A(n5975), 
        .ZN(U2820) );
  OAI21_X1 U7014 ( .B1(n5997), .B2(n6528), .A(n5976), .ZN(n5977) );
  AOI21_X1 U7015 ( .B1(EBX_REG_6__SCAN_IN), .B2(n6018), .A(n5977), .ZN(n5985)
         );
  AOI21_X1 U7016 ( .B1(n5978), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6002), 
        .ZN(n5979) );
  OAI21_X1 U7017 ( .B1(n6009), .B2(n5980), .A(n5979), .ZN(n5981) );
  AOI21_X1 U7018 ( .B1(n5983), .B2(n5982), .A(n5981), .ZN(n5984) );
  OAI211_X1 U7019 ( .C1(n5986), .C2(n6022), .A(n5985), .B(n5984), .ZN(U2821)
         );
  AOI21_X1 U7020 ( .B1(n6005), .B2(n5987), .A(REIP_REG_5__SCAN_IN), .ZN(n5998)
         );
  INV_X1 U7021 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5988) );
  OAI22_X1 U7022 ( .A1(n6009), .A2(n5989), .B1(n5988), .B2(n6023), .ZN(n5990)
         );
  AOI211_X1 U7023 ( .C1(n6018), .C2(EBX_REG_5__SCAN_IN), .A(n6002), .B(n5990), 
        .ZN(n5996) );
  INV_X1 U7024 ( .A(n5991), .ZN(n5994) );
  AOI22_X1 U7025 ( .A1(n5994), .A2(n6030), .B1(n5993), .B2(n5992), .ZN(n5995)
         );
  OAI211_X1 U7026 ( .C1(n5998), .C2(n5997), .A(n5996), .B(n5995), .ZN(U2822)
         );
  NAND2_X1 U7027 ( .A1(n6005), .A2(n6003), .ZN(n6035) );
  AND2_X1 U7028 ( .A1(n6035), .A2(n5999), .ZN(n6028) );
  OAI22_X1 U7029 ( .A1(n6028), .A2(n6525), .B1(n6000), .B2(n6023), .ZN(n6001)
         );
  AOI211_X1 U7030 ( .C1(n6018), .C2(EBX_REG_4__SCAN_IN), .A(n6002), .B(n6001), 
        .ZN(n6014) );
  NOR2_X1 U7031 ( .A1(n6003), .A2(REIP_REG_4__SCAN_IN), .ZN(n6004) );
  NAND2_X1 U7032 ( .A1(n6005), .A2(n6004), .ZN(n6008) );
  NAND2_X1 U7033 ( .A1(n6026), .A2(n6006), .ZN(n6007) );
  OAI211_X1 U7034 ( .C1(n6010), .C2(n6009), .A(n6008), .B(n6007), .ZN(n6011)
         );
  AOI21_X1 U7035 ( .B1(n6012), .B2(n6030), .A(n6011), .ZN(n6013) );
  OAI211_X1 U7036 ( .C1(n6015), .C2(n6022), .A(n6014), .B(n6013), .ZN(U2823)
         );
  OR2_X1 U7037 ( .A1(n6017), .A2(n6016), .ZN(n6034) );
  AOI22_X1 U7038 ( .A1(n6020), .A2(n6019), .B1(n6018), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n6033) );
  INV_X1 U7039 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6523) );
  INV_X1 U7040 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6024) );
  OAI22_X1 U7041 ( .A1(n6024), .A2(n6023), .B1(n6022), .B2(n6021), .ZN(n6025)
         );
  AOI21_X1 U7042 ( .B1(n6026), .B2(n6277), .A(n6025), .ZN(n6027) );
  OAI21_X1 U7043 ( .B1(n6028), .B2(n6523), .A(n6027), .ZN(n6029) );
  AOI21_X1 U7044 ( .B1(n6031), .B2(n6030), .A(n6029), .ZN(n6032) );
  OAI211_X1 U7045 ( .C1(n6035), .C2(n6034), .A(n6033), .B(n6032), .ZN(U2824)
         );
  AOI22_X1 U7046 ( .A1(n6036), .A2(n6043), .B1(n6042), .B2(DATAI_18_), .ZN(
        n6038) );
  AOI22_X1 U7047 ( .A1(n6046), .A2(DATAI_2_), .B1(n6045), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U7048 ( .A1(n6038), .A2(n6037), .ZN(U2873) );
  AOI22_X1 U7049 ( .A1(n6039), .A2(n6043), .B1(n6042), .B2(DATAI_17_), .ZN(
        n6041) );
  AOI22_X1 U7050 ( .A1(n6046), .A2(DATAI_1_), .B1(n6045), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7051 ( .A1(n6041), .A2(n6040), .ZN(U2874) );
  AOI22_X1 U7052 ( .A1(n6044), .A2(n6043), .B1(n6042), .B2(DATAI_16_), .ZN(
        n6048) );
  AOI22_X1 U7053 ( .A1(n6046), .A2(DATAI_0_), .B1(n6045), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6047) );
  NAND2_X1 U7054 ( .A1(n6048), .A2(n6047), .ZN(U2875) );
  INV_X1 U7055 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6155) );
  AOI22_X1 U7056 ( .A1(n6067), .A2(LWORD_REG_15__SCAN_IN), .B1(n6062), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6050) );
  OAI21_X1 U7057 ( .B1(n6155), .B2(n6069), .A(n6050), .ZN(U2908) );
  INV_X1 U7058 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6150) );
  AOI22_X1 U7059 ( .A1(n6067), .A2(LWORD_REG_14__SCAN_IN), .B1(n6062), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6051) );
  OAI21_X1 U7060 ( .B1(n6150), .B2(n6069), .A(n6051), .ZN(U2909) );
  AOI22_X1 U7061 ( .A1(n6067), .A2(LWORD_REG_13__SCAN_IN), .B1(n6062), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6052) );
  OAI21_X1 U7062 ( .B1(n6147), .B2(n6069), .A(n6052), .ZN(U2910) );
  AOI22_X1 U7063 ( .A1(n6067), .A2(LWORD_REG_12__SCAN_IN), .B1(n6062), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6053) );
  OAI21_X1 U7064 ( .B1(n3737), .B2(n6069), .A(n6053), .ZN(U2911) );
  AOI22_X1 U7065 ( .A1(n6067), .A2(LWORD_REG_11__SCAN_IN), .B1(n6066), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6054) );
  OAI21_X1 U7066 ( .B1(n6142), .B2(n6069), .A(n6054), .ZN(U2912) );
  AOI22_X1 U7067 ( .A1(n6067), .A2(LWORD_REG_10__SCAN_IN), .B1(n6062), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6055) );
  OAI21_X1 U7068 ( .B1(n6139), .B2(n6069), .A(n6055), .ZN(U2913) );
  AOI22_X1 U7069 ( .A1(n6067), .A2(LWORD_REG_9__SCAN_IN), .B1(n6062), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6056) );
  OAI21_X1 U7070 ( .B1(n6136), .B2(n6069), .A(n6056), .ZN(U2914) );
  AOI22_X1 U7071 ( .A1(n6067), .A2(LWORD_REG_8__SCAN_IN), .B1(n6062), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6057) );
  OAI21_X1 U7072 ( .B1(n6133), .B2(n6069), .A(n6057), .ZN(U2915) );
  AOI22_X1 U7073 ( .A1(n6067), .A2(LWORD_REG_7__SCAN_IN), .B1(n6062), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6058) );
  OAI21_X1 U7074 ( .B1(n6130), .B2(n6069), .A(n6058), .ZN(U2916) );
  AOI22_X1 U7075 ( .A1(n6067), .A2(LWORD_REG_6__SCAN_IN), .B1(n6062), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6059) );
  OAI21_X1 U7076 ( .B1(n4904), .B2(n6069), .A(n6059), .ZN(U2917) );
  AOI22_X1 U7077 ( .A1(n6067), .A2(LWORD_REG_5__SCAN_IN), .B1(n6062), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6060) );
  OAI21_X1 U7078 ( .B1(n6125), .B2(n6069), .A(n6060), .ZN(U2918) );
  INV_X1 U7079 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6122) );
  AOI22_X1 U7080 ( .A1(n6067), .A2(LWORD_REG_4__SCAN_IN), .B1(n6062), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6061) );
  OAI21_X1 U7081 ( .B1(n6122), .B2(n6069), .A(n6061), .ZN(U2919) );
  AOI22_X1 U7082 ( .A1(n6067), .A2(LWORD_REG_3__SCAN_IN), .B1(n6062), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6063) );
  OAI21_X1 U7083 ( .B1(n6119), .B2(n6069), .A(n6063), .ZN(U2920) );
  AOI22_X1 U7084 ( .A1(n6067), .A2(LWORD_REG_2__SCAN_IN), .B1(n6066), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6064) );
  OAI21_X1 U7085 ( .B1(n6116), .B2(n6069), .A(n6064), .ZN(U2921) );
  AOI22_X1 U7086 ( .A1(n6067), .A2(LWORD_REG_1__SCAN_IN), .B1(n6066), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6065) );
  OAI21_X1 U7087 ( .B1(n6113), .B2(n6069), .A(n6065), .ZN(U2922) );
  AOI22_X1 U7088 ( .A1(n6067), .A2(LWORD_REG_0__SCAN_IN), .B1(n6066), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6068) );
  OAI21_X1 U7089 ( .B1(n6110), .B2(n6069), .A(n6068), .ZN(U2923) );
  NAND2_X2 U7090 ( .A1(n6071), .A2(n6070), .ZN(n6154) );
  INV_X1 U7091 ( .A(n6072), .ZN(n6073) );
  AND2_X1 U7092 ( .A1(n6151), .A2(DATAI_0_), .ZN(n6108) );
  AOI21_X1 U7093 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n6088), .A(n6108), .ZN(n6074) );
  OAI21_X1 U7094 ( .B1(n6075), .B2(n6154), .A(n6074), .ZN(U2924) );
  AND2_X1 U7095 ( .A1(n6151), .A2(DATAI_1_), .ZN(n6111) );
  AOI21_X1 U7096 ( .B1(UWORD_REG_1__SCAN_IN), .B2(n6088), .A(n6111), .ZN(n6076) );
  OAI21_X1 U7097 ( .B1(n6077), .B2(n6154), .A(n6076), .ZN(U2925) );
  AND2_X1 U7098 ( .A1(n6151), .A2(DATAI_2_), .ZN(n6114) );
  AOI21_X1 U7099 ( .B1(UWORD_REG_2__SCAN_IN), .B2(n6152), .A(n6114), .ZN(n6078) );
  OAI21_X1 U7100 ( .B1(n6079), .B2(n6154), .A(n6078), .ZN(U2926) );
  AND2_X1 U7101 ( .A1(n6151), .A2(DATAI_3_), .ZN(n6117) );
  AOI21_X1 U7102 ( .B1(UWORD_REG_3__SCAN_IN), .B2(n6088), .A(n6117), .ZN(n6080) );
  OAI21_X1 U7103 ( .B1(n6081), .B2(n6154), .A(n6080), .ZN(U2927) );
  INV_X1 U7104 ( .A(DATAI_4_), .ZN(n6082) );
  NOR2_X1 U7105 ( .A1(n6105), .A2(n6082), .ZN(n6120) );
  AOI21_X1 U7106 ( .B1(UWORD_REG_4__SCAN_IN), .B2(n6088), .A(n6120), .ZN(n6083) );
  OAI21_X1 U7107 ( .B1(n6084), .B2(n6154), .A(n6083), .ZN(U2928) );
  AND2_X1 U7108 ( .A1(n6151), .A2(DATAI_5_), .ZN(n6123) );
  AOI21_X1 U7109 ( .B1(UWORD_REG_5__SCAN_IN), .B2(n6152), .A(n6123), .ZN(n6085) );
  OAI21_X1 U7110 ( .B1(n6086), .B2(n6154), .A(n6085), .ZN(U2929) );
  NOR2_X1 U7111 ( .A1(n6105), .A2(n6087), .ZN(n6126) );
  AOI21_X1 U7112 ( .B1(UWORD_REG_6__SCAN_IN), .B2(n6088), .A(n6126), .ZN(n6089) );
  OAI21_X1 U7113 ( .B1(n6090), .B2(n6154), .A(n6089), .ZN(U2930) );
  AND2_X1 U7114 ( .A1(n6151), .A2(DATAI_7_), .ZN(n6128) );
  AOI21_X1 U7115 ( .B1(UWORD_REG_7__SCAN_IN), .B2(n6152), .A(n6128), .ZN(n6091) );
  OAI21_X1 U7116 ( .B1(n6092), .B2(n6154), .A(n6091), .ZN(U2931) );
  AND2_X1 U7117 ( .A1(n6151), .A2(DATAI_8_), .ZN(n6131) );
  AOI21_X1 U7118 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n6152), .A(n6131), .ZN(n6093) );
  OAI21_X1 U7119 ( .B1(n3972), .B2(n6154), .A(n6093), .ZN(U2932) );
  AND2_X1 U7120 ( .A1(n6151), .A2(DATAI_9_), .ZN(n6134) );
  AOI21_X1 U7121 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6152), .A(n6134), .ZN(n6094) );
  OAI21_X1 U7122 ( .B1(n6095), .B2(n6154), .A(n6094), .ZN(U2933) );
  AND2_X1 U7123 ( .A1(n6151), .A2(DATAI_10_), .ZN(n6137) );
  AOI21_X1 U7124 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n6152), .A(n6137), .ZN(
        n6096) );
  OAI21_X1 U7125 ( .B1(n6097), .B2(n6154), .A(n6096), .ZN(U2934) );
  AND2_X1 U7126 ( .A1(n6151), .A2(DATAI_11_), .ZN(n6140) );
  AOI21_X1 U7127 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n6152), .A(n6140), .ZN(
        n6098) );
  OAI21_X1 U7128 ( .B1(n6099), .B2(n6154), .A(n6098), .ZN(U2935) );
  AND2_X1 U7129 ( .A1(n6151), .A2(DATAI_12_), .ZN(n6143) );
  AOI21_X1 U7130 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6152), .A(n6143), .ZN(
        n6100) );
  OAI21_X1 U7131 ( .B1(n6101), .B2(n6154), .A(n6100), .ZN(U2936) );
  AND2_X1 U7132 ( .A1(n6151), .A2(DATAI_13_), .ZN(n6145) );
  AOI21_X1 U7133 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n6152), .A(n6145), .ZN(
        n6102) );
  OAI21_X1 U7134 ( .B1(n6103), .B2(n6154), .A(n6102), .ZN(U2937) );
  INV_X1 U7135 ( .A(DATAI_14_), .ZN(n6104) );
  NOR2_X1 U7136 ( .A1(n6105), .A2(n6104), .ZN(n6148) );
  AOI21_X1 U7137 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6152), .A(n6148), .ZN(
        n6106) );
  OAI21_X1 U7138 ( .B1(n6107), .B2(n6154), .A(n6106), .ZN(U2938) );
  AOI21_X1 U7139 ( .B1(LWORD_REG_0__SCAN_IN), .B2(n6152), .A(n6108), .ZN(n6109) );
  OAI21_X1 U7140 ( .B1(n6110), .B2(n6154), .A(n6109), .ZN(U2939) );
  AOI21_X1 U7141 ( .B1(LWORD_REG_1__SCAN_IN), .B2(n6152), .A(n6111), .ZN(n6112) );
  OAI21_X1 U7142 ( .B1(n6113), .B2(n6154), .A(n6112), .ZN(U2940) );
  AOI21_X1 U7143 ( .B1(LWORD_REG_2__SCAN_IN), .B2(n6152), .A(n6114), .ZN(n6115) );
  OAI21_X1 U7144 ( .B1(n6116), .B2(n6154), .A(n6115), .ZN(U2941) );
  AOI21_X1 U7145 ( .B1(LWORD_REG_3__SCAN_IN), .B2(n6152), .A(n6117), .ZN(n6118) );
  OAI21_X1 U7146 ( .B1(n6119), .B2(n6154), .A(n6118), .ZN(U2942) );
  AOI21_X1 U7147 ( .B1(LWORD_REG_4__SCAN_IN), .B2(n6152), .A(n6120), .ZN(n6121) );
  OAI21_X1 U7148 ( .B1(n6122), .B2(n6154), .A(n6121), .ZN(U2943) );
  AOI21_X1 U7149 ( .B1(LWORD_REG_5__SCAN_IN), .B2(n6152), .A(n6123), .ZN(n6124) );
  OAI21_X1 U7150 ( .B1(n6125), .B2(n6154), .A(n6124), .ZN(U2944) );
  AOI21_X1 U7151 ( .B1(LWORD_REG_6__SCAN_IN), .B2(n6152), .A(n6126), .ZN(n6127) );
  OAI21_X1 U7152 ( .B1(n4904), .B2(n6154), .A(n6127), .ZN(U2945) );
  AOI21_X1 U7153 ( .B1(LWORD_REG_7__SCAN_IN), .B2(n6152), .A(n6128), .ZN(n6129) );
  OAI21_X1 U7154 ( .B1(n6130), .B2(n6154), .A(n6129), .ZN(U2946) );
  AOI21_X1 U7155 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n6152), .A(n6131), .ZN(n6132) );
  OAI21_X1 U7156 ( .B1(n6133), .B2(n6154), .A(n6132), .ZN(U2947) );
  AOI21_X1 U7157 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n6152), .A(n6134), .ZN(n6135) );
  OAI21_X1 U7158 ( .B1(n6136), .B2(n6154), .A(n6135), .ZN(U2948) );
  AOI21_X1 U7159 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6152), .A(n6137), .ZN(
        n6138) );
  OAI21_X1 U7160 ( .B1(n6139), .B2(n6154), .A(n6138), .ZN(U2949) );
  AOI21_X1 U7161 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n6152), .A(n6140), .ZN(
        n6141) );
  OAI21_X1 U7162 ( .B1(n6142), .B2(n6154), .A(n6141), .ZN(U2950) );
  AOI21_X1 U7163 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n6152), .A(n6143), .ZN(
        n6144) );
  OAI21_X1 U7164 ( .B1(n3737), .B2(n6154), .A(n6144), .ZN(U2951) );
  AOI21_X1 U7165 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n6152), .A(n6145), .ZN(
        n6146) );
  OAI21_X1 U7166 ( .B1(n6147), .B2(n6154), .A(n6146), .ZN(U2952) );
  AOI21_X1 U7167 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6152), .A(n6148), .ZN(
        n6149) );
  OAI21_X1 U7168 ( .B1(n6150), .B2(n6154), .A(n6149), .ZN(U2953) );
  AOI22_X1 U7169 ( .A1(n6152), .A2(LWORD_REG_15__SCAN_IN), .B1(n6151), .B2(
        DATAI_15_), .ZN(n6153) );
  OAI21_X1 U7170 ( .B1(n6155), .B2(n6154), .A(n6153), .ZN(U2954) );
  AOI22_X1 U7171 ( .A1(n6215), .A2(REIP_REG_2__SCAN_IN), .B1(n6156), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6164) );
  NAND2_X1 U7172 ( .A1(n6159), .A2(n6158), .ZN(n6160) );
  XOR2_X1 U7173 ( .A(n2994), .B(n6160), .Z(n6214) );
  AOI22_X1 U7174 ( .A1(n6162), .A2(n6161), .B1(n6214), .B2(n6173), .ZN(n6163)
         );
  OAI211_X1 U7175 ( .C1(n6166), .C2(n6165), .A(n6164), .B(n6163), .ZN(U2984)
         );
  INV_X1 U7176 ( .A(n6167), .ZN(n6169) );
  AOI21_X1 U7177 ( .B1(n6169), .B2(n6232), .A(n6168), .ZN(n6228) );
  NAND2_X1 U7178 ( .A1(n6171), .A2(n6170), .ZN(n6172) );
  AOI22_X1 U7179 ( .A1(n6228), .A2(n6173), .B1(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6172), .ZN(n6174) );
  NAND2_X1 U7180 ( .A1(n6215), .A2(REIP_REG_0__SCAN_IN), .ZN(n6222) );
  OAI211_X1 U7181 ( .C1(n6176), .C2(n6175), .A(n6174), .B(n6222), .ZN(U2986)
         );
  INV_X1 U7182 ( .A(n6177), .ZN(n6185) );
  INV_X1 U7183 ( .A(n6178), .ZN(n6180) );
  AOI21_X1 U7184 ( .B1(n6210), .B2(n6180), .A(n6179), .ZN(n6184) );
  AOI22_X1 U7185 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6182), .B1(n6227), .B2(n6181), .ZN(n6183) );
  OAI211_X1 U7186 ( .C1(INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n6185), .A(n6184), .B(n6183), .ZN(U3007) );
  INV_X1 U7187 ( .A(n6186), .ZN(n6195) );
  INV_X1 U7188 ( .A(n6187), .ZN(n6189) );
  AOI21_X1 U7189 ( .B1(n6210), .B2(n6189), .A(n6188), .ZN(n6193) );
  AOI22_X1 U7190 ( .A1(n6191), .A2(n6227), .B1(n6190), .B2(n6194), .ZN(n6192)
         );
  OAI211_X1 U7191 ( .C1(n6195), .C2(n6194), .A(n6193), .B(n6192), .ZN(U3009)
         );
  AOI21_X1 U7192 ( .B1(n6210), .B2(n6197), .A(n6196), .ZN(n6198) );
  OAI21_X1 U7193 ( .B1(n6199), .B2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6198), 
        .ZN(n6200) );
  AOI21_X1 U7194 ( .B1(n6201), .B2(n6227), .A(n6200), .ZN(n6202) );
  OAI21_X1 U7195 ( .B1(n6204), .B2(n6203), .A(n6202), .ZN(U3011) );
  INV_X1 U7196 ( .A(n6205), .ZN(n6211) );
  OAI21_X1 U7197 ( .B1(n6207), .B2(n6216), .A(n6206), .ZN(n6208) );
  AOI22_X1 U7198 ( .A1(n6211), .A2(n6210), .B1(n6209), .B2(n6208), .ZN(n6221)
         );
  INV_X1 U7199 ( .A(n6212), .ZN(n6213) );
  AOI22_X1 U7200 ( .A1(n6214), .A2(n6227), .B1(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6213), .ZN(n6220) );
  NAND2_X1 U7201 ( .A1(n6215), .A2(REIP_REG_2__SCAN_IN), .ZN(n6219) );
  NAND3_X1 U7202 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6217), .A3(n6216), 
        .ZN(n6218) );
  NAND4_X1 U7203 ( .A1(n6221), .A2(n6220), .A3(n6219), .A4(n6218), .ZN(U3016)
         );
  OAI211_X1 U7204 ( .C1(n6225), .C2(n6224), .A(n6223), .B(n6222), .ZN(n6226)
         );
  AOI21_X1 U7205 ( .B1(n6228), .B2(n6227), .A(n6226), .ZN(n6229) );
  OAI221_X1 U7206 ( .B1(n6232), .B2(n6231), .C1(n6232), .C2(n6230), .A(n6229), 
        .ZN(U3018) );
  NOR2_X1 U7207 ( .A1(n6234), .A2(n6233), .ZN(U3019) );
  NOR3_X1 U7208 ( .A1(n6237), .A2(n6236), .A3(n6235), .ZN(n6238) );
  NOR2_X1 U7209 ( .A1(n6238), .A2(n6586), .ZN(n6245) );
  NAND2_X1 U7210 ( .A1(n6239), .A2(n6370), .ZN(n6241) );
  INV_X1 U7211 ( .A(n6372), .ZN(n6240) );
  NAND2_X1 U7212 ( .A1(n6240), .A2(n6468), .ZN(n6244) );
  NAND2_X1 U7213 ( .A1(n6241), .A2(n6244), .ZN(n6248) );
  AOI22_X1 U7214 ( .A1(n6245), .A2(n6248), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6242), .ZN(n6270) );
  INV_X1 U7215 ( .A(n6244), .ZN(n6264) );
  AOI22_X1 U7216 ( .A1(n6265), .A2(n6384), .B1(n6375), .B2(n6264), .ZN(n6251)
         );
  INV_X1 U7217 ( .A(n6245), .ZN(n6249) );
  AOI21_X1 U7218 ( .B1(n6586), .B2(n6246), .A(n6379), .ZN(n6247) );
  AOI22_X1 U7219 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6267), .B1(n6376), 
        .B2(n6266), .ZN(n6250) );
  OAI211_X1 U7220 ( .C1(n6270), .C2(n6387), .A(n6251), .B(n6250), .ZN(U3044)
         );
  AOI22_X1 U7221 ( .A1(n6265), .A2(n6390), .B1(n6388), .B2(n6264), .ZN(n6253)
         );
  AOI22_X1 U7222 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6267), .B1(n6389), 
        .B2(n6266), .ZN(n6252) );
  OAI211_X1 U7223 ( .C1(n6270), .C2(n6393), .A(n6253), .B(n6252), .ZN(U3045)
         );
  AOI22_X1 U7224 ( .A1(n6265), .A2(n6394), .B1(n6430), .B2(n6264), .ZN(n6255)
         );
  AOI22_X1 U7225 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6267), .B1(n6432), 
        .B2(n6266), .ZN(n6254) );
  OAI211_X1 U7226 ( .C1(n6270), .C2(n6397), .A(n6255), .B(n6254), .ZN(U3046)
         );
  AOI22_X1 U7227 ( .A1(n6265), .A2(n6399), .B1(n6398), .B2(n6264), .ZN(n6257)
         );
  AOI22_X1 U7228 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6267), .B1(n6400), 
        .B2(n6266), .ZN(n6256) );
  OAI211_X1 U7229 ( .C1(n6270), .C2(n6403), .A(n6257), .B(n6256), .ZN(U3047)
         );
  AOI22_X1 U7230 ( .A1(n6265), .A2(n6404), .B1(n6436), .B2(n6264), .ZN(n6259)
         );
  AOI22_X1 U7231 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6267), .B1(n6438), 
        .B2(n6266), .ZN(n6258) );
  OAI211_X1 U7232 ( .C1(n6270), .C2(n6407), .A(n6259), .B(n6258), .ZN(U3048)
         );
  AOI22_X1 U7233 ( .A1(n6265), .A2(n6410), .B1(n6408), .B2(n6264), .ZN(n6261)
         );
  AOI22_X1 U7234 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6267), .B1(n6409), 
        .B2(n6266), .ZN(n6260) );
  OAI211_X1 U7235 ( .C1(n6270), .C2(n6413), .A(n6261), .B(n6260), .ZN(U3049)
         );
  AOI22_X1 U7236 ( .A1(n6265), .A2(n6415), .B1(n6414), .B2(n6264), .ZN(n6263)
         );
  AOI22_X1 U7237 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6267), .B1(n6416), 
        .B2(n6266), .ZN(n6262) );
  OAI211_X1 U7238 ( .C1(n6270), .C2(n6419), .A(n6263), .B(n6262), .ZN(U3050)
         );
  AOI22_X1 U7239 ( .A1(n6265), .A2(n6423), .B1(n6443), .B2(n6264), .ZN(n6269)
         );
  AOI22_X1 U7240 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6267), .B1(n6447), 
        .B2(n6266), .ZN(n6268) );
  OAI211_X1 U7241 ( .C1(n6270), .C2(n6427), .A(n6269), .B(n6268), .ZN(U3051)
         );
  INV_X1 U7242 ( .A(n6273), .ZN(n6278) );
  NAND3_X1 U7243 ( .A1(n6275), .A2(n6274), .A3(n6468), .ZN(n6276) );
  OAI21_X1 U7244 ( .B1(n6278), .B2(n6277), .A(n6276), .ZN(n6313) );
  NAND2_X1 U7245 ( .A1(n6454), .A2(n6329), .ZN(n6284) );
  INV_X1 U7246 ( .A(n6284), .ZN(n6312) );
  AOI22_X1 U7247 ( .A1(n6279), .A2(n6313), .B1(n6375), .B2(n6312), .ZN(n6289)
         );
  NOR3_X1 U7248 ( .A1(n6345), .A2(n6314), .A3(n6586), .ZN(n6281) );
  NOR2_X1 U7249 ( .A1(n6281), .A2(n6280), .ZN(n6287) );
  NOR2_X1 U7250 ( .A1(n6283), .A2(n6282), .ZN(n6322) );
  AOI21_X1 U7251 ( .B1(n6284), .B2(STATE2_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6285) );
  OAI211_X1 U7252 ( .C1(n6287), .C2(n6322), .A(n6286), .B(n6285), .ZN(n6315)
         );
  AOI22_X1 U7253 ( .A1(n6315), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6384), 
        .B2(n6314), .ZN(n6288) );
  OAI211_X1 U7254 ( .C1(n6290), .C2(n6318), .A(n6289), .B(n6288), .ZN(U3068)
         );
  AOI22_X1 U7255 ( .A1(n6291), .A2(n6313), .B1(n6388), .B2(n6312), .ZN(n6293)
         );
  AOI22_X1 U7256 ( .A1(n6315), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6390), 
        .B2(n6314), .ZN(n6292) );
  OAI211_X1 U7257 ( .C1(n6294), .C2(n6318), .A(n6293), .B(n6292), .ZN(U3069)
         );
  AOI22_X1 U7258 ( .A1(n6431), .A2(n6313), .B1(n6430), .B2(n6312), .ZN(n6296)
         );
  AOI22_X1 U7259 ( .A1(n6315), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6394), 
        .B2(n6314), .ZN(n6295) );
  OAI211_X1 U7260 ( .C1(n6297), .C2(n6318), .A(n6296), .B(n6295), .ZN(U3070)
         );
  AOI22_X1 U7261 ( .A1(n6298), .A2(n6313), .B1(n6398), .B2(n6312), .ZN(n6300)
         );
  AOI22_X1 U7262 ( .A1(n6315), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6399), 
        .B2(n6314), .ZN(n6299) );
  OAI211_X1 U7263 ( .C1(n6301), .C2(n6318), .A(n6300), .B(n6299), .ZN(U3071)
         );
  AOI22_X1 U7264 ( .A1(n6437), .A2(n6313), .B1(n6436), .B2(n6312), .ZN(n6303)
         );
  AOI22_X1 U7265 ( .A1(n6315), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6404), 
        .B2(n6314), .ZN(n6302) );
  OAI211_X1 U7266 ( .C1(n6304), .C2(n6318), .A(n6303), .B(n6302), .ZN(U3072)
         );
  AOI22_X1 U7267 ( .A1(n6305), .A2(n6313), .B1(n6408), .B2(n6312), .ZN(n6307)
         );
  AOI22_X1 U7268 ( .A1(n6315), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6410), 
        .B2(n6314), .ZN(n6306) );
  OAI211_X1 U7269 ( .C1(n6308), .C2(n6318), .A(n6307), .B(n6306), .ZN(U3073)
         );
  AOI22_X1 U7270 ( .A1(n6356), .A2(n6313), .B1(n6414), .B2(n6312), .ZN(n6310)
         );
  AOI22_X1 U7271 ( .A1(n6315), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6415), 
        .B2(n6314), .ZN(n6309) );
  OAI211_X1 U7272 ( .C1(n6311), .C2(n6318), .A(n6310), .B(n6309), .ZN(U3074)
         );
  AOI22_X1 U7273 ( .A1(n6445), .A2(n6313), .B1(n6443), .B2(n6312), .ZN(n6317)
         );
  AOI22_X1 U7274 ( .A1(n6315), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6423), 
        .B2(n6314), .ZN(n6316) );
  OAI211_X1 U7275 ( .C1(n6319), .C2(n6318), .A(n6317), .B(n6316), .ZN(U3075)
         );
  AND2_X1 U7276 ( .A1(n6320), .A2(n6328), .ZN(n6325) );
  INV_X1 U7277 ( .A(n6321), .ZN(n6344) );
  AOI21_X1 U7278 ( .B1(n6322), .B2(n6370), .A(n6344), .ZN(n6324) );
  INV_X1 U7279 ( .A(n6324), .ZN(n6323) );
  AOI22_X1 U7280 ( .A1(n6325), .A2(n6323), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6329), .ZN(n6350) );
  AOI22_X1 U7281 ( .A1(n6346), .A2(n6376), .B1(n6344), .B2(n6375), .ZN(n6331)
         );
  NAND2_X1 U7282 ( .A1(n6325), .A2(n6324), .ZN(n6327) );
  OAI211_X1 U7283 ( .C1(n6329), .C2(n6328), .A(n6327), .B(n6326), .ZN(n6347)
         );
  AOI22_X1 U7284 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6347), .B1(n6384), 
        .B2(n6345), .ZN(n6330) );
  OAI211_X1 U7285 ( .C1(n6350), .C2(n6387), .A(n6331), .B(n6330), .ZN(U3076)
         );
  AOI22_X1 U7286 ( .A1(n6346), .A2(n6389), .B1(n6344), .B2(n6388), .ZN(n6333)
         );
  AOI22_X1 U7287 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6347), .B1(n6390), 
        .B2(n6345), .ZN(n6332) );
  OAI211_X1 U7288 ( .C1(n6350), .C2(n6393), .A(n6333), .B(n6332), .ZN(U3077)
         );
  AOI22_X1 U7289 ( .A1(n6345), .A2(n6394), .B1(n6344), .B2(n6430), .ZN(n6335)
         );
  AOI22_X1 U7290 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6347), .B1(n6432), 
        .B2(n6346), .ZN(n6334) );
  OAI211_X1 U7291 ( .C1(n6350), .C2(n6397), .A(n6335), .B(n6334), .ZN(U3078)
         );
  AOI22_X1 U7292 ( .A1(n6345), .A2(n6399), .B1(n6344), .B2(n6398), .ZN(n6337)
         );
  AOI22_X1 U7293 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6347), .B1(n6400), 
        .B2(n6346), .ZN(n6336) );
  OAI211_X1 U7294 ( .C1(n6350), .C2(n6403), .A(n6337), .B(n6336), .ZN(U3079)
         );
  AOI22_X1 U7295 ( .A1(n6345), .A2(n6404), .B1(n6344), .B2(n6436), .ZN(n6339)
         );
  AOI22_X1 U7296 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6347), .B1(n6438), 
        .B2(n6346), .ZN(n6338) );
  OAI211_X1 U7297 ( .C1(n6350), .C2(n6407), .A(n6339), .B(n6338), .ZN(U3080)
         );
  AOI22_X1 U7298 ( .A1(n6345), .A2(n6410), .B1(n6344), .B2(n6408), .ZN(n6341)
         );
  AOI22_X1 U7299 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6347), .B1(n6409), 
        .B2(n6346), .ZN(n6340) );
  OAI211_X1 U7300 ( .C1(n6350), .C2(n6413), .A(n6341), .B(n6340), .ZN(U3081)
         );
  AOI22_X1 U7301 ( .A1(n6346), .A2(n6416), .B1(n6344), .B2(n6414), .ZN(n6343)
         );
  AOI22_X1 U7302 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6347), .B1(n6415), 
        .B2(n6345), .ZN(n6342) );
  OAI211_X1 U7303 ( .C1(n6350), .C2(n6419), .A(n6343), .B(n6342), .ZN(U3082)
         );
  AOI22_X1 U7304 ( .A1(n6345), .A2(n6423), .B1(n6344), .B2(n6443), .ZN(n6349)
         );
  AOI22_X1 U7305 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6347), .B1(n6447), 
        .B2(n6346), .ZN(n6348) );
  OAI211_X1 U7306 ( .C1(n6350), .C2(n6427), .A(n6349), .B(n6348), .ZN(U3083)
         );
  INV_X1 U7307 ( .A(n6351), .ZN(n6361) );
  AOI22_X1 U7308 ( .A1(n6431), .A2(n6361), .B1(n6430), .B2(n6360), .ZN(n6353)
         );
  AOI22_X1 U7309 ( .A1(n6363), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6432), 
        .B2(n6362), .ZN(n6352) );
  OAI211_X1 U7310 ( .C1(n6435), .C2(n6366), .A(n6353), .B(n6352), .ZN(U3086)
         );
  AOI22_X1 U7311 ( .A1(n6437), .A2(n6361), .B1(n6436), .B2(n6360), .ZN(n6355)
         );
  AOI22_X1 U7312 ( .A1(n6363), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6438), 
        .B2(n6362), .ZN(n6354) );
  OAI211_X1 U7313 ( .C1(n6441), .C2(n6366), .A(n6355), .B(n6354), .ZN(U3088)
         );
  AOI22_X1 U7314 ( .A1(n6356), .A2(n6361), .B1(n6414), .B2(n6360), .ZN(n6358)
         );
  AOI22_X1 U7315 ( .A1(n6363), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6416), 
        .B2(n6362), .ZN(n6357) );
  OAI211_X1 U7316 ( .C1(n6359), .C2(n6366), .A(n6358), .B(n6357), .ZN(U3090)
         );
  AOI22_X1 U7317 ( .A1(n6445), .A2(n6361), .B1(n6443), .B2(n6360), .ZN(n6365)
         );
  AOI22_X1 U7318 ( .A1(n6363), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6447), 
        .B2(n6362), .ZN(n6364) );
  OAI211_X1 U7319 ( .C1(n6452), .C2(n6366), .A(n6365), .B(n6364), .ZN(U3091)
         );
  INV_X1 U7320 ( .A(n6367), .ZN(n6369) );
  AOI21_X1 U7321 ( .B1(n6369), .B2(n6368), .A(n6586), .ZN(n6377) );
  NAND2_X1 U7322 ( .A1(n6371), .A2(n6370), .ZN(n6374) );
  NOR2_X1 U7323 ( .A1(n6372), .A2(n6468), .ZN(n6420) );
  INV_X1 U7324 ( .A(n6420), .ZN(n6373) );
  NAND2_X1 U7325 ( .A1(n6374), .A2(n6373), .ZN(n6382) );
  AOI22_X1 U7326 ( .A1(n6377), .A2(n6382), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6378), .ZN(n6428) );
  AOI22_X1 U7327 ( .A1(n6421), .A2(n6376), .B1(n6375), .B2(n6420), .ZN(n6386)
         );
  INV_X1 U7328 ( .A(n6377), .ZN(n6383) );
  INV_X1 U7329 ( .A(n6378), .ZN(n6380) );
  AOI21_X1 U7330 ( .B1(n6586), .B2(n6380), .A(n6379), .ZN(n6381) );
  OAI21_X1 U7331 ( .B1(n6383), .B2(n6382), .A(n6381), .ZN(n6424) );
  AOI22_X1 U7332 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6424), .B1(n6384), 
        .B2(n6422), .ZN(n6385) );
  OAI211_X1 U7333 ( .C1(n6428), .C2(n6387), .A(n6386), .B(n6385), .ZN(U3108)
         );
  AOI22_X1 U7334 ( .A1(n6421), .A2(n6389), .B1(n6388), .B2(n6420), .ZN(n6392)
         );
  AOI22_X1 U7335 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6424), .B1(n6390), 
        .B2(n6422), .ZN(n6391) );
  OAI211_X1 U7336 ( .C1(n6428), .C2(n6393), .A(n6392), .B(n6391), .ZN(U3109)
         );
  AOI22_X1 U7337 ( .A1(n6422), .A2(n6394), .B1(n6430), .B2(n6420), .ZN(n6396)
         );
  AOI22_X1 U7338 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6424), .B1(n6432), 
        .B2(n6421), .ZN(n6395) );
  OAI211_X1 U7339 ( .C1(n6428), .C2(n6397), .A(n6396), .B(n6395), .ZN(U3110)
         );
  AOI22_X1 U7340 ( .A1(n6422), .A2(n6399), .B1(n6398), .B2(n6420), .ZN(n6402)
         );
  AOI22_X1 U7341 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6424), .B1(n6400), 
        .B2(n6421), .ZN(n6401) );
  OAI211_X1 U7342 ( .C1(n6428), .C2(n6403), .A(n6402), .B(n6401), .ZN(U3111)
         );
  AOI22_X1 U7343 ( .A1(n6422), .A2(n6404), .B1(n6436), .B2(n6420), .ZN(n6406)
         );
  AOI22_X1 U7344 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6424), .B1(n6438), 
        .B2(n6421), .ZN(n6405) );
  OAI211_X1 U7345 ( .C1(n6428), .C2(n6407), .A(n6406), .B(n6405), .ZN(U3112)
         );
  AOI22_X1 U7346 ( .A1(n6421), .A2(n6409), .B1(n6408), .B2(n6420), .ZN(n6412)
         );
  AOI22_X1 U7347 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6424), .B1(n6410), 
        .B2(n6422), .ZN(n6411) );
  OAI211_X1 U7348 ( .C1(n6428), .C2(n6413), .A(n6412), .B(n6411), .ZN(U3113)
         );
  AOI22_X1 U7349 ( .A1(n6422), .A2(n6415), .B1(n6414), .B2(n6420), .ZN(n6418)
         );
  AOI22_X1 U7350 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6424), .B1(n6416), 
        .B2(n6421), .ZN(n6417) );
  OAI211_X1 U7351 ( .C1(n6428), .C2(n6419), .A(n6418), .B(n6417), .ZN(U3114)
         );
  AOI22_X1 U7352 ( .A1(n6421), .A2(n6447), .B1(n6443), .B2(n6420), .ZN(n6426)
         );
  AOI22_X1 U7353 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6424), .B1(n6423), 
        .B2(n6422), .ZN(n6425) );
  OAI211_X1 U7354 ( .C1(n6428), .C2(n6427), .A(n6426), .B(n6425), .ZN(U3115)
         );
  INV_X1 U7355 ( .A(n6429), .ZN(n6444) );
  AOI22_X1 U7356 ( .A1(n6431), .A2(n6444), .B1(n6430), .B2(n6442), .ZN(n6434)
         );
  AOI22_X1 U7357 ( .A1(n6448), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n6432), 
        .B2(n6446), .ZN(n6433) );
  OAI211_X1 U7358 ( .C1(n6435), .C2(n6451), .A(n6434), .B(n6433), .ZN(U3118)
         );
  AOI22_X1 U7359 ( .A1(n6437), .A2(n6444), .B1(n6436), .B2(n6442), .ZN(n6440)
         );
  AOI22_X1 U7360 ( .A1(n6448), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n6438), 
        .B2(n6446), .ZN(n6439) );
  OAI211_X1 U7361 ( .C1(n6441), .C2(n6451), .A(n6440), .B(n6439), .ZN(U3120)
         );
  AOI22_X1 U7362 ( .A1(n6445), .A2(n6444), .B1(n6443), .B2(n6442), .ZN(n6450)
         );
  AOI22_X1 U7363 ( .A1(n6448), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n6447), 
        .B2(n6446), .ZN(n6449) );
  OAI211_X1 U7364 ( .C1(n6452), .C2(n6451), .A(n6450), .B(n6449), .ZN(U3123)
         );
  INV_X1 U7365 ( .A(n6463), .ZN(n6465) );
  INV_X1 U7366 ( .A(n6453), .ZN(n6456) );
  NOR3_X1 U7367 ( .A1(n6456), .A2(n6455), .A3(n6454), .ZN(n6460) );
  INV_X1 U7368 ( .A(n6457), .ZN(n6458) );
  OAI22_X1 U7369 ( .A1(n6460), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n6459), .B2(n6458), .ZN(n6462) );
  NAND2_X1 U7370 ( .A1(n6460), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6461) );
  OAI211_X1 U7371 ( .C1(n6463), .C2(n4695), .A(n6462), .B(n6461), .ZN(n6464)
         );
  OAI21_X1 U7372 ( .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6465), .A(n6464), 
        .ZN(n6466) );
  AOI222_X1 U7373 ( .A1(n6468), .A2(n6467), .B1(n6468), .B2(n6466), .C1(n6467), 
        .C2(n6466), .ZN(n6477) );
  INV_X1 U7374 ( .A(MORE_REG_SCAN_IN), .ZN(n6470) );
  AOI21_X1 U7375 ( .B1(n6674), .B2(n6470), .A(n6469), .ZN(n6472) );
  NOR4_X1 U7376 ( .A1(n6474), .A2(n6473), .A3(n6472), .A4(n6471), .ZN(n6475)
         );
  OAI211_X1 U7377 ( .C1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n6477), .A(n6476), .B(n6475), .ZN(n6487) );
  OAI21_X1 U7378 ( .B1(n6493), .B2(n6728), .A(n6490), .ZN(n6478) );
  OAI211_X1 U7379 ( .C1(n6480), .C2(n6479), .A(STATE2_REG_2__SCAN_IN), .B(
        n6478), .ZN(n6482) );
  AOI221_X1 U7380 ( .B1(STATE2_REG_1__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(n6487), .C2(STATE2_REG_0__SCAN_IN), .A(n6482), .ZN(n6569) );
  AOI21_X1 U7381 ( .B1(READY_N), .B2(n6481), .A(n6569), .ZN(n6494) );
  OAI211_X1 U7382 ( .C1(n6583), .C2(n6483), .A(n6490), .B(n6482), .ZN(n6484)
         );
  INV_X1 U7383 ( .A(n6484), .ZN(n6485) );
  AOI211_X1 U7384 ( .C1(n6491), .C2(n6487), .A(n6486), .B(n6485), .ZN(n6488)
         );
  OAI221_X1 U7385 ( .B1(n6490), .B2(n6494), .C1(n6490), .C2(n6489), .A(n6488), 
        .ZN(U3148) );
  AOI21_X1 U7386 ( .B1(n6492), .B2(n6728), .A(n6491), .ZN(n6498) );
  NOR3_X1 U7387 ( .A1(n6494), .A2(n6493), .A3(n6501), .ZN(n6496) );
  NOR2_X1 U7388 ( .A1(n6496), .A2(n6495), .ZN(n6497) );
  OAI21_X1 U7389 ( .B1(n6569), .B2(n6498), .A(n6497), .ZN(U3149) );
  OAI211_X1 U7390 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6728), .A(n6570), .B(
        n6583), .ZN(n6500) );
  OAI21_X1 U7391 ( .B1(n6501), .B2(n6500), .A(n6499), .ZN(U3150) );
  AND2_X1 U7392 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6503), .ZN(U3151) );
  AND2_X1 U7393 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6503), .ZN(U3152) );
  AND2_X1 U7394 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6503), .ZN(U3153) );
  AND2_X1 U7395 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6503), .ZN(U3154) );
  AND2_X1 U7396 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6503), .ZN(U3155) );
  AND2_X1 U7397 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6503), .ZN(U3156) );
  AND2_X1 U7398 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6503), .ZN(U3157) );
  AND2_X1 U7399 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6503), .ZN(U3158) );
  AND2_X1 U7400 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6503), .ZN(U3159) );
  AND2_X1 U7401 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6503), .ZN(U3160) );
  AND2_X1 U7402 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6503), .ZN(U3161) );
  AND2_X1 U7403 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6503), .ZN(U3162) );
  AND2_X1 U7404 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6503), .ZN(U3163) );
  AND2_X1 U7405 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6503), .ZN(U3164) );
  AND2_X1 U7406 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6503), .ZN(U3165) );
  AND2_X1 U7407 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6503), .ZN(U3166) );
  AND2_X1 U7408 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6503), .ZN(U3167) );
  AND2_X1 U7409 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6502), .ZN(U3168) );
  AND2_X1 U7410 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6502), .ZN(U3169) );
  AND2_X1 U7411 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6502), .ZN(U3170) );
  AND2_X1 U7412 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6502), .ZN(U3171) );
  AND2_X1 U7413 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6502), .ZN(U3172) );
  AND2_X1 U7414 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6502), .ZN(U3173) );
  AND2_X1 U7415 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6502), .ZN(U3174) );
  AND2_X1 U7416 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6502), .ZN(U3175) );
  AND2_X1 U7417 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6502), .ZN(U3176) );
  AND2_X1 U7418 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6502), .ZN(U3177) );
  AND2_X1 U7419 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6502), .ZN(U3178) );
  AND2_X1 U7420 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6502), .ZN(U3179) );
  AND2_X1 U7421 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6503), .ZN(U3180) );
  INV_X1 U7422 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6511) );
  NOR2_X1 U7423 ( .A1(n6511), .A2(n6519), .ZN(n6514) );
  NAND2_X1 U7424 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6505) );
  NAND2_X1 U7425 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6510) );
  INV_X1 U7426 ( .A(HOLD), .ZN(n6731) );
  NOR2_X1 U7427 ( .A1(n6511), .A2(n6731), .ZN(n6506) );
  INV_X1 U7428 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6715) );
  INV_X1 U7429 ( .A(NA_N), .ZN(n6688) );
  AOI221_X1 U7430 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6688), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6517) );
  AOI221_X1 U7431 ( .B1(n6506), .B2(n6788), .C1(n6715), .C2(n6788), .A(n6517), 
        .ZN(n6504) );
  OAI221_X1 U7432 ( .B1(n6514), .B2(n6505), .C1(n6514), .C2(n6510), .A(n6504), 
        .ZN(U3181) );
  NOR2_X1 U7433 ( .A1(n4126), .A2(n6715), .ZN(n6507) );
  OAI21_X1 U7434 ( .B1(n6507), .B2(n6506), .A(n6505), .ZN(n6508) );
  NAND3_X1 U7435 ( .A1(n6509), .A2(n6510), .A3(n6508), .ZN(U3182) );
  INV_X1 U7436 ( .A(n6510), .ZN(n6515) );
  OAI221_X1 U7437 ( .B1(n6511), .B2(READY_N), .C1(n6511), .C2(n6688), .A(n6715), .ZN(n6512) );
  AOI21_X1 U7438 ( .B1(n6519), .B2(n6512), .A(n6731), .ZN(n6513) );
  AOI211_X1 U7439 ( .C1(n6515), .C2(n6514), .A(n4126), .B(n6513), .ZN(n6518)
         );
  NAND4_X1 U7440 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(STATE_REG_0__SCAN_IN), 
        .A3(n6515), .A4(n6688), .ZN(n6516) );
  OAI21_X1 U7441 ( .B1(n6518), .B2(n6517), .A(n6516), .ZN(U3183) );
  NOR2_X2 U7442 ( .A1(n6519), .A2(n6788), .ZN(n6562) );
  NAND2_X1 U7443 ( .A1(n6519), .A2(n6789), .ZN(n6564) );
  AOI22_X1 U7444 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6788), .ZN(n6520) );
  OAI21_X1 U7445 ( .B1(n5085), .B2(n6561), .A(n6520), .ZN(U3184) );
  AOI22_X1 U7446 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6788), .ZN(n6521) );
  OAI21_X1 U7447 ( .B1(n6523), .B2(n6564), .A(n6521), .ZN(U3185) );
  AOI22_X1 U7448 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6788), .ZN(n6522) );
  OAI21_X1 U7449 ( .B1(n6523), .B2(n6561), .A(n6522), .ZN(U3186) );
  AOI22_X1 U7450 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6788), .ZN(n6524) );
  OAI21_X1 U7451 ( .B1(n6525), .B2(n6561), .A(n6524), .ZN(U3187) );
  AOI22_X1 U7452 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6788), .ZN(n6526) );
  OAI21_X1 U7453 ( .B1(n6528), .B2(n6564), .A(n6526), .ZN(U3188) );
  AOI22_X1 U7454 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6788), .ZN(n6527) );
  OAI21_X1 U7455 ( .B1(n6528), .B2(n6561), .A(n6527), .ZN(U3189) );
  AOI22_X1 U7456 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6788), .ZN(n6529) );
  OAI21_X1 U7457 ( .B1(n6530), .B2(n6561), .A(n6529), .ZN(U3190) );
  AOI22_X1 U7458 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6788), .ZN(n6531) );
  OAI21_X1 U7459 ( .B1(n6533), .B2(n6564), .A(n6531), .ZN(U3191) );
  AOI22_X1 U7460 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6788), .ZN(n6532) );
  OAI21_X1 U7461 ( .B1(n6533), .B2(n6561), .A(n6532), .ZN(U3192) );
  AOI22_X1 U7462 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6788), .ZN(n6534) );
  OAI21_X1 U7463 ( .B1(n6535), .B2(n6561), .A(n6534), .ZN(U3193) );
  AOI22_X1 U7464 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6788), .ZN(n6536) );
  OAI21_X1 U7465 ( .B1(n6538), .B2(n6564), .A(n6536), .ZN(U3194) );
  AOI22_X1 U7466 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6788), .ZN(n6537) );
  OAI21_X1 U7467 ( .B1(n6538), .B2(n6561), .A(n6537), .ZN(U3195) );
  AOI22_X1 U7468 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6788), .ZN(n6539) );
  OAI21_X1 U7469 ( .B1(n6540), .B2(n6564), .A(n6539), .ZN(U3196) );
  AOI22_X1 U7470 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6788), .ZN(n6541) );
  OAI21_X1 U7471 ( .B1(n5639), .B2(n6564), .A(n6541), .ZN(U3197) );
  AOI22_X1 U7472 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6788), .ZN(n6542) );
  OAI21_X1 U7473 ( .B1(n5639), .B2(n6561), .A(n6542), .ZN(U3198) );
  AOI22_X1 U7474 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6788), .ZN(n6543) );
  OAI21_X1 U7475 ( .B1(n6544), .B2(n6564), .A(n6543), .ZN(U3199) );
  AOI22_X1 U7476 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6788), .ZN(n6545) );
  OAI21_X1 U7477 ( .B1(n6547), .B2(n6564), .A(n6545), .ZN(U3200) );
  AOI22_X1 U7478 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6788), .ZN(n6546) );
  OAI21_X1 U7479 ( .B1(n6547), .B2(n6561), .A(n6546), .ZN(U3201) );
  AOI22_X1 U7480 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6788), .ZN(n6548) );
  OAI21_X1 U7481 ( .B1(n6756), .B2(n6564), .A(n6548), .ZN(U3202) );
  AOI22_X1 U7482 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6788), .ZN(n6549) );
  OAI21_X1 U7483 ( .B1(n6734), .B2(n6564), .A(n6549), .ZN(U3203) );
  AOI22_X1 U7484 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6788), .ZN(n6550) );
  OAI21_X1 U7485 ( .B1(n6734), .B2(n6561), .A(n6550), .ZN(U3204) );
  AOI22_X1 U7486 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6788), .ZN(n6551) );
  OAI21_X1 U7487 ( .B1(n6552), .B2(n6561), .A(n6551), .ZN(U3205) );
  AOI22_X1 U7488 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6788), .ZN(n6553) );
  OAI21_X1 U7489 ( .B1(n6718), .B2(n6561), .A(n6553), .ZN(U3206) );
  AOI22_X1 U7490 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6788), .ZN(n6554) );
  OAI21_X1 U7491 ( .B1(n6687), .B2(n6561), .A(n6554), .ZN(U3207) );
  AOI22_X1 U7492 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6788), .ZN(n6555) );
  OAI21_X1 U7493 ( .B1(n6660), .B2(n6564), .A(n6555), .ZN(U3208) );
  AOI22_X1 U7494 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6788), .ZN(n6556) );
  OAI21_X1 U7495 ( .B1(n6660), .B2(n6561), .A(n6556), .ZN(U3209) );
  AOI22_X1 U7496 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6788), .ZN(n6557) );
  OAI21_X1 U7497 ( .B1(n6626), .B2(n6564), .A(n6557), .ZN(U3210) );
  AOI22_X1 U7498 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6788), .ZN(n6558) );
  OAI21_X1 U7499 ( .B1(n6626), .B2(n6561), .A(n6558), .ZN(U3211) );
  AOI22_X1 U7500 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6788), .ZN(n6560) );
  OAI21_X1 U7501 ( .B1(n6733), .B2(n6561), .A(n6560), .ZN(U3212) );
  AOI22_X1 U7502 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6788), .ZN(n6563) );
  OAI21_X1 U7503 ( .B1(n6691), .B2(n6564), .A(n6563), .ZN(U3213) );
  MUX2_X1 U7504 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6788), .Z(U3446) );
  MUX2_X1 U7505 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6788), .Z(U3447) );
  MUX2_X1 U7506 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6788), .Z(U3448) );
  OAI21_X1 U7507 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6568), .A(n6566), .ZN(
        n6565) );
  INV_X1 U7508 ( .A(n6565), .ZN(U3451) );
  OAI21_X1 U7509 ( .B1(n6568), .B2(n6567), .A(n6566), .ZN(U3452) );
  INV_X1 U7510 ( .A(n6569), .ZN(n6572) );
  OAI211_X1 U7511 ( .C1(n6573), .C2(n6572), .A(n6571), .B(n6570), .ZN(U3453)
         );
  AOI21_X1 U7512 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6574) );
  AOI22_X1 U7513 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6574), .B2(n5085), .ZN(n6576) );
  INV_X1 U7514 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6754) );
  AOI22_X1 U7515 ( .A1(n6578), .A2(n6576), .B1(n6754), .B2(n6575), .ZN(U3468)
         );
  INV_X1 U7516 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6630) );
  OAI21_X1 U7517 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6578), .ZN(n6577) );
  OAI21_X1 U7518 ( .B1(n6578), .B2(n6630), .A(n6577), .ZN(U3469) );
  OAI22_X1 U7519 ( .A1(n6788), .A2(n6673), .B1(W_R_N_REG_SCAN_IN), .B2(n6789), 
        .ZN(n6579) );
  INV_X1 U7520 ( .A(n6579), .ZN(U3470) );
  OAI211_X1 U7521 ( .C1(n6580), .C2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .B(n6728), .ZN(n6581) );
  OAI21_X1 U7522 ( .B1(n6582), .B2(n6581), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n6584) );
  NAND2_X1 U7523 ( .A1(n6584), .A2(n6583), .ZN(n6592) );
  INV_X1 U7524 ( .A(n6585), .ZN(n6590) );
  OAI211_X1 U7525 ( .C1(READY_N), .C2(n6588), .A(n6587), .B(n6586), .ZN(n6589)
         );
  NOR2_X1 U7526 ( .A1(n6590), .A2(n6589), .ZN(n6591) );
  MUX2_X1 U7527 ( .A(n6592), .B(REQUESTPENDING_REG_SCAN_IN), .S(n6591), .Z(
        U3472) );
  OAI22_X1 U7528 ( .A1(n6788), .A2(MEMORYFETCH_REG_SCAN_IN), .B1(
        M_IO_N_REG_SCAN_IN), .B2(n6789), .ZN(n6593) );
  INV_X1 U7529 ( .A(n6593), .ZN(U3473) );
  AOI22_X1 U7530 ( .A1(DATAI_6_), .A2(keyinput_f25), .B1(DATAI_29_), .B2(
        keyinput_f2), .ZN(n6594) );
  OAI221_X1 U7531 ( .B1(DATAI_6_), .B2(keyinput_f25), .C1(DATAI_29_), .C2(
        keyinput_f2), .A(n6594), .ZN(n6653) );
  AOI22_X1 U7532 ( .A1(DATAI_4_), .A2(keyinput_f27), .B1(REIP_REG_19__SCAN_IN), 
        .B2(keyinput_f63), .ZN(n6595) );
  OAI221_X1 U7533 ( .B1(DATAI_4_), .B2(keyinput_f27), .C1(REIP_REG_19__SCAN_IN), .C2(keyinput_f63), .A(n6595), .ZN(n6652) );
  AOI22_X1 U7534 ( .A1(keyinput_f49), .A2(BYTEENABLE_REG_2__SCAN_IN), .B1(
        REIP_REG_24__SCAN_IN), .B2(keyinput_f58), .ZN(n6596) );
  OAI221_X1 U7535 ( .B1(keyinput_f49), .B2(BYTEENABLE_REG_2__SCAN_IN), .C1(
        REIP_REG_24__SCAN_IN), .C2(keyinput_f58), .A(n6596), .ZN(n6603) );
  AOI22_X1 U7536 ( .A1(keyinput_f38), .A2(ADS_N_REG_SCAN_IN), .B1(DATAI_1_), 
        .B2(keyinput_f30), .ZN(n6597) );
  OAI221_X1 U7537 ( .B1(keyinput_f38), .B2(ADS_N_REG_SCAN_IN), .C1(DATAI_1_), 
        .C2(keyinput_f30), .A(n6597), .ZN(n6602) );
  AOI22_X1 U7538 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_f32), .B1(
        DATAI_22_), .B2(keyinput_f9), .ZN(n6598) );
  OAI221_X1 U7539 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_f32), .C1(
        DATAI_22_), .C2(keyinput_f9), .A(n6598), .ZN(n6601) );
  AOI22_X1 U7540 ( .A1(DATAI_25_), .A2(keyinput_f6), .B1(DATAI_30_), .B2(
        keyinput_f1), .ZN(n6599) );
  OAI221_X1 U7541 ( .B1(DATAI_25_), .B2(keyinput_f6), .C1(DATAI_30_), .C2(
        keyinput_f1), .A(n6599), .ZN(n6600) );
  NOR4_X1 U7542 ( .A1(n6603), .A2(n6602), .A3(n6601), .A4(n6600), .ZN(n6607)
         );
  AOI22_X1 U7543 ( .A1(DATAI_16_), .A2(keyinput_f15), .B1(DATAI_31_), .B2(
        keyinput_f0), .ZN(n6604) );
  OAI221_X1 U7544 ( .B1(DATAI_16_), .B2(keyinput_f15), .C1(DATAI_31_), .C2(
        keyinput_f0), .A(n6604), .ZN(n6605) );
  AOI21_X1 U7545 ( .B1(keyinput_f59), .B2(n6718), .A(n6605), .ZN(n6606) );
  OAI211_X1 U7546 ( .C1(keyinput_f59), .C2(n6718), .A(n6607), .B(n6606), .ZN(
        n6651) );
  AOI22_X1 U7547 ( .A1(DATAI_7_), .A2(keyinput_f24), .B1(DATAI_28_), .B2(
        keyinput_f3), .ZN(n6608) );
  OAI221_X1 U7548 ( .B1(DATAI_7_), .B2(keyinput_f24), .C1(DATAI_28_), .C2(
        keyinput_f3), .A(n6608), .ZN(n6615) );
  AOI22_X1 U7549 ( .A1(DATAI_9_), .A2(keyinput_f22), .B1(REIP_REG_25__SCAN_IN), 
        .B2(keyinput_f57), .ZN(n6609) );
  OAI221_X1 U7550 ( .B1(DATAI_9_), .B2(keyinput_f22), .C1(REIP_REG_25__SCAN_IN), .C2(keyinput_f57), .A(n6609), .ZN(n6614) );
  AOI22_X1 U7551 ( .A1(DATAI_13_), .A2(keyinput_f18), .B1(REIP_REG_29__SCAN_IN), .B2(keyinput_f53), .ZN(n6610) );
  OAI221_X1 U7552 ( .B1(DATAI_13_), .B2(keyinput_f18), .C1(
        REIP_REG_29__SCAN_IN), .C2(keyinput_f53), .A(n6610), .ZN(n6613) );
  AOI22_X1 U7553 ( .A1(DATAI_18_), .A2(keyinput_f13), .B1(DATAI_19_), .B2(
        keyinput_f12), .ZN(n6611) );
  OAI221_X1 U7554 ( .B1(DATAI_18_), .B2(keyinput_f13), .C1(DATAI_19_), .C2(
        keyinput_f12), .A(n6611), .ZN(n6612) );
  NOR4_X1 U7555 ( .A1(n6615), .A2(n6614), .A3(n6613), .A4(n6612), .ZN(n6649)
         );
  AOI22_X1 U7556 ( .A1(DATAI_27_), .A2(keyinput_f4), .B1(REIP_REG_22__SCAN_IN), 
        .B2(keyinput_f60), .ZN(n6616) );
  OAI221_X1 U7557 ( .B1(DATAI_27_), .B2(keyinput_f4), .C1(REIP_REG_22__SCAN_IN), .C2(keyinput_f60), .A(n6616), .ZN(n6623) );
  AOI22_X1 U7558 ( .A1(keyinput_f36), .A2(HOLD), .B1(MORE_REG_SCAN_IN), .B2(
        keyinput_f44), .ZN(n6617) );
  OAI221_X1 U7559 ( .B1(keyinput_f36), .B2(HOLD), .C1(MORE_REG_SCAN_IN), .C2(
        keyinput_f44), .A(n6617), .ZN(n6622) );
  AOI22_X1 U7560 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(keyinput_f39), .B1(
        REIP_REG_31__SCAN_IN), .B2(keyinput_f51), .ZN(n6618) );
  OAI221_X1 U7561 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput_f39), .C1(
        REIP_REG_31__SCAN_IN), .C2(keyinput_f51), .A(n6618), .ZN(n6621) );
  AOI22_X1 U7562 ( .A1(DATAI_20_), .A2(keyinput_f11), .B1(REIP_REG_27__SCAN_IN), .B2(keyinput_f55), .ZN(n6619) );
  OAI221_X1 U7563 ( .B1(DATAI_20_), .B2(keyinput_f11), .C1(
        REIP_REG_27__SCAN_IN), .C2(keyinput_f55), .A(n6619), .ZN(n6620) );
  NOR4_X1 U7564 ( .A1(n6623), .A2(n6622), .A3(n6621), .A4(n6620), .ZN(n6648)
         );
  AOI22_X1 U7565 ( .A1(n6626), .A2(keyinput_f54), .B1(keyinput_f19), .B2(n6625), .ZN(n6624) );
  OAI221_X1 U7566 ( .B1(n6626), .B2(keyinput_f54), .C1(n6625), .C2(
        keyinput_f19), .A(n6624), .ZN(n6636) );
  AOI22_X1 U7567 ( .A1(n6628), .A2(keyinput_f31), .B1(keyinput_f42), .B2(n6715), .ZN(n6627) );
  OAI221_X1 U7568 ( .B1(n6628), .B2(keyinput_f31), .C1(n6715), .C2(
        keyinput_f42), .A(n6627), .ZN(n6635) );
  AOI22_X1 U7569 ( .A1(n6631), .A2(keyinput_f20), .B1(keyinput_f47), .B2(n6630), .ZN(n6629) );
  OAI221_X1 U7570 ( .B1(n6631), .B2(keyinput_f20), .C1(n6630), .C2(
        keyinput_f47), .A(n6629), .ZN(n6634) );
  INV_X1 U7571 ( .A(DATAI_15_), .ZN(n6727) );
  AOI22_X1 U7572 ( .A1(n6721), .A2(keyinput_f29), .B1(keyinput_f16), .B2(n6727), .ZN(n6632) );
  OAI221_X1 U7573 ( .B1(n6721), .B2(keyinput_f29), .C1(n6727), .C2(
        keyinput_f16), .A(n6632), .ZN(n6633) );
  NOR4_X1 U7574 ( .A1(n6636), .A2(n6635), .A3(n6634), .A4(n6633), .ZN(n6647)
         );
  AOI22_X1 U7575 ( .A1(keyinput_f40), .A2(M_IO_N_REG_SCAN_IN), .B1(DATAI_24_), 
        .B2(keyinput_f7), .ZN(n6637) );
  OAI221_X1 U7576 ( .B1(keyinput_f40), .B2(M_IO_N_REG_SCAN_IN), .C1(DATAI_24_), 
        .C2(keyinput_f7), .A(n6637), .ZN(n6645) );
  AOI22_X1 U7577 ( .A1(keyinput_f46), .A2(W_R_N_REG_SCAN_IN), .B1(
        REIP_REG_30__SCAN_IN), .B2(keyinput_f52), .ZN(n6638) );
  OAI221_X1 U7578 ( .B1(keyinput_f46), .B2(W_R_N_REG_SCAN_IN), .C1(
        REIP_REG_30__SCAN_IN), .C2(keyinput_f52), .A(n6638), .ZN(n6644) );
  AOI22_X1 U7579 ( .A1(n6640), .A2(keyinput_f21), .B1(n6756), .B2(keyinput_f62), .ZN(n6639) );
  OAI221_X1 U7580 ( .B1(n6640), .B2(keyinput_f21), .C1(n6756), .C2(
        keyinput_f62), .A(n6639), .ZN(n6643) );
  AOI22_X1 U7581 ( .A1(n6728), .A2(keyinput_f35), .B1(keyinput_f61), .B2(n6734), .ZN(n6641) );
  OAI221_X1 U7582 ( .B1(n6728), .B2(keyinput_f35), .C1(n6734), .C2(
        keyinput_f61), .A(n6641), .ZN(n6642) );
  NOR4_X1 U7583 ( .A1(n6645), .A2(n6644), .A3(n6643), .A4(n6642), .ZN(n6646)
         );
  NAND4_X1 U7584 ( .A1(n6649), .A2(n6648), .A3(n6647), .A4(n6646), .ZN(n6650)
         );
  NOR4_X1 U7585 ( .A1(n6653), .A2(n6652), .A3(n6651), .A4(n6650), .ZN(n6685)
         );
  INV_X1 U7586 ( .A(keyinput_f33), .ZN(n6655) );
  AOI22_X1 U7587 ( .A1(n6656), .A2(keyinput_f43), .B1(NA_N), .B2(n6655), .ZN(
        n6654) );
  OAI221_X1 U7588 ( .B1(n6656), .B2(keyinput_f43), .C1(n6655), .C2(NA_N), .A(
        n6654), .ZN(n6682) );
  AOI22_X1 U7589 ( .A1(n6658), .A2(keyinput_f28), .B1(n4544), .B2(keyinput_f10), .ZN(n6657) );
  OAI221_X1 U7590 ( .B1(n6658), .B2(keyinput_f28), .C1(n4544), .C2(
        keyinput_f10), .A(n6657), .ZN(n6681) );
  XNOR2_X1 U7591 ( .A(n6704), .B(keyinput_f41), .ZN(n6663) );
  AOI22_X1 U7592 ( .A1(n6661), .A2(keyinput_f23), .B1(n6660), .B2(keyinput_f56), .ZN(n6659) );
  OAI221_X1 U7593 ( .B1(n6661), .B2(keyinput_f23), .C1(n6660), .C2(
        keyinput_f56), .A(n6659), .ZN(n6662) );
  AOI211_X1 U7594 ( .C1(n6706), .C2(keyinput_f48), .A(n6663), .B(n6662), .ZN(
        n6664) );
  OAI21_X1 U7595 ( .B1(n6706), .B2(keyinput_f48), .A(n6664), .ZN(n6680) );
  INV_X1 U7596 ( .A(BS16_N), .ZN(n6666) );
  OAI22_X1 U7597 ( .A1(n6104), .A2(keyinput_f17), .B1(n6666), .B2(keyinput_f34), .ZN(n6665) );
  AOI221_X1 U7598 ( .B1(n6104), .B2(keyinput_f17), .C1(keyinput_f34), .C2(
        n6666), .A(n6665), .ZN(n6678) );
  INV_X1 U7599 ( .A(DATAI_17_), .ZN(n6668) );
  OAI22_X1 U7600 ( .A1(n4540), .A2(keyinput_f8), .B1(n6668), .B2(keyinput_f14), 
        .ZN(n6667) );
  AOI221_X1 U7601 ( .B1(n4540), .B2(keyinput_f8), .C1(keyinput_f14), .C2(n6668), .A(n6667), .ZN(n6677) );
  INV_X1 U7602 ( .A(DATAI_26_), .ZN(n6671) );
  OAI22_X1 U7603 ( .A1(n6671), .A2(keyinput_f5), .B1(n6670), .B2(keyinput_f50), 
        .ZN(n6669) );
  AOI221_X1 U7604 ( .B1(n6671), .B2(keyinput_f5), .C1(keyinput_f50), .C2(n6670), .A(n6669), .ZN(n6676) );
  OAI22_X1 U7605 ( .A1(n6674), .A2(keyinput_f45), .B1(n6673), .B2(keyinput_f37), .ZN(n6672) );
  AOI221_X1 U7606 ( .B1(n6674), .B2(keyinput_f45), .C1(keyinput_f37), .C2(
        n6673), .A(n6672), .ZN(n6675) );
  NAND4_X1 U7607 ( .A1(n6678), .A2(n6677), .A3(n6676), .A4(n6675), .ZN(n6679)
         );
  NOR4_X1 U7608 ( .A1(n6682), .A2(n6681), .A3(n6680), .A4(n6679), .ZN(n6684)
         );
  NOR2_X1 U7609 ( .A1(n6787), .A2(keyinput_f26), .ZN(n6683) );
  AOI221_X1 U7610 ( .B1(n6685), .B2(n6684), .C1(keyinput_f26), .C2(n6787), .A(
        n6683), .ZN(n6786) );
  AOI22_X1 U7611 ( .A1(n6688), .A2(keyinput_g33), .B1(n6687), .B2(keyinput_g58), .ZN(n6686) );
  OAI221_X1 U7612 ( .B1(n6688), .B2(keyinput_g33), .C1(n6687), .C2(
        keyinput_g58), .A(n6686), .ZN(n6699) );
  AOI22_X1 U7613 ( .A1(n6691), .A2(keyinput_g51), .B1(keyinput_g57), .B2(n6690), .ZN(n6689) );
  OAI221_X1 U7614 ( .B1(n6691), .B2(keyinput_g51), .C1(n6690), .C2(
        keyinput_g57), .A(n6689), .ZN(n6698) );
  AOI22_X1 U7615 ( .A1(n6104), .A2(keyinput_g17), .B1(keyinput_g6), .B2(n6693), 
        .ZN(n6692) );
  OAI221_X1 U7616 ( .B1(n6104), .B2(keyinput_g17), .C1(n6693), .C2(keyinput_g6), .A(n6692), .ZN(n6697) );
  AOI22_X1 U7617 ( .A1(n6695), .A2(keyinput_g7), .B1(keyinput_g15), .B2(n4547), 
        .ZN(n6694) );
  OAI221_X1 U7618 ( .B1(n6695), .B2(keyinput_g7), .C1(n4547), .C2(keyinput_g15), .A(n6694), .ZN(n6696) );
  NOR4_X1 U7619 ( .A1(n6699), .A2(n6698), .A3(n6697), .A4(n6696), .ZN(n6745)
         );
  AOI22_X1 U7620 ( .A1(DATAI_3_), .A2(keyinput_g28), .B1(DATAI_23_), .B2(
        keyinput_g8), .ZN(n6700) );
  OAI221_X1 U7621 ( .B1(DATAI_3_), .B2(keyinput_g28), .C1(DATAI_23_), .C2(
        keyinput_g8), .A(n6700), .ZN(n6710) );
  AOI22_X1 U7622 ( .A1(DATAI_26_), .A2(keyinput_g5), .B1(DATAI_28_), .B2(
        keyinput_g3), .ZN(n6701) );
  OAI221_X1 U7623 ( .B1(DATAI_26_), .B2(keyinput_g5), .C1(DATAI_28_), .C2(
        keyinput_g3), .A(n6701), .ZN(n6709) );
  AOI22_X1 U7624 ( .A1(n6704), .A2(keyinput_g41), .B1(n6703), .B2(keyinput_g1), 
        .ZN(n6702) );
  OAI221_X1 U7625 ( .B1(n6704), .B2(keyinput_g41), .C1(n6703), .C2(keyinput_g1), .A(n6702), .ZN(n6708) );
  AOI22_X1 U7626 ( .A1(DATAI_4_), .A2(keyinput_g27), .B1(n6706), .B2(
        keyinput_g48), .ZN(n6705) );
  OAI221_X1 U7627 ( .B1(DATAI_4_), .B2(keyinput_g27), .C1(n6706), .C2(
        keyinput_g48), .A(n6705), .ZN(n6707) );
  NOR4_X1 U7628 ( .A1(n6710), .A2(n6709), .A3(n6708), .A4(n6707), .ZN(n6744)
         );
  INV_X1 U7629 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6712) );
  AOI22_X1 U7630 ( .A1(n6713), .A2(keyinput_g39), .B1(keyinput_g40), .B2(n6712), .ZN(n6711) );
  OAI221_X1 U7631 ( .B1(n6713), .B2(keyinput_g39), .C1(n6712), .C2(
        keyinput_g40), .A(n6711), .ZN(n6725) );
  AOI22_X1 U7632 ( .A1(n6716), .A2(keyinput_g38), .B1(n6715), .B2(keyinput_g42), .ZN(n6714) );
  OAI221_X1 U7633 ( .B1(n6716), .B2(keyinput_g38), .C1(n6715), .C2(
        keyinput_g42), .A(n6714), .ZN(n6724) );
  AOI22_X1 U7634 ( .A1(n6718), .A2(keyinput_g59), .B1(keyinput_g13), .B2(n4536), .ZN(n6717) );
  OAI221_X1 U7635 ( .B1(n6718), .B2(keyinput_g59), .C1(n4536), .C2(
        keyinput_g13), .A(n6717), .ZN(n6723) );
  AOI22_X1 U7636 ( .A1(n6721), .A2(keyinput_g29), .B1(n6720), .B2(keyinput_g18), .ZN(n6719) );
  OAI221_X1 U7637 ( .B1(n6721), .B2(keyinput_g29), .C1(n6720), .C2(
        keyinput_g18), .A(n6719), .ZN(n6722) );
  NOR4_X1 U7638 ( .A1(n6725), .A2(n6724), .A3(n6723), .A4(n6722), .ZN(n6743)
         );
  AOI22_X1 U7639 ( .A1(n6728), .A2(keyinput_g35), .B1(keyinput_g16), .B2(n6727), .ZN(n6726) );
  OAI221_X1 U7640 ( .B1(n6728), .B2(keyinput_g35), .C1(n6727), .C2(
        keyinput_g16), .A(n6726), .ZN(n6741) );
  AOI22_X1 U7641 ( .A1(n6731), .A2(keyinput_g36), .B1(n6730), .B2(keyinput_g4), 
        .ZN(n6729) );
  OAI221_X1 U7642 ( .B1(n6731), .B2(keyinput_g36), .C1(n6730), .C2(keyinput_g4), .A(n6729), .ZN(n6740) );
  AOI22_X1 U7643 ( .A1(n6734), .A2(keyinput_g61), .B1(n6733), .B2(keyinput_g53), .ZN(n6732) );
  OAI221_X1 U7644 ( .B1(n6734), .B2(keyinput_g61), .C1(n6733), .C2(
        keyinput_g53), .A(n6732), .ZN(n6739) );
  AOI22_X1 U7645 ( .A1(n6737), .A2(keyinput_g30), .B1(n6736), .B2(keyinput_g2), 
        .ZN(n6735) );
  OAI221_X1 U7646 ( .B1(n6737), .B2(keyinput_g30), .C1(n6736), .C2(keyinput_g2), .A(n6735), .ZN(n6738) );
  NOR4_X1 U7647 ( .A1(n6741), .A2(n6740), .A3(n6739), .A4(n6738), .ZN(n6742)
         );
  NAND4_X1 U7648 ( .A1(n6745), .A2(n6744), .A3(n6743), .A4(n6742), .ZN(n6784)
         );
  AOI22_X1 U7649 ( .A1(FLUSH_REG_SCAN_IN), .A2(keyinput_g45), .B1(
        REIP_REG_22__SCAN_IN), .B2(keyinput_g60), .ZN(n6746) );
  OAI221_X1 U7650 ( .B1(FLUSH_REG_SCAN_IN), .B2(keyinput_g45), .C1(
        REIP_REG_22__SCAN_IN), .C2(keyinput_g60), .A(n6746), .ZN(n6753) );
  AOI22_X1 U7651 ( .A1(DATAI_20_), .A2(keyinput_g11), .B1(DATAI_31_), .B2(
        keyinput_g0), .ZN(n6747) );
  OAI221_X1 U7652 ( .B1(DATAI_20_), .B2(keyinput_g11), .C1(DATAI_31_), .C2(
        keyinput_g0), .A(n6747), .ZN(n6752) );
  AOI22_X1 U7653 ( .A1(MORE_REG_SCAN_IN), .A2(keyinput_g44), .B1(
        REIP_REG_26__SCAN_IN), .B2(keyinput_g56), .ZN(n6748) );
  OAI221_X1 U7654 ( .B1(MORE_REG_SCAN_IN), .B2(keyinput_g44), .C1(
        REIP_REG_26__SCAN_IN), .C2(keyinput_g56), .A(n6748), .ZN(n6751) );
  AOI22_X1 U7655 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_g32), .B1(
        DATAI_0_), .B2(keyinput_g31), .ZN(n6749) );
  OAI221_X1 U7656 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_g32), .C1(
        DATAI_0_), .C2(keyinput_g31), .A(n6749), .ZN(n6750) );
  NOR4_X1 U7657 ( .A1(n6753), .A2(n6752), .A3(n6751), .A4(n6750), .ZN(n6782)
         );
  XOR2_X1 U7658 ( .A(n6754), .B(keyinput_g49), .Z(n6762) );
  AOI22_X1 U7659 ( .A1(BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput_g47), .B1(
        n6756), .B2(keyinput_g62), .ZN(n6755) );
  OAI221_X1 U7660 ( .B1(BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_g47), .C1(
        n6756), .C2(keyinput_g62), .A(n6755), .ZN(n6761) );
  AOI22_X1 U7661 ( .A1(DATAI_7_), .A2(keyinput_g24), .B1(DATAI_10_), .B2(
        keyinput_g21), .ZN(n6757) );
  OAI221_X1 U7662 ( .B1(DATAI_7_), .B2(keyinput_g24), .C1(DATAI_10_), .C2(
        keyinput_g21), .A(n6757), .ZN(n6760) );
  AOI22_X1 U7663 ( .A1(DATAI_6_), .A2(keyinput_g25), .B1(DATAI_9_), .B2(
        keyinput_g22), .ZN(n6758) );
  OAI221_X1 U7664 ( .B1(DATAI_6_), .B2(keyinput_g25), .C1(DATAI_9_), .C2(
        keyinput_g22), .A(n6758), .ZN(n6759) );
  NOR4_X1 U7665 ( .A1(n6762), .A2(n6761), .A3(n6760), .A4(n6759), .ZN(n6781)
         );
  AOI22_X1 U7666 ( .A1(BS16_N), .A2(keyinput_g34), .B1(REIP_REG_30__SCAN_IN), 
        .B2(keyinput_g52), .ZN(n6763) );
  OAI221_X1 U7667 ( .B1(BS16_N), .B2(keyinput_g34), .C1(REIP_REG_30__SCAN_IN), 
        .C2(keyinput_g52), .A(n6763), .ZN(n6770) );
  AOI22_X1 U7668 ( .A1(REIP_REG_19__SCAN_IN), .A2(keyinput_g63), .B1(
        STATEBS16_REG_SCAN_IN), .B2(keyinput_g43), .ZN(n6764) );
  OAI221_X1 U7669 ( .B1(REIP_REG_19__SCAN_IN), .B2(keyinput_g63), .C1(
        STATEBS16_REG_SCAN_IN), .C2(keyinput_g43), .A(n6764), .ZN(n6769) );
  AOI22_X1 U7670 ( .A1(W_R_N_REG_SCAN_IN), .A2(keyinput_g46), .B1(DATAI_17_), 
        .B2(keyinput_g14), .ZN(n6765) );
  OAI221_X1 U7671 ( .B1(W_R_N_REG_SCAN_IN), .B2(keyinput_g46), .C1(DATAI_17_), 
        .C2(keyinput_g14), .A(n6765), .ZN(n6768) );
  AOI22_X1 U7672 ( .A1(DATAI_22_), .A2(keyinput_g9), .B1(DATAI_11_), .B2(
        keyinput_g20), .ZN(n6766) );
  OAI221_X1 U7673 ( .B1(DATAI_22_), .B2(keyinput_g9), .C1(DATAI_11_), .C2(
        keyinput_g20), .A(n6766), .ZN(n6767) );
  NOR4_X1 U7674 ( .A1(n6770), .A2(n6769), .A3(n6768), .A4(n6767), .ZN(n6780)
         );
  AOI22_X1 U7675 ( .A1(DATAI_8_), .A2(keyinput_g23), .B1(REIP_REG_27__SCAN_IN), 
        .B2(keyinput_g55), .ZN(n6771) );
  OAI221_X1 U7676 ( .B1(DATAI_8_), .B2(keyinput_g23), .C1(REIP_REG_27__SCAN_IN), .C2(keyinput_g55), .A(n6771), .ZN(n6778) );
  AOI22_X1 U7677 ( .A1(DATAI_19_), .A2(keyinput_g12), .B1(REIP_REG_28__SCAN_IN), .B2(keyinput_g54), .ZN(n6772) );
  OAI221_X1 U7678 ( .B1(DATAI_19_), .B2(keyinput_g12), .C1(
        REIP_REG_28__SCAN_IN), .C2(keyinput_g54), .A(n6772), .ZN(n6777) );
  AOI22_X1 U7679 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_g50), .B1(
        READREQUEST_REG_SCAN_IN), .B2(keyinput_g37), .ZN(n6773) );
  OAI221_X1 U7680 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_g50), .C1(
        READREQUEST_REG_SCAN_IN), .C2(keyinput_g37), .A(n6773), .ZN(n6776) );
  AOI22_X1 U7681 ( .A1(DATAI_21_), .A2(keyinput_g10), .B1(DATAI_12_), .B2(
        keyinput_g19), .ZN(n6774) );
  OAI221_X1 U7682 ( .B1(DATAI_21_), .B2(keyinput_g10), .C1(DATAI_12_), .C2(
        keyinput_g19), .A(n6774), .ZN(n6775) );
  NOR4_X1 U7683 ( .A1(n6778), .A2(n6777), .A3(n6776), .A4(n6775), .ZN(n6779)
         );
  NAND4_X1 U7684 ( .A1(n6782), .A2(n6781), .A3(n6780), .A4(n6779), .ZN(n6783)
         );
  OAI22_X1 U7685 ( .A1(keyinput_g26), .A2(n6787), .B1(n6784), .B2(n6783), .ZN(
        n6785) );
  AOI211_X1 U7686 ( .C1(keyinput_g26), .C2(n6787), .A(n6786), .B(n6785), .ZN(
        n6791) );
  AOI22_X1 U7687 ( .A1(n6789), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n6788), .ZN(n6790) );
  XNOR2_X1 U7688 ( .A(n6791), .B(n6790), .ZN(U3445) );
  XNOR2_X1 U3476 ( .A(n3399), .B(n4503), .ZN(n3629) );
  XNOR2_X1 U3610 ( .A(n3769), .B(n3770), .ZN(n5214) );
  CLKBUF_X1 U34480 ( .A(n3406), .Z(n2988) );
  CLKBUF_X2 U3458 ( .A(n3201), .Z(n3016) );
  CLKBUF_X1 U34620 ( .A(n3170), .Z(n3546) );
  NAND2_X1 U3467 ( .A1(n3355), .A2(n3427), .ZN(n3399) );
  AND2_X2 U3477 ( .A1(n5439), .A2(n5441), .ZN(n2984) );
  CLKBUF_X1 U3484 ( .A(n6066), .Z(n6062) );
  CLKBUF_X1 U3724 ( .A(n3234), .Z(n5343) );
endmodule

