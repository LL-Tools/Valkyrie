

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput63, keyinput62, keyinput61, 
        keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, 
        keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, 
        keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, 
        keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, 
        keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, 
        keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, 
        keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, 
        keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, 
        keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, 
        keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, 
        keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput63, keyinput62,
         keyinput61, keyinput60, keyinput59, keyinput58, keyinput57,
         keyinput56, keyinput55, keyinput54, keyinput53, keyinput52,
         keyinput51, keyinput50, keyinput49, keyinput48, keyinput47,
         keyinput46, keyinput45, keyinput44, keyinput43, keyinput42,
         keyinput41, keyinput40, keyinput39, keyinput38, keyinput37,
         keyinput36, keyinput35, keyinput34, keyinput33, keyinput32,
         keyinput31, keyinput30, keyinput29, keyinput28, keyinput27,
         keyinput26, keyinput25, keyinput24, keyinput23, keyinput22,
         keyinput21, keyinput20, keyinput19, keyinput18, keyinput17,
         keyinput16, keyinput15, keyinput14, keyinput13, keyinput12,
         keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6,
         keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2952, n2953, n2954, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614;

  NAND2_X1 U3400 ( .A1(n3877), .A2(n4162), .ZN(n5013) );
  INV_X2 U3401 ( .A(n5292), .ZN(n5298) );
  OAI21_X1 U3402 ( .B1(n3328), .B2(n3327), .A(n3329), .ZN(n3323) );
  CLKBUF_X2 U3403 ( .A(n3274), .Z(n2953) );
  CLKBUF_X2 U3404 ( .A(n3249), .Z(n3855) );
  CLKBUF_X1 U3405 ( .A(n3198), .Z(n4527) );
  CLKBUF_X2 U3406 ( .A(n3128), .Z(n2976) );
  AND2_X1 U3407 ( .A1(n4425), .A2(n4416), .ZN(n3249) );
  AND2_X2 U3408 ( .A1(n4975), .A2(n4416), .ZN(n3128) );
  AND2_X2 U3409 ( .A1(n4974), .A2(n4416), .ZN(n3273) );
  CLKBUF_X3 U3410 ( .A(n3128), .Z(n2975) );
  AND4_X1 U3411 ( .A1(n3093), .A2(n3092), .A3(n3091), .A4(n3090), .ZN(n3094)
         );
  NAND2_X1 U3412 ( .A1(n3323), .A2(n3322), .ZN(n3374) );
  NAND2_X1 U3413 ( .A1(n3880), .A2(n4715), .ZN(n4030) );
  BUF_X1 U3415 ( .A(n3944), .Z(n4517) );
  INV_X1 U3416 ( .A(n5292), .ZN(n5808) );
  INV_X1 U3417 ( .A(n3951), .ZN(n4236) );
  OR2_X2 U3418 ( .A1(n3105), .A2(n3104), .ZN(n4501) );
  NAND2_X1 U3419 ( .A1(n2969), .A2(n4396), .ZN(n4395) );
  AND2_X1 U3420 ( .A1(n4666), .A2(n4667), .ZN(n4665) );
  INV_X1 U3421 ( .A(n5745), .ZN(n5717) );
  INV_X1 U3422 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3063) );
  OR2_X1 U3423 ( .A1(n4419), .A2(n4288), .ZN(n2952) );
  NAND2_X2 U3424 ( .A1(n3240), .A2(n3239), .ZN(n3353) );
  AND2_X4 U3425 ( .A1(n3068), .A2(n4457), .ZN(n3280) );
  NAND2_X4 U3426 ( .A1(n3085), .A2(n3084), .ZN(n3178) );
  AND4_X2 U3427 ( .A1(n3089), .A2(n3088), .A3(n3087), .A4(n3086), .ZN(n3095)
         );
  XNOR2_X2 U3428 ( .A(n4083), .B(n5903), .ZN(n4737) );
  NAND2_X2 U3429 ( .A1(n3011), .A2(n4082), .ZN(n4083) );
  XNOR2_X1 U3430 ( .A(n4227), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5050)
         );
  AOI21_X1 U3431 ( .B1(n3023), .B2(n3019), .A(n3017), .ZN(n3016) );
  NAND2_X1 U3432 ( .A1(n3444), .A2(n3443), .ZN(n4122) );
  AOI21_X1 U3433 ( .B1(n4367), .B2(n4368), .A(n4071), .ZN(n5833) );
  NAND2_X1 U3434 ( .A1(n3372), .A2(n3371), .ZN(n4470) );
  NAND2_X1 U3436 ( .A1(n3181), .A2(n4249), .ZN(n4420) );
  NOR2_X2 U3437 ( .A1(n3951), .A2(n3969), .ZN(n3961) );
  BUF_X4 U3438 ( .A(n3224), .Z(n2954) );
  INV_X2 U3439 ( .A(n4715), .ZN(n3192) );
  AND2_X2 U3440 ( .A1(n3075), .A2(n3074), .ZN(n3176) );
  BUF_X2 U3441 ( .A(n3273), .Z(n3821) );
  CLKBUF_X2 U3442 ( .A(n3152), .Z(n3833) );
  BUF_X2 U3443 ( .A(n3272), .Z(n3822) );
  CLKBUF_X2 U3444 ( .A(n3244), .Z(n3731) );
  BUF_X2 U34450 ( .A(n3157), .Z(n3820) );
  CLKBUF_X2 U34460 ( .A(n3304), .Z(n3860) );
  CLKBUF_X2 U34470 ( .A(n3275), .Z(n3861) );
  BUF_X2 U34480 ( .A(n3298), .Z(n3750) );
  OR2_X1 U3449 ( .A1(n4157), .A2(n4156), .ZN(n5032) );
  NAND2_X1 U3450 ( .A1(n5312), .A2(n5313), .ZN(n5311) );
  NAND2_X1 U34510 ( .A1(n3031), .A2(n3034), .ZN(n5279) );
  NAND2_X1 U34520 ( .A1(n5287), .A2(n4143), .ZN(n4144) );
  CLKBUF_X1 U34530 ( .A(n2965), .Z(n2963) );
  AOI21_X1 U3454 ( .B1(n3016), .B2(n3018), .A(n2983), .ZN(n3014) );
  NAND2_X1 U34550 ( .A1(n4665), .A2(n3040), .ZN(n4861) );
  AOI21_X1 U34560 ( .B1(n3028), .B2(n3030), .A(n3027), .ZN(n3026) );
  NOR2_X1 U3457 ( .A1(n3021), .A2(n4944), .ZN(n3020) );
  AND2_X1 U3458 ( .A1(n4666), .A2(n4667), .ZN(n2967) );
  OR2_X1 U34590 ( .A1(n5062), .A2(n5887), .ZN(n5058) );
  XNOR2_X1 U34600 ( .A(n4122), .B(n3447), .ZN(n4111) );
  NAND2_X1 U34610 ( .A1(n4122), .A2(n4121), .ZN(n4130) );
  NAND2_X1 U34620 ( .A1(n3350), .A2(n3349), .ZN(n4397) );
  XNOR2_X1 U34630 ( .A(n3416), .B(n3420), .ZN(n4093) );
  NAND2_X1 U34640 ( .A1(n3341), .A2(n3340), .ZN(n6143) );
  NAND2_X1 U34650 ( .A1(n5248), .A2(n4321), .ZN(n5534) );
  AND2_X1 U3466 ( .A1(n3321), .A2(n3337), .ZN(n3329) );
  NAND2_X1 U3467 ( .A1(n3039), .A2(n2984), .ZN(n3258) );
  NOR2_X1 U34680 ( .A1(n4518), .A2(n4894), .ZN(n6238) );
  NAND2_X2 U34690 ( .A1(n4244), .A2(n4249), .ZN(n4323) );
  AND2_X2 U34710 ( .A1(n5817), .A2(n4166), .ZN(n5823) );
  NAND2_X1 U34720 ( .A1(n3358), .A2(n3357), .ZN(n6103) );
  NAND2_X1 U34730 ( .A1(n3292), .A2(n3291), .ZN(n3296) );
  CLKBUF_X1 U34740 ( .A(n3234), .Z(n2959) );
  OAI211_X1 U3475 ( .C1(n4177), .C2(n3182), .A(n2952), .B(n4420), .ZN(n3183)
         );
  NAND2_X1 U3476 ( .A1(n3207), .A2(n3206), .ZN(n3234) );
  AND2_X1 U3477 ( .A1(n3219), .A2(n3218), .ZN(n3888) );
  INV_X1 U3478 ( .A(n4179), .ZN(n3181) );
  NOR2_X1 U3479 ( .A1(n3879), .A2(n3054), .ZN(n3203) );
  AND2_X1 U3480 ( .A1(n3196), .A2(n3195), .ZN(n3228) );
  NAND2_X1 U3481 ( .A1(n3190), .A2(n4290), .ZN(n3879) );
  INV_X2 U3482 ( .A(n3176), .ZN(n3193) );
  OR2_X1 U3483 ( .A1(n3944), .A2(n4198), .ZN(n3191) );
  OR2_X1 U3484 ( .A1(n3286), .A2(n3285), .ZN(n4123) );
  OR2_X1 U3485 ( .A1(n3270), .A2(n3269), .ZN(n4064) );
  NAND4_X2 U3486 ( .A1(n3174), .A2(n3173), .A3(n3172), .A4(n3171), .ZN(n3944)
         );
  AND4_X1 U3487 ( .A1(n3156), .A2(n3155), .A3(n3154), .A4(n3153), .ZN(n3174)
         );
  AND4_X1 U3488 ( .A1(n3132), .A2(n3131), .A3(n3130), .A4(n3129), .ZN(n3150)
         );
  AND4_X1 U3489 ( .A1(n3110), .A2(n3109), .A3(n3108), .A4(n3107), .ZN(n3115)
         );
  AND4_X1 U3490 ( .A1(n3073), .A2(n3072), .A3(n3071), .A4(n3070), .ZN(n3074)
         );
  AND4_X1 U3491 ( .A1(n3162), .A2(n3161), .A3(n3160), .A4(n3159), .ZN(n3173)
         );
  AND4_X1 U3492 ( .A1(n3146), .A2(n3145), .A3(n3144), .A4(n3143), .ZN(n3147)
         );
  AND4_X1 U3493 ( .A1(n3136), .A2(n3135), .A3(n3134), .A4(n3133), .ZN(n3149)
         );
  AND4_X1 U3494 ( .A1(n3067), .A2(n3066), .A3(n3065), .A4(n3064), .ZN(n3075)
         );
  AND4_X1 U3495 ( .A1(n3083), .A2(n3082), .A3(n3081), .A4(n3080), .ZN(n3084)
         );
  AND4_X1 U3496 ( .A1(n3166), .A2(n3165), .A3(n3164), .A4(n3163), .ZN(n3172)
         );
  INV_X2 U3497 ( .A(n6440), .ZN(n4387) );
  BUF_X4 U3498 ( .A(n3815), .Z(n2972) );
  AND2_X2 U3499 ( .A1(n4974), .A2(n3068), .ZN(n3274) );
  AND2_X2 U3500 ( .A1(n3068), .A2(n4425), .ZN(n3244) );
  AND2_X2 U3501 ( .A1(n4425), .A2(n3069), .ZN(n3298) );
  BUF_X4 U3502 ( .A(n3815), .Z(n2973) );
  AND2_X2 U3503 ( .A1(n3063), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3068)
         );
  AND2_X2 U3504 ( .A1(n3062), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4974)
         );
  AND2_X2 U3505 ( .A1(n3038), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4975)
         );
  AND2_X2 U3506 ( .A1(n4457), .A2(n4426), .ZN(n3815) );
  NOR2_X2 U3507 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4426) );
  AND2_X2 U3508 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4425) );
  CLKBUF_X1 U3510 ( .A(n4405), .Z(n2956) );
  NOR2_X2 U3512 ( .A1(n4395), .A2(n4486), .ZN(n4405) );
  NAND3_X1 U3513 ( .A1(n4405), .A2(n4404), .A3(n3440), .ZN(n4614) );
  CLKBUF_X1 U3514 ( .A(n5824), .Z(n2958) );
  OAI21_X2 U3517 ( .B1(n5348), .B2(n4136), .A(n4135), .ZN(n2962) );
  NAND2_X1 U3518 ( .A1(n3013), .A2(n3014), .ZN(n5348) );
  OAI21_X1 U3519 ( .B1(n5348), .B2(n4136), .A(n4135), .ZN(n5341) );
  OAI21_X1 U3520 ( .B1(n2962), .B2(n4138), .A(n4137), .ZN(n2965) );
  NAND2_X1 U3521 ( .A1(n5287), .A2(n4143), .ZN(n2964) );
  OR2_X1 U3522 ( .A1(n2964), .A2(n3036), .ZN(n3031) );
  OAI21_X1 U3523 ( .B1(n5341), .B2(n4138), .A(n4137), .ZN(n5333) );
  OR2_X1 U3524 ( .A1(n2965), .A2(n4140), .ZN(n2966) );
  AND3_X1 U3525 ( .A1(n3187), .A2(n4715), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3905) );
  AND2_X1 U3526 ( .A1(n3904), .A2(n3194), .ZN(n3216) );
  AND2_X2 U3527 ( .A1(n2967), .A2(n2968), .ZN(n3534) );
  AND2_X1 U3528 ( .A1(n3528), .A2(n3040), .ZN(n2968) );
  AOI21_X1 U3529 ( .B1(n4077), .B2(n3574), .A(n3381), .ZN(n3382) );
  AND2_X2 U3530 ( .A1(n3351), .A2(n4397), .ZN(n2969) );
  AND2_X1 U3531 ( .A1(n3193), .A2(n3944), .ZN(n3904) );
  XNOR2_X1 U3532 ( .A(n3330), .B(n3329), .ZN(n4471) );
  AOI21_X2 U3533 ( .B1(n5321), .B2(n5320), .A(n5290), .ZN(n5312) );
  XNOR2_X1 U3534 ( .A(n3353), .B(n6103), .ZN(n4417) );
  OR2_X2 U3535 ( .A1(n3210), .A2(n3186), .ZN(n2982) );
  AND2_X2 U3536 ( .A1(n3012), .A2(n3403), .ZN(n4077) );
  OR2_X1 U3537 ( .A1(n3217), .A2(n3216), .ZN(n3219) );
  OAI22_X2 U3538 ( .A1(n5299), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5306), .B2(n5293), .ZN(n5294) );
  OAI21_X2 U3539 ( .B1(n5292), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5311), 
        .ZN(n5306) );
  NAND2_X4 U3540 ( .A1(n3095), .A2(n3094), .ZN(n3187) );
  NAND2_X1 U3541 ( .A1(n3176), .A2(n3178), .ZN(n3943) );
  NOR2_X2 U3542 ( .A1(n4614), .A2(n4615), .ZN(n4666) );
  AND2_X2 U3543 ( .A1(n5085), .A2(n3052), .ZN(n4160) );
  NOR2_X2 U3544 ( .A1(n5133), .A2(n5134), .ZN(n5135) );
  OR2_X1 U3545 ( .A1(n5146), .A2(n5155), .ZN(n5487) );
  NOR2_X2 U3546 ( .A1(n5112), .A2(n3044), .ZN(n5146) );
  NOR2_X2 U3547 ( .A1(n5185), .A2(n5187), .ZN(n5178) );
  AND2_X4 U3548 ( .A1(n4975), .A2(n3068), .ZN(n3137) );
  AND2_X2 U3549 ( .A1(n4457), .A2(n4416), .ZN(n2978) );
  AND2_X1 U3550 ( .A1(n4457), .A2(n4416), .ZN(n3158) );
  AND2_X1 U3552 ( .A1(n4457), .A2(n4416), .ZN(n2977) );
  CLKBUF_X1 U3553 ( .A(n4245), .Z(n4246) );
  AND2_X1 U3554 ( .A1(n4466), .A2(n6332), .ZN(n4291) );
  NAND2_X1 U3555 ( .A1(n3905), .A2(n2970), .ZN(n3939) );
  NOR2_X2 U3556 ( .A1(n3944), .A2(n4715), .ZN(n4749) );
  NAND3_X1 U3557 ( .A1(n4437), .A2(n4291), .A3(n6345), .ZN(n4317) );
  OR2_X1 U3558 ( .A1(n5115), .A2(n5170), .ZN(n3009) );
  AOI21_X1 U3559 ( .B1(n3020), .B2(n3055), .A(n2989), .ZN(n3019) );
  INV_X1 U3560 ( .A(n4133), .ZN(n3021) );
  INV_X1 U3561 ( .A(n4944), .ZN(n3024) );
  NAND2_X1 U3562 ( .A1(n4294), .A2(n4293), .ZN(n4307) );
  INV_X1 U3563 ( .A(n4501), .ZN(n5228) );
  OAI211_X1 U3564 ( .C1(n3178), .C2(n3194), .A(n4290), .B(n3943), .ZN(n3179)
         );
  INV_X1 U3565 ( .A(n3178), .ZN(n3180) );
  NAND2_X1 U3566 ( .A1(n3423), .A2(n3422), .ZN(n3441) );
  AND2_X1 U3567 ( .A1(n3421), .A2(n3420), .ZN(n3422) );
  OR2_X1 U3568 ( .A1(n3903), .A2(n4183), .ZN(n3930) );
  NAND2_X1 U3569 ( .A1(n4501), .A2(n3180), .ZN(n3197) );
  OR2_X1 U3570 ( .A1(n3370), .A2(n3369), .ZN(n4086) );
  NAND2_X1 U3571 ( .A1(n2986), .A2(n3047), .ZN(n3046) );
  INV_X1 U3572 ( .A(n5160), .ZN(n3047) );
  NOR2_X1 U3573 ( .A1(n4976), .A2(n3297), .ZN(n3847) );
  AND2_X1 U3574 ( .A1(n3042), .A2(n3041), .ZN(n3040) );
  INV_X1 U3575 ( .A(n4862), .ZN(n3041) );
  NAND2_X1 U3576 ( .A1(n3033), .A2(n2990), .ZN(n4224) );
  NAND2_X1 U3577 ( .A1(n3036), .A2(n3034), .ZN(n3032) );
  NOR2_X1 U3578 ( .A1(n4732), .A2(n3002), .ZN(n3001) );
  INV_X1 U3579 ( .A(n4671), .ZN(n3002) );
  OR2_X1 U3580 ( .A1(n4030), .A2(n4236), .ZN(n4009) );
  NAND2_X1 U3581 ( .A1(n4236), .A2(n3969), .ZN(n4035) );
  INV_X1 U3582 ( .A(n3198), .ZN(n4290) );
  NAND2_X1 U3583 ( .A1(n3314), .A2(n3313), .ZN(n3335) );
  NAND2_X1 U3584 ( .A1(n3312), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3313) );
  NAND2_X1 U3585 ( .A1(n3342), .A2(n3297), .ZN(n3314) );
  INV_X1 U3586 ( .A(n3905), .ZN(n3931) );
  OAI21_X2 U3587 ( .B1(n4496), .B2(STATE2_REG_0__SCAN_IN), .A(n3271), .ZN(
        n3328) );
  CLKBUF_X1 U3588 ( .A(n4179), .Z(n4278) );
  OAI21_X1 U3589 ( .B1(n6445), .B2(n4479), .A(n6415), .ZN(n4500) );
  NAND2_X1 U3590 ( .A1(n5735), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4754) );
  NAND2_X1 U3591 ( .A1(n4030), .A2(n3969), .ZN(n4303) );
  NAND2_X1 U3592 ( .A1(n4314), .A2(n4313), .ZN(n4436) );
  OR2_X1 U3593 ( .A1(n4423), .A2(n4311), .ZN(n4314) );
  INV_X1 U3594 ( .A(n3745), .ZN(n4173) );
  NOR2_X1 U3595 ( .A1(n3852), .A2(n4169), .ZN(n4188) );
  AND2_X1 U3596 ( .A1(n5085), .A2(n3049), .ZN(n4176) );
  AND2_X1 U3597 ( .A1(n3051), .A2(n3050), .ZN(n3049) );
  INV_X1 U3598 ( .A(n3878), .ZN(n3050) );
  NAND2_X1 U3599 ( .A1(n3772), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3807)
         );
  NOR2_X1 U3600 ( .A1(n3511), .A2(n5670), .ZN(n3529) );
  AND2_X1 U3601 ( .A1(n3436), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3462)
         );
  NOR2_X1 U3602 ( .A1(n5157), .A2(n5149), .ZN(n5151) );
  NOR3_X1 U3603 ( .A1(n5116), .A2(n3010), .A3(n3009), .ZN(n5165) );
  AND2_X1 U3604 ( .A1(n4022), .A2(n4021), .ZN(n5170) );
  NOR3_X1 U3605 ( .A1(n5223), .A2(n3005), .A3(n3003), .ZN(n5180) );
  OR2_X1 U3606 ( .A1(n5125), .A2(n3004), .ZN(n3003) );
  INV_X1 U3607 ( .A(n5192), .ZN(n3004) );
  NAND2_X1 U3608 ( .A1(n5292), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4132) );
  INV_X1 U3609 ( .A(n4866), .ZN(n3027) );
  NAND2_X1 U3610 ( .A1(n4794), .A2(n4793), .ZN(n4792) );
  AND2_X1 U3611 ( .A1(n5463), .A2(n4961), .ZN(n5878) );
  OR2_X1 U3612 ( .A1(n4424), .A2(n4300), .ZN(n4996) );
  NAND2_X1 U3613 ( .A1(n3941), .A2(n3940), .ZN(n4466) );
  OR2_X1 U3614 ( .A1(n3939), .A2(n4185), .ZN(n3940) );
  INV_X1 U3615 ( .A(n6143), .ZN(n6101) );
  NAND2_X1 U3616 ( .A1(n4472), .A2(n6101), .ZN(n6064) );
  NAND2_X1 U3617 ( .A1(n3297), .A2(n4500), .ZN(n4894) );
  AND2_X1 U3618 ( .A1(n6538), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3948) );
  INV_X1 U3619 ( .A(n5741), .ZN(n5746) );
  NAND2_X1 U3620 ( .A1(n6452), .A2(n4187), .ZN(n5735) );
  AND3_X1 U3621 ( .A1(n6328), .A2(n6336), .A3(n5885), .ZN(n4187) );
  NAND2_X1 U3622 ( .A1(n5763), .A2(n4501), .ZN(n5759) );
  AND2_X1 U3623 ( .A1(n5248), .A2(n5019), .ZN(n5770) );
  AND2_X1 U3624 ( .A1(n5248), .A2(n5020), .ZN(n5774) );
  INV_X1 U3625 ( .A(n5248), .ZN(n5773) );
  NAND2_X1 U3626 ( .A1(n5248), .A2(n4322), .ZN(n5249) );
  INV_X1 U3627 ( .A(n5840), .ZN(n5558) );
  INV_X1 U3628 ( .A(n5823), .ZN(n5323) );
  NAND2_X1 U3629 ( .A1(n4307), .A2(n4302), .ZN(n5887) );
  INV_X1 U3630 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6311) );
  INV_X1 U3631 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6538) );
  OR2_X1 U3632 ( .A1(n5991), .A2(n6064), .ZN(n6063) );
  INV_X1 U3633 ( .A(n3403), .ZN(n3423) );
  OR2_X1 U3634 ( .A1(n3413), .A2(n3412), .ZN(n4103) );
  OR2_X1 U3635 ( .A1(n3433), .A2(n3432), .ZN(n4113) );
  OR2_X1 U3636 ( .A1(n3392), .A2(n3391), .ZN(n4102) );
  AND2_X1 U3637 ( .A1(n4501), .A2(n3188), .ZN(n3189) );
  NAND2_X1 U3638 ( .A1(n3106), .A2(n4501), .ZN(n3882) );
  OR2_X1 U3639 ( .A1(n3187), .A2(n3297), .ZN(n3359) );
  AOI22_X1 U3640 ( .A1(n3304), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3142), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3120) );
  OAI21_X1 U3641 ( .B1(n3225), .B2(n3199), .A(n4527), .ZN(n3200) );
  NOR2_X1 U3642 ( .A1(n4418), .A2(n3889), .ZN(n4298) );
  AOI22_X1 U3643 ( .A1(n3272), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3067) );
  AOI22_X1 U3644 ( .A1(n3274), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3072) );
  AOI22_X1 U3645 ( .A1(n3152), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3128), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3071) );
  AND2_X1 U3646 ( .A1(n3052), .A2(n4161), .ZN(n3051) );
  NOR2_X1 U3647 ( .A1(n5075), .A2(n3053), .ZN(n3052) );
  INV_X1 U3648 ( .A(n5087), .ZN(n3053) );
  NOR2_X1 U3649 ( .A1(n4777), .A2(n3043), .ZN(n3042) );
  INV_X1 U3650 ( .A(n4678), .ZN(n3043) );
  XNOR2_X1 U3651 ( .A(n3403), .B(n3421), .ZN(n4085) );
  OAI211_X1 U3652 ( .C1(n3397), .C2(n3063), .A(n3326), .B(n3325), .ZN(n3348)
         );
  NOR2_X1 U3653 ( .A1(n5105), .A2(n5090), .ZN(n2995) );
  NOR2_X1 U3654 ( .A1(n5808), .A2(n3037), .ZN(n3036) );
  NOR2_X1 U3655 ( .A1(n4145), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3037)
         );
  NAND2_X1 U3656 ( .A1(n5808), .A2(n3035), .ZN(n3034) );
  INV_X1 U3657 ( .A(n5001), .ZN(n3035) );
  OR2_X1 U3658 ( .A1(n3006), .A2(n5138), .ZN(n3005) );
  INV_X1 U3659 ( .A(n5561), .ZN(n3017) );
  INV_X1 U3660 ( .A(n3019), .ZN(n3018) );
  INV_X1 U3661 ( .A(n4128), .ZN(n3030) );
  INV_X1 U3662 ( .A(n3029), .ZN(n3028) );
  OAI21_X1 U3663 ( .B1(n4793), .B2(n3030), .A(n4865), .ZN(n3029) );
  INV_X1 U3664 ( .A(n4413), .ZN(n2996) );
  NOR2_X1 U3665 ( .A1(n4401), .A2(n2999), .ZN(n2998) );
  INV_X1 U3666 ( .A(n4490), .ZN(n2999) );
  INV_X1 U3667 ( .A(n4410), .ZN(n2997) );
  NAND2_X1 U3668 ( .A1(n4077), .A2(n2970), .ZN(n3011) );
  NAND2_X1 U3669 ( .A1(n3178), .A2(n4501), .ZN(n4288) );
  INV_X1 U3670 ( .A(n3938), .ZN(n4185) );
  NAND2_X1 U3671 ( .A1(n3360), .A2(n3359), .ZN(n3919) );
  AND2_X1 U3672 ( .A1(n3897), .A2(n3901), .ZN(n3938) );
  OR2_X1 U3673 ( .A1(n3902), .A2(n3896), .ZN(n3897) );
  AND2_X1 U3674 ( .A1(n6311), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3896)
         );
  AND2_X1 U3675 ( .A1(n3931), .A2(n3930), .ZN(n3932) );
  AOI21_X1 U3676 ( .B1(n2959), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3238), 
        .ZN(n3241) );
  INV_X1 U3677 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U3678 ( .A1(n3157), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3132) );
  AOI22_X1 U3679 ( .A1(n3128), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3274), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3092) );
  AOI22_X1 U3680 ( .A1(n2974), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3274), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3098) );
  AOI22_X1 U3681 ( .A1(n3137), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3099) );
  INV_X1 U3682 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6305) );
  NOR2_X1 U3683 ( .A1(n5627), .A2(n4202), .ZN(n5494) );
  INV_X1 U3684 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5670) );
  INV_X1 U3685 ( .A(n5711), .ZN(n5734) );
  OAI22_X1 U3686 ( .A1(n2980), .A2(n5181), .B1(n5014), .B2(n5078), .ZN(n5018)
         );
  NOR2_X1 U3687 ( .A1(n3960), .A2(n3959), .ZN(n4409) );
  AND2_X1 U3688 ( .A1(n3957), .A2(n3956), .ZN(n4305) );
  AND3_X1 U3689 ( .A1(n4251), .A2(n6346), .A3(n4291), .ZN(n5777) );
  INV_X1 U3690 ( .A(n3944), .ZN(n4249) );
  OAI21_X1 U3691 ( .B1(n3876), .B2(n5064), .A(n3875), .ZN(n3878) );
  OAI21_X1 U3692 ( .B1(n3876), .B2(n5273), .A(n3790), .ZN(n5101) );
  AND2_X1 U3693 ( .A1(n3769), .A2(n3768), .ZN(n5147) );
  NOR2_X1 U3694 ( .A1(n3744), .A2(n5502), .ZN(n3767) );
  OR2_X1 U3695 ( .A1(n3048), .A2(n3046), .ZN(n3044) );
  INV_X1 U3696 ( .A(n5154), .ZN(n3048) );
  NAND2_X1 U3697 ( .A1(n3045), .A2(n2986), .ZN(n5159) );
  INV_X1 U3698 ( .A(n5112), .ZN(n3045) );
  AND2_X1 U3699 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3699), .ZN(n3700)
         );
  INV_X1 U3700 ( .A(n3698), .ZN(n3699) );
  AND2_X1 U3701 ( .A1(n3651), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3653)
         );
  NAND2_X1 U3702 ( .A1(n3653), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3698)
         );
  NOR2_X1 U3703 ( .A1(n3613), .A2(n5124), .ZN(n3614) );
  AND2_X1 U3704 ( .A1(n3614), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3651)
         );
  NAND2_X1 U3705 ( .A1(n3595), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3613)
         );
  NOR2_X1 U3706 ( .A1(n3581), .A2(n3565), .ZN(n3595) );
  NAND2_X1 U3707 ( .A1(n3564), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3581)
         );
  INV_X1 U3708 ( .A(n3563), .ZN(n3564) );
  AND2_X1 U3709 ( .A1(n3529), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3530)
         );
  INV_X1 U3710 ( .A(n4933), .ZN(n3546) );
  AND2_X1 U3711 ( .A1(n3527), .A2(n3526), .ZN(n4872) );
  AND3_X1 U3712 ( .A1(n3510), .A2(n3509), .A3(n3508), .ZN(n4862) );
  NAND2_X1 U3713 ( .A1(PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n3482), .ZN(n3511)
         );
  NAND2_X1 U3714 ( .A1(n3477), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3478)
         );
  AND2_X1 U3715 ( .A1(n3462), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3477)
         );
  NAND2_X1 U3716 ( .A1(n4682), .A2(n4681), .ZN(n4680) );
  AOI21_X1 U3717 ( .B1(n4111), .B2(n3574), .A(n3451), .ZN(n4615) );
  AOI21_X1 U3718 ( .B1(n4101), .B2(n3574), .A(n3439), .ZN(n4549) );
  NAND2_X1 U3719 ( .A1(n3399), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3435)
         );
  INV_X1 U3720 ( .A(n3376), .ZN(n3377) );
  AND2_X1 U3721 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3377), .ZN(n3399)
         );
  NAND2_X1 U3722 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3376) );
  AND2_X1 U3723 ( .A1(n4277), .A2(n4159), .ZN(n4238) );
  NOR2_X1 U3724 ( .A1(n4154), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4988)
         );
  NAND2_X1 U3725 ( .A1(n2995), .A2(n2994), .ZN(n5078) );
  INV_X1 U3726 ( .A(n5076), .ZN(n2994) );
  INV_X1 U3727 ( .A(n2995), .ZN(n5092) );
  OR2_X1 U3728 ( .A1(n5116), .A2(n3007), .ZN(n5157) );
  INV_X1 U3729 ( .A(n3009), .ZN(n3008) );
  AND2_X1 U3730 ( .A1(n4012), .A2(n5191), .ZN(n5189) );
  AND2_X1 U3731 ( .A1(n5335), .A2(n4142), .ZN(n4143) );
  NOR3_X1 U3732 ( .A1(n5223), .A2(n3005), .A3(n5125), .ZN(n5198) );
  OR2_X1 U3733 ( .A1(n5298), .A2(n5349), .ZN(n4135) );
  NOR2_X1 U3734 ( .A1(n3195), .A2(n4120), .ZN(n4121) );
  NOR2_X1 U3735 ( .A1(n4937), .A2(n4938), .ZN(n5221) );
  AND2_X1 U3736 ( .A1(n4670), .A2(n2991), .ZN(n5665) );
  INV_X1 U3737 ( .A(n5667), .ZN(n3000) );
  NAND2_X1 U3738 ( .A1(n4670), .A2(n2987), .ZN(n5666) );
  AND2_X1 U3739 ( .A1(n4670), .A2(n3001), .ZN(n4730) );
  NAND2_X1 U3740 ( .A1(n4670), .A2(n4671), .ZN(n4731) );
  AND2_X1 U3741 ( .A1(n5912), .A2(n4808), .ZN(n4956) );
  NAND2_X1 U3742 ( .A1(n2997), .A2(n2998), .ZN(n4491) );
  NOR2_X1 U3743 ( .A1(n4410), .A2(n4401), .ZN(n4489) );
  AND2_X1 U3744 ( .A1(n4301), .A2(n4996), .ZN(n5459) );
  AND2_X1 U3745 ( .A1(n4556), .A2(n6232), .ZN(n4558) );
  INV_X1 U3746 ( .A(n4472), .ZN(n4687) );
  AND2_X1 U3747 ( .A1(n6409), .A2(n4500), .ZN(n4540) );
  OR2_X1 U3748 ( .A1(n6144), .A2(n6101), .ZN(n6108) );
  OR2_X1 U3749 ( .A1(n6224), .A2(n4472), .ZN(n6144) );
  INV_X2 U3750 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6442) );
  INV_X1 U3751 ( .A(n4230), .ZN(n4244) );
  INV_X1 U3752 ( .A(n5755), .ZN(n5698) );
  INV_X1 U3753 ( .A(n5525), .ZN(n5737) );
  XNOR2_X1 U3754 ( .A(n3958), .B(n4305), .ZN(n5756) );
  AND2_X1 U3755 ( .A1(n5711), .A2(n5735), .ZN(n5525) );
  OR2_X1 U3756 ( .A1(n4754), .A2(n4717), .ZN(n5741) );
  OR3_X1 U3757 ( .A1(n4754), .A2(n3951), .A3(n4197), .ZN(n5755) );
  NAND2_X1 U3758 ( .A1(n3949), .A2(n6332), .ZN(n4939) );
  INV_X1 U3759 ( .A(n5225), .ZN(n4940) );
  INV_X1 U3760 ( .A(n5759), .ZN(n5211) );
  INV_X2 U3761 ( .A(n4939), .ZN(n5763) );
  INV_X1 U3762 ( .A(n5534), .ZN(n5771) );
  NAND2_X1 U3763 ( .A1(n4318), .A2(n4317), .ZN(n5248) );
  OAI21_X1 U3764 ( .B1(n4436), .B2(n4316), .A(n6332), .ZN(n4318) );
  CLKBUF_X1 U3765 ( .A(n4259), .Z(n4358) );
  XNOR2_X1 U3766 ( .A(n4190), .B(n4214), .ZN(n4719) );
  OR2_X1 U3767 ( .A1(n4189), .A2(n5065), .ZN(n4190) );
  OR2_X1 U3768 ( .A1(n5406), .A2(n4997), .ZN(n5393) );
  AND2_X1 U3769 ( .A1(n5001), .A2(n5443), .ZN(n5386) );
  NOR2_X1 U3770 ( .A1(n5116), .A2(n3009), .ZN(n5163) );
  NAND2_X1 U3771 ( .A1(n3015), .A2(n3019), .ZN(n5562) );
  NAND2_X1 U3772 ( .A1(n5807), .A2(n3022), .ZN(n3015) );
  NAND2_X1 U3773 ( .A1(n4792), .A2(n4128), .ZN(n4868) );
  INV_X1 U3774 ( .A(n5887), .ZN(n5908) );
  INV_X1 U3775 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6138) );
  INV_X1 U3777 ( .A(n3296), .ZN(n3260) );
  CLKBUF_X1 U3778 ( .A(n4468), .Z(n4469) );
  AND2_X1 U3779 ( .A1(n4472), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6067) );
  NAND2_X1 U3780 ( .A1(n2960), .A2(n3243), .ZN(n4447) );
  INV_X1 U3781 ( .A(n6232), .ZN(n6221) );
  OAI21_X1 U3782 ( .B1(n4467), .B2(n6410), .A(n4894), .ZN(n5921) );
  AND2_X1 U3783 ( .A1(n4466), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6323) );
  NAND2_X1 U3784 ( .A1(n6413), .A2(n6538), .ZN(n6425) );
  INV_X1 U3785 ( .A(n6323), .ZN(n6415) );
  INV_X1 U3786 ( .A(n6423), .ZN(n6418) );
  NOR2_X1 U3787 ( .A1(n2960), .A2(n5995), .ZN(n4459) );
  OR2_X1 U3788 ( .A1(n4561), .A2(n6143), .ZN(n4850) );
  INV_X1 U3789 ( .A(n5982), .ZN(n5965) );
  INV_X1 U3790 ( .A(n5990), .ZN(n5977) );
  AND2_X1 U3791 ( .A1(n4502), .A2(n6143), .ZN(n5986) );
  OR2_X1 U3792 ( .A1(n4896), .A2(n4895), .ZN(n6060) );
  INV_X1 U3793 ( .A(n6096), .ZN(n6087) );
  INV_X1 U3794 ( .A(n6108), .ZN(n6179) );
  INV_X1 U3795 ( .A(n4909), .ZN(n6223) );
  INV_X1 U3796 ( .A(n4905), .ZN(n6239) );
  INV_X1 U3797 ( .A(n6160), .ZN(n6245) );
  INV_X1 U3798 ( .A(n4914), .ZN(n6244) );
  INV_X1 U3799 ( .A(n4901), .ZN(n6251) );
  INV_X1 U3800 ( .A(n6168), .ZN(n6257) );
  INV_X1 U3801 ( .A(n4897), .ZN(n6256) );
  INV_X1 U3802 ( .A(n6172), .ZN(n6263) );
  INV_X1 U3803 ( .A(n4919), .ZN(n6262) );
  INV_X1 U3804 ( .A(n6176), .ZN(n6269) );
  INV_X1 U3805 ( .A(n6216), .ZN(n6278) );
  INV_X1 U3806 ( .A(n4837), .ZN(n6277) );
  AND2_X1 U3807 ( .A1(n6316), .A2(n6315), .ZN(n6331) );
  AND2_X1 U3808 ( .A1(n3948), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6332) );
  INV_X1 U3809 ( .A(n6338), .ZN(n6412) );
  INV_X1 U3810 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6413) );
  INV_X1 U3811 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6351) );
  AND2_X1 U3812 ( .A1(STATE_REG_1__SCAN_IN), .A2(n6351), .ZN(n6449) );
  OR2_X1 U3813 ( .A1(n5070), .A2(n5225), .ZN(n4051) );
  NAND2_X1 U3814 ( .A1(n5032), .A2(n5835), .ZN(n4172) );
  AND2_X1 U3815 ( .A1(n5058), .A2(n5057), .ZN(n5059) );
  NAND2_X1 U3816 ( .A1(n4665), .A2(n4678), .ZN(n4677) );
  AND2_X1 U3817 ( .A1(n2998), .A2(n2996), .ZN(n2979) );
  OR2_X1 U3818 ( .A1(n5078), .A2(n5015), .ZN(n2980) );
  NOR2_X1 U3819 ( .A1(n5112), .A2(n3046), .ZN(n2981) );
  AND2_X1 U3821 ( .A1(n5298), .A2(n4134), .ZN(n2983) );
  INV_X1 U3822 ( .A(n3023), .ZN(n3022) );
  NAND2_X1 U3823 ( .A1(n3055), .A2(n3024), .ZN(n3023) );
  OR2_X1 U3824 ( .A1(n4078), .A2(n3359), .ZN(n2984) );
  NAND2_X1 U3825 ( .A1(n3943), .A2(n3194), .ZN(n3199) );
  NAND2_X1 U3826 ( .A1(n3205), .A2(n3188), .ZN(n3223) );
  NOR2_X2 U3827 ( .A1(n6144), .A2(n6143), .ZN(n2985) );
  INV_X1 U3828 ( .A(n4236), .ZN(n4043) );
  NOR2_X1 U3829 ( .A1(n5168), .A2(n5167), .ZN(n2986) );
  NAND2_X1 U3830 ( .A1(n2956), .A2(n4404), .ZN(n4403) );
  AND2_X1 U3831 ( .A1(n3001), .A2(n4778), .ZN(n2987) );
  OAI21_X1 U3832 ( .B1(n5807), .B2(n4133), .A(n3055), .ZN(n4943) );
  OR2_X1 U3833 ( .A1(n5116), .A2(n5115), .ZN(n2988) );
  AND2_X1 U3834 ( .A1(n5298), .A2(n4968), .ZN(n2989) );
  AND2_X1 U3835 ( .A1(n3032), .A2(n5278), .ZN(n2990) );
  NAND2_X1 U3836 ( .A1(n4665), .A2(n3042), .ZN(n4775) );
  AND2_X1 U3837 ( .A1(n2987), .A2(n3000), .ZN(n2991) );
  INV_X1 U3838 ( .A(n3434), .ZN(n3513) );
  INV_X1 U3839 ( .A(n3513), .ZN(n4174) );
  NAND2_X1 U3840 ( .A1(n4238), .A2(n4291), .ZN(n5817) );
  INV_X1 U3841 ( .A(n5817), .ZN(n5835) );
  AND2_X1 U3842 ( .A1(n2997), .A2(n2979), .ZN(n2992) );
  OR2_X1 U3843 ( .A1(n5223), .A2(n3005), .ZN(n2993) );
  INV_X1 U3844 ( .A(n5162), .ZN(n3010) );
  AND3_X1 U3845 ( .A1(n4025), .A2(n4024), .A3(n4023), .ZN(n5162) );
  AND2_X2 U3846 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4416) );
  NAND3_X1 U3847 ( .A1(n2997), .A2(n2979), .A3(n4548), .ZN(n4617) );
  NOR2_X1 U3848 ( .A1(n5223), .A2(n5138), .ZN(n5207) );
  INV_X1 U3849 ( .A(n5208), .ZN(n3006) );
  NAND3_X1 U3850 ( .A1(n5162), .A2(n3008), .A3(n5156), .ZN(n3007) );
  NAND3_X1 U3851 ( .A1(n3375), .A2(n4470), .A3(n3374), .ZN(n3403) );
  NAND2_X1 U3852 ( .A1(n4473), .A2(n3373), .ZN(n3012) );
  NAND2_X1 U3853 ( .A1(n5807), .A2(n3016), .ZN(n3013) );
  NAND2_X1 U3854 ( .A1(n4794), .A2(n3028), .ZN(n3025) );
  NAND2_X1 U3855 ( .A1(n3025), .A2(n3026), .ZN(n4923) );
  NAND2_X1 U3856 ( .A1(n4144), .A2(n3034), .ZN(n3033) );
  OR2_X1 U3857 ( .A1(n4144), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5286)
         );
  INV_X1 U3858 ( .A(n2964), .ZN(n5327) );
  AND2_X2 U3859 ( .A1(n3069), .A2(n4457), .ZN(n3157) );
  NOR2_X4 U3860 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4457) );
  AND2_X2 U3861 ( .A1(n3061), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3069)
         );
  INV_X1 U3862 ( .A(n3882), .ZN(n3127) );
  NAND2_X1 U3863 ( .A1(n3882), .A2(n3224), .ZN(n3196) );
  AOI22_X1 U3864 ( .A1(n3272), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3123) );
  INV_X1 U3865 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3038) );
  NAND3_X1 U3866 ( .A1(n3353), .A2(n3297), .A3(n3243), .ZN(n3039) );
  NAND2_X1 U3867 ( .A1(n5085), .A2(n5087), .ZN(n5074) );
  NAND2_X1 U3868 ( .A1(n5085), .A2(n3051), .ZN(n3877) );
  CLKBUF_X1 U3869 ( .A(n4224), .Z(n5277) );
  OAI21_X2 U3870 ( .B1(n6143), .B2(n4060), .A(n4059), .ZN(n4275) );
  CLKBUF_X1 U3871 ( .A(n3220), .Z(n3222) );
  INV_X1 U3872 ( .A(n3199), .ZN(n3106) );
  XNOR2_X1 U3873 ( .A(n4176), .B(n4175), .ZN(n5230) );
  NAND2_X1 U3874 ( .A1(n3534), .A2(n3533), .ZN(n3548) );
  NAND2_X1 U3875 ( .A1(n5826), .A2(n5825), .ZN(n5824) );
  OR2_X1 U3876 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3876) );
  INV_X1 U3877 ( .A(n3876), .ZN(n3870) );
  AND2_X1 U3878 ( .A1(n3191), .A2(n3176), .ZN(n3054) );
  AND2_X1 U3879 ( .A1(n5806), .A2(n4132), .ZN(n3055) );
  OR2_X1 U3880 ( .A1(n5763), .A2(n4050), .ZN(n3056) );
  INV_X1 U3881 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4990) );
  AND4_X1 U3882 ( .A1(n3114), .A2(n3113), .A3(n3112), .A4(n3111), .ZN(n3057)
         );
  INV_X1 U3883 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6568) );
  OR2_X2 U3884 ( .A1(n5013), .A2(n6225), .ZN(n3058) );
  INV_X1 U3885 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4460) );
  NAND2_X1 U3886 ( .A1(n4163), .A2(n6232), .ZN(n6225) );
  AND2_X1 U3887 ( .A1(n4051), .A2(n3056), .ZN(n3059) );
  AND3_X1 U3888 ( .A1(n3106), .A2(n3197), .A3(n3192), .ZN(n3060) );
  NOR2_X1 U3889 ( .A1(n4749), .A2(n3909), .ZN(n3915) );
  AND2_X1 U3890 ( .A1(n6138), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3912)
         );
  INV_X1 U3891 ( .A(n5122), .ZN(n3611) );
  INV_X1 U3892 ( .A(n4872), .ZN(n3528) );
  INV_X1 U3893 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n3297) );
  AOI22_X1 U3894 ( .A1(n3137), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3091) );
  NAND2_X1 U3895 ( .A1(n3192), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3360) );
  INV_X1 U3896 ( .A(n5195), .ZN(n3632) );
  NAND2_X1 U3897 ( .A1(n4935), .A2(n3548), .ZN(n5216) );
  INV_X1 U3898 ( .A(n3348), .ZN(n3349) );
  INV_X1 U3899 ( .A(n3441), .ZN(n3444) );
  AND2_X1 U3900 ( .A1(n3771), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3772)
         );
  OR2_X1 U3901 ( .A1(n3205), .A2(n3590), .ZN(n4976) );
  OR2_X1 U3902 ( .A1(n3311), .A2(n3310), .ZN(n4057) );
  AND4_X1 U3903 ( .A1(n4444), .A2(n4443), .A3(n4442), .A4(n4441), .ZN(n4445)
         );
  AOI22_X1 U3904 ( .A1(n3851), .A2(n3850), .B1(n3870), .B2(n5023), .ZN(n4161)
         );
  AND4_X1 U3905 ( .A1(n3170), .A2(n3169), .A3(n3168), .A4(n3167), .ZN(n3171)
         );
  AND2_X1 U3906 ( .A1(n3808), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3809)
         );
  INV_X1 U3907 ( .A(n3847), .ZN(n3873) );
  NOR2_X1 U3908 ( .A1(n5292), .A2(n6476), .ZN(n4150) );
  INV_X1 U3909 ( .A(n5311), .ZN(n5291) );
  NOR2_X1 U3910 ( .A1(n5000), .A2(n5571), .ZN(n5443) );
  AND2_X1 U3911 ( .A1(n4299), .A2(n4307), .ZN(n4625) );
  INV_X1 U3912 ( .A(n6192), .ZN(n6219) );
  OR2_X1 U3913 ( .A1(n6425), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4164) );
  OR2_X1 U3914 ( .A1(n5096), .A2(n4211), .ZN(n5066) );
  OR2_X1 U3915 ( .A1(n5480), .A2(n4208), .ZN(n5096) );
  INV_X1 U3916 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5124) );
  AND4_X1 U3917 ( .A1(REIP_REG_14__SCAN_IN), .A2(n4879), .A3(
        REIP_REG_13__SCAN_IN), .A4(REIP_REG_12__SCAN_IN), .ZN(n5139) );
  OR3_X1 U3918 ( .A1(n4754), .A2(n4287), .A3(n4200), .ZN(n5711) );
  AND2_X1 U3919 ( .A1(n4719), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4720) );
  NOR2_X2 U3920 ( .A1(n3178), .A2(n6442), .ZN(n3574) );
  AND4_X1 U3921 ( .A1(n3141), .A2(n3140), .A3(n3139), .A4(n3138), .ZN(n3148)
         );
  NAND2_X1 U3922 ( .A1(n3809), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3852)
         );
  NOR2_X1 U3923 ( .A1(n6568), .A2(n3478), .ZN(n3482) );
  NOR2_X1 U3924 ( .A1(n3435), .A2(n4745), .ZN(n3436) );
  AND2_X1 U3925 ( .A1(n4076), .A2(n4075), .ZN(n4735) );
  OR2_X1 U3926 ( .A1(n6425), .A2(n6339), .ZN(n5885) );
  AND2_X1 U3927 ( .A1(n6189), .A2(n4819), .ZN(n5954) );
  AND2_X1 U3928 ( .A1(n4469), .A2(n4495), .ZN(n4502) );
  NAND2_X1 U3929 ( .A1(n4502), .A2(n6101), .ZN(n6002) );
  AND2_X1 U3930 ( .A1(n6066), .A2(n3237), .ZN(n4589) );
  INV_X1 U3931 ( .A(n4469), .ZN(n4553) );
  INV_X1 U3932 ( .A(n4689), .ZN(n6231) );
  NAND2_X1 U3933 ( .A1(n4178), .A2(n4291), .ZN(n4230) );
  OAI21_X1 U3934 ( .B1(n5062), .B2(n5755), .A(n4218), .ZN(n4219) );
  NAND2_X1 U3935 ( .A1(n3700), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3744)
         );
  AND2_X1 U3936 ( .A1(n5735), .A2(n4191), .ZN(n5692) );
  AND2_X1 U3937 ( .A1(n5735), .A2(n4720), .ZN(n5745) );
  AND2_X1 U3938 ( .A1(n5735), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5743) );
  INV_X1 U3939 ( .A(n5249), .ZN(n5250) );
  NOR2_X1 U3940 ( .A1(n4387), .A2(n5777), .ZN(n5803) );
  INV_X1 U3941 ( .A(n4317), .ZN(n4342) );
  AND2_X1 U3942 ( .A1(n5186), .A2(n5196), .ZN(n5764) );
  NAND2_X1 U3943 ( .A1(n3530), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3563)
         );
  AOI21_X1 U3944 ( .B1(n5056), .B2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5055), 
        .ZN(n5057) );
  OR2_X1 U3945 ( .A1(n5393), .A2(n4998), .ZN(n5372) );
  NAND2_X1 U3946 ( .A1(n4622), .A2(n4621), .ZN(n4624) );
  INV_X1 U3947 ( .A(n5846), .ZN(n5914) );
  INV_X1 U3948 ( .A(n4996), .ZN(n5912) );
  INV_X1 U3949 ( .A(n4850), .ZN(n4857) );
  OAI221_X1 U3950 ( .B1(n4824), .B2(n6413), .C1(n4824), .C2(n4823), .A(n4822), 
        .ZN(n4854) );
  INV_X1 U3951 ( .A(n2971), .ZN(n6189) );
  INV_X1 U3952 ( .A(n6002), .ZN(n6019) );
  INV_X1 U3953 ( .A(n6063), .ZN(n6047) );
  OAI211_X1 U3954 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6442), .A(n4822), .B(n4637), .ZN(n4659) );
  OR2_X1 U3955 ( .A1(n6107), .A2(n6106), .ZN(n6132) );
  NAND2_X1 U3956 ( .A1(n4077), .A2(n4553), .ZN(n6065) );
  INV_X1 U3957 ( .A(n4894), .ZN(n4634) );
  NOR2_X1 U3958 ( .A1(n6464), .A2(n4894), .ZN(n6222) );
  NOR2_X1 U3959 ( .A1(n6459), .A2(n4894), .ZN(n6250) );
  INV_X1 U3960 ( .A(n4842), .ZN(n6268) );
  NOR2_X1 U3961 ( .A1(n6538), .A2(n6442), .ZN(n4479) );
  AND2_X1 U3962 ( .A1(n4230), .A2(n4231), .ZN(n6452) );
  INV_X1 U3963 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6455) );
  INV_X1 U3964 ( .A(n4219), .ZN(n4220) );
  INV_X1 U3965 ( .A(n5743), .ZN(n5678) );
  INV_X1 U3966 ( .A(n5692), .ZN(n5673) );
  INV_X1 U3967 ( .A(n4940), .ZN(n5758) );
  NAND2_X1 U3968 ( .A1(n5228), .A2(n5763), .ZN(n5225) );
  INV_X1 U3969 ( .A(n5777), .ZN(n5805) );
  OR2_X1 U3970 ( .A1(n5823), .A2(n4363), .ZN(n5840) );
  XNOR2_X1 U3971 ( .A(n4991), .B(n4990), .ZN(n5012) );
  NAND2_X1 U3972 ( .A1(n4307), .A2(n4297), .ZN(n5846) );
  INV_X1 U3973 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6313) );
  OR2_X1 U3974 ( .A1(n5602), .A2(n6409), .ZN(n6423) );
  AND2_X1 U3975 ( .A1(n4826), .A2(n4825), .ZN(n4860) );
  NAND2_X1 U3976 ( .A1(n4818), .A2(n4817), .ZN(n5982) );
  INV_X1 U3977 ( .A(n5986), .ZN(n4613) );
  OR2_X1 U3978 ( .A1(n5991), .A2(n6185), .ZN(n6053) );
  INV_X1 U3979 ( .A(n6059), .ZN(n4913) );
  OR2_X1 U3980 ( .A1(n6065), .A2(n4631), .ZN(n4713) );
  OR2_X1 U3981 ( .A1(n6065), .A2(n6185), .ZN(n6096) );
  OR2_X1 U3982 ( .A1(n6065), .A2(n6064), .ZN(n6135) );
  OR2_X1 U3983 ( .A1(n6224), .A2(n6185), .ZN(n6216) );
  OR2_X1 U3984 ( .A1(n6224), .A2(n6064), .ZN(n6283) );
  AND2_X1 U3985 ( .A1(n6322), .A2(n6321), .ZN(n6338) );
  INV_X1 U3986 ( .A(n6408), .ZN(n6406) );
  INV_X1 U3987 ( .A(READY_N), .ZN(n6345) );
  INV_X1 U3988 ( .A(n6608), .ZN(n6398) );
  INV_X1 U3989 ( .A(n6609), .ZN(n6403) );
  OAI21_X1 U3990 ( .B1(n5235), .B2(n5759), .A(n3059), .ZN(U2829) );
  INV_X1 U3991 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3061) );
  INV_X1 U3992 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3062) );
  AND2_X2 U3993 ( .A1(n3069), .A2(n4974), .ZN(n3272) );
  AND2_X2 U3994 ( .A1(n4974), .A2(n4426), .ZN(n3304) );
  AOI22_X1 U3995 ( .A1(n3137), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3066) );
  AOI22_X1 U3996 ( .A1(n3273), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3065) );
  AOI22_X1 U3997 ( .A1(n3298), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n2978), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3064) );
  AOI22_X1 U3998 ( .A1(n3280), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3073) );
  AND2_X2 U3999 ( .A1(n4975), .A2(n3069), .ZN(n3152) );
  AND2_X2 U4000 ( .A1(n4975), .A2(n4426), .ZN(n3275) );
  AND2_X2 U4001 ( .A1(n4426), .A2(n4425), .ZN(n3142) );
  AOI22_X1 U4002 ( .A1(n3275), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3142), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3070) );
  AOI22_X1 U4003 ( .A1(n3304), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3079) );
  AOI22_X1 U4004 ( .A1(n3272), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3078) );
  AOI22_X1 U4005 ( .A1(n3298), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n2978), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3077) );
  AOI22_X1 U4006 ( .A1(n3128), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3076) );
  AND4_X2 U4007 ( .A1(n3079), .A2(n3078), .A3(n3077), .A4(n3076), .ZN(n3085)
         );
  AOI22_X1 U4008 ( .A1(n3152), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3083) );
  AOI22_X1 U4009 ( .A1(n3275), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3082) );
  AOI22_X1 U4010 ( .A1(n3142), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3081) );
  AOI22_X1 U4011 ( .A1(n3274), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3080) );
  AOI22_X1 U4012 ( .A1(n3273), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3089) );
  AOI22_X1 U4013 ( .A1(n3275), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3088) );
  AOI22_X1 U4014 ( .A1(n3280), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3087) );
  AOI22_X1 U4015 ( .A1(n3272), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3142), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3086) );
  AOI22_X1 U4016 ( .A1(n3152), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3093) );
  AOI22_X1 U4017 ( .A1(n3298), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n2977), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3090) );
  INV_X2 U4018 ( .A(n3187), .ZN(n3194) );
  AOI22_X1 U4019 ( .A1(n3152), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3097) );
  AOI22_X1 U4020 ( .A1(n3298), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n2977), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3096) );
  NAND4_X1 U4021 ( .A1(n3099), .A2(n3098), .A3(n3097), .A4(n3096), .ZN(n3105)
         );
  AOI22_X1 U4022 ( .A1(n3275), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n2972), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3103) );
  AOI22_X1 U4023 ( .A1(n3273), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3102) );
  AOI22_X1 U4024 ( .A1(n3272), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3142), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3101) );
  AOI22_X1 U4025 ( .A1(n3280), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3100) );
  NAND4_X1 U4026 ( .A1(n3103), .A2(n3102), .A3(n3101), .A4(n3100), .ZN(n3104)
         );
  AOI22_X1 U4027 ( .A1(n3137), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3110) );
  AOI22_X1 U4028 ( .A1(n2975), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3274), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3109) );
  AOI22_X1 U4029 ( .A1(n3298), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n2977), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3108) );
  AOI22_X1 U4030 ( .A1(n3152), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3107) );
  AOI22_X1 U4031 ( .A1(n3275), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n2972), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3114) );
  AOI22_X1 U4032 ( .A1(n3273), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3113) );
  AOI22_X1 U4033 ( .A1(n3272), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3142), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3112) );
  AOI22_X1 U4034 ( .A1(n3280), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3111) );
  NAND2_X1 U4035 ( .A1(n3115), .A2(n3057), .ZN(n3198) );
  AOI22_X1 U4036 ( .A1(n3152), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3119) );
  AOI22_X1 U4037 ( .A1(n2976), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3274), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3118) );
  AOI22_X1 U4038 ( .A1(n3273), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3117) );
  AOI22_X1 U4039 ( .A1(n3298), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n2978), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3116) );
  NAND4_X1 U4040 ( .A1(n3119), .A2(n3118), .A3(n3117), .A4(n3116), .ZN(n3125)
         );
  AOI22_X1 U4041 ( .A1(n3137), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3122) );
  AOI22_X1 U4042 ( .A1(n3275), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3121) );
  NAND4_X1 U4043 ( .A1(n3123), .A2(n3122), .A3(n3121), .A4(n3120), .ZN(n3124)
         );
  OR2_X2 U4044 ( .A1(n3125), .A2(n3124), .ZN(n3188) );
  AND3_X1 U4045 ( .A1(n4290), .A2(n3176), .A3(n3188), .ZN(n3126) );
  NAND2_X1 U4046 ( .A1(n3127), .A2(n3126), .ZN(n4245) );
  INV_X1 U4047 ( .A(n4245), .ZN(n3151) );
  NAND2_X1 U4048 ( .A1(n3152), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3131) );
  NAND2_X1 U4049 ( .A1(n3128), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3130)
         );
  NAND2_X1 U4050 ( .A1(n3274), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3129) );
  NAND2_X1 U4051 ( .A1(n3273), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3136)
         );
  NAND2_X1 U4052 ( .A1(n3275), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3135) );
  NAND2_X1 U4053 ( .A1(n3304), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3134) );
  NAND2_X1 U4054 ( .A1(n2972), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3133) );
  NAND2_X1 U4055 ( .A1(n3137), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3141)
         );
  NAND2_X1 U4056 ( .A1(n3298), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3140) );
  NAND2_X1 U4057 ( .A1(n3244), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3139)
         );
  NAND2_X1 U4058 ( .A1(n2978), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3138)
         );
  NAND2_X1 U4059 ( .A1(n3272), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3146) );
  NAND2_X1 U4060 ( .A1(n3280), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3145) );
  NAND2_X1 U4061 ( .A1(n3249), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3144)
         );
  NAND2_X1 U4062 ( .A1(n3142), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3143) );
  NAND4_X4 U4063 ( .A1(n3150), .A2(n3149), .A3(n3148), .A4(n3147), .ZN(n4715)
         );
  NAND2_X1 U4064 ( .A1(n3151), .A2(n4715), .ZN(n4177) );
  NAND2_X1 U4065 ( .A1(n2976), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3156)
         );
  NAND2_X1 U4066 ( .A1(n3152), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3155) );
  NAND2_X1 U4067 ( .A1(n3137), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3154)
         );
  NAND2_X1 U4068 ( .A1(n3244), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3153)
         );
  NAND2_X1 U4069 ( .A1(n3274), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3162) );
  NAND2_X1 U4070 ( .A1(n3157), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3161) );
  NAND2_X1 U4071 ( .A1(n3298), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3160) );
  NAND2_X1 U4072 ( .A1(n2977), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3159)
         );
  NAND2_X1 U4073 ( .A1(n3272), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3166) );
  NAND2_X1 U4074 ( .A1(n3280), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3165) );
  NAND2_X1 U4075 ( .A1(n3273), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3164)
         );
  NAND2_X1 U4076 ( .A1(n3142), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3163) );
  NAND2_X1 U4077 ( .A1(n3275), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3170) );
  NAND2_X1 U4078 ( .A1(n3304), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3169) );
  NAND2_X1 U4079 ( .A1(n2973), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3168) );
  NAND2_X1 U4080 ( .A1(n3249), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3167)
         );
  INV_X1 U4081 ( .A(STATE_REG_2__SCAN_IN), .ZN(n3175) );
  XNOR2_X1 U4082 ( .A(n3175), .B(STATE_REG_1__SCAN_IN), .ZN(n4198) );
  INV_X1 U4083 ( .A(n3191), .ZN(n3182) );
  NOR2_X1 U4084 ( .A1(n3193), .A2(n3188), .ZN(n3177) );
  NAND3_X1 U4085 ( .A1(n3177), .A2(n4749), .A3(n4290), .ZN(n4419) );
  NAND2_X2 U4086 ( .A1(n3193), .A2(n3180), .ZN(n3205) );
  AND3_X2 U4087 ( .A1(n3179), .A2(n3223), .A3(n4501), .ZN(n3201) );
  NAND2_X1 U4088 ( .A1(n3201), .A2(n3060), .ZN(n4179) );
  NAND2_X1 U4089 ( .A1(n3183), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3210) );
  INV_X1 U4090 ( .A(n4164), .ZN(n3211) );
  XNOR2_X1 U4091 ( .A(n6138), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6186)
         );
  INV_X1 U4092 ( .A(n3948), .ZN(n3212) );
  AND2_X1 U4093 ( .A1(n3212), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3184)
         );
  AOI21_X1 U4094 ( .B1(n3211), .B2(n6186), .A(n3184), .ZN(n3208) );
  INV_X1 U4095 ( .A(n3208), .ZN(n3185) );
  NOR2_X1 U4096 ( .A1(n3185), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3186)
         );
  OAI211_X1 U4097 ( .C1(n3205), .C2(n3187), .A(n3189), .B(n3943), .ZN(n3220)
         );
  INV_X1 U4098 ( .A(n3220), .ZN(n3190) );
  NOR2_X2 U4099 ( .A1(n3944), .A2(n3192), .ZN(n3224) );
  INV_X1 U4100 ( .A(n3216), .ZN(n3195) );
  INV_X1 U4101 ( .A(n3197), .ZN(n3225) );
  NAND3_X1 U4102 ( .A1(n3201), .A2(n4249), .A3(n3200), .ZN(n3202) );
  NAND2_X1 U4103 ( .A1(n3202), .A2(n3192), .ZN(n3217) );
  NAND3_X1 U4104 ( .A1(n3217), .A2(n3228), .A3(n3203), .ZN(n3204) );
  NAND2_X1 U4105 ( .A1(n3204), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3207) );
  NAND2_X1 U4106 ( .A1(n3205), .A2(n3905), .ZN(n3206) );
  NAND2_X1 U4107 ( .A1(n3234), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3209) );
  NAND3_X1 U4108 ( .A1(n3210), .A2(n3209), .A3(n3208), .ZN(n3232) );
  AND2_X2 U4109 ( .A1(n2982), .A2(n3232), .ZN(n3259) );
  NAND2_X1 U4110 ( .A1(n3234), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3215) );
  MUX2_X1 U4111 ( .A(n3212), .B(n3211), .S(n6138), .Z(n3213) );
  INV_X1 U4112 ( .A(n3213), .ZN(n3214) );
  NAND2_X1 U4113 ( .A1(n3215), .A2(n3214), .ZN(n3292) );
  NAND2_X1 U4114 ( .A1(n4527), .A2(n4715), .ZN(n3218) );
  AND2_X1 U4115 ( .A1(n3205), .A2(n3187), .ZN(n3221) );
  OAI21_X1 U4116 ( .B1(n3222), .B2(n3221), .A(n4517), .ZN(n3227) );
  NOR2_X1 U4117 ( .A1(n6425), .A2(n3297), .ZN(n6333) );
  NAND2_X1 U4118 ( .A1(n3223), .A2(n2954), .ZN(n3226) );
  NOR2_X1 U4119 ( .A1(n4527), .A2(n3188), .ZN(n3945) );
  NAND4_X1 U4120 ( .A1(n3225), .A2(n3192), .A3(n3945), .A4(n3187), .ZN(n4450)
         );
  NAND4_X1 U4121 ( .A1(n3227), .A2(n6333), .A3(n3226), .A4(n4450), .ZN(n3230)
         );
  INV_X1 U4122 ( .A(n3228), .ZN(n3229) );
  NOR2_X1 U4123 ( .A1(n3230), .A2(n3229), .ZN(n3231) );
  NAND2_X1 U4124 ( .A1(n3888), .A2(n3231), .ZN(n3291) );
  NAND2_X1 U4125 ( .A1(n3259), .A2(n3296), .ZN(n3233) );
  NAND2_X1 U4126 ( .A1(n3233), .A2(n3232), .ZN(n3242) );
  INV_X1 U4127 ( .A(n3242), .ZN(n3240) );
  AND2_X1 U4128 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3235) );
  NAND2_X1 U4129 ( .A1(n3235), .A2(n6305), .ZN(n6066) );
  INV_X1 U4130 ( .A(n3235), .ZN(n3236) );
  NAND2_X1 U4131 ( .A1(n3236), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3237) );
  OAI22_X1 U4132 ( .A1(n4589), .A2(n4164), .B1(n3948), .B2(n6305), .ZN(n3238)
         );
  INV_X1 U4133 ( .A(n3241), .ZN(n3239) );
  NAND2_X1 U4134 ( .A1(n3242), .A2(n3241), .ZN(n3243) );
  AOI22_X1 U4135 ( .A1(n3833), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3820), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3248) );
  AOI22_X1 U4136 ( .A1(n2975), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3247) );
  AOI22_X1 U4137 ( .A1(n3834), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3246) );
  AOI22_X1 U4138 ( .A1(n3750), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n2977), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3245) );
  NAND4_X1 U4139 ( .A1(n3248), .A2(n3247), .A3(n3246), .A4(n3245), .ZN(n3255)
         );
  AOI22_X1 U4140 ( .A1(n3821), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3253) );
  AOI22_X1 U4141 ( .A1(n3861), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3252) );
  CLKBUF_X2 U4142 ( .A(n3142), .Z(n3305) );
  AOI22_X1 U4143 ( .A1(n3822), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3251) );
  AOI22_X1 U4144 ( .A1(n3303), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3250) );
  NAND4_X1 U4145 ( .A1(n3253), .A2(n3252), .A3(n3251), .A4(n3250), .ZN(n3254)
         );
  NOR2_X1 U4146 ( .A1(n3255), .A2(n3254), .ZN(n4078) );
  INV_X1 U4147 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3256) );
  OAI22_X1 U4148 ( .A1(n3360), .A2(n4078), .B1(n3931), .B2(n3256), .ZN(n3257)
         );
  XNOR2_X2 U4149 ( .A(n3258), .B(n3257), .ZN(n3352) );
  XNOR2_X2 U4150 ( .A(n3259), .B(n3260), .ZN(n4496) );
  INV_X1 U4151 ( .A(n3359), .ZN(n3316) );
  AOI22_X1 U4152 ( .A1(n2953), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3820), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3264) );
  AOI22_X1 U4153 ( .A1(n3834), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3750), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3263) );
  AOI22_X1 U4154 ( .A1(n3833), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3821), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3262) );
  AOI22_X1 U4155 ( .A1(n3860), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3261) );
  NAND4_X1 U4156 ( .A1(n3264), .A2(n3263), .A3(n3262), .A4(n3261), .ZN(n3270)
         );
  AOI22_X1 U4157 ( .A1(n3822), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3303), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3268) );
  AOI22_X1 U4158 ( .A1(n3861), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3267) );
  AOI22_X1 U4159 ( .A1(n2975), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n2972), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3266) );
  AOI22_X1 U4160 ( .A1(n3731), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n2978), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3265) );
  NAND4_X1 U4161 ( .A1(n3268), .A2(n3267), .A3(n3266), .A4(n3265), .ZN(n3269)
         );
  NAND2_X1 U4162 ( .A1(n3316), .A2(n4064), .ZN(n3271) );
  INV_X1 U4163 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3290) );
  AOI22_X1 U4164 ( .A1(n3822), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3821), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3279) );
  AOI22_X1 U4165 ( .A1(n2975), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3820), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3278) );
  AOI22_X1 U4166 ( .A1(n2953), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3277) );
  AOI22_X1 U4167 ( .A1(n3275), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n2972), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3276) );
  NAND4_X1 U4168 ( .A1(n3279), .A2(n3278), .A3(n3277), .A4(n3276), .ZN(n3286)
         );
  AOI22_X1 U4169 ( .A1(n3833), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3284) );
  AOI22_X1 U4170 ( .A1(n3860), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3283) );
  AOI22_X1 U4171 ( .A1(n3750), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n2977), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3282) );
  BUF_X1 U4172 ( .A(n3280), .Z(n3303) );
  AOI22_X1 U4173 ( .A1(n3303), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3281) );
  NAND4_X1 U4174 ( .A1(n3284), .A2(n3283), .A3(n3282), .A4(n3281), .ZN(n3285)
         );
  NOR2_X1 U4175 ( .A1(n3359), .A2(n4123), .ZN(n3315) );
  INV_X1 U4176 ( .A(n3315), .ZN(n3289) );
  INV_X1 U4177 ( .A(n3360), .ZN(n3287) );
  NAND2_X1 U4178 ( .A1(n3287), .A2(n4064), .ZN(n3288) );
  OAI211_X1 U4179 ( .C1(n3290), .C2(n3931), .A(n3289), .B(n3288), .ZN(n3327)
         );
  INV_X1 U4180 ( .A(n3291), .ZN(n3294) );
  INV_X1 U4181 ( .A(n3292), .ZN(n3293) );
  NAND2_X1 U4182 ( .A1(n3294), .A2(n3293), .ZN(n3295) );
  NAND2_X2 U4183 ( .A1(n3296), .A2(n3295), .ZN(n3342) );
  AOI22_X1 U4184 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n2975), .B1(n3861), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4185 ( .A1(n3834), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3750), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4186 ( .A1(n2953), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U4187 ( .A1(n3821), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3299) );
  NAND4_X1 U4188 ( .A1(n3302), .A2(n3301), .A3(n3300), .A4(n3299), .ZN(n3311)
         );
  AOI22_X1 U4189 ( .A1(n3822), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3303), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4190 ( .A1(n3860), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4191 ( .A1(n3833), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3307) );
  AOI22_X1 U4192 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n3820), .B1(n2978), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3306) );
  NAND4_X1 U4193 ( .A1(n3309), .A2(n3308), .A3(n3307), .A4(n3306), .ZN(n3310)
         );
  INV_X1 U4194 ( .A(n4057), .ZN(n4065) );
  NAND2_X1 U4195 ( .A1(n3194), .A2(n4065), .ZN(n3312) );
  NAND2_X1 U4196 ( .A1(n3315), .A2(n4057), .ZN(n3338) );
  AND2_X1 U4197 ( .A1(n3338), .A2(n3359), .ZN(n3317) );
  NAND2_X1 U4198 ( .A1(n3335), .A2(n3317), .ZN(n3321) );
  INV_X1 U4199 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3320) );
  AOI21_X1 U4200 ( .B1(n3194), .B2(n4123), .A(n3297), .ZN(n3319) );
  NAND2_X1 U4201 ( .A1(n3192), .A2(n4057), .ZN(n3318) );
  OAI211_X1 U4202 ( .C1(n3931), .C2(n3320), .A(n3319), .B(n3318), .ZN(n3337)
         );
  NAND2_X1 U4203 ( .A1(n3328), .A2(n3327), .ZN(n3322) );
  XNOR2_X2 U4204 ( .A(n3352), .B(n3374), .ZN(n4468) );
  NAND2_X1 U4205 ( .A1(n4468), .A2(n3574), .ZN(n3324) );
  NAND2_X1 U4206 ( .A1(n6442), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3745) );
  NAND2_X1 U4207 ( .A1(n3324), .A2(n3745), .ZN(n3347) );
  INV_X1 U4208 ( .A(n4288), .ZN(n5019) );
  NAND2_X1 U4209 ( .A1(n5019), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3397) );
  OAI21_X1 U4210 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3376), .ZN(n5839) );
  AOI22_X1 U4211 ( .A1(n4173), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n3870), 
        .B2(n5839), .ZN(n3326) );
  NOR2_X2 U4212 ( .A1(n4501), .A2(n6442), .ZN(n3434) );
  NAND2_X1 U4213 ( .A1(n4174), .A2(EAX_REG_2__SCAN_IN), .ZN(n3325) );
  NAND2_X1 U4214 ( .A1(n3347), .A2(n3348), .ZN(n3346) );
  XNOR2_X1 U4215 ( .A(n3328), .B(n3327), .ZN(n3330) );
  NAND2_X1 U4216 ( .A1(n4471), .A2(n3574), .ZN(n3334) );
  AOI22_X1 U4217 ( .A1(n4174), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6442), .ZN(n3332) );
  INV_X1 U4218 ( .A(n3397), .ZN(n3343) );
  NAND2_X1 U4219 ( .A1(n3343), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3331) );
  AND2_X1 U4220 ( .A1(n3332), .A2(n3331), .ZN(n3333) );
  NAND2_X1 U4221 ( .A1(n3334), .A2(n3333), .ZN(n4390) );
  NAND2_X1 U4222 ( .A1(n3335), .A2(n3338), .ZN(n3336) );
  NAND2_X1 U4223 ( .A1(n3336), .A2(n3337), .ZN(n3341) );
  INV_X1 U4224 ( .A(n3337), .ZN(n3339) );
  NAND2_X1 U4225 ( .A1(n3339), .A2(n3338), .ZN(n3340) );
  AOI21_X1 U4226 ( .B1(n6143), .B2(n3225), .A(n6442), .ZN(n4320) );
  INV_X1 U4227 ( .A(n3574), .ZN(n3562) );
  AOI22_X1 U4228 ( .A1(n4174), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6442), .ZN(n3345) );
  NAND2_X1 U4229 ( .A1(n3343), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3344) );
  OAI211_X1 U4230 ( .C1(n3342), .C2(n3562), .A(n3345), .B(n3344), .ZN(n4319)
         );
  MUX2_X1 U4231 ( .A(n3870), .B(n4320), .S(n4319), .Z(n4391) );
  NAND2_X1 U4232 ( .A1(n4390), .A2(n4391), .ZN(n4398) );
  NAND2_X1 U4233 ( .A1(n3346), .A2(n4398), .ZN(n3351) );
  INV_X1 U4234 ( .A(n3347), .ZN(n3350) );
  INV_X1 U4235 ( .A(n3352), .ZN(n3375) );
  NAND2_X1 U4236 ( .A1(n3375), .A2(n3374), .ZN(n3373) );
  NAND2_X1 U4237 ( .A1(n2959), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3358) );
  NAND3_X1 U4238 ( .A1(n6313), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6031) );
  INV_X1 U4239 ( .A(n6031), .ZN(n3354) );
  NAND2_X1 U4240 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3354), .ZN(n6026) );
  NAND2_X1 U4241 ( .A1(n6313), .A2(n6026), .ZN(n3355) );
  NAND3_X1 U4242 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6220) );
  INV_X1 U4243 ( .A(n6220), .ZN(n6233) );
  NAND2_X1 U4244 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6233), .ZN(n6217) );
  NAND2_X1 U4245 ( .A1(n3355), .A2(n6217), .ZN(n4888) );
  OAI22_X1 U4246 ( .A1(n4164), .A2(n4888), .B1(n3948), .B2(n6313), .ZN(n3356)
         );
  INV_X1 U4247 ( .A(n3356), .ZN(n3357) );
  NAND2_X1 U4248 ( .A1(n4417), .A2(n3297), .ZN(n3372) );
  AOI22_X1 U4249 ( .A1(n3833), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3820), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3364) );
  INV_X1 U4250 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n6593) );
  AOI22_X1 U4251 ( .A1(n2975), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3363) );
  AOI22_X1 U4252 ( .A1(n3834), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3362) );
  AOI22_X1 U4253 ( .A1(n3750), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n2978), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3361) );
  NAND4_X1 U4254 ( .A1(n3364), .A2(n3363), .A3(n3362), .A4(n3361), .ZN(n3370)
         );
  AOI22_X1 U4255 ( .A1(n3821), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4256 ( .A1(n3861), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4257 ( .A1(n3822), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4258 ( .A1(n3303), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3365) );
  NAND4_X1 U4259 ( .A1(n3368), .A2(n3367), .A3(n3366), .A4(n3365), .ZN(n3369)
         );
  AOI22_X1 U4260 ( .A1(n3919), .A2(n4086), .B1(n3905), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3371) );
  INV_X1 U4261 ( .A(n4470), .ZN(n4473) );
  NOR2_X1 U4262 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3377), .ZN(n3378)
         );
  NOR2_X1 U4263 ( .A1(n3399), .A2(n3378), .ZN(n5725) );
  INV_X1 U4264 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4738) );
  OAI22_X1 U4265 ( .A1(n5725), .A2(n3876), .B1(n3745), .B2(n4738), .ZN(n3379)
         );
  AOI21_X1 U4266 ( .B1(n3434), .B2(EAX_REG_3__SCAN_IN), .A(n3379), .ZN(n3380)
         );
  OAI21_X1 U4267 ( .B1(n3061), .B2(n3397), .A(n3380), .ZN(n3381) );
  INV_X1 U4268 ( .A(n3382), .ZN(n4396) );
  AOI22_X1 U4269 ( .A1(n3834), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3750), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3386) );
  AOI22_X1 U4270 ( .A1(n2974), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3385) );
  AOI22_X1 U4271 ( .A1(n3833), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3384) );
  AOI22_X1 U4272 ( .A1(n3861), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3383) );
  NAND4_X1 U4273 ( .A1(n3386), .A2(n3385), .A3(n3384), .A4(n3383), .ZN(n3392)
         );
  AOI22_X1 U4274 ( .A1(n3822), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3390) );
  AOI22_X1 U4275 ( .A1(n3820), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3821), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3389) );
  AOI22_X1 U4276 ( .A1(n3303), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3388) );
  AOI22_X1 U4277 ( .A1(n2953), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n2978), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3387) );
  NAND4_X1 U4278 ( .A1(n3390), .A2(n3389), .A3(n3388), .A4(n3387), .ZN(n3391)
         );
  NAND2_X1 U4279 ( .A1(n3919), .A2(n4102), .ZN(n3394) );
  NAND2_X1 U4280 ( .A1(n3905), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3393) );
  NAND2_X1 U4281 ( .A1(n3394), .A2(n3393), .ZN(n3421) );
  NAND2_X1 U4282 ( .A1(n6442), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3396)
         );
  NAND2_X1 U4283 ( .A1(n4174), .A2(EAX_REG_4__SCAN_IN), .ZN(n3395) );
  OAI211_X1 U4284 ( .C1(n3397), .C2(n4460), .A(n3396), .B(n3395), .ZN(n3398)
         );
  NAND2_X1 U4285 ( .A1(n3398), .A2(n3876), .ZN(n3401) );
  OAI21_X1 U4286 ( .B1(n3399), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3435), 
        .ZN(n5831) );
  NAND2_X1 U4287 ( .A1(n5831), .A2(n3870), .ZN(n3400) );
  NAND2_X1 U4288 ( .A1(n3401), .A2(n3400), .ZN(n3402) );
  AOI21_X1 U4289 ( .B1(n4085), .B2(n3574), .A(n3402), .ZN(n4486) );
  NAND2_X1 U4290 ( .A1(n3423), .A2(n3421), .ZN(n3416) );
  AOI22_X1 U4291 ( .A1(n3833), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3820), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3407) );
  AOI22_X1 U4292 ( .A1(n2975), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3406) );
  AOI22_X1 U4293 ( .A1(n3834), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3405) );
  INV_X1 U4294 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n6594) );
  AOI22_X1 U4295 ( .A1(n3750), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n2978), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3404) );
  NAND4_X1 U4296 ( .A1(n3407), .A2(n3406), .A3(n3405), .A4(n3404), .ZN(n3413)
         );
  AOI22_X1 U4297 ( .A1(n3821), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3411) );
  AOI22_X1 U4298 ( .A1(n3861), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n2972), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3410) );
  AOI22_X1 U4299 ( .A1(n3822), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3409) );
  AOI22_X1 U4300 ( .A1(n3303), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3408) );
  NAND4_X1 U4301 ( .A1(n3411), .A2(n3410), .A3(n3409), .A4(n3408), .ZN(n3412)
         );
  NAND2_X1 U4302 ( .A1(n3919), .A2(n4103), .ZN(n3415) );
  NAND2_X1 U4303 ( .A1(n3905), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3414) );
  NAND2_X1 U4304 ( .A1(n3415), .A2(n3414), .ZN(n3420) );
  NAND2_X1 U4305 ( .A1(n4093), .A2(n3574), .ZN(n3419) );
  XNOR2_X1 U4306 ( .A(n3435), .B(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5700) );
  INV_X1 U4307 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4745) );
  OAI22_X1 U4308 ( .A1(n5700), .A2(n3876), .B1(n3745), .B2(n4745), .ZN(n3417)
         );
  AOI21_X1 U4309 ( .B1(n3434), .B2(EAX_REG_5__SCAN_IN), .A(n3417), .ZN(n3418)
         );
  NAND2_X1 U4310 ( .A1(n3419), .A2(n3418), .ZN(n4404) );
  AOI22_X1 U4311 ( .A1(n3833), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3820), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3427) );
  AOI22_X1 U4312 ( .A1(n2975), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3426) );
  AOI22_X1 U4313 ( .A1(n3834), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3425) );
  AOI22_X1 U4314 ( .A1(n3750), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n2978), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3424) );
  NAND4_X1 U4315 ( .A1(n3427), .A2(n3426), .A3(n3425), .A4(n3424), .ZN(n3433)
         );
  AOI22_X1 U4316 ( .A1(n3821), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4317 ( .A1(n3861), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4318 ( .A1(n3822), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4319 ( .A1(n3303), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3428) );
  NAND4_X1 U4320 ( .A1(n3431), .A2(n3430), .A3(n3429), .A4(n3428), .ZN(n3432)
         );
  AOI22_X1 U4321 ( .A1(n3919), .A2(n4113), .B1(n3905), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3442) );
  NAND2_X1 U4322 ( .A1(n3441), .A2(n3442), .ZN(n4101) );
  INV_X1 U4323 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4551) );
  NOR2_X1 U4324 ( .A1(n3436), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3437)
         );
  OR2_X1 U4325 ( .A1(n3462), .A2(n3437), .ZN(n5822) );
  AOI22_X1 U4326 ( .A1(n5822), .A2(n3870), .B1(n4173), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3438) );
  OAI21_X1 U4327 ( .B1(n3513), .B2(n4551), .A(n3438), .ZN(n3439) );
  INV_X1 U4328 ( .A(n4549), .ZN(n3440) );
  INV_X1 U4329 ( .A(n3442), .ZN(n3443) );
  INV_X1 U4330 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3446) );
  NAND2_X1 U4331 ( .A1(n3919), .A2(n4123), .ZN(n3445) );
  OAI21_X1 U4332 ( .B1(n3446), .B2(n3931), .A(n3445), .ZN(n3447) );
  INV_X1 U4333 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3450) );
  XNOR2_X1 U4334 ( .A(n3462), .B(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4769) );
  NAND2_X1 U4335 ( .A1(n4769), .A2(n3870), .ZN(n3449) );
  NAND2_X1 U4336 ( .A1(n4173), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3448)
         );
  OAI211_X1 U4337 ( .C1(n3513), .C2(n3450), .A(n3449), .B(n3448), .ZN(n3451)
         );
  AOI22_X1 U4338 ( .A1(n3822), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3303), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4339 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n3833), .B1(n3861), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4340 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n2974), .B1(n2953), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3453) );
  AOI22_X1 U4341 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n3750), .B1(n3731), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3452) );
  NAND4_X1 U4342 ( .A1(n3455), .A2(n3454), .A3(n3453), .A4(n3452), .ZN(n3461)
         );
  AOI22_X1 U4343 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n3821), .B1(n3860), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3459) );
  AOI22_X1 U4344 ( .A1(n3820), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3458) );
  AOI22_X1 U4345 ( .A1(n3834), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3457) );
  AOI22_X1 U4346 ( .A1(n3305), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3456) );
  NAND4_X1 U4347 ( .A1(n3459), .A2(n3458), .A3(n3457), .A4(n3456), .ZN(n3460)
         );
  OAI21_X1 U4348 ( .B1(n3461), .B2(n3460), .A(n3574), .ZN(n3466) );
  NAND2_X1 U4349 ( .A1(n3434), .A2(EAX_REG_8__SCAN_IN), .ZN(n3465) );
  XNOR2_X1 U4350 ( .A(n3477), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4798) );
  NAND2_X1 U4351 ( .A1(n4798), .A2(n3870), .ZN(n3464) );
  NAND2_X1 U4352 ( .A1(n4173), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3463)
         );
  NAND4_X1 U4353 ( .A1(n3466), .A2(n3465), .A3(n3464), .A4(n3463), .ZN(n4667)
         );
  AOI22_X1 U4354 ( .A1(n3821), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3470) );
  AOI22_X1 U4355 ( .A1(n2975), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3820), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3469) );
  AOI22_X1 U4356 ( .A1(n2953), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3468) );
  AOI22_X1 U4357 ( .A1(n3861), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3467) );
  NAND4_X1 U4358 ( .A1(n3470), .A2(n3469), .A3(n3468), .A4(n3467), .ZN(n3476)
         );
  AOI22_X1 U4359 ( .A1(n3833), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3834), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3474) );
  AOI22_X1 U4360 ( .A1(n3822), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3473) );
  AOI22_X1 U4361 ( .A1(n3750), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3472) );
  AOI22_X1 U4362 ( .A1(n3303), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3471) );
  NAND4_X1 U4363 ( .A1(n3474), .A2(n3473), .A3(n3472), .A4(n3471), .ZN(n3475)
         );
  NOR2_X1 U4364 ( .A1(n3476), .A2(n3475), .ZN(n3481) );
  AOI21_X1 U4365 ( .B1(n6568), .B2(n3478), .A(n3482), .ZN(n5682) );
  OR2_X1 U4366 ( .A1(n5682), .A2(n3876), .ZN(n3480) );
  AOI22_X1 U4367 ( .A1(n4174), .A2(EAX_REG_9__SCAN_IN), .B1(n4173), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3479) );
  OAI211_X1 U4368 ( .C1(n3481), .C2(n3562), .A(n3480), .B(n3479), .ZN(n4678)
         );
  OR2_X1 U4369 ( .A1(n3482), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3483)
         );
  NAND2_X1 U4370 ( .A1(n3483), .A2(n3511), .ZN(n4927) );
  AOI22_X1 U4371 ( .A1(n2975), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3820), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3487) );
  AOI22_X1 U4372 ( .A1(n3834), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3486) );
  AOI22_X1 U4373 ( .A1(n3860), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3485) );
  AOI22_X1 U4374 ( .A1(n3833), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n2972), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3484) );
  NAND4_X1 U4375 ( .A1(n3487), .A2(n3486), .A3(n3485), .A4(n3484), .ZN(n3493)
         );
  AOI22_X1 U4376 ( .A1(n3822), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3303), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3491) );
  AOI22_X1 U4377 ( .A1(n3861), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3490) );
  AOI22_X1 U4378 ( .A1(n3821), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3489) );
  AOI22_X1 U4379 ( .A1(n3750), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3488) );
  NAND4_X1 U4380 ( .A1(n3491), .A2(n3490), .A3(n3489), .A4(n3488), .ZN(n3492)
         );
  OAI21_X1 U4381 ( .B1(n3493), .B2(n3492), .A(n3574), .ZN(n3496) );
  NAND2_X1 U4382 ( .A1(n3434), .A2(EAX_REG_10__SCAN_IN), .ZN(n3495) );
  NAND2_X1 U4383 ( .A1(n4173), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3494)
         );
  NAND3_X1 U4384 ( .A1(n3496), .A2(n3495), .A3(n3494), .ZN(n3497) );
  AOI21_X1 U4385 ( .B1(n4927), .B2(n3870), .A(n3497), .ZN(n4777) );
  AOI22_X1 U4386 ( .A1(n3833), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3501) );
  AOI22_X1 U4387 ( .A1(n3820), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3500) );
  AOI22_X1 U4388 ( .A1(n3834), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3750), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3499) );
  AOI22_X1 U4389 ( .A1(n3303), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3498) );
  NAND4_X1 U4390 ( .A1(n3501), .A2(n3500), .A3(n3499), .A4(n3498), .ZN(n3507)
         );
  AOI22_X1 U4391 ( .A1(n3861), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3821), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3505) );
  AOI22_X1 U4392 ( .A1(n3860), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3504) );
  AOI22_X1 U4393 ( .A1(n2975), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n2972), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3503) );
  AOI22_X1 U4394 ( .A1(n3731), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3502) );
  NAND4_X1 U4395 ( .A1(n3505), .A2(n3504), .A3(n3503), .A4(n3502), .ZN(n3506)
         );
  OAI21_X1 U4396 ( .B1(n3507), .B2(n3506), .A(n3574), .ZN(n3510) );
  XOR2_X1 U4397 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3511), .Z(n5811) );
  AOI22_X1 U4398 ( .A1(n4173), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .B1(n3870), 
        .B2(n5811), .ZN(n3509) );
  NAND2_X1 U4399 ( .A1(n3434), .A2(EAX_REG_11__SCAN_IN), .ZN(n3508) );
  XNOR2_X1 U4400 ( .A(n3529), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4948)
         );
  INV_X1 U4401 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3512) );
  AOI21_X1 U4402 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n3512), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3515) );
  AND2_X1 U4403 ( .A1(n3434), .A2(EAX_REG_12__SCAN_IN), .ZN(n3514) );
  OAI22_X1 U4404 ( .A1(n4948), .A2(n3876), .B1(n3515), .B2(n3514), .ZN(n3527)
         );
  AOI22_X1 U4405 ( .A1(n3821), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3519) );
  AOI22_X1 U4406 ( .A1(n2975), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3518) );
  AOI22_X1 U4407 ( .A1(n3834), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3517) );
  AOI22_X1 U4408 ( .A1(n3303), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3516) );
  NAND4_X1 U4409 ( .A1(n3519), .A2(n3518), .A3(n3517), .A4(n3516), .ZN(n3525)
         );
  AOI22_X1 U4410 ( .A1(n3833), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3523) );
  AOI22_X1 U4411 ( .A1(n3861), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3522) );
  AOI22_X1 U4412 ( .A1(n3750), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3521) );
  AOI22_X1 U4413 ( .A1(n3822), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3520) );
  NAND4_X1 U4414 ( .A1(n3523), .A2(n3522), .A3(n3521), .A4(n3520), .ZN(n3524)
         );
  OAI21_X1 U4415 ( .B1(n3525), .B2(n3524), .A(n3574), .ZN(n3526) );
  NAND2_X1 U4416 ( .A1(n4174), .A2(EAX_REG_13__SCAN_IN), .ZN(n3532) );
  OAI21_X1 U4417 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3530), .A(n3563), 
        .ZN(n5662) );
  AOI22_X1 U4418 ( .A1(n3870), .A2(n5662), .B1(n4173), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3531) );
  NAND2_X1 U4419 ( .A1(n3532), .A2(n3531), .ZN(n3533) );
  OAI21_X1 U4420 ( .B1(n3534), .B2(n3533), .A(n3548), .ZN(n4932) );
  INV_X1 U4421 ( .A(n4932), .ZN(n3547) );
  AOI22_X1 U4422 ( .A1(n3861), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3833), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3538) );
  AOI22_X1 U4423 ( .A1(n2975), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4424 ( .A1(n3822), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3821), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3536) );
  AOI22_X1 U4425 ( .A1(n3303), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3535) );
  NAND4_X1 U4426 ( .A1(n3538), .A2(n3537), .A3(n3536), .A4(n3535), .ZN(n3544)
         );
  AOI22_X1 U4427 ( .A1(n3834), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4428 ( .A1(n3860), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4429 ( .A1(n3820), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n2972), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4430 ( .A1(n3750), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3539) );
  NAND4_X1 U4431 ( .A1(n3542), .A2(n3541), .A3(n3540), .A4(n3539), .ZN(n3543)
         );
  OR2_X1 U4432 ( .A1(n3544), .A2(n3543), .ZN(n3545) );
  NAND2_X1 U4433 ( .A1(n3574), .A2(n3545), .ZN(n4933) );
  NAND2_X1 U4434 ( .A1(n3547), .A2(n3546), .ZN(n4935) );
  AOI22_X1 U4435 ( .A1(n3861), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3552) );
  AOI22_X1 U4436 ( .A1(n3833), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3551) );
  AOI22_X1 U4437 ( .A1(n3280), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4438 ( .A1(n3731), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3549) );
  NAND4_X1 U4439 ( .A1(n3552), .A2(n3551), .A3(n3550), .A4(n3549), .ZN(n3558)
         );
  AOI22_X1 U4440 ( .A1(n2975), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3820), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3556) );
  AOI22_X1 U4441 ( .A1(n3834), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3750), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3555) );
  AOI22_X1 U4442 ( .A1(n3860), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4443 ( .A1(n3821), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n2972), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3553) );
  NAND4_X1 U4444 ( .A1(n3556), .A2(n3555), .A3(n3554), .A4(n3553), .ZN(n3557)
         );
  NOR2_X1 U4445 ( .A1(n3558), .A2(n3557), .ZN(n3561) );
  XNOR2_X1 U4446 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3563), .ZN(n5648)
         );
  INV_X1 U4447 ( .A(n5648), .ZN(n5353) );
  AOI22_X1 U4448 ( .A1(n4173), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n3870), 
        .B2(n5353), .ZN(n3560) );
  NAND2_X1 U4449 ( .A1(n4174), .A2(EAX_REG_14__SCAN_IN), .ZN(n3559) );
  OAI211_X1 U4450 ( .C1(n3562), .C2(n3561), .A(n3560), .B(n3559), .ZN(n5217)
         );
  NAND2_X1 U4451 ( .A1(n5216), .A2(n5217), .ZN(n5133) );
  INV_X1 U4452 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3565) );
  XNOR2_X1 U4453 ( .A(n3581), .B(n3565), .ZN(n5343) );
  AOI22_X1 U4454 ( .A1(n3861), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3821), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3569) );
  AOI22_X1 U4455 ( .A1(n2974), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3568) );
  AOI22_X1 U4456 ( .A1(n3833), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n2972), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3567) );
  AOI22_X1 U4457 ( .A1(n3860), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3566) );
  NAND4_X1 U4458 ( .A1(n3569), .A2(n3568), .A3(n3567), .A4(n3566), .ZN(n3576)
         );
  AOI22_X1 U4459 ( .A1(n3137), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3573) );
  AOI22_X1 U4460 ( .A1(n3822), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3303), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3572) );
  AOI22_X1 U4461 ( .A1(n3820), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3571) );
  AOI22_X1 U4462 ( .A1(n3750), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3570) );
  NAND4_X1 U4463 ( .A1(n3573), .A2(n3572), .A3(n3571), .A4(n3570), .ZN(n3575)
         );
  OAI21_X1 U4464 ( .B1(n3576), .B2(n3575), .A(n3574), .ZN(n3579) );
  NAND2_X1 U4465 ( .A1(n4174), .A2(EAX_REG_15__SCAN_IN), .ZN(n3578) );
  NAND2_X1 U4466 ( .A1(n4173), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3577)
         );
  NAND3_X1 U4467 ( .A1(n3579), .A2(n3578), .A3(n3577), .ZN(n3580) );
  AOI21_X1 U4468 ( .B1(n5343), .B2(n3870), .A(n3580), .ZN(n5134) );
  XOR2_X1 U4469 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3595), .Z(n5641) );
  AOI22_X1 U4470 ( .A1(n4174), .A2(EAX_REG_16__SCAN_IN), .B1(n4173), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3594) );
  AOI22_X1 U4471 ( .A1(n2953), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3750), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4472 ( .A1(n3821), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n2972), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3584) );
  AOI22_X1 U4473 ( .A1(n3860), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3583) );
  AOI22_X1 U4474 ( .A1(n3822), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3582) );
  NAND4_X1 U4475 ( .A1(n3585), .A2(n3584), .A3(n3583), .A4(n3582), .ZN(n3592)
         );
  AOI22_X1 U4476 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n3861), .B1(n3303), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3589) );
  AOI22_X1 U4477 ( .A1(n3833), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3820), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3588) );
  AOI22_X1 U4478 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n2975), .B1(n3731), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4479 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n3834), .B1(n3158), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3586) );
  NAND4_X1 U4480 ( .A1(n3589), .A2(n3588), .A3(n3587), .A4(n3586), .ZN(n3591)
         );
  NAND2_X1 U4481 ( .A1(n3187), .A2(n4501), .ZN(n3590) );
  OAI21_X1 U4482 ( .B1(n3592), .B2(n3591), .A(n3847), .ZN(n3593) );
  OAI211_X1 U4483 ( .C1(n5641), .C2(n3876), .A(n3594), .B(n3593), .ZN(n5205)
         );
  NAND2_X1 U4484 ( .A1(n5135), .A2(n5205), .ZN(n5120) );
  INV_X1 U4485 ( .A(n5120), .ZN(n3612) );
  XNOR2_X1 U4486 ( .A(n3613), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5557)
         );
  NAND2_X1 U4487 ( .A1(n5557), .A2(n3870), .ZN(n3610) );
  AOI22_X1 U4488 ( .A1(n2976), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3820), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3599) );
  AOI22_X1 U4489 ( .A1(n3137), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4490 ( .A1(n3861), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4491 ( .A1(n3822), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3596) );
  NAND4_X1 U4492 ( .A1(n3599), .A2(n3598), .A3(n3597), .A4(n3596), .ZN(n3605)
         );
  AOI22_X1 U4493 ( .A1(n3833), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3603) );
  AOI22_X1 U4494 ( .A1(n3821), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3602) );
  AOI22_X1 U4495 ( .A1(n3750), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3601) );
  AOI22_X1 U4496 ( .A1(n3303), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3600) );
  NAND4_X1 U4497 ( .A1(n3603), .A2(n3602), .A3(n3601), .A4(n3600), .ZN(n3604)
         );
  NOR2_X1 U4498 ( .A1(n3605), .A2(n3604), .ZN(n3608) );
  AOI21_X1 U4499 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5124), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3606) );
  AOI21_X1 U4500 ( .B1(n3434), .B2(EAX_REG_17__SCAN_IN), .A(n3606), .ZN(n3607)
         );
  OAI21_X1 U4501 ( .B1(n3873), .B2(n3608), .A(n3607), .ZN(n3609) );
  NAND2_X1 U4502 ( .A1(n3610), .A2(n3609), .ZN(n5122) );
  NAND2_X1 U4503 ( .A1(n3612), .A2(n3611), .ZN(n5194) );
  INV_X1 U4504 ( .A(n5194), .ZN(n3633) );
  INV_X1 U4505 ( .A(n3651), .ZN(n3616) );
  OR2_X1 U4506 ( .A1(n3614), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3615)
         );
  NAND2_X1 U4507 ( .A1(n3616), .A2(n3615), .ZN(n5632) );
  AOI22_X1 U4508 ( .A1(n3833), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3820), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4509 ( .A1(n3834), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3750), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3619) );
  AOI22_X1 U4510 ( .A1(n3280), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4511 ( .A1(n3861), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3617) );
  NAND4_X1 U4512 ( .A1(n3620), .A2(n3619), .A3(n3618), .A4(n3617), .ZN(n3626)
         );
  AOI22_X1 U4513 ( .A1(n2975), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4514 ( .A1(n3821), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3623) );
  AOI22_X1 U4515 ( .A1(n3822), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4516 ( .A1(n3731), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3621) );
  NAND4_X1 U4517 ( .A1(n3624), .A2(n3623), .A3(n3622), .A4(n3621), .ZN(n3625)
         );
  NOR2_X1 U4518 ( .A1(n3626), .A2(n3625), .ZN(n3627) );
  NOR2_X1 U4519 ( .A1(n3873), .A2(n3627), .ZN(n3631) );
  INV_X1 U4520 ( .A(EAX_REG_18__SCAN_IN), .ZN(n3629) );
  NAND2_X1 U4521 ( .A1(n6442), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3628)
         );
  OAI211_X1 U4522 ( .C1(n3513), .C2(n3629), .A(n3876), .B(n3628), .ZN(n3630)
         );
  OAI22_X1 U4523 ( .A1(n5632), .A2(n3876), .B1(n3631), .B2(n3630), .ZN(n5195)
         );
  NAND2_X1 U4524 ( .A1(n3633), .A2(n3632), .ZN(n5185) );
  INV_X1 U4525 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3634) );
  XNOR2_X1 U4526 ( .A(n3651), .B(n3634), .ZN(n5528) );
  NAND2_X1 U4527 ( .A1(n5528), .A2(n3870), .ZN(n3650) );
  AOI22_X1 U4528 ( .A1(n3833), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3638) );
  AOI22_X1 U4529 ( .A1(n2976), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3820), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3637) );
  AOI22_X1 U4530 ( .A1(n2953), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3636) );
  AOI22_X1 U4531 ( .A1(n3750), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3635) );
  NAND4_X1 U4532 ( .A1(n3638), .A2(n3637), .A3(n3636), .A4(n3635), .ZN(n3644)
         );
  AOI22_X1 U4533 ( .A1(n3861), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3821), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4534 ( .A1(n3834), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4535 ( .A1(n3822), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4536 ( .A1(n3280), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3639) );
  NAND4_X1 U4537 ( .A1(n3642), .A2(n3641), .A3(n3640), .A4(n3639), .ZN(n3643)
         );
  NOR2_X1 U4538 ( .A1(n3644), .A2(n3643), .ZN(n3648) );
  NAND2_X1 U4539 ( .A1(n6442), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3645)
         );
  NAND2_X1 U4540 ( .A1(n3876), .A2(n3645), .ZN(n3646) );
  AOI21_X1 U4541 ( .B1(n3434), .B2(EAX_REG_19__SCAN_IN), .A(n3646), .ZN(n3647)
         );
  OAI21_X1 U4542 ( .B1(n3873), .B2(n3648), .A(n3647), .ZN(n3649) );
  NAND2_X1 U4543 ( .A1(n3650), .A2(n3649), .ZN(n5187) );
  INV_X1 U4544 ( .A(n3653), .ZN(n3652) );
  INV_X1 U4545 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U4546 ( .A1(n3652), .A2(n5322), .ZN(n3654) );
  AND2_X1 U4547 ( .A1(n3654), .A2(n3698), .ZN(n5514) );
  AOI22_X1 U4548 ( .A1(n3861), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4549 ( .A1(n2975), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3137), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3657) );
  AOI22_X1 U4550 ( .A1(n3833), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4551 ( .A1(n3750), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3655) );
  NAND4_X1 U4552 ( .A1(n3658), .A2(n3657), .A3(n3656), .A4(n3655), .ZN(n3664)
         );
  AOI22_X1 U4553 ( .A1(n2953), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U4554 ( .A1(n3821), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3661) );
  AOI22_X1 U4555 ( .A1(n3860), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3660) );
  AOI22_X1 U4556 ( .A1(n3303), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3659) );
  NAND4_X1 U4557 ( .A1(n3662), .A2(n3661), .A3(n3660), .A4(n3659), .ZN(n3663)
         );
  OR2_X1 U4558 ( .A1(n3664), .A2(n3663), .ZN(n3667) );
  INV_X1 U4559 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4386) );
  OAI21_X1 U4560 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6455), .A(n6442), 
        .ZN(n3665) );
  OAI21_X1 U4561 ( .B1(n3513), .B2(n4386), .A(n3665), .ZN(n3666) );
  AOI21_X1 U4562 ( .B1(n3847), .B2(n3667), .A(n3666), .ZN(n3668) );
  AOI21_X1 U4563 ( .B1(n5514), .B2(n3870), .A(n3668), .ZN(n5179) );
  NAND2_X1 U4564 ( .A1(n5178), .A2(n5179), .ZN(n5112) );
  AOI22_X1 U4565 ( .A1(n3822), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4566 ( .A1(n3820), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3750), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4567 ( .A1(n3861), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3821), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4568 ( .A1(n3833), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n2972), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3669) );
  NAND4_X1 U4569 ( .A1(n3672), .A2(n3671), .A3(n3670), .A4(n3669), .ZN(n3678)
         );
  AOI22_X1 U4570 ( .A1(n2974), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3676) );
  AOI22_X1 U4571 ( .A1(n2953), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3675) );
  AOI22_X1 U4572 ( .A1(n3305), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3674) );
  AOI22_X1 U4573 ( .A1(n3137), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3673) );
  NAND4_X1 U4574 ( .A1(n3676), .A2(n3675), .A3(n3674), .A4(n3673), .ZN(n3677)
         );
  NOR2_X1 U4575 ( .A1(n3678), .A2(n3677), .ZN(n3681) );
  INV_X1 U4576 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5314) );
  OAI21_X1 U4577 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5314), .A(n3876), .ZN(
        n3679) );
  AOI21_X1 U4578 ( .B1(n3434), .B2(EAX_REG_21__SCAN_IN), .A(n3679), .ZN(n3680)
         );
  OAI21_X1 U4579 ( .B1(n3873), .B2(n3681), .A(n3680), .ZN(n3683) );
  XNOR2_X1 U4580 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n3698), .ZN(n5316)
         );
  NAND2_X1 U4581 ( .A1(n3870), .A2(n5316), .ZN(n3682) );
  NAND2_X1 U4582 ( .A1(n3683), .A2(n3682), .ZN(n5168) );
  AOI22_X1 U4583 ( .A1(n3820), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4584 ( .A1(n3137), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3750), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4585 ( .A1(n3822), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3303), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4586 ( .A1(n3833), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3684) );
  NAND4_X1 U4587 ( .A1(n3687), .A2(n3686), .A3(n3685), .A4(n3684), .ZN(n3693)
         );
  AOI22_X1 U4588 ( .A1(n3861), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3821), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4589 ( .A1(n2975), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4590 ( .A1(n3731), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4591 ( .A1(n3860), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3688) );
  NAND4_X1 U4592 ( .A1(n3691), .A2(n3690), .A3(n3689), .A4(n3688), .ZN(n3692)
         );
  NOR2_X1 U4593 ( .A1(n3693), .A2(n3692), .ZN(n3697) );
  OAI21_X1 U4594 ( .B1(PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6455), .A(n6442), 
        .ZN(n3694) );
  INV_X1 U4595 ( .A(n3694), .ZN(n3695) );
  AOI21_X1 U4596 ( .B1(n3434), .B2(EAX_REG_22__SCAN_IN), .A(n3695), .ZN(n3696)
         );
  OAI21_X1 U4597 ( .B1(n3873), .B2(n3697), .A(n3696), .ZN(n3702) );
  OAI21_X1 U4598 ( .B1(n3700), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n3744), 
        .ZN(n5513) );
  OR2_X1 U4599 ( .A1(n5513), .A2(n3876), .ZN(n3701) );
  NAND2_X1 U4600 ( .A1(n3702), .A2(n3701), .ZN(n5167) );
  AOI22_X1 U4601 ( .A1(n3833), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3820), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4602 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n2976), .B1(n2953), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4603 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n3834), .B1(n3731), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4604 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n3750), .B1(n3158), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3703) );
  NAND4_X1 U4605 ( .A1(n3706), .A2(n3705), .A3(n3704), .A4(n3703), .ZN(n3712)
         );
  AOI22_X1 U4606 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n3860), .B1(n3821), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4607 ( .A1(n3861), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3709) );
  AOI22_X1 U4608 ( .A1(n3822), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3708) );
  AOI22_X1 U4609 ( .A1(n3303), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3707) );
  NAND4_X1 U4610 ( .A1(n3710), .A2(n3709), .A3(n3708), .A4(n3707), .ZN(n3711)
         );
  OR2_X1 U4611 ( .A1(n3712), .A2(n3711), .ZN(n3730) );
  AOI22_X1 U4612 ( .A1(n3833), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3820), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4613 ( .A1(n2975), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3715) );
  AOI22_X1 U4614 ( .A1(n3834), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3714) );
  AOI22_X1 U4615 ( .A1(n3750), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3713) );
  NAND4_X1 U4616 ( .A1(n3716), .A2(n3715), .A3(n3714), .A4(n3713), .ZN(n3722)
         );
  AOI22_X1 U4617 ( .A1(n3821), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4618 ( .A1(n3861), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n2972), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4619 ( .A1(n3822), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4620 ( .A1(n3303), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3717) );
  NAND4_X1 U4621 ( .A1(n3720), .A2(n3719), .A3(n3718), .A4(n3717), .ZN(n3721)
         );
  OR2_X1 U4622 ( .A1(n3722), .A2(n3721), .ZN(n3729) );
  XNOR2_X1 U4623 ( .A(n3730), .B(n3729), .ZN(n3726) );
  NAND2_X1 U4624 ( .A1(n6442), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3723)
         );
  NAND2_X1 U4625 ( .A1(n3876), .A2(n3723), .ZN(n3724) );
  AOI21_X1 U4626 ( .B1(n3434), .B2(EAX_REG_23__SCAN_IN), .A(n3724), .ZN(n3725)
         );
  OAI21_X1 U4627 ( .B1(n3873), .B2(n3726), .A(n3725), .ZN(n3728) );
  XNOR2_X1 U4628 ( .A(n3744), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5493)
         );
  NAND2_X1 U4629 ( .A1(n5493), .A2(n3870), .ZN(n3727) );
  NAND2_X1 U4630 ( .A1(n3728), .A2(n3727), .ZN(n5160) );
  NAND2_X1 U4631 ( .A1(n3730), .A2(n3729), .ZN(n3761) );
  INV_X1 U4632 ( .A(n3761), .ZN(n3742) );
  AOI22_X1 U4633 ( .A1(n3833), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3820), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4634 ( .A1(n2976), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3734) );
  AOI22_X1 U4635 ( .A1(n3834), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3733) );
  AOI22_X1 U4636 ( .A1(n3750), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3732) );
  NAND4_X1 U4637 ( .A1(n3735), .A2(n3734), .A3(n3733), .A4(n3732), .ZN(n3741)
         );
  AOI22_X1 U4638 ( .A1(n3821), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4639 ( .A1(n3861), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4640 ( .A1(n3822), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4641 ( .A1(n3280), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3736) );
  NAND4_X1 U4642 ( .A1(n3739), .A2(n3738), .A3(n3737), .A4(n3736), .ZN(n3740)
         );
  NOR2_X1 U4643 ( .A1(n3741), .A2(n3740), .ZN(n3762) );
  XNOR2_X1 U4644 ( .A(n3742), .B(n3762), .ZN(n3743) );
  NAND2_X1 U4645 ( .A1(n3847), .A2(n3743), .ZN(n3749) );
  INV_X1 U4646 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5502) );
  INV_X1 U4647 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5492) );
  XNOR2_X1 U4648 ( .A(n3767), .B(n5492), .ZN(n5485) );
  NOR2_X1 U4649 ( .A1(n5485), .A2(n3876), .ZN(n3747) );
  NOR2_X1 U4650 ( .A1(n3745), .A2(n5492), .ZN(n3746) );
  AOI211_X1 U4651 ( .C1(n3434), .C2(EAX_REG_24__SCAN_IN), .A(n3747), .B(n3746), 
        .ZN(n3748) );
  NAND2_X1 U4652 ( .A1(n3749), .A2(n3748), .ZN(n5154) );
  AOI22_X1 U4653 ( .A1(n3833), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3820), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3754) );
  AOI22_X1 U4654 ( .A1(n2976), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4655 ( .A1(n3834), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4656 ( .A1(n3750), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3751) );
  NAND4_X1 U4657 ( .A1(n3754), .A2(n3753), .A3(n3752), .A4(n3751), .ZN(n3760)
         );
  AOI22_X1 U4658 ( .A1(n3821), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3758) );
  AOI22_X1 U4659 ( .A1(n3861), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n2972), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4660 ( .A1(n3822), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4661 ( .A1(n3303), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3755) );
  NAND4_X1 U4662 ( .A1(n3758), .A2(n3757), .A3(n3756), .A4(n3755), .ZN(n3759)
         );
  OR2_X1 U4663 ( .A1(n3760), .A2(n3759), .ZN(n3775) );
  NOR2_X1 U4664 ( .A1(n3762), .A2(n3761), .ZN(n3776) );
  XNOR2_X1 U4665 ( .A(n3775), .B(n3776), .ZN(n3766) );
  INV_X1 U4666 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3763) );
  AOI21_X1 U4667 ( .B1(n3763), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3764) );
  AOI21_X1 U4668 ( .B1(n3434), .B2(EAX_REG_25__SCAN_IN), .A(n3764), .ZN(n3765)
         );
  OAI21_X1 U4669 ( .B1(n3873), .B2(n3766), .A(n3765), .ZN(n3769) );
  NAND2_X1 U4670 ( .A1(n3767), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3770)
         );
  XNOR2_X1 U4671 ( .A(n3770), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5477)
         );
  NAND2_X1 U4672 ( .A1(n5477), .A2(n3870), .ZN(n3768) );
  NAND2_X1 U4673 ( .A1(n5146), .A2(n5147), .ZN(n5100) );
  INV_X1 U4674 ( .A(n3770), .ZN(n3771) );
  INV_X1 U4675 ( .A(n3772), .ZN(n3773) );
  INV_X1 U4676 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5102) );
  NAND2_X1 U4677 ( .A1(n3773), .A2(n5102), .ZN(n3774) );
  NAND2_X1 U4678 ( .A1(n3807), .A2(n3774), .ZN(n5273) );
  NAND2_X1 U4679 ( .A1(n3776), .A2(n3775), .ZN(n3801) );
  AOI22_X1 U4680 ( .A1(n3861), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3820), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4681 ( .A1(n3821), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4682 ( .A1(n3822), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4683 ( .A1(n2953), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3777) );
  NAND4_X1 U4684 ( .A1(n3780), .A2(n3779), .A3(n3778), .A4(n3777), .ZN(n3786)
         );
  AOI22_X1 U4685 ( .A1(n3137), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3750), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4686 ( .A1(n2976), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4687 ( .A1(n3833), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n2972), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4688 ( .A1(n3280), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3781) );
  NAND4_X1 U4689 ( .A1(n3784), .A2(n3783), .A3(n3782), .A4(n3781), .ZN(n3785)
         );
  NOR2_X1 U4690 ( .A1(n3786), .A2(n3785), .ZN(n3802) );
  XNOR2_X1 U4691 ( .A(n3801), .B(n3802), .ZN(n3789) );
  AOI21_X1 U4692 ( .B1(PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6442), .A(n3870), 
        .ZN(n3788) );
  NAND2_X1 U4693 ( .A1(n4174), .A2(EAX_REG_26__SCAN_IN), .ZN(n3787) );
  OAI211_X1 U4694 ( .C1(n3789), .C2(n3873), .A(n3788), .B(n3787), .ZN(n3790)
         );
  NOR2_X2 U4695 ( .A1(n5100), .A2(n5101), .ZN(n5085) );
  AOI22_X1 U4696 ( .A1(n3833), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3820), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4697 ( .A1(n2976), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4698 ( .A1(n3834), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4699 ( .A1(n3750), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3791) );
  NAND4_X1 U4700 ( .A1(n3794), .A2(n3793), .A3(n3792), .A4(n3791), .ZN(n3800)
         );
  AOI22_X1 U4701 ( .A1(n3821), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4702 ( .A1(n3861), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n2972), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4703 ( .A1(n3822), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4704 ( .A1(n3280), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3795) );
  NAND4_X1 U4705 ( .A1(n3798), .A2(n3797), .A3(n3796), .A4(n3795), .ZN(n3799)
         );
  OR2_X1 U4706 ( .A1(n3800), .A2(n3799), .ZN(n3813) );
  NOR2_X1 U4707 ( .A1(n3802), .A2(n3801), .ZN(n3814) );
  XOR2_X1 U4708 ( .A(n3813), .B(n3814), .Z(n3803) );
  NAND2_X1 U4709 ( .A1(n3803), .A2(n3847), .ZN(n3806) );
  INV_X1 U4710 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5089) );
  NOR2_X1 U4711 ( .A1(n5089), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3804) );
  AOI211_X1 U4712 ( .C1(n3434), .C2(EAX_REG_27__SCAN_IN), .A(n3870), .B(n3804), 
        .ZN(n3805) );
  XNOR2_X1 U4713 ( .A(n3807), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5088)
         );
  AOI22_X1 U4714 ( .A1(n3806), .A2(n3805), .B1(n3870), .B2(n5088), .ZN(n5087)
         );
  INV_X1 U4715 ( .A(n3807), .ZN(n3808) );
  INV_X1 U4716 ( .A(n3809), .ZN(n3811) );
  INV_X1 U4717 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3810) );
  NAND2_X1 U4718 ( .A1(n3811), .A2(n3810), .ZN(n3812) );
  NAND2_X1 U4719 ( .A1(n3852), .A2(n3812), .ZN(n5257) );
  NAND2_X1 U4720 ( .A1(n3814), .A2(n3813), .ZN(n3845) );
  AOI22_X1 U4721 ( .A1(n3860), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4722 ( .A1(n2953), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n2972), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4723 ( .A1(n3731), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4724 ( .A1(n3303), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3816) );
  NAND4_X1 U4725 ( .A1(n3819), .A2(n3818), .A3(n3817), .A4(n3816), .ZN(n3828)
         );
  AOI22_X1 U4726 ( .A1(n3833), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3861), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4727 ( .A1(n2976), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3820), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4728 ( .A1(n3137), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3750), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4729 ( .A1(n3822), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3821), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3823) );
  NAND4_X1 U4730 ( .A1(n3826), .A2(n3825), .A3(n3824), .A4(n3823), .ZN(n3827)
         );
  NOR2_X1 U4731 ( .A1(n3828), .A2(n3827), .ZN(n3846) );
  XNOR2_X1 U4732 ( .A(n3845), .B(n3846), .ZN(n3831) );
  AOI21_X1 U4733 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6442), .A(n3870), 
        .ZN(n3830) );
  NAND2_X1 U4734 ( .A1(n4174), .A2(EAX_REG_28__SCAN_IN), .ZN(n3829) );
  OAI211_X1 U4735 ( .C1(n3831), .C2(n3873), .A(n3830), .B(n3829), .ZN(n3832)
         );
  OAI21_X1 U4736 ( .B1(n3876), .B2(n5257), .A(n3832), .ZN(n5075) );
  AOI22_X1 U4737 ( .A1(n3833), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4738 ( .A1(n2975), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4739 ( .A1(n3834), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4740 ( .A1(n3750), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3835) );
  NAND4_X1 U4741 ( .A1(n3838), .A2(n3837), .A3(n3836), .A4(n3835), .ZN(n3844)
         );
  AOI22_X1 U4742 ( .A1(n3821), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4743 ( .A1(n3861), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4744 ( .A1(n3822), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4745 ( .A1(n3303), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3839) );
  NAND4_X1 U4746 ( .A1(n3842), .A2(n3841), .A3(n3840), .A4(n3839), .ZN(n3843)
         );
  OR2_X1 U4747 ( .A1(n3844), .A2(n3843), .ZN(n3853) );
  NOR2_X1 U4748 ( .A1(n3846), .A2(n3845), .ZN(n3854) );
  XOR2_X1 U4749 ( .A(n3853), .B(n3854), .Z(n3848) );
  NAND2_X1 U4750 ( .A1(n3848), .A2(n3847), .ZN(n3851) );
  INV_X1 U4751 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4169) );
  AOI21_X1 U4752 ( .B1(n4169), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3849) );
  AOI21_X1 U4753 ( .B1(n3434), .B2(EAX_REG_29__SCAN_IN), .A(n3849), .ZN(n3850)
         );
  XNOR2_X1 U4754 ( .A(n3852), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5023)
         );
  XNOR2_X1 U4755 ( .A(n4188), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5064)
         );
  NAND2_X1 U4756 ( .A1(n3854), .A2(n3853), .ZN(n3869) );
  AOI22_X1 U4757 ( .A1(n2953), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3731), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4758 ( .A1(n2972), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4759 ( .A1(n3137), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4760 ( .A1(n3822), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3856) );
  NAND4_X1 U4761 ( .A1(n3859), .A2(n3858), .A3(n3857), .A4(n3856), .ZN(n3867)
         );
  AOI22_X1 U4762 ( .A1(n3280), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4763 ( .A1(n3152), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4764 ( .A1(n2976), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3750), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4765 ( .A1(n3861), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3821), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3862) );
  NAND4_X1 U4766 ( .A1(n3865), .A2(n3864), .A3(n3863), .A4(n3862), .ZN(n3866)
         );
  NOR2_X1 U4767 ( .A1(n3867), .A2(n3866), .ZN(n3868) );
  XNOR2_X1 U4768 ( .A(n3869), .B(n3868), .ZN(n3874) );
  AOI21_X1 U4769 ( .B1(PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6442), .A(n3870), 
        .ZN(n3872) );
  NAND2_X1 U4770 ( .A1(n4174), .A2(EAX_REG_30__SCAN_IN), .ZN(n3871) );
  OAI211_X1 U4771 ( .C1(n3874), .C2(n3873), .A(n3872), .B(n3871), .ZN(n3875)
         );
  AOI21_X1 U4772 ( .B1(n3877), .B2(n3878), .A(n4176), .ZN(n5010) );
  INV_X1 U4773 ( .A(n5010), .ZN(n5235) );
  INV_X1 U4774 ( .A(n3188), .ZN(n3880) );
  NAND2_X2 U4775 ( .A1(n4517), .A2(n3188), .ZN(n3969) );
  NAND2_X1 U4776 ( .A1(n3192), .A2(n4517), .ZN(n4753) );
  OR2_X1 U4777 ( .A1(n4753), .A2(n4527), .ZN(n4442) );
  OAI21_X1 U4778 ( .B1(n5019), .B2(n4290), .A(n4442), .ZN(n3881) );
  AOI21_X1 U4779 ( .B1(n3879), .B2(n4303), .A(n3881), .ZN(n3886) );
  NAND3_X1 U4780 ( .A1(n3882), .A2(n4715), .A3(n3205), .ZN(n3885) );
  INV_X1 U4781 ( .A(n3205), .ZN(n3883) );
  NAND2_X1 U4782 ( .A1(n3883), .A2(n2954), .ZN(n3884) );
  AND2_X1 U4783 ( .A1(n3885), .A2(n3884), .ZN(n4276) );
  AND2_X1 U4784 ( .A1(n3886), .A2(n4276), .ZN(n3887) );
  NAND2_X1 U4785 ( .A1(n3888), .A2(n3887), .ZN(n4418) );
  INV_X1 U4786 ( .A(n4450), .ZN(n3889) );
  NOR2_X1 U4787 ( .A1(n4976), .A2(n4249), .ZN(n4280) );
  NAND2_X1 U4788 ( .A1(n4298), .A2(n4280), .ZN(n4424) );
  XNOR2_X1 U4789 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3911) );
  NAND2_X1 U4790 ( .A1(n3912), .A2(n3911), .ZN(n3891) );
  NAND2_X1 U4791 ( .A1(n6301), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3890) );
  NAND2_X1 U4792 ( .A1(n3891), .A2(n3890), .ZN(n3908) );
  XNOR2_X1 U4793 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3906) );
  NAND2_X1 U4794 ( .A1(n3908), .A2(n3906), .ZN(n3893) );
  NAND2_X1 U4795 ( .A1(n6305), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3892) );
  NAND2_X1 U4796 ( .A1(n3893), .A2(n3892), .ZN(n3900) );
  XNOR2_X1 U4797 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3898) );
  NAND2_X1 U4798 ( .A1(n3900), .A2(n3898), .ZN(n3895) );
  NAND2_X1 U4799 ( .A1(n6313), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3894) );
  NAND2_X1 U4800 ( .A1(n3895), .A2(n3894), .ZN(n3902) );
  NAND2_X1 U4801 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4460), .ZN(n3901) );
  NAND2_X1 U4802 ( .A1(n3919), .A2(n3938), .ZN(n3937) );
  INV_X1 U4803 ( .A(n3898), .ZN(n3899) );
  XNOR2_X1 U4804 ( .A(n3900), .B(n3899), .ZN(n4180) );
  INV_X1 U4805 ( .A(n4180), .ZN(n3903) );
  NOR2_X1 U4806 ( .A1(n3902), .A2(n3901), .ZN(n4183) );
  INV_X1 U4807 ( .A(n3930), .ZN(n3934) );
  INV_X1 U4808 ( .A(n3906), .ZN(n3907) );
  XNOR2_X1 U4809 ( .A(n3908), .B(n3907), .ZN(n4181) );
  NAND2_X1 U4810 ( .A1(n3919), .A2(n4181), .ZN(n3910) );
  INV_X1 U4811 ( .A(n3910), .ZN(n3929) );
  AND2_X1 U4812 ( .A1(n4249), .A2(n3193), .ZN(n3909) );
  INV_X1 U4813 ( .A(n3915), .ZN(n3928) );
  OAI211_X1 U4814 ( .C1(n4181), .C2(n3931), .A(n3915), .B(n3910), .ZN(n3927)
         );
  AOI21_X1 U4815 ( .B1(n3919), .B2(n4517), .A(n3176), .ZN(n3925) );
  XOR2_X1 U4816 ( .A(n3912), .B(n3911), .Z(n4182) );
  NAND2_X1 U4817 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4182), .ZN(n3924) );
  INV_X1 U4818 ( .A(n4182), .ZN(n3917) );
  AND2_X1 U4819 ( .A1(n3194), .A2(n3193), .ZN(n4159) );
  INV_X1 U4820 ( .A(n3912), .ZN(n3913) );
  OAI21_X1 U4821 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6138), .A(n3913), 
        .ZN(n3918) );
  OAI21_X1 U4822 ( .B1(n4159), .B2(n3918), .A(n4715), .ZN(n3914) );
  AOI22_X1 U4823 ( .A1(n3915), .A2(n3914), .B1(n3925), .B2(n3924), .ZN(n3920)
         );
  INV_X1 U4824 ( .A(n3939), .ZN(n3916) );
  OAI21_X1 U4825 ( .B1(n3917), .B2(n3920), .A(n3916), .ZN(n3923) );
  INV_X1 U4826 ( .A(n3918), .ZN(n3921) );
  NAND3_X1 U4827 ( .A1(n3921), .A2(n3920), .A3(n3919), .ZN(n3922) );
  OAI211_X1 U4828 ( .C1(n3925), .C2(n3924), .A(n3923), .B(n3922), .ZN(n3926)
         );
  AOI22_X1 U4829 ( .A1(n3929), .A2(n3928), .B1(n3927), .B2(n3926), .ZN(n3933)
         );
  OAI22_X1 U4830 ( .A1(n3934), .A2(n3939), .B1(n3933), .B2(n3932), .ZN(n3935)
         );
  AOI21_X1 U4831 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n3297), .A(n3935), 
        .ZN(n3936) );
  NAND2_X1 U4832 ( .A1(n3937), .A2(n3936), .ZN(n3941) );
  OR2_X1 U4833 ( .A1(n4424), .A2(n4466), .ZN(n4446) );
  NAND2_X1 U4834 ( .A1(n3194), .A2(n5228), .ZN(n3942) );
  OR2_X1 U4835 ( .A1(n3943), .A2(n3942), .ZN(n4315) );
  INV_X1 U4836 ( .A(n4315), .ZN(n3946) );
  NAND2_X1 U4837 ( .A1(n4715), .A2(n3944), .ZN(n3951) );
  NAND3_X1 U4838 ( .A1(n3946), .A2(n3945), .A3(n4236), .ZN(n3947) );
  NAND2_X1 U4839 ( .A1(n4446), .A2(n3947), .ZN(n3949) );
  INV_X1 U4840 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4402) );
  INV_X1 U4841 ( .A(n4303), .ZN(n3982) );
  INV_X1 U4842 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5903) );
  INV_X1 U4843 ( .A(n4035), .ZN(n3981) );
  AOI22_X1 U4844 ( .A1(n3982), .A2(n5903), .B1(n3981), .B2(n4402), .ZN(n3950)
         );
  OAI21_X1 U4845 ( .B1(n3969), .B2(n4402), .A(n3950), .ZN(n4401) );
  INV_X1 U4846 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3952) );
  NAND2_X1 U4847 ( .A1(n3961), .A2(n3952), .ZN(n3955) );
  OR2_X1 U4848 ( .A1(n4030), .A2(n3952), .ZN(n3954) );
  NAND2_X1 U4849 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4043), .ZN(n3953)
         );
  NAND4_X1 U4850 ( .A1(n3955), .A2(n4009), .A3(n3954), .A4(n3953), .ZN(n3958)
         );
  NAND2_X1 U4851 ( .A1(n4030), .A2(EBX_REG_0__SCAN_IN), .ZN(n3957) );
  INV_X1 U4852 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4752) );
  NAND2_X1 U4853 ( .A1(n3969), .A2(n4752), .ZN(n3956) );
  NOR2_X1 U4854 ( .A1(n5756), .A2(n4043), .ZN(n3960) );
  INV_X1 U4855 ( .A(n3958), .ZN(n3959) );
  INV_X1 U4856 ( .A(EBX_REG_2__SCAN_IN), .ZN(n3962) );
  NAND2_X1 U4857 ( .A1(n3961), .A2(n3962), .ZN(n3965) );
  OR2_X1 U4858 ( .A1(n4030), .A2(n3962), .ZN(n3964) );
  NAND2_X1 U4859 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n4043), .ZN(n3963)
         );
  NAND4_X1 U4860 ( .A1(n3965), .A2(n4009), .A3(n3964), .A4(n3963), .ZN(n4408)
         );
  NAND2_X1 U4861 ( .A1(n4409), .A2(n4408), .ZN(n4410) );
  INV_X1 U4862 ( .A(EBX_REG_4__SCAN_IN), .ZN(n5706) );
  NAND2_X1 U4863 ( .A1(n3961), .A2(n5706), .ZN(n3968) );
  INV_X1 U4864 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U4865 ( .A1(n4030), .A2(n5894), .ZN(n3966) );
  OAI211_X1 U4866 ( .C1(n4043), .C2(EBX_REG_4__SCAN_IN), .A(n3966), .B(n3969), 
        .ZN(n3967) );
  NAND2_X1 U4867 ( .A1(n3968), .A2(n3967), .ZN(n4490) );
  INV_X1 U4868 ( .A(n3969), .ZN(n5181) );
  NAND2_X1 U4869 ( .A1(n5181), .A2(EBX_REG_5__SCAN_IN), .ZN(n3971) );
  OR2_X1 U4870 ( .A1(n4303), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3970)
         );
  OAI211_X1 U4871 ( .C1(n4035), .C2(EBX_REG_5__SCAN_IN), .A(n3971), .B(n3970), 
        .ZN(n4413) );
  INV_X1 U4872 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4550) );
  NAND2_X1 U4873 ( .A1(n3961), .A2(n4550), .ZN(n3974) );
  OR2_X1 U4874 ( .A1(n4030), .A2(n4550), .ZN(n3973) );
  NAND2_X1 U4875 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4043), .ZN(n3972)
         );
  NAND4_X1 U4876 ( .A1(n3974), .A2(n4009), .A3(n3973), .A4(n3972), .ZN(n4548)
         );
  NAND2_X1 U4877 ( .A1(n5181), .A2(EBX_REG_7__SCAN_IN), .ZN(n3976) );
  OR2_X1 U4878 ( .A1(n4303), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3975)
         );
  OAI211_X1 U4879 ( .C1(n4035), .C2(EBX_REG_7__SCAN_IN), .A(n3976), .B(n3975), 
        .ZN(n4618) );
  NOR2_X2 U4880 ( .A1(n4617), .A2(n4618), .ZN(n4670) );
  INV_X1 U4881 ( .A(n3961), .ZN(n3980) );
  INV_X1 U4882 ( .A(n4030), .ZN(n4039) );
  INV_X1 U4883 ( .A(n4009), .ZN(n3977) );
  AOI21_X1 U4884 ( .B1(n4039), .B2(EBX_REG_8__SCAN_IN), .A(n3977), .ZN(n3979)
         );
  NAND2_X1 U4885 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n4043), .ZN(n3978)
         );
  OAI211_X1 U4886 ( .C1(EBX_REG_8__SCAN_IN), .C2(n3980), .A(n3979), .B(n3978), 
        .ZN(n4671) );
  INV_X1 U4887 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4733) );
  INV_X1 U4888 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6461) );
  AOI22_X1 U4889 ( .A1(n3982), .A2(n6461), .B1(n3981), .B2(n4733), .ZN(n3983)
         );
  OAI21_X1 U4890 ( .B1(n3969), .B2(n4733), .A(n3983), .ZN(n4732) );
  INV_X1 U4891 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4789) );
  NAND2_X1 U4892 ( .A1(n3961), .A2(n4789), .ZN(n3986) );
  INV_X1 U4893 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4129) );
  NAND2_X1 U4894 ( .A1(n4030), .A2(n4129), .ZN(n3984) );
  OAI211_X1 U4895 ( .C1(n4043), .C2(EBX_REG_10__SCAN_IN), .A(n3984), .B(n3969), 
        .ZN(n3985) );
  NAND2_X1 U4896 ( .A1(n3986), .A2(n3985), .ZN(n4778) );
  OR2_X1 U4897 ( .A1(n4035), .A2(EBX_REG_11__SCAN_IN), .ZN(n3989) );
  NAND2_X1 U4898 ( .A1(n3969), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3987) );
  OAI211_X1 U4899 ( .C1(n3951), .C2(EBX_REG_11__SCAN_IN), .A(n4030), .B(n3987), 
        .ZN(n3988) );
  NAND2_X1 U4900 ( .A1(n3989), .A2(n3988), .ZN(n5667) );
  INV_X1 U4901 ( .A(EBX_REG_12__SCAN_IN), .ZN(n4878) );
  NAND2_X1 U4902 ( .A1(n3961), .A2(n4878), .ZN(n3992) );
  INV_X1 U4903 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4968) );
  NAND2_X1 U4904 ( .A1(n4030), .A2(n4968), .ZN(n3990) );
  OAI211_X1 U4905 ( .C1(n3951), .C2(EBX_REG_12__SCAN_IN), .A(n3990), .B(n3969), 
        .ZN(n3991) );
  NAND2_X1 U4906 ( .A1(n3992), .A2(n3991), .ZN(n4873) );
  NAND2_X1 U4907 ( .A1(n5665), .A2(n4873), .ZN(n4937) );
  NAND2_X1 U4908 ( .A1(n5181), .A2(EBX_REG_13__SCAN_IN), .ZN(n3994) );
  OR2_X1 U4909 ( .A1(n4035), .A2(EBX_REG_13__SCAN_IN), .ZN(n3993) );
  OAI211_X1 U4910 ( .C1(n4303), .C2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(n3994), .B(n3993), .ZN(n4938) );
  INV_X1 U4911 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U4912 ( .A1(n3961), .A2(n5227), .ZN(n3997) );
  INV_X1 U4913 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U4914 ( .A1(n4030), .A2(n5349), .ZN(n3995) );
  OAI211_X1 U4915 ( .C1(EBX_REG_14__SCAN_IN), .C2(n3951), .A(n3995), .B(n3969), 
        .ZN(n3996) );
  NAND2_X1 U4916 ( .A1(n3997), .A2(n3996), .ZN(n5222) );
  NAND2_X1 U4917 ( .A1(n5221), .A2(n5222), .ZN(n5223) );
  OR2_X1 U4918 ( .A1(n4035), .A2(EBX_REG_15__SCAN_IN), .ZN(n4000) );
  NAND2_X1 U4919 ( .A1(n3969), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3998) );
  OAI211_X1 U4920 ( .C1(n3951), .C2(EBX_REG_15__SCAN_IN), .A(n4030), .B(n3998), 
        .ZN(n3999) );
  NAND2_X1 U4921 ( .A1(n4000), .A2(n3999), .ZN(n5138) );
  INV_X1 U4922 ( .A(EBX_REG_16__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U4923 ( .A1(n3961), .A2(n6556), .ZN(n4003) );
  INV_X1 U4924 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U4925 ( .A1(n4030), .A2(n5582), .ZN(n4001) );
  OAI211_X1 U4926 ( .C1(n3951), .C2(EBX_REG_16__SCAN_IN), .A(n4001), .B(n3969), 
        .ZN(n4002) );
  NAND2_X1 U4927 ( .A1(n4003), .A2(n4002), .ZN(n5208) );
  OR2_X1 U4928 ( .A1(n4035), .A2(EBX_REG_17__SCAN_IN), .ZN(n4006) );
  NAND2_X1 U4929 ( .A1(n3969), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4004) );
  OAI211_X1 U4930 ( .C1(n3951), .C2(EBX_REG_17__SCAN_IN), .A(n4030), .B(n4004), 
        .ZN(n4005) );
  NAND2_X1 U4931 ( .A1(n4006), .A2(n4005), .ZN(n5125) );
  INV_X1 U4932 ( .A(EBX_REG_19__SCAN_IN), .ZN(n4007) );
  NAND2_X1 U4933 ( .A1(n3961), .A2(n4007), .ZN(n4011) );
  NAND2_X1 U4934 ( .A1(n4039), .A2(EBX_REG_19__SCAN_IN), .ZN(n4010) );
  NAND2_X1 U4935 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n4043), .ZN(n4008) );
  NAND4_X1 U4936 ( .A1(n4011), .A2(n4010), .A3(n4009), .A4(n4008), .ZN(n5192)
         );
  OR2_X1 U4937 ( .A1(n4303), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4012)
         );
  OR2_X1 U4938 ( .A1(n4043), .A2(EBX_REG_18__SCAN_IN), .ZN(n5191) );
  OAI22_X1 U4939 ( .A1(n4303), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n3951), .ZN(n5183) );
  NAND2_X1 U4940 ( .A1(n5189), .A2(n5183), .ZN(n4014) );
  NAND2_X1 U4941 ( .A1(n5181), .A2(EBX_REG_20__SCAN_IN), .ZN(n4013) );
  OAI211_X1 U4942 ( .C1(n5189), .C2(n5181), .A(n4014), .B(n4013), .ZN(n4015)
         );
  INV_X1 U4943 ( .A(n4015), .ZN(n4016) );
  NAND2_X1 U4944 ( .A1(n5180), .A2(n4016), .ZN(n5116) );
  OR2_X1 U4945 ( .A1(n4035), .A2(EBX_REG_21__SCAN_IN), .ZN(n4019) );
  NAND2_X1 U4946 ( .A1(n3969), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4017) );
  OAI211_X1 U4947 ( .C1(n3951), .C2(EBX_REG_21__SCAN_IN), .A(n4030), .B(n4017), 
        .ZN(n4018) );
  NAND2_X1 U4948 ( .A1(n4019), .A2(n4018), .ZN(n5115) );
  INV_X1 U4949 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U4950 ( .A1(n3961), .A2(n5503), .ZN(n4022) );
  INV_X1 U4951 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U4952 ( .A1(n4030), .A2(n5417), .ZN(n4020) );
  OAI211_X1 U4953 ( .C1(n3951), .C2(EBX_REG_22__SCAN_IN), .A(n4020), .B(n3969), 
        .ZN(n4021) );
  OR2_X1 U4954 ( .A1(n4035), .A2(EBX_REG_23__SCAN_IN), .ZN(n4025) );
  OR2_X1 U4955 ( .A1(n4303), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4024)
         );
  NAND2_X1 U4956 ( .A1(n5181), .A2(EBX_REG_23__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U4957 ( .A1(n4039), .A2(EBX_REG_24__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n3951), .ZN(n4028) );
  INV_X1 U4958 ( .A(EBX_REG_24__SCAN_IN), .ZN(n4026) );
  NAND2_X1 U4959 ( .A1(n3961), .A2(n4026), .ZN(n4027) );
  NAND2_X1 U4960 ( .A1(n4028), .A2(n4027), .ZN(n5156) );
  OR2_X1 U4961 ( .A1(n4035), .A2(EBX_REG_25__SCAN_IN), .ZN(n4032) );
  NAND2_X1 U4962 ( .A1(n3969), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4029) );
  OAI211_X1 U4963 ( .C1(n4043), .C2(EBX_REG_25__SCAN_IN), .A(n4030), .B(n4029), 
        .ZN(n4031) );
  NAND2_X1 U4964 ( .A1(n4032), .A2(n4031), .ZN(n5149) );
  AOI22_X1 U4965 ( .A1(n4039), .A2(EBX_REG_26__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n3951), .ZN(n4034) );
  INV_X1 U4966 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5145) );
  NAND2_X1 U4967 ( .A1(n3961), .A2(n5145), .ZN(n4033) );
  NAND2_X1 U4968 ( .A1(n4034), .A2(n4033), .ZN(n5103) );
  NAND2_X1 U4969 ( .A1(n5151), .A2(n5103), .ZN(n5105) );
  INV_X1 U4970 ( .A(EBX_REG_27__SCAN_IN), .ZN(n4038) );
  OR2_X1 U4971 ( .A1(n4035), .A2(EBX_REG_27__SCAN_IN), .ZN(n4037) );
  OR2_X1 U4972 ( .A1(n4303), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4036)
         );
  OAI211_X1 U4973 ( .C1(n4038), .C2(n3969), .A(n4037), .B(n4036), .ZN(n5090)
         );
  AOI22_X1 U4974 ( .A1(n4039), .A2(EBX_REG_28__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n3951), .ZN(n4041) );
  INV_X1 U4975 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5144) );
  NAND2_X1 U4976 ( .A1(n3961), .A2(n5144), .ZN(n4040) );
  AND2_X1 U4977 ( .A1(n4041), .A2(n4040), .ZN(n5076) );
  OAI22_X1 U4978 ( .A1(n4303), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n3951), .ZN(n5015) );
  NAND2_X1 U4979 ( .A1(n2980), .A2(n3969), .ZN(n4193) );
  INV_X1 U4980 ( .A(n5078), .ZN(n4042) );
  NAND2_X1 U4981 ( .A1(n2980), .A2(n4042), .ZN(n4045) );
  AND2_X1 U4982 ( .A1(n4043), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4044)
         );
  AOI21_X1 U4983 ( .B1(n4303), .B2(EBX_REG_30__SCAN_IN), .A(n4044), .ZN(n4192)
         );
  INV_X1 U4984 ( .A(n4192), .ZN(n4046) );
  NAND3_X1 U4985 ( .A1(n4193), .A2(n4045), .A3(n4046), .ZN(n4049) );
  AOI21_X1 U4986 ( .B1(n5078), .B2(n5181), .A(n4046), .ZN(n4047) );
  NAND2_X1 U4987 ( .A1(n4047), .A2(n2980), .ZN(n4048) );
  NAND2_X1 U4988 ( .A1(n4049), .A2(n4048), .ZN(n5070) );
  INV_X1 U4989 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4050) );
  NAND2_X1 U4990 ( .A1(n4468), .A2(n2970), .ZN(n4054) );
  NAND2_X1 U4991 ( .A1(n4057), .A2(n4064), .ZN(n4079) );
  XNOR2_X1 U4992 ( .A(n4079), .B(n4078), .ZN(n4052) );
  AND2_X1 U4993 ( .A1(n3192), .A2(n3188), .ZN(n4055) );
  AOI21_X1 U4994 ( .B1(n4052), .B2(n2954), .A(n4055), .ZN(n4053) );
  NAND2_X1 U4995 ( .A1(n4054), .A2(n4053), .ZN(n5832) );
  NAND2_X1 U4996 ( .A1(n5832), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4072)
         );
  INV_X1 U4997 ( .A(n2970), .ZN(n4060) );
  INV_X1 U4998 ( .A(n2954), .ZN(n4248) );
  INV_X1 U4999 ( .A(n4055), .ZN(n4056) );
  OAI21_X1 U5000 ( .B1(n4248), .B2(n4057), .A(n4056), .ZN(n4058) );
  INV_X1 U5001 ( .A(n4058), .ZN(n4059) );
  NAND2_X1 U5002 ( .A1(n4275), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4061)
         );
  INV_X1 U5003 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4980) );
  NAND2_X1 U5004 ( .A1(n4061), .A2(n4980), .ZN(n4063) );
  AND2_X1 U5005 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4062) );
  NAND2_X1 U5006 ( .A1(n4275), .A2(n4062), .ZN(n4070) );
  AND2_X1 U5007 ( .A1(n4063), .A2(n4070), .ZN(n4367) );
  NAND2_X1 U5008 ( .A1(n4471), .A2(n2970), .ZN(n4069) );
  XNOR2_X1 U5009 ( .A(n4065), .B(n4064), .ZN(n4067) );
  NAND3_X1 U5010 ( .A1(n4290), .A2(n3193), .A3(n3188), .ZN(n4066) );
  AOI21_X1 U5011 ( .B1(n4067), .B2(n2954), .A(n4066), .ZN(n4068) );
  NAND2_X1 U5012 ( .A1(n4069), .A2(n4068), .ZN(n4368) );
  INV_X1 U5013 ( .A(n4070), .ZN(n4071) );
  NAND2_X1 U5014 ( .A1(n4072), .A2(n5833), .ZN(n4076) );
  INV_X1 U5015 ( .A(n5832), .ZN(n4074) );
  INV_X1 U5016 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4073) );
  NAND2_X1 U5017 ( .A1(n4074), .A2(n4073), .ZN(n4075) );
  NAND2_X1 U5018 ( .A1(n4079), .A2(n4078), .ZN(n4087) );
  INV_X1 U5019 ( .A(n4086), .ZN(n4080) );
  XNOR2_X1 U5020 ( .A(n4087), .B(n4080), .ZN(n4081) );
  NAND2_X1 U5021 ( .A1(n4081), .A2(n2954), .ZN(n4082) );
  NAND2_X1 U5022 ( .A1(n4735), .A2(n4737), .ZN(n4736) );
  NAND2_X1 U5023 ( .A1(n4083), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4084)
         );
  NAND2_X1 U5024 ( .A1(n4736), .A2(n4084), .ZN(n5826) );
  NAND2_X1 U5025 ( .A1(n4085), .A2(n2970), .ZN(n4090) );
  NAND2_X1 U5026 ( .A1(n4087), .A2(n4086), .ZN(n4105) );
  XNOR2_X1 U5027 ( .A(n4105), .B(n4102), .ZN(n4088) );
  NAND2_X1 U5028 ( .A1(n4088), .A2(n2954), .ZN(n4089) );
  NAND2_X1 U5029 ( .A1(n4090), .A2(n4089), .ZN(n4091) );
  XNOR2_X1 U5030 ( .A(n4091), .B(n5894), .ZN(n5825) );
  NAND2_X1 U5031 ( .A1(n4091), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4092)
         );
  NAND2_X1 U5032 ( .A1(n5824), .A2(n4092), .ZN(n4744) );
  NAND2_X1 U5033 ( .A1(n4093), .A2(n2970), .ZN(n4098) );
  INV_X1 U5034 ( .A(n4102), .ZN(n4094) );
  OR2_X1 U5035 ( .A1(n4105), .A2(n4094), .ZN(n4095) );
  XNOR2_X1 U5036 ( .A(n4095), .B(n4103), .ZN(n4096) );
  NAND2_X1 U5037 ( .A1(n4096), .A2(n2954), .ZN(n4097) );
  NAND2_X1 U5038 ( .A1(n4098), .A2(n4097), .ZN(n4099) );
  INV_X1 U5039 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4806) );
  XNOR2_X1 U5040 ( .A(n4099), .B(n4806), .ZN(n4743) );
  NAND2_X1 U5041 ( .A1(n4744), .A2(n4743), .ZN(n4742) );
  NAND2_X1 U5042 ( .A1(n4099), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4100)
         );
  NAND2_X1 U5043 ( .A1(n4742), .A2(n4100), .ZN(n4622) );
  NAND3_X1 U5044 ( .A1(n4122), .A2(n2970), .A3(n4101), .ZN(n4108) );
  NAND2_X1 U5045 ( .A1(n4103), .A2(n4102), .ZN(n4104) );
  OR2_X1 U5046 ( .A1(n4105), .A2(n4104), .ZN(n4112) );
  XNOR2_X1 U5047 ( .A(n4112), .B(n4113), .ZN(n4106) );
  NAND2_X1 U5048 ( .A1(n4106), .A2(n2954), .ZN(n4107) );
  NAND2_X1 U5049 ( .A1(n4108), .A2(n4107), .ZN(n4109) );
  INV_X1 U5050 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4805) );
  XNOR2_X1 U5051 ( .A(n4109), .B(n4805), .ZN(n4621) );
  NAND2_X1 U5052 ( .A1(n4109), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4110)
         );
  NAND2_X1 U5053 ( .A1(n4624), .A2(n4110), .ZN(n4682) );
  NAND2_X1 U5054 ( .A1(n4111), .A2(n2970), .ZN(n4117) );
  INV_X1 U5055 ( .A(n4112), .ZN(n4114) );
  NAND2_X1 U5056 ( .A1(n4114), .A2(n4113), .ZN(n4125) );
  XNOR2_X1 U5057 ( .A(n4125), .B(n4123), .ZN(n4115) );
  NAND2_X1 U5058 ( .A1(n4115), .A2(n2954), .ZN(n4116) );
  NAND2_X1 U5059 ( .A1(n4117), .A2(n4116), .ZN(n4118) );
  INV_X1 U5060 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4955) );
  XNOR2_X1 U5061 ( .A(n4118), .B(n4955), .ZN(n4681) );
  NAND2_X1 U5062 ( .A1(n4118), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4119)
         );
  NAND2_X1 U5063 ( .A1(n4680), .A2(n4119), .ZN(n4794) );
  NAND2_X1 U5064 ( .A1(n4123), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4120) );
  INV_X1 U5065 ( .A(n4123), .ZN(n4124) );
  OR3_X1 U5066 ( .A1(n4125), .A2(n4124), .A3(n4248), .ZN(n4126) );
  NAND2_X1 U5067 ( .A1(n4130), .A2(n4126), .ZN(n4127) );
  INV_X1 U5068 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6492) );
  XNOR2_X1 U5069 ( .A(n4127), .B(n6492), .ZN(n4793) );
  NAND2_X1 U5070 ( .A1(n4127), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4128)
         );
  INV_X2 U5071 ( .A(n4130), .ZN(n5292) );
  NAND2_X1 U5072 ( .A1(n5298), .A2(n6461), .ZN(n4865) );
  OR2_X1 U5073 ( .A1(n5298), .A2(n6461), .ZN(n4866) );
  NAND2_X1 U5074 ( .A1(n5298), .A2(n4129), .ZN(n4924) );
  NAND2_X2 U5075 ( .A1(n4923), .A2(n4924), .ZN(n5807) );
  INV_X1 U5076 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4131) );
  AND2_X1 U5077 ( .A1(n5298), .A2(n4131), .ZN(n4133) );
  OR2_X1 U5078 ( .A1(n5298), .A2(n4129), .ZN(n5806) );
  NOR2_X1 U5079 ( .A1(n5808), .A2(n4968), .ZN(n4944) );
  XNOR2_X1 U5080 ( .A(n5808), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5561)
         );
  INV_X1 U5081 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4134) );
  AND2_X1 U5082 ( .A1(n5298), .A2(n5349), .ZN(n4136) );
  INV_X1 U5083 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5591) );
  NOR2_X1 U5084 ( .A1(n5808), .A2(n5591), .ZN(n4138) );
  NAND2_X1 U5085 ( .A1(n5298), .A2(n5591), .ZN(n4137) );
  NAND2_X1 U5086 ( .A1(n5298), .A2(n5582), .ZN(n5334) );
  NAND2_X1 U5087 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5000) );
  NAND2_X1 U5088 ( .A1(n5298), .A2(n5000), .ZN(n4139) );
  NAND2_X1 U5089 ( .A1(n5334), .A2(n4139), .ZN(n4140) );
  OR2_X2 U5090 ( .A1(n5333), .A2(n4140), .ZN(n5287) );
  OR2_X1 U5091 ( .A1(n5298), .A2(n5582), .ZN(n5335) );
  NOR2_X1 U5092 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4141) );
  OR2_X1 U5093 ( .A1(n5298), .A2(n4141), .ZN(n4142) );
  INV_X1 U5094 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5442) );
  NOR2_X1 U5095 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5411) );
  NOR2_X1 U5096 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5395) );
  INV_X1 U5097 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5289) );
  NAND3_X1 U5098 ( .A1(n5411), .A2(n5395), .A3(n5289), .ZN(n4145) );
  AND2_X1 U5099 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5410) );
  AND2_X1 U5100 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5435) );
  AND2_X1 U5101 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4995) );
  AND3_X1 U5102 ( .A1(n5410), .A2(n5435), .A3(n4995), .ZN(n5001) );
  XNOR2_X1 U5103 ( .A(n5808), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5278)
         );
  INV_X1 U5104 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U5105 ( .A1(n5298), .A2(n5385), .ZN(n4146) );
  NAND2_X1 U5106 ( .A1(n4224), .A2(n4146), .ZN(n4149) );
  INV_X1 U5107 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5367) );
  INV_X1 U5108 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4147) );
  NAND2_X1 U5109 ( .A1(n5367), .A2(n4147), .ZN(n5359) );
  OR3_X1 U5110 ( .A1(n5808), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n5359), 
        .ZN(n4225) );
  INV_X1 U5111 ( .A(n4225), .ZN(n4148) );
  NAND2_X1 U5112 ( .A1(n4149), .A2(n4148), .ZN(n4154) );
  INV_X1 U5113 ( .A(n4988), .ZN(n4153) );
  INV_X1 U5114 ( .A(n4149), .ZN(n4151) );
  INV_X1 U5115 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6476) );
  NAND2_X1 U5116 ( .A1(n4151), .A2(n4150), .ZN(n5262) );
  NAND2_X1 U5117 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5358) );
  NOR2_X2 U5118 ( .A1(n5262), .A2(n5358), .ZN(n4989) );
  INV_X1 U5119 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5035) );
  NAND2_X1 U5120 ( .A1(n4989), .A2(n5035), .ZN(n4152) );
  NAND2_X1 U5121 ( .A1(n4153), .A2(n4152), .ZN(n4157) );
  INV_X1 U5122 ( .A(n4154), .ZN(n4155) );
  NOR3_X1 U5123 ( .A1(n4989), .A2(n4155), .A3(n5035), .ZN(n4156) );
  AND2_X1 U5124 ( .A1(n4976), .A2(n3192), .ZN(n4158) );
  NOR2_X1 U5125 ( .A1(n3879), .A2(n4158), .ZN(n4277) );
  NAND3_X1 U5127 ( .A1(n3297), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6340) );
  INV_X1 U5128 ( .A(n6340), .ZN(n4163) );
  NOR2_X2 U5129 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6232) );
  AND2_X1 U5130 ( .A1(n4164), .A2(n6221), .ZN(n6439) );
  INV_X1 U5131 ( .A(n6439), .ZN(n4165) );
  NAND2_X1 U5132 ( .A1(n4165), .A2(n3297), .ZN(n4166) );
  NAND2_X1 U5133 ( .A1(n3297), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4168) );
  NAND2_X1 U5134 ( .A1(n6455), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4167) );
  AND2_X1 U5135 ( .A1(n4168), .A2(n4167), .ZN(n4363) );
  NAND2_X1 U5136 ( .A1(n3297), .A2(n6442), .ZN(n6339) );
  INV_X2 U5137 ( .A(n5885), .ZN(n5910) );
  NAND2_X1 U5138 ( .A1(n5910), .A2(REIP_REG_29__SCAN_IN), .ZN(n5033) );
  OAI21_X1 U5139 ( .B1(n5323), .B2(n4169), .A(n5033), .ZN(n4170) );
  AOI21_X1 U5140 ( .B1(n5558), .B2(n5023), .A(n4170), .ZN(n4171) );
  NAND3_X1 U5141 ( .A1(n4172), .A2(n3058), .A3(n4171), .ZN(U2957) );
  AOI22_X1 U5142 ( .A1(n4174), .A2(EAX_REG_31__SCAN_IN), .B1(n4173), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4175) );
  INV_X1 U5143 ( .A(n4177), .ZN(n4178) );
  NAND3_X1 U5144 ( .A1(n4182), .A2(n4181), .A3(n4180), .ZN(n4184) );
  AOI21_X1 U5145 ( .B1(n4185), .B2(n4184), .A(n4183), .ZN(n4282) );
  NOR2_X1 U5146 ( .A1(n4278), .A2(n4282), .ZN(n4233) );
  NAND2_X1 U5147 ( .A1(n4233), .A2(n6332), .ZN(n4231) );
  NOR2_X1 U5148 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6445) );
  NAND3_X1 U5149 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), 
        .A3(n6445), .ZN(n6328) );
  INV_X1 U5150 ( .A(n6339), .ZN(n4186) );
  NAND3_X1 U5151 ( .A1(n4186), .A2(STATE2_REG_1__SCAN_IN), .A3(n6455), .ZN(
        n6336) );
  INV_X1 U5152 ( .A(n4188), .ZN(n4189) );
  INV_X1 U5153 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5065) );
  INV_X1 U5154 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4214) );
  NOR2_X1 U5155 ( .A1(n4719), .A2(n6538), .ZN(n4191) );
  NAND2_X1 U5156 ( .A1(n5230), .A2(n5692), .ZN(n4221) );
  INV_X1 U5157 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5026) );
  NAND2_X1 U5158 ( .A1(n3961), .A2(n5026), .ZN(n5014) );
  NAND2_X1 U5159 ( .A1(n5018), .A2(n4192), .ZN(n4194) );
  NAND2_X1 U5160 ( .A1(n4194), .A2(n4193), .ZN(n4196) );
  OAI22_X1 U5161 ( .A1(n4303), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n3951), .ZN(n4195) );
  XNOR2_X1 U5162 ( .A(n4196), .B(n4195), .ZN(n5062) );
  NAND2_X1 U5163 ( .A1(n6345), .A2(n6455), .ZN(n4714) );
  NAND2_X1 U5164 ( .A1(n4714), .A2(EBX_REG_31__SCAN_IN), .ZN(n4197) );
  NAND2_X1 U5165 ( .A1(n4198), .A2(n6351), .ZN(n4281) );
  INV_X1 U5166 ( .A(n4281), .ZN(n6346) );
  NOR2_X1 U5167 ( .A1(n4517), .A2(n6346), .ZN(n4287) );
  INV_X1 U5168 ( .A(n4714), .ZN(n4199) );
  NAND2_X1 U5169 ( .A1(n4715), .A2(n4199), .ZN(n4200) );
  INV_X1 U5170 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6381) );
  INV_X1 U5171 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6373) );
  INV_X1 U5172 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6369) );
  INV_X1 U5173 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6367) );
  INV_X1 U5174 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6362) );
  NAND3_X1 U5175 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5710) );
  NOR2_X1 U5176 ( .A1(n6362), .A2(n5710), .ZN(n4761) );
  NAND2_X1 U5177 ( .A1(REIP_REG_5__SCAN_IN), .A2(n4761), .ZN(n4765) );
  NOR3_X1 U5178 ( .A1(n6369), .A2(n6367), .A3(n4765), .ZN(n4718) );
  NAND2_X1 U5179 ( .A1(REIP_REG_8__SCAN_IN), .A2(n4718), .ZN(n4781) );
  NAND2_X1 U5180 ( .A1(REIP_REG_9__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .ZN(
        n5663) );
  NOR3_X1 U5181 ( .A1(n6373), .A2(n4781), .A3(n5663), .ZN(n4879) );
  AND2_X1 U5182 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5139), .ZN(n5637) );
  NAND2_X1 U5183 ( .A1(REIP_REG_16__SCAN_IN), .A2(n5637), .ZN(n5123) );
  NOR2_X1 U5184 ( .A1(n6381), .A2(n5123), .ZN(n4201) );
  NAND2_X1 U5185 ( .A1(n5734), .A2(n4201), .ZN(n5627) );
  NAND3_X1 U5186 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n4202) );
  AND3_X1 U5187 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4205) );
  NAND2_X1 U5188 ( .A1(n5494), .A2(n4205), .ZN(n5480) );
  NAND3_X1 U5189 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4208) );
  NAND2_X1 U5190 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4211) );
  NOR2_X1 U5191 ( .A1(n5066), .A2(REIP_REG_29__SCAN_IN), .ZN(n5029) );
  AND2_X1 U5192 ( .A1(n5735), .A2(n4201), .ZN(n5524) );
  INV_X1 U5193 ( .A(n4202), .ZN(n4203) );
  NAND2_X1 U5194 ( .A1(n5524), .A2(n4203), .ZN(n4204) );
  NAND2_X1 U5195 ( .A1(n5737), .A2(n4204), .ZN(n5522) );
  INV_X1 U5196 ( .A(n4205), .ZN(n4206) );
  NAND2_X1 U5197 ( .A1(n5734), .A2(n4206), .ZN(n4207) );
  NAND2_X1 U5198 ( .A1(n5522), .A2(n4207), .ZN(n5499) );
  INV_X1 U5199 ( .A(n4208), .ZN(n4209) );
  NOR2_X1 U5200 ( .A1(n5525), .A2(n4209), .ZN(n4210) );
  NOR2_X1 U5201 ( .A1(n5499), .A2(n4210), .ZN(n5111) );
  NAND2_X1 U5202 ( .A1(n5734), .A2(n4211), .ZN(n4212) );
  NAND2_X1 U5203 ( .A1(n5111), .A2(n4212), .ZN(n5081) );
  NOR2_X1 U5204 ( .A1(n5029), .A2(n5081), .ZN(n5063) );
  OAI21_X1 U5205 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5711), .A(n5063), .ZN(n4217) );
  INV_X1 U5206 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6539) );
  INV_X1 U5207 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6401) );
  NOR4_X1 U5208 ( .A1(n5066), .A2(REIP_REG_31__SCAN_IN), .A3(n6539), .A4(n6401), .ZN(n4216) );
  OR3_X1 U5209 ( .A1(n4281), .A2(READY_N), .A3(STATEBS16_REG_SCAN_IN), .ZN(
        n6319) );
  NAND3_X1 U5210 ( .A1(n2954), .A2(EBX_REG_31__SCAN_IN), .A3(n6319), .ZN(n4213) );
  OAI22_X1 U5211 ( .A1(n5678), .A2(n4214), .B1(n4754), .B2(n4213), .ZN(n4215)
         );
  AOI211_X1 U5212 ( .C1(n4217), .C2(REIP_REG_31__SCAN_IN), .A(n4216), .B(n4215), .ZN(n4218) );
  NAND2_X1 U5213 ( .A1(n4221), .A2(n4220), .ZN(U2796) );
  INV_X2 U5214 ( .A(n6225), .ZN(n5563) );
  NAND2_X1 U5215 ( .A1(n5910), .A2(REIP_REG_31__SCAN_IN), .ZN(n5053) );
  NAND2_X1 U5216 ( .A1(n5823), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4222)
         );
  OAI211_X1 U5217 ( .C1(n5840), .C2(n4719), .A(n5053), .B(n4222), .ZN(n4223)
         );
  AOI21_X1 U5218 ( .B1(n5230), .B2(n5563), .A(n4223), .ZN(n4229) );
  AND2_X1 U5219 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5051) );
  NOR4_X1 U5220 ( .A1(n5277), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n4225), .ZN(n4226) );
  AOI21_X1 U5221 ( .B1(n4989), .B2(n5051), .A(n4226), .ZN(n4227) );
  NAND2_X1 U5222 ( .A1(n5050), .A2(n5835), .ZN(n4228) );
  NAND2_X1 U5223 ( .A1(n4229), .A2(n4228), .ZN(U2955) );
  AND2_X1 U5224 ( .A1(n6232), .A2(n6538), .ZN(n6450) );
  AOI211_X1 U5225 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4231), .A(n6450), .B(
        n4244), .ZN(n4232) );
  INV_X1 U5226 ( .A(n4232), .ZN(U2788) );
  INV_X1 U5227 ( .A(n4233), .ZN(n4235) );
  NOR2_X1 U5228 ( .A1(n4466), .A2(n4749), .ZN(n4234) );
  AOI21_X1 U5229 ( .B1(n4235), .B2(n4177), .A(n4234), .ZN(n5607) );
  NOR2_X1 U5230 ( .A1(n4749), .A2(n4236), .ZN(n6453) );
  NAND2_X1 U5231 ( .A1(n6453), .A2(n4281), .ZN(n4237) );
  NAND2_X1 U5232 ( .A1(n4237), .A2(n6345), .ZN(n6441) );
  NAND2_X1 U5233 ( .A1(n5607), .A2(n6441), .ZN(n6287) );
  AND2_X1 U5234 ( .A1(n6287), .A2(n6332), .ZN(n5614) );
  INV_X1 U5235 ( .A(MORE_REG_SCAN_IN), .ZN(n4243) );
  INV_X1 U5236 ( .A(n4466), .ZN(n4311) );
  OR2_X1 U5237 ( .A1(n4424), .A2(n4311), .ZN(n4241) );
  INV_X1 U5238 ( .A(n4238), .ZN(n6285) );
  NAND2_X1 U5239 ( .A1(n4277), .A2(n4749), .ZN(n4423) );
  NAND3_X1 U5240 ( .A1(n6285), .A2(n4177), .A3(n4423), .ZN(n4239) );
  AOI22_X1 U5241 ( .A1(n4239), .A2(n4311), .B1(n3181), .B2(n4282), .ZN(n4240)
         );
  NAND2_X1 U5242 ( .A1(n4241), .A2(n4240), .ZN(n6289) );
  NAND2_X1 U5243 ( .A1(n6289), .A2(n5614), .ZN(n4242) );
  OAI21_X1 U5244 ( .B1(n5614), .B2(n4243), .A(n4242), .ZN(U3471) );
  OAI21_X1 U5245 ( .B1(n2954), .B2(n6345), .A(n4244), .ZN(n4259) );
  NAND2_X1 U5246 ( .A1(n4358), .A2(UWORD_REG_4__SCAN_IN), .ZN(n4247) );
  NOR2_X1 U5247 ( .A1(n4246), .A2(n3951), .ZN(n4437) );
  NAND2_X1 U5248 ( .A1(n4342), .A2(DATAI_4_), .ZN(n4263) );
  OAI211_X1 U5249 ( .C1(n4323), .C2(n4386), .A(n4247), .B(n4263), .ZN(U2928)
         );
  INV_X1 U5250 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4351) );
  OR2_X1 U5251 ( .A1(n4246), .A2(n4248), .ZN(n6320) );
  INV_X1 U5252 ( .A(n6320), .ZN(n4250) );
  NOR2_X1 U5253 ( .A1(n4278), .A2(n4249), .ZN(n6297) );
  OR2_X1 U5254 ( .A1(n4250), .A2(n6297), .ZN(n4251) );
  NAND2_X1 U5255 ( .A1(n5777), .A2(n4715), .ZN(n4389) );
  NAND2_X1 U5256 ( .A1(n3297), .A2(n4479), .ZN(n6440) );
  AOI22_X1 U5257 ( .A1(n4387), .A2(UWORD_REG_9__SCAN_IN), .B1(n5803), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4252) );
  OAI21_X1 U5258 ( .B1(n4351), .B2(n4389), .A(n4252), .ZN(U2898) );
  INV_X1 U5259 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4354) );
  AOI22_X1 U5260 ( .A1(n4387), .A2(UWORD_REG_10__SCAN_IN), .B1(n5803), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4253) );
  OAI21_X1 U5261 ( .B1(n4354), .B2(n4389), .A(n4253), .ZN(U2897) );
  INV_X1 U5262 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4348) );
  AOI22_X1 U5263 ( .A1(n4387), .A2(UWORD_REG_8__SCAN_IN), .B1(n5803), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4254) );
  OAI21_X1 U5264 ( .B1(n4348), .B2(n4389), .A(n4254), .ZN(U2899) );
  INV_X1 U5265 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4361) );
  AOI22_X1 U5266 ( .A1(n4387), .A2(UWORD_REG_12__SCAN_IN), .B1(n5803), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4255) );
  OAI21_X1 U5267 ( .B1(n4361), .B2(n4389), .A(n4255), .ZN(U2895) );
  INV_X1 U5268 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6456) );
  AOI22_X1 U5269 ( .A1(n4387), .A2(UWORD_REG_13__SCAN_IN), .B1(n5803), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4256) );
  OAI21_X1 U5270 ( .B1(n6456), .B2(n4389), .A(n4256), .ZN(U2894) );
  INV_X1 U5271 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4357) );
  AOI22_X1 U5272 ( .A1(n4387), .A2(UWORD_REG_11__SCAN_IN), .B1(n5803), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4257) );
  OAI21_X1 U5273 ( .B1(n4357), .B2(n4389), .A(n4257), .ZN(U2896) );
  INV_X1 U5274 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4339) );
  AOI22_X1 U5275 ( .A1(n4387), .A2(UWORD_REG_14__SCAN_IN), .B1(n5803), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4258) );
  OAI21_X1 U5276 ( .B1(n4339), .B2(n4389), .A(n4258), .ZN(U2893) );
  INV_X1 U5277 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6508) );
  NAND2_X1 U5278 ( .A1(n4358), .A2(LWORD_REG_14__SCAN_IN), .ZN(n4260) );
  NAND2_X1 U5279 ( .A1(n4342), .A2(DATAI_14_), .ZN(n4337) );
  OAI211_X1 U5280 ( .C1(n4323), .C2(n6508), .A(n4260), .B(n4337), .ZN(U2953)
         );
  NAND2_X1 U5281 ( .A1(n4358), .A2(LWORD_REG_7__SCAN_IN), .ZN(n4261) );
  NAND2_X1 U5282 ( .A1(n4342), .A2(DATAI_7_), .ZN(n4340) );
  OAI211_X1 U5283 ( .C1(n4323), .C2(n3450), .A(n4261), .B(n4340), .ZN(U2946)
         );
  INV_X1 U5284 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6489) );
  NAND2_X1 U5285 ( .A1(n4358), .A2(LWORD_REG_8__SCAN_IN), .ZN(n4262) );
  NAND2_X1 U5286 ( .A1(n4342), .A2(DATAI_8_), .ZN(n4346) );
  OAI211_X1 U5287 ( .C1(n4323), .C2(n6489), .A(n4262), .B(n4346), .ZN(U2947)
         );
  INV_X1 U5288 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6496) );
  NAND2_X1 U5289 ( .A1(n4259), .A2(LWORD_REG_4__SCAN_IN), .ZN(n4264) );
  OAI211_X1 U5290 ( .C1(n4323), .C2(n6496), .A(n4264), .B(n4263), .ZN(U2943)
         );
  INV_X1 U5291 ( .A(EAX_REG_10__SCAN_IN), .ZN(n5787) );
  NAND2_X1 U5292 ( .A1(n4259), .A2(LWORD_REG_10__SCAN_IN), .ZN(n4265) );
  NAND2_X1 U5293 ( .A1(n4342), .A2(DATAI_10_), .ZN(n4352) );
  OAI211_X1 U5294 ( .C1(n4323), .C2(n5787), .A(n4265), .B(n4352), .ZN(U2949)
         );
  INV_X1 U5295 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4384) );
  NAND2_X1 U5296 ( .A1(n4259), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4266) );
  NAND2_X1 U5297 ( .A1(n4342), .A2(DATAI_0_), .ZN(n4329) );
  OAI211_X1 U5298 ( .C1(n4323), .C2(n4384), .A(n4266), .B(n4329), .ZN(U2924)
         );
  INV_X1 U5299 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5781) );
  NAND2_X1 U5300 ( .A1(n4259), .A2(LWORD_REG_13__SCAN_IN), .ZN(n4267) );
  NAND2_X1 U5301 ( .A1(n4342), .A2(DATAI_13_), .ZN(n4324) );
  OAI211_X1 U5302 ( .C1(n4323), .C2(n5781), .A(n4267), .B(n4324), .ZN(U2952)
         );
  INV_X1 U5303 ( .A(EAX_REG_5__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U5304 ( .A1(n4259), .A2(LWORD_REG_5__SCAN_IN), .ZN(n4268) );
  NAND2_X1 U5305 ( .A1(n4342), .A2(DATAI_5_), .ZN(n4326) );
  OAI211_X1 U5306 ( .C1(n4323), .C2(n5794), .A(n4268), .B(n4326), .ZN(U2944)
         );
  INV_X1 U5307 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U5308 ( .A1(n4259), .A2(LWORD_REG_12__SCAN_IN), .ZN(n4269) );
  NAND2_X1 U5309 ( .A1(n4342), .A2(DATAI_12_), .ZN(n4359) );
  OAI211_X1 U5310 ( .C1(n4323), .C2(n5783), .A(n4269), .B(n4359), .ZN(U2951)
         );
  INV_X1 U5311 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U5312 ( .A1(n4259), .A2(LWORD_REG_11__SCAN_IN), .ZN(n4270) );
  NAND2_X1 U5313 ( .A1(n4342), .A2(DATAI_11_), .ZN(n4355) );
  OAI211_X1 U5314 ( .C1(n4323), .C2(n5785), .A(n4270), .B(n4355), .ZN(U2950)
         );
  INV_X1 U5315 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6574) );
  AOI22_X1 U5316 ( .A1(n4259), .A2(LWORD_REG_15__SCAN_IN), .B1(n4342), .B2(
        DATAI_15_), .ZN(n4271) );
  OAI21_X1 U5317 ( .B1(n6574), .B2(n4323), .A(n4271), .ZN(U2954) );
  INV_X1 U5318 ( .A(DATAI_6_), .ZN(n4552) );
  NOR2_X1 U5319 ( .A1(n4317), .A2(n4552), .ZN(n4273) );
  AOI21_X1 U5320 ( .B1(LWORD_REG_6__SCAN_IN), .B2(n4259), .A(n4273), .ZN(n4272) );
  OAI21_X1 U5321 ( .B1(n4551), .B2(n4323), .A(n4272), .ZN(U2945) );
  INV_X1 U5322 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6523) );
  AOI21_X1 U5323 ( .B1(UWORD_REG_6__SCAN_IN), .B2(n4259), .A(n4273), .ZN(n4274) );
  OAI21_X1 U5324 ( .B1(n6523), .B2(n4323), .A(n4274), .ZN(U2930) );
  XOR2_X1 U5325 ( .A(n4275), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n4362) );
  INV_X1 U5326 ( .A(n4362), .ZN(n4310) );
  NAND2_X1 U5327 ( .A1(n4277), .A2(n4276), .ZN(n4279) );
  NAND2_X1 U5328 ( .A1(n4279), .A2(n4278), .ZN(n4443) );
  NAND2_X1 U5329 ( .A1(n4311), .A2(n4280), .ZN(n4285) );
  NAND2_X1 U5330 ( .A1(n4517), .A2(n4281), .ZN(n4283) );
  NOR2_X1 U5331 ( .A1(n4282), .A2(READY_N), .ZN(n4312) );
  NAND3_X1 U5332 ( .A1(n4283), .A2(n4312), .A3(n4527), .ZN(n4284) );
  NAND3_X1 U5333 ( .A1(n4443), .A2(n4285), .A3(n4284), .ZN(n4286) );
  NAND2_X1 U5334 ( .A1(n4286), .A2(n6332), .ZN(n4294) );
  OR3_X1 U5335 ( .A1(n4246), .A2(n4287), .A3(READY_N), .ZN(n4289) );
  NAND3_X1 U5336 ( .A1(n4289), .A2(n4715), .A3(n4288), .ZN(n4292) );
  NAND3_X1 U5337 ( .A1(n4292), .A2(n4291), .A3(n4290), .ZN(n4293) );
  NOR2_X1 U5338 ( .A1(n2952), .A2(n3194), .ZN(n4295) );
  NOR2_X1 U5339 ( .A1(n4437), .A2(n4295), .ZN(n4296) );
  NAND4_X1 U5340 ( .A1(n4420), .A2(n4296), .A3(n6285), .A4(n4423), .ZN(n4297)
         );
  INV_X1 U5341 ( .A(n4298), .ZN(n4299) );
  INV_X1 U5342 ( .A(n4625), .ZN(n4301) );
  INV_X1 U5343 ( .A(n4307), .ZN(n4300) );
  NOR2_X1 U5344 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5459), .ZN(n4370)
         );
  OAI21_X1 U5345 ( .B1(n2952), .B2(n3187), .A(n6320), .ZN(n4302) );
  NOR2_X1 U5346 ( .A1(n4303), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4304)
         );
  OR2_X1 U5347 ( .A1(n4305), .A2(n4304), .ZN(n4755) );
  NOR2_X1 U5348 ( .A1(n5887), .A2(n4755), .ZN(n4306) );
  AOI211_X1 U5349 ( .C1(n5910), .C2(REIP_REG_0__SCAN_IN), .A(n4370), .B(n4306), 
        .ZN(n4309) );
  NAND2_X1 U5350 ( .A1(n4307), .A2(n6297), .ZN(n5463) );
  INV_X1 U5351 ( .A(n5463), .ZN(n4960) );
  NOR2_X1 U5352 ( .A1(n5910), .A2(n4307), .ZN(n4369) );
  OAI21_X1 U5353 ( .B1(n4960), .B2(n4369), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4308) );
  OAI211_X1 U5354 ( .C1(n4310), .C2(n5846), .A(n4309), .B(n4308), .ZN(U3018)
         );
  INV_X1 U5355 ( .A(n4420), .ZN(n5604) );
  NAND2_X1 U5356 ( .A1(n5604), .A2(n4312), .ZN(n4313) );
  NOR2_X1 U5357 ( .A1(n4419), .A2(n4315), .ZN(n4316) );
  NAND2_X1 U5358 ( .A1(n3205), .A2(n4501), .ZN(n4321) );
  XNOR2_X1 U5359 ( .A(n4320), .B(n4319), .ZN(n4760) );
  INV_X1 U5360 ( .A(n4321), .ZN(n4322) );
  INV_X1 U5361 ( .A(DATAI_0_), .ZN(n6464) );
  INV_X1 U5362 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6554) );
  OAI222_X1 U5363 ( .A1(n5534), .A2(n4760), .B1(n5249), .B2(n6464), .C1(n5248), 
        .C2(n6554), .ZN(U2891) );
  NAND2_X1 U5364 ( .A1(n4358), .A2(UWORD_REG_13__SCAN_IN), .ZN(n4325) );
  OAI211_X1 U5365 ( .C1(n4323), .C2(n6456), .A(n4325), .B(n4324), .ZN(U2937)
         );
  INV_X1 U5366 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4375) );
  NAND2_X1 U5367 ( .A1(n4358), .A2(UWORD_REG_5__SCAN_IN), .ZN(n4327) );
  OAI211_X1 U5368 ( .C1(n4323), .C2(n4375), .A(n4327), .B(n4326), .ZN(U2929)
         );
  INV_X1 U5369 ( .A(EAX_REG_1__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U5370 ( .A1(n4358), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4328) );
  NAND2_X1 U5371 ( .A1(n4342), .A2(DATAI_1_), .ZN(n4332) );
  OAI211_X1 U5372 ( .C1(n4323), .C2(n5802), .A(n4328), .B(n4332), .ZN(U2940)
         );
  NAND2_X1 U5373 ( .A1(n4358), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4330) );
  OAI211_X1 U5374 ( .C1(n4323), .C2(n6554), .A(n4330), .B(n4329), .ZN(U2939)
         );
  INV_X1 U5375 ( .A(EAX_REG_3__SCAN_IN), .ZN(n5798) );
  NAND2_X1 U5376 ( .A1(n4358), .A2(LWORD_REG_3__SCAN_IN), .ZN(n4331) );
  NAND2_X1 U5377 ( .A1(n4342), .A2(DATAI_3_), .ZN(n4335) );
  OAI211_X1 U5378 ( .C1(n4323), .C2(n5798), .A(n4331), .B(n4335), .ZN(U2942)
         );
  INV_X1 U5379 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4380) );
  NAND2_X1 U5380 ( .A1(n4358), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4333) );
  OAI211_X1 U5381 ( .C1(n4323), .C2(n4380), .A(n4333), .B(n4332), .ZN(U2925)
         );
  NAND2_X1 U5382 ( .A1(n4358), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4334) );
  NAND2_X1 U5383 ( .A1(n4342), .A2(DATAI_2_), .ZN(n4344) );
  OAI211_X1 U5384 ( .C1(n4323), .C2(n3629), .A(n4334), .B(n4344), .ZN(U2926)
         );
  INV_X1 U5385 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4378) );
  NAND2_X1 U5386 ( .A1(n4259), .A2(UWORD_REG_3__SCAN_IN), .ZN(n4336) );
  OAI211_X1 U5387 ( .C1(n4323), .C2(n4378), .A(n4336), .B(n4335), .ZN(U2927)
         );
  NAND2_X1 U5388 ( .A1(n4358), .A2(UWORD_REG_14__SCAN_IN), .ZN(n4338) );
  OAI211_X1 U5389 ( .C1(n4323), .C2(n4339), .A(n4338), .B(n4337), .ZN(U2938)
         );
  INV_X1 U5390 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4382) );
  NAND2_X1 U5391 ( .A1(n4358), .A2(UWORD_REG_7__SCAN_IN), .ZN(n4341) );
  OAI211_X1 U5392 ( .C1(n4323), .C2(n4382), .A(n4341), .B(n4340), .ZN(U2931)
         );
  INV_X1 U5393 ( .A(EAX_REG_9__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U5394 ( .A1(n4358), .A2(LWORD_REG_9__SCAN_IN), .ZN(n4343) );
  NAND2_X1 U5395 ( .A1(n4342), .A2(DATAI_9_), .ZN(n4349) );
  OAI211_X1 U5396 ( .C1(n4323), .C2(n5789), .A(n4343), .B(n4349), .ZN(U2948)
         );
  INV_X1 U5397 ( .A(EAX_REG_2__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U5398 ( .A1(n4358), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4345) );
  OAI211_X1 U5399 ( .C1(n4323), .C2(n5800), .A(n4345), .B(n4344), .ZN(U2941)
         );
  NAND2_X1 U5400 ( .A1(n4358), .A2(UWORD_REG_8__SCAN_IN), .ZN(n4347) );
  OAI211_X1 U5401 ( .C1(n4323), .C2(n4348), .A(n4347), .B(n4346), .ZN(U2932)
         );
  NAND2_X1 U5402 ( .A1(n4358), .A2(UWORD_REG_9__SCAN_IN), .ZN(n4350) );
  OAI211_X1 U5403 ( .C1(n4323), .C2(n4351), .A(n4350), .B(n4349), .ZN(U2933)
         );
  NAND2_X1 U5404 ( .A1(n4358), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4353) );
  OAI211_X1 U5405 ( .C1(n4323), .C2(n4354), .A(n4353), .B(n4352), .ZN(U2934)
         );
  NAND2_X1 U5406 ( .A1(n4358), .A2(UWORD_REG_11__SCAN_IN), .ZN(n4356) );
  OAI211_X1 U5407 ( .C1(n4323), .C2(n4357), .A(n4356), .B(n4355), .ZN(U2935)
         );
  NAND2_X1 U5408 ( .A1(n4358), .A2(UWORD_REG_12__SCAN_IN), .ZN(n4360) );
  OAI211_X1 U5409 ( .C1(n4323), .C2(n4361), .A(n4360), .B(n4359), .ZN(U2936)
         );
  NAND2_X1 U5410 ( .A1(n4362), .A2(n5835), .ZN(n4366) );
  NAND2_X1 U5411 ( .A1(n5323), .A2(n4363), .ZN(n4364) );
  AOI22_X1 U5412 ( .A1(n4364), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .B1(n5910), 
        .B2(REIP_REG_0__SCAN_IN), .ZN(n4365) );
  OAI211_X1 U5413 ( .C1(n4760), .C2(n6225), .A(n4366), .B(n4365), .ZN(U2986)
         );
  XNOR2_X1 U5414 ( .A(n4368), .B(n4367), .ZN(n4676) );
  XNOR2_X1 U5415 ( .A(n5756), .B(n3951), .ZN(n4483) );
  INV_X1 U5416 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6429) );
  NOR2_X1 U5417 ( .A1(n5885), .A2(n6429), .ZN(n4672) );
  NOR2_X1 U5418 ( .A1(n4370), .A2(n4369), .ZN(n4807) );
  NOR2_X1 U5419 ( .A1(n4980), .A2(n4807), .ZN(n4371) );
  AOI211_X1 U5420 ( .C1(n5908), .C2(n4483), .A(n4672), .B(n4371), .ZN(n4373)
         );
  NAND2_X1 U5421 ( .A1(n4625), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4961)
         );
  INV_X1 U5422 ( .A(n5878), .ZN(n5916) );
  INV_X1 U5423 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5043) );
  NOR2_X1 U5424 ( .A1(n4996), .A2(n5043), .ZN(n5907) );
  OAI21_X1 U5425 ( .B1(n5916), .B2(n5907), .A(n4980), .ZN(n4372) );
  OAI211_X1 U5426 ( .C1(n4676), .C2(n5846), .A(n4373), .B(n4372), .ZN(U3017)
         );
  OAI222_X1 U5427 ( .A1(n4755), .A2(n5225), .B1(n5763), .B2(n4752), .C1(n5759), 
        .C2(n4760), .ZN(U2859) );
  AOI22_X1 U5428 ( .A1(n4387), .A2(UWORD_REG_5__SCAN_IN), .B1(n5795), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4374) );
  OAI21_X1 U5429 ( .B1(n4375), .B2(n4389), .A(n4374), .ZN(U2902) );
  AOI22_X1 U5430 ( .A1(n4387), .A2(UWORD_REG_2__SCAN_IN), .B1(n5795), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4376) );
  OAI21_X1 U5431 ( .B1(n3629), .B2(n4389), .A(n4376), .ZN(U2905) );
  AOI22_X1 U5432 ( .A1(n4387), .A2(UWORD_REG_3__SCAN_IN), .B1(n5795), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4377) );
  OAI21_X1 U5433 ( .B1(n4378), .B2(n4389), .A(n4377), .ZN(U2904) );
  AOI22_X1 U5434 ( .A1(n4387), .A2(UWORD_REG_1__SCAN_IN), .B1(n5795), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4379) );
  OAI21_X1 U5435 ( .B1(n4380), .B2(n4389), .A(n4379), .ZN(U2906) );
  AOI22_X1 U5436 ( .A1(n4387), .A2(UWORD_REG_7__SCAN_IN), .B1(n5795), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4381) );
  OAI21_X1 U5437 ( .B1(n4382), .B2(n4389), .A(n4381), .ZN(U2900) );
  AOI22_X1 U5438 ( .A1(n4387), .A2(UWORD_REG_0__SCAN_IN), .B1(n5795), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4383) );
  OAI21_X1 U5439 ( .B1(n4384), .B2(n4389), .A(n4383), .ZN(U2907) );
  AOI22_X1 U5440 ( .A1(n4387), .A2(UWORD_REG_4__SCAN_IN), .B1(n5795), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4385) );
  OAI21_X1 U5441 ( .B1(n4386), .B2(n4389), .A(n4385), .ZN(U2903) );
  AOI22_X1 U5442 ( .A1(n4387), .A2(UWORD_REG_6__SCAN_IN), .B1(n5795), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4388) );
  OAI21_X1 U5443 ( .B1(n6523), .B2(n4389), .A(n4388), .ZN(U2901) );
  INV_X1 U5444 ( .A(n4390), .ZN(n4393) );
  INV_X1 U5445 ( .A(n4391), .ZN(n4392) );
  NAND2_X1 U5446 ( .A1(n4393), .A2(n4392), .ZN(n4394) );
  AND2_X1 U5447 ( .A1(n4394), .A2(n4398), .ZN(n5752) );
  INV_X1 U5448 ( .A(n5752), .ZN(n4484) );
  INV_X1 U5449 ( .A(DATAI_1_), .ZN(n4518) );
  OAI222_X1 U5450 ( .A1(n4484), .A2(n5534), .B1(n5249), .B2(n4518), .C1(n5248), 
        .C2(n5802), .ZN(U2890) );
  OAI21_X1 U5451 ( .B1(n2969), .B2(n4396), .A(n4395), .ZN(n5723) );
  INV_X1 U5452 ( .A(DATAI_3_), .ZN(n6459) );
  OAI222_X1 U5453 ( .A1(n5723), .A2(n5534), .B1(n5249), .B2(n6459), .C1(n5248), 
        .C2(n5798), .ZN(U2888) );
  INV_X1 U5454 ( .A(n4397), .ZN(n4399) );
  AOI21_X1 U5455 ( .B1(n4399), .B2(n4398), .A(n2969), .ZN(n5836) );
  INV_X1 U5456 ( .A(n5836), .ZN(n4412) );
  INV_X1 U5457 ( .A(DATAI_2_), .ZN(n4400) );
  OAI222_X1 U5458 ( .A1(n4412), .A2(n5534), .B1(n5249), .B2(n4400), .C1(n5248), 
        .C2(n5800), .ZN(U2889) );
  AOI21_X1 U5459 ( .B1(n4401), .B2(n4410), .A(n4489), .ZN(n5897) );
  INV_X1 U5460 ( .A(n5897), .ZN(n5719) );
  OAI222_X1 U5461 ( .A1(n5719), .A2(n5225), .B1(n4402), .B2(n5763), .C1(n5723), 
        .C2(n5759), .ZN(U2856) );
  OR2_X1 U5462 ( .A1(n2956), .A2(n4404), .ZN(n4406) );
  NAND2_X1 U5463 ( .A1(n4403), .A2(n4406), .ZN(n5699) );
  INV_X1 U5464 ( .A(DATAI_5_), .ZN(n4407) );
  OAI222_X1 U5465 ( .A1(n5699), .A2(n5534), .B1(n5249), .B2(n4407), .C1(n5248), 
        .C2(n5794), .ZN(U2886) );
  OR2_X1 U5466 ( .A1(n4409), .A2(n4408), .ZN(n4411) );
  NAND2_X1 U5467 ( .A1(n4411), .A2(n4410), .ZN(n5905) );
  OAI222_X1 U5468 ( .A1(n5905), .A2(n5225), .B1(n5763), .B2(n3962), .C1(n4412), 
        .C2(n5759), .ZN(U2857) );
  AOI21_X1 U5469 ( .B1(n4413), .B2(n4491), .A(n2992), .ZN(n5875) );
  INV_X1 U5470 ( .A(n5875), .ZN(n4415) );
  INV_X1 U5471 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4414) );
  OAI222_X1 U5472 ( .A1(n4415), .A2(n5225), .B1(n4414), .B2(n5763), .C1(n5699), 
        .C2(n5759), .ZN(U2854) );
  INV_X1 U5473 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5613) );
  NAND2_X1 U5474 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5613), .ZN(n4463) );
  INV_X1 U5475 ( .A(n4416), .ZN(n4456) );
  INV_X1 U5476 ( .A(n4418), .ZN(n4422) );
  AND3_X1 U5477 ( .A1(n4420), .A2(n4419), .A3(n4246), .ZN(n4421) );
  NAND2_X1 U5478 ( .A1(n4422), .A2(n4421), .ZN(n6295) );
  NAND2_X1 U5479 ( .A1(n2971), .A2(n6295), .ZN(n4435) );
  NAND2_X1 U5480 ( .A1(n4424), .A2(n4423), .ZN(n4453) );
  MUX2_X1 U5481 ( .A(n4426), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4425), 
        .Z(n4427) );
  NOR2_X1 U5482 ( .A1(n4427), .A2(n4416), .ZN(n4433) );
  AOI21_X1 U5483 ( .B1(n4425), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3061), 
        .ZN(n4428) );
  NOR2_X1 U5484 ( .A1(n3750), .A2(n4428), .ZN(n6416) );
  NAND2_X1 U5485 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4429) );
  XNOR2_X1 U5486 ( .A(n4429), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4430)
         );
  NAND2_X1 U5487 ( .A1(n6297), .A2(n4430), .ZN(n4431) );
  OAI21_X1 U5488 ( .B1(n6416), .B2(n4450), .A(n4431), .ZN(n4432) );
  AOI21_X1 U5489 ( .B1(n4453), .B2(n4433), .A(n4432), .ZN(n4434) );
  NAND2_X1 U5490 ( .A1(n4435), .A2(n4434), .ZN(n6414) );
  INV_X1 U5491 ( .A(n4436), .ZN(n4444) );
  OAI21_X1 U5492 ( .B1(n6297), .B2(n3151), .A(n6346), .ZN(n4439) );
  INV_X1 U5493 ( .A(n4437), .ZN(n4438) );
  NAND2_X1 U5494 ( .A1(n4439), .A2(n4438), .ZN(n4440) );
  NAND3_X1 U5495 ( .A1(n4440), .A2(n4466), .A3(n6345), .ZN(n4441) );
  NAND2_X1 U5496 ( .A1(n4446), .A2(n4445), .ZN(n6298) );
  MUX2_X1 U5497 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6414), .S(n6298), 
        .Z(n6314) );
  INV_X1 U5498 ( .A(n6295), .ZN(n4979) );
  XNOR2_X1 U5499 ( .A(n4425), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4452)
         );
  XNOR2_X1 U5500 ( .A(n3062), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4448)
         );
  NAND2_X1 U5501 ( .A1(n6297), .A2(n4448), .ZN(n4449) );
  OAI21_X1 U5502 ( .B1(n4452), .B2(n4450), .A(n4449), .ZN(n4451) );
  AOI21_X1 U5503 ( .B1(n4453), .B2(n4452), .A(n4451), .ZN(n4454) );
  OAI21_X1 U5504 ( .B1(n4447), .B2(n4979), .A(n4454), .ZN(n5047) );
  MUX2_X1 U5505 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n5047), .S(n6298), 
        .Z(n6308) );
  NAND3_X1 U5506 ( .A1(n6314), .A2(n6308), .A3(n6538), .ZN(n4455) );
  OAI21_X1 U5507 ( .B1(n4463), .B2(n4456), .A(n4455), .ZN(n6293) );
  INV_X1 U5508 ( .A(n4457), .ZN(n4458) );
  NAND2_X1 U5509 ( .A1(n6293), .A2(n4458), .ZN(n4480) );
  INV_X1 U5510 ( .A(n6103), .ZN(n5995) );
  XNOR2_X1 U5511 ( .A(n4459), .B(n4460), .ZN(n5709) );
  NAND2_X1 U5512 ( .A1(n5709), .A2(n5604), .ZN(n4462) );
  OR2_X1 U5513 ( .A1(n6298), .A2(n4460), .ZN(n4461) );
  NAND2_X1 U5514 ( .A1(n4462), .A2(n4461), .ZN(n4465) );
  NOR2_X1 U5515 ( .A1(n4463), .A2(n4460), .ZN(n4464) );
  AOI21_X1 U5516 ( .B1(n4465), .B2(n6538), .A(n4464), .ZN(n6291) );
  AND3_X1 U5517 ( .A1(n4480), .A2(n6291), .A3(n5613), .ZN(n4467) );
  NAND2_X1 U5518 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4479), .ZN(n6410) );
  NAND2_X1 U5519 ( .A1(n4469), .A2(n4470), .ZN(n6224) );
  NOR2_X1 U5520 ( .A1(n6144), .A2(n6455), .ZN(n6137) );
  NAND2_X1 U5521 ( .A1(n4469), .A2(n4473), .ZN(n5991) );
  INV_X1 U5522 ( .A(n5991), .ZN(n4474) );
  NAND2_X1 U5523 ( .A1(n4474), .A2(n6067), .ZN(n6029) );
  NAND2_X1 U5524 ( .A1(n6029), .A2(n6065), .ZN(n4475) );
  OAI21_X1 U5525 ( .B1(n6137), .B2(n4475), .A(n6232), .ZN(n5953) );
  INV_X1 U5526 ( .A(n5953), .ZN(n4477) );
  INV_X1 U5527 ( .A(n4077), .ZN(n4554) );
  NOR2_X1 U5528 ( .A1(n6221), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6228) );
  INV_X1 U5529 ( .A(n6228), .ZN(n4891) );
  AND2_X1 U5530 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6413), .ZN(n5473) );
  OAI22_X1 U5531 ( .A1(n4554), .A2(n4891), .B1(n6189), .B2(n5473), .ZN(n4476)
         );
  OAI21_X1 U5532 ( .B1(n4477), .B2(n4476), .A(n5921), .ZN(n4478) );
  OAI21_X1 U5533 ( .B1(n5921), .B2(n6313), .A(n4478), .ZN(U3462) );
  AND3_X1 U5534 ( .A1(n4480), .A2(n6291), .A3(n4479), .ZN(n6325) );
  OAI22_X1 U5535 ( .A1(n6143), .A2(n6221), .B1(n3342), .B2(n5473), .ZN(n4481)
         );
  OAI21_X1 U5536 ( .B1(n6325), .B2(n4481), .A(n5921), .ZN(n4482) );
  OAI21_X1 U5537 ( .B1(n5921), .B2(n6138), .A(n4482), .ZN(U3465) );
  INV_X1 U5538 ( .A(n4483), .ZN(n4485) );
  OAI222_X1 U5539 ( .A1(n4485), .A2(n5758), .B1(n5763), .B2(n3952), .C1(n4484), 
        .C2(n5759), .ZN(U2858) );
  XOR2_X1 U5540 ( .A(n4395), .B(n4486), .Z(n5828) );
  INV_X1 U5541 ( .A(n5828), .ZN(n4488) );
  INV_X1 U5542 ( .A(DATAI_4_), .ZN(n4487) );
  OAI222_X1 U5543 ( .A1(n5534), .A2(n4488), .B1(n5249), .B2(n4487), .C1(n5248), 
        .C2(n6496), .ZN(U2887) );
  OR2_X1 U5544 ( .A1(n4490), .A2(n4489), .ZN(n4492) );
  NAND2_X1 U5545 ( .A1(n4492), .A2(n4491), .ZN(n5886) );
  OAI22_X1 U5546 ( .A1(n5758), .A2(n5886), .B1(n5763), .B2(n5706), .ZN(n4493)
         );
  AOI21_X1 U5547 ( .B1(n5828), .B2(n5211), .A(n4493), .ZN(n4494) );
  INV_X1 U5548 ( .A(n4494), .ZN(U2855) );
  OAI21_X1 U5549 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6413), .A(n4634), 
        .ZN(n4689) );
  NOR2_X1 U5550 ( .A1(n4470), .A2(n4472), .ZN(n4495) );
  AOI21_X1 U5551 ( .B1(n4502), .B2(STATEBS16_REG_SCAN_IN), .A(n6221), .ZN(
        n4503) );
  INV_X1 U5552 ( .A(n4496), .ZN(n5992) );
  NOR2_X1 U5553 ( .A1(n4447), .A2(n5992), .ZN(n6139) );
  NAND2_X1 U5554 ( .A1(n6139), .A2(n5995), .ZN(n4584) );
  OR2_X1 U5555 ( .A1(n4584), .A2(n3342), .ZN(n4498) );
  NOR2_X1 U5556 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6305), .ZN(n6142)
         );
  NAND2_X1 U5557 ( .A1(n6142), .A2(n6313), .ZN(n4581) );
  NOR2_X1 U5558 ( .A1(n6138), .A2(n4581), .ZN(n4541) );
  INV_X1 U5559 ( .A(n4541), .ZN(n4497) );
  AND2_X1 U5560 ( .A1(n4498), .A2(n4497), .ZN(n4504) );
  AOI22_X1 U5561 ( .A1(n4503), .A2(n4504), .B1(n4581), .B2(n6221), .ZN(n4499)
         );
  NAND2_X1 U5562 ( .A1(n6231), .A2(n4499), .ZN(n4546) );
  NAND2_X1 U5563 ( .A1(n5563), .A2(DATAI_23_), .ZN(n6284) );
  NOR2_X1 U5564 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6413), .ZN(n6409) );
  NAND2_X1 U5565 ( .A1(n4540), .A2(n4501), .ZN(n4837) );
  AND2_X1 U5566 ( .A1(n5563), .A2(DATAI_31_), .ZN(n6279) );
  AOI22_X1 U5567 ( .A1(n6277), .A2(n4541), .B1(n6279), .B2(n5986), .ZN(n4510)
         );
  INV_X1 U5568 ( .A(n4503), .ZN(n4505) );
  OR2_X1 U5569 ( .A1(n4505), .A2(n4504), .ZN(n4508) );
  INV_X1 U5570 ( .A(n4581), .ZN(n4506) );
  NAND2_X1 U5571 ( .A1(n4506), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4507) );
  NAND2_X1 U5572 ( .A1(n4508), .A2(n4507), .ZN(n4542) );
  INV_X1 U5573 ( .A(DATAI_7_), .ZN(n4616) );
  NOR2_X2 U5574 ( .A1(n4616), .A2(n4894), .ZN(n6275) );
  NAND2_X1 U5575 ( .A1(n4542), .A2(n6275), .ZN(n4509) );
  OAI211_X1 U5576 ( .C1(n6002), .C2(n6284), .A(n4510), .B(n4509), .ZN(n4511)
         );
  AOI21_X1 U5577 ( .B1(n4546), .B2(INSTQUEUE_REG_5__7__SCAN_IN), .A(n4511), 
        .ZN(n4512) );
  INV_X1 U5578 ( .A(n4512), .ZN(U3067) );
  NAND2_X1 U5579 ( .A1(n5563), .A2(DATAI_16_), .ZN(n6237) );
  NAND2_X1 U5580 ( .A1(n4540), .A2(n4715), .ZN(n4909) );
  AND2_X1 U5581 ( .A1(n5563), .A2(DATAI_24_), .ZN(n6234) );
  AOI22_X1 U5582 ( .A1(n6223), .A2(n4541), .B1(n6234), .B2(n5986), .ZN(n4514)
         );
  NAND2_X1 U5583 ( .A1(n4542), .A2(n6222), .ZN(n4513) );
  OAI211_X1 U5584 ( .C1(n6002), .C2(n6237), .A(n4514), .B(n4513), .ZN(n4515)
         );
  AOI21_X1 U5585 ( .B1(n4546), .B2(INSTQUEUE_REG_5__0__SCAN_IN), .A(n4515), 
        .ZN(n4516) );
  INV_X1 U5586 ( .A(n4516), .ZN(U3060) );
  NAND2_X1 U5587 ( .A1(n5563), .A2(DATAI_17_), .ZN(n6243) );
  NAND2_X1 U5588 ( .A1(n4540), .A2(n4517), .ZN(n4905) );
  AND2_X1 U5589 ( .A1(n5563), .A2(DATAI_25_), .ZN(n6240) );
  AOI22_X1 U5590 ( .A1(n6239), .A2(n4541), .B1(n6240), .B2(n5986), .ZN(n4520)
         );
  NAND2_X1 U5591 ( .A1(n4542), .A2(n6238), .ZN(n4519) );
  OAI211_X1 U5592 ( .C1(n6002), .C2(n6243), .A(n4520), .B(n4519), .ZN(n4521)
         );
  AOI21_X1 U5593 ( .B1(n4546), .B2(INSTQUEUE_REG_5__1__SCAN_IN), .A(n4521), 
        .ZN(n4522) );
  INV_X1 U5594 ( .A(n4522), .ZN(U3061) );
  NAND2_X1 U5595 ( .A1(n5563), .A2(DATAI_19_), .ZN(n6255) );
  NAND2_X1 U5596 ( .A1(n4540), .A2(n3188), .ZN(n4901) );
  AND2_X1 U5597 ( .A1(n5563), .A2(DATAI_27_), .ZN(n6252) );
  AOI22_X1 U5598 ( .A1(n6251), .A2(n4541), .B1(n6252), .B2(n5986), .ZN(n4524)
         );
  NAND2_X1 U5599 ( .A1(n4542), .A2(n6250), .ZN(n4523) );
  OAI211_X1 U5600 ( .C1(n6002), .C2(n6255), .A(n4524), .B(n4523), .ZN(n4525)
         );
  AOI21_X1 U5601 ( .B1(n4546), .B2(INSTQUEUE_REG_5__3__SCAN_IN), .A(n4525), 
        .ZN(n4526) );
  INV_X1 U5602 ( .A(n4526), .ZN(U3063) );
  NAND2_X1 U5603 ( .A1(n5563), .A2(DATAI_18_), .ZN(n6249) );
  NAND2_X1 U5604 ( .A1(n4540), .A2(n4527), .ZN(n4914) );
  AND2_X1 U5605 ( .A1(n5563), .A2(DATAI_26_), .ZN(n6246) );
  AOI22_X1 U5606 ( .A1(n6244), .A2(n4541), .B1(n6246), .B2(n5986), .ZN(n4529)
         );
  NAND2_X1 U5607 ( .A1(DATAI_2_), .A2(n4634), .ZN(n6160) );
  NAND2_X1 U5608 ( .A1(n6245), .A2(n4542), .ZN(n4528) );
  OAI211_X1 U5609 ( .C1(n6002), .C2(n6249), .A(n4529), .B(n4528), .ZN(n4530)
         );
  AOI21_X1 U5610 ( .B1(n4546), .B2(INSTQUEUE_REG_5__2__SCAN_IN), .A(n4530), 
        .ZN(n4531) );
  INV_X1 U5611 ( .A(n4531), .ZN(U3062) );
  NAND2_X1 U5612 ( .A1(n5563), .A2(DATAI_20_), .ZN(n6261) );
  NAND2_X1 U5613 ( .A1(n4540), .A2(n3187), .ZN(n4897) );
  AND2_X1 U5614 ( .A1(n5563), .A2(DATAI_28_), .ZN(n6258) );
  AOI22_X1 U5615 ( .A1(n6256), .A2(n4541), .B1(n6258), .B2(n5986), .ZN(n4533)
         );
  NAND2_X1 U5616 ( .A1(DATAI_4_), .A2(n4634), .ZN(n6168) );
  NAND2_X1 U5617 ( .A1(n6257), .A2(n4542), .ZN(n4532) );
  OAI211_X1 U5618 ( .C1(n6002), .C2(n6261), .A(n4533), .B(n4532), .ZN(n4534)
         );
  AOI21_X1 U5619 ( .B1(n4546), .B2(INSTQUEUE_REG_5__4__SCAN_IN), .A(n4534), 
        .ZN(n4535) );
  INV_X1 U5620 ( .A(n4535), .ZN(U3064) );
  NAND2_X1 U5621 ( .A1(n5563), .A2(DATAI_21_), .ZN(n6267) );
  NAND2_X1 U5622 ( .A1(n4540), .A2(n3193), .ZN(n4919) );
  AND2_X1 U5623 ( .A1(n5563), .A2(DATAI_29_), .ZN(n6264) );
  AOI22_X1 U5624 ( .A1(n6262), .A2(n4541), .B1(n6264), .B2(n5986), .ZN(n4537)
         );
  NAND2_X1 U5625 ( .A1(DATAI_5_), .A2(n4634), .ZN(n6172) );
  NAND2_X1 U5626 ( .A1(n6263), .A2(n4542), .ZN(n4536) );
  OAI211_X1 U5627 ( .C1(n6002), .C2(n6267), .A(n4537), .B(n4536), .ZN(n4538)
         );
  AOI21_X1 U5628 ( .B1(n4546), .B2(INSTQUEUE_REG_5__5__SCAN_IN), .A(n4538), 
        .ZN(n4539) );
  INV_X1 U5629 ( .A(n4539), .ZN(U3065) );
  NAND2_X1 U5630 ( .A1(n5563), .A2(DATAI_22_), .ZN(n6273) );
  NAND2_X1 U5631 ( .A1(n4540), .A2(n3178), .ZN(n4842) );
  AND2_X1 U5632 ( .A1(n5563), .A2(DATAI_30_), .ZN(n6270) );
  AOI22_X1 U5633 ( .A1(n6268), .A2(n4541), .B1(n6270), .B2(n5986), .ZN(n4544)
         );
  NAND2_X1 U5634 ( .A1(DATAI_6_), .A2(n4634), .ZN(n6176) );
  NAND2_X1 U5635 ( .A1(n6269), .A2(n4542), .ZN(n4543) );
  OAI211_X1 U5636 ( .C1(n6002), .C2(n6273), .A(n4544), .B(n4543), .ZN(n4545)
         );
  AOI21_X1 U5637 ( .B1(n4546), .B2(INSTQUEUE_REG_5__6__SCAN_IN), .A(n4545), 
        .ZN(n4547) );
  INV_X1 U5638 ( .A(n4547), .ZN(U3066) );
  OAI21_X1 U5639 ( .B1(n4548), .B2(n2992), .A(n4617), .ZN(n5690) );
  XNOR2_X1 U5640 ( .A(n4403), .B(n4549), .ZN(n5816) );
  OAI222_X1 U5641 ( .A1(n5758), .A2(n5690), .B1(n4550), .B2(n5763), .C1(n5759), 
        .C2(n5816), .ZN(U2853) );
  OAI222_X1 U5642 ( .A1(n4552), .A2(n5249), .B1(n5534), .B2(n5816), .C1(n4551), 
        .C2(n5248), .ZN(U2885) );
  NAND3_X1 U5643 ( .A1(n4554), .A2(n4553), .A3(n4687), .ZN(n4561) );
  AND2_X1 U5644 ( .A1(n4447), .A2(n4496), .ZN(n4886) );
  NAND2_X1 U5645 ( .A1(n6189), .A2(n4886), .ZN(n5927) );
  INV_X1 U5646 ( .A(n5927), .ZN(n4555) );
  INV_X1 U5647 ( .A(n3342), .ZN(n6296) );
  NAND3_X1 U5648 ( .A1(n6313), .A2(n6305), .A3(n6301), .ZN(n5922) );
  NOR2_X1 U5649 ( .A1(n6138), .A2(n5922), .ZN(n4578) );
  AOI21_X1 U5650 ( .B1(n4555), .B2(n6296), .A(n4578), .ZN(n4559) );
  OR2_X1 U5651 ( .A1(n4561), .A2(n6455), .ZN(n4556) );
  AOI22_X1 U5652 ( .A1(n4559), .A2(n4558), .B1(n6221), .B2(n5922), .ZN(n4557)
         );
  NAND2_X1 U5653 ( .A1(n6231), .A2(n4557), .ZN(n4577) );
  INV_X1 U5654 ( .A(n4558), .ZN(n4560) );
  OAI22_X1 U5655 ( .A1(n4560), .A2(n4559), .B1(n6442), .B2(n5922), .ZN(n4576)
         );
  AOI22_X1 U5656 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4577), .B1(n6263), 
        .B2(n4576), .ZN(n4563) );
  NOR2_X2 U5657 ( .A1(n4561), .A2(n6101), .ZN(n5947) );
  AOI22_X1 U5658 ( .A1(n5947), .A2(n6264), .B1(n6262), .B2(n4578), .ZN(n4562)
         );
  OAI211_X1 U5659 ( .C1(n6267), .C2(n4850), .A(n4563), .B(n4562), .ZN(U3033)
         );
  AOI22_X1 U5660 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4577), .B1(n6257), 
        .B2(n4576), .ZN(n4565) );
  AOI22_X1 U5661 ( .A1(n5947), .A2(n6258), .B1(n6256), .B2(n4578), .ZN(n4564)
         );
  OAI211_X1 U5662 ( .C1(n6261), .C2(n4850), .A(n4565), .B(n4564), .ZN(U3032)
         );
  AOI22_X1 U5663 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4577), .B1(n6245), 
        .B2(n4576), .ZN(n4567) );
  AOI22_X1 U5664 ( .A1(n5947), .A2(n6246), .B1(n6244), .B2(n4578), .ZN(n4566)
         );
  OAI211_X1 U5665 ( .C1(n6249), .C2(n4850), .A(n4567), .B(n4566), .ZN(U3030)
         );
  AOI22_X1 U5666 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4577), .B1(n6269), 
        .B2(n4576), .ZN(n4569) );
  AOI22_X1 U5667 ( .A1(n5947), .A2(n6270), .B1(n6268), .B2(n4578), .ZN(n4568)
         );
  OAI211_X1 U5668 ( .C1(n6273), .C2(n4850), .A(n4569), .B(n4568), .ZN(U3034)
         );
  AOI22_X1 U5669 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4577), .B1(n6238), 
        .B2(n4576), .ZN(n4571) );
  AOI22_X1 U5670 ( .A1(n5947), .A2(n6240), .B1(n6239), .B2(n4578), .ZN(n4570)
         );
  OAI211_X1 U5671 ( .C1(n6243), .C2(n4850), .A(n4571), .B(n4570), .ZN(U3029)
         );
  AOI22_X1 U5672 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4577), .B1(n6250), 
        .B2(n4576), .ZN(n4573) );
  AOI22_X1 U5673 ( .A1(n5947), .A2(n6252), .B1(n6251), .B2(n4578), .ZN(n4572)
         );
  OAI211_X1 U5674 ( .C1(n6255), .C2(n4850), .A(n4573), .B(n4572), .ZN(U3031)
         );
  AOI22_X1 U5675 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4577), .B1(n6222), 
        .B2(n4576), .ZN(n4575) );
  AOI22_X1 U5676 ( .A1(n5947), .A2(n6234), .B1(n6223), .B2(n4578), .ZN(n4574)
         );
  OAI211_X1 U5677 ( .C1(n6237), .C2(n4850), .A(n4575), .B(n4574), .ZN(U3028)
         );
  AOI22_X1 U5678 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4577), .B1(n6275), 
        .B2(n4576), .ZN(n4580) );
  AOI22_X1 U5679 ( .A1(n5947), .A2(n6279), .B1(n6277), .B2(n4578), .ZN(n4579)
         );
  OAI211_X1 U5680 ( .C1(n6284), .C2(n4850), .A(n4580), .B(n4579), .ZN(U3035)
         );
  NOR2_X1 U5681 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4581), .ZN(n5984)
         );
  INV_X1 U5682 ( .A(n5984), .ZN(n4609) );
  AND2_X1 U5683 ( .A1(n4589), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5997) );
  INV_X1 U5684 ( .A(n4888), .ZN(n4582) );
  OR2_X1 U5685 ( .A1(n6186), .A2(n4582), .ZN(n5923) );
  INV_X1 U5686 ( .A(n5923), .ZN(n4590) );
  OAI21_X1 U5687 ( .B1(n4590), .B2(n6442), .A(n4634), .ZN(n5924) );
  AOI211_X1 U5688 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4609), .A(n5997), .B(
        n5924), .ZN(n4587) );
  NOR2_X1 U5689 ( .A1(n4077), .A2(n4469), .ZN(n4818) );
  INV_X1 U5690 ( .A(n6064), .ZN(n4583) );
  NAND2_X1 U5691 ( .A1(n4818), .A2(n4583), .ZN(n5990) );
  NOR3_X1 U5692 ( .A1(n5977), .A2(n5986), .A3(n6221), .ZN(n4585) );
  OAI21_X1 U5693 ( .B1(n4585), .B2(n6228), .A(n4584), .ZN(n4586) );
  NAND2_X1 U5694 ( .A1(n4587), .A2(n4586), .ZN(n5987) );
  NAND2_X1 U5695 ( .A1(n5987), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4593) );
  INV_X1 U5696 ( .A(n6139), .ZN(n4588) );
  NOR2_X1 U5697 ( .A1(n4588), .A2(n6221), .ZN(n6097) );
  NOR2_X1 U5698 ( .A1(n4589), .A2(n6442), .ZN(n6187) );
  AOI22_X1 U5699 ( .A1(n6097), .A2(n6189), .B1(n6187), .B2(n4590), .ZN(n5983)
         );
  INV_X1 U5700 ( .A(n6275), .ZN(n6183) );
  OAI22_X1 U5701 ( .A1(n4837), .A2(n4609), .B1(n5983), .B2(n6183), .ZN(n4591)
         );
  AOI21_X1 U5702 ( .B1(n6279), .B2(n5977), .A(n4591), .ZN(n4592) );
  OAI211_X1 U5703 ( .C1(n4613), .C2(n6284), .A(n4593), .B(n4592), .ZN(U3059)
         );
  NAND2_X1 U5704 ( .A1(n5987), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4596) );
  INV_X1 U5705 ( .A(n6249), .ZN(n6157) );
  INV_X1 U5706 ( .A(n6246), .ZN(n6117) );
  OAI22_X1 U5707 ( .A1(n6117), .A2(n5990), .B1(n4914), .B2(n4609), .ZN(n4594)
         );
  AOI21_X1 U5708 ( .B1(n6157), .B2(n5986), .A(n4594), .ZN(n4595) );
  OAI211_X1 U5709 ( .C1(n5983), .C2(n6160), .A(n4596), .B(n4595), .ZN(U3054)
         );
  NAND2_X1 U5710 ( .A1(n5987), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4599) );
  INV_X1 U5711 ( .A(n6261), .ZN(n6165) );
  INV_X1 U5712 ( .A(n6258), .ZN(n6123) );
  OAI22_X1 U5713 ( .A1(n6123), .A2(n5990), .B1(n4897), .B2(n4609), .ZN(n4597)
         );
  AOI21_X1 U5714 ( .B1(n6165), .B2(n5986), .A(n4597), .ZN(n4598) );
  OAI211_X1 U5715 ( .C1(n5983), .C2(n6168), .A(n4599), .B(n4598), .ZN(U3056)
         );
  NAND2_X1 U5716 ( .A1(n5987), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4602) );
  INV_X1 U5717 ( .A(n6238), .ZN(n6156) );
  OAI22_X1 U5718 ( .A1(n4905), .A2(n4609), .B1(n5983), .B2(n6156), .ZN(n4600)
         );
  AOI21_X1 U5719 ( .B1(n6240), .B2(n5977), .A(n4600), .ZN(n4601) );
  OAI211_X1 U5720 ( .C1(n4613), .C2(n6243), .A(n4602), .B(n4601), .ZN(U3053)
         );
  NAND2_X1 U5721 ( .A1(n5987), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4605) );
  INV_X1 U5722 ( .A(n6267), .ZN(n6169) );
  INV_X1 U5723 ( .A(n6264), .ZN(n6126) );
  OAI22_X1 U5724 ( .A1(n6126), .A2(n5990), .B1(n4919), .B2(n4609), .ZN(n4603)
         );
  AOI21_X1 U5725 ( .B1(n6169), .B2(n5986), .A(n4603), .ZN(n4604) );
  OAI211_X1 U5726 ( .C1(n5983), .C2(n6172), .A(n4605), .B(n4604), .ZN(U3057)
         );
  NAND2_X1 U5727 ( .A1(n5987), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4608) );
  INV_X1 U5728 ( .A(n6222), .ZN(n6152) );
  OAI22_X1 U5729 ( .A1(n4909), .A2(n4609), .B1(n5983), .B2(n6152), .ZN(n4606)
         );
  AOI21_X1 U5730 ( .B1(n6234), .B2(n5977), .A(n4606), .ZN(n4607) );
  OAI211_X1 U5731 ( .C1(n4613), .C2(n6237), .A(n4608), .B(n4607), .ZN(U3052)
         );
  NAND2_X1 U5732 ( .A1(n5987), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4612) );
  INV_X1 U5733 ( .A(n6250), .ZN(n6164) );
  OAI22_X1 U5734 ( .A1(n4901), .A2(n4609), .B1(n5983), .B2(n6164), .ZN(n4610)
         );
  AOI21_X1 U5735 ( .B1(n6252), .B2(n5977), .A(n4610), .ZN(n4611) );
  OAI211_X1 U5736 ( .C1(n4613), .C2(n6255), .A(n4612), .B(n4611), .ZN(U3055)
         );
  XNOR2_X1 U5737 ( .A(n4614), .B(n4615), .ZN(n4774) );
  OAI222_X1 U5738 ( .A1(n5534), .A2(n4774), .B1(n5249), .B2(n4616), .C1(n5248), 
        .C2(n3450), .ZN(U2884) );
  AOI21_X1 U5739 ( .B1(n4618), .B2(n4617), .A(n4670), .ZN(n5869) );
  INV_X1 U5740 ( .A(n5869), .ZN(n4620) );
  INV_X1 U5741 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4619) );
  OAI222_X1 U5742 ( .A1(n4620), .A2(n5225), .B1(n4619), .B2(n5763), .C1(n5759), 
        .C2(n4774), .ZN(U2852) );
  OR2_X1 U5743 ( .A1(n4622), .A2(n4621), .ZN(n4623) );
  NAND2_X1 U5744 ( .A1(n4624), .A2(n4623), .ZN(n5818) );
  NOR2_X1 U5745 ( .A1(n5887), .A2(n5690), .ZN(n4629) );
  AOI21_X1 U5746 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n5911) );
  NAND2_X1 U5747 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5891) );
  NOR2_X1 U5748 ( .A1(n5911), .A2(n5891), .ZN(n5872) );
  NAND2_X1 U5749 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n5872), .ZN(n4803)
         );
  NOR2_X1 U5750 ( .A1(n4073), .A2(n4980), .ZN(n5906) );
  AOI21_X1 U5751 ( .B1(n5916), .B2(n5906), .A(n5912), .ZN(n5890) );
  NOR2_X1 U5752 ( .A1(n4803), .A2(n5890), .ZN(n4627) );
  NAND2_X1 U5753 ( .A1(n5459), .A2(n5463), .ZN(n5848) );
  NOR2_X1 U5754 ( .A1(n4625), .A2(n4960), .ZN(n5430) );
  OAI22_X1 U5755 ( .A1(n5430), .A2(n5906), .B1(n5912), .B2(n4807), .ZN(n5913)
         );
  AOI21_X1 U5756 ( .B1(n4803), .B2(n5848), .A(n5913), .ZN(n5884) );
  INV_X1 U5757 ( .A(n5884), .ZN(n4626) );
  MUX2_X1 U5758 ( .A(n4627), .B(n4626), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n4628) );
  AOI211_X1 U5759 ( .C1(n5910), .C2(REIP_REG_6__SCAN_IN), .A(n4629), .B(n4628), 
        .ZN(n4630) );
  OAI21_X1 U5760 ( .B1(n5846), .B2(n5818), .A(n4630), .ZN(U3012) );
  NAND2_X1 U5761 ( .A1(n4472), .A2(n6143), .ZN(n6185) );
  NAND2_X1 U5762 ( .A1(n4687), .A2(n6101), .ZN(n4631) );
  NAND2_X1 U5763 ( .A1(n6096), .A2(n4713), .ZN(n4632) );
  AOI21_X1 U5764 ( .B1(n4632), .B2(STATEBS16_REG_SCAN_IN), .A(n6221), .ZN(
        n4636) );
  AND2_X1 U5765 ( .A1(n4447), .A2(n5992), .ZN(n4819) );
  AND2_X1 U5766 ( .A1(n4819), .A2(n2971), .ZN(n6069) );
  INV_X1 U5767 ( .A(n5997), .ZN(n6105) );
  NOR2_X1 U5768 ( .A1(n6105), .A2(n6313), .ZN(n4633) );
  AOI22_X1 U5769 ( .A1(n4636), .A2(n6069), .B1(n6186), .B2(n4633), .ZN(n4664)
         );
  OAI21_X1 U5770 ( .B1(n6186), .B2(n6442), .A(n4634), .ZN(n5996) );
  NOR2_X1 U5771 ( .A1(n6187), .A2(n5996), .ZN(n4822) );
  INV_X1 U5772 ( .A(n6069), .ZN(n4635) );
  NAND3_X1 U5773 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6305), .ZN(n6072) );
  OR2_X1 U5774 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6072), .ZN(n4660)
         );
  AOI22_X1 U5775 ( .A1(n4636), .A2(n4635), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n4660), .ZN(n4637) );
  NAND2_X1 U5776 ( .A1(n4659), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4640)
         );
  INV_X1 U5777 ( .A(n6237), .ZN(n6145) );
  INV_X1 U5778 ( .A(n6234), .ZN(n6111) );
  OAI22_X1 U5779 ( .A1(n4660), .A2(n4909), .B1(n4713), .B2(n6111), .ZN(n4638)
         );
  AOI21_X1 U5780 ( .B1(n6087), .B2(n6145), .A(n4638), .ZN(n4639) );
  OAI211_X1 U5781 ( .C1(n4664), .C2(n6152), .A(n4640), .B(n4639), .ZN(U3100)
         );
  NAND2_X1 U5782 ( .A1(n4659), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4643)
         );
  INV_X1 U5783 ( .A(n6284), .ZN(n6178) );
  INV_X1 U5784 ( .A(n6279), .ZN(n6136) );
  OAI22_X1 U5785 ( .A1(n4660), .A2(n4837), .B1(n4713), .B2(n6136), .ZN(n4641)
         );
  AOI21_X1 U5786 ( .B1(n6087), .B2(n6178), .A(n4641), .ZN(n4642) );
  OAI211_X1 U5787 ( .C1(n4664), .C2(n6183), .A(n4643), .B(n4642), .ZN(U3107)
         );
  NAND2_X1 U5788 ( .A1(n4659), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4646)
         );
  OAI22_X1 U5789 ( .A1(n4660), .A2(n4919), .B1(n4713), .B2(n6126), .ZN(n4644)
         );
  AOI21_X1 U5790 ( .B1(n6087), .B2(n6169), .A(n4644), .ZN(n4645) );
  OAI211_X1 U5791 ( .C1(n4664), .C2(n6172), .A(n4646), .B(n4645), .ZN(U3105)
         );
  NAND2_X1 U5792 ( .A1(n4659), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4649)
         );
  OAI22_X1 U5793 ( .A1(n4660), .A2(n4897), .B1(n4713), .B2(n6123), .ZN(n4647)
         );
  AOI21_X1 U5794 ( .B1(n6087), .B2(n6165), .A(n4647), .ZN(n4648) );
  OAI211_X1 U5795 ( .C1(n4664), .C2(n6168), .A(n4649), .B(n4648), .ZN(U3104)
         );
  NAND2_X1 U5796 ( .A1(n4659), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4652)
         );
  INV_X1 U5797 ( .A(n6273), .ZN(n6173) );
  INV_X1 U5798 ( .A(n6270), .ZN(n6129) );
  OAI22_X1 U5799 ( .A1(n4660), .A2(n4842), .B1(n4713), .B2(n6129), .ZN(n4650)
         );
  AOI21_X1 U5800 ( .B1(n6087), .B2(n6173), .A(n4650), .ZN(n4651) );
  OAI211_X1 U5801 ( .C1(n4664), .C2(n6176), .A(n4652), .B(n4651), .ZN(U3106)
         );
  NAND2_X1 U5802 ( .A1(n4659), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4655)
         );
  INV_X1 U5803 ( .A(n6243), .ZN(n6153) );
  INV_X1 U5804 ( .A(n6240), .ZN(n6114) );
  OAI22_X1 U5805 ( .A1(n4660), .A2(n4905), .B1(n4713), .B2(n6114), .ZN(n4653)
         );
  AOI21_X1 U5806 ( .B1(n6087), .B2(n6153), .A(n4653), .ZN(n4654) );
  OAI211_X1 U5807 ( .C1(n4664), .C2(n6156), .A(n4655), .B(n4654), .ZN(U3101)
         );
  NAND2_X1 U5808 ( .A1(n4659), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4658)
         );
  OAI22_X1 U5809 ( .A1(n4660), .A2(n4914), .B1(n4713), .B2(n6117), .ZN(n4656)
         );
  AOI21_X1 U5810 ( .B1(n6087), .B2(n6157), .A(n4656), .ZN(n4657) );
  OAI211_X1 U5811 ( .C1(n4664), .C2(n6160), .A(n4658), .B(n4657), .ZN(U3102)
         );
  NAND2_X1 U5812 ( .A1(n4659), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4663)
         );
  INV_X1 U5813 ( .A(n6255), .ZN(n6161) );
  INV_X1 U5814 ( .A(n6252), .ZN(n6120) );
  OAI22_X1 U5815 ( .A1(n4660), .A2(n4901), .B1(n4713), .B2(n6120), .ZN(n4661)
         );
  AOI21_X1 U5816 ( .B1(n6087), .B2(n6161), .A(n4661), .ZN(n4662) );
  OAI211_X1 U5817 ( .C1(n4664), .C2(n6164), .A(n4663), .B(n4662), .ZN(U3103)
         );
  NOR2_X1 U5818 ( .A1(n4666), .A2(n4667), .ZN(n4668) );
  OR2_X1 U5819 ( .A1(n4665), .A2(n4668), .ZN(n4795) );
  INV_X1 U5820 ( .A(DATAI_8_), .ZN(n4669) );
  OAI222_X1 U5821 ( .A1(n4795), .A2(n5534), .B1(n5249), .B2(n4669), .C1(n5248), 
        .C2(n6489), .ZN(U2883) );
  INV_X1 U5822 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6571) );
  OAI21_X1 U5823 ( .B1(n4671), .B2(n4670), .A(n4731), .ZN(n4802) );
  OAI222_X1 U5824 ( .A1(n4795), .A2(n5759), .B1(n5763), .B2(n6571), .C1(n4802), 
        .C2(n5225), .ZN(U2851) );
  AOI21_X1 U5825 ( .B1(n5823), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4672), 
        .ZN(n4673) );
  OAI21_X1 U5826 ( .B1(n5840), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4673), 
        .ZN(n4674) );
  AOI21_X1 U5827 ( .B1(n5752), .B2(n5563), .A(n4674), .ZN(n4675) );
  OAI21_X1 U5828 ( .B1(n4676), .B2(n5817), .A(n4675), .ZN(U2985) );
  OAI21_X1 U5829 ( .B1(n4665), .B2(n4678), .A(n4677), .ZN(n5681) );
  AOI22_X1 U5830 ( .A1(n5250), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n5773), .ZN(n4679) );
  OAI21_X1 U5831 ( .B1(n5681), .B2(n5534), .A(n4679), .ZN(U2882) );
  OAI21_X1 U5832 ( .B1(n4682), .B2(n4681), .A(n4680), .ZN(n5864) );
  INV_X1 U5833 ( .A(n4774), .ZN(n4685) );
  AOI22_X1 U5834 ( .A1(n5823), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .B1(n5910), 
        .B2(REIP_REG_7__SCAN_IN), .ZN(n4683) );
  OAI21_X1 U5835 ( .B1(n5840), .B2(n4769), .A(n4683), .ZN(n4684) );
  AOI21_X1 U5836 ( .B1(n4685), .B2(n5563), .A(n4684), .ZN(n4686) );
  OAI21_X1 U5837 ( .B1(n5864), .B2(n5817), .A(n4686), .ZN(U2979) );
  INV_X1 U5838 ( .A(n6065), .ZN(n6068) );
  NAND3_X1 U5839 ( .A1(n6068), .A2(n4687), .A3(STATEBS16_REG_SCAN_IN), .ZN(
        n4688) );
  NAND2_X1 U5840 ( .A1(n4688), .A2(n6232), .ZN(n4692) );
  AND2_X1 U5841 ( .A1(n2971), .A2(n6296), .ZN(n6218) );
  NAND3_X1 U5842 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6305), .A3(n6301), .ZN(n4893) );
  NOR2_X1 U5843 ( .A1(n6138), .A2(n4893), .ZN(n4710) );
  AOI21_X1 U5844 ( .B1(n6218), .B2(n4886), .A(n4710), .ZN(n4693) );
  INV_X1 U5845 ( .A(n4693), .ZN(n4691) );
  AOI21_X1 U5846 ( .B1(n6221), .B2(n4893), .A(n4689), .ZN(n4690) );
  OAI21_X1 U5847 ( .B1(n4692), .B2(n4691), .A(n4690), .ZN(n4709) );
  OAI22_X1 U5848 ( .A1(n4693), .A2(n4692), .B1(n6442), .B2(n4893), .ZN(n4708)
         );
  AOI22_X1 U5849 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4709), .B1(n6238), 
        .B2(n4708), .ZN(n4695) );
  NOR3_X4 U5850 ( .A1(n6065), .A2(n6101), .A3(n4472), .ZN(n6059) );
  AOI22_X1 U5851 ( .A1(n6059), .A2(n6240), .B1(n6239), .B2(n4710), .ZN(n4694)
         );
  OAI211_X1 U5852 ( .C1(n4713), .C2(n6243), .A(n4695), .B(n4694), .ZN(U3093)
         );
  AOI22_X1 U5853 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4709), .B1(n6257), 
        .B2(n4708), .ZN(n4697) );
  AOI22_X1 U5854 ( .A1(n6059), .A2(n6258), .B1(n6256), .B2(n4710), .ZN(n4696)
         );
  OAI211_X1 U5855 ( .C1(n4713), .C2(n6261), .A(n4697), .B(n4696), .ZN(U3096)
         );
  AOI22_X1 U5856 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4709), .B1(n6263), 
        .B2(n4708), .ZN(n4699) );
  AOI22_X1 U5857 ( .A1(n6059), .A2(n6264), .B1(n6262), .B2(n4710), .ZN(n4698)
         );
  OAI211_X1 U5858 ( .C1(n4713), .C2(n6267), .A(n4699), .B(n4698), .ZN(U3097)
         );
  AOI22_X1 U5859 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4709), .B1(n6269), 
        .B2(n4708), .ZN(n4701) );
  AOI22_X1 U5860 ( .A1(n6059), .A2(n6270), .B1(n6268), .B2(n4710), .ZN(n4700)
         );
  OAI211_X1 U5861 ( .C1(n4713), .C2(n6273), .A(n4701), .B(n4700), .ZN(U3098)
         );
  AOI22_X1 U5862 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4709), .B1(n6275), 
        .B2(n4708), .ZN(n4703) );
  AOI22_X1 U5863 ( .A1(n6059), .A2(n6279), .B1(n6277), .B2(n4710), .ZN(n4702)
         );
  OAI211_X1 U5864 ( .C1(n4713), .C2(n6284), .A(n4703), .B(n4702), .ZN(U3099)
         );
  AOI22_X1 U5865 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4709), .B1(n6222), 
        .B2(n4708), .ZN(n4705) );
  AOI22_X1 U5866 ( .A1(n6059), .A2(n6234), .B1(n6223), .B2(n4710), .ZN(n4704)
         );
  OAI211_X1 U5867 ( .C1(n4713), .C2(n6237), .A(n4705), .B(n4704), .ZN(U3092)
         );
  AOI22_X1 U5868 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4709), .B1(n6245), 
        .B2(n4708), .ZN(n4707) );
  AOI22_X1 U5869 ( .A1(n6059), .A2(n6246), .B1(n6244), .B2(n4710), .ZN(n4706)
         );
  OAI211_X1 U5870 ( .C1(n4713), .C2(n6249), .A(n4707), .B(n4706), .ZN(U3094)
         );
  AOI22_X1 U5871 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4709), .B1(n6250), 
        .B2(n4708), .ZN(n4712) );
  AOI22_X1 U5872 ( .A1(n6059), .A2(n6252), .B1(n6251), .B2(n4710), .ZN(n4711)
         );
  OAI211_X1 U5873 ( .C1(n4713), .C2(n6255), .A(n4712), .B(n4711), .ZN(U3095)
         );
  INV_X1 U5874 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5061) );
  AND3_X1 U5875 ( .A1(n4715), .A2(n5061), .A3(n4714), .ZN(n4716) );
  AOI21_X1 U5876 ( .B1(n2954), .B2(n6319), .A(n4716), .ZN(n4717) );
  NAND2_X1 U5877 ( .A1(n4718), .A2(n4781), .ZN(n4723) );
  INV_X1 U5878 ( .A(n4798), .ZN(n4721) );
  NAND2_X1 U5879 ( .A1(n5745), .A2(n4721), .ZN(n4722) );
  OAI21_X1 U5880 ( .B1(n5711), .B2(n4723), .A(n4722), .ZN(n4728) );
  NAND2_X1 U5881 ( .A1(n5734), .A2(n4781), .ZN(n4724) );
  AND2_X1 U5882 ( .A1(n4724), .A2(n5735), .ZN(n5679) );
  INV_X1 U5883 ( .A(n5679), .ZN(n4725) );
  AOI22_X1 U5884 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n5743), .B1(
        REIP_REG_8__SCAN_IN), .B2(n4725), .ZN(n4726) );
  NAND2_X1 U5885 ( .A1(n6450), .A2(n5735), .ZN(n5702) );
  OAI211_X1 U5886 ( .C1(n5755), .C2(n4802), .A(n4726), .B(n5702), .ZN(n4727)
         );
  AOI211_X1 U5887 ( .C1(EBX_REG_8__SCAN_IN), .C2(n5746), .A(n4728), .B(n4727), 
        .ZN(n4729) );
  OAI21_X1 U5888 ( .B1(n5673), .B2(n4795), .A(n4729), .ZN(U2819) );
  AOI21_X1 U5889 ( .B1(n4732), .B2(n4731), .A(n4730), .ZN(n5858) );
  INV_X1 U5890 ( .A(n5858), .ZN(n4734) );
  OAI222_X1 U5891 ( .A1(n4734), .A2(n5225), .B1(n4733), .B2(n5763), .C1(n5681), 
        .C2(n5759), .ZN(U2850) );
  OAI21_X1 U5892 ( .B1(n4735), .B2(n4737), .A(n4736), .ZN(n5898) );
  NAND2_X1 U5893 ( .A1(n5910), .A2(REIP_REG_3__SCAN_IN), .ZN(n5895) );
  OAI21_X1 U5894 ( .B1(n5323), .B2(n4738), .A(n5895), .ZN(n4740) );
  NOR2_X1 U5895 ( .A1(n5723), .A2(n6225), .ZN(n4739) );
  AOI211_X1 U5896 ( .C1(n5558), .C2(n5725), .A(n4740), .B(n4739), .ZN(n4741)
         );
  OAI21_X1 U5897 ( .B1(n5817), .B2(n5898), .A(n4741), .ZN(U2983) );
  OAI21_X1 U5898 ( .B1(n4744), .B2(n4743), .A(n4742), .ZN(n5876) );
  NAND2_X1 U5899 ( .A1(n5910), .A2(REIP_REG_5__SCAN_IN), .ZN(n5873) );
  OAI21_X1 U5900 ( .B1(n5323), .B2(n4745), .A(n5873), .ZN(n4747) );
  NOR2_X1 U5901 ( .A1(n5699), .A2(n6225), .ZN(n4746) );
  AOI211_X1 U5902 ( .C1(n5558), .C2(n5700), .A(n4747), .B(n4746), .ZN(n4748)
         );
  OAI21_X1 U5903 ( .B1(n5817), .B2(n5876), .A(n4748), .ZN(U2981) );
  INV_X1 U5904 ( .A(n4749), .ZN(n4750) );
  NOR2_X1 U5905 ( .A1(n4754), .A2(n4750), .ZN(n4751) );
  OR2_X1 U5906 ( .A1(n4751), .A2(n5692), .ZN(n5751) );
  INV_X1 U5907 ( .A(n5751), .ZN(n5722) );
  NAND2_X1 U5908 ( .A1(n5678), .A2(n5717), .ZN(n4758) );
  INV_X1 U5909 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6436) );
  OAI22_X1 U5910 ( .A1(n5525), .A2(n6436), .B1(n5741), .B2(n4752), .ZN(n4757)
         );
  NOR2_X1 U5911 ( .A1(n4754), .A2(n4753), .ZN(n5730) );
  INV_X1 U5912 ( .A(n5730), .ZN(n5749) );
  OAI22_X1 U5913 ( .A1(n5749), .A2(n3342), .B1(n5755), .B2(n4755), .ZN(n4756)
         );
  AOI211_X1 U5914 ( .C1(PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n4758), .A(n4757), 
        .B(n4756), .ZN(n4759) );
  OAI21_X1 U5915 ( .B1(n4760), .B2(n5722), .A(n4759), .ZN(U2827) );
  NAND2_X1 U5916 ( .A1(n5734), .A2(n4761), .ZN(n5695) );
  INV_X1 U5917 ( .A(n5695), .ZN(n4762) );
  NAND2_X1 U5918 ( .A1(n4762), .A2(REIP_REG_5__SCAN_IN), .ZN(n4767) );
  NOR3_X1 U5919 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6367), .A3(n4767), .ZN(n4772)
         );
  INV_X1 U5920 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4764) );
  AOI22_X1 U5921 ( .A1(EBX_REG_7__SCAN_IN), .A2(n5746), .B1(n5698), .B2(n5869), 
        .ZN(n4763) );
  OAI211_X1 U5922 ( .C1(n5678), .C2(n4764), .A(n4763), .B(n5702), .ZN(n4771)
         );
  INV_X1 U5923 ( .A(n4765), .ZN(n4766) );
  OAI21_X1 U5924 ( .B1(n5711), .B2(n4766), .A(n5735), .ZN(n5697) );
  NOR2_X1 U5925 ( .A1(REIP_REG_6__SCAN_IN), .A2(n4767), .ZN(n5687) );
  OAI21_X1 U5926 ( .B1(n5697), .B2(n5687), .A(REIP_REG_7__SCAN_IN), .ZN(n4768)
         );
  OAI21_X1 U5927 ( .B1(n5717), .B2(n4769), .A(n4768), .ZN(n4770) );
  NOR3_X1 U5928 ( .A1(n4772), .A2(n4771), .A3(n4770), .ZN(n4773) );
  OAI21_X1 U5929 ( .B1(n4774), .B2(n5673), .A(n4773), .ZN(U2820) );
  INV_X1 U5930 ( .A(n4775), .ZN(n4776) );
  AOI21_X1 U5931 ( .B1(n4777), .B2(n4677), .A(n4776), .ZN(n4929) );
  INV_X1 U5932 ( .A(n4929), .ZN(n4788) );
  INV_X1 U5933 ( .A(n4927), .ZN(n4785) );
  INV_X1 U5934 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6371) );
  INV_X1 U5935 ( .A(n5702), .ZN(n5708) );
  INV_X1 U5936 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6471) );
  OR2_X1 U5937 ( .A1(n4778), .A2(n4730), .ZN(n4779) );
  NAND2_X1 U5938 ( .A1(n4779), .A2(n5666), .ZN(n5849) );
  OAI22_X1 U5939 ( .A1(n6471), .A2(n5678), .B1(n5755), .B2(n5849), .ZN(n4780)
         );
  AOI211_X1 U5940 ( .C1(EBX_REG_10__SCAN_IN), .C2(n5746), .A(n5708), .B(n4780), 
        .ZN(n4783) );
  NOR2_X1 U5941 ( .A1(n5711), .A2(n4781), .ZN(n5677) );
  OAI211_X1 U5942 ( .C1(REIP_REG_9__SCAN_IN), .C2(REIP_REG_10__SCAN_IN), .A(
        n5677), .B(n5663), .ZN(n4782) );
  OAI211_X1 U5943 ( .C1(n5679), .C2(n6371), .A(n4783), .B(n4782), .ZN(n4784)
         );
  AOI21_X1 U5944 ( .B1(n5745), .B2(n4785), .A(n4784), .ZN(n4786) );
  OAI21_X1 U5945 ( .B1(n4788), .B2(n5673), .A(n4786), .ZN(U2817) );
  AOI22_X1 U5946 ( .A1(n5250), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n5773), .ZN(n4787) );
  OAI21_X1 U5947 ( .B1(n4788), .B2(n5534), .A(n4787), .ZN(U2881) );
  OAI22_X1 U5948 ( .A1(n5758), .A2(n5849), .B1(n5763), .B2(n4789), .ZN(n4790)
         );
  AOI21_X1 U5949 ( .B1(n4929), .B2(n5211), .A(n4790), .ZN(n4791) );
  INV_X1 U5950 ( .A(n4791), .ZN(U2849) );
  OAI21_X1 U5951 ( .B1(n4794), .B2(n4793), .A(n4792), .ZN(n4816) );
  INV_X1 U5952 ( .A(n4795), .ZN(n4800) );
  INV_X1 U5953 ( .A(REIP_REG_8__SCAN_IN), .ZN(n4796) );
  NOR2_X1 U5954 ( .A1(n5885), .A2(n4796), .ZN(n4813) );
  AOI21_X1 U5955 ( .B1(n5823), .B2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n4813), 
        .ZN(n4797) );
  OAI21_X1 U5956 ( .B1(n5840), .B2(n4798), .A(n4797), .ZN(n4799) );
  AOI21_X1 U5957 ( .B1(n4800), .B2(n5563), .A(n4799), .ZN(n4801) );
  OAI21_X1 U5958 ( .B1(n4816), .B2(n5817), .A(n4801), .ZN(U2978) );
  INV_X1 U5959 ( .A(n4802), .ZN(n4814) );
  NOR2_X1 U5960 ( .A1(n4805), .A2(n4803), .ZN(n4808) );
  INV_X1 U5961 ( .A(n5890), .ZN(n4804) );
  NAND2_X1 U5962 ( .A1(n4808), .A2(n4804), .ZN(n5852) );
  NOR2_X1 U5963 ( .A1(n4955), .A2(n5852), .ZN(n4811) );
  NOR2_X1 U5964 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n5852), .ZN(n5867)
         );
  NAND3_X1 U5965 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n5906), .ZN(n5877) );
  NOR3_X1 U5966 ( .A1(n4806), .A2(n4805), .A3(n5877), .ZN(n4958) );
  NAND2_X1 U5967 ( .A1(n4807), .A2(n4996), .ZN(n5432) );
  INV_X1 U5968 ( .A(n5432), .ZN(n4809) );
  OAI22_X1 U5969 ( .A1(n5430), .A2(n4958), .B1(n4809), .B2(n4956), .ZN(n5865)
         );
  OR2_X1 U5970 ( .A1(n5867), .A2(n5865), .ZN(n4810) );
  MUX2_X1 U5971 ( .A(n4811), .B(n4810), .S(INSTADDRPOINTER_REG_8__SCAN_IN), 
        .Z(n4812) );
  AOI211_X1 U5972 ( .C1(n5908), .C2(n4814), .A(n4813), .B(n4812), .ZN(n4815)
         );
  OAI21_X1 U5973 ( .B1(n5846), .B2(n4816), .A(n4815), .ZN(U3010) );
  NAND3_X1 U5974 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6313), .A3(n6305), .ZN(n5958) );
  NOR2_X1 U5975 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5958), .ZN(n4824)
         );
  INV_X1 U5976 ( .A(n6185), .ZN(n4817) );
  OAI21_X1 U5977 ( .B1(n4857), .B2(n5965), .A(n4891), .ZN(n4821) );
  INV_X1 U5978 ( .A(n5954), .ZN(n4820) );
  NAND2_X1 U5979 ( .A1(n4821), .A2(n4820), .ZN(n4823) );
  NAND2_X1 U5980 ( .A1(n4854), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4829) );
  INV_X1 U5981 ( .A(n4824), .ZN(n4855) );
  NAND2_X1 U5982 ( .A1(n5954), .A2(n6232), .ZN(n4826) );
  NAND3_X1 U5983 ( .A1(n5997), .A2(n6186), .A3(n6313), .ZN(n4825) );
  OAI22_X1 U5984 ( .A1(n4909), .A2(n4855), .B1(n4860), .B2(n6152), .ZN(n4827)
         );
  AOI21_X1 U5985 ( .B1(n6145), .B2(n5965), .A(n4827), .ZN(n4828) );
  OAI211_X1 U5986 ( .C1(n6111), .C2(n4850), .A(n4829), .B(n4828), .ZN(U3036)
         );
  NAND2_X1 U5987 ( .A1(n4854), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4833) );
  OAI22_X1 U5988 ( .A1(n4901), .A2(n4855), .B1(n4860), .B2(n6164), .ZN(n4831)
         );
  NOR2_X1 U5989 ( .A1(n5982), .A2(n6255), .ZN(n4830) );
  NOR2_X1 U5990 ( .A1(n4831), .A2(n4830), .ZN(n4832) );
  OAI211_X1 U5991 ( .C1(n4850), .C2(n6120), .A(n4833), .B(n4832), .ZN(U3039)
         );
  NAND2_X1 U5992 ( .A1(n4854), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4836) );
  OAI22_X1 U5993 ( .A1(n6267), .A2(n5982), .B1(n4919), .B2(n4855), .ZN(n4834)
         );
  AOI21_X1 U5994 ( .B1(n6264), .B2(n4857), .A(n4834), .ZN(n4835) );
  OAI211_X1 U5995 ( .C1(n4860), .C2(n6172), .A(n4836), .B(n4835), .ZN(U3041)
         );
  NAND2_X1 U5996 ( .A1(n4854), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4841) );
  OAI22_X1 U5997 ( .A1(n4837), .A2(n4855), .B1(n4860), .B2(n6183), .ZN(n4839)
         );
  NOR2_X1 U5998 ( .A1(n5982), .A2(n6284), .ZN(n4838) );
  NOR2_X1 U5999 ( .A1(n4839), .A2(n4838), .ZN(n4840) );
  OAI211_X1 U6000 ( .C1(n4850), .C2(n6136), .A(n4841), .B(n4840), .ZN(U3043)
         );
  NAND2_X1 U6001 ( .A1(n4854), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4845) );
  OAI22_X1 U6002 ( .A1(n6273), .A2(n5982), .B1(n4842), .B2(n4855), .ZN(n4843)
         );
  AOI21_X1 U6003 ( .B1(n6270), .B2(n4857), .A(n4843), .ZN(n4844) );
  OAI211_X1 U6004 ( .C1(n4860), .C2(n6176), .A(n4845), .B(n4844), .ZN(U3042)
         );
  NAND2_X1 U6005 ( .A1(n4854), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4849) );
  OAI22_X1 U6006 ( .A1(n4905), .A2(n4855), .B1(n4860), .B2(n6156), .ZN(n4847)
         );
  NOR2_X1 U6007 ( .A1(n5982), .A2(n6243), .ZN(n4846) );
  NOR2_X1 U6008 ( .A1(n4847), .A2(n4846), .ZN(n4848) );
  OAI211_X1 U6009 ( .C1(n4850), .C2(n6114), .A(n4849), .B(n4848), .ZN(U3037)
         );
  NAND2_X1 U6010 ( .A1(n4854), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4853) );
  OAI22_X1 U6011 ( .A1(n6261), .A2(n5982), .B1(n4897), .B2(n4855), .ZN(n4851)
         );
  AOI21_X1 U6012 ( .B1(n6258), .B2(n4857), .A(n4851), .ZN(n4852) );
  OAI211_X1 U6013 ( .C1(n4860), .C2(n6168), .A(n4853), .B(n4852), .ZN(U3040)
         );
  NAND2_X1 U6014 ( .A1(n4854), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4859) );
  OAI22_X1 U6015 ( .A1(n6249), .A2(n5982), .B1(n4914), .B2(n4855), .ZN(n4856)
         );
  AOI21_X1 U6016 ( .B1(n6246), .B2(n4857), .A(n4856), .ZN(n4858) );
  OAI211_X1 U6017 ( .C1(n4860), .C2(n6160), .A(n4859), .B(n4858), .ZN(U3038)
         );
  NAND2_X1 U6018 ( .A1(n4775), .A2(n4862), .ZN(n4863) );
  NAND2_X1 U6019 ( .A1(n4861), .A2(n4863), .ZN(n5812) );
  AOI22_X1 U6020 ( .A1(n5250), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n5773), .ZN(n4864) );
  OAI21_X1 U6021 ( .B1(n5812), .B2(n5534), .A(n4864), .ZN(U2880) );
  NAND2_X1 U6022 ( .A1(n4866), .A2(n4865), .ZN(n4867) );
  XNOR2_X1 U6023 ( .A(n4868), .B(n4867), .ZN(n5860) );
  NAND2_X1 U6024 ( .A1(n5860), .A2(n5835), .ZN(n4871) );
  NAND2_X1 U6025 ( .A1(n5910), .A2(REIP_REG_9__SCAN_IN), .ZN(n5856) );
  OAI21_X1 U6026 ( .B1(n5323), .B2(n6568), .A(n5856), .ZN(n4869) );
  AOI21_X1 U6027 ( .B1(n5558), .B2(n5682), .A(n4869), .ZN(n4870) );
  OAI211_X1 U6028 ( .C1(n6225), .C2(n5681), .A(n4871), .B(n4870), .ZN(U2977)
         );
  XOR2_X1 U6029 ( .A(n4872), .B(n4861), .Z(n4950) );
  OR2_X1 U6030 ( .A1(n4873), .A2(n5665), .ZN(n4874) );
  NAND2_X1 U6031 ( .A1(n4874), .A2(n4937), .ZN(n4952) );
  OAI22_X1 U6032 ( .A1(n5758), .A2(n4952), .B1(n5763), .B2(n4878), .ZN(n4875)
         );
  AOI21_X1 U6033 ( .B1(n4950), .B2(n5211), .A(n4875), .ZN(n4876) );
  INV_X1 U6034 ( .A(n4876), .ZN(U2847) );
  INV_X1 U6035 ( .A(n4950), .ZN(n4885) );
  AOI22_X1 U6036 ( .A1(n5250), .A2(DATAI_12_), .B1(EAX_REG_12__SCAN_IN), .B2(
        n5773), .ZN(n4877) );
  OAI21_X1 U6037 ( .B1(n4885), .B2(n5534), .A(n4877), .ZN(U2879) );
  INV_X1 U6038 ( .A(n4948), .ZN(n4883) );
  NAND2_X1 U6039 ( .A1(n5734), .A2(n4879), .ZN(n5656) );
  OAI22_X1 U6040 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5656), .B1(n5741), .B2(
        n4878), .ZN(n4882) );
  OAI21_X1 U6041 ( .B1(n5711), .B2(n4879), .A(n5735), .ZN(n5668) );
  AOI22_X1 U6042 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n5743), .B1(
        REIP_REG_12__SCAN_IN), .B2(n5668), .ZN(n4880) );
  OAI211_X1 U6043 ( .C1(n5755), .C2(n4952), .A(n4880), .B(n5702), .ZN(n4881)
         );
  AOI211_X1 U6044 ( .C1(n5745), .C2(n4883), .A(n4882), .B(n4881), .ZN(n4884)
         );
  OAI21_X1 U6045 ( .B1(n4885), .B2(n5673), .A(n4884), .ZN(U2815) );
  INV_X1 U6046 ( .A(n4886), .ZN(n4887) );
  NOR2_X1 U6047 ( .A1(n4887), .A2(n6189), .ZN(n4890) );
  OR2_X1 U6048 ( .A1(n6186), .A2(n4888), .ZN(n6099) );
  INV_X1 U6049 ( .A(n6099), .ZN(n4889) );
  AOI22_X1 U6050 ( .A1(n4890), .A2(n6232), .B1(n5997), .B2(n4889), .ZN(n6054)
         );
  NAND3_X1 U6051 ( .A1(n4913), .A2(n6232), .A3(n6063), .ZN(n4892) );
  AOI21_X1 U6052 ( .B1(n4892), .B2(n4891), .A(n4890), .ZN(n4896) );
  NOR2_X1 U6053 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4893), .ZN(n6058)
         );
  INV_X1 U6054 ( .A(n6187), .ZN(n6098) );
  AOI21_X1 U6055 ( .B1(n6099), .B2(STATE2_REG_2__SCAN_IN), .A(n4894), .ZN(
        n6104) );
  OAI211_X1 U6056 ( .C1(n6413), .C2(n6058), .A(n6098), .B(n6104), .ZN(n4895)
         );
  NAND2_X1 U6057 ( .A1(n6060), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4900) );
  INV_X1 U6058 ( .A(n6058), .ZN(n4918) );
  OAI22_X1 U6059 ( .A1(n4897), .A2(n4918), .B1(n6123), .B2(n6063), .ZN(n4898)
         );
  AOI21_X1 U6060 ( .B1(n6059), .B2(n6165), .A(n4898), .ZN(n4899) );
  OAI211_X1 U6061 ( .C1(n6054), .C2(n6168), .A(n4900), .B(n4899), .ZN(U3088)
         );
  NAND2_X1 U6062 ( .A1(n6060), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4904) );
  OAI22_X1 U6063 ( .A1(n4901), .A2(n4918), .B1(n6054), .B2(n6164), .ZN(n4902)
         );
  AOI21_X1 U6064 ( .B1(n6252), .B2(n6047), .A(n4902), .ZN(n4903) );
  OAI211_X1 U6065 ( .C1(n4913), .C2(n6255), .A(n4904), .B(n4903), .ZN(U3087)
         );
  NAND2_X1 U6066 ( .A1(n6060), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4908) );
  OAI22_X1 U6067 ( .A1(n4905), .A2(n4918), .B1(n6054), .B2(n6156), .ZN(n4906)
         );
  AOI21_X1 U6068 ( .B1(n6240), .B2(n6047), .A(n4906), .ZN(n4907) );
  OAI211_X1 U6069 ( .C1(n4913), .C2(n6243), .A(n4908), .B(n4907), .ZN(U3085)
         );
  NAND2_X1 U6070 ( .A1(n6060), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4912) );
  OAI22_X1 U6071 ( .A1(n4909), .A2(n4918), .B1(n6054), .B2(n6152), .ZN(n4910)
         );
  AOI21_X1 U6072 ( .B1(n6234), .B2(n6047), .A(n4910), .ZN(n4911) );
  OAI211_X1 U6073 ( .C1(n4913), .C2(n6237), .A(n4912), .B(n4911), .ZN(U3084)
         );
  NAND2_X1 U6074 ( .A1(n6060), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4917) );
  OAI22_X1 U6075 ( .A1(n4914), .A2(n4918), .B1(n6117), .B2(n6063), .ZN(n4915)
         );
  AOI21_X1 U6076 ( .B1(n6059), .B2(n6157), .A(n4915), .ZN(n4916) );
  OAI211_X1 U6077 ( .C1(n6054), .C2(n6160), .A(n4917), .B(n4916), .ZN(U3086)
         );
  NAND2_X1 U6078 ( .A1(n6060), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4922) );
  OAI22_X1 U6079 ( .A1(n4919), .A2(n4918), .B1(n6126), .B2(n6063), .ZN(n4920)
         );
  AOI21_X1 U6080 ( .B1(n6059), .B2(n6169), .A(n4920), .ZN(n4921) );
  OAI211_X1 U6081 ( .C1(n6054), .C2(n6172), .A(n4922), .B(n4921), .ZN(U3089)
         );
  NAND2_X1 U6082 ( .A1(n5806), .A2(n4924), .ZN(n4925) );
  XNOR2_X1 U6083 ( .A(n4923), .B(n4925), .ZN(n5851) );
  INV_X1 U6084 ( .A(n5851), .ZN(n4931) );
  AOI22_X1 U6085 ( .A1(n5823), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n5910), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n4926) );
  OAI21_X1 U6086 ( .B1(n5840), .B2(n4927), .A(n4926), .ZN(n4928) );
  AOI21_X1 U6087 ( .B1(n4929), .B2(n5563), .A(n4928), .ZN(n4930) );
  OAI21_X1 U6088 ( .B1(n4931), .B2(n5817), .A(n4930), .ZN(U2976) );
  NAND2_X1 U6089 ( .A1(n4932), .A2(n4933), .ZN(n4934) );
  AND2_X1 U6090 ( .A1(n4935), .A2(n4934), .ZN(n5659) );
  INV_X1 U6091 ( .A(n5659), .ZN(n4942) );
  AOI22_X1 U6092 ( .A1(n5250), .A2(DATAI_13_), .B1(EAX_REG_13__SCAN_IN), .B2(
        n5773), .ZN(n4936) );
  OAI21_X1 U6093 ( .B1(n4942), .B2(n5534), .A(n4936), .ZN(U2878) );
  AOI21_X1 U6094 ( .B1(n4938), .B2(n4937), .A(n5221), .ZN(n5653) );
  AOI22_X1 U6095 ( .A1(n4940), .A2(n5653), .B1(EBX_REG_13__SCAN_IN), .B2(n4939), .ZN(n4941) );
  OAI21_X1 U6096 ( .B1(n4942), .B2(n5759), .A(n4941), .ZN(U2846) );
  NOR2_X1 U6097 ( .A1(n4944), .A2(n2989), .ZN(n4945) );
  XNOR2_X1 U6098 ( .A(n4943), .B(n4945), .ZN(n4973) );
  INV_X1 U6099 ( .A(REIP_REG_12__SCAN_IN), .ZN(n4946) );
  NOR2_X1 U6100 ( .A1(n5885), .A2(n4946), .ZN(n4953) );
  AOI21_X1 U6101 ( .B1(n5823), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n4953), 
        .ZN(n4947) );
  OAI21_X1 U6102 ( .B1(n5840), .B2(n4948), .A(n4947), .ZN(n4949) );
  AOI21_X1 U6103 ( .B1(n4950), .B2(n5563), .A(n4949), .ZN(n4951) );
  OAI21_X1 U6104 ( .B1(n4973), .B2(n5817), .A(n4951), .ZN(U2974) );
  INV_X1 U6105 ( .A(n4952), .ZN(n4954) );
  AOI21_X1 U6106 ( .B1(n5908), .B2(n4954), .A(n4953), .ZN(n4972) );
  NOR4_X1 U6107 ( .A1(n4955), .A2(n6492), .A3(n6461), .A4(n4129), .ZN(n4957)
         );
  NAND2_X1 U6108 ( .A1(n4957), .A2(n4956), .ZN(n4964) );
  NAND2_X1 U6109 ( .A1(n5432), .A2(n4964), .ZN(n5427) );
  NAND2_X1 U6110 ( .A1(n4958), .A2(n4957), .ZN(n4962) );
  INV_X1 U6111 ( .A(n4962), .ZN(n5429) );
  OR2_X1 U6112 ( .A1(n5430), .A2(n5429), .ZN(n4959) );
  NAND2_X1 U6113 ( .A1(n5427), .A2(n4959), .ZN(n5843) );
  NAND2_X1 U6114 ( .A1(n4960), .A2(n5429), .ZN(n4967) );
  INV_X1 U6115 ( .A(n4967), .ZN(n5595) );
  NOR2_X1 U6116 ( .A1(n4962), .A2(n4961), .ZN(n4965) );
  OR3_X1 U6117 ( .A1(n5912), .A2(n5595), .A3(n4965), .ZN(n4963) );
  NAND2_X1 U6118 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5593) );
  AND2_X1 U6119 ( .A1(n4963), .A2(n5593), .ZN(n4970) );
  INV_X1 U6120 ( .A(n4964), .ZN(n4966) );
  NOR2_X1 U6121 ( .A1(n4966), .A2(n4965), .ZN(n5460) );
  NAND2_X1 U6122 ( .A1(n5460), .A2(n4967), .ZN(n5842) );
  INV_X1 U6123 ( .A(n5842), .ZN(n5586) );
  OAI21_X1 U6124 ( .B1(n5586), .B2(n4131), .A(n4968), .ZN(n4969) );
  OAI21_X1 U6125 ( .B1(n5843), .B2(n4970), .A(n4969), .ZN(n4971) );
  OAI211_X1 U6126 ( .C1(n4973), .C2(n5846), .A(n4972), .B(n4971), .ZN(U3006)
         );
  NAND2_X1 U6127 ( .A1(n6297), .A2(n3062), .ZN(n4978) );
  INV_X1 U6128 ( .A(n4976), .ZN(n6294) );
  OAI21_X1 U6129 ( .B1(n4974), .B2(n4975), .A(n6294), .ZN(n4977) );
  OAI211_X1 U6130 ( .C1(n4496), .C2(n4979), .A(n4978), .B(n4977), .ZN(n6299)
         );
  INV_X1 U6131 ( .A(n6425), .ZN(n5603) );
  INV_X1 U6132 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4981) );
  AOI22_X1 U6133 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4981), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4980), .ZN(n5042) );
  NOR2_X1 U6134 ( .A1(n6538), .A2(n5043), .ZN(n4982) );
  AOI222_X1 U6135 ( .A1(n6299), .A2(n5603), .B1(n5042), .B2(n4982), .C1(n4974), 
        .C2(n6323), .ZN(n4987) );
  NAND2_X1 U6136 ( .A1(n6298), .A2(n6332), .ZN(n4985) );
  INV_X1 U6137 ( .A(n6410), .ZN(n4983) );
  NAND2_X1 U6138 ( .A1(n4983), .A2(FLUSH_REG_SCAN_IN), .ZN(n4984) );
  NAND2_X1 U6139 ( .A1(n4985), .A2(n4984), .ZN(n5602) );
  OAI21_X1 U6140 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6415), .A(n6423), 
        .ZN(n6421) );
  INV_X1 U6141 ( .A(n6421), .ZN(n4986) );
  OAI22_X1 U6142 ( .A1(n4987), .A2(n6418), .B1(n3062), .B2(n4986), .ZN(U3460)
         );
  AOI21_X1 U6143 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n4989), .A(n4988), 
        .ZN(n4991) );
  INV_X1 U6144 ( .A(n5848), .ZN(n5434) );
  NOR2_X1 U6145 ( .A1(n4134), .A2(n5593), .ZN(n5464) );
  NAND2_X1 U6146 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5464), .ZN(n5585) );
  NAND2_X1 U6147 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5579) );
  NOR2_X1 U6148 ( .A1(n5585), .A2(n5579), .ZN(n5428) );
  INV_X1 U6149 ( .A(n5000), .ZN(n5433) );
  NAND3_X1 U6150 ( .A1(n5428), .A2(n5433), .A3(n5435), .ZN(n4992) );
  AND2_X1 U6151 ( .A1(n5848), .A2(n4992), .ZN(n4993) );
  NOR2_X1 U6152 ( .A1(n5843), .A2(n4993), .ZN(n5426) );
  INV_X1 U6153 ( .A(n5410), .ZN(n5392) );
  NAND2_X1 U6154 ( .A1(n5848), .A2(n5392), .ZN(n4994) );
  NAND2_X1 U6155 ( .A1(n5426), .A2(n4994), .ZN(n5406) );
  AOI21_X1 U6156 ( .B1(n5878), .B2(n4996), .A(n4995), .ZN(n4997) );
  NAND2_X1 U6157 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5377) );
  AND2_X1 U6158 ( .A1(n5848), .A2(n5377), .ZN(n4998) );
  AND2_X1 U6159 ( .A1(n5848), .A2(n5358), .ZN(n4999) );
  NOR2_X1 U6160 ( .A1(n5372), .A2(n4999), .ZN(n5036) );
  OAI21_X1 U6161 ( .B1(n5051), .B2(n5434), .A(n5036), .ZN(n5056) );
  NOR2_X1 U6162 ( .A1(n5885), .A2(n6539), .ZN(n5007) );
  INV_X1 U6163 ( .A(n5007), .ZN(n5004) );
  NAND2_X1 U6164 ( .A1(n5428), .A2(n5842), .ZN(n5571) );
  INV_X1 U6165 ( .A(n5377), .ZN(n5002) );
  NAND2_X1 U6166 ( .A1(n5386), .A2(n5002), .ZN(n5357) );
  NOR2_X1 U6167 ( .A1(n5357), .A2(n5358), .ZN(n5052) );
  NAND3_X1 U6168 ( .A1(n5052), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n4990), .ZN(n5003) );
  OAI211_X1 U6169 ( .C1(n5070), .C2(n5887), .A(n5004), .B(n5003), .ZN(n5005)
         );
  AOI21_X1 U6170 ( .B1(n5056), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5005), 
        .ZN(n5006) );
  OAI21_X1 U6171 ( .B1(n5012), .B2(n5846), .A(n5006), .ZN(U2988) );
  AOI21_X1 U6172 ( .B1(n5823), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5007), 
        .ZN(n5008) );
  OAI21_X1 U6173 ( .B1(n5840), .B2(n5064), .A(n5008), .ZN(n5009) );
  AOI21_X1 U6174 ( .B1(n5010), .B2(n5563), .A(n5009), .ZN(n5011) );
  OAI21_X1 U6175 ( .B1(n5012), .B2(n5817), .A(n5011), .ZN(U2956) );
  OAI211_X1 U6176 ( .C1(n5181), .C2(n5015), .A(n5078), .B(n5014), .ZN(n5016)
         );
  INV_X1 U6177 ( .A(n5016), .ZN(n5017) );
  OR2_X1 U6178 ( .A1(n5018), .A2(n5017), .ZN(n5028) );
  OAI222_X1 U6179 ( .A1(n5759), .A2(n5013), .B1(n5026), .B2(n5763), .C1(n5028), 
        .C2(n5758), .ZN(U2830) );
  AOI22_X1 U6180 ( .A1(n5770), .A2(DATAI_29_), .B1(n5773), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5022) );
  AND2_X1 U6181 ( .A1(n3176), .A2(n4501), .ZN(n5020) );
  NAND2_X1 U6182 ( .A1(n5774), .A2(DATAI_13_), .ZN(n5021) );
  OAI211_X1 U6183 ( .C1(n5013), .C2(n5534), .A(n5022), .B(n5021), .ZN(U2862)
         );
  NAND2_X1 U6184 ( .A1(n5743), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5025)
         );
  NAND2_X1 U6185 ( .A1(n5745), .A2(n5023), .ZN(n5024) );
  OAI211_X1 U6186 ( .C1(n5741), .C2(n5026), .A(n5025), .B(n5024), .ZN(n5027)
         );
  AOI21_X1 U6187 ( .B1(n5081), .B2(REIP_REG_29__SCAN_IN), .A(n5027), .ZN(n5031) );
  INV_X1 U6188 ( .A(n5028), .ZN(n5039) );
  AOI21_X1 U6189 ( .B1(n5039), .B2(n5698), .A(n5029), .ZN(n5030) );
  OAI211_X1 U6190 ( .C1(n5013), .C2(n5673), .A(n5031), .B(n5030), .ZN(U2798)
         );
  INV_X1 U6191 ( .A(n5032), .ZN(n5041) );
  INV_X1 U6192 ( .A(n5052), .ZN(n5034) );
  OAI21_X1 U6193 ( .B1(n5034), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5033), 
        .ZN(n5038) );
  NOR2_X1 U6194 ( .A1(n5036), .A2(n5035), .ZN(n5037) );
  AOI211_X1 U6195 ( .C1(n5908), .C2(n5039), .A(n5038), .B(n5037), .ZN(n5040)
         );
  OAI21_X1 U6196 ( .B1(n5041), .B2(n5846), .A(n5040), .ZN(U2989) );
  INV_X1 U6197 ( .A(n4425), .ZN(n5044) );
  AOI21_X1 U6198 ( .B1(n6323), .B2(n5044), .A(n6418), .ZN(n5049) );
  NOR3_X1 U6199 ( .A1(n6538), .A2(n5043), .A3(n5042), .ZN(n5046) );
  NOR3_X1 U6200 ( .A1(n6415), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n5044), 
        .ZN(n5045) );
  AOI211_X1 U6201 ( .C1(n5047), .C2(n5603), .A(n5046), .B(n5045), .ZN(n5048)
         );
  OAI22_X1 U6202 ( .A1(n5049), .A2(n3063), .B1(n5048), .B2(n6418), .ZN(U3459)
         );
  INV_X1 U6203 ( .A(n5050), .ZN(n5060) );
  NAND3_X1 U6204 ( .A1(n5052), .A2(n5051), .A3(n4981), .ZN(n5054) );
  NAND2_X1 U6205 ( .A1(n5054), .A2(n5053), .ZN(n5055) );
  OAI21_X1 U6206 ( .B1(n5060), .B2(n5846), .A(n5059), .ZN(U2987) );
  OAI22_X1 U6207 ( .A1(n5062), .A2(n5758), .B1(n5763), .B2(n5061), .ZN(U2828)
         );
  INV_X1 U6208 ( .A(n5063), .ZN(n5072) );
  OAI22_X1 U6209 ( .A1(n5065), .A2(n5678), .B1(n5717), .B2(n5064), .ZN(n5068)
         );
  NOR3_X1 U6210 ( .A1(n5066), .A2(REIP_REG_30__SCAN_IN), .A3(n6401), .ZN(n5067) );
  AOI211_X1 U6211 ( .C1(EBX_REG_30__SCAN_IN), .C2(n5746), .A(n5068), .B(n5067), 
        .ZN(n5069) );
  OAI21_X1 U6212 ( .B1(n5070), .B2(n5755), .A(n5069), .ZN(n5071) );
  AOI21_X1 U6213 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5072), .A(n5071), .ZN(n5073) );
  OAI21_X1 U6214 ( .B1(n5235), .B2(n5673), .A(n5073), .ZN(U2797) );
  AOI21_X1 U6215 ( .B1(n5075), .B2(n5074), .A(n4160), .ZN(n5259) );
  INV_X1 U6216 ( .A(n5259), .ZN(n5238) );
  OAI22_X1 U6217 ( .A1(n3810), .A2(n5678), .B1(n5717), .B2(n5257), .ZN(n5080)
         );
  NAND2_X1 U6218 ( .A1(n5092), .A2(n5076), .ZN(n5077) );
  NAND2_X1 U6219 ( .A1(n5078), .A2(n5077), .ZN(n5362) );
  NOR2_X1 U6220 ( .A1(n5362), .A2(n5755), .ZN(n5079) );
  AOI211_X1 U6221 ( .C1(EBX_REG_28__SCAN_IN), .C2(n5746), .A(n5080), .B(n5079), 
        .ZN(n5084) );
  INV_X1 U6222 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6396) );
  NOR2_X1 U6223 ( .A1(n5096), .A2(n6396), .ZN(n5082) );
  OAI21_X1 U6224 ( .B1(n5082), .B2(REIP_REG_28__SCAN_IN), .A(n5081), .ZN(n5083) );
  OAI211_X1 U6225 ( .C1(n5238), .C2(n5673), .A(n5084), .B(n5083), .ZN(U2799)
         );
  OAI21_X1 U6227 ( .B1(n5086), .B2(n5087), .A(n5074), .ZN(n5264) );
  INV_X1 U6228 ( .A(n5111), .ZN(n5098) );
  INV_X1 U6229 ( .A(n5088), .ZN(n5266) );
  OAI22_X1 U6230 ( .A1(n5089), .A2(n5678), .B1(n5717), .B2(n5266), .ZN(n5094)
         );
  NAND2_X1 U6231 ( .A1(n5105), .A2(n5090), .ZN(n5091) );
  NAND2_X1 U6232 ( .A1(n5092), .A2(n5091), .ZN(n5370) );
  NOR2_X1 U6233 ( .A1(n5370), .A2(n5755), .ZN(n5093) );
  AOI211_X1 U6234 ( .C1(n5746), .C2(EBX_REG_27__SCAN_IN), .A(n5094), .B(n5093), 
        .ZN(n5095) );
  OAI21_X1 U6235 ( .B1(REIP_REG_27__SCAN_IN), .B2(n5096), .A(n5095), .ZN(n5097) );
  AOI21_X1 U6236 ( .B1(REIP_REG_27__SCAN_IN), .B2(n5098), .A(n5097), .ZN(n5099) );
  OAI21_X1 U6237 ( .B1(n5264), .B2(n5673), .A(n5099), .ZN(U2800) );
  INV_X1 U6238 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6393) );
  NOR2_X1 U6239 ( .A1(n6393), .A2(n5480), .ZN(n5476) );
  AOI21_X1 U6240 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5476), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5110) );
  AOI21_X1 U6241 ( .B1(n5101), .B2(n2957), .A(n5086), .ZN(n5275) );
  NAND2_X1 U6242 ( .A1(n5275), .A2(n5692), .ZN(n5109) );
  OAI22_X1 U6243 ( .A1(n5102), .A2(n5678), .B1(n5717), .B2(n5273), .ZN(n5107)
         );
  OR2_X1 U6244 ( .A1(n5151), .A2(n5103), .ZN(n5104) );
  NAND2_X1 U6245 ( .A1(n5105), .A2(n5104), .ZN(n5380) );
  NOR2_X1 U6246 ( .A1(n5380), .A2(n5755), .ZN(n5106) );
  AOI211_X1 U6247 ( .C1(EBX_REG_26__SCAN_IN), .C2(n5746), .A(n5107), .B(n5106), 
        .ZN(n5108) );
  OAI211_X1 U6248 ( .C1(n5111), .C2(n5110), .A(n5109), .B(n5108), .ZN(U2801)
         );
  XNOR2_X1 U6250 ( .A(n5113), .B(n5168), .ZN(n5319) );
  INV_X1 U6251 ( .A(n5522), .ZN(n5510) );
  INV_X1 U6252 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6388) );
  AND2_X1 U6253 ( .A1(n6388), .A2(n5494), .ZN(n5509) );
  INV_X1 U6254 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5174) );
  OAI22_X1 U6255 ( .A1(n5741), .A2(n5174), .B1(n5314), .B2(n5678), .ZN(n5114)
         );
  AOI211_X1 U6256 ( .C1(n5510), .C2(REIP_REG_21__SCAN_IN), .A(n5509), .B(n5114), .ZN(n5119) );
  NAND2_X1 U6257 ( .A1(n5116), .A2(n5115), .ZN(n5117) );
  AND2_X1 U6258 ( .A1(n2988), .A2(n5117), .ZN(n5422) );
  AOI22_X1 U6259 ( .A1(n5698), .A2(n5422), .B1(n5745), .B2(n5316), .ZN(n5118)
         );
  OAI211_X1 U6260 ( .C1(n5319), .C2(n5673), .A(n5119), .B(n5118), .ZN(U2806)
         );
  BUF_X1 U6261 ( .A(n5120), .Z(n5121) );
  XOR2_X1 U6262 ( .A(n5122), .B(n5121), .Z(n5767) );
  INV_X1 U6263 ( .A(n5767), .ZN(n5132) );
  NOR2_X1 U6264 ( .A1(n5525), .A2(n5524), .ZN(n5629) );
  OAI21_X1 U6265 ( .B1(n5711), .B2(n5123), .A(n6381), .ZN(n5130) );
  INV_X1 U6266 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5202) );
  OAI22_X1 U6267 ( .A1(n5741), .A2(n5202), .B1(n5124), .B2(n5678), .ZN(n5129)
         );
  AND2_X1 U6268 ( .A1(n5125), .A2(n2993), .ZN(n5126) );
  OR2_X1 U6269 ( .A1(n5126), .A2(n5198), .ZN(n5566) );
  NAND2_X1 U6270 ( .A1(n5557), .A2(n5745), .ZN(n5127) );
  OAI211_X1 U6271 ( .C1(n5566), .C2(n5755), .A(n5127), .B(n5702), .ZN(n5128)
         );
  AOI211_X1 U6272 ( .C1(n5629), .C2(n5130), .A(n5129), .B(n5128), .ZN(n5131)
         );
  OAI21_X1 U6273 ( .B1(n5132), .B2(n5673), .A(n5131), .ZN(U2810) );
  AND2_X1 U6274 ( .A1(n5133), .A2(n5134), .ZN(n5136) );
  OR2_X1 U6275 ( .A1(n5136), .A2(n5135), .ZN(n5347) );
  OAI21_X1 U6276 ( .B1(n5711), .B2(n5139), .A(n5735), .ZN(n5646) );
  INV_X1 U6277 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5137) );
  OAI22_X1 U6278 ( .A1(n5717), .A2(n5343), .B1(n5741), .B2(n5137), .ZN(n5142)
         );
  AOI21_X1 U6279 ( .B1(n5138), .B2(n5223), .A(n5207), .ZN(n5584) );
  NOR2_X1 U6280 ( .A1(n5711), .A2(REIP_REG_15__SCAN_IN), .ZN(n5636) );
  AOI22_X1 U6281 ( .A1(n5698), .A2(n5584), .B1(n5139), .B2(n5636), .ZN(n5140)
         );
  OAI211_X1 U6282 ( .C1(n5678), .C2(n3565), .A(n5140), .B(n5702), .ZN(n5141)
         );
  AOI211_X1 U6283 ( .C1(REIP_REG_15__SCAN_IN), .C2(n5646), .A(n5142), .B(n5141), .ZN(n5143) );
  OAI21_X1 U6284 ( .B1(n5347), .B2(n5673), .A(n5143), .ZN(U2812) );
  OAI222_X1 U6285 ( .A1(n5759), .A2(n5238), .B1(n5144), .B2(n5763), .C1(n5362), 
        .C2(n5225), .ZN(U2831) );
  OAI222_X1 U6286 ( .A1(n5759), .A2(n5264), .B1(n5763), .B2(n4038), .C1(n5370), 
        .C2(n5225), .ZN(U2832) );
  INV_X1 U6287 ( .A(n5275), .ZN(n5243) );
  OAI222_X1 U6288 ( .A1(n5759), .A2(n5243), .B1(n5145), .B2(n5763), .C1(n5380), 
        .C2(n5225), .ZN(U2833) );
  OR2_X1 U6289 ( .A1(n5146), .A2(n5147), .ZN(n5148) );
  AND2_X1 U6290 ( .A1(n2957), .A2(n5148), .ZN(n5535) );
  AND2_X1 U6291 ( .A1(n5157), .A2(n5149), .ZN(n5150) );
  OR2_X1 U6292 ( .A1(n5151), .A2(n5150), .ZN(n5478) );
  INV_X1 U6293 ( .A(EBX_REG_25__SCAN_IN), .ZN(n6551) );
  OAI22_X1 U6294 ( .A1(n5478), .A2(n5225), .B1(n6551), .B2(n5763), .ZN(n5152)
         );
  AOI21_X1 U6295 ( .B1(n5535), .B2(n5211), .A(n5152), .ZN(n5153) );
  INV_X1 U6296 ( .A(n5153), .ZN(U2834) );
  NOR2_X1 U6297 ( .A1(n2981), .A2(n5154), .ZN(n5155) );
  OR2_X1 U6298 ( .A1(n5165), .A2(n5156), .ZN(n5158) );
  AND2_X1 U6299 ( .A1(n5158), .A2(n5157), .ZN(n5399) );
  INV_X1 U6300 ( .A(n5399), .ZN(n5486) );
  OAI222_X1 U6301 ( .A1(n5759), .A2(n5487), .B1(n5763), .B2(n4026), .C1(n5486), 
        .C2(n5225), .ZN(U2835) );
  AND2_X1 U6302 ( .A1(n5159), .A2(n5160), .ZN(n5161) );
  OR2_X1 U6303 ( .A1(n5161), .A2(n2981), .ZN(n5496) );
  INV_X1 U6304 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5166) );
  NOR2_X1 U6305 ( .A1(n5163), .A2(n5162), .ZN(n5164) );
  OR2_X1 U6306 ( .A1(n5165), .A2(n5164), .ZN(n5495) );
  OAI222_X1 U6307 ( .A1(n5759), .A2(n5496), .B1(n5763), .B2(n5166), .C1(n5495), 
        .C2(n5225), .ZN(U2836) );
  OAI21_X1 U6308 ( .B1(n5113), .B2(n5168), .A(n5167), .ZN(n5169) );
  NAND2_X1 U6309 ( .A1(n5169), .A2(n5159), .ZN(n5506) );
  INV_X1 U6310 ( .A(n5506), .ZN(n5538) );
  INV_X1 U6311 ( .A(n5170), .ZN(n5171) );
  XNOR2_X1 U6312 ( .A(n2988), .B(n5171), .ZN(n5414) );
  INV_X1 U6313 ( .A(n5414), .ZN(n5505) );
  OAI22_X1 U6314 ( .A1(n5758), .A2(n5505), .B1(n5503), .B2(n5763), .ZN(n5172)
         );
  AOI21_X1 U6315 ( .B1(n5538), .B2(n5211), .A(n5172), .ZN(n5173) );
  INV_X1 U6316 ( .A(n5173), .ZN(U2837) );
  INV_X1 U6317 ( .A(n5319), .ZN(n5541) );
  INV_X1 U6318 ( .A(n5422), .ZN(n5175) );
  OAI22_X1 U6319 ( .A1(n5225), .A2(n5175), .B1(n5174), .B2(n5763), .ZN(n5176)
         );
  AOI21_X1 U6320 ( .B1(n5541), .B2(n5211), .A(n5176), .ZN(n5177) );
  INV_X1 U6321 ( .A(n5177), .ZN(U2838) );
  OAI21_X1 U6322 ( .B1(n5178), .B2(n5179), .A(n5113), .ZN(n5517) );
  INV_X1 U6323 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5184) );
  MUX2_X1 U6324 ( .A(n5181), .B(n5189), .S(n5180), .Z(n5182) );
  XOR2_X1 U6325 ( .A(n5183), .B(n5182), .Z(n5518) );
  OAI222_X1 U6326 ( .A1(n5759), .A2(n5517), .B1(n5184), .B2(n5763), .C1(n5225), 
        .C2(n5518), .ZN(U2839) );
  AND2_X1 U6328 ( .A1(n5186), .A2(n5187), .ZN(n5188) );
  NOR2_X1 U6329 ( .A1(n5178), .A2(n5188), .ZN(n5547) );
  INV_X1 U6330 ( .A(n5547), .ZN(n5193) );
  NAND2_X1 U6331 ( .A1(n5189), .A2(n3969), .ZN(n5190) );
  OAI21_X1 U6332 ( .B1(n5191), .B2(n3969), .A(n5190), .ZN(n5199) );
  NAND2_X1 U6333 ( .A1(n5199), .A2(n5198), .ZN(n5197) );
  XOR2_X1 U6334 ( .A(n5192), .B(n5197), .Z(n5533) );
  OAI222_X1 U6335 ( .A1(n5193), .A2(n5759), .B1(n5763), .B2(n4007), .C1(n5758), 
        .C2(n5533), .ZN(U2840) );
  NAND2_X1 U6336 ( .A1(n5194), .A2(n5195), .ZN(n5196) );
  INV_X1 U6337 ( .A(n5764), .ZN(n5201) );
  INV_X1 U6338 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5200) );
  OAI21_X1 U6339 ( .B1(n5199), .B2(n5198), .A(n5197), .ZN(n5635) );
  OAI222_X1 U6340 ( .A1(n5201), .A2(n5759), .B1(n5200), .B2(n5763), .C1(n5758), 
        .C2(n5635), .ZN(U2841) );
  OAI22_X1 U6341 ( .A1(n5225), .A2(n5566), .B1(n5202), .B2(n5763), .ZN(n5203)
         );
  AOI21_X1 U6342 ( .B1(n5767), .B2(n5211), .A(n5203), .ZN(n5204) );
  INV_X1 U6343 ( .A(n5204), .ZN(U2842) );
  OR2_X1 U6344 ( .A1(n5135), .A2(n5205), .ZN(n5206) );
  AND2_X1 U6345 ( .A1(n5121), .A2(n5206), .ZN(n5772) );
  OR2_X1 U6346 ( .A1(n5208), .A2(n5207), .ZN(n5209) );
  NAND2_X1 U6347 ( .A1(n5209), .A2(n2993), .ZN(n5644) );
  OAI22_X1 U6348 ( .A1(n5225), .A2(n5644), .B1(n5763), .B2(n6556), .ZN(n5210)
         );
  AOI21_X1 U6349 ( .B1(n5772), .B2(n5211), .A(n5210), .ZN(n5212) );
  INV_X1 U6350 ( .A(n5212), .ZN(U2843) );
  INV_X1 U6351 ( .A(n5584), .ZN(n5213) );
  OAI22_X1 U6352 ( .A1(n5758), .A2(n5213), .B1(n5763), .B2(n5137), .ZN(n5214)
         );
  INV_X1 U6353 ( .A(n5214), .ZN(n5215) );
  OAI21_X1 U6354 ( .B1(n5347), .B2(n5759), .A(n5215), .ZN(U2844) );
  INV_X1 U6355 ( .A(n5216), .ZN(n5219) );
  INV_X1 U6356 ( .A(n5217), .ZN(n5218) );
  NAND2_X1 U6357 ( .A1(n5219), .A2(n5218), .ZN(n5220) );
  AND2_X1 U6358 ( .A1(n5220), .A2(n5133), .ZN(n5649) );
  INV_X1 U6359 ( .A(n5649), .ZN(n5252) );
  OR2_X1 U6360 ( .A1(n5222), .A2(n5221), .ZN(n5224) );
  AND2_X1 U6361 ( .A1(n5224), .A2(n5223), .ZN(n5647) );
  INV_X1 U6362 ( .A(n5647), .ZN(n5226) );
  OAI222_X1 U6363 ( .A1(n5252), .A2(n5759), .B1(n5227), .B2(n5763), .C1(n5226), 
        .C2(n5225), .ZN(U2845) );
  AND2_X1 U6364 ( .A1(n5248), .A2(n5228), .ZN(n5229) );
  NAND2_X1 U6365 ( .A1(n5230), .A2(n5229), .ZN(n5232) );
  AOI22_X1 U6366 ( .A1(n5770), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5773), .ZN(n5231) );
  NAND2_X1 U6367 ( .A1(n5232), .A2(n5231), .ZN(U2860) );
  AOI22_X1 U6368 ( .A1(n5770), .A2(DATAI_30_), .B1(n5773), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5234) );
  NAND2_X1 U6369 ( .A1(n5774), .A2(DATAI_14_), .ZN(n5233) );
  OAI211_X1 U6370 ( .C1(n5235), .C2(n5534), .A(n5234), .B(n5233), .ZN(U2861)
         );
  AOI22_X1 U6371 ( .A1(n5770), .A2(DATAI_28_), .B1(n5773), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U6372 ( .A1(n5774), .A2(DATAI_12_), .ZN(n5236) );
  OAI211_X1 U6373 ( .C1(n5238), .C2(n5534), .A(n5237), .B(n5236), .ZN(U2863)
         );
  AOI22_X1 U6374 ( .A1(n5770), .A2(DATAI_27_), .B1(n5773), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U6375 ( .A1(n5774), .A2(DATAI_11_), .ZN(n5239) );
  OAI211_X1 U6376 ( .C1(n5264), .C2(n5534), .A(n5240), .B(n5239), .ZN(U2864)
         );
  AOI22_X1 U6377 ( .A1(n5770), .A2(DATAI_26_), .B1(n5773), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5242) );
  NAND2_X1 U6378 ( .A1(n5774), .A2(DATAI_10_), .ZN(n5241) );
  OAI211_X1 U6379 ( .C1(n5243), .C2(n5534), .A(n5242), .B(n5241), .ZN(U2865)
         );
  AOI22_X1 U6380 ( .A1(n5770), .A2(DATAI_24_), .B1(n5773), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5245) );
  NAND2_X1 U6381 ( .A1(n5774), .A2(DATAI_8_), .ZN(n5244) );
  OAI211_X1 U6382 ( .C1(n5487), .C2(n5534), .A(n5245), .B(n5244), .ZN(U2867)
         );
  AOI22_X1 U6383 ( .A1(n5770), .A2(DATAI_23_), .B1(n5773), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5247) );
  NAND2_X1 U6384 ( .A1(n5774), .A2(DATAI_7_), .ZN(n5246) );
  OAI211_X1 U6385 ( .C1(n5496), .C2(n5534), .A(n5247), .B(n5246), .ZN(U2868)
         );
  INV_X1 U6386 ( .A(DATAI_15_), .ZN(n6566) );
  OAI222_X1 U6387 ( .A1(n5347), .A2(n5534), .B1(n5249), .B2(n6566), .C1(n5248), 
        .C2(n6574), .ZN(U2876) );
  AOI22_X1 U6388 ( .A1(n5250), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n5773), .ZN(n5251) );
  OAI21_X1 U6389 ( .B1(n5252), .B2(n5534), .A(n5251), .ZN(U2877) );
  NAND3_X1 U6390 ( .A1(n4151), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5298), .ZN(n5254) );
  NAND2_X1 U6391 ( .A1(n6476), .A2(n5385), .ZN(n5376) );
  NOR2_X1 U6392 ( .A1(n5808), .A2(n5376), .ZN(n5253) );
  NAND2_X1 U6393 ( .A1(n5279), .A2(n5253), .ZN(n5261) );
  AOI22_X1 U6394 ( .A1(n5254), .A2(n5261), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n6476), .ZN(n5255) );
  XNOR2_X1 U6395 ( .A(n5255), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5365)
         );
  INV_X1 U6396 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6399) );
  NOR2_X1 U6397 ( .A1(n5885), .A2(n6399), .ZN(n5356) );
  AOI21_X1 U6398 ( .B1(n5823), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5356), 
        .ZN(n5256) );
  OAI21_X1 U6399 ( .B1(n5840), .B2(n5257), .A(n5256), .ZN(n5258) );
  AOI21_X1 U6400 ( .B1(n5259), .B2(n5563), .A(n5258), .ZN(n5260) );
  OAI21_X1 U6401 ( .B1(n5817), .B2(n5365), .A(n5260), .ZN(U2958) );
  NAND2_X1 U6402 ( .A1(n5262), .A2(n5261), .ZN(n5263) );
  XNOR2_X1 U6403 ( .A(n5263), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5374)
         );
  INV_X1 U6404 ( .A(n5264), .ZN(n5268) );
  NOR2_X1 U6405 ( .A1(n5885), .A2(n6396), .ZN(n5366) );
  AOI21_X1 U6406 ( .B1(n5823), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5366), 
        .ZN(n5265) );
  OAI21_X1 U6407 ( .B1(n5840), .B2(n5266), .A(n5265), .ZN(n5267) );
  AOI21_X1 U6408 ( .B1(n5268), .B2(n5563), .A(n5267), .ZN(n5269) );
  OAI21_X1 U6409 ( .B1(n5374), .B2(n5817), .A(n5269), .ZN(U2959) );
  XNOR2_X1 U6410 ( .A(n5298), .B(n6476), .ZN(n5270) );
  XNOR2_X1 U6411 ( .A(n4149), .B(n5270), .ZN(n5383) );
  INV_X1 U6412 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5271) );
  NOR2_X1 U6413 ( .A1(n5885), .A2(n5271), .ZN(n5375) );
  AOI21_X1 U6414 ( .B1(n5823), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5375), 
        .ZN(n5272) );
  OAI21_X1 U6415 ( .B1(n5840), .B2(n5273), .A(n5272), .ZN(n5274) );
  AOI21_X1 U6416 ( .B1(n5275), .B2(n5563), .A(n5274), .ZN(n5276) );
  OAI21_X1 U6417 ( .B1(n5817), .B2(n5383), .A(n5276), .ZN(U2960) );
  OAI21_X1 U6418 ( .B1(n5279), .B2(n5278), .A(n5277), .ZN(n5280) );
  INV_X1 U6419 ( .A(n5280), .ZN(n5390) );
  INV_X1 U6420 ( .A(n5477), .ZN(n5283) );
  INV_X1 U6421 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5281) );
  NOR2_X1 U6422 ( .A1(n5885), .A2(n5281), .ZN(n5384) );
  AOI21_X1 U6423 ( .B1(n5823), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5384), 
        .ZN(n5282) );
  OAI21_X1 U6424 ( .B1(n5840), .B2(n5283), .A(n5282), .ZN(n5284) );
  AOI21_X1 U6425 ( .B1(n5535), .B2(n5563), .A(n5284), .ZN(n5285) );
  OAI21_X1 U6426 ( .B1(n5390), .B2(n5817), .A(n5285), .ZN(U2961) );
  OAI21_X1 U6427 ( .B1(n2966), .B2(n5442), .A(n5808), .ZN(n5288) );
  AND2_X2 U6428 ( .A1(n5286), .A2(n5288), .ZN(n5321) );
  XNOR2_X1 U6429 ( .A(n5298), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5320)
         );
  NOR2_X1 U6430 ( .A1(n5298), .A2(n5289), .ZN(n5290) );
  XNOR2_X1 U6431 ( .A(n5808), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5313)
         );
  NOR2_X1 U6432 ( .A1(n5808), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5305)
         );
  NAND2_X1 U6433 ( .A1(n5291), .A2(n5305), .ZN(n5299) );
  NAND3_X1 U6434 ( .A1(n5298), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5293) );
  XNOR2_X1 U6435 ( .A(n5294), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5401)
         );
  NAND2_X1 U6436 ( .A1(n5910), .A2(REIP_REG_24__SCAN_IN), .ZN(n5391) );
  OAI21_X1 U6437 ( .B1(n5323), .B2(n5492), .A(n5391), .ZN(n5296) );
  NOR2_X1 U6438 ( .A1(n5487), .A2(n6225), .ZN(n5295) );
  AOI211_X1 U6439 ( .C1(n5558), .C2(n5485), .A(n5296), .B(n5295), .ZN(n5297)
         );
  OAI21_X1 U6440 ( .B1(n5401), .B2(n5817), .A(n5297), .ZN(U2962) );
  NAND3_X1 U6441 ( .A1(n5298), .A2(n5410), .A3(n5435), .ZN(n5300) );
  OAI21_X1 U6442 ( .B1(n2966), .B2(n5300), .A(n5299), .ZN(n5301) );
  XNOR2_X1 U6443 ( .A(n5301), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5408)
         );
  NAND2_X1 U6444 ( .A1(n5910), .A2(REIP_REG_23__SCAN_IN), .ZN(n5402) );
  OAI21_X1 U6445 ( .B1(n5323), .B2(n5502), .A(n5402), .ZN(n5303) );
  NOR2_X1 U6446 ( .A1(n5496), .A2(n6225), .ZN(n5302) );
  AOI211_X1 U6447 ( .C1(n5558), .C2(n5493), .A(n5303), .B(n5302), .ZN(n5304)
         );
  OAI21_X1 U6448 ( .B1(n5408), .B2(n5817), .A(n5304), .ZN(U2963) );
  AOI21_X1 U6449 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5808), .A(n5305), 
        .ZN(n5307) );
  XOR2_X1 U6450 ( .A(n5307), .B(n5306), .Z(n5409) );
  NAND2_X1 U6451 ( .A1(n5409), .A2(n5835), .ZN(n5310) );
  AND2_X1 U6452 ( .A1(n5910), .A2(REIP_REG_22__SCAN_IN), .ZN(n5413) );
  NOR2_X1 U6453 ( .A1(n5840), .A2(n5513), .ZN(n5308) );
  AOI211_X1 U6454 ( .C1(n5823), .C2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5413), 
        .B(n5308), .ZN(n5309) );
  OAI211_X1 U6455 ( .C1(n6225), .C2(n5506), .A(n5310), .B(n5309), .ZN(U2964)
         );
  OAI21_X1 U6456 ( .B1(n5313), .B2(n5312), .A(n5311), .ZN(n5418) );
  NAND2_X1 U6457 ( .A1(n5418), .A2(n5835), .ZN(n5318) );
  NAND2_X1 U6458 ( .A1(n5910), .A2(REIP_REG_21__SCAN_IN), .ZN(n5419) );
  OAI21_X1 U6459 ( .B1(n5323), .B2(n5314), .A(n5419), .ZN(n5315) );
  AOI21_X1 U6460 ( .B1(n5558), .B2(n5316), .A(n5315), .ZN(n5317) );
  OAI211_X1 U6461 ( .C1(n6225), .C2(n5319), .A(n5318), .B(n5317), .ZN(U2965)
         );
  XNOR2_X1 U6462 ( .A(n5321), .B(n5320), .ZN(n5441) );
  NAND2_X1 U6463 ( .A1(n5910), .A2(REIP_REG_20__SCAN_IN), .ZN(n5438) );
  OAI21_X1 U6464 ( .B1(n5323), .B2(n5322), .A(n5438), .ZN(n5325) );
  NOR2_X1 U6465 ( .A1(n5517), .A2(n6225), .ZN(n5324) );
  AOI211_X1 U6466 ( .C1(n5558), .C2(n5514), .A(n5325), .B(n5324), .ZN(n5326)
         );
  OAI21_X1 U6467 ( .B1(n5817), .B2(n5441), .A(n5326), .ZN(U2966) );
  OAI21_X1 U6468 ( .B1(n5327), .B2(n5442), .A(n5286), .ZN(n5328) );
  XNOR2_X1 U6469 ( .A(n5328), .B(n4130), .ZN(n5449) );
  INV_X1 U6470 ( .A(n5528), .ZN(n5330) );
  NAND2_X1 U6471 ( .A1(n5910), .A2(REIP_REG_19__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U6472 ( .A1(n5823), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5329)
         );
  OAI211_X1 U6473 ( .C1(n5330), .C2(n5840), .A(n5445), .B(n5329), .ZN(n5331)
         );
  AOI21_X1 U6474 ( .B1(n5547), .B2(n5563), .A(n5331), .ZN(n5332) );
  OAI21_X1 U6475 ( .B1(n5449), .B2(n5817), .A(n5332), .ZN(U2967) );
  NAND2_X1 U6476 ( .A1(n5335), .A2(n5334), .ZN(n5336) );
  XNOR2_X1 U6477 ( .A(n2963), .B(n5336), .ZN(n5576) );
  INV_X1 U6478 ( .A(n5641), .ZN(n5338) );
  AOI22_X1 U6479 ( .A1(n5823), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n5910), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5337) );
  OAI21_X1 U6480 ( .B1(n5338), .B2(n5840), .A(n5337), .ZN(n5339) );
  AOI21_X1 U6481 ( .B1(n5772), .B2(n5563), .A(n5339), .ZN(n5340) );
  OAI21_X1 U6482 ( .B1(n5576), .B2(n5817), .A(n5340), .ZN(U2970) );
  XNOR2_X1 U6483 ( .A(n5298), .B(n5591), .ZN(n5342) );
  XNOR2_X1 U6484 ( .A(n2962), .B(n5342), .ZN(n5588) );
  NAND2_X1 U6485 ( .A1(n5588), .A2(n5835), .ZN(n5346) );
  AND2_X1 U6486 ( .A1(n5910), .A2(REIP_REG_15__SCAN_IN), .ZN(n5583) );
  NOR2_X1 U6487 ( .A1(n5840), .A2(n5343), .ZN(n5344) );
  AOI211_X1 U6488 ( .C1(n5823), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5583), 
        .B(n5344), .ZN(n5345) );
  OAI211_X1 U6489 ( .C1(n6225), .C2(n5347), .A(n5346), .B(n5345), .ZN(U2971)
         );
  XNOR2_X1 U6490 ( .A(n4130), .B(n5349), .ZN(n5350) );
  XNOR2_X1 U6491 ( .A(n2961), .B(n5350), .ZN(n5470) );
  NAND2_X1 U6492 ( .A1(n5910), .A2(REIP_REG_14__SCAN_IN), .ZN(n5465) );
  INV_X1 U6493 ( .A(n5465), .ZN(n5351) );
  AOI21_X1 U6494 ( .B1(n5823), .B2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5351), 
        .ZN(n5352) );
  OAI21_X1 U6495 ( .B1(n5840), .B2(n5353), .A(n5352), .ZN(n5354) );
  AOI21_X1 U6496 ( .B1(n5649), .B2(n5563), .A(n5354), .ZN(n5355) );
  OAI21_X1 U6497 ( .B1(n5470), .B2(n5817), .A(n5355), .ZN(U2972) );
  INV_X1 U6498 ( .A(n5356), .ZN(n5361) );
  INV_X1 U6499 ( .A(n5357), .ZN(n5368) );
  NAND3_X1 U6500 ( .A1(n5368), .A2(n5359), .A3(n5358), .ZN(n5360) );
  OAI211_X1 U6501 ( .C1(n5362), .C2(n5887), .A(n5361), .B(n5360), .ZN(n5363)
         );
  AOI21_X1 U6502 ( .B1(n5372), .B2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n5363), 
        .ZN(n5364) );
  OAI21_X1 U6503 ( .B1(n5365), .B2(n5846), .A(n5364), .ZN(U2990) );
  AOI21_X1 U6504 ( .B1(n5368), .B2(n5367), .A(n5366), .ZN(n5369) );
  OAI21_X1 U6505 ( .B1(n5370), .B2(n5887), .A(n5369), .ZN(n5371) );
  AOI21_X1 U6506 ( .B1(n5372), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5371), 
        .ZN(n5373) );
  OAI21_X1 U6507 ( .B1(n5374), .B2(n5846), .A(n5373), .ZN(U2991) );
  INV_X1 U6508 ( .A(n5375), .ZN(n5379) );
  NAND3_X1 U6509 ( .A1(n5386), .A2(n5377), .A3(n5376), .ZN(n5378) );
  OAI211_X1 U6510 ( .C1(n5380), .C2(n5887), .A(n5379), .B(n5378), .ZN(n5381)
         );
  AOI21_X1 U6511 ( .B1(n5393), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5381), 
        .ZN(n5382) );
  OAI21_X1 U6512 ( .B1(n5383), .B2(n5846), .A(n5382), .ZN(U2992) );
  AOI21_X1 U6513 ( .B1(n5386), .B2(n5385), .A(n5384), .ZN(n5387) );
  OAI21_X1 U6514 ( .B1(n5478), .B2(n5887), .A(n5387), .ZN(n5388) );
  AOI21_X1 U6515 ( .B1(n5393), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5388), 
        .ZN(n5389) );
  OAI21_X1 U6516 ( .B1(n5390), .B2(n5846), .A(n5389), .ZN(U2993) );
  INV_X1 U6517 ( .A(n5391), .ZN(n5398) );
  INV_X1 U6518 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5396) );
  NAND2_X1 U6519 ( .A1(n5443), .A2(n5435), .ZN(n5420) );
  OR2_X1 U6520 ( .A1(n5420), .A2(n5392), .ZN(n5403) );
  INV_X1 U6521 ( .A(n5393), .ZN(n5394) );
  AOI211_X1 U6522 ( .C1(n5396), .C2(n5403), .A(n5395), .B(n5394), .ZN(n5397)
         );
  AOI211_X1 U6523 ( .C1(n5908), .C2(n5399), .A(n5398), .B(n5397), .ZN(n5400)
         );
  OAI21_X1 U6524 ( .B1(n5401), .B2(n5846), .A(n5400), .ZN(U2994) );
  NOR2_X1 U6525 ( .A1(n5495), .A2(n5887), .ZN(n5405) );
  OAI21_X1 U6526 ( .B1(n5403), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5402), 
        .ZN(n5404) );
  AOI211_X1 U6527 ( .C1(n5406), .C2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5405), .B(n5404), .ZN(n5407) );
  OAI21_X1 U6528 ( .B1(n5408), .B2(n5846), .A(n5407), .ZN(U2995) );
  NAND2_X1 U6529 ( .A1(n5409), .A2(n5914), .ZN(n5416) );
  NOR3_X1 U6530 ( .A1(n5420), .A2(n5411), .A3(n5410), .ZN(n5412) );
  AOI211_X1 U6531 ( .C1(n5908), .C2(n5414), .A(n5413), .B(n5412), .ZN(n5415)
         );
  OAI211_X1 U6532 ( .C1(n5426), .C2(n5417), .A(n5416), .B(n5415), .ZN(U2996)
         );
  INV_X1 U6533 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5425) );
  NAND2_X1 U6534 ( .A1(n5418), .A2(n5914), .ZN(n5424) );
  OAI21_X1 U6535 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5420), .A(n5419), 
        .ZN(n5421) );
  AOI21_X1 U6536 ( .B1(n5908), .B2(n5422), .A(n5421), .ZN(n5423) );
  OAI211_X1 U6537 ( .C1(n5426), .C2(n5425), .A(n5424), .B(n5423), .ZN(U2997)
         );
  NAND2_X1 U6538 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5428), .ZN(n5452) );
  OAI221_X1 U6539 ( .B1(n5430), .B2(n5429), .C1(n5430), .C2(n5428), .A(n5427), 
        .ZN(n5431) );
  AOI21_X1 U6540 ( .B1(n5452), .B2(n5432), .A(n5431), .ZN(n5567) );
  OAI21_X1 U6541 ( .B1(n5434), .B2(n5433), .A(n5567), .ZN(n5447) );
  INV_X1 U6542 ( .A(n5435), .ZN(n5436) );
  OAI211_X1 U6543 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5443), .B(n5436), .ZN(n5437) );
  OAI211_X1 U6544 ( .C1(n5518), .C2(n5887), .A(n5438), .B(n5437), .ZN(n5439)
         );
  AOI21_X1 U6545 ( .B1(n5447), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5439), 
        .ZN(n5440) );
  OAI21_X1 U6546 ( .B1(n5441), .B2(n5846), .A(n5440), .ZN(U2998) );
  NAND2_X1 U6547 ( .A1(n5443), .A2(n5442), .ZN(n5444) );
  OAI211_X1 U6548 ( .C1(n5533), .C2(n5887), .A(n5445), .B(n5444), .ZN(n5446)
         );
  AOI21_X1 U6549 ( .B1(n5447), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5446), 
        .ZN(n5448) );
  OAI21_X1 U6550 ( .B1(n5449), .B2(n5846), .A(n5448), .ZN(U2999) );
  NOR3_X1 U6551 ( .A1(n2963), .A2(n5292), .A3(n5582), .ZN(n5553) );
  NAND3_X1 U6552 ( .A1(n2963), .A2(n5292), .A3(n5582), .ZN(n5554) );
  NOR2_X1 U6553 ( .A1(n5554), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5450)
         );
  AOI21_X1 U6554 ( .B1(n5553), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5450), 
        .ZN(n5451) );
  XNOR2_X1 U6555 ( .A(n5451), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5550)
         );
  INV_X1 U6556 ( .A(n5550), .ZN(n5458) );
  NOR2_X1 U6557 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5452), .ZN(n5456)
         );
  OAI21_X1 U6558 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5878), .A(n5567), 
        .ZN(n5453) );
  AOI22_X1 U6559 ( .A1(n5910), .A2(REIP_REG_18__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5453), .ZN(n5454) );
  OAI21_X1 U6560 ( .B1(n5887), .B2(n5635), .A(n5454), .ZN(n5455) );
  AOI21_X1 U6561 ( .B1(n5842), .B2(n5456), .A(n5455), .ZN(n5457) );
  OAI21_X1 U6562 ( .B1(n5458), .B2(n5846), .A(n5457), .ZN(U3000) );
  INV_X1 U6563 ( .A(n5459), .ZN(n5461) );
  NOR3_X1 U6564 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5460), .A3(n5593), 
        .ZN(n5598) );
  AOI211_X1 U6565 ( .C1(n5461), .C2(n5593), .A(n5598), .B(n5843), .ZN(n5462)
         );
  OAI21_X1 U6566 ( .B1(n5464), .B2(n5463), .A(n5462), .ZN(n5597) );
  NAND2_X1 U6567 ( .A1(n5464), .A2(n5842), .ZN(n5467) );
  NAND2_X1 U6568 ( .A1(n5908), .A2(n5647), .ZN(n5466) );
  OAI211_X1 U6569 ( .C1(n5467), .C2(INSTADDRPOINTER_REG_14__SCAN_IN), .A(n5466), .B(n5465), .ZN(n5468) );
  AOI21_X1 U6570 ( .B1(n5597), .B2(INSTADDRPOINTER_REG_14__SCAN_IN), .A(n5468), 
        .ZN(n5469) );
  OAI21_X1 U6571 ( .B1(n5470), .B2(n5846), .A(n5469), .ZN(U3004) );
  INV_X1 U6572 ( .A(n6067), .ZN(n5951) );
  OAI211_X1 U6573 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n4472), .A(n5951), .B(
        n6232), .ZN(n5471) );
  OAI21_X1 U6574 ( .B1(n5473), .B2(n4496), .A(n5471), .ZN(n5472) );
  MUX2_X1 U6575 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5472), .S(n5921), 
        .Z(U3464) );
  XNOR2_X1 U6576 ( .A(n4469), .B(n6067), .ZN(n5474) );
  OAI22_X1 U6577 ( .A1(n5474), .A2(n6221), .B1(n4447), .B2(n5473), .ZN(n5475)
         );
  MUX2_X1 U6578 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5475), .S(n5921), 
        .Z(U3463) );
  AND2_X1 U6579 ( .A1(n5795), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U6580 ( .A1(EBX_REG_25__SCAN_IN), .A2(n5746), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n5743), .ZN(n5484) );
  AOI22_X1 U6581 ( .A1(n5477), .A2(n5745), .B1(n5476), .B2(n5281), .ZN(n5483)
         );
  NOR2_X1 U6582 ( .A1(n5478), .A2(n5755), .ZN(n5479) );
  AOI21_X1 U6583 ( .B1(n5535), .B2(n5692), .A(n5479), .ZN(n5482) );
  NOR2_X1 U6584 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5480), .ZN(n5489) );
  OAI21_X1 U6585 ( .B1(n5489), .B2(n5499), .A(REIP_REG_25__SCAN_IN), .ZN(n5481) );
  NAND4_X1 U6586 ( .A1(n5484), .A2(n5483), .A3(n5482), .A4(n5481), .ZN(U2802)
         );
  AOI22_X1 U6587 ( .A1(EBX_REG_24__SCAN_IN), .A2(n5746), .B1(n5485), .B2(n5745), .ZN(n5491) );
  OAI22_X1 U6588 ( .A1(n5487), .A2(n5673), .B1(n5486), .B2(n5755), .ZN(n5488)
         );
  AOI211_X1 U6589 ( .C1(REIP_REG_24__SCAN_IN), .C2(n5499), .A(n5489), .B(n5488), .ZN(n5490) );
  OAI211_X1 U6590 ( .C1(n5492), .C2(n5678), .A(n5491), .B(n5490), .ZN(U2803)
         );
  AOI22_X1 U6591 ( .A1(EBX_REG_23__SCAN_IN), .A2(n5746), .B1(n5493), .B2(n5745), .ZN(n5501) );
  INV_X1 U6592 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6390) );
  NAND2_X1 U6593 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5494), .ZN(n5504) );
  INV_X1 U6594 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6392) );
  OAI21_X1 U6595 ( .B1(n6390), .B2(n5504), .A(n6392), .ZN(n5498) );
  OAI22_X1 U6596 ( .A1(n5496), .A2(n5673), .B1(n5495), .B2(n5755), .ZN(n5497)
         );
  AOI21_X1 U6597 ( .B1(n5499), .B2(n5498), .A(n5497), .ZN(n5500) );
  OAI211_X1 U6598 ( .C1(n5502), .C2(n5678), .A(n5501), .B(n5500), .ZN(U2804)
         );
  OAI22_X1 U6599 ( .A1(REIP_REG_22__SCAN_IN), .A2(n5504), .B1(n5741), .B2(
        n5503), .ZN(n5508) );
  OAI22_X1 U6600 ( .A1(n5506), .A2(n5673), .B1(n5505), .B2(n5755), .ZN(n5507)
         );
  AOI211_X1 U6601 ( .C1(PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n5743), .A(n5508), 
        .B(n5507), .ZN(n5512) );
  OAI21_X1 U6602 ( .B1(n5510), .B2(n5509), .A(REIP_REG_22__SCAN_IN), .ZN(n5511) );
  OAI211_X1 U6603 ( .C1(n5717), .C2(n5513), .A(n5512), .B(n5511), .ZN(U2805)
         );
  INV_X1 U6604 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6383) );
  NOR2_X1 U6605 ( .A1(n6383), .A2(n5627), .ZN(n5527) );
  AOI21_X1 U6606 ( .B1(REIP_REG_19__SCAN_IN), .B2(n5527), .A(
        REIP_REG_20__SCAN_IN), .ZN(n5523) );
  AOI22_X1 U6607 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n5743), .B1(n5514), 
        .B2(n5745), .ZN(n5515) );
  INV_X1 U6608 ( .A(n5515), .ZN(n5516) );
  AOI21_X1 U6609 ( .B1(EBX_REG_20__SCAN_IN), .B2(n5746), .A(n5516), .ZN(n5521)
         );
  INV_X1 U6610 ( .A(n5517), .ZN(n5544) );
  INV_X1 U6611 ( .A(n5518), .ZN(n5519) );
  AOI22_X1 U6612 ( .A1(n5544), .A2(n5692), .B1(n5698), .B2(n5519), .ZN(n5520)
         );
  OAI211_X1 U6613 ( .C1(n5523), .C2(n5522), .A(n5521), .B(n5520), .ZN(U2807)
         );
  OAI22_X1 U6614 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5627), .B1(n5525), .B2(
        n5524), .ZN(n5526) );
  AOI22_X1 U6615 ( .A1(EBX_REG_19__SCAN_IN), .A2(n5746), .B1(
        REIP_REG_19__SCAN_IN), .B2(n5526), .ZN(n5532) );
  INV_X1 U6616 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6386) );
  AOI22_X1 U6617 ( .A1(n5528), .A2(n5745), .B1(n5527), .B2(n6386), .ZN(n5529)
         );
  OAI211_X1 U6618 ( .C1(n3634), .C2(n5678), .A(n5529), .B(n5702), .ZN(n5530)
         );
  AOI21_X1 U6619 ( .B1(n5547), .B2(n5692), .A(n5530), .ZN(n5531) );
  OAI211_X1 U6620 ( .C1(n5533), .C2(n5755), .A(n5532), .B(n5531), .ZN(U2808)
         );
  AOI22_X1 U6621 ( .A1(n5535), .A2(n5771), .B1(n5770), .B2(DATAI_25_), .ZN(
        n5537) );
  AOI22_X1 U6622 ( .A1(n5774), .A2(DATAI_9_), .B1(n5773), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U6623 ( .A1(n5537), .A2(n5536), .ZN(U2866) );
  AOI22_X1 U6624 ( .A1(n5538), .A2(n5771), .B1(n5770), .B2(DATAI_22_), .ZN(
        n5540) );
  AOI22_X1 U6625 ( .A1(n5774), .A2(DATAI_6_), .B1(n5773), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5539) );
  NAND2_X1 U6626 ( .A1(n5540), .A2(n5539), .ZN(U2869) );
  AOI22_X1 U6627 ( .A1(n5541), .A2(n5771), .B1(n5770), .B2(DATAI_21_), .ZN(
        n5543) );
  AOI22_X1 U6628 ( .A1(n5774), .A2(DATAI_5_), .B1(n5773), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5542) );
  NAND2_X1 U6629 ( .A1(n5543), .A2(n5542), .ZN(U2870) );
  AOI22_X1 U6630 ( .A1(n5544), .A2(n5771), .B1(n5770), .B2(DATAI_20_), .ZN(
        n5546) );
  AOI22_X1 U6631 ( .A1(n5774), .A2(DATAI_4_), .B1(n5773), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U6632 ( .A1(n5546), .A2(n5545), .ZN(U2871) );
  AOI22_X1 U6633 ( .A1(n5547), .A2(n5771), .B1(n5770), .B2(DATAI_19_), .ZN(
        n5549) );
  AOI22_X1 U6634 ( .A1(n5774), .A2(DATAI_3_), .B1(n5773), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U6635 ( .A1(n5549), .A2(n5548), .ZN(U2872) );
  AOI22_X1 U6636 ( .A1(n5910), .A2(REIP_REG_18__SCAN_IN), .B1(n5823), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5552) );
  AOI22_X1 U6637 ( .A1(n5550), .A2(n5835), .B1(n5563), .B2(n5764), .ZN(n5551)
         );
  OAI211_X1 U6638 ( .C1(n5840), .C2(n5632), .A(n5552), .B(n5551), .ZN(U2968)
         );
  INV_X1 U6639 ( .A(n5553), .ZN(n5555) );
  NAND2_X1 U6640 ( .A1(n5555), .A2(n5554), .ZN(n5556) );
  XNOR2_X1 U6641 ( .A(n5556), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5575)
         );
  AOI22_X1 U6642 ( .A1(n5910), .A2(REIP_REG_17__SCAN_IN), .B1(n5823), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5560) );
  AOI22_X1 U6643 ( .A1(n5767), .A2(n5563), .B1(n5558), .B2(n5557), .ZN(n5559)
         );
  OAI211_X1 U6644 ( .C1(n5575), .C2(n5817), .A(n5560), .B(n5559), .ZN(U2969)
         );
  AOI22_X1 U6645 ( .A1(n5910), .A2(REIP_REG_13__SCAN_IN), .B1(n5823), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5565) );
  XNOR2_X1 U6646 ( .A(n5562), .B(n5561), .ZN(n5596) );
  AOI22_X1 U6647 ( .A1(n5596), .A2(n5835), .B1(n5563), .B2(n5659), .ZN(n5564)
         );
  OAI211_X1 U6648 ( .C1(n5840), .C2(n5662), .A(n5565), .B(n5564), .ZN(U2973)
         );
  INV_X1 U6649 ( .A(n5566), .ZN(n5573) );
  NAND2_X1 U6650 ( .A1(n5910), .A2(REIP_REG_17__SCAN_IN), .ZN(n5570) );
  INV_X1 U6651 ( .A(n5567), .ZN(n5568) );
  NAND2_X1 U6652 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5568), .ZN(n5569) );
  OAI211_X1 U6653 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5571), .A(n5570), .B(n5569), .ZN(n5572) );
  AOI21_X1 U6654 ( .B1(n5908), .B2(n5573), .A(n5572), .ZN(n5574) );
  OAI21_X1 U6655 ( .B1(n5575), .B2(n5846), .A(n5574), .ZN(U3001) );
  AOI21_X1 U6656 ( .B1(n5848), .B2(n5585), .A(n5843), .ZN(n5592) );
  AOI211_X1 U6657 ( .C1(n5591), .C2(n5582), .A(n5586), .B(n5585), .ZN(n5580)
         );
  INV_X1 U6658 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6379) );
  NOR2_X1 U6659 ( .A1(n5885), .A2(n6379), .ZN(n5578) );
  OAI22_X1 U6660 ( .A1(n5576), .A2(n5846), .B1(n5887), .B2(n5644), .ZN(n5577)
         );
  AOI211_X1 U6661 ( .C1(n5580), .C2(n5579), .A(n5578), .B(n5577), .ZN(n5581)
         );
  OAI21_X1 U6662 ( .B1(n5592), .B2(n5582), .A(n5581), .ZN(U3002) );
  AOI21_X1 U6663 ( .B1(n5908), .B2(n5584), .A(n5583), .ZN(n5590) );
  NOR2_X1 U6664 ( .A1(n5586), .A2(n5585), .ZN(n5587) );
  AOI22_X1 U6665 ( .A1(n5588), .A2(n5914), .B1(n5587), .B2(n5591), .ZN(n5589)
         );
  OAI211_X1 U6666 ( .C1(n5592), .C2(n5591), .A(n5590), .B(n5589), .ZN(U3003)
         );
  NOR2_X1 U6667 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5593), .ZN(n5594)
         );
  AOI22_X1 U6668 ( .A1(n5910), .A2(REIP_REG_13__SCAN_IN), .B1(n5595), .B2(
        n5594), .ZN(n5601) );
  AOI22_X1 U6669 ( .A1(n5596), .A2(n5914), .B1(n5908), .B2(n5653), .ZN(n5600)
         );
  OAI21_X1 U6670 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5598), .A(n5597), 
        .ZN(n5599) );
  NAND3_X1 U6671 ( .A1(n5601), .A2(n5600), .A3(n5599), .ZN(U3005) );
  NAND4_X1 U6672 ( .A1(n5709), .A2(n5604), .A3(n5603), .A4(n5602), .ZN(n5605)
         );
  OAI21_X1 U6673 ( .B1(n6423), .B2(n4460), .A(n5605), .ZN(U3455) );
  NOR2_X1 U6674 ( .A1(n6351), .A2(ADS_N_REG_SCAN_IN), .ZN(n5606) );
  NAND2_X1 U6675 ( .A1(STATE_REG_1__SCAN_IN), .A2(n3175), .ZN(n6349) );
  AOI21_X1 U6676 ( .B1(n5606), .B2(n6349), .A(n6449), .ZN(U2789) );
  INV_X1 U6677 ( .A(n6333), .ZN(n5610) );
  INV_X1 U6678 ( .A(n5607), .ZN(n5608) );
  INV_X1 U6679 ( .A(n6332), .ZN(n6330) );
  OAI21_X1 U6680 ( .B1(n5608), .B2(n6330), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5609) );
  OAI21_X1 U6681 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5610), .A(n5609), .ZN(
        U2790) );
  INV_X2 U6682 ( .A(n6449), .ZN(n6610) );
  NOR2_X1 U6683 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5612) );
  OAI21_X1 U6684 ( .B1(n5612), .B2(D_C_N_REG_SCAN_IN), .A(n6610), .ZN(n5611)
         );
  OAI21_X1 U6685 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6610), .A(n5611), .ZN(
        U2791) );
  AOI21_X1 U6686 ( .B1(STATE_REG_0__SCAN_IN), .B2(n6349), .A(n6449), .ZN(n6408) );
  OAI21_X1 U6687 ( .B1(n5612), .B2(BS16_N), .A(n6408), .ZN(n6407) );
  OAI21_X1 U6688 ( .B1(n6408), .B2(n6455), .A(n6407), .ZN(U2792) );
  OAI21_X1 U6689 ( .B1(n5614), .B2(n5613), .A(n5817), .ZN(U2793) );
  NOR4_X1 U6690 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_21__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n5618) );
  NOR4_X1 U6691 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_17__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n5617) );
  NOR4_X1 U6692 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5616) );
  NOR4_X1 U6693 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5615) );
  NAND4_X1 U6694 ( .A1(n5618), .A2(n5617), .A3(n5616), .A4(n5615), .ZN(n5624)
         );
  NOR4_X1 U6695 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), 
        .A3(DATAWIDTH_REG_4__SCAN_IN), .A4(DATAWIDTH_REG_5__SCAN_IN), .ZN(
        n5622) );
  AOI211_X1 U6696 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_16__SCAN_IN), .B(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n5621) );
  NOR4_X1 U6697 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_12__SCAN_IN), .A4(
        DATAWIDTH_REG_13__SCAN_IN), .ZN(n5620) );
  NOR4_X1 U6698 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_9__SCAN_IN), .ZN(
        n5619) );
  NAND4_X1 U6699 ( .A1(n5622), .A2(n5621), .A3(n5620), .A4(n5619), .ZN(n5623)
         );
  NOR2_X1 U6700 ( .A1(n5624), .A2(n5623), .ZN(n6431) );
  INV_X1 U6701 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6404) );
  INV_X1 U6702 ( .A(n6431), .ZN(n6435) );
  INV_X1 U6703 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6427) );
  INV_X1 U6704 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6428) );
  NAND4_X1 U6705 ( .A1(n6431), .A2(n6436), .A3(n6427), .A4(n6428), .ZN(n5625)
         );
  OAI221_X1 U6706 ( .B1(n6431), .B2(n6404), .C1(n6435), .C2(n6429), .A(n5625), 
        .ZN(U2794) );
  NOR2_X1 U6707 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6435), .ZN(n6437) );
  AOI22_X1 U6708 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(n6435), .B1(n6437), 
        .B2(n6427), .ZN(n5626) );
  NAND2_X1 U6709 ( .A1(n5626), .A2(n5625), .ZN(U2795) );
  NOR2_X1 U6710 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5627), .ZN(n5628) );
  AOI211_X1 U6711 ( .C1(n5743), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5628), 
        .B(n5708), .ZN(n5631) );
  AOI22_X1 U6712 ( .A1(EBX_REG_18__SCAN_IN), .A2(n5746), .B1(
        REIP_REG_18__SCAN_IN), .B2(n5629), .ZN(n5630) );
  OAI211_X1 U6713 ( .C1(n5632), .C2(n5717), .A(n5631), .B(n5630), .ZN(n5633)
         );
  AOI21_X1 U6714 ( .B1(n5764), .B2(n5692), .A(n5633), .ZN(n5634) );
  OAI21_X1 U6715 ( .B1(n5755), .B2(n5635), .A(n5634), .ZN(U2809) );
  OAI21_X1 U6716 ( .B1(n5646), .B2(n5636), .A(REIP_REG_16__SCAN_IN), .ZN(n5639) );
  NAND3_X1 U6717 ( .A1(n5734), .A2(n6379), .A3(n5637), .ZN(n5638) );
  OAI211_X1 U6718 ( .C1(n5741), .C2(n6556), .A(n5639), .B(n5638), .ZN(n5640)
         );
  AOI211_X1 U6719 ( .C1(n5743), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5708), 
        .B(n5640), .ZN(n5643) );
  AOI22_X1 U6720 ( .A1(n5772), .A2(n5692), .B1(n5745), .B2(n5641), .ZN(n5642)
         );
  OAI211_X1 U6721 ( .C1(n5755), .C2(n5644), .A(n5643), .B(n5642), .ZN(U2811)
         );
  NAND2_X1 U6722 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n5654) );
  INV_X1 U6723 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6377) );
  OAI21_X1 U6724 ( .B1(n5654), .B2(n5656), .A(n6377), .ZN(n5645) );
  AOI22_X1 U6725 ( .A1(EBX_REG_14__SCAN_IN), .A2(n5746), .B1(n5646), .B2(n5645), .ZN(n5652) );
  AOI22_X1 U6726 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n5743), .B1(n5698), 
        .B2(n5647), .ZN(n5651) );
  AOI22_X1 U6727 ( .A1(n5649), .A2(n5692), .B1(n5745), .B2(n5648), .ZN(n5650)
         );
  NAND4_X1 U6728 ( .A1(n5652), .A2(n5651), .A3(n5650), .A4(n5702), .ZN(U2813)
         );
  AOI22_X1 U6729 ( .A1(EBX_REG_13__SCAN_IN), .A2(n5746), .B1(n5698), .B2(n5653), .ZN(n5661) );
  OAI21_X1 U6730 ( .B1(REIP_REG_13__SCAN_IN), .B2(REIP_REG_12__SCAN_IN), .A(
        n5654), .ZN(n5657) );
  AOI22_X1 U6731 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n5743), .B1(
        REIP_REG_13__SCAN_IN), .B2(n5668), .ZN(n5655) );
  OAI211_X1 U6732 ( .C1(n5657), .C2(n5656), .A(n5655), .B(n5702), .ZN(n5658)
         );
  AOI21_X1 U6733 ( .B1(n5659), .B2(n5692), .A(n5658), .ZN(n5660) );
  OAI211_X1 U6734 ( .C1(n5662), .C2(n5717), .A(n5661), .B(n5660), .ZN(U2814)
         );
  INV_X1 U6735 ( .A(n5677), .ZN(n5664) );
  NOR3_X1 U6736 ( .A1(n5664), .A2(REIP_REG_11__SCAN_IN), .A3(n5663), .ZN(n5672) );
  AOI21_X1 U6737 ( .B1(n5667), .B2(n5666), .A(n5665), .ZN(n5841) );
  AOI22_X1 U6738 ( .A1(n5698), .A2(n5841), .B1(REIP_REG_11__SCAN_IN), .B2(
        n5668), .ZN(n5669) );
  OAI211_X1 U6739 ( .C1(n5678), .C2(n5670), .A(n5669), .B(n5702), .ZN(n5671)
         );
  AOI211_X1 U6740 ( .C1(EBX_REG_11__SCAN_IN), .C2(n5746), .A(n5672), .B(n5671), 
        .ZN(n5676) );
  OAI22_X1 U6741 ( .A1(n5812), .A2(n5673), .B1(n5717), .B2(n5811), .ZN(n5674)
         );
  INV_X1 U6742 ( .A(n5674), .ZN(n5675) );
  NAND2_X1 U6743 ( .A1(n5676), .A2(n5675), .ZN(U2816) );
  INV_X1 U6744 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6502) );
  AOI22_X1 U6745 ( .A1(EBX_REG_9__SCAN_IN), .A2(n5746), .B1(n5677), .B2(n6502), 
        .ZN(n5686) );
  OAI22_X1 U6746 ( .A1(n5679), .A2(n6502), .B1(n6568), .B2(n5678), .ZN(n5680)
         );
  AOI211_X1 U6747 ( .C1(n5698), .C2(n5858), .A(n5708), .B(n5680), .ZN(n5685)
         );
  INV_X1 U6748 ( .A(n5681), .ZN(n5683) );
  AOI22_X1 U6749 ( .A1(n5683), .A2(n5692), .B1(n5745), .B2(n5682), .ZN(n5684)
         );
  NAND3_X1 U6750 ( .A1(n5686), .A2(n5685), .A3(n5684), .ZN(U2818) );
  INV_X1 U6751 ( .A(n5816), .ZN(n5693) );
  AOI211_X1 U6752 ( .C1(n5743), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n5708), 
        .B(n5687), .ZN(n5689) );
  AOI22_X1 U6753 ( .A1(EBX_REG_6__SCAN_IN), .A2(n5746), .B1(
        REIP_REG_6__SCAN_IN), .B2(n5697), .ZN(n5688) );
  OAI211_X1 U6754 ( .C1(n5755), .C2(n5690), .A(n5689), .B(n5688), .ZN(n5691)
         );
  AOI21_X1 U6755 ( .B1(n5693), .B2(n5692), .A(n5691), .ZN(n5694) );
  OAI21_X1 U6756 ( .B1(n5822), .B2(n5717), .A(n5694), .ZN(U2821) );
  INV_X1 U6757 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6364) );
  NAND2_X1 U6758 ( .A1(n6364), .A2(n5695), .ZN(n5696) );
  AOI22_X1 U6759 ( .A1(EBX_REG_5__SCAN_IN), .A2(n5746), .B1(n5697), .B2(n5696), 
        .ZN(n5705) );
  AOI22_X1 U6760 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n5743), .B1(n5698), 
        .B2(n5875), .ZN(n5704) );
  INV_X1 U6761 ( .A(n5699), .ZN(n5701) );
  AOI22_X1 U6762 ( .A1(n5701), .A2(n5751), .B1(n5700), .B2(n5745), .ZN(n5703)
         );
  NAND4_X1 U6763 ( .A1(n5705), .A2(n5704), .A3(n5703), .A4(n5702), .ZN(U2822)
         );
  OAI22_X1 U6764 ( .A1(n5741), .A2(n5706), .B1(n5755), .B2(n5886), .ZN(n5707)
         );
  AOI211_X1 U6765 ( .C1(n5743), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5708), 
        .B(n5707), .ZN(n5716) );
  INV_X1 U6766 ( .A(n5735), .ZN(n5742) );
  OAI21_X1 U6767 ( .B1(n5742), .B2(n5710), .A(n5737), .ZN(n5728) );
  NAND2_X1 U6768 ( .A1(n5709), .A2(n5730), .ZN(n5713) );
  OR3_X1 U6769 ( .A1(n5711), .A2(n5710), .A3(REIP_REG_4__SCAN_IN), .ZN(n5712)
         );
  OAI211_X1 U6770 ( .C1(n6362), .C2(n5728), .A(n5713), .B(n5712), .ZN(n5714)
         );
  AOI21_X1 U6771 ( .B1(n5828), .B2(n5751), .A(n5714), .ZN(n5715) );
  OAI211_X1 U6772 ( .C1(n5831), .C2(n5717), .A(n5716), .B(n5715), .ZN(U2823)
         );
  INV_X1 U6773 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6360) );
  NAND2_X1 U6774 ( .A1(n5734), .A2(n6429), .ZN(n5747) );
  NAND3_X1 U6775 ( .A1(n5747), .A2(REIP_REG_2__SCAN_IN), .A3(n5735), .ZN(n5727) );
  AOI22_X1 U6776 ( .A1(n5746), .A2(EBX_REG_3__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n5743), .ZN(n5718) );
  OAI21_X1 U6777 ( .B1(n5755), .B2(n5719), .A(n5718), .ZN(n5720) );
  AOI21_X1 U6778 ( .B1(n5730), .B2(n2971), .A(n5720), .ZN(n5721) );
  OAI21_X1 U6779 ( .B1(n5723), .B2(n5722), .A(n5721), .ZN(n5724) );
  AOI21_X1 U6780 ( .B1(n5725), .B2(n5745), .A(n5724), .ZN(n5726) );
  OAI221_X1 U6781 ( .B1(n5728), .B2(n6360), .C1(n5728), .C2(n5727), .A(n5726), 
        .ZN(U2824) );
  INV_X1 U6782 ( .A(n5839), .ZN(n5729) );
  AOI22_X1 U6783 ( .A1(n5743), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n5745), 
        .B2(n5729), .ZN(n5732) );
  INV_X1 U6784 ( .A(n4447), .ZN(n5993) );
  NAND2_X1 U6785 ( .A1(n5993), .A2(n5730), .ZN(n5731) );
  OAI211_X1 U6786 ( .C1(n5905), .C2(n5755), .A(n5732), .B(n5731), .ZN(n5733)
         );
  AOI21_X1 U6787 ( .B1(n5836), .B2(n5751), .A(n5733), .ZN(n5740) );
  AND2_X1 U6788 ( .A1(n5734), .A2(REIP_REG_1__SCAN_IN), .ZN(n5738) );
  NAND3_X1 U6789 ( .A1(n5735), .A2(REIP_REG_1__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5736) );
  OAI211_X1 U6790 ( .C1(n5738), .C2(REIP_REG_2__SCAN_IN), .A(n5737), .B(n5736), 
        .ZN(n5739) );
  OAI211_X1 U6791 ( .C1(n5741), .C2(n3962), .A(n5740), .B(n5739), .ZN(U2825)
         );
  AOI22_X1 U6792 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n5743), .B1(n5742), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5754) );
  INV_X1 U6793 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5744) );
  AOI22_X1 U6794 ( .A1(n5746), .A2(EBX_REG_1__SCAN_IN), .B1(n5745), .B2(n5744), 
        .ZN(n5748) );
  OAI211_X1 U6795 ( .C1(n5749), .C2(n4496), .A(n5748), .B(n5747), .ZN(n5750)
         );
  AOI21_X1 U6796 ( .B1(n5752), .B2(n5751), .A(n5750), .ZN(n5753) );
  OAI211_X1 U6797 ( .C1(n5756), .C2(n5755), .A(n5754), .B(n5753), .ZN(U2826)
         );
  INV_X1 U6798 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5762) );
  INV_X1 U6799 ( .A(n5841), .ZN(n5757) );
  OAI22_X1 U6800 ( .A1(n5812), .A2(n5759), .B1(n5758), .B2(n5757), .ZN(n5760)
         );
  INV_X1 U6801 ( .A(n5760), .ZN(n5761) );
  OAI21_X1 U6802 ( .B1(n5763), .B2(n5762), .A(n5761), .ZN(U2848) );
  AOI22_X1 U6803 ( .A1(n5764), .A2(n5771), .B1(n5770), .B2(DATAI_18_), .ZN(
        n5766) );
  AOI22_X1 U6804 ( .A1(n5774), .A2(DATAI_2_), .B1(n5773), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U6805 ( .A1(n5766), .A2(n5765), .ZN(U2873) );
  AOI22_X1 U6806 ( .A1(n5767), .A2(n5771), .B1(n5770), .B2(DATAI_17_), .ZN(
        n5769) );
  AOI22_X1 U6807 ( .A1(n5774), .A2(DATAI_1_), .B1(n5773), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5768) );
  NAND2_X1 U6808 ( .A1(n5769), .A2(n5768), .ZN(U2874) );
  AOI22_X1 U6809 ( .A1(n5772), .A2(n5771), .B1(n5770), .B2(DATAI_16_), .ZN(
        n5776) );
  AOI22_X1 U6810 ( .A1(n5774), .A2(DATAI_0_), .B1(n5773), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5775) );
  NAND2_X1 U6811 ( .A1(n5776), .A2(n5775), .ZN(U2875) );
  AOI22_X1 U6812 ( .A1(n4387), .A2(LWORD_REG_15__SCAN_IN), .B1(n5795), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n5778) );
  OAI21_X1 U6813 ( .B1(n6574), .B2(n5805), .A(n5778), .ZN(U2908) );
  AOI22_X1 U6814 ( .A1(n4387), .A2(LWORD_REG_14__SCAN_IN), .B1(n5795), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n5779) );
  OAI21_X1 U6815 ( .B1(n6508), .B2(n5805), .A(n5779), .ZN(U2909) );
  AOI22_X1 U6816 ( .A1(n4387), .A2(LWORD_REG_13__SCAN_IN), .B1(n5795), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n5780) );
  OAI21_X1 U6817 ( .B1(n5781), .B2(n5805), .A(n5780), .ZN(U2910) );
  AOI22_X1 U6818 ( .A1(n4387), .A2(LWORD_REG_12__SCAN_IN), .B1(n5795), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n5782) );
  OAI21_X1 U6819 ( .B1(n5783), .B2(n5805), .A(n5782), .ZN(U2911) );
  AOI22_X1 U6820 ( .A1(n4387), .A2(LWORD_REG_11__SCAN_IN), .B1(n5795), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n5784) );
  OAI21_X1 U6821 ( .B1(n5785), .B2(n5805), .A(n5784), .ZN(U2912) );
  AOI22_X1 U6822 ( .A1(n4387), .A2(LWORD_REG_10__SCAN_IN), .B1(n5795), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n5786) );
  OAI21_X1 U6823 ( .B1(n5787), .B2(n5805), .A(n5786), .ZN(U2913) );
  AOI22_X1 U6824 ( .A1(n4387), .A2(LWORD_REG_9__SCAN_IN), .B1(n5795), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n5788) );
  OAI21_X1 U6825 ( .B1(n5789), .B2(n5805), .A(n5788), .ZN(U2914) );
  AOI22_X1 U6826 ( .A1(n4387), .A2(LWORD_REG_8__SCAN_IN), .B1(n5795), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n5790) );
  OAI21_X1 U6827 ( .B1(n6489), .B2(n5805), .A(n5790), .ZN(U2915) );
  AOI22_X1 U6828 ( .A1(n4387), .A2(LWORD_REG_7__SCAN_IN), .B1(n5795), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n5791) );
  OAI21_X1 U6829 ( .B1(n3450), .B2(n5805), .A(n5791), .ZN(U2916) );
  AOI22_X1 U6830 ( .A1(n4387), .A2(LWORD_REG_6__SCAN_IN), .B1(n5795), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5792) );
  OAI21_X1 U6831 ( .B1(n4551), .B2(n5805), .A(n5792), .ZN(U2917) );
  AOI22_X1 U6832 ( .A1(n4387), .A2(LWORD_REG_5__SCAN_IN), .B1(n5795), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n5793) );
  OAI21_X1 U6833 ( .B1(n5794), .B2(n5805), .A(n5793), .ZN(U2918) );
  AOI22_X1 U6834 ( .A1(n4387), .A2(LWORD_REG_4__SCAN_IN), .B1(n5795), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n5796) );
  OAI21_X1 U6835 ( .B1(n6496), .B2(n5805), .A(n5796), .ZN(U2919) );
  AOI22_X1 U6836 ( .A1(n4387), .A2(LWORD_REG_3__SCAN_IN), .B1(n5803), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n5797) );
  OAI21_X1 U6837 ( .B1(n5798), .B2(n5805), .A(n5797), .ZN(U2920) );
  AOI22_X1 U6838 ( .A1(n4387), .A2(LWORD_REG_2__SCAN_IN), .B1(n5803), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n5799) );
  OAI21_X1 U6839 ( .B1(n5800), .B2(n5805), .A(n5799), .ZN(U2921) );
  AOI22_X1 U6840 ( .A1(n4387), .A2(LWORD_REG_1__SCAN_IN), .B1(n5803), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n5801) );
  OAI21_X1 U6841 ( .B1(n5802), .B2(n5805), .A(n5801), .ZN(U2922) );
  AOI22_X1 U6842 ( .A1(n4387), .A2(LWORD_REG_0__SCAN_IN), .B1(n5803), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n5804) );
  OAI21_X1 U6843 ( .B1(n6554), .B2(n5805), .A(n5804), .ZN(U2923) );
  NAND2_X1 U6844 ( .A1(n5807), .A2(n5806), .ZN(n5810) );
  XNOR2_X1 U6845 ( .A(n5808), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5809)
         );
  XNOR2_X1 U6846 ( .A(n5810), .B(n5809), .ZN(n5847) );
  AOI22_X1 U6847 ( .A1(n5910), .A2(REIP_REG_11__SCAN_IN), .B1(n5823), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5815) );
  OAI22_X1 U6848 ( .A1(n5812), .A2(n6225), .B1(n5840), .B2(n5811), .ZN(n5813)
         );
  INV_X1 U6849 ( .A(n5813), .ZN(n5814) );
  OAI211_X1 U6850 ( .C1(n5847), .C2(n5817), .A(n5815), .B(n5814), .ZN(U2975)
         );
  AOI22_X1 U6851 ( .A1(n5910), .A2(REIP_REG_6__SCAN_IN), .B1(n5823), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5821) );
  OAI22_X1 U6852 ( .A1(n5818), .A2(n5817), .B1(n5816), .B2(n6225), .ZN(n5819)
         );
  INV_X1 U6853 ( .A(n5819), .ZN(n5820) );
  OAI211_X1 U6854 ( .C1(n5840), .C2(n5822), .A(n5821), .B(n5820), .ZN(U2980)
         );
  AOI22_X1 U6855 ( .A1(n5910), .A2(REIP_REG_4__SCAN_IN), .B1(n5823), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5830) );
  OAI21_X1 U6856 ( .B1(n5826), .B2(n5825), .A(n2958), .ZN(n5827) );
  INV_X1 U6857 ( .A(n5827), .ZN(n5889) );
  AOI22_X1 U6858 ( .A1(n5835), .A2(n5889), .B1(n5828), .B2(n5563), .ZN(n5829)
         );
  OAI211_X1 U6859 ( .C1(n5840), .C2(n5831), .A(n5830), .B(n5829), .ZN(U2982)
         );
  AOI22_X1 U6860 ( .A1(n5910), .A2(REIP_REG_2__SCAN_IN), .B1(n5823), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5838) );
  XOR2_X1 U6861 ( .A(n5832), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n5834) );
  XNOR2_X1 U6862 ( .A(n5834), .B(n5833), .ZN(n5915) );
  AOI22_X1 U6863 ( .A1(n5836), .A2(n5563), .B1(n5915), .B2(n5835), .ZN(n5837)
         );
  OAI211_X1 U6864 ( .C1(n5840), .C2(n5839), .A(n5838), .B(n5837), .ZN(U2984)
         );
  AOI22_X1 U6865 ( .A1(n5908), .A2(n5841), .B1(n5910), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n5845) );
  AOI22_X1 U6866 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n5843), .B1(n5842), .B2(n4131), .ZN(n5844) );
  OAI211_X1 U6867 ( .C1(n5847), .C2(n5846), .A(n5845), .B(n5844), .ZN(U3007)
         );
  NAND2_X1 U6868 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5853) );
  AOI21_X1 U6869 ( .B1(n5853), .B2(n5848), .A(n5865), .ZN(n5863) );
  OAI22_X1 U6870 ( .A1(n5887), .A2(n5849), .B1(n6371), .B2(n5885), .ZN(n5850)
         );
  AOI21_X1 U6871 ( .B1(n5851), .B2(n5914), .A(n5850), .ZN(n5855) );
  NOR2_X1 U6872 ( .A1(n5853), .A2(n5852), .ZN(n5859) );
  OAI221_X1 U6873 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n6461), .C2(n4129), .A(n5859), 
        .ZN(n5854) );
  OAI211_X1 U6874 ( .C1(n5863), .C2(n4129), .A(n5855), .B(n5854), .ZN(U3008)
         );
  INV_X1 U6875 ( .A(n5856), .ZN(n5857) );
  AOI21_X1 U6876 ( .B1(n5908), .B2(n5858), .A(n5857), .ZN(n5862) );
  AOI22_X1 U6877 ( .A1(n5860), .A2(n5914), .B1(n5859), .B2(n6461), .ZN(n5861)
         );
  OAI211_X1 U6878 ( .C1(n5863), .C2(n6461), .A(n5862), .B(n5861), .ZN(U3009)
         );
  INV_X1 U6879 ( .A(n5864), .ZN(n5866) );
  AOI22_X1 U6880 ( .A1(n5866), .A2(n5914), .B1(INSTADDRPOINTER_REG_7__SCAN_IN), 
        .B2(n5865), .ZN(n5871) );
  NOR2_X1 U6881 ( .A1(n5885), .A2(n6369), .ZN(n5868) );
  AOI211_X1 U6882 ( .C1(n5869), .C2(n5908), .A(n5868), .B(n5867), .ZN(n5870)
         );
  NAND2_X1 U6883 ( .A1(n5871), .A2(n5870), .ZN(U3011) );
  AOI21_X1 U6884 ( .B1(n5912), .B2(n5872), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n5883) );
  INV_X1 U6885 ( .A(n5873), .ZN(n5874) );
  AOI21_X1 U6886 ( .B1(n5908), .B2(n5875), .A(n5874), .ZN(n5882) );
  INV_X1 U6887 ( .A(n5876), .ZN(n5880) );
  NOR3_X1 U6888 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n5878), .A3(n5877), 
        .ZN(n5879) );
  AOI21_X1 U6889 ( .B1(n5880), .B2(n5914), .A(n5879), .ZN(n5881) );
  OAI211_X1 U6890 ( .C1(n5884), .C2(n5883), .A(n5882), .B(n5881), .ZN(U3013)
         );
  AOI21_X1 U6891 ( .B1(n5912), .B2(n5911), .A(n5913), .ZN(n5904) );
  OAI22_X1 U6892 ( .A1(n5887), .A2(n5886), .B1(n6362), .B2(n5885), .ZN(n5888)
         );
  AOI21_X1 U6893 ( .B1(n5889), .B2(n5914), .A(n5888), .ZN(n5893) );
  NOR2_X1 U6894 ( .A1(n5911), .A2(n5890), .ZN(n5900) );
  OAI211_X1 U6895 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n5900), .B(n5891), .ZN(n5892) );
  OAI211_X1 U6896 ( .C1(n5904), .C2(n5894), .A(n5893), .B(n5892), .ZN(U3014)
         );
  INV_X1 U6897 ( .A(n5895), .ZN(n5896) );
  AOI21_X1 U6898 ( .B1(n5908), .B2(n5897), .A(n5896), .ZN(n5902) );
  INV_X1 U6899 ( .A(n5898), .ZN(n5899) );
  AOI22_X1 U6900 ( .A1(n5900), .A2(n5903), .B1(n5899), .B2(n5914), .ZN(n5901)
         );
  OAI211_X1 U6901 ( .C1(n5904), .C2(n5903), .A(n5902), .B(n5901), .ZN(U3015)
         );
  INV_X1 U6902 ( .A(n5905), .ZN(n5909) );
  AOI22_X1 U6903 ( .A1(n5909), .A2(n5908), .B1(n5907), .B2(n5906), .ZN(n5920)
         );
  AOI22_X1 U6904 ( .A1(n5912), .A2(n5911), .B1(n5910), .B2(REIP_REG_2__SCAN_IN), .ZN(n5919) );
  AOI22_X1 U6905 ( .A1(n5915), .A2(n5914), .B1(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n5913), .ZN(n5918) );
  NAND3_X1 U6906 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4073), .A3(n5916), 
        .ZN(n5917) );
  NAND4_X1 U6907 ( .A1(n5920), .A2(n5919), .A3(n5918), .A4(n5917), .ZN(U3016)
         );
  NOR2_X1 U6908 ( .A1(n6311), .A2(n5921), .ZN(U3019) );
  NOR2_X1 U6909 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5922), .ZN(n5946)
         );
  OAI22_X1 U6910 ( .A1(n5927), .A2(n6221), .B1(n6105), .B2(n5923), .ZN(n5945)
         );
  AOI22_X1 U6911 ( .A1(n6223), .A2(n5946), .B1(n6222), .B2(n5945), .ZN(n5932)
         );
  INV_X1 U6912 ( .A(n5946), .ZN(n5925) );
  AOI211_X1 U6913 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5925), .A(n6187), .B(
        n5924), .ZN(n5930) );
  INV_X1 U6914 ( .A(n6283), .ZN(n5926) );
  OAI21_X1 U6915 ( .B1(n5947), .B2(n5926), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5928) );
  NAND3_X1 U6916 ( .A1(n5928), .A2(n6232), .A3(n5927), .ZN(n5929) );
  NAND2_X1 U6917 ( .A1(n5930), .A2(n5929), .ZN(n5948) );
  AOI22_X1 U6918 ( .A1(n5948), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n6145), 
        .B2(n5947), .ZN(n5931) );
  OAI211_X1 U6919 ( .C1(n6111), .C2(n6283), .A(n5932), .B(n5931), .ZN(U3020)
         );
  AOI22_X1 U6920 ( .A1(n6239), .A2(n5946), .B1(n6238), .B2(n5945), .ZN(n5934)
         );
  AOI22_X1 U6921 ( .A1(n5948), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n6153), 
        .B2(n5947), .ZN(n5933) );
  OAI211_X1 U6922 ( .C1(n6114), .C2(n6283), .A(n5934), .B(n5933), .ZN(U3021)
         );
  AOI22_X1 U6923 ( .A1(n6245), .A2(n5945), .B1(n6244), .B2(n5946), .ZN(n5936)
         );
  AOI22_X1 U6924 ( .A1(n5948), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n6157), 
        .B2(n5947), .ZN(n5935) );
  OAI211_X1 U6925 ( .C1(n6117), .C2(n6283), .A(n5936), .B(n5935), .ZN(U3022)
         );
  AOI22_X1 U6926 ( .A1(n6251), .A2(n5946), .B1(n6250), .B2(n5945), .ZN(n5938)
         );
  AOI22_X1 U6927 ( .A1(n5948), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n6161), 
        .B2(n5947), .ZN(n5937) );
  OAI211_X1 U6928 ( .C1(n6120), .C2(n6283), .A(n5938), .B(n5937), .ZN(U3023)
         );
  AOI22_X1 U6929 ( .A1(n6257), .A2(n5945), .B1(n6256), .B2(n5946), .ZN(n5940)
         );
  AOI22_X1 U6930 ( .A1(n5948), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n6165), 
        .B2(n5947), .ZN(n5939) );
  OAI211_X1 U6931 ( .C1(n6123), .C2(n6283), .A(n5940), .B(n5939), .ZN(U3024)
         );
  AOI22_X1 U6932 ( .A1(n6263), .A2(n5945), .B1(n6262), .B2(n5946), .ZN(n5942)
         );
  AOI22_X1 U6933 ( .A1(n5948), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n6169), 
        .B2(n5947), .ZN(n5941) );
  OAI211_X1 U6934 ( .C1(n6126), .C2(n6283), .A(n5942), .B(n5941), .ZN(U3025)
         );
  AOI22_X1 U6935 ( .A1(n6269), .A2(n5945), .B1(n6268), .B2(n5946), .ZN(n5944)
         );
  AOI22_X1 U6936 ( .A1(n5948), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n6173), 
        .B2(n5947), .ZN(n5943) );
  OAI211_X1 U6937 ( .C1(n6129), .C2(n6283), .A(n5944), .B(n5943), .ZN(U3026)
         );
  AOI22_X1 U6938 ( .A1(n6277), .A2(n5946), .B1(n6275), .B2(n5945), .ZN(n5950)
         );
  AOI22_X1 U6939 ( .A1(n5948), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n6178), 
        .B2(n5947), .ZN(n5949) );
  OAI211_X1 U6940 ( .C1(n6136), .C2(n6283), .A(n5950), .B(n5949), .ZN(U3027)
         );
  NOR2_X1 U6941 ( .A1(n6066), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5976)
         );
  AOI22_X1 U6942 ( .A1(n6234), .A2(n5965), .B1(n6223), .B2(n5976), .ZN(n5962)
         );
  INV_X1 U6943 ( .A(n5958), .ZN(n5956) );
  OAI21_X1 U6944 ( .B1(n4469), .B2(n5951), .A(n6232), .ZN(n5952) );
  NAND2_X1 U6945 ( .A1(n5953), .A2(n5952), .ZN(n5957) );
  AOI21_X1 U6946 ( .B1(n5954), .B2(n6296), .A(n5976), .ZN(n5959) );
  NAND2_X1 U6947 ( .A1(n5957), .A2(n5959), .ZN(n5955) );
  OAI211_X1 U6948 ( .C1(n6232), .C2(n5956), .A(n5955), .B(n6231), .ZN(n5979)
         );
  INV_X1 U6949 ( .A(n5957), .ZN(n5960) );
  OAI22_X1 U6950 ( .A1(n5960), .A2(n5959), .B1(n5958), .B2(n6442), .ZN(n5978)
         );
  AOI22_X1 U6951 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n5979), .B1(n6222), 
        .B2(n5978), .ZN(n5961) );
  OAI211_X1 U6952 ( .C1(n6237), .C2(n5990), .A(n5962), .B(n5961), .ZN(U3044)
         );
  AOI22_X1 U6953 ( .A1(n6153), .A2(n5977), .B1(n6239), .B2(n5976), .ZN(n5964)
         );
  AOI22_X1 U6954 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n5979), .B1(n6238), 
        .B2(n5978), .ZN(n5963) );
  OAI211_X1 U6955 ( .C1(n5982), .C2(n6114), .A(n5964), .B(n5963), .ZN(U3045)
         );
  AOI22_X1 U6956 ( .A1(n6246), .A2(n5965), .B1(n6244), .B2(n5976), .ZN(n5967)
         );
  AOI22_X1 U6957 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n5979), .B1(n6245), 
        .B2(n5978), .ZN(n5966) );
  OAI211_X1 U6958 ( .C1(n6249), .C2(n5990), .A(n5967), .B(n5966), .ZN(U3046)
         );
  AOI22_X1 U6959 ( .A1(n6161), .A2(n5977), .B1(n6251), .B2(n5976), .ZN(n5969)
         );
  AOI22_X1 U6960 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n5979), .B1(n6250), 
        .B2(n5978), .ZN(n5968) );
  OAI211_X1 U6961 ( .C1(n5982), .C2(n6120), .A(n5969), .B(n5968), .ZN(U3047)
         );
  AOI22_X1 U6962 ( .A1(n6165), .A2(n5977), .B1(n6256), .B2(n5976), .ZN(n5971)
         );
  AOI22_X1 U6963 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n5979), .B1(n6257), 
        .B2(n5978), .ZN(n5970) );
  OAI211_X1 U6964 ( .C1(n5982), .C2(n6123), .A(n5971), .B(n5970), .ZN(U3048)
         );
  AOI22_X1 U6965 ( .A1(n6169), .A2(n5977), .B1(n6262), .B2(n5976), .ZN(n5973)
         );
  AOI22_X1 U6966 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n5979), .B1(n6263), 
        .B2(n5978), .ZN(n5972) );
  OAI211_X1 U6967 ( .C1(n5982), .C2(n6126), .A(n5973), .B(n5972), .ZN(U3049)
         );
  AOI22_X1 U6968 ( .A1(n6173), .A2(n5977), .B1(n6268), .B2(n5976), .ZN(n5975)
         );
  AOI22_X1 U6969 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n5979), .B1(n6269), 
        .B2(n5978), .ZN(n5974) );
  OAI211_X1 U6970 ( .C1(n5982), .C2(n6129), .A(n5975), .B(n5974), .ZN(U3050)
         );
  AOI22_X1 U6971 ( .A1(n6178), .A2(n5977), .B1(n6277), .B2(n5976), .ZN(n5981)
         );
  AOI22_X1 U6972 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n5979), .B1(n6275), 
        .B2(n5978), .ZN(n5980) );
  OAI211_X1 U6973 ( .C1(n5982), .C2(n6136), .A(n5981), .B(n5980), .ZN(U3051)
         );
  INV_X1 U6974 ( .A(n5983), .ZN(n5985) );
  AOI22_X1 U6975 ( .A1(n6269), .A2(n5985), .B1(n6268), .B2(n5984), .ZN(n5989)
         );
  AOI22_X1 U6976 ( .A1(n5987), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n6173), 
        .B2(n5986), .ZN(n5988) );
  OAI211_X1 U6977 ( .C1(n6129), .C2(n5990), .A(n5989), .B(n5988), .ZN(U3058)
         );
  NOR2_X1 U6978 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6031), .ZN(n6018)
         );
  NAND2_X1 U6979 ( .A1(n5993), .A2(n5992), .ZN(n6192) );
  NAND2_X1 U6980 ( .A1(n6219), .A2(n6232), .ZN(n6190) );
  NAND3_X1 U6981 ( .A1(n6187), .A2(n6186), .A3(n6313), .ZN(n5994) );
  OAI21_X1 U6982 ( .B1(n6190), .B2(n2971), .A(n5994), .ZN(n6017) );
  AOI22_X1 U6983 ( .A1(n6223), .A2(n6018), .B1(n6222), .B2(n6017), .ZN(n6004)
         );
  AOI21_X1 U6984 ( .B1(n6002), .B2(n6053), .A(n6455), .ZN(n6001) );
  NAND2_X1 U6985 ( .A1(n6219), .A2(n5995), .ZN(n6027) );
  NAND2_X1 U6986 ( .A1(n6027), .A2(n6232), .ZN(n6000) );
  NOR2_X1 U6987 ( .A1(n5997), .A2(n5996), .ZN(n6195) );
  INV_X1 U6988 ( .A(n6018), .ZN(n5998) );
  AOI21_X1 U6989 ( .B1(n5998), .B2(STATE2_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5999) );
  OAI211_X1 U6990 ( .C1(n6001), .C2(n6000), .A(n6195), .B(n5999), .ZN(n6020)
         );
  AOI22_X1 U6991 ( .A1(n6020), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6234), 
        .B2(n6019), .ZN(n6003) );
  OAI211_X1 U6992 ( .C1(n6237), .C2(n6053), .A(n6004), .B(n6003), .ZN(U3068)
         );
  AOI22_X1 U6993 ( .A1(n6239), .A2(n6018), .B1(n6238), .B2(n6017), .ZN(n6006)
         );
  AOI22_X1 U6994 ( .A1(n6020), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6240), 
        .B2(n6019), .ZN(n6005) );
  OAI211_X1 U6995 ( .C1(n6243), .C2(n6053), .A(n6006), .B(n6005), .ZN(U3069)
         );
  AOI22_X1 U6996 ( .A1(n6245), .A2(n6017), .B1(n6244), .B2(n6018), .ZN(n6008)
         );
  AOI22_X1 U6997 ( .A1(n6020), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6246), 
        .B2(n6019), .ZN(n6007) );
  OAI211_X1 U6998 ( .C1(n6249), .C2(n6053), .A(n6008), .B(n6007), .ZN(U3070)
         );
  AOI22_X1 U6999 ( .A1(n6251), .A2(n6018), .B1(n6250), .B2(n6017), .ZN(n6010)
         );
  AOI22_X1 U7000 ( .A1(n6020), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6252), 
        .B2(n6019), .ZN(n6009) );
  OAI211_X1 U7001 ( .C1(n6255), .C2(n6053), .A(n6010), .B(n6009), .ZN(U3071)
         );
  AOI22_X1 U7002 ( .A1(n6257), .A2(n6017), .B1(n6256), .B2(n6018), .ZN(n6012)
         );
  AOI22_X1 U7003 ( .A1(n6020), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6258), 
        .B2(n6019), .ZN(n6011) );
  OAI211_X1 U7004 ( .C1(n6261), .C2(n6053), .A(n6012), .B(n6011), .ZN(U3072)
         );
  AOI22_X1 U7005 ( .A1(n6263), .A2(n6017), .B1(n6262), .B2(n6018), .ZN(n6014)
         );
  AOI22_X1 U7006 ( .A1(n6020), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6264), 
        .B2(n6019), .ZN(n6013) );
  OAI211_X1 U7007 ( .C1(n6267), .C2(n6053), .A(n6014), .B(n6013), .ZN(U3073)
         );
  AOI22_X1 U7008 ( .A1(n6269), .A2(n6017), .B1(n6268), .B2(n6018), .ZN(n6016)
         );
  AOI22_X1 U7009 ( .A1(n6020), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6270), 
        .B2(n6019), .ZN(n6015) );
  OAI211_X1 U7010 ( .C1(n6273), .C2(n6053), .A(n6016), .B(n6015), .ZN(U3074)
         );
  AOI22_X1 U7011 ( .A1(n6277), .A2(n6018), .B1(n6275), .B2(n6017), .ZN(n6022)
         );
  AOI22_X1 U7012 ( .A1(n6020), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6279), 
        .B2(n6019), .ZN(n6021) );
  OAI211_X1 U7013 ( .C1(n6284), .C2(n6053), .A(n6022), .B(n6021), .ZN(U3075)
         );
  INV_X1 U7014 ( .A(n6026), .ZN(n6048) );
  AOI22_X1 U7015 ( .A1(n6223), .A2(n6048), .B1(n6047), .B2(n6145), .ZN(n6033)
         );
  INV_X1 U7016 ( .A(n6029), .ZN(n6023) );
  NAND2_X1 U7017 ( .A1(n6232), .A2(n6023), .ZN(n6024) );
  NAND2_X1 U7018 ( .A1(n6024), .A2(n6031), .ZN(n6025) );
  NAND2_X1 U7019 ( .A1(n6231), .A2(n6025), .ZN(n6050) );
  OAI21_X1 U7020 ( .B1(n6027), .B2(n3342), .A(n6026), .ZN(n6028) );
  NAND3_X1 U7021 ( .A1(n6029), .A2(n6232), .A3(n6028), .ZN(n6030) );
  OAI21_X1 U7022 ( .B1(n6031), .B2(n6442), .A(n6030), .ZN(n6049) );
  AOI22_X1 U7023 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6050), .B1(n6222), 
        .B2(n6049), .ZN(n6032) );
  OAI211_X1 U7024 ( .C1(n6111), .C2(n6053), .A(n6033), .B(n6032), .ZN(U3076)
         );
  AOI22_X1 U7025 ( .A1(n6239), .A2(n6048), .B1(n6047), .B2(n6153), .ZN(n6035)
         );
  AOI22_X1 U7026 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6050), .B1(n6238), 
        .B2(n6049), .ZN(n6034) );
  OAI211_X1 U7027 ( .C1(n6114), .C2(n6053), .A(n6035), .B(n6034), .ZN(U3077)
         );
  AOI22_X1 U7028 ( .A1(n6244), .A2(n6048), .B1(n6047), .B2(n6157), .ZN(n6037)
         );
  AOI22_X1 U7029 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6050), .B1(n6245), 
        .B2(n6049), .ZN(n6036) );
  OAI211_X1 U7030 ( .C1(n6117), .C2(n6053), .A(n6037), .B(n6036), .ZN(U3078)
         );
  INV_X1 U7031 ( .A(n6053), .ZN(n6042) );
  AOI22_X1 U7032 ( .A1(n6251), .A2(n6048), .B1(n6042), .B2(n6252), .ZN(n6039)
         );
  AOI22_X1 U7033 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6050), .B1(n6250), 
        .B2(n6049), .ZN(n6038) );
  OAI211_X1 U7034 ( .C1(n6255), .C2(n6063), .A(n6039), .B(n6038), .ZN(U3079)
         );
  AOI22_X1 U7035 ( .A1(n6256), .A2(n6048), .B1(n6047), .B2(n6165), .ZN(n6041)
         );
  AOI22_X1 U7036 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6050), .B1(n6257), 
        .B2(n6049), .ZN(n6040) );
  OAI211_X1 U7037 ( .C1(n6123), .C2(n6053), .A(n6041), .B(n6040), .ZN(U3080)
         );
  AOI22_X1 U7038 ( .A1(n6262), .A2(n6048), .B1(n6042), .B2(n6264), .ZN(n6044)
         );
  AOI22_X1 U7039 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6050), .B1(n6263), 
        .B2(n6049), .ZN(n6043) );
  OAI211_X1 U7040 ( .C1(n6267), .C2(n6063), .A(n6044), .B(n6043), .ZN(U3081)
         );
  AOI22_X1 U7041 ( .A1(n6268), .A2(n6048), .B1(n6047), .B2(n6173), .ZN(n6046)
         );
  AOI22_X1 U7042 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6050), .B1(n6269), 
        .B2(n6049), .ZN(n6045) );
  OAI211_X1 U7043 ( .C1(n6129), .C2(n6053), .A(n6046), .B(n6045), .ZN(U3082)
         );
  AOI22_X1 U7044 ( .A1(n6277), .A2(n6048), .B1(n6047), .B2(n6178), .ZN(n6052)
         );
  AOI22_X1 U7045 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6050), .B1(n6275), 
        .B2(n6049), .ZN(n6051) );
  OAI211_X1 U7046 ( .C1(n6136), .C2(n6053), .A(n6052), .B(n6051), .ZN(U3083)
         );
  INV_X1 U7047 ( .A(n6054), .ZN(n6057) );
  AOI22_X1 U7048 ( .A1(n6269), .A2(n6057), .B1(n6268), .B2(n6058), .ZN(n6056)
         );
  AOI22_X1 U7049 ( .A1(n6060), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6173), 
        .B2(n6059), .ZN(n6055) );
  OAI211_X1 U7050 ( .C1(n6129), .C2(n6063), .A(n6056), .B(n6055), .ZN(U3090)
         );
  AOI22_X1 U7051 ( .A1(n6277), .A2(n6058), .B1(n6275), .B2(n6057), .ZN(n6062)
         );
  AOI22_X1 U7052 ( .A1(n6060), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6178), 
        .B2(n6059), .ZN(n6061) );
  OAI211_X1 U7053 ( .C1(n6136), .C2(n6063), .A(n6062), .B(n6061), .ZN(U3091)
         );
  NOR2_X1 U7054 ( .A1(n6066), .A2(n6313), .ZN(n6090) );
  AOI22_X1 U7055 ( .A1(n6087), .A2(n6234), .B1(n6223), .B2(n6090), .ZN(n6076)
         );
  AOI21_X1 U7056 ( .B1(n6068), .B2(n6067), .A(n6221), .ZN(n6071) );
  AOI21_X1 U7057 ( .B1(n6069), .B2(n6296), .A(n6090), .ZN(n6073) );
  AOI22_X1 U7058 ( .A1(n6071), .A2(n6073), .B1(n6072), .B2(n6221), .ZN(n6070)
         );
  NAND2_X1 U7059 ( .A1(n6231), .A2(n6070), .ZN(n6093) );
  INV_X1 U7060 ( .A(n6071), .ZN(n6074) );
  OAI22_X1 U7061 ( .A1(n6074), .A2(n6073), .B1(n6072), .B2(n6442), .ZN(n6092)
         );
  AOI22_X1 U7062 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6093), .B1(n6222), 
        .B2(n6092), .ZN(n6075) );
  OAI211_X1 U7063 ( .C1(n6237), .C2(n6135), .A(n6076), .B(n6075), .ZN(U3108)
         );
  AOI22_X1 U7064 ( .A1(n6087), .A2(n6240), .B1(n6239), .B2(n6090), .ZN(n6078)
         );
  AOI22_X1 U7065 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6093), .B1(n6238), 
        .B2(n6092), .ZN(n6077) );
  OAI211_X1 U7066 ( .C1(n6243), .C2(n6135), .A(n6078), .B(n6077), .ZN(U3109)
         );
  AOI22_X1 U7067 ( .A1(n6087), .A2(n6246), .B1(n6244), .B2(n6090), .ZN(n6080)
         );
  AOI22_X1 U7068 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6093), .B1(n6245), 
        .B2(n6092), .ZN(n6079) );
  OAI211_X1 U7069 ( .C1(n6249), .C2(n6135), .A(n6080), .B(n6079), .ZN(U3110)
         );
  INV_X1 U7070 ( .A(n6135), .ZN(n6091) );
  AOI22_X1 U7071 ( .A1(n6161), .A2(n6091), .B1(n6251), .B2(n6090), .ZN(n6082)
         );
  AOI22_X1 U7072 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6093), .B1(n6250), 
        .B2(n6092), .ZN(n6081) );
  OAI211_X1 U7073 ( .C1(n6120), .C2(n6096), .A(n6082), .B(n6081), .ZN(U3111)
         );
  AOI22_X1 U7074 ( .A1(n6087), .A2(n6258), .B1(n6256), .B2(n6090), .ZN(n6084)
         );
  AOI22_X1 U7075 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6093), .B1(n6257), 
        .B2(n6092), .ZN(n6083) );
  OAI211_X1 U7076 ( .C1(n6261), .C2(n6135), .A(n6084), .B(n6083), .ZN(U3112)
         );
  AOI22_X1 U7077 ( .A1(n6169), .A2(n6091), .B1(n6262), .B2(n6090), .ZN(n6086)
         );
  AOI22_X1 U7078 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6093), .B1(n6263), 
        .B2(n6092), .ZN(n6085) );
  OAI211_X1 U7079 ( .C1(n6126), .C2(n6096), .A(n6086), .B(n6085), .ZN(U3113)
         );
  AOI22_X1 U7080 ( .A1(n6087), .A2(n6270), .B1(n6268), .B2(n6090), .ZN(n6089)
         );
  AOI22_X1 U7081 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6093), .B1(n6269), 
        .B2(n6092), .ZN(n6088) );
  OAI211_X1 U7082 ( .C1(n6273), .C2(n6135), .A(n6089), .B(n6088), .ZN(U3114)
         );
  AOI22_X1 U7083 ( .A1(n6178), .A2(n6091), .B1(n6277), .B2(n6090), .ZN(n6095)
         );
  AOI22_X1 U7084 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6093), .B1(n6275), 
        .B2(n6092), .ZN(n6094) );
  OAI211_X1 U7085 ( .C1(n6136), .C2(n6096), .A(n6095), .B(n6094), .ZN(U3115)
         );
  NAND2_X1 U7086 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6142), .ZN(n6146) );
  NOR2_X1 U7087 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6146), .ZN(n6131)
         );
  INV_X1 U7088 ( .A(n6097), .ZN(n6100) );
  OAI22_X1 U7089 ( .A1(n6100), .A2(n6189), .B1(n6099), .B2(n6098), .ZN(n6130)
         );
  AOI22_X1 U7090 ( .A1(n6223), .A2(n6131), .B1(n6222), .B2(n6130), .ZN(n6110)
         );
  AOI21_X1 U7091 ( .B1(n6108), .B2(n6135), .A(n6455), .ZN(n6102) );
  AOI211_X1 U7092 ( .C1(n6139), .C2(n6103), .A(n6221), .B(n6102), .ZN(n6107)
         );
  OAI211_X1 U7093 ( .C1(n6413), .C2(n6131), .A(n6105), .B(n6104), .ZN(n6106)
         );
  AOI22_X1 U7094 ( .A1(n6132), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n6145), 
        .B2(n6179), .ZN(n6109) );
  OAI211_X1 U7095 ( .C1(n6111), .C2(n6135), .A(n6110), .B(n6109), .ZN(U3116)
         );
  AOI22_X1 U7096 ( .A1(n6239), .A2(n6131), .B1(n6238), .B2(n6130), .ZN(n6113)
         );
  AOI22_X1 U7097 ( .A1(n6132), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n6153), 
        .B2(n6179), .ZN(n6112) );
  OAI211_X1 U7098 ( .C1(n6114), .C2(n6135), .A(n6113), .B(n6112), .ZN(U3117)
         );
  AOI22_X1 U7099 ( .A1(n6245), .A2(n6130), .B1(n6244), .B2(n6131), .ZN(n6116)
         );
  AOI22_X1 U7100 ( .A1(n6132), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n6157), 
        .B2(n6179), .ZN(n6115) );
  OAI211_X1 U7101 ( .C1(n6117), .C2(n6135), .A(n6116), .B(n6115), .ZN(U3118)
         );
  AOI22_X1 U7102 ( .A1(n6251), .A2(n6131), .B1(n6250), .B2(n6130), .ZN(n6119)
         );
  AOI22_X1 U7103 ( .A1(n6132), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n6161), 
        .B2(n6179), .ZN(n6118) );
  OAI211_X1 U7104 ( .C1(n6120), .C2(n6135), .A(n6119), .B(n6118), .ZN(U3119)
         );
  AOI22_X1 U7105 ( .A1(n6257), .A2(n6130), .B1(n6256), .B2(n6131), .ZN(n6122)
         );
  AOI22_X1 U7106 ( .A1(n6132), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n6165), 
        .B2(n6179), .ZN(n6121) );
  OAI211_X1 U7107 ( .C1(n6123), .C2(n6135), .A(n6122), .B(n6121), .ZN(U3120)
         );
  AOI22_X1 U7108 ( .A1(n6263), .A2(n6130), .B1(n6262), .B2(n6131), .ZN(n6125)
         );
  AOI22_X1 U7109 ( .A1(n6132), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n6169), 
        .B2(n6179), .ZN(n6124) );
  OAI211_X1 U7110 ( .C1(n6126), .C2(n6135), .A(n6125), .B(n6124), .ZN(U3121)
         );
  AOI22_X1 U7111 ( .A1(n6269), .A2(n6130), .B1(n6268), .B2(n6131), .ZN(n6128)
         );
  AOI22_X1 U7112 ( .A1(n6132), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n6173), 
        .B2(n6179), .ZN(n6127) );
  OAI211_X1 U7113 ( .C1(n6129), .C2(n6135), .A(n6128), .B(n6127), .ZN(U3122)
         );
  AOI22_X1 U7114 ( .A1(n6277), .A2(n6131), .B1(n6275), .B2(n6130), .ZN(n6134)
         );
  AOI22_X1 U7115 ( .A1(n6132), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n6178), 
        .B2(n6179), .ZN(n6133) );
  OAI211_X1 U7116 ( .C1(n6136), .C2(n6135), .A(n6134), .B(n6133), .ZN(U3123)
         );
  NOR2_X1 U7117 ( .A1(n6442), .A2(n6313), .ZN(n6141) );
  NOR2_X1 U7118 ( .A1(n6137), .A2(n6221), .ZN(n6147) );
  NOR2_X1 U7119 ( .A1(n6138), .A2(n6146), .ZN(n6177) );
  AOI21_X1 U7120 ( .B1(n6218), .B2(n6139), .A(n6177), .ZN(n6148) );
  INV_X1 U7121 ( .A(n6148), .ZN(n6140) );
  AOI22_X1 U7122 ( .A1(n6142), .A2(n6141), .B1(n6147), .B2(n6140), .ZN(n6184)
         );
  AOI22_X1 U7123 ( .A1(n6145), .A2(n2985), .B1(n6223), .B2(n6177), .ZN(n6151)
         );
  AOI22_X1 U7124 ( .A1(n6148), .A2(n6147), .B1(n6221), .B2(n6146), .ZN(n6149)
         );
  NAND2_X1 U7125 ( .A1(n6231), .A2(n6149), .ZN(n6180) );
  AOI22_X1 U7126 ( .A1(n6180), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n6234), 
        .B2(n6179), .ZN(n6150) );
  OAI211_X1 U7127 ( .C1(n6184), .C2(n6152), .A(n6151), .B(n6150), .ZN(U3124)
         );
  AOI22_X1 U7128 ( .A1(n6153), .A2(n2985), .B1(n6239), .B2(n6177), .ZN(n6155)
         );
  AOI22_X1 U7129 ( .A1(n6180), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n6240), 
        .B2(n6179), .ZN(n6154) );
  OAI211_X1 U7130 ( .C1(n6184), .C2(n6156), .A(n6155), .B(n6154), .ZN(U3125)
         );
  AOI22_X1 U7131 ( .A1(n6157), .A2(n2985), .B1(n6244), .B2(n6177), .ZN(n6159)
         );
  AOI22_X1 U7132 ( .A1(n6180), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n6246), 
        .B2(n6179), .ZN(n6158) );
  OAI211_X1 U7133 ( .C1(n6184), .C2(n6160), .A(n6159), .B(n6158), .ZN(U3126)
         );
  AOI22_X1 U7134 ( .A1(n6161), .A2(n2985), .B1(n6251), .B2(n6177), .ZN(n6163)
         );
  AOI22_X1 U7135 ( .A1(n6180), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n6252), 
        .B2(n6179), .ZN(n6162) );
  OAI211_X1 U7136 ( .C1(n6184), .C2(n6164), .A(n6163), .B(n6162), .ZN(U3127)
         );
  AOI22_X1 U7137 ( .A1(n6258), .A2(n6179), .B1(n6256), .B2(n6177), .ZN(n6167)
         );
  AOI22_X1 U7138 ( .A1(n6180), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n6165), 
        .B2(n2985), .ZN(n6166) );
  OAI211_X1 U7139 ( .C1(n6184), .C2(n6168), .A(n6167), .B(n6166), .ZN(U3128)
         );
  AOI22_X1 U7140 ( .A1(n6264), .A2(n6179), .B1(n6262), .B2(n6177), .ZN(n6171)
         );
  AOI22_X1 U7141 ( .A1(n6180), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n6169), 
        .B2(n2985), .ZN(n6170) );
  OAI211_X1 U7142 ( .C1(n6184), .C2(n6172), .A(n6171), .B(n6170), .ZN(U3129)
         );
  AOI22_X1 U7143 ( .A1(n6173), .A2(n2985), .B1(n6268), .B2(n6177), .ZN(n6175)
         );
  AOI22_X1 U7144 ( .A1(n6180), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n6270), 
        .B2(n6179), .ZN(n6174) );
  OAI211_X1 U7145 ( .C1(n6184), .C2(n6176), .A(n6175), .B(n6174), .ZN(U3130)
         );
  AOI22_X1 U7146 ( .A1(n6178), .A2(n2985), .B1(n6277), .B2(n6177), .ZN(n6182)
         );
  AOI22_X1 U7147 ( .A1(n6180), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n6279), 
        .B2(n6179), .ZN(n6181) );
  OAI211_X1 U7148 ( .C1(n6184), .C2(n6183), .A(n6182), .B(n6181), .ZN(U3131)
         );
  NOR2_X1 U7149 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6220), .ZN(n6212)
         );
  NAND3_X1 U7150 ( .A1(n6187), .A2(n6186), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6188) );
  OAI21_X1 U7151 ( .B1(n6190), .B2(n6189), .A(n6188), .ZN(n6211) );
  AOI22_X1 U7152 ( .A1(n6223), .A2(n6212), .B1(n6222), .B2(n6211), .ZN(n6198)
         );
  OAI21_X1 U7153 ( .B1(n2985), .B2(n6278), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6191) );
  NAND3_X1 U7154 ( .A1(n6192), .A2(n6232), .A3(n6191), .ZN(n6196) );
  OAI21_X1 U7155 ( .B1(n6413), .B2(n6212), .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .ZN(n6193) );
  INV_X1 U7156 ( .A(n6193), .ZN(n6194) );
  NAND3_X1 U7157 ( .A1(n6196), .A2(n6195), .A3(n6194), .ZN(n6213) );
  AOI22_X1 U7158 ( .A1(n6213), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n6234), 
        .B2(n2985), .ZN(n6197) );
  OAI211_X1 U7159 ( .C1(n6237), .C2(n6216), .A(n6198), .B(n6197), .ZN(U3132)
         );
  AOI22_X1 U7160 ( .A1(n6239), .A2(n6212), .B1(n6238), .B2(n6211), .ZN(n6200)
         );
  AOI22_X1 U7161 ( .A1(n6213), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n6240), 
        .B2(n2985), .ZN(n6199) );
  OAI211_X1 U7162 ( .C1(n6243), .C2(n6216), .A(n6200), .B(n6199), .ZN(U3133)
         );
  AOI22_X1 U7163 ( .A1(n6245), .A2(n6211), .B1(n6244), .B2(n6212), .ZN(n6202)
         );
  AOI22_X1 U7164 ( .A1(n6213), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n6246), 
        .B2(n2985), .ZN(n6201) );
  OAI211_X1 U7165 ( .C1(n6249), .C2(n6216), .A(n6202), .B(n6201), .ZN(U3134)
         );
  AOI22_X1 U7166 ( .A1(n6251), .A2(n6212), .B1(n6250), .B2(n6211), .ZN(n6204)
         );
  AOI22_X1 U7167 ( .A1(n6213), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n6252), 
        .B2(n2985), .ZN(n6203) );
  OAI211_X1 U7168 ( .C1(n6255), .C2(n6216), .A(n6204), .B(n6203), .ZN(U3135)
         );
  AOI22_X1 U7169 ( .A1(n6257), .A2(n6211), .B1(n6256), .B2(n6212), .ZN(n6206)
         );
  AOI22_X1 U7170 ( .A1(n6213), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n6258), 
        .B2(n2985), .ZN(n6205) );
  OAI211_X1 U7171 ( .C1(n6261), .C2(n6216), .A(n6206), .B(n6205), .ZN(U3136)
         );
  AOI22_X1 U7172 ( .A1(n6263), .A2(n6211), .B1(n6262), .B2(n6212), .ZN(n6208)
         );
  AOI22_X1 U7173 ( .A1(n6213), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n6264), 
        .B2(n2985), .ZN(n6207) );
  OAI211_X1 U7174 ( .C1(n6267), .C2(n6216), .A(n6208), .B(n6207), .ZN(U3137)
         );
  AOI22_X1 U7175 ( .A1(n6269), .A2(n6211), .B1(n6268), .B2(n6212), .ZN(n6210)
         );
  AOI22_X1 U7176 ( .A1(n6213), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n6270), 
        .B2(n2985), .ZN(n6209) );
  OAI211_X1 U7177 ( .C1(n6273), .C2(n6216), .A(n6210), .B(n6209), .ZN(U3138)
         );
  AOI22_X1 U7178 ( .A1(n6277), .A2(n6212), .B1(n6275), .B2(n6211), .ZN(n6215)
         );
  AOI22_X1 U7179 ( .A1(n6213), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n6279), 
        .B2(n2985), .ZN(n6214) );
  OAI211_X1 U7180 ( .C1(n6284), .C2(n6216), .A(n6215), .B(n6214), .ZN(U3139)
         );
  INV_X1 U7181 ( .A(n6217), .ZN(n6276) );
  AOI21_X1 U7182 ( .B1(n6219), .B2(n6218), .A(n6276), .ZN(n6227) );
  OAI22_X1 U7183 ( .A1(n6227), .A2(n6221), .B1(n6220), .B2(n6442), .ZN(n6274)
         );
  AOI22_X1 U7184 ( .A1(n6223), .A2(n6276), .B1(n6222), .B2(n6274), .ZN(n6236)
         );
  INV_X1 U7185 ( .A(n6224), .ZN(n6226) );
  AOI21_X1 U7186 ( .B1(n6226), .B2(n4472), .A(n6225), .ZN(n6229) );
  OAI21_X1 U7187 ( .B1(n6229), .B2(n6228), .A(n6227), .ZN(n6230) );
  OAI211_X1 U7188 ( .C1(n6233), .C2(n6232), .A(n6231), .B(n6230), .ZN(n6280)
         );
  AOI22_X1 U7189 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n6280), .B1(n6234), 
        .B2(n6278), .ZN(n6235) );
  OAI211_X1 U7190 ( .C1(n6237), .C2(n6283), .A(n6236), .B(n6235), .ZN(U3140)
         );
  AOI22_X1 U7191 ( .A1(n6239), .A2(n6276), .B1(n6238), .B2(n6274), .ZN(n6242)
         );
  AOI22_X1 U7192 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n6280), .B1(n6240), 
        .B2(n6278), .ZN(n6241) );
  OAI211_X1 U7193 ( .C1(n6243), .C2(n6283), .A(n6242), .B(n6241), .ZN(U3141)
         );
  AOI22_X1 U7194 ( .A1(n6245), .A2(n6274), .B1(n6276), .B2(n6244), .ZN(n6248)
         );
  AOI22_X1 U7195 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n6280), .B1(n6246), 
        .B2(n6278), .ZN(n6247) );
  OAI211_X1 U7196 ( .C1(n6249), .C2(n6283), .A(n6248), .B(n6247), .ZN(U3142)
         );
  AOI22_X1 U7197 ( .A1(n6251), .A2(n6276), .B1(n6250), .B2(n6274), .ZN(n6254)
         );
  AOI22_X1 U7198 ( .A1(INSTQUEUE_REG_15__3__SCAN_IN), .A2(n6280), .B1(n6252), 
        .B2(n6278), .ZN(n6253) );
  OAI211_X1 U7199 ( .C1(n6255), .C2(n6283), .A(n6254), .B(n6253), .ZN(U3143)
         );
  AOI22_X1 U7200 ( .A1(n6257), .A2(n6274), .B1(n6276), .B2(n6256), .ZN(n6260)
         );
  AOI22_X1 U7201 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n6280), .B1(n6258), 
        .B2(n6278), .ZN(n6259) );
  OAI211_X1 U7202 ( .C1(n6261), .C2(n6283), .A(n6260), .B(n6259), .ZN(U3144)
         );
  AOI22_X1 U7203 ( .A1(n6263), .A2(n6274), .B1(n6276), .B2(n6262), .ZN(n6266)
         );
  AOI22_X1 U7204 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n6280), .B1(n6264), 
        .B2(n6278), .ZN(n6265) );
  OAI211_X1 U7205 ( .C1(n6267), .C2(n6283), .A(n6266), .B(n6265), .ZN(U3145)
         );
  AOI22_X1 U7206 ( .A1(n6269), .A2(n6274), .B1(n6276), .B2(n6268), .ZN(n6272)
         );
  AOI22_X1 U7207 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n6280), .B1(n6270), 
        .B2(n6278), .ZN(n6271) );
  OAI211_X1 U7208 ( .C1(n6273), .C2(n6283), .A(n6272), .B(n6271), .ZN(U3146)
         );
  AOI22_X1 U7209 ( .A1(n6277), .A2(n6276), .B1(n6275), .B2(n6274), .ZN(n6282)
         );
  AOI22_X1 U7210 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n6280), .B1(n6279), 
        .B2(n6278), .ZN(n6281) );
  OAI211_X1 U7211 ( .C1(n6284), .C2(n6283), .A(n6282), .B(n6281), .ZN(U3147)
         );
  NOR2_X1 U7212 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6286) );
  OAI21_X1 U7213 ( .B1(n6287), .B2(n6286), .A(n6285), .ZN(n6288) );
  NOR2_X1 U7214 ( .A1(n6289), .A2(n6288), .ZN(n6290) );
  NAND2_X1 U7215 ( .A1(n6291), .A2(n6290), .ZN(n6292) );
  NOR2_X1 U7216 ( .A1(n6293), .A2(n6292), .ZN(n6316) );
  NAND2_X1 U7217 ( .A1(n6314), .A2(n6313), .ZN(n6310) );
  AOI22_X1 U7218 ( .A1(n6296), .A2(n6295), .B1(n6294), .B2(n3038), .ZN(n6420)
         );
  NAND2_X1 U7219 ( .A1(n6297), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6426) );
  NAND3_X1 U7220 ( .A1(n6420), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6426), .ZN(n6300) );
  OAI211_X1 U7221 ( .C1(n6301), .C2(n6300), .A(n6299), .B(n6298), .ZN(n6303)
         );
  NAND2_X1 U7222 ( .A1(n6301), .A2(n6300), .ZN(n6302) );
  NAND2_X1 U7223 ( .A1(n6303), .A2(n6302), .ZN(n6306) );
  INV_X1 U7224 ( .A(n6306), .ZN(n6304) );
  NOR2_X1 U7225 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6304), .ZN(n6307)
         );
  OAI22_X1 U7226 ( .A1(n6308), .A2(n6307), .B1(n6306), .B2(n6305), .ZN(n6309)
         );
  NAND2_X1 U7227 ( .A1(n6310), .A2(n6309), .ZN(n6312) );
  OAI211_X1 U7228 ( .C1(n6314), .C2(n6313), .A(n6312), .B(n6311), .ZN(n6315)
         );
  NAND2_X1 U7229 ( .A1(n6331), .A2(n6332), .ZN(n6318) );
  NAND2_X1 U7230 ( .A1(n4387), .A2(READY_N), .ZN(n6317) );
  NAND2_X1 U7231 ( .A1(n6318), .A2(n6317), .ZN(n6322) );
  OR2_X1 U7232 ( .A1(n6320), .A2(n6319), .ZN(n6321) );
  AOI21_X1 U7233 ( .B1(n6323), .B2(n6445), .A(n6338), .ZN(n6324) );
  INV_X1 U7234 ( .A(n6324), .ZN(n6327) );
  OAI21_X1 U7235 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6345), .A(n6412), .ZN(
        n6334) );
  NOR2_X1 U7236 ( .A1(n6325), .A2(n6334), .ZN(n6326) );
  MUX2_X1 U7237 ( .A(n6327), .B(n6326), .S(STATE2_REG_0__SCAN_IN), .Z(n6329)
         );
  OAI211_X1 U7238 ( .C1(n6331), .C2(n6330), .A(n6329), .B(n6328), .ZN(U3148)
         );
  AOI21_X1 U7239 ( .B1(n6333), .B2(n6345), .A(n6332), .ZN(n6337) );
  NAND3_X1 U7240 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6339), .A3(n6334), .ZN(
        n6335) );
  OAI211_X1 U7241 ( .C1(n6338), .C2(n6337), .A(n6336), .B(n6335), .ZN(U3149)
         );
  OAI211_X1 U7242 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6345), .A(n6410), .B(
        n6339), .ZN(n6341) );
  OAI21_X1 U7243 ( .B1(n6445), .B2(n6341), .A(n6340), .ZN(U3150) );
  AND2_X1 U7244 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6406), .ZN(U3151) );
  AND2_X1 U7245 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6406), .ZN(U3152) );
  AND2_X1 U7246 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6406), .ZN(U3153) );
  AND2_X1 U7247 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6406), .ZN(U3154) );
  AND2_X1 U7248 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6406), .ZN(U3155) );
  AND2_X1 U7249 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6406), .ZN(U3156) );
  AND2_X1 U7250 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6406), .ZN(U3157) );
  AND2_X1 U7251 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6406), .ZN(U3158) );
  INV_X1 U7252 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6573) );
  NOR2_X1 U7253 ( .A1(n6408), .A2(n6573), .ZN(U3159) );
  AND2_X1 U7254 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6406), .ZN(U3160) );
  AND2_X1 U7255 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6406), .ZN(U3161) );
  AND2_X1 U7256 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6406), .ZN(U3162) );
  AND2_X1 U7257 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6406), .ZN(U3163) );
  AND2_X1 U7258 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6406), .ZN(U3164) );
  AND2_X1 U7259 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6406), .ZN(U3165) );
  INV_X1 U7260 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6540) );
  NOR2_X1 U7261 ( .A1(n6408), .A2(n6540), .ZN(U3166) );
  AND2_X1 U7262 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6406), .ZN(U3167) );
  AND2_X1 U7263 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6406), .ZN(U3168) );
  AND2_X1 U7264 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6406), .ZN(U3169) );
  AND2_X1 U7265 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6406), .ZN(U3170) );
  AND2_X1 U7266 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6406), .ZN(U3171) );
  AND2_X1 U7267 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6406), .ZN(U3172) );
  AND2_X1 U7268 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6406), .ZN(U3173) );
  AND2_X1 U7269 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6406), .ZN(U3174) );
  AND2_X1 U7270 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6406), .ZN(U3175) );
  AND2_X1 U7271 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6406), .ZN(U3176) );
  AND2_X1 U7272 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6406), .ZN(U3177) );
  AND2_X1 U7273 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6406), .ZN(U3178) );
  AND2_X1 U7274 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6406), .ZN(U3179) );
  AND2_X1 U7275 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6406), .ZN(U3180) );
  NOR2_X1 U7276 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6342) );
  INV_X1 U7277 ( .A(HOLD), .ZN(n6348) );
  OAI21_X1 U7278 ( .B1(n6342), .B2(n6348), .A(REQUESTPENDING_REG_SCAN_IN), 
        .ZN(n6343) );
  INV_X1 U7279 ( .A(NA_N), .ZN(n6527) );
  AOI221_X1 U7280 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6527), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6356) );
  AOI21_X1 U7281 ( .B1(n6610), .B2(n6343), .A(n6356), .ZN(n6344) );
  OAI21_X1 U7282 ( .B1(n6345), .B2(n6349), .A(n6344), .ZN(U3181) );
  INV_X1 U7283 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6447) );
  NOR2_X1 U7284 ( .A1(n6351), .A2(n6447), .ZN(n6353) );
  AOI221_X1 U7285 ( .B1(n3175), .B2(n6353), .C1(n6348), .C2(n6353), .A(n6346), 
        .ZN(n6347) );
  NAND2_X1 U7286 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6354) );
  OAI211_X1 U7287 ( .C1(n6349), .C2(n6348), .A(n6347), .B(n6354), .ZN(U3182)
         );
  AOI21_X1 U7288 ( .B1(READY_N), .B2(n6527), .A(n6349), .ZN(n6350) );
  AOI21_X1 U7289 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(n3175), .A(n6350), 
        .ZN(n6352) );
  AOI21_X1 U7290 ( .B1(HOLD), .B2(n6352), .A(n6351), .ZN(n6357) );
  AOI21_X1 U7291 ( .B1(n6353), .B2(n6527), .A(STATE_REG_2__SCAN_IN), .ZN(n6355) );
  OAI22_X1 U7292 ( .A1(n6357), .A2(n6356), .B1(n6355), .B2(n6354), .ZN(U3183)
         );
  NOR2_X2 U7293 ( .A1(n3175), .A2(n6610), .ZN(n6609) );
  NOR2_X2 U7294 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6610), .ZN(n6608) );
  AOI22_X1 U7295 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6608), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6610), .ZN(n6358) );
  OAI21_X1 U7296 ( .B1(n6429), .B2(n6403), .A(n6358), .ZN(U3184) );
  AOI22_X1 U7297 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6610), .ZN(n6359) );
  OAI21_X1 U7298 ( .B1(n6360), .B2(n6398), .A(n6359), .ZN(U3185) );
  AOI22_X1 U7299 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6610), .ZN(n6361) );
  OAI21_X1 U7300 ( .B1(n6362), .B2(n6398), .A(n6361), .ZN(U3186) );
  AOI22_X1 U7301 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6610), .ZN(n6363) );
  OAI21_X1 U7302 ( .B1(n6364), .B2(n6398), .A(n6363), .ZN(U3187) );
  AOI22_X1 U7303 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6610), .ZN(n6365) );
  OAI21_X1 U7304 ( .B1(n6367), .B2(n6398), .A(n6365), .ZN(U3188) );
  AOI22_X1 U7305 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6608), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6610), .ZN(n6366) );
  OAI21_X1 U7306 ( .B1(n6367), .B2(n6403), .A(n6366), .ZN(U3189) );
  AOI22_X1 U7307 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6608), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6610), .ZN(n6368) );
  OAI21_X1 U7308 ( .B1(n6369), .B2(n6403), .A(n6368), .ZN(U3190) );
  AOI22_X1 U7309 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6610), .ZN(n6370) );
  OAI21_X1 U7310 ( .B1(n6502), .B2(n6398), .A(n6370), .ZN(U3191) );
  INV_X1 U7311 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n6529) );
  OAI222_X1 U7312 ( .A1(n6398), .A2(n6371), .B1(n6529), .B2(n6449), .C1(n6502), 
        .C2(n6403), .ZN(U3192) );
  INV_X1 U7313 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n6462) );
  OAI222_X1 U7314 ( .A1(n6403), .A2(n6371), .B1(n6462), .B2(n6449), .C1(n6373), 
        .C2(n6398), .ZN(U3193) );
  AOI22_X1 U7315 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6608), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6610), .ZN(n6372) );
  OAI21_X1 U7316 ( .B1(n6373), .B2(n6403), .A(n6372), .ZN(U3194) );
  AOI22_X1 U7317 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6608), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6610), .ZN(n6374) );
  OAI21_X1 U7318 ( .B1(n4946), .B2(n6403), .A(n6374), .ZN(U3195) );
  AOI22_X1 U7319 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6610), .ZN(n6375) );
  OAI21_X1 U7320 ( .B1(n6377), .B2(n6398), .A(n6375), .ZN(U3196) );
  AOI22_X1 U7321 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6608), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6610), .ZN(n6376) );
  OAI21_X1 U7322 ( .B1(n6377), .B2(n6403), .A(n6376), .ZN(U3197) );
  AOI22_X1 U7323 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6610), .ZN(n6378) );
  OAI21_X1 U7324 ( .B1(n6379), .B2(n6398), .A(n6378), .ZN(U3198) );
  AOI22_X1 U7325 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6610), .ZN(n6380) );
  OAI21_X1 U7326 ( .B1(n6381), .B2(n6398), .A(n6380), .ZN(U3199) );
  AOI22_X1 U7327 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6610), .ZN(n6382) );
  OAI21_X1 U7328 ( .B1(n6383), .B2(n6398), .A(n6382), .ZN(U3200) );
  AOI22_X1 U7329 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6610), .ZN(n6384) );
  OAI21_X1 U7330 ( .B1(n6386), .B2(n6398), .A(n6384), .ZN(U3201) );
  AOI22_X1 U7331 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6608), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6610), .ZN(n6385) );
  OAI21_X1 U7332 ( .B1(n6386), .B2(n6403), .A(n6385), .ZN(U3202) );
  AOI22_X1 U7333 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6610), .ZN(n6387) );
  OAI21_X1 U7334 ( .B1(n6388), .B2(n6398), .A(n6387), .ZN(U3203) );
  AOI22_X1 U7335 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6610), .ZN(n6389) );
  OAI21_X1 U7336 ( .B1(n6390), .B2(n6398), .A(n6389), .ZN(U3204) );
  AOI22_X1 U7337 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6608), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6610), .ZN(n6391) );
  OAI21_X1 U7338 ( .B1(n6392), .B2(n6403), .A(n6391), .ZN(U3206) );
  INV_X1 U7339 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6546) );
  OAI222_X1 U7340 ( .A1(n6398), .A2(n5281), .B1(n6546), .B2(n6449), .C1(n6393), 
        .C2(n6403), .ZN(U3207) );
  AOI22_X1 U7341 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6608), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6610), .ZN(n6394) );
  OAI21_X1 U7342 ( .B1(n5281), .B2(n6403), .A(n6394), .ZN(U3208) );
  AOI22_X1 U7343 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6610), .ZN(n6395) );
  OAI21_X1 U7344 ( .B1(n6396), .B2(n6398), .A(n6395), .ZN(U3209) );
  AOI22_X1 U7345 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6610), .ZN(n6397) );
  OAI21_X1 U7346 ( .B1(n6399), .B2(n6398), .A(n6397), .ZN(U3210) );
  INV_X1 U7347 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6524) );
  OAI222_X1 U7348 ( .A1(n6403), .A2(n6399), .B1(n6524), .B2(n6449), .C1(n6401), 
        .C2(n6398), .ZN(U3211) );
  AOI22_X1 U7349 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6608), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6610), .ZN(n6400) );
  OAI21_X1 U7350 ( .B1(n6401), .B2(n6403), .A(n6400), .ZN(U3212) );
  AOI22_X1 U7351 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6608), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6610), .ZN(n6402) );
  OAI21_X1 U7352 ( .B1(n6539), .B2(n6403), .A(n6402), .ZN(U3213) );
  MUX2_X1 U7353 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6449), .Z(U3445) );
  MUX2_X1 U7354 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6449), .Z(U3446) );
  INV_X1 U7355 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n6504) );
  AOI22_X1 U7356 ( .A1(n6449), .A2(n6404), .B1(n6504), .B2(n6610), .ZN(U3447)
         );
  MUX2_X1 U7357 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6449), .Z(U3448) );
  INV_X1 U7358 ( .A(n6407), .ZN(n6405) );
  AOI21_X1 U7359 ( .B1(n6428), .B2(n6406), .A(n6405), .ZN(U3451) );
  OAI21_X1 U7360 ( .B1(n6408), .B2(n6427), .A(n6407), .ZN(U3452) );
  INV_X1 U7361 ( .A(n6409), .ZN(n6411) );
  OAI211_X1 U7362 ( .C1(n6413), .C2(n6412), .A(n6411), .B(n6410), .ZN(U3453)
         );
  INV_X1 U7363 ( .A(n6414), .ZN(n6417) );
  OAI22_X1 U7364 ( .A1(n6417), .A2(n6425), .B1(n6416), .B2(n6415), .ZN(n6419)
         );
  MUX2_X1 U7365 ( .A(n6419), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6418), 
        .Z(U3456) );
  OAI22_X1 U7366 ( .A1(n6420), .A2(n6425), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6538), .ZN(n6422) );
  OAI22_X1 U7367 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6423), .B1(n6422), .B2(n6421), .ZN(n6424) );
  OAI21_X1 U7368 ( .B1(n6426), .B2(n6425), .A(n6424), .ZN(U3461) );
  OAI211_X1 U7369 ( .C1(n6428), .C2(n6436), .A(n6427), .B(n6437), .ZN(n6433)
         );
  OAI21_X1 U7370 ( .B1(n6436), .B2(n6429), .A(n6431), .ZN(n6430) );
  OAI21_X1 U7371 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(n6431), .A(n6430), .ZN(
        n6432) );
  NAND2_X1 U7372 ( .A1(n6433), .A2(n6432), .ZN(U3468) );
  INV_X1 U7373 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6434) );
  AOI22_X1 U7374 ( .A1(n6437), .A2(n6436), .B1(n6435), .B2(n6434), .ZN(U3469)
         );
  NAND2_X1 U7375 ( .A1(n6610), .A2(W_R_N_REG_SCAN_IN), .ZN(n6438) );
  OAI21_X1 U7376 ( .B1(n6610), .B2(READREQUEST_REG_SCAN_IN), .A(n6438), .ZN(
        U3470) );
  OAI211_X1 U7377 ( .C1(READY_N), .C2(n6440), .A(n6439), .B(n6452), .ZN(n6448)
         );
  AOI211_X1 U7378 ( .C1(n2954), .C2(n6455), .A(n6442), .B(n6441), .ZN(n6443)
         );
  NOR2_X1 U7379 ( .A1(n6443), .A2(n3297), .ZN(n6444) );
  OAI21_X1 U7380 ( .B1(n6445), .B2(n6444), .A(n6448), .ZN(n6446) );
  OAI21_X1 U7381 ( .B1(n6448), .B2(n6447), .A(n6446), .ZN(U3472) );
  MUX2_X1 U7382 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6449), .Z(U3473) );
  OAI21_X1 U7383 ( .B1(n6450), .B2(READREQUEST_REG_SCAN_IN), .A(n6452), .ZN(
        n6451) );
  OAI21_X1 U7384 ( .B1(n6453), .B2(n6452), .A(n6451), .ZN(U3474) );
  AOI22_X1 U7385 ( .A1(n6456), .A2(keyinput0), .B1(n6455), .B2(keyinput43), 
        .ZN(n6454) );
  OAI221_X1 U7386 ( .B1(n6456), .B2(keyinput0), .C1(n6455), .C2(keyinput43), 
        .A(n6454), .ZN(n6469) );
  INV_X1 U7387 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n6458) );
  AOI22_X1 U7388 ( .A1(n6459), .A2(keyinput24), .B1(keyinput32), .B2(n6458), 
        .ZN(n6457) );
  OAI221_X1 U7389 ( .B1(n6459), .B2(keyinput24), .C1(n6458), .C2(keyinput32), 
        .A(n6457), .ZN(n6468) );
  AOI22_X1 U7390 ( .A1(n6462), .A2(keyinput49), .B1(n6461), .B2(keyinput46), 
        .ZN(n6460) );
  OAI221_X1 U7391 ( .B1(n6462), .B2(keyinput49), .C1(n6461), .C2(keyinput46), 
        .A(n6460), .ZN(n6467) );
  INV_X1 U7392 ( .A(DATAI_17_), .ZN(n6465) );
  AOI22_X1 U7393 ( .A1(n6465), .A2(keyinput29), .B1(keyinput19), .B2(n6464), 
        .ZN(n6463) );
  OAI221_X1 U7394 ( .B1(n6465), .B2(keyinput29), .C1(n6464), .C2(keyinput19), 
        .A(n6463), .ZN(n6466) );
  NOR4_X1 U7395 ( .A1(n6469), .A2(n6468), .A3(n6467), .A4(n6466), .ZN(n6518)
         );
  AOI22_X1 U7396 ( .A1(n6594), .A2(keyinput33), .B1(keyinput56), .B2(n6471), 
        .ZN(n6470) );
  OAI221_X1 U7397 ( .B1(n6594), .B2(keyinput33), .C1(n6471), .C2(keyinput56), 
        .A(n6470), .ZN(n6484) );
  INV_X1 U7398 ( .A(DATAI_21_), .ZN(n6474) );
  INV_X1 U7399 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6473) );
  AOI22_X1 U7400 ( .A1(n6474), .A2(keyinput48), .B1(n6473), .B2(keyinput10), 
        .ZN(n6472) );
  OAI221_X1 U7401 ( .B1(n6474), .B2(keyinput48), .C1(n6473), .C2(keyinput10), 
        .A(n6472), .ZN(n6483) );
  INV_X1 U7402 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n6477) );
  AOI22_X1 U7403 ( .A1(n6477), .A2(keyinput18), .B1(keyinput55), .B2(n6476), 
        .ZN(n6475) );
  OAI221_X1 U7404 ( .B1(n6477), .B2(keyinput18), .C1(n6476), .C2(keyinput55), 
        .A(n6475), .ZN(n6482) );
  INV_X1 U7405 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n6478) );
  XOR2_X1 U7406 ( .A(n6478), .B(keyinput21), .Z(n6480) );
  XNOR2_X1 U7407 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .B(keyinput60), .ZN(n6479) );
  NAND2_X1 U7408 ( .A1(n6480), .A2(n6479), .ZN(n6481) );
  NOR4_X1 U7409 ( .A1(n6484), .A2(n6483), .A3(n6482), .A4(n6481), .ZN(n6517)
         );
  INV_X1 U7410 ( .A(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n6487) );
  INV_X1 U7411 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n6486) );
  AOI22_X1 U7412 ( .A1(n6487), .A2(keyinput3), .B1(n6486), .B2(keyinput16), 
        .ZN(n6485) );
  OAI221_X1 U7413 ( .B1(n6487), .B2(keyinput3), .C1(n6486), .C2(keyinput16), 
        .A(n6485), .ZN(n6500) );
  INV_X1 U7414 ( .A(UWORD_REG_10__SCAN_IN), .ZN(n6490) );
  AOI22_X1 U7415 ( .A1(n6490), .A2(keyinput27), .B1(n6489), .B2(keyinput54), 
        .ZN(n6488) );
  OAI221_X1 U7416 ( .B1(n6490), .B2(keyinput27), .C1(n6489), .C2(keyinput54), 
        .A(n6488), .ZN(n6499) );
  INV_X1 U7417 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6493) );
  AOI22_X1 U7418 ( .A1(n6493), .A2(keyinput14), .B1(keyinput12), .B2(n6492), 
        .ZN(n6491) );
  OAI221_X1 U7419 ( .B1(n6493), .B2(keyinput14), .C1(n6492), .C2(keyinput12), 
        .A(n6491), .ZN(n6498) );
  INV_X1 U7420 ( .A(DATAI_28_), .ZN(n6495) );
  AOI22_X1 U7421 ( .A1(n6496), .A2(keyinput13), .B1(keyinput1), .B2(n6495), 
        .ZN(n6494) );
  OAI221_X1 U7422 ( .B1(n6496), .B2(keyinput13), .C1(n6495), .C2(keyinput1), 
        .A(n6494), .ZN(n6497) );
  NOR4_X1 U7423 ( .A1(n6500), .A2(n6499), .A3(n6498), .A4(n6497), .ZN(n6516)
         );
  AOI22_X1 U7424 ( .A1(n6502), .A2(keyinput35), .B1(n3810), .B2(keyinput6), 
        .ZN(n6501) );
  OAI221_X1 U7425 ( .B1(n6502), .B2(keyinput35), .C1(n3810), .C2(keyinput6), 
        .A(n6501), .ZN(n6514) );
  INV_X1 U7426 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n6505) );
  AOI22_X1 U7427 ( .A1(n6505), .A2(keyinput63), .B1(keyinput28), .B2(n6504), 
        .ZN(n6503) );
  OAI221_X1 U7428 ( .B1(n6505), .B2(keyinput63), .C1(n6504), .C2(keyinput28), 
        .A(n6503), .ZN(n6513) );
  INV_X1 U7429 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n6507) );
  AOI22_X1 U7430 ( .A1(n6508), .A2(keyinput15), .B1(n6507), .B2(keyinput40), 
        .ZN(n6506) );
  OAI221_X1 U7431 ( .B1(n6508), .B2(keyinput15), .C1(n6507), .C2(keyinput40), 
        .A(n6506), .ZN(n6512) );
  XNOR2_X1 U7432 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .B(keyinput31), .ZN(n6510)
         );
  XNOR2_X1 U7433 ( .A(keyinput36), .B(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U7434 ( .A1(n6510), .A2(n6509), .ZN(n6511) );
  NOR4_X1 U7435 ( .A1(n6514), .A2(n6513), .A3(n6512), .A4(n6511), .ZN(n6515)
         );
  NAND4_X1 U7436 ( .A1(n6518), .A2(n6517), .A3(n6516), .A4(n6515), .ZN(n6584)
         );
  INV_X1 U7437 ( .A(LWORD_REG_11__SCAN_IN), .ZN(n6521) );
  INV_X1 U7438 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6520) );
  AOI22_X1 U7439 ( .A1(n6521), .A2(keyinput2), .B1(keyinput42), .B2(n6520), 
        .ZN(n6519) );
  OAI221_X1 U7440 ( .B1(n6521), .B2(keyinput2), .C1(n6520), .C2(keyinput42), 
        .A(n6519), .ZN(n6533) );
  AOI22_X1 U7441 ( .A1(n6524), .A2(keyinput34), .B1(n6523), .B2(keyinput17), 
        .ZN(n6522) );
  OAI221_X1 U7442 ( .B1(n6524), .B2(keyinput34), .C1(n6523), .C2(keyinput17), 
        .A(n6522), .ZN(n6532) );
  INV_X1 U7443 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n6526) );
  AOI22_X1 U7444 ( .A1(n6527), .A2(keyinput23), .B1(n6526), .B2(keyinput44), 
        .ZN(n6525) );
  OAI221_X1 U7445 ( .B1(n6527), .B2(keyinput23), .C1(n6526), .C2(keyinput44), 
        .A(n6525), .ZN(n6531) );
  AOI22_X1 U7446 ( .A1(n6529), .A2(keyinput25), .B1(n4619), .B2(keyinput20), 
        .ZN(n6528) );
  OAI221_X1 U7447 ( .B1(n6529), .B2(keyinput25), .C1(n4619), .C2(keyinput20), 
        .A(n6528), .ZN(n6530) );
  NOR4_X1 U7448 ( .A1(n6533), .A2(n6532), .A3(n6531), .A4(n6530), .ZN(n6582)
         );
  INV_X1 U7449 ( .A(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n6536) );
  INV_X1 U7450 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n6535) );
  AOI22_X1 U7451 ( .A1(n6536), .A2(keyinput30), .B1(keyinput47), .B2(n6535), 
        .ZN(n6534) );
  OAI221_X1 U7452 ( .B1(n6536), .B2(keyinput30), .C1(n6535), .C2(keyinput47), 
        .A(n6534), .ZN(n6549) );
  AOI22_X1 U7453 ( .A1(n6539), .A2(keyinput11), .B1(n6538), .B2(keyinput50), 
        .ZN(n6537) );
  OAI221_X1 U7454 ( .B1(n6539), .B2(keyinput11), .C1(n6538), .C2(keyinput50), 
        .A(n6537), .ZN(n6543) );
  XNOR2_X1 U7455 ( .A(n6540), .B(keyinput53), .ZN(n6542) );
  XOR2_X1 U7456 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .B(keyinput4), .Z(n6541) );
  OR3_X1 U7457 ( .A1(n6543), .A2(n6542), .A3(n6541), .ZN(n6548) );
  INV_X1 U7458 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n6545) );
  AOI22_X1 U7459 ( .A1(n6546), .A2(keyinput7), .B1(n6545), .B2(keyinput51), 
        .ZN(n6544) );
  OAI221_X1 U7460 ( .B1(n6546), .B2(keyinput7), .C1(n6545), .C2(keyinput51), 
        .A(n6544), .ZN(n6547) );
  NOR3_X1 U7461 ( .A1(n6549), .A2(n6548), .A3(n6547), .ZN(n6581) );
  INV_X1 U7462 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n6552) );
  AOI22_X1 U7463 ( .A1(n6552), .A2(keyinput38), .B1(keyinput22), .B2(n6551), 
        .ZN(n6550) );
  OAI221_X1 U7464 ( .B1(n6552), .B2(keyinput38), .C1(n6551), .C2(keyinput22), 
        .A(n6550), .ZN(n6564) );
  AOI22_X1 U7465 ( .A1(n4073), .A2(keyinput52), .B1(keyinput8), .B2(n6554), 
        .ZN(n6553) );
  OAI221_X1 U7466 ( .B1(n4073), .B2(keyinput52), .C1(n6554), .C2(keyinput8), 
        .A(n6553), .ZN(n6563) );
  INV_X1 U7467 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n6557) );
  AOI22_X1 U7468 ( .A1(n6557), .A2(keyinput37), .B1(n6556), .B2(keyinput26), 
        .ZN(n6555) );
  OAI221_X1 U7469 ( .B1(n6557), .B2(keyinput37), .C1(n6556), .C2(keyinput26), 
        .A(n6555), .ZN(n6562) );
  INV_X1 U7470 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n6560) );
  INV_X1 U7471 ( .A(LWORD_REG_12__SCAN_IN), .ZN(n6559) );
  AOI22_X1 U7472 ( .A1(n6560), .A2(keyinput41), .B1(keyinput58), .B2(n6559), 
        .ZN(n6558) );
  OAI221_X1 U7473 ( .B1(n6560), .B2(keyinput41), .C1(n6559), .C2(keyinput58), 
        .A(n6558), .ZN(n6561) );
  NOR4_X1 U7474 ( .A1(n6564), .A2(n6563), .A3(n6562), .A4(n6561), .ZN(n6580)
         );
  AOI22_X1 U7475 ( .A1(n4007), .A2(keyinput59), .B1(keyinput45), .B2(n6566), 
        .ZN(n6565) );
  OAI221_X1 U7476 ( .B1(n4007), .B2(keyinput59), .C1(n6566), .C2(keyinput45), 
        .A(n6565), .ZN(n6578) );
  AOI22_X1 U7477 ( .A1(n4414), .A2(keyinput57), .B1(keyinput5), .B2(n6568), 
        .ZN(n6567) );
  OAI221_X1 U7478 ( .B1(n4414), .B2(keyinput57), .C1(n6568), .C2(keyinput5), 
        .A(n6567), .ZN(n6577) );
  INV_X1 U7479 ( .A(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n6570) );
  AOI22_X1 U7480 ( .A1(n6571), .A2(keyinput61), .B1(n6570), .B2(keyinput62), 
        .ZN(n6569) );
  OAI221_X1 U7481 ( .B1(n6571), .B2(keyinput61), .C1(n6570), .C2(keyinput62), 
        .A(n6569), .ZN(n6576) );
  AOI22_X1 U7482 ( .A1(n6574), .A2(keyinput39), .B1(keyinput9), .B2(n6573), 
        .ZN(n6572) );
  OAI221_X1 U7483 ( .B1(n6574), .B2(keyinput39), .C1(n6573), .C2(keyinput9), 
        .A(n6572), .ZN(n6575) );
  NOR4_X1 U7484 ( .A1(n6578), .A2(n6577), .A3(n6576), .A4(n6575), .ZN(n6579)
         );
  NAND4_X1 U7485 ( .A1(n6582), .A2(n6581), .A3(n6580), .A4(n6579), .ZN(n6583)
         );
  NOR2_X1 U7486 ( .A1(n6584), .A2(n6583), .ZN(n6614) );
  NAND4_X1 U7487 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_23__SCAN_IN), .A4(
        ADDRESS_REG_9__SCAN_IN), .ZN(n6588) );
  NAND4_X1 U7488 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(EAX_REG_0__SCAN_IN), .A3(EAX_REG_4__SCAN_IN), .A4(LWORD_REG_11__SCAN_IN), .ZN(n6587) );
  NAND4_X1 U7489 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .A3(DATAO_REG_27__SCAN_IN), .A4(
        LWORD_REG_12__SCAN_IN), .ZN(n6586) );
  NAND4_X1 U7490 ( .A1(STATE2_REG_1__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .A3(
        DATAI_17_), .A4(DATAO_REG_28__SCAN_IN), .ZN(n6585) );
  NOR4_X1 U7491 ( .A1(n6588), .A2(n6587), .A3(n6586), .A4(n6585), .ZN(n6607)
         );
  NOR4_X1 U7492 ( .A1(ADDRESS_REG_8__SCAN_IN), .A2(BE_N_REG_1__SCAN_IN), .A3(
        ADDRESS_REG_23__SCAN_IN), .A4(ADDRESS_REG_21__SCAN_IN), .ZN(n6592) );
  NOR4_X1 U7493 ( .A1(STATEBS16_REG_SCAN_IN), .A2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .A3(EAX_REG_8__SCAN_IN), .A4(NA_N), 
        .ZN(n6591) );
  NOR4_X1 U7494 ( .A1(EAX_REG_14__SCAN_IN), .A2(DATAI_15_), .A3(
        DATAO_REG_26__SCAN_IN), .A4(UWORD_REG_10__SCAN_IN), .ZN(n6590) );
  NOR4_X1 U7495 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(EBX_REG_5__SCAN_IN), 
        .A3(EAX_REG_15__SCAN_IN), .A4(DATAI_0_), .ZN(n6589) );
  NAND4_X1 U7496 ( .A1(n6592), .A2(n6591), .A3(n6590), .A4(n6589), .ZN(n6600)
         );
  NAND3_X1 U7497 ( .A1(n6594), .A2(n6593), .A3(n3810), .ZN(n6599) );
  NOR4_X1 U7498 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(
        INSTQUEUE_REG_7__2__SCAN_IN), .A3(INSTQUEUE_REG_5__2__SCAN_IN), .A4(
        EBX_REG_8__SCAN_IN), .ZN(n6597) );
  NOR4_X1 U7499 ( .A1(INSTQUEUE_REG_2__6__SCAN_IN), .A2(
        INSTQUEUE_REG_8__7__SCAN_IN), .A3(EAX_REG_22__SCAN_IN), .A4(DATAI_3_), 
        .ZN(n6596) );
  NOR3_X1 U7500 ( .A1(EBX_REG_25__SCAN_IN), .A2(EAX_REG_29__SCAN_IN), .A3(
        DATAI_28_), .ZN(n6595) );
  NAND4_X1 U7501 ( .A1(n6597), .A2(n6596), .A3(ADDRESS_REG_27__SCAN_IN), .A4(
        n6595), .ZN(n6598) );
  NOR4_X1 U7502 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n6600), .A3(n6599), 
        .A4(n6598), .ZN(n6606) );
  NAND4_X1 U7503 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A3(EBX_REG_7__SCAN_IN), .A4(
        EBX_REG_16__SCAN_IN), .ZN(n6604) );
  NAND4_X1 U7504 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(
        INSTQUEUE_REG_12__4__SCAN_IN), .A3(INSTQUEUE_REG_8__4__SCAN_IN), .A4(
        INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n6603) );
  NAND4_X1 U7505 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(
        INSTQUEUE_REG_5__6__SCAN_IN), .A3(INSTQUEUE_REG_10__3__SCAN_IN), .A4(
        DATAI_21_), .ZN(n6602) );
  NAND4_X1 U7506 ( .A1(INSTQUEUE_REG_2__7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_2__SCAN_IN), .A3(EBX_REG_19__SCAN_IN), .A4(
        REIP_REG_30__SCAN_IN), .ZN(n6601) );
  NOR4_X1 U7507 ( .A1(n6604), .A2(n6603), .A3(n6602), .A4(n6601), .ZN(n6605)
         );
  NAND3_X1 U7508 ( .A1(n6607), .A2(n6606), .A3(n6605), .ZN(n6612) );
  AOI222_X1 U7509 ( .A1(n6610), .A2(ADDRESS_REG_21__SCAN_IN), .B1(
        REIP_REG_22__SCAN_IN), .B2(n6609), .C1(REIP_REG_23__SCAN_IN), .C2(
        n6608), .ZN(n6611) );
  XNOR2_X1 U7510 ( .A(n6612), .B(n6611), .ZN(n6613) );
  XNOR2_X1 U7511 ( .A(n6614), .B(n6613), .ZN(U3205) );
  OR2_X1 U5126 ( .A1(n4160), .A2(n4161), .ZN(n4162) );
  CLKBUF_X1 U3414 ( .A(n3128), .Z(n2974) );
  CLKBUF_X1 U3435 ( .A(n3904), .Z(n2970) );
  CLKBUF_X1 U34700 ( .A(n5100), .Z(n2957) );
  CLKBUF_X1 U3509 ( .A(n5185), .Z(n5186) );
  CLKBUF_X1 U3511 ( .A(n3353), .Z(n2960) );
  CLKBUF_X1 U3515 ( .A(n4417), .Z(n2971) );
  CLKBUF_X1 U3516 ( .A(n4471), .Z(n4472) );
  CLKBUF_X1 U3551 ( .A(n5085), .Z(n5086) );
  CLKBUF_X1 U3776 ( .A(n5112), .Z(n5113) );
  CLKBUF_X1 U3820 ( .A(n5348), .Z(n2961) );
  CLKBUF_X1 U6226 ( .A(n5803), .Z(n5795) );
  CLKBUF_X1 U6249 ( .A(n3137), .Z(n3834) );
endmodule

