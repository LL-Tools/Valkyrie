

module b21_C_gen_AntiSAT_k_128_8 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2, 
        keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7, 
        keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12, 
        keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17, 
        keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22, 
        keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27, 
        keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32, 
        keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37, 
        keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42, 
        keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47, 
        keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52, 
        keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57, 
        keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62, 
        keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3, 
        keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8, 
        keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13, 
        keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18, 
        keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23, 
        keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28, 
        keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33, 
        keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38, 
        keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43, 
        keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48, 
        keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53, 
        keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58, 
        keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63, 
        ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, 
        ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, 
        ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, 
        ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, 
        U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, 
        P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, 
        P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, 
        P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, 
        P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, 
        P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, 
        P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, 
        P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, 
        P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, 
        P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, 
        P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, 
        P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, 
        P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, 
        P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, 
        P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, 
        P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, 
        P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223;

  INV_X2 U4817 ( .A(n8721), .ZN(n8689) );
  NAND3_X1 U4819 ( .A1(n5603), .A2(n5602), .A3(n5601), .ZN(n6385) );
  INV_X1 U4820 ( .A(n4312), .ZN(n5904) );
  NAND4_X2 U4821 ( .A1(n4894), .A2(n4893), .A3(n4892), .A4(n4891), .ZN(n9331)
         );
  AND2_X1 U4822 ( .A1(n4866), .A2(n4867), .ZN(n4933) );
  AND2_X2 U4823 ( .A1(n9219), .A2(n9214), .ZN(n5872) );
  AND4_X1 U4824 ( .A1(n5522), .A2(n5521), .A3(n5520), .A4(n5519), .ZN(n4839)
         );
  NAND2_X2 U4825 ( .A1(n4674), .A2(n4673), .ZN(n4928) );
  INV_X1 U4826 ( .A(n8631), .ZN(n8606) );
  INV_X1 U4827 ( .A(n4314), .ZN(n5979) );
  INV_X1 U4828 ( .A(n6498), .ZN(n6884) );
  INV_X1 U4829 ( .A(n8952), .ZN(n5892) );
  INV_X2 U4830 ( .A(n4313), .ZN(n4318) );
  NAND2_X1 U4831 ( .A1(n5958), .A2(n8093), .ZN(n8207) );
  XNOR2_X1 U4832 ( .A(n5545), .B(n5544), .ZN(n5547) );
  NAND2_X1 U4833 ( .A1(n5948), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5949) );
  INV_X1 U4834 ( .A(n4932), .ZN(n5993) );
  OR2_X1 U4835 ( .A1(n4874), .A2(n4736), .ZN(n4864) );
  NAND2_X1 U4836 ( .A1(n5540), .A2(n5525), .ZN(n6293) );
  INV_X1 U4837 ( .A(n4933), .ZN(n5997) );
  AND4_X1 U4838 ( .A1(n4919), .A2(n4918), .A3(n4917), .A4(n4916), .ZN(n7095)
         );
  NAND2_X1 U4839 ( .A1(n5396), .A2(n5395), .ZN(n9401) );
  XNOR2_X1 U4840 ( .A(n5392), .B(n5391), .ZN(n7940) );
  NAND4_X1 U4841 ( .A1(n5613), .A2(n5612), .A3(n5611), .A4(n5610), .ZN(n5620)
         );
  INV_X1 U4843 ( .A(n7098), .ZN(n6798) );
  NAND4_X2 U4844 ( .A1(n4872), .A2(n4871), .A3(n4870), .A4(n4869), .ZN(n6423)
         );
  NAND2_X1 U4845 ( .A1(n5547), .A2(n9219), .ZN(n4312) );
  NAND2_X1 U4846 ( .A1(n9214), .A2(n5546), .ZN(n4313) );
  MUX2_X2 U4847 ( .A(n8318), .B(n8317), .S(n8415), .Z(n8328) );
  OAI21_X2 U4848 ( .B1(n7815), .B2(n7814), .A(n7823), .ZN(n7992) );
  NAND2_X2 U4849 ( .A1(n7681), .A2(n7680), .ZN(n7815) );
  XNOR2_X2 U4850 ( .A(n5949), .B(P2_IR_REG_20__SCAN_IN), .ZN(n8238) );
  NOR2_X2 U4852 ( .A1(n7718), .A2(n7719), .ZN(n7717) );
  OAI21_X2 U4853 ( .B1(n7622), .B2(n8221), .A(n8139), .ZN(n7718) );
  XNOR2_X2 U4854 ( .A(n9329), .B(n6494), .ZN(n6638) );
  INV_X2 U4855 ( .A(n5952), .ZN(n10055) );
  OAI21_X2 U4856 ( .B1(n5135), .B2(n4691), .A(n4689), .ZN(n5194) );
  NAND2_X4 U4857 ( .A1(n4868), .A2(n4867), .ZN(n4989) );
  NAND2_X1 U4858 ( .A1(n6463), .A2(n6379), .ZN(n6375) );
  INV_X2 U4859 ( .A(n6692), .ZN(n6463) );
  BUF_X1 U4861 ( .A(n4320), .Z(n4316) );
  BUF_X1 U4862 ( .A(n4320), .Z(n4317) );
  AND2_X1 U4863 ( .A1(n5547), .A2(n5546), .ZN(n5598) );
  INV_X1 U4864 ( .A(n4319), .ZN(n4320) );
  INV_X1 U4865 ( .A(n5598), .ZN(n4319) );
  INV_X1 U4866 ( .A(n6949), .ZN(n10086) );
  XNOR2_X2 U4867 ( .A(n4642), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8591) );
  AND2_X1 U4868 ( .A1(n5600), .A2(n5599), .ZN(n5603) );
  NAND2_X1 U4869 ( .A1(n8660), .A2(n8659), .ZN(n9299) );
  OR2_X1 U4870 ( .A1(n5849), .A2(n8759), .ZN(n5861) );
  AND2_X1 U4871 ( .A1(n6470), .A2(n6487), .ZN(n6473) );
  NAND2_X1 U4872 ( .A1(n6380), .A2(n6375), .ZN(n6951) );
  NAND2_X1 U4873 ( .A1(n5650), .A2(n5649), .ZN(n6736) );
  INV_X2 U4874 ( .A(n6498), .ZN(n8706) );
  INV_X1 U4875 ( .A(n6910), .ZN(n6379) );
  NAND2_X2 U4876 ( .A1(n5953), .A2(n8242), .ZN(n10081) );
  NAND2_X2 U4877 ( .A1(n6293), .A2(n8246), .ZN(n5576) );
  CLKBUF_X3 U4878 ( .A(n4928), .Z(n6066) );
  AND2_X1 U4879 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7612) );
  AND2_X1 U4880 ( .A1(n4452), .A2(n4449), .ZN(n8595) );
  AOI21_X1 U4881 ( .B1(n5977), .B2(n10049), .A(n5976), .ZN(n9130) );
  AND2_X1 U4882 ( .A1(n4664), .A2(n4666), .ZN(n9314) );
  XNOR2_X1 U4883 ( .A(n4808), .B(n8205), .ZN(n9131) );
  NOR2_X1 U4884 ( .A1(n8765), .A2(n8618), .ZN(n8619) );
  NOR2_X1 U4885 ( .A1(n4585), .A2(n4584), .ZN(n8963) );
  NAND2_X1 U4886 ( .A1(n9025), .A2(n4592), .ZN(n4588) );
  OAI22_X1 U4887 ( .A1(n9108), .A2(n5801), .B1(n9115), .B2(n7956), .ZN(n9092)
         );
  NAND2_X1 U4888 ( .A1(n4590), .A2(n8175), .ZN(n4584) );
  AND2_X1 U4889 ( .A1(n4810), .A2(n4377), .ZN(n7908) );
  NAND2_X1 U4890 ( .A1(n5848), .A2(n5847), .ZN(n9146) );
  NAND2_X1 U4891 ( .A1(n4764), .A2(n4766), .ZN(n8788) );
  OR2_X1 U4892 ( .A1(n5839), .A2(n8771), .ZN(n5849) );
  NAND2_X1 U4893 ( .A1(n5138), .A2(n5137), .ZN(n7932) );
  NAND2_X1 U4894 ( .A1(n5078), .A2(n5077), .ZN(n9845) );
  NAND2_X1 U4895 ( .A1(n5718), .A2(n5717), .ZN(n10141) );
  AND2_X1 U4896 ( .A1(n8114), .A2(n8113), .ZN(n8215) );
  INV_X2 U4897 ( .A(n9049), .ZN(n10070) );
  AND2_X2 U4898 ( .A1(n6922), .A2(n9598), .ZN(n9939) );
  AND2_X1 U4899 ( .A1(n8485), .A2(n8477), .ZN(n8430) );
  AND3_X1 U4900 ( .A1(n5586), .A2(n5585), .A3(n5584), .ZN(n6692) );
  NAND2_X2 U4901 ( .A1(n6419), .A2(n6418), .ZN(n8721) );
  OAI211_X2 U4902 ( .C1(n6067), .C2(n5642), .A(n5581), .B(n5580), .ZN(n6910)
         );
  NAND4_X1 U4903 ( .A1(n4904), .A2(n4903), .A3(n4902), .A4(n4901), .ZN(n9329)
         );
  OAI211_X1 U4904 ( .C1(n6078), .C2(n5642), .A(n5607), .B(n5606), .ZN(n6949)
         );
  OAI211_X1 U4905 ( .C1(n6076), .C2(n5642), .A(n5619), .B(n5618), .ZN(n10056)
         );
  OR2_X1 U4906 ( .A1(n4989), .A2(n6835), .ZN(n4869) );
  AND2_X1 U4907 ( .A1(n8583), .A2(n9408), .ZN(n5477) );
  NAND2_X1 U4908 ( .A1(n4866), .A2(n9779), .ZN(n4932) );
  NAND2_X1 U4909 ( .A1(n4879), .A2(n4878), .ZN(n8588) );
  OR2_X1 U4910 ( .A1(n9769), .A2(n5181), .ZN(n4863) );
  NAND2_X1 U4911 ( .A1(n4864), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4540) );
  MUX2_X1 U4912 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5524), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n5525) );
  OR2_X1 U4913 ( .A1(n4877), .A2(n5181), .ZN(n4616) );
  OR2_X1 U4914 ( .A1(n5543), .A2(n5765), .ZN(n5545) );
  XNOR2_X1 U4915 ( .A(n4980), .B(n4966), .ZN(n4978) );
  OAI21_X1 U4916 ( .B1(n4770), .B2(n4366), .A(n4323), .ZN(n8246) );
  OR2_X1 U4917 ( .A1(n5020), .A2(n5019), .ZN(n5043) );
  AOI21_X1 U4918 ( .B1(n5526), .B2(P2_IR_REG_31__SCAN_IN), .A(n4828), .ZN(
        n4770) );
  OR2_X2 U4919 ( .A1(n6066), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9221) );
  AND2_X1 U4920 ( .A1(n5917), .A2(n4611), .ZN(n4610) );
  NOR2_X1 U4921 ( .A1(n4827), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4614) );
  CLKBUF_X1 U4922 ( .A(n5571), .Z(n5614) );
  NOR2_X1 U4923 ( .A1(n4970), .A2(n4969), .ZN(n4987) );
  AND4_X1 U4924 ( .A1(n5177), .A2(n5406), .A3(n5198), .A4(n4855), .ZN(n4856)
         );
  AND4_X1 U4925 ( .A1(n5513), .A2(n5512), .A3(n5511), .A4(n5510), .ZN(n5518)
         );
  AND4_X1 U4926 ( .A1(n5515), .A2(n5644), .A3(n5514), .A4(n5572), .ZN(n5517)
         );
  AND2_X1 U4927 ( .A1(n5604), .A2(n5516), .ZN(n5571) );
  NAND2_X1 U4928 ( .A1(n4881), .A2(n7612), .ZN(n4673) );
  NOR2_X1 U4929 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4854) );
  NOR2_X1 U4930 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4853) );
  NOR2_X1 U4931 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4851) );
  NOR2_X1 U4932 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4852) );
  INV_X1 U4933 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5644) );
  NOR2_X1 U4934 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5604) );
  NOR2_X1 U4935 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4905) );
  INV_X4 U4936 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X2 U4937 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NOR2_X2 U4938 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7613) );
  NOR2_X1 U4939 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5510) );
  NOR2_X1 U4940 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5511) );
  NOR2_X1 U4941 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5512) );
  INV_X1 U4942 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5177) );
  NOR2_X1 U4943 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5515) );
  NOR3_X1 U4944 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5522) );
  INV_X1 U4945 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5406) );
  INV_X1 U4946 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5198) );
  INV_X1 U4947 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5453) );
  AND2_X1 U4948 ( .A1(n6384), .A2(n6919), .ZN(n6376) );
  NAND2_X1 U4949 ( .A1(n6385), .A2(n10086), .ZN(n8093) );
  OAI21_X1 U4950 ( .B1(n8742), .B2(n8615), .A(n8614), .ZN(n8620) );
  INV_X4 U4951 ( .A(n4312), .ZN(n4321) );
  AND2_X4 U4952 ( .A1(n5576), .A2(n6066), .ZN(n5630) );
  AND2_X1 U4953 ( .A1(n9437), .A2(n4709), .ZN(n4708) );
  NAND2_X1 U4954 ( .A1(n4342), .A2(n5335), .ZN(n4709) );
  NAND2_X1 U4955 ( .A1(n5272), .A2(n5271), .ZN(n4717) );
  NAND2_X1 U4956 ( .A1(n4798), .A2(n4797), .ZN(n8981) );
  AOI21_X1 U4957 ( .B1(n4799), .B2(n4800), .A(n8986), .ZN(n4797) );
  OR2_X1 U4958 ( .A1(n7716), .A2(n4813), .ZN(n4810) );
  NAND2_X1 U4959 ( .A1(n4814), .A2(n7719), .ZN(n4813) );
  NAND2_X1 U4960 ( .A1(n4999), .A2(n5376), .ZN(n4982) );
  AOI21_X1 U4961 ( .B1(n8331), .B2(n8402), .A(n9836), .ZN(n4431) );
  NAND2_X1 U4962 ( .A1(n8332), .A2(n8415), .ZN(n4432) );
  INV_X1 U4963 ( .A(n8198), .ZN(n8201) );
  NOR2_X1 U4964 ( .A1(n8734), .A2(n4761), .ZN(n4760) );
  INV_X1 U4965 ( .A(n8802), .ZN(n4761) );
  NOR2_X1 U4966 ( .A1(n9127), .A2(n5912), .ZN(n8189) );
  NOR2_X1 U4967 ( .A1(n9005), .A2(n4804), .ZN(n4801) );
  INV_X1 U4968 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5516) );
  INV_X1 U4969 ( .A(n6622), .ZN(n4641) );
  INV_X1 U4970 ( .A(n8467), .ZN(n4583) );
  NOR2_X1 U4971 ( .A1(n9575), .A2(n9566), .ZN(n9539) );
  NOR2_X1 U4972 ( .A1(n5147), .A2(n4726), .ZN(n4725) );
  INV_X1 U4973 ( .A(n4728), .ZN(n4726) );
  INV_X1 U4974 ( .A(n4866), .ZN(n4868) );
  INV_X1 U4975 ( .A(n9779), .ZN(n4867) );
  NAND2_X1 U4976 ( .A1(n8037), .A2(n8036), .ZN(n8042) );
  OAI21_X1 U4977 ( .B1(n5358), .B2(n5357), .A(n5356), .ZN(n5373) );
  AND4_X1 U4978 ( .A1(n4856), .A2(n4859), .A3(n4561), .A4(n4374), .ZN(n4558)
         );
  INV_X1 U4979 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4734) );
  OAI21_X1 U4980 ( .B1(n5194), .B2(n4478), .A(n4476), .ZN(n5233) );
  INV_X1 U4981 ( .A(n4479), .ZN(n4478) );
  AOI21_X1 U4982 ( .B1(n4477), .B2(n4479), .A(n4385), .ZN(n4476) );
  NOR2_X1 U4983 ( .A1(n5213), .A2(n4480), .ZN(n4479) );
  INV_X1 U4984 ( .A(n4690), .ZN(n4689) );
  OAI21_X1 U4985 ( .B1(n4693), .B2(n4691), .A(n5171), .ZN(n4690) );
  NAND2_X1 U4986 ( .A1(n4692), .A2(n5151), .ZN(n4691) );
  NAND2_X1 U4987 ( .A1(n4860), .A2(n5136), .ZN(n5180) );
  OAI21_X1 U4988 ( .B1(n5113), .B2(n5112), .A(n5111), .ZN(n5133) );
  INV_X1 U4989 ( .A(n4775), .ZN(n4774) );
  OAI21_X1 U4990 ( .B1(n4341), .B2(n4776), .A(n7970), .ZN(n4775) );
  OAI22_X1 U4991 ( .A1(n8734), .A2(n4762), .B1(n8628), .B2(n8629), .ZN(n4759)
         );
  INV_X1 U4992 ( .A(n4749), .ZN(n4745) );
  XNOR2_X1 U4993 ( .A(n8606), .B(n6902), .ZN(n6663) );
  NAND2_X1 U4994 ( .A1(n10015), .A2(n10010), .ZN(n4763) );
  NAND2_X1 U4995 ( .A1(n8621), .A2(n4750), .ZN(n4749) );
  INV_X1 U4996 ( .A(n8622), .ZN(n4750) );
  XNOR2_X1 U4997 ( .A(n8053), .B(n5979), .ZN(n4594) );
  OAI21_X1 U4998 ( .B1(n8052), .B2(n8236), .A(n8199), .ZN(n8053) );
  INV_X1 U4999 ( .A(n5872), .ZN(n5911) );
  OAI21_X1 U5000 ( .B1(n6368), .B2(n10161), .A(n4399), .ZN(n6364) );
  NAND2_X1 U5001 ( .A1(n6368), .A2(n10161), .ZN(n4399) );
  AND2_X1 U5002 ( .A1(n4393), .A2(n4392), .ZN(n6550) );
  NAND2_X1 U5003 ( .A1(n6547), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4392) );
  OR2_X1 U5004 ( .A1(n9135), .A2(n8966), .ZN(n5879) );
  XNOR2_X1 U5005 ( .A(n9135), .B(n8057), .ZN(n8945) );
  NAND2_X1 U5006 ( .A1(n5868), .A2(n8989), .ZN(n5869) );
  NOR2_X1 U5007 ( .A1(n9161), .A2(n9063), .ZN(n5836) );
  INV_X1 U5008 ( .A(n8225), .ZN(n4809) );
  NAND2_X1 U5009 ( .A1(n7010), .A2(n8211), .ZN(n4830) );
  NAND2_X1 U5010 ( .A1(n5576), .A2(n5527), .ZN(n5642) );
  AND2_X1 U5011 ( .A1(n6322), .A2(n6321), .ZN(n6326) );
  AND2_X1 U5012 ( .A1(n4667), .A2(n4665), .ZN(n4664) );
  INV_X1 U5013 ( .A(n9317), .ZN(n4665) );
  NAND2_X1 U5014 ( .A1(n5405), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5409) );
  AND2_X1 U5015 ( .A1(n9731), .A2(n8411), .ZN(n8420) );
  OR2_X1 U5016 ( .A1(n6000), .A2(n8409), .ZN(n6013) );
  NOR2_X1 U5017 ( .A1(n8463), .A2(n8575), .ZN(n8453) );
  NAND2_X1 U5018 ( .A1(n4704), .A2(n4703), .ZN(n5493) );
  AOI21_X1 U5019 ( .B1(n4368), .B2(n4705), .A(n4329), .ZN(n4703) );
  NAND2_X1 U5020 ( .A1(n4711), .A2(n4710), .ZN(n9468) );
  AOI21_X1 U5021 ( .B1(n4328), .B2(n4715), .A(n4358), .ZN(n4710) );
  AOI21_X1 U5022 ( .B1(n9612), .B2(n5170), .A(n5169), .ZN(n9594) );
  NAND2_X1 U5023 ( .A1(n6828), .A2(n4899), .ZN(n6637) );
  INV_X1 U5024 ( .A(n8397), .ZN(n5244) );
  INV_X1 U5025 ( .A(n4999), .ZN(n6058) );
  XNOR2_X1 U5026 ( .A(n5233), .B(n5231), .ZN(n6974) );
  NAND2_X1 U5027 ( .A1(n5504), .A2(n5503), .ZN(n9406) );
  AND2_X1 U5028 ( .A1(n5502), .A2(n5501), .ZN(n5503) );
  NAND2_X2 U5029 ( .A1(n5383), .A2(n5382), .ZN(n5390) );
  NAND2_X1 U5030 ( .A1(n7940), .A2(n4998), .ZN(n5383) );
  INV_X1 U5031 ( .A(n8080), .ZN(n4537) );
  INV_X1 U5032 ( .A(n8108), .ZN(n4538) );
  INV_X1 U5033 ( .A(n8349), .ZN(n4428) );
  NAND2_X1 U5034 ( .A1(n4430), .A2(n8343), .ZN(n4429) );
  NAND2_X1 U5035 ( .A1(n4432), .A2(n4431), .ZN(n4430) );
  AOI21_X1 U5036 ( .B1(n8155), .B2(n4517), .A(n4516), .ZN(n4515) );
  INV_X1 U5037 ( .A(n8156), .ZN(n4516) );
  INV_X1 U5038 ( .A(n4518), .ZN(n4517) );
  INV_X1 U5039 ( .A(n8173), .ZN(n4687) );
  OAI21_X1 U5040 ( .B1(n4523), .B2(n4522), .A(n4683), .ZN(n4682) );
  INV_X1 U5041 ( .A(n4684), .ZN(n4683) );
  NAND2_X1 U5042 ( .A1(n8986), .A2(n8174), .ZN(n4522) );
  AOI21_X1 U5043 ( .B1(n8171), .B2(n4353), .A(n4524), .ZN(n4523) );
  NAND2_X1 U5044 ( .A1(n4423), .A2(n4422), .ZN(n4483) );
  AND2_X1 U5045 ( .A1(n8518), .A2(n8415), .ZN(n4422) );
  NAND2_X1 U5046 ( .A1(n4424), .A2(n8508), .ZN(n4423) );
  OR2_X1 U5047 ( .A1(n8368), .A2(n8367), .ZN(n4424) );
  OAI21_X1 U5048 ( .B1(n8386), .B2(n4440), .A(n8378), .ZN(n8389) );
  INV_X1 U5049 ( .A(n4792), .ZN(n4791) );
  OAI21_X1 U5050 ( .B1(n4794), .B2(n4793), .A(n8749), .ZN(n4792) );
  INV_X1 U5051 ( .A(n8600), .ZN(n4793) );
  INV_X1 U5052 ( .A(n8192), .ZN(n4513) );
  OAI21_X1 U5053 ( .B1(n8196), .B2(n8191), .A(n4510), .ZN(n4507) );
  AND2_X1 U5054 ( .A1(n4675), .A2(n4511), .ZN(n4510) );
  NAND2_X1 U5055 ( .A1(n8197), .A2(n8186), .ZN(n4511) );
  NOR2_X1 U5056 ( .A1(n9135), .A2(n9140), .ZN(n4489) );
  INV_X1 U5057 ( .A(n6385), .ZN(n5608) );
  NAND2_X1 U5058 ( .A1(n5523), .A2(n4828), .ZN(n4827) );
  NOR2_X1 U5059 ( .A1(n9752), .A2(n9533), .ZN(n4620) );
  NOR2_X1 U5060 ( .A1(n4994), .A2(n4445), .ZN(n4444) );
  INV_X1 U5061 ( .A(n4978), .ZN(n4445) );
  INV_X1 U5062 ( .A(n4981), .ZN(n4447) );
  NOR2_X1 U5063 ( .A1(n8640), .A2(n4488), .ZN(n4487) );
  INV_X1 U5064 ( .A(n4489), .ZN(n4488) );
  NOR2_X1 U5065 ( .A1(n9164), .A2(n4492), .ZN(n4491) );
  INV_X1 U5066 ( .A(n4493), .ZN(n4492) );
  NOR2_X1 U5067 ( .A1(n9171), .A2(n9177), .ZN(n4493) );
  AND2_X1 U5068 ( .A1(n9177), .A2(n9075), .ZN(n8158) );
  INV_X1 U5069 ( .A(n4609), .ZN(n4608) );
  NAND2_X1 U5070 ( .A1(n4607), .A2(n8066), .ZN(n4606) );
  NAND2_X1 U5071 ( .A1(n8154), .A2(n8150), .ZN(n4607) );
  OR2_X1 U5072 ( .A1(n9191), .A2(n7955), .ZN(n8151) );
  OR2_X1 U5073 ( .A1(n7727), .A2(n7891), .ZN(n8142) );
  NOR2_X1 U5074 ( .A1(n7727), .A2(n7048), .ZN(n4499) );
  NAND2_X1 U5075 ( .A1(n8215), .A2(n8110), .ZN(n4601) );
  NAND2_X1 U5076 ( .A1(n8248), .A2(n5979), .ZN(n8239) );
  NOR2_X1 U5077 ( .A1(n8676), .A2(n9279), .ZN(n4832) );
  INV_X1 U5078 ( .A(n4417), .ZN(n7213) );
  NOR2_X1 U5079 ( .A1(n4628), .A2(n5390), .ZN(n4627) );
  INV_X1 U5080 ( .A(n4629), .ZN(n4628) );
  NAND2_X1 U5081 ( .A1(n5390), .A2(n9418), .ZN(n8466) );
  OR2_X1 U5082 ( .A1(n9427), .A2(n9440), .ZN(n8570) );
  NOR2_X1 U5083 ( .A1(n5355), .A2(n9427), .ZN(n4629) );
  OR2_X1 U5084 ( .A1(n5355), .A2(n9419), .ZN(n9414) );
  NAND2_X1 U5085 ( .A1(n5355), .A2(n9419), .ZN(n8567) );
  OR2_X1 U5086 ( .A1(n9667), .A2(n9452), .ZN(n8519) );
  NOR2_X1 U5087 ( .A1(n9502), .A2(n4619), .ZN(n4618) );
  INV_X1 U5088 ( .A(n4620), .ZN(n4619) );
  OR2_X1 U5089 ( .A1(n9502), .A2(n9528), .ZN(n8511) );
  NOR2_X1 U5090 ( .A1(n4551), .A2(n4548), .ZN(n4547) );
  INV_X1 U5091 ( .A(n8514), .ZN(n4548) );
  INV_X1 U5092 ( .A(n9547), .ZN(n4551) );
  INV_X1 U5093 ( .A(n8498), .ZN(n4544) );
  OR2_X1 U5094 ( .A1(n7932), .A2(n7855), .ZN(n8495) );
  NAND2_X1 U5095 ( .A1(n5027), .A2(n8490), .ZN(n4573) );
  NOR2_X1 U5096 ( .A1(n9968), .A2(n7288), .ZN(n4624) );
  INV_X1 U5097 ( .A(n7283), .ZN(n5442) );
  NOR2_X1 U5098 ( .A1(n4849), .A2(n9667), .ZN(n9475) );
  NOR2_X1 U5099 ( .A1(n9533), .A2(n5424), .ZN(n9505) );
  NAND2_X1 U5100 ( .A1(n6010), .A2(n6009), .ZN(n8037) );
  NAND2_X1 U5101 ( .A1(n6006), .A2(n6005), .ZN(n6010) );
  AND2_X1 U5102 ( .A1(n4858), .A2(n4857), .ZN(n4561) );
  NOR2_X1 U5103 ( .A1(n5290), .A2(n4701), .ZN(n4700) );
  INV_X1 U5104 ( .A(n5275), .ZN(n4701) );
  OAI21_X1 U5105 ( .B1(n5256), .B2(n5257), .A(n5258), .ZN(n5274) );
  NOR2_X1 U5106 ( .A1(n5152), .A2(n4694), .ZN(n4693) );
  INV_X1 U5107 ( .A(n5134), .ZN(n4694) );
  INV_X1 U5108 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4560) );
  INV_X1 U5109 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4559) );
  AOI21_X1 U5110 ( .B1(n4324), .B2(n4681), .A(n4367), .ZN(n4676) );
  NAND2_X1 U5111 ( .A1(n5031), .A2(n4471), .ZN(n4469) );
  AND2_X1 U5112 ( .A1(n5073), .A2(n5059), .ZN(n5071) );
  NAND2_X1 U5113 ( .A1(n4470), .A2(n4467), .ZN(n5055) );
  INV_X1 U5114 ( .A(n4473), .ZN(n4467) );
  NAND2_X1 U5115 ( .A1(n5029), .A2(n5012), .ZN(n5030) );
  OAI21_X1 U5116 ( .B1(n4928), .B2(n4442), .A(n4441), .ZN(n4925) );
  INV_X1 U5117 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4442) );
  NAND2_X1 U5118 ( .A1(n4928), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4441) );
  NOR2_X1 U5119 ( .A1(n7205), .A2(n4783), .ZN(n4782) );
  INV_X1 U5120 ( .A(n4787), .ZN(n4783) );
  NAND2_X1 U5121 ( .A1(n8776), .A2(n8610), .ZN(n8616) );
  INV_X1 U5122 ( .A(n6805), .ZN(n4768) );
  NOR2_X1 U5123 ( .A1(n4760), .A2(n8634), .ZN(n4752) );
  AND2_X1 U5124 ( .A1(n8758), .A2(n4749), .ZN(n4744) );
  NOR2_X1 U5125 ( .A1(n8634), .A2(n4754), .ZN(n4753) );
  INV_X1 U5126 ( .A(n4759), .ZN(n4754) );
  NOR2_X1 U5127 ( .A1(n4359), .A2(n4748), .ZN(n4747) );
  AND2_X1 U5128 ( .A1(n8758), .A2(n4749), .ZN(n4748) );
  INV_X1 U5129 ( .A(n8634), .ZN(n4756) );
  OR2_X1 U5130 ( .A1(n6683), .A2(n6682), .ZN(n4765) );
  NAND2_X1 U5131 ( .A1(n8612), .A2(n8611), .ZN(n8615) );
  NAND2_X1 U5132 ( .A1(n8768), .A2(n8988), .ZN(n8612) );
  OR2_X1 U5133 ( .A1(n8616), .A2(n4846), .ZN(n8765) );
  XOR2_X1 U5134 ( .A(n8631), .B(n9149), .Z(n8768) );
  NAND2_X1 U5135 ( .A1(n6670), .A2(n6671), .ZN(n10010) );
  AND2_X1 U5136 ( .A1(n8243), .A2(n8242), .ZN(n4535) );
  NAND2_X1 U5137 ( .A1(n6362), .A2(n6259), .ZN(n8851) );
  NOR2_X1 U5138 ( .A1(n8285), .A2(n8284), .ZN(n8283) );
  OR2_X1 U5139 ( .A1(n8274), .A2(n8273), .ZN(n4393) );
  NOR2_X1 U5140 ( .A1(n6550), .A2(n6549), .ZN(n6598) );
  NAND2_X1 U5141 ( .A1(n6938), .A2(n6939), .ZN(n7266) );
  NAND2_X1 U5142 ( .A1(n5560), .A2(n5561), .ZN(n5778) );
  NAND2_X1 U5143 ( .A1(n6028), .A2(n4807), .ZN(n4806) );
  INV_X1 U5144 ( .A(n5879), .ZN(n4807) );
  NOR2_X1 U5145 ( .A1(n8189), .A2(n8186), .ZN(n8205) );
  NOR2_X1 U5146 ( .A1(n4589), .A2(n4587), .ZN(n4586) );
  NAND2_X1 U5147 ( .A1(n8964), .A2(n8175), .ZN(n4587) );
  AOI21_X1 U5148 ( .B1(n4801), .B2(n9026), .A(n4336), .ZN(n4799) );
  INV_X1 U5149 ( .A(n4801), .ZN(n4800) );
  AND2_X1 U5150 ( .A1(n8172), .A2(n8173), .ZN(n9005) );
  NAND2_X1 U5151 ( .A1(n9154), .A2(n9009), .ZN(n9006) );
  NOR2_X1 U5152 ( .A1(n9154), .A2(n9043), .ZN(n9019) );
  NAND2_X1 U5153 ( .A1(n9018), .A2(n9017), .ZN(n9016) );
  AND2_X1 U5154 ( .A1(n9036), .A2(n9037), .ZN(n5967) );
  INV_X1 U5155 ( .A(n4820), .ZN(n9033) );
  NAND2_X1 U5156 ( .A1(n4824), .A2(n4826), .ZN(n4821) );
  OR2_X1 U5157 ( .A1(n9171), .A2(n8752), .ZN(n9059) );
  OR2_X1 U5158 ( .A1(n9086), .A2(n8752), .ZN(n4837) );
  AND2_X1 U5159 ( .A1(n8166), .A2(n9037), .ZN(n9060) );
  OR2_X1 U5160 ( .A1(n9188), .A2(n9119), .ZN(n5789) );
  NAND2_X1 U5161 ( .A1(n8147), .A2(n8151), .ZN(n4609) );
  INV_X1 U5162 ( .A(n4812), .ZN(n4811) );
  OAI21_X1 U5163 ( .B1(n8223), .B2(n4816), .A(n4815), .ZN(n4812) );
  NOR2_X1 U5164 ( .A1(n7890), .A2(n4814), .ZN(n7889) );
  NAND2_X1 U5165 ( .A1(n9808), .A2(n7891), .ZN(n4816) );
  OR2_X1 U5166 ( .A1(n9816), .A2(n7720), .ZN(n4834) );
  OR2_X1 U5167 ( .A1(n7716), .A2(n8224), .ZN(n4817) );
  AND2_X1 U5168 ( .A1(n8118), .A2(n8116), .ZN(n8216) );
  NOR2_X1 U5169 ( .A1(n4505), .A2(n7011), .ZN(n7137) );
  OR2_X1 U5170 ( .A1(n6684), .A2(n7013), .ZN(n4505) );
  OAI22_X1 U5171 ( .A1(n6896), .A2(n5664), .B1(n6902), .B2(n8828), .ZN(n7010)
         );
  INV_X1 U5172 ( .A(n8936), .ZN(n6039) );
  NAND2_X1 U5173 ( .A1(n8640), .A2(n10142), .ZN(n6038) );
  AOI21_X1 U5174 ( .B1(n5540), .B2(n4819), .A(n5541), .ZN(n4818) );
  NOR2_X1 U5175 ( .A1(n5542), .A2(n5765), .ZN(n4819) );
  NOR2_X1 U5176 ( .A1(n4334), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n4528) );
  AND2_X1 U5177 ( .A1(n5715), .A2(n5705), .ZN(n6547) );
  NAND2_X1 U5178 ( .A1(n7078), .A2(n7079), .ZN(n4655) );
  NOR2_X1 U5179 ( .A1(n4832), .A2(n9243), .ZN(n4660) );
  INV_X1 U5180 ( .A(n4832), .ZN(n4659) );
  INV_X1 U5181 ( .A(n4655), .ZN(n4650) );
  INV_X1 U5182 ( .A(n4652), .ZN(n4651) );
  OAI21_X1 U5183 ( .B1(n4656), .B2(n4653), .A(n7238), .ZN(n4652) );
  INV_X1 U5184 ( .A(n4649), .ZN(n4648) );
  OAI21_X1 U5185 ( .B1(n4656), .B2(n4650), .A(n7239), .ZN(n4649) );
  AND2_X1 U5186 ( .A1(n6625), .A2(n6355), .ZN(n6825) );
  AOI21_X1 U5187 ( .B1(n4669), .B2(n4327), .A(n4361), .ZN(n4667) );
  XNOR2_X1 U5188 ( .A(n8709), .B(n8721), .ZN(n8712) );
  NOR2_X1 U5189 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4876) );
  NAND2_X1 U5190 ( .A1(n8537), .A2(n6837), .ZN(n4450) );
  NOR2_X1 U5191 ( .A1(n9896), .A2(n4380), .ZN(n6243) );
  OR2_X1 U5192 ( .A1(n6243), .A2(n6242), .ZN(n4411) );
  NOR2_X1 U5193 ( .A1(n8452), .A2(n6013), .ZN(n9380) );
  AND2_X1 U5194 ( .A1(n5429), .A2(n8453), .ZN(n4579) );
  OAI22_X1 U5195 ( .A1(n4577), .A2(n4580), .B1(n4582), .B2(n8453), .ZN(n4576)
         );
  NOR2_X1 U5196 ( .A1(n5429), .A2(n8453), .ZN(n4580) );
  INV_X1 U5197 ( .A(n8453), .ZN(n4581) );
  OR2_X1 U5198 ( .A1(n5390), .A2(n9418), .ZN(n8526) );
  INV_X1 U5199 ( .A(n4708), .ZN(n4707) );
  AOI21_X1 U5200 ( .B1(n4708), .B2(n4706), .A(n4362), .ZN(n4705) );
  INV_X1 U5201 ( .A(n5335), .ZN(n4706) );
  OAI21_X1 U5202 ( .B1(n9468), .B2(n5319), .A(n5318), .ZN(n9450) );
  AOI21_X1 U5203 ( .B1(n4326), .B2(n4714), .A(n4357), .ZN(n4713) );
  INV_X1 U5204 ( .A(n5271), .ZN(n4714) );
  INV_X1 U5205 ( .A(n4326), .ZN(n4715) );
  NAND2_X1 U5206 ( .A1(n5255), .A2(n5254), .ZN(n9521) );
  AND4_X1 U5207 ( .A1(n5192), .A2(n5191), .A3(n5190), .A4(n5189), .ZN(n9586)
         );
  AOI21_X1 U5208 ( .B1(n5131), .B2(n4729), .A(n4382), .ZN(n4728) );
  INV_X1 U5209 ( .A(n5110), .ZN(n4729) );
  INV_X1 U5210 ( .A(n5131), .ZN(n4730) );
  AND4_X1 U5211 ( .A1(n4993), .A2(n4992), .A3(n4991), .A4(n4990), .ZN(n7292)
         );
  AND2_X1 U5212 ( .A1(n8490), .A2(n8319), .ZN(n8436) );
  OAI21_X1 U5213 ( .B1(n7105), .B2(n7107), .A(n8435), .ZN(n7169) );
  NOR2_X1 U5214 ( .A1(n8429), .A2(n4721), .ZN(n4720) );
  INV_X1 U5215 ( .A(n4950), .ZN(n4721) );
  NAND2_X1 U5216 ( .A1(n4719), .A2(n4718), .ZN(n7281) );
  NOR2_X1 U5217 ( .A1(n4845), .A2(n8309), .ZN(n4718) );
  NAND2_X1 U5218 ( .A1(n8399), .A2(n8398), .ZN(n8413) );
  INV_X1 U5219 ( .A(n9454), .ZN(n9660) );
  OR2_X1 U5220 ( .A1(n8415), .A2(n6837), .ZN(n9787) );
  NAND2_X1 U5221 ( .A1(n4930), .A2(n4434), .ZN(n7124) );
  INV_X1 U5222 ( .A(n4435), .ZN(n4434) );
  OAI22_X1 U5223 ( .A1(n8397), .A2(n6077), .B1(n4999), .B2(n6173), .ZN(n4435)
         );
  AND4_X1 U5224 ( .A1(n4940), .A2(n4939), .A3(n4938), .A4(n4937), .ZN(n6855)
         );
  NAND2_X1 U5225 ( .A1(n4873), .A2(n4862), .ZN(n4736) );
  NAND2_X1 U5226 ( .A1(n5375), .A2(n5374), .ZN(n5392) );
  XNOR2_X1 U5227 ( .A(n5373), .B(n5372), .ZN(n7901) );
  OAI21_X1 U5228 ( .B1(n5276), .B2(n4698), .A(n4696), .ZN(n5321) );
  INV_X1 U5229 ( .A(n4697), .ZN(n4696) );
  OAI21_X1 U5230 ( .B1(n4700), .B2(n4698), .A(n5302), .ZN(n4697) );
  NAND2_X1 U5231 ( .A1(n4699), .A2(n5289), .ZN(n4698) );
  NAND2_X1 U5232 ( .A1(n5404), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5408) );
  NAND2_X1 U5233 ( .A1(n4481), .A2(n5195), .ZN(n5214) );
  NAND2_X1 U5234 ( .A1(n4448), .A2(n4981), .ZN(n4996) );
  NAND2_X1 U5235 ( .A1(n4979), .A2(n4978), .ZN(n4448) );
  NAND2_X1 U5236 ( .A1(n4416), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4921) );
  INV_X1 U5237 ( .A(n4905), .ZN(n4416) );
  AOI21_X1 U5238 ( .B1(n8803), .B2(n8802), .A(n8626), .ZN(n8735) );
  XNOR2_X1 U5239 ( .A(n8616), .B(n4846), .ZN(n8742) );
  OAI22_X1 U5240 ( .A1(n6562), .A2(n6561), .B1(n6560), .B2(n6559), .ZN(n6708)
         );
  NAND2_X1 U5241 ( .A1(n4772), .A2(n4771), .ZN(n7984) );
  AOI21_X1 U5242 ( .B1(n4774), .B2(n4776), .A(n4379), .ZN(n4771) );
  NOR2_X1 U5243 ( .A1(n4757), .A2(n4745), .ZN(n4742) );
  AND2_X1 U5244 ( .A1(n6667), .A2(n6666), .ZN(n10015) );
  INV_X1 U5245 ( .A(n6663), .ZN(n6664) );
  NAND2_X1 U5246 ( .A1(n4533), .A2(n4532), .ZN(n4531) );
  OAI21_X1 U5247 ( .B1(n8241), .B2(n4535), .A(n4534), .ZN(n4533) );
  NAND2_X1 U5248 ( .A1(n4594), .A2(n4390), .ZN(n4532) );
  NAND2_X1 U5249 ( .A1(n8245), .A2(n8244), .ZN(n4534) );
  OR2_X1 U5250 ( .A1(n8635), .A2(n5911), .ZN(n5891) );
  NAND2_X1 U5251 ( .A1(n8049), .A2(n8048), .ZN(n9795) );
  NAND2_X1 U5252 ( .A1(n6029), .A2(n6028), .ZN(n6027) );
  NAND2_X1 U5253 ( .A1(n4638), .A2(n6621), .ZN(n4635) );
  NAND2_X1 U5254 ( .A1(n5218), .A2(n5217), .ZN(n9566) );
  NAND2_X1 U5255 ( .A1(n5162), .A2(n5161), .ZN(n9624) );
  NAND2_X1 U5256 ( .A1(n4643), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4642) );
  INV_X1 U5257 ( .A(n7293), .ZN(n9326) );
  OR2_X1 U5258 ( .A1(n4932), .A2(n4890), .ZN(n4891) );
  NAND2_X1 U5259 ( .A1(n4933), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4892) );
  NAND2_X1 U5260 ( .A1(n5042), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n4894) );
  OAI21_X1 U5261 ( .B1(n6150), .B2(P1_REG2_REG_1__SCAN_IN), .A(n4412), .ZN(
        n6188) );
  NAND2_X1 U5262 ( .A1(n6150), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4412) );
  AND2_X1 U5263 ( .A1(n5986), .A2(n5403), .ZN(n9391) );
  OR2_X1 U5264 ( .A1(n4932), .A2(n4865), .ZN(n4871) );
  AND2_X1 U5265 ( .A1(n9389), .A2(n9382), .ZN(n6024) );
  AOI21_X1 U5266 ( .B1(n8020), .B2(n9992), .A(n6003), .ZN(n6055) );
  NAND2_X1 U5267 ( .A1(n5880), .A2(n4998), .ZN(n5396) );
  NOR2_X1 U5268 ( .A1(n5505), .A2(n9406), .ZN(n9638) );
  NAND2_X1 U5269 ( .A1(n5495), .A2(n5494), .ZN(n5505) );
  INV_X1 U5270 ( .A(n9409), .ZN(n5494) );
  OAI21_X1 U5271 ( .B1(n8102), .B2(n8081), .A(n4536), .ZN(n8082) );
  NOR2_X1 U5272 ( .A1(n4538), .A2(n4537), .ZN(n4536) );
  AND2_X1 U5273 ( .A1(n8154), .A2(n8152), .ZN(n4518) );
  NAND2_X1 U5274 ( .A1(n4425), .A2(n8350), .ZN(n8353) );
  NAND2_X1 U5275 ( .A1(n4429), .A2(n4426), .ZN(n4425) );
  NOR2_X1 U5276 ( .A1(n4428), .A2(n4427), .ZN(n4426) );
  OAI211_X1 U5277 ( .C1(n8153), .C2(n4370), .A(n4335), .B(n4322), .ZN(n4520)
         );
  AND2_X1 U5278 ( .A1(n8166), .A2(n9059), .ZN(n4519) );
  NOR2_X1 U5279 ( .A1(n8424), .A2(n4461), .ZN(n4460) );
  NAND2_X1 U5280 ( .A1(n4685), .A2(n4686), .ZN(n4524) );
  AOI21_X1 U5281 ( .B1(n8063), .B2(n8201), .A(n4687), .ZN(n4686) );
  NAND2_X1 U5282 ( .A1(n8064), .A2(n8198), .ZN(n4685) );
  OAI21_X1 U5283 ( .B1(n8175), .B2(n8201), .A(n8182), .ZN(n4684) );
  NAND2_X1 U5284 ( .A1(n4682), .A2(n8177), .ZN(n8180) );
  INV_X1 U5285 ( .A(n8377), .ZN(n4484) );
  OAI211_X1 U5286 ( .C1(n8369), .C2(n8415), .A(n4483), .B(n8371), .ZN(n4482)
         );
  NOR2_X1 U5287 ( .A1(n8236), .A2(n8201), .ZN(n4675) );
  OR2_X1 U5288 ( .A1(n9795), .A2(n8051), .ZN(n8200) );
  NAND2_X1 U5289 ( .A1(n8391), .A2(n8392), .ZN(n4439) );
  INV_X1 U5290 ( .A(n5195), .ZN(n4480) );
  INV_X1 U5291 ( .A(n5193), .ZN(n4477) );
  INV_X1 U5292 ( .A(n5172), .ZN(n4692) );
  AND2_X1 U5293 ( .A1(n4324), .A2(n4465), .ZN(n4471) );
  NAND2_X1 U5294 ( .A1(n5093), .A2(n7578), .ZN(n5111) );
  NAND2_X1 U5295 ( .A1(n4475), .A2(n5052), .ZN(n4473) );
  INV_X1 U5296 ( .A(n4760), .ZN(n4755) );
  NAND2_X1 U5297 ( .A1(n4789), .A2(n4788), .ZN(n8607) );
  AOI21_X1 U5298 ( .B1(n4791), .B2(n4793), .A(n4349), .ZN(n4788) );
  AND4_X1 U5299 ( .A1(n4509), .A2(n4508), .A3(n4512), .A4(n4507), .ZN(n8240)
         );
  NAND2_X1 U5300 ( .A1(n4346), .A2(n4513), .ZN(n4508) );
  INV_X1 U5301 ( .A(n8204), .ZN(n4512) );
  OR2_X1 U5302 ( .A1(n8640), .A2(n5892), .ZN(n8059) );
  AND2_X1 U5303 ( .A1(n8986), .A2(n5968), .ZN(n4592) );
  AND2_X1 U5304 ( .A1(n9005), .A2(n9006), .ZN(n5968) );
  AND2_X1 U5305 ( .A1(n5824), .A2(n9080), .ZN(n4824) );
  NAND2_X1 U5306 ( .A1(n5824), .A2(n4823), .ZN(n4822) );
  INV_X1 U5307 ( .A(n4837), .ZN(n4823) );
  AND2_X1 U5308 ( .A1(n9177), .A2(n9120), .ZN(n5802) );
  NAND2_X1 U5309 ( .A1(n5535), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5796) );
  INV_X1 U5310 ( .A(n5784), .ZN(n5535) );
  OR2_X1 U5311 ( .A1(n5771), .A2(n7566), .ZN(n5784) );
  NAND2_X1 U5312 ( .A1(n5534), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5771) );
  INV_X1 U5313 ( .A(n5759), .ZN(n5534) );
  NOR2_X1 U5314 ( .A1(n7895), .A2(n4498), .ZN(n4497) );
  INV_X1 U5315 ( .A(n4499), .ZN(n4498) );
  OR2_X1 U5316 ( .A1(n5708), .A2(n8271), .ZN(n5720) );
  OR2_X1 U5317 ( .A1(n10132), .A2(n5714), .ZN(n8119) );
  INV_X1 U5318 ( .A(n8113), .ZN(n4600) );
  INV_X1 U5319 ( .A(n4601), .ZN(n4598) );
  NOR2_X1 U5320 ( .A1(n6684), .A2(n4502), .ZN(n4501) );
  NAND2_X1 U5321 ( .A1(n10125), .A2(n4503), .ZN(n4502) );
  INV_X1 U5322 ( .A(n7011), .ZN(n4504) );
  NAND2_X1 U5323 ( .A1(n5531), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5708) );
  INV_X1 U5324 ( .A(n5695), .ZN(n5531) );
  NAND2_X1 U5325 ( .A1(n6962), .A2(n6736), .ZN(n8080) );
  OR2_X1 U5326 ( .A1(n10057), .A2(n10056), .ZN(n10058) );
  INV_X1 U5327 ( .A(n4827), .ZN(n4611) );
  OR2_X1 U5328 ( .A1(n5654), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U5329 ( .A1(n7613), .A2(n4880), .ZN(n4674) );
  INV_X1 U5330 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4880) );
  INV_X1 U5331 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4881) );
  NAND2_X1 U5332 ( .A1(n6868), .A2(n4333), .ZN(n4639) );
  OR2_X1 U5333 ( .A1(n8452), .A2(n8451), .ZN(n8456) );
  NAND2_X1 U5334 ( .A1(n4437), .A2(n4436), .ZN(n8405) );
  NAND2_X1 U5335 ( .A1(n8409), .A2(n8415), .ZN(n4436) );
  OAI21_X1 U5336 ( .B1(n8410), .B2(n8396), .A(n4438), .ZN(n4437) );
  NOR2_X1 U5337 ( .A1(n8409), .A2(n9397), .ZN(n8463) );
  AND2_X1 U5338 ( .A1(n8409), .A2(n9397), .ZN(n8575) );
  OR2_X1 U5339 ( .A1(n9401), .A2(n9228), .ZN(n8461) );
  NAND2_X1 U5340 ( .A1(n9401), .A2(n9228), .ZN(n8467) );
  NOR2_X1 U5341 ( .A1(n4567), .A2(n4565), .ZN(n4564) );
  INV_X1 U5342 ( .A(n8334), .ZN(n4565) );
  INV_X1 U5343 ( .A(n8443), .ZN(n4567) );
  NAND2_X1 U5344 ( .A1(n8443), .A2(n8333), .ZN(n4566) );
  OR2_X1 U5345 ( .A1(n7859), .A2(n4632), .ZN(n4631) );
  OR2_X1 U5346 ( .A1(n7799), .A2(n9845), .ZN(n4632) );
  INV_X1 U5347 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n4969) );
  NOR2_X1 U5348 ( .A1(n9401), .A2(n4626), .ZN(n4625) );
  INV_X1 U5349 ( .A(n4627), .ZN(n4626) );
  NAND2_X1 U5350 ( .A1(n9503), .A2(n5425), .ZN(n9507) );
  NAND2_X1 U5351 ( .A1(n5901), .A2(n5900), .ZN(n6006) );
  NAND2_X1 U5352 ( .A1(n5896), .A2(n5895), .ZN(n5901) );
  OAI21_X1 U5353 ( .B1(n5341), .B2(n5340), .A(n5339), .ZN(n5358) );
  INV_X1 U5354 ( .A(n5303), .ZN(n4699) );
  NAND2_X1 U5355 ( .A1(n5236), .A2(n5235), .ZN(n5256) );
  AOI21_X1 U5356 ( .B1(n5071), .B2(n4680), .A(n4679), .ZN(n4678) );
  INV_X1 U5357 ( .A(n5073), .ZN(n4679) );
  INV_X1 U5358 ( .A(n5054), .ZN(n4680) );
  INV_X1 U5359 ( .A(n5071), .ZN(n4681) );
  XNOR2_X1 U5360 ( .A(n5007), .B(SI_7_), .ZN(n5004) );
  AOI21_X1 U5361 ( .B1(n4995), .B2(n4447), .A(n4360), .ZN(n4446) );
  NAND2_X1 U5362 ( .A1(n4763), .A2(n6666), .ZN(n6699) );
  OR2_X1 U5363 ( .A1(n7201), .A2(n7200), .ZN(n4787) );
  NAND2_X1 U5364 ( .A1(n4786), .A2(n4785), .ZN(n4784) );
  INV_X1 U5365 ( .A(n7203), .ZN(n4786) );
  OR2_X1 U5366 ( .A1(n5796), .A2(n5795), .ZN(n5798) );
  NAND2_X1 U5367 ( .A1(n5536), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5806) );
  INV_X1 U5368 ( .A(n5798), .ZN(n5536) );
  INV_X1 U5369 ( .A(n4778), .ZN(n4776) );
  OR2_X1 U5370 ( .A1(n5681), .A2(n8878), .ZN(n5695) );
  OR2_X1 U5371 ( .A1(n5806), .A2(n8004), .ZN(n5816) );
  NOR2_X1 U5372 ( .A1(n8601), .A2(n4795), .ZN(n4794) );
  INV_X1 U5373 ( .A(n8002), .ZN(n4795) );
  NAND2_X1 U5374 ( .A1(n5532), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5730) );
  INV_X1 U5375 ( .A(n5720), .ZN(n5532) );
  OR2_X1 U5376 ( .A1(n5730), .A2(n7059), .ZN(n5745) );
  AND2_X1 U5377 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5636) );
  NAND2_X1 U5378 ( .A1(n6806), .A2(n6805), .ZN(n4769) );
  INV_X1 U5379 ( .A(n7732), .ZN(n4777) );
  OR2_X1 U5380 ( .A1(n7803), .A2(n7802), .ZN(n4778) );
  NAND2_X1 U5381 ( .A1(n4779), .A2(n4780), .ZN(n7701) );
  AOI21_X1 U5382 ( .B1(n4782), .B2(n7202), .A(n4781), .ZN(n4780) );
  INV_X1 U5383 ( .A(n7377), .ZN(n4781) );
  NAND2_X1 U5384 ( .A1(n6363), .A2(n6364), .ZN(n6362) );
  NAND2_X1 U5385 ( .A1(n8852), .A2(n8851), .ZN(n8850) );
  NAND2_X1 U5386 ( .A1(n6516), .A2(n6517), .ZN(n6515) );
  NOR2_X1 U5387 ( .A1(n6540), .A2(n4396), .ZN(n8880) );
  AND2_X1 U5388 ( .A1(n6541), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4396) );
  OR2_X1 U5389 ( .A1(n8880), .A2(n8881), .ZN(n4395) );
  AND2_X1 U5390 ( .A1(n4395), .A2(n4394), .ZN(n8285) );
  NAND2_X1 U5391 ( .A1(n8874), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4394) );
  AND2_X1 U5392 ( .A1(n6606), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4391) );
  NAND2_X1 U5393 ( .A1(n6776), .A2(n4398), .ZN(n6778) );
  OR2_X1 U5394 ( .A1(n6777), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4398) );
  NAND2_X1 U5395 ( .A1(n6778), .A2(n6779), .ZN(n6936) );
  NAND2_X1 U5396 ( .A1(n6936), .A2(n4397), .ZN(n6938) );
  OR2_X1 U5397 ( .A1(n6937), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4397) );
  NOR2_X1 U5398 ( .A1(n7874), .A2(n7875), .ZN(n8890) );
  NAND2_X1 U5399 ( .A1(n8890), .A2(n8889), .ZN(n8888) );
  NAND2_X1 U5400 ( .A1(n8888), .A2(n4400), .ZN(n8265) );
  OR2_X1 U5401 ( .A1(n8895), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4400) );
  NOR2_X1 U5402 ( .A1(n8265), .A2(n8264), .ZN(n8263) );
  NAND2_X1 U5403 ( .A1(n8990), .A2(n4487), .ZN(n6035) );
  AND2_X1 U5404 ( .A1(n8990), .A2(n4337), .ZN(n8930) );
  INV_X1 U5405 ( .A(n8945), .ZN(n8949) );
  INV_X1 U5406 ( .A(n5861), .ZN(n5860) );
  OR2_X1 U5407 ( .A1(n9146), .A2(n8965), .ZN(n5857) );
  NOR2_X1 U5408 ( .A1(n9146), .A2(n8999), .ZN(n8990) );
  NAND2_X1 U5409 ( .A1(n8990), .A2(n5868), .ZN(n8971) );
  INV_X1 U5410 ( .A(n8172), .ZN(n4591) );
  INV_X1 U5411 ( .A(n4588), .ZN(n4585) );
  OR2_X1 U5412 ( .A1(n9149), .A2(n8988), .ZN(n8172) );
  OR2_X1 U5413 ( .A1(n9161), .A2(n8751), .ZN(n9024) );
  NAND2_X1 U5414 ( .A1(n9110), .A2(n4330), .ZN(n9043) );
  NAND2_X1 U5415 ( .A1(n5537), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5827) );
  INV_X1 U5416 ( .A(n5816), .ZN(n5537) );
  OR2_X1 U5417 ( .A1(n5827), .A2(n8780), .ZN(n5829) );
  INV_X1 U5418 ( .A(n5966), .ZN(n9036) );
  NAND2_X1 U5419 ( .A1(n9110), .A2(n4491), .ZN(n9052) );
  AND2_X1 U5420 ( .A1(n9069), .A2(n9070), .ZN(n5965) );
  NAND2_X1 U5421 ( .A1(n9110), .A2(n9099), .ZN(n9093) );
  NAND2_X1 U5422 ( .A1(n4604), .A2(n4602), .ZN(n9117) );
  AND2_X1 U5423 ( .A1(n4606), .A2(n4603), .ZN(n4602) );
  NAND2_X1 U5424 ( .A1(n4345), .A2(n4814), .ZN(n4603) );
  AND2_X1 U5425 ( .A1(n9109), .A2(n9115), .ZN(n9110) );
  AND2_X1 U5426 ( .A1(n8159), .A2(n8156), .ZN(n9118) );
  AND2_X1 U5427 ( .A1(n7964), .A2(n7963), .ZN(n9109) );
  AND2_X1 U5428 ( .A1(n9191), .A2(n8818), .ZN(n5777) );
  AND2_X1 U5429 ( .A1(n7627), .A2(n4495), .ZN(n7964) );
  AND2_X1 U5430 ( .A1(n4497), .A2(n4496), .ZN(n4495) );
  NAND2_X1 U5431 ( .A1(n7627), .A2(n4497), .ZN(n7910) );
  NAND2_X1 U5432 ( .A1(n5533), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5759) );
  INV_X1 U5433 ( .A(n5747), .ZN(n5533) );
  NAND2_X1 U5434 ( .A1(n7627), .A2(n9816), .ZN(n7723) );
  AND2_X1 U5435 ( .A1(n7328), .A2(n10151), .ZN(n7627) );
  NAND2_X1 U5436 ( .A1(n8134), .A2(n8132), .ZN(n8220) );
  NOR2_X1 U5437 ( .A1(n7254), .A2(n10141), .ZN(n7328) );
  NAND2_X1 U5438 ( .A1(n8130), .A2(n8070), .ZN(n8219) );
  AND2_X1 U5439 ( .A1(n7186), .A2(n8217), .ZN(n7249) );
  AOI21_X1 U5440 ( .B1(n4597), .B2(n4596), .A(n4595), .ZN(n7186) );
  INV_X1 U5441 ( .A(n4599), .ZN(n4595) );
  AND2_X1 U5442 ( .A1(n4598), .A2(n8216), .ZN(n4596) );
  AOI21_X1 U5443 ( .B1(n8216), .B2(n4600), .A(n5962), .ZN(n4599) );
  NAND2_X1 U5444 ( .A1(n4504), .A2(n4501), .ZN(n7190) );
  AND2_X1 U5445 ( .A1(n5688), .A2(n5676), .ZN(n4829) );
  INV_X1 U5446 ( .A(n8215), .ZN(n5688) );
  NOR2_X1 U5447 ( .A1(n7015), .A2(n5961), .ZN(n6984) );
  AND2_X1 U5448 ( .A1(n5636), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U5449 ( .A1(n5656), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5670) );
  OAI21_X1 U5450 ( .B1(n6959), .B2(n8208), .A(n8098), .ZN(n6732) );
  AND2_X1 U5451 ( .A1(n8080), .A2(n8100), .ZN(n6731) );
  NAND2_X1 U5452 ( .A1(n6946), .A2(n10086), .ZN(n10057) );
  NOR2_X1 U5453 ( .A1(n6910), .A2(n6919), .ZN(n6946) );
  INV_X1 U5454 ( .A(n6384), .ZN(n6914) );
  NAND2_X1 U5455 ( .A1(n8031), .A2(n8030), .ZN(n9800) );
  AND2_X1 U5456 ( .A1(n4614), .A2(n4613), .ZN(n4612) );
  AND2_X1 U5457 ( .A1(n5917), .A2(n5542), .ZN(n4613) );
  AND2_X1 U5458 ( .A1(n4839), .A2(n5917), .ZN(n4615) );
  NAND2_X1 U5459 ( .A1(n4525), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5943) );
  AND2_X1 U5460 ( .A1(n4528), .A2(n4527), .ZN(n4526) );
  NAND2_X1 U5461 ( .A1(n5920), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5947) );
  NAND2_X1 U5462 ( .A1(n5780), .A2(n5562), .ZN(n5920) );
  OR3_X1 U5463 ( .A1(n5702), .A2(P2_IR_REG_10__SCAN_IN), .A3(
        P2_IR_REG_11__SCAN_IN), .ZN(n5726) );
  OR2_X1 U5464 ( .A1(n5665), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5677) );
  NOR2_X1 U5465 ( .A1(n4641), .A2(n4639), .ZN(n4638) );
  INV_X1 U5466 ( .A(n5311), .ZN(n5312) );
  INV_X1 U5467 ( .A(n5247), .ZN(n5248) );
  NAND2_X1 U5468 ( .A1(n5248), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5265) );
  OR2_X1 U5469 ( .A1(n7078), .A2(n7079), .ZN(n4656) );
  NAND2_X1 U5470 ( .A1(n6422), .A2(n6421), .ZN(n6430) );
  OAI21_X1 U5471 ( .B1(n6621), .B2(n4637), .A(n4636), .ZN(n6997) );
  AOI21_X1 U5472 ( .B1(n6755), .B2(n4641), .A(n4640), .ZN(n4636) );
  INV_X1 U5473 ( .A(n6755), .ZN(n4637) );
  OAI22_X1 U5474 ( .A1(n6855), .A2(n6498), .B1(n6798), .B2(n8718), .ZN(n6751)
         );
  INV_X1 U5475 ( .A(n5265), .ZN(n5266) );
  NOR2_X1 U5476 ( .A1(n5280), .A2(n9252), .ZN(n5297) );
  NOR2_X1 U5477 ( .A1(n8591), .A2(n8586), .ZN(n6320) );
  NOR2_X1 U5478 ( .A1(n5365), .A2(n5364), .ZN(n5384) );
  INV_X1 U5479 ( .A(n8420), .ZN(n8406) );
  NAND2_X1 U5480 ( .A1(n8591), .A2(n9408), .ZN(n6419) );
  AND4_X1 U5481 ( .A1(n5109), .A2(n5108), .A3(n5107), .A4(n5106), .ZN(n7688)
         );
  AND4_X1 U5482 ( .A1(n5069), .A2(n5068), .A3(n5067), .A4(n5066), .ZN(n7339)
         );
  OR2_X1 U5483 ( .A1(n4989), .A2(n6123), .ZN(n4893) );
  NAND2_X1 U5484 ( .A1(n5461), .A2(n5455), .ZN(n6624) );
  AND2_X1 U5485 ( .A1(n6177), .A2(n6137), .ZN(n6331) );
  OR2_X1 U5486 ( .A1(n6207), .A2(n6206), .ZN(n6220) );
  AND2_X1 U5487 ( .A1(n4411), .A2(n4410), .ZN(n9341) );
  NAND2_X1 U5488 ( .A1(n6450), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4410) );
  NAND2_X1 U5489 ( .A1(n9341), .A2(n9342), .ZN(n9340) );
  OR2_X1 U5490 ( .A1(n7072), .A2(n4418), .ZN(n4417) );
  NOR2_X1 U5491 ( .A1(n4420), .A2(n4419), .ZN(n4418) );
  INV_X1 U5492 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n4419) );
  NOR2_X1 U5493 ( .A1(n9362), .A2(n4404), .ZN(n9908) );
  AND2_X1 U5494 ( .A1(n9367), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4404) );
  NOR2_X1 U5495 ( .A1(n9908), .A2(n9909), .ZN(n9907) );
  AND2_X1 U5496 ( .A1(n8461), .A2(n8467), .ZN(n8395) );
  OR2_X1 U5497 ( .A1(n5402), .A2(n8395), .ZN(n5986) );
  INV_X1 U5498 ( .A(n8395), .ZN(n8450) );
  OR2_X1 U5499 ( .A1(n5496), .A2(n4440), .ZN(n5497) );
  AND4_X1 U5500 ( .A1(n5389), .A2(n5388), .A3(n5387), .A4(n5386), .ZN(n9418)
         );
  AND4_X1 U5501 ( .A1(n5354), .A2(n5353), .A3(n5352), .A4(n5351), .ZN(n9419)
         );
  NAND2_X1 U5502 ( .A1(n9460), .A2(n4629), .ZN(n9425) );
  AND2_X1 U5503 ( .A1(n9475), .A2(n9660), .ZN(n9460) );
  NAND2_X1 U5504 ( .A1(n9460), .A2(n9651), .ZN(n9439) );
  AOI21_X1 U5505 ( .B1(n8518), .B2(n8361), .A(n4555), .ZN(n4554) );
  INV_X1 U5506 ( .A(n8423), .ZN(n4555) );
  OR2_X1 U5507 ( .A1(n9469), .A2(n8422), .ZN(n9470) );
  NAND2_X1 U5508 ( .A1(n9507), .A2(n8364), .ZN(n9484) );
  NAND2_X1 U5509 ( .A1(n9539), .A2(n4331), .ZN(n4849) );
  NAND2_X1 U5510 ( .A1(n9539), .A2(n4618), .ZN(n9511) );
  AOI21_X1 U5511 ( .B1(n9547), .B2(n4550), .A(n4461), .ZN(n4549) );
  INV_X1 U5512 ( .A(n8359), .ZN(n4550) );
  OR2_X1 U5513 ( .A1(n9505), .A2(n8424), .ZN(n9520) );
  AND2_X1 U5514 ( .A1(n5230), .A2(n5229), .ZN(n9536) );
  OR2_X1 U5515 ( .A1(n5187), .A2(n5186), .ZN(n5204) );
  NOR2_X1 U5516 ( .A1(n5204), .A2(n5203), .ZN(n5219) );
  AOI21_X1 U5517 ( .B1(n8501), .B2(n4544), .A(n4543), .ZN(n4542) );
  INV_X1 U5518 ( .A(n8501), .ZN(n4545) );
  INV_X1 U5519 ( .A(n8502), .ZN(n4543) );
  NAND2_X1 U5520 ( .A1(n4724), .A2(n4723), .ZN(n9612) );
  AOI21_X1 U5521 ( .B1(n4725), .B2(n4730), .A(n4384), .ZN(n4723) );
  NOR2_X1 U5522 ( .A1(n9623), .A2(n9624), .ZN(n9621) );
  NAND2_X1 U5523 ( .A1(n5443), .A2(n4630), .ZN(n9623) );
  NOR2_X1 U5524 ( .A1(n4631), .A2(n7932), .ZN(n4630) );
  NAND2_X1 U5525 ( .A1(n4568), .A2(n8338), .ZN(n7848) );
  NAND2_X1 U5526 ( .A1(n7785), .A2(n8334), .ZN(n4568) );
  NAND2_X1 U5527 ( .A1(n7848), .A2(n8443), .ZN(n7926) );
  NOR2_X1 U5528 ( .A1(n7384), .A2(n4632), .ZN(n7856) );
  AND4_X1 U5529 ( .A1(n5086), .A2(n5085), .A3(n5084), .A4(n5083), .ZN(n7794)
         );
  NAND2_X1 U5530 ( .A1(n7169), .A2(n4572), .ZN(n4571) );
  NOR2_X1 U5531 ( .A1(n7384), .A2(n9845), .ZN(n9846) );
  NAND2_X1 U5532 ( .A1(n4733), .A2(n4731), .ZN(n9833) );
  NOR2_X1 U5533 ( .A1(n9835), .A2(n4732), .ZN(n4731) );
  INV_X1 U5534 ( .A(n5070), .ZN(n4732) );
  AND2_X1 U5535 ( .A1(n5064), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5080) );
  NOR2_X1 U5536 ( .A1(n5043), .A2(n7242), .ZN(n5064) );
  NAND2_X1 U5537 ( .A1(n7170), .A2(n8490), .ZN(n7303) );
  AND2_X1 U5538 ( .A1(n5442), .A2(n4375), .ZN(n7305) );
  OR2_X1 U5539 ( .A1(n7169), .A2(n5027), .ZN(n7170) );
  NAND2_X1 U5540 ( .A1(n4541), .A2(n5417), .ZN(n7105) );
  NAND2_X1 U5541 ( .A1(n5442), .A2(n9958), .ZN(n7284) );
  AND2_X1 U5542 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n4951) );
  NAND2_X1 U5543 ( .A1(n4951), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n4970) );
  AND2_X1 U5544 ( .A1(n6789), .A2(n6798), .ZN(n6858) );
  INV_X1 U5545 ( .A(n8430), .ZN(n4433) );
  NAND2_X1 U5546 ( .A1(n6715), .A2(n4433), .ZN(n6714) );
  NOR2_X1 U5547 ( .A1(n6716), .A2(n7124), .ZN(n6789) );
  INV_X1 U5548 ( .A(n6637), .ZN(n4702) );
  NAND2_X1 U5549 ( .A1(n6925), .A2(n4617), .ZN(n6716) );
  AND2_X1 U5550 ( .A1(n9943), .A2(n8427), .ZN(n4617) );
  NAND2_X1 U5551 ( .A1(n6827), .A2(n6829), .ZN(n6828) );
  AND4_X1 U5552 ( .A1(n5026), .A2(n5025), .A3(n5024), .A4(n5023), .ZN(n9963)
         );
  AND4_X1 U5553 ( .A1(n4975), .A2(n4974), .A3(n4973), .A4(n4972), .ZN(n9965)
         );
  AND4_X1 U5554 ( .A1(n4956), .A2(n4955), .A3(n4954), .A4(n4953), .ZN(n7293)
         );
  AND2_X1 U5555 ( .A1(n6825), .A2(n5458), .ZN(n6352) );
  NAND2_X1 U5556 ( .A1(n4860), .A2(n4840), .ZN(n5456) );
  XNOR2_X1 U5557 ( .A(n8046), .B(n8045), .ZN(n9210) );
  XNOR2_X1 U5558 ( .A(n8037), .B(n8036), .ZN(n8732) );
  XNOR2_X1 U5559 ( .A(n6006), .B(n6005), .ZN(n9217) );
  NAND2_X1 U5560 ( .A1(n5394), .A2(n5393), .ZN(n5896) );
  NAND2_X1 U5561 ( .A1(n5392), .A2(n5391), .ZN(n5394) );
  AND3_X1 U5562 ( .A1(n4856), .A2(n4859), .A3(n4561), .ZN(n4840) );
  NAND2_X1 U5563 ( .A1(n4695), .A2(n5289), .ZN(n5304) );
  AND2_X1 U5564 ( .A1(n4671), .A2(n5242), .ZN(n4670) );
  NOR2_X1 U5565 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(n4841), .ZN(n4671) );
  OR2_X1 U5566 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n4841) );
  NAND2_X1 U5567 ( .A1(n5197), .A2(n5196), .ZN(n5240) );
  NAND2_X1 U5568 ( .A1(n4688), .A2(n5151), .ZN(n5173) );
  XNOR2_X1 U5569 ( .A(n5091), .B(n5088), .ZN(n6115) );
  NAND2_X1 U5570 ( .A1(n4677), .A2(n4678), .ZN(n5091) );
  OR2_X1 U5571 ( .A1(n5055), .A2(n4681), .ZN(n4677) );
  NAND2_X1 U5572 ( .A1(n5055), .A2(n5054), .ZN(n5072) );
  OR2_X1 U5573 ( .A1(n5036), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5038) );
  OR2_X1 U5574 ( .A1(n5038), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5075) );
  NAND2_X1 U5575 ( .A1(n4474), .A2(n5029), .ZN(n5053) );
  OR2_X1 U5576 ( .A1(n4959), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5098) );
  XNOR2_X1 U5577 ( .A(n4963), .B(n7511), .ZN(n4961) );
  XNOR2_X1 U5578 ( .A(n4925), .B(n4911), .ZN(n4923) );
  OAI21_X1 U5579 ( .B1(n6066), .B2(n6062), .A(n4885), .ZN(n4906) );
  NAND2_X1 U5580 ( .A1(n6066), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4885) );
  NAND2_X1 U5581 ( .A1(n5871), .A2(n5870), .ZN(n9135) );
  NAND2_X1 U5582 ( .A1(n7940), .A2(n8047), .ZN(n5871) );
  NAND2_X1 U5583 ( .A1(n4784), .A2(n4787), .ZN(n7204) );
  NAND2_X1 U5584 ( .A1(n5578), .A2(n5577), .ZN(n7727) );
  NAND2_X1 U5585 ( .A1(n5529), .A2(n5528), .ZN(n9154) );
  AOI21_X1 U5586 ( .B1(n4373), .B2(n4768), .A(n4767), .ZN(n4766) );
  INV_X1 U5587 ( .A(n7023), .ZN(n4767) );
  AOI22_X1 U5588 ( .A1(n4747), .A2(n4745), .B1(n4758), .B2(n4744), .ZN(n4743)
         );
  NOR2_X1 U5589 ( .A1(n4759), .A2(n4752), .ZN(n4751) );
  INV_X1 U5590 ( .A(n4747), .ZN(n4746) );
  NAND2_X1 U5591 ( .A1(n4790), .A2(n8600), .ZN(n8748) );
  NAND2_X1 U5592 ( .A1(n8003), .A2(n4794), .ZN(n4790) );
  NAND2_X1 U5593 ( .A1(n5729), .A2(n5728), .ZN(n7330) );
  AND2_X1 U5594 ( .A1(n8768), .A2(n8617), .ZN(n8618) );
  NAND2_X1 U5595 ( .A1(n7733), .A2(n7732), .ZN(n7805) );
  NAND2_X1 U5596 ( .A1(n5783), .A2(n5782), .ZN(n9188) );
  INV_X1 U5597 ( .A(n5620), .ZN(n6961) );
  AND2_X1 U5598 ( .A1(n4769), .A2(n4343), .ZN(n6814) );
  NAND2_X1 U5599 ( .A1(n8003), .A2(n8002), .ZN(n8602) );
  NAND2_X1 U5600 ( .A1(n5805), .A2(n5804), .ZN(n9171) );
  NAND2_X1 U5601 ( .A1(n4773), .A2(n4778), .ZN(n7971) );
  NAND2_X1 U5602 ( .A1(n7733), .A2(n4341), .ZN(n4773) );
  NAND2_X1 U5603 ( .A1(n5794), .A2(n5793), .ZN(n9182) );
  INV_X1 U5604 ( .A(n4763), .ZN(n10011) );
  OR2_X1 U5605 ( .A1(n8637), .A2(n9076), .ZN(n8781) );
  INV_X1 U5606 ( .A(n8251), .ZN(n4530) );
  NAND4_X1 U5607 ( .A1(n5663), .A2(n5662), .A3(n5661), .A4(n5660), .ZN(n8828)
         );
  NAND2_X1 U5608 ( .A1(n5872), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5602) );
  NAND2_X1 U5609 ( .A1(n4318), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5601) );
  NOR2_X1 U5610 ( .A1(n6302), .A2(n6301), .ZN(n6300) );
  AND2_X1 U5611 ( .A1(n6515), .A2(n6264), .ZN(n6302) );
  INV_X1 U5612 ( .A(n4395), .ZN(n8883) );
  INV_X1 U5613 ( .A(n4393), .ZN(n8272) );
  INV_X1 U5614 ( .A(n5975), .ZN(n5976) );
  OAI21_X1 U5615 ( .B1(n8944), .B2(n8232), .A(n4805), .ZN(n4808) );
  AND2_X1 U5616 ( .A1(n4806), .A2(n5894), .ZN(n4805) );
  NAND2_X1 U5617 ( .A1(n4796), .A2(n4799), .ZN(n8983) );
  OR2_X1 U5618 ( .A1(n9018), .A2(n4800), .ZN(n4796) );
  NAND2_X1 U5619 ( .A1(n9016), .A2(n4803), .ZN(n8998) );
  NAND2_X1 U5620 ( .A1(n9169), .A2(n4837), .ZN(n9051) );
  NAND2_X1 U5621 ( .A1(n9081), .A2(n9080), .ZN(n9169) );
  OAI21_X1 U5622 ( .B1(n7889), .B2(n4609), .A(n8150), .ZN(n4605) );
  NOR2_X1 U5623 ( .A1(n7889), .A2(n5964), .ZN(n7904) );
  NAND2_X1 U5624 ( .A1(n4810), .A2(n4811), .ZN(n7909) );
  AND2_X1 U5625 ( .A1(n4817), .A2(n4816), .ZN(n7888) );
  NAND2_X1 U5626 ( .A1(n6983), .A2(n8113), .ZN(n7133) );
  NOR2_X1 U5627 ( .A1(n7011), .A2(n7013), .ZN(n6989) );
  OAI211_X1 U5628 ( .C1(n4740), .C2(n4739), .A(n4738), .B(n4737), .ZN(n6902)
         );
  NAND2_X1 U5629 ( .A1(n5630), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n4737) );
  OAI21_X1 U5630 ( .B1(n5576), .B2(n10037), .A(n4485), .ZN(n6919) );
  NAND2_X1 U5631 ( .A1(n5576), .A2(n9222), .ZN(n4485) );
  INV_X1 U5632 ( .A(n10054), .ZN(n8926) );
  AOI211_X1 U5633 ( .C1(n10142), .C2(n9795), .A(n9799), .B(n9794), .ZN(n9823)
         );
  NOR2_X1 U5634 ( .A1(n8941), .A2(n6040), .ZN(n6041) );
  NAND2_X1 U5635 ( .A1(n6039), .A2(n6038), .ZN(n6040) );
  NAND2_X1 U5636 ( .A1(n5780), .A2(n4528), .ZN(n5944) );
  NAND2_X1 U5637 ( .A1(n4401), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5605) );
  INV_X1 U5638 ( .A(n5604), .ZN(n4401) );
  INV_X1 U5639 ( .A(n4668), .ZN(n9226) );
  AOI21_X1 U5640 ( .B1(n4664), .B2(n9259), .A(n8713), .ZN(n4662) );
  INV_X1 U5641 ( .A(n4664), .ZN(n4663) );
  NAND2_X1 U5642 ( .A1(n5310), .A2(n5309), .ZN(n9667) );
  NAND2_X1 U5643 ( .A1(n8661), .A2(n9299), .ZN(n9244) );
  NAND2_X1 U5644 ( .A1(n4647), .A2(n4655), .ZN(n7240) );
  NAND2_X1 U5645 ( .A1(n7080), .A2(n4656), .ZN(n4647) );
  NAND2_X1 U5646 ( .A1(n4659), .A2(n4355), .ZN(n4658) );
  NAND2_X1 U5647 ( .A1(n5184), .A2(n5183), .ZN(n9715) );
  NAND2_X1 U5648 ( .A1(n5202), .A2(n5201), .ZN(n9706) );
  AOI22_X1 U5649 ( .A1(n4651), .A2(n4653), .B1(n4648), .B2(n4650), .ZN(n4644)
         );
  OR2_X1 U5650 ( .A1(n4651), .A2(n4648), .ZN(n4646) );
  CLKBUF_X1 U5651 ( .A(n9310), .Z(n9302) );
  NAND2_X1 U5652 ( .A1(n5363), .A2(n5362), .ZN(n9427) );
  NAND2_X1 U5653 ( .A1(n7901), .A2(n4998), .ZN(n5363) );
  NAND2_X1 U5654 ( .A1(n4666), .A2(n4667), .ZN(n9316) );
  OR2_X1 U5655 ( .A1(n4875), .A2(n4862), .ZN(n4879) );
  NAND2_X1 U5656 ( .A1(n4874), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4875) );
  AOI21_X1 U5657 ( .B1(n4454), .B2(n4451), .A(n4450), .ZN(n4449) );
  NAND2_X1 U5658 ( .A1(n4453), .A2(n9513), .ZN(n4452) );
  NOR2_X1 U5659 ( .A1(n8420), .A2(n4389), .ZN(n4451) );
  INV_X1 U5660 ( .A(n9418), .ZN(n9395) );
  INV_X1 U5661 ( .A(n6855), .ZN(n9327) );
  INV_X1 U5662 ( .A(n7095), .ZN(n9328) );
  NAND2_X1 U5663 ( .A1(n6188), .A2(n6319), .ZN(n6187) );
  INV_X1 U5664 ( .A(n4411), .ZN(n6449) );
  NOR2_X1 U5665 ( .A1(n6654), .A2(n4421), .ZN(n6658) );
  AND2_X1 U5666 ( .A1(n6655), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4421) );
  NOR2_X1 U5667 ( .A1(n6658), .A2(n6657), .ZN(n7072) );
  XNOR2_X1 U5668 ( .A(n4417), .B(n7220), .ZN(n7074) );
  OAI21_X1 U5669 ( .B1(n7216), .B2(n4406), .A(n4405), .ZN(n9354) );
  NAND2_X1 U5670 ( .A1(n4409), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4406) );
  NAND2_X1 U5671 ( .A1(n7664), .A2(n4409), .ZN(n4405) );
  INV_X1 U5672 ( .A(n7666), .ZN(n4409) );
  INV_X1 U5673 ( .A(n7664), .ZN(n4407) );
  XNOR2_X1 U5674 ( .A(n4402), .B(n9541), .ZN(n9374) );
  OR2_X1 U5675 ( .A1(n9907), .A2(n4403), .ZN(n4402) );
  AND2_X1 U5676 ( .A1(n9368), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4403) );
  NOR2_X1 U5677 ( .A1(n9381), .A2(n9622), .ZN(n9635) );
  AOI21_X1 U5678 ( .B1(n5999), .B2(n9693), .A(n5998), .ZN(n8029) );
  AND2_X1 U5679 ( .A1(n6020), .A2(n9322), .ZN(n5998) );
  OAI21_X1 U5680 ( .B1(n9450), .B2(n4707), .A(n4705), .ZN(n9424) );
  OAI21_X1 U5681 ( .B1(n9450), .B2(n4342), .A(n5335), .ZN(n9436) );
  NAND2_X1 U5682 ( .A1(n5325), .A2(n5324), .ZN(n9454) );
  NAND2_X1 U5683 ( .A1(n4712), .A2(n4713), .ZN(n9489) );
  OR2_X1 U5684 ( .A1(n9521), .A2(n4715), .ZN(n4712) );
  NAND2_X1 U5685 ( .A1(n4716), .A2(n5271), .ZN(n9499) );
  OR2_X1 U5686 ( .A1(n9521), .A2(n5272), .ZN(n4716) );
  NAND2_X1 U5687 ( .A1(n5264), .A2(n5263), .ZN(n9533) );
  NAND2_X1 U5688 ( .A1(n4552), .A2(n8359), .ZN(n9548) );
  NAND2_X1 U5689 ( .A1(n9553), .A2(n8514), .ZN(n4552) );
  NAND2_X1 U5690 ( .A1(n9614), .A2(n8498), .ZN(n9591) );
  NAND2_X1 U5691 ( .A1(n4727), .A2(n4728), .ZN(n7930) );
  OR2_X1 U5692 ( .A1(n7788), .A2(n4730), .ZN(n4727) );
  NAND2_X1 U5693 ( .A1(n7788), .A2(n5110), .ZN(n7850) );
  NAND2_X1 U5694 ( .A1(n7106), .A2(n5003), .ZN(n7168) );
  AND2_X1 U5695 ( .A1(n4719), .A2(n4722), .ZN(n7282) );
  NAND2_X1 U5696 ( .A1(n6787), .A2(n4950), .ZN(n6852) );
  OAI21_X1 U5697 ( .B1(n6715), .B2(n4433), .A(n6714), .ZN(n7129) );
  INV_X1 U5698 ( .A(n9589), .ZN(n9595) );
  OR3_X1 U5699 ( .A1(n9787), .A2(n8589), .A3(n5410), .ZN(n9598) );
  INV_X1 U5700 ( .A(n9943), .ZN(n6839) );
  INV_X1 U5701 ( .A(n9628), .ZN(n9844) );
  INV_X1 U5702 ( .A(n8413), .ZN(n9731) );
  AOI211_X1 U5703 ( .C1(n9644), .C2(n9992), .A(n9643), .B(n9642), .ZN(n9732)
         );
  INV_X1 U5704 ( .A(n6494), .ZN(n6925) );
  INV_X1 U5705 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4539) );
  XNOR2_X1 U5706 ( .A(n5896), .B(n5895), .ZN(n5880) );
  NAND2_X1 U5707 ( .A1(n5449), .A2(n4874), .ZN(n7903) );
  XNOR2_X1 U5708 ( .A(n5321), .B(n5320), .ZN(n7659) );
  XNOR2_X1 U5709 ( .A(n4414), .B(n4922), .ZN(n6173) );
  NAND2_X1 U5710 ( .A1(n4415), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4414) );
  NAND2_X1 U5711 ( .A1(n4921), .A2(n4920), .ZN(n4415) );
  XNOR2_X1 U5712 ( .A(n4413), .B(n4886), .ZN(n6150) );
  NAND2_X1 U5713 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4413) );
  NAND2_X1 U5714 ( .A1(n4529), .A2(n4593), .ZN(P2_U3244) );
  OR2_X1 U5715 ( .A1(n8250), .A2(n8249), .ZN(n4593) );
  NAND2_X1 U5716 ( .A1(n4531), .A2(n4530), .ZN(n4529) );
  NAND2_X1 U5717 ( .A1(n8452), .A2(n5490), .ZN(n6021) );
  MUX2_X1 U5718 ( .A(n9639), .B(n9638), .S(n10007), .Z(n9640) );
  NAND2_X1 U5719 ( .A1(n8452), .A2(n5507), .ZN(n6025) );
  INV_X1 U5720 ( .A(n6053), .ZN(n6054) );
  OAI21_X1 U5721 ( .B1(n4438), .B2(n9767), .A(n6052), .ZN(n6053) );
  AOI21_X1 U5722 ( .B1(n9401), .B2(n5507), .A(n5479), .ZN(n5480) );
  OR2_X1 U5723 ( .A1(n5487), .A2(n9994), .ZN(n5481) );
  OR2_X1 U5724 ( .A1(n4515), .A2(n8161), .ZN(n4322) );
  INV_X2 U5725 ( .A(n6498), .ZN(n8716) );
  NAND2_X1 U5726 ( .A1(n5346), .A2(n5345), .ZN(n5355) );
  NAND3_X1 U5727 ( .A1(n5560), .A2(n4839), .A3(n4610), .ZN(n4323) );
  OR2_X1 U5728 ( .A1(n9146), .A2(n9010), .ZN(n8175) );
  AND2_X1 U5729 ( .A1(n4678), .A2(n5088), .ZN(n4324) );
  AND2_X1 U5730 ( .A1(n9539), .A2(n5444), .ZN(n4325) );
  AND2_X1 U5731 ( .A1(n9504), .A2(n4717), .ZN(n4326) );
  AND2_X1 U5732 ( .A1(n8699), .A2(n8700), .ZN(n4327) );
  AND2_X1 U5733 ( .A1(n4713), .A2(n4354), .ZN(n4328) );
  AND2_X1 U5734 ( .A1(n9427), .A2(n9647), .ZN(n4329) );
  AND2_X1 U5735 ( .A1(n5846), .A2(n5845), .ZN(n8988) );
  AND2_X1 U5736 ( .A1(n4491), .A2(n4490), .ZN(n4330) );
  AND2_X1 U5737 ( .A1(n4618), .A2(n4621), .ZN(n4331) );
  NOR2_X1 U5738 ( .A1(n6807), .A2(n8825), .ZN(n4332) );
  AND2_X1 U5739 ( .A1(n8142), .A2(n8143), .ZN(n8224) );
  NAND2_X1 U5740 ( .A1(n6873), .A2(n7001), .ZN(n4333) );
  NAND2_X1 U5741 ( .A1(n5946), .A2(n5921), .ZN(n4334) );
  AND2_X1 U5742 ( .A1(n8162), .A2(n9070), .ZN(n4335) );
  AND2_X1 U5743 ( .A1(n9127), .A2(n5912), .ZN(n8186) );
  AND2_X1 U5744 ( .A1(n9533), .A2(n5424), .ZN(n8424) );
  NAND2_X1 U5745 ( .A1(n8175), .A2(n8176), .ZN(n8982) );
  INV_X1 U5746 ( .A(n8982), .ZN(n8986) );
  AND2_X1 U5747 ( .A1(n4802), .A2(n8988), .ZN(n4336) );
  AND2_X1 U5748 ( .A1(n4487), .A2(n4486), .ZN(n4337) );
  AND2_X1 U5749 ( .A1(n5027), .A2(n5003), .ZN(n4338) );
  NAND2_X1 U5750 ( .A1(n7627), .A2(n4499), .ZN(n4500) );
  INV_X1 U5751 ( .A(n7177), .ZN(n4623) );
  NAND2_X1 U5752 ( .A1(n6621), .A2(n6622), .ZN(n6756) );
  INV_X2 U5753 ( .A(n6615), .ZN(n6498) );
  OR2_X1 U5754 ( .A1(n9427), .A2(n9647), .ZN(n4339) );
  INV_X1 U5755 ( .A(n5653), .ZN(n4739) );
  AND2_X1 U5756 ( .A1(n9460), .A2(n4627), .ZN(n4340) );
  NOR2_X1 U5757 ( .A1(n7804), .A2(n4777), .ZN(n4341) );
  OR2_X1 U5758 ( .A1(n9188), .A2(n7907), .ZN(n8066) );
  AND2_X1 U5759 ( .A1(n9454), .A2(n9648), .ZN(n4342) );
  XNOR2_X1 U5760 ( .A(n5943), .B(n5942), .ZN(n5953) );
  NAND2_X1 U5761 ( .A1(n6804), .A2(n6803), .ZN(n4343) );
  NOR2_X1 U5762 ( .A1(n9266), .A2(n4327), .ZN(n4344) );
  INV_X1 U5763 ( .A(n4605), .ZN(n7953) );
  AND2_X1 U5764 ( .A1(n8066), .A2(n4608), .ZN(n4345) );
  NOR2_X1 U5765 ( .A1(n8234), .A2(n8198), .ZN(n4346) );
  AOI21_X1 U5766 ( .B1(n5429), .B2(n4440), .A(n4583), .ZN(n4582) );
  NAND2_X1 U5767 ( .A1(n5988), .A2(n5987), .ZN(n8409) );
  INV_X1 U5768 ( .A(n8409), .ZN(n4438) );
  NAND2_X1 U5769 ( .A1(n5565), .A2(n5564), .ZN(n9177) );
  NAND2_X1 U5770 ( .A1(n8059), .A2(n8188), .ZN(n6028) );
  NAND2_X1 U5771 ( .A1(n9025), .A2(n5968), .ZN(n9008) );
  NAND2_X1 U5772 ( .A1(n8062), .A2(n9006), .ZN(n9017) );
  INV_X1 U5773 ( .A(n9017), .ZN(n9026) );
  INV_X1 U5774 ( .A(n7202), .ZN(n4785) );
  AND3_X1 U5775 ( .A1(n4560), .A2(n4559), .A3(n4957), .ZN(n4347) );
  NAND3_X1 U5776 ( .A1(n5591), .A2(n5590), .A3(n5589), .ZN(n6384) );
  NAND2_X1 U5777 ( .A1(n5246), .A2(n5245), .ZN(n9752) );
  NOR2_X1 U5778 ( .A1(n8787), .A2(n7036), .ZN(n4348) );
  NAND2_X1 U5779 ( .A1(n5279), .A2(n5278), .ZN(n9502) );
  NAND2_X1 U5780 ( .A1(n5882), .A2(n5881), .ZN(n8640) );
  AND2_X1 U5781 ( .A1(n8605), .A2(n8604), .ZN(n4349) );
  NOR2_X1 U5782 ( .A1(n4999), .A2(n6150), .ZN(n4350) );
  INV_X1 U5783 ( .A(n8518), .ZN(n4556) );
  NAND2_X1 U5784 ( .A1(n5815), .A2(n5814), .ZN(n9164) );
  INV_X1 U5785 ( .A(n9243), .ZN(n4661) );
  INV_X1 U5786 ( .A(n9401), .ZN(n8720) );
  NAND2_X1 U5787 ( .A1(n4558), .A2(n4860), .ZN(n4351) );
  NOR2_X1 U5788 ( .A1(n6598), .A2(n4391), .ZN(n4352) );
  XNOR2_X1 U5789 ( .A(n5089), .B(SI_11_), .ZN(n5088) );
  NAND2_X1 U5790 ( .A1(n5757), .A2(n5756), .ZN(n7895) );
  XNOR2_X1 U5791 ( .A(n4997), .B(SI_6_), .ZN(n4994) );
  AND2_X1 U5792 ( .A1(n8170), .A2(n9026), .ZN(n4353) );
  NAND2_X1 U5793 ( .A1(n9491), .A2(n9510), .ZN(n4354) );
  INV_X1 U5794 ( .A(n9613), .ZN(n4427) );
  INV_X1 U5795 ( .A(n9140), .ZN(n5868) );
  NAND2_X1 U5796 ( .A1(n5859), .A2(n5858), .ZN(n9140) );
  NAND2_X1 U5797 ( .A1(n9276), .A2(n8673), .ZN(n4355) );
  INV_X1 U5798 ( .A(n4804), .ZN(n4803) );
  NAND2_X1 U5799 ( .A1(n9164), .A2(n9038), .ZN(n4356) );
  AND2_X1 U5800 ( .A1(n8479), .A2(n8307), .ZN(n8429) );
  AND2_X1 U5801 ( .A1(n9502), .A2(n9682), .ZN(n4357) );
  NOR2_X1 U5802 ( .A1(n9491), .A2(n9510), .ZN(n4358) );
  INV_X1 U5803 ( .A(n4826), .ZN(n4825) );
  NAND2_X1 U5804 ( .A1(n9099), .A2(n9075), .ZN(n4826) );
  AND2_X1 U5805 ( .A1(n4905), .A2(n4854), .ZN(n4941) );
  INV_X1 U5806 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5181) );
  OR2_X1 U5807 ( .A1(n4756), .A2(n4755), .ZN(n4359) );
  AND2_X1 U5808 ( .A1(n4997), .A2(SI_6_), .ZN(n4360) );
  NOR2_X1 U5809 ( .A1(n8705), .A2(n8704), .ZN(n4361) );
  NOR2_X1 U5810 ( .A1(n5355), .A2(n9656), .ZN(n4362) );
  AND2_X1 U5811 ( .A1(n8526), .A2(n8466), .ZN(n8571) );
  INV_X1 U5812 ( .A(n8571), .ZN(n4440) );
  NAND3_X1 U5813 ( .A1(n4860), .A2(n4840), .A3(n4735), .ZN(n4363) );
  NAND2_X1 U5814 ( .A1(n5197), .A2(n4671), .ZN(n4364) );
  OR2_X1 U5815 ( .A1(n4736), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n4365) );
  AND2_X1 U5816 ( .A1(n8147), .A2(n8146), .ZN(n8223) );
  INV_X1 U5817 ( .A(n8223), .ZN(n4814) );
  AND2_X1 U5818 ( .A1(n4828), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4366) );
  AND2_X1 U5819 ( .A1(n5090), .A2(SI_11_), .ZN(n4367) );
  AND2_X1 U5820 ( .A1(n4707), .A2(n4339), .ZN(n4368) );
  INV_X1 U5821 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4828) );
  INV_X1 U5822 ( .A(n4860), .ZN(n5118) );
  AND3_X1 U5823 ( .A1(n5096), .A2(n4347), .A3(n4941), .ZN(n4860) );
  OR2_X1 U5824 ( .A1(n7895), .A2(n7906), .ZN(n8147) );
  OR2_X1 U5825 ( .A1(n4753), .A2(n4751), .ZN(n4369) );
  NAND2_X1 U5826 ( .A1(n8155), .A2(n4521), .ZN(n4370) );
  INV_X1 U5827 ( .A(n6868), .ZN(n4640) );
  INV_X1 U5828 ( .A(n4758), .ZN(n4757) );
  NOR2_X1 U5829 ( .A1(n4759), .A2(n8634), .ZN(n4758) );
  INV_X1 U5830 ( .A(n4590), .ZN(n4589) );
  NAND2_X1 U5831 ( .A1(n8986), .A2(n4591), .ZN(n4590) );
  NAND2_X1 U5832 ( .A1(n9008), .A2(n8172), .ZN(n8985) );
  AND2_X1 U5833 ( .A1(n5425), .A2(n8518), .ZN(n4371) );
  AND2_X1 U5834 ( .A1(n4705), .A2(n4339), .ZN(n4372) );
  AND2_X1 U5835 ( .A1(n6813), .A2(n4343), .ZN(n4373) );
  NAND2_X1 U5836 ( .A1(n5121), .A2(n5120), .ZN(n7859) );
  AND3_X1 U5837 ( .A1(n4735), .A2(n5453), .A3(n4734), .ZN(n4374) );
  AND2_X1 U5838 ( .A1(n4624), .A2(n4623), .ZN(n4375) );
  NAND2_X1 U5839 ( .A1(n5101), .A2(n5100), .ZN(n7799) );
  AND2_X1 U5840 ( .A1(n4369), .A2(n4743), .ZN(n4376) );
  AND2_X1 U5841 ( .A1(n4811), .A2(n4809), .ZN(n4377) );
  AND2_X1 U5842 ( .A1(n4822), .A2(n4356), .ZN(n4378) );
  OR2_X1 U5843 ( .A1(n10081), .A2(n8238), .ZN(n7025) );
  NAND2_X1 U5844 ( .A1(n6012), .A2(n6011), .ZN(n8452) );
  INV_X1 U5845 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4527) );
  AND2_X1 U5846 ( .A1(n9621), .A2(n9607), .ZN(n9574) );
  NAND2_X1 U5847 ( .A1(n5838), .A2(n5837), .ZN(n9149) );
  INV_X1 U5848 ( .A(n9149), .ZN(n4802) );
  INV_X1 U5849 ( .A(n8509), .ZN(n4461) );
  OR2_X1 U5850 ( .A1(n7177), .A2(n9963), .ZN(n8490) );
  INV_X1 U5851 ( .A(n8490), .ZN(n4574) );
  NAND2_X1 U5852 ( .A1(n4733), .A2(n5070), .ZN(n9832) );
  AND3_X1 U5853 ( .A1(n4853), .A2(n4851), .A3(n4852), .ZN(n5096) );
  NAND2_X1 U5854 ( .A1(n5903), .A2(n5902), .ZN(n9127) );
  INV_X1 U5855 ( .A(n9127), .ZN(n4486) );
  AND2_X1 U5856 ( .A1(n7974), .A2(n7973), .ZN(n4379) );
  AND2_X1 U5857 ( .A1(n6240), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4380) );
  NAND2_X1 U5858 ( .A1(n9110), .A2(n4493), .ZN(n4494) );
  AND2_X1 U5859 ( .A1(n4408), .A2(n4407), .ZN(n4381) );
  AND2_X1 U5860 ( .A1(n7859), .A2(n9854), .ZN(n4382) );
  AND2_X1 U5861 ( .A1(n4784), .A2(n4782), .ZN(n4383) );
  OR2_X1 U5862 ( .A1(n7216), .A2(n7217), .ZN(n4408) );
  NOR2_X1 U5863 ( .A1(n7932), .A2(n9615), .ZN(n4384) );
  NAND2_X1 U5864 ( .A1(n9539), .A2(n4620), .ZN(n4622) );
  AND2_X1 U5865 ( .A1(n5212), .A2(SI_17_), .ZN(n4385) );
  INV_X1 U5866 ( .A(n8626), .ZN(n4762) );
  AND2_X1 U5867 ( .A1(n8625), .A2(n8624), .ZN(n8626) );
  NAND2_X1 U5868 ( .A1(n9752), .A2(n9681), .ZN(n4386) );
  NAND2_X1 U5869 ( .A1(n5296), .A2(n5295), .ZN(n9491) );
  INV_X1 U5870 ( .A(n9491), .ZN(n4621) );
  NAND2_X1 U5871 ( .A1(n4645), .A2(n4644), .ZN(n7645) );
  NAND2_X1 U5872 ( .A1(n4615), .A2(n5560), .ZN(n5913) );
  NAND2_X1 U5873 ( .A1(n5826), .A2(n5825), .ZN(n9161) );
  INV_X1 U5874 ( .A(n9161), .ZN(n4490) );
  AND2_X1 U5875 ( .A1(n5442), .A2(n4624), .ZN(n4387) );
  NOR2_X1 U5876 ( .A1(n7385), .A2(n9785), .ZN(n5443) );
  INV_X1 U5877 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4735) );
  NOR2_X1 U5878 ( .A1(n7016), .A2(n8211), .ZN(n7015) );
  INV_X1 U5879 ( .A(n7015), .ZN(n4597) );
  NAND2_X1 U5880 ( .A1(n5770), .A2(n5769), .ZN(n9191) );
  INV_X1 U5881 ( .A(n9191), .ZN(n4496) );
  OAI21_X1 U5882 ( .B1(n6897), .B2(n8212), .A(n8108), .ZN(n7016) );
  OR2_X1 U5883 ( .A1(n7384), .A2(n4631), .ZN(n4388) );
  OR2_X1 U5884 ( .A1(n7015), .A2(n4601), .ZN(n6983) );
  NAND2_X1 U5885 ( .A1(n4769), .A2(n4373), .ZN(n7024) );
  NAND2_X1 U5886 ( .A1(n4830), .A2(n5676), .ZN(n6978) );
  NAND2_X1 U5887 ( .A1(n5560), .A2(n4839), .ZN(n5916) );
  INV_X1 U5888 ( .A(n4845), .ZN(n4722) );
  INV_X1 U5889 ( .A(n7013), .ZN(n4503) );
  AND2_X1 U5890 ( .A1(n5953), .A2(n8056), .ZN(n8198) );
  NAND2_X1 U5891 ( .A1(n5707), .A2(n5706), .ZN(n10132) );
  INV_X1 U5892 ( .A(n10132), .ZN(n4506) );
  INV_X1 U5893 ( .A(n9408), .ZN(n9513) );
  OR2_X1 U5894 ( .A1(n8458), .A2(n8591), .ZN(n4389) );
  OR2_X1 U5895 ( .A1(n8055), .A2(n5952), .ZN(n4390) );
  INV_X1 U5896 ( .A(n6277), .ZN(n4740) );
  INV_X1 U5897 ( .A(n7073), .ZN(n4420) );
  XNOR2_X1 U5898 ( .A(n5947), .B(n5946), .ZN(n8916) );
  INV_X1 U5899 ( .A(n5547), .ZN(n9214) );
  NOR2_X1 U5900 ( .A1(n4874), .A2(n4365), .ZN(n9769) );
  OR2_X1 U5901 ( .A1(n10072), .A2(n6482), .ZN(n8975) );
  OR3_X2 U5902 ( .A1(n6357), .A2(n9969), .A3(n6356), .ZN(n9315) );
  AND2_X1 U5903 ( .A1(n9931), .A2(n8586), .ZN(n9969) );
  NOR2_X4 U5904 ( .A1(n7653), .A2(n9988), .ZN(n9320) );
  NAND2_X1 U5905 ( .A1(n8866), .A2(n6262), .ZN(n6516) );
  XNOR2_X1 U5906 ( .A(n7663), .B(n7668), .ZN(n7216) );
  INV_X1 U5907 ( .A(n7124), .ZN(n6726) );
  NAND2_X2 U5908 ( .A1(n4999), .A2(n5527), .ZN(n8397) );
  AOI21_X2 U5909 ( .B1(n4439), .B2(n8395), .A(n8394), .ZN(n8410) );
  NAND2_X2 U5910 ( .A1(n4482), .A2(n4484), .ZN(n8386) );
  NAND2_X1 U5911 ( .A1(n4979), .A2(n4444), .ZN(n4443) );
  NAND2_X1 U5912 ( .A1(n4443), .A2(n4446), .ZN(n5006) );
  OAI21_X2 U5913 ( .B1(n4454), .B2(n8460), .A(n8534), .ZN(n4453) );
  OR2_X2 U5914 ( .A1(n8419), .A2(n8418), .ZN(n4454) );
  NAND2_X1 U5915 ( .A1(n4458), .A2(n4455), .ZN(n8368) );
  NAND2_X1 U5916 ( .A1(n4456), .A2(n8415), .ZN(n4455) );
  NAND2_X1 U5917 ( .A1(n4457), .A2(n8512), .ZN(n4456) );
  NAND2_X1 U5918 ( .A1(n4464), .A2(n8510), .ZN(n4457) );
  NAND2_X1 U5919 ( .A1(n4459), .A2(n8402), .ZN(n4458) );
  NAND2_X1 U5920 ( .A1(n4462), .A2(n4460), .ZN(n4459) );
  NAND2_X1 U5921 ( .A1(n4464), .A2(n4463), .ZN(n4462) );
  AND2_X1 U5922 ( .A1(n8357), .A2(n8356), .ZN(n4463) );
  NAND2_X1 U5923 ( .A1(n8354), .A2(n8355), .ZN(n4464) );
  NAND3_X1 U5924 ( .A1(n4324), .A2(n4473), .A3(n4465), .ZN(n4468) );
  NAND2_X1 U5925 ( .A1(n4466), .A2(n4475), .ZN(n4465) );
  AND2_X1 U5926 ( .A1(n5052), .A2(n4472), .ZN(n4466) );
  NAND2_X1 U5927 ( .A1(n5030), .A2(n5029), .ZN(n4475) );
  NAND3_X1 U5928 ( .A1(n4469), .A2(n4676), .A3(n4468), .ZN(n5113) );
  NAND2_X1 U5929 ( .A1(n5031), .A2(n5029), .ZN(n4470) );
  INV_X1 U5930 ( .A(n5029), .ZN(n4472) );
  OR2_X1 U5931 ( .A1(n5031), .A2(n5030), .ZN(n4474) );
  NAND2_X1 U5932 ( .A1(n5194), .A2(n5193), .ZN(n4481) );
  AND2_X1 U5933 ( .A1(n8990), .A2(n4489), .ZN(n8955) );
  INV_X1 U5934 ( .A(n4494), .ZN(n9083) );
  INV_X1 U5935 ( .A(n4500), .ZN(n7724) );
  NAND3_X1 U5936 ( .A1(n4504), .A2(n4501), .A3(n4506), .ZN(n7254) );
  NAND3_X1 U5937 ( .A1(n4346), .A2(n8190), .A3(n8193), .ZN(n4509) );
  NAND2_X1 U5938 ( .A1(n8153), .A2(n4518), .ZN(n4514) );
  NAND2_X1 U5939 ( .A1(n4514), .A2(n8155), .ZN(n8160) );
  NAND2_X1 U5940 ( .A1(n4520), .A2(n4519), .ZN(n8157) );
  INV_X1 U5941 ( .A(n8161), .ZN(n4521) );
  NAND2_X1 U5942 ( .A1(n5780), .A2(n4526), .ZN(n4525) );
  MUX2_X1 U5943 ( .A(n8076), .B(n8077), .S(n8198), .Z(n8102) );
  NAND2_X4 U5944 ( .A1(n4868), .A2(n9779), .ZN(n4936) );
  XNOR2_X2 U5945 ( .A(n4540), .B(n4539), .ZN(n9779) );
  NAND2_X1 U5946 ( .A1(n8301), .A2(n8551), .ZN(n4541) );
  NAND2_X1 U5947 ( .A1(n8300), .A2(n8486), .ZN(n8301) );
  NAND2_X1 U5948 ( .A1(n5415), .A2(n8477), .ZN(n8300) );
  OAI21_X1 U5949 ( .B1(n9614), .B2(n4545), .A(n4542), .ZN(n9584) );
  INV_X1 U5950 ( .A(n9584), .ZN(n5421) );
  NAND2_X1 U5951 ( .A1(n9553), .A2(n4547), .ZN(n4546) );
  NAND2_X1 U5952 ( .A1(n4546), .A2(n4549), .ZN(n9519) );
  NAND2_X1 U5953 ( .A1(n9503), .A2(n4371), .ZN(n4553) );
  NAND2_X1 U5954 ( .A1(n4553), .A2(n4554), .ZN(n9469) );
  AND4_X2 U5956 ( .A1(n5096), .A2(n4347), .A3(n4941), .A4(n4861), .ZN(n4557)
         );
  NAND2_X1 U5957 ( .A1(n7785), .A2(n4564), .ZN(n4563) );
  AND2_X1 U5958 ( .A1(n5420), .A2(n4566), .ZN(n4562) );
  NAND2_X1 U5959 ( .A1(n4563), .A2(n4562), .ZN(n7924) );
  NAND2_X1 U5960 ( .A1(n4571), .A2(n4569), .ZN(n9837) );
  INV_X1 U5961 ( .A(n4570), .ZN(n4569) );
  OAI21_X1 U5962 ( .B1(n8491), .B2(n4573), .A(n8471), .ZN(n4570) );
  NOR2_X1 U5963 ( .A1(n8491), .A2(n4574), .ZN(n4572) );
  INV_X1 U5964 ( .A(n9837), .ZN(n5418) );
  OAI211_X1 U5965 ( .C1(n5496), .C2(n4578), .A(n4576), .B(n4575), .ZN(n5999)
         );
  NAND2_X1 U5966 ( .A1(n5496), .A2(n4579), .ZN(n4575) );
  INV_X1 U5967 ( .A(n4582), .ZN(n4577) );
  NAND2_X1 U5968 ( .A1(n4582), .A2(n4581), .ZN(n4578) );
  NAND2_X1 U5969 ( .A1(n5497), .A2(n5429), .ZN(n5990) );
  NAND2_X1 U5970 ( .A1(n4588), .A2(n4586), .ZN(n8962) );
  NAND2_X1 U5971 ( .A1(n7890), .A2(n4345), .ZN(n4604) );
  NAND4_X1 U5972 ( .A1(n5560), .A2(n4839), .A3(n4614), .A4(n5917), .ZN(n5540)
         );
  NAND2_X1 U5974 ( .A1(n9035), .A2(n5967), .ZN(n9034) );
  AOI21_X1 U5975 ( .B1(n6032), .B2(n8232), .A(n5969), .ZN(n5970) );
  NOR3_X1 U5976 ( .A1(n7249), .A2(n7248), .A3(n8219), .ZN(n7317) );
  OAI21_X1 U5977 ( .B1(n7317), .B2(n8127), .A(n8134), .ZN(n7622) );
  AOI22_X1 U5978 ( .A1(n8035), .A2(n8034), .B1(n8191), .B2(n8033), .ZN(n8052)
         );
  NOR2_X2 U5979 ( .A1(n7717), .A2(n5963), .ZN(n7890) );
  NAND2_X1 U5980 ( .A1(n9068), .A2(n5965), .ZN(n9058) );
  NAND2_X1 U5981 ( .A1(n8950), .A2(n8949), .ZN(n8948) );
  OR2_X1 U5982 ( .A1(n5487), .A2(n10005), .ZN(n5492) );
  NOR2_X1 U5983 ( .A1(n9331), .A2(n8427), .ZN(n8428) );
  NOR2_X1 U5984 ( .A1(n9455), .A2(n5426), .ZN(n9438) );
  NAND2_X1 U5985 ( .A1(n5959), .A2(n10041), .ZN(n10044) );
  NAND2_X1 U5986 ( .A1(n6914), .A2(n6919), .ZN(n6691) );
  NAND2_X1 U5987 ( .A1(n5970), .A2(n8205), .ZN(n8035) );
  NAND2_X1 U5988 ( .A1(n9100), .A2(n9101), .ZN(n9068) );
  INV_X1 U5989 ( .A(n8207), .ZN(n5956) );
  NAND2_X1 U5990 ( .A1(n5957), .A2(n5956), .ZN(n6950) );
  AND3_X4 U5991 ( .A1(n5518), .A2(n5517), .A3(n5571), .ZN(n5560) );
  INV_X2 U5992 ( .A(n5576), .ZN(n5653) );
  INV_X1 U5993 ( .A(n10042), .ZN(n10041) );
  NAND2_X1 U5994 ( .A1(n9211), .A2(n4818), .ZN(n5546) );
  NAND2_X1 U5995 ( .A1(n10044), .A2(n8078), .ZN(n6959) );
  NAND2_X2 U5996 ( .A1(n5433), .A2(n8588), .ZN(n4999) );
  XNOR2_X2 U5997 ( .A(n4616), .B(n4873), .ZN(n5433) );
  INV_X1 U5998 ( .A(n4622), .ZN(n9529) );
  NAND2_X1 U5999 ( .A1(n9460), .A2(n4625), .ZN(n6000) );
  NAND2_X1 U6000 ( .A1(n4635), .A2(n4633), .ZN(n6883) );
  INV_X1 U6001 ( .A(n4634), .ZN(n4633) );
  OAI21_X1 U6002 ( .B1(n6755), .B2(n4639), .A(n4850), .ZN(n4634) );
  NAND2_X1 U6003 ( .A1(n6756), .A2(n6755), .ZN(n6869) );
  NAND2_X1 U6004 ( .A1(n5409), .A2(n5406), .ZN(n4643) );
  NAND2_X1 U6005 ( .A1(n7080), .A2(n4646), .ZN(n4645) );
  NAND2_X1 U6006 ( .A1(n4655), .A2(n4654), .ZN(n4653) );
  INV_X1 U6007 ( .A(n7239), .ZN(n4654) );
  NAND3_X1 U6008 ( .A1(n8661), .A2(n9299), .A3(n4660), .ZN(n4657) );
  NAND2_X1 U6009 ( .A1(n4657), .A2(n4658), .ZN(n9251) );
  NAND3_X1 U6010 ( .A1(n8661), .A2(n9299), .A3(n4661), .ZN(n9277) );
  OAI21_X1 U6011 ( .B1(n9266), .B2(n4663), .A(n4662), .ZN(n4668) );
  NAND2_X1 U6012 ( .A1(n9266), .A2(n4669), .ZN(n4666) );
  INV_X1 U6013 ( .A(n9259), .ZN(n4669) );
  NAND2_X1 U6014 ( .A1(n5197), .A2(n4670), .ZN(n5404) );
  OAI21_X2 U6015 ( .B1(n7992), .B2(n7991), .A(n7990), .ZN(n8646) );
  NAND2_X2 U6016 ( .A1(n4672), .A2(n5008), .ZN(n5031) );
  NAND2_X1 U6017 ( .A1(n5006), .A2(n5005), .ZN(n4672) );
  NAND3_X1 U6018 ( .A1(n4674), .A2(n4673), .A3(n4882), .ZN(n5595) );
  NAND2_X1 U6019 ( .A1(n5135), .A2(n4693), .ZN(n4688) );
  NAND2_X1 U6020 ( .A1(n5135), .A2(n5134), .ZN(n5153) );
  NAND2_X1 U6021 ( .A1(n5276), .A2(n4700), .ZN(n4695) );
  NAND2_X1 U6022 ( .A1(n5276), .A2(n5275), .ZN(n5291) );
  NAND2_X1 U6023 ( .A1(n4702), .A2(n8433), .ZN(n6635) );
  NAND2_X1 U6024 ( .A1(n9450), .A2(n4372), .ZN(n4704) );
  NAND2_X1 U6025 ( .A1(n9521), .A2(n4328), .ZN(n4711) );
  NAND2_X1 U6026 ( .A1(n4720), .A2(n6787), .ZN(n4719) );
  NAND2_X1 U6027 ( .A1(n7788), .A2(n4725), .ZN(n4724) );
  NAND2_X1 U6028 ( .A1(n7383), .A2(n8439), .ZN(n4733) );
  NAND4_X1 U6029 ( .A1(n4860), .A2(n4840), .A3(n4735), .A4(n5453), .ZN(n5450)
         );
  NAND2_X1 U6030 ( .A1(n7106), .A2(n4338), .ZN(n7166) );
  NAND2_X1 U6031 ( .A1(n7166), .A2(n5028), .ZN(n7301) );
  NOR2_X1 U6032 ( .A1(n4874), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n4877) );
  NAND2_X1 U6033 ( .A1(n6080), .A2(n8047), .ZN(n4738) );
  NAND2_X1 U6034 ( .A1(n8757), .A2(n4742), .ZN(n4741) );
  OAI21_X1 U6035 ( .B1(n8757), .B2(n8758), .A(n4749), .ZN(n8803) );
  OAI211_X1 U6036 ( .C1(n8757), .C2(n4746), .A(n4376), .B(n4741), .ZN(n8642)
         );
  NAND2_X1 U6037 ( .A1(n4765), .A2(n6681), .ZN(n6806) );
  NAND3_X1 U6038 ( .A1(n4765), .A2(n6681), .A3(n4373), .ZN(n4764) );
  NAND2_X1 U6039 ( .A1(n7733), .A2(n4774), .ZN(n4772) );
  NAND2_X1 U6040 ( .A1(n7203), .A2(n4782), .ZN(n4779) );
  XNOR2_X2 U6041 ( .A(n7701), .B(n7702), .ZN(n7700) );
  NAND2_X1 U6042 ( .A1(n8003), .A2(n4791), .ZN(n4789) );
  NAND4_X1 U6043 ( .A1(n5560), .A2(n4839), .A3(n5523), .A4(n5917), .ZN(n5526)
         );
  NAND2_X1 U6044 ( .A1(n9018), .A2(n4799), .ZN(n4798) );
  NOR2_X1 U6045 ( .A1(n9023), .A2(n9009), .ZN(n4804) );
  NAND2_X1 U6046 ( .A1(n8944), .A2(n5879), .ZN(n6029) );
  INV_X1 U6047 ( .A(n4817), .ZN(n7715) );
  OR2_X1 U6048 ( .A1(n7895), .A2(n8819), .ZN(n4815) );
  NOR2_X1 U6050 ( .A1(n5803), .A2(n4825), .ZN(n9081) );
  OAI21_X1 U6051 ( .B1(n5803), .B2(n4821), .A(n4378), .ZN(n4820) );
  NAND2_X1 U6052 ( .A1(n4830), .A2(n4829), .ZN(n6980) );
  XNOR2_X1 U6053 ( .A(n5493), .B(n8571), .ZN(n9410) );
  NAND2_X1 U6054 ( .A1(n9410), .A2(n9992), .ZN(n5495) );
  OR2_X1 U6055 ( .A1(n8943), .A2(n10146), .ZN(n6042) );
  INV_X1 U6056 ( .A(n8657), .ZN(n8660) );
  CLKBUF_X1 U6057 ( .A(n6683), .Z(n10009) );
  INV_X1 U6058 ( .A(n6507), .ZN(n6504) );
  NAND2_X1 U6059 ( .A1(n6463), .A2(n7025), .ZN(n6469) );
  AND2_X1 U6060 ( .A1(n9331), .A2(n9932), .ZN(n6829) );
  NAND2_X1 U6061 ( .A1(n6692), .A2(n6910), .ZN(n8092) );
  OR2_X1 U6062 ( .A1(n4936), .A2(n6131), .ZN(n4870) );
  NAND2_X1 U6063 ( .A1(n8778), .A2(n8777), .ZN(n8776) );
  NAND2_X1 U6064 ( .A1(n7620), .A2(n4834), .ZN(n7716) );
  AND2_X1 U6065 ( .A1(n9060), .A2(n9059), .ZN(n4831) );
  INV_X1 U6066 ( .A(n8424), .ZN(n5422) );
  NAND2_X1 U6067 ( .A1(n9706), .A2(n9712), .ZN(n4833) );
  OR2_X1 U6068 ( .A1(n4438), .A2(n9728), .ZN(n4835) );
  AND2_X1 U6069 ( .A1(n9026), .A2(n9024), .ZN(n4836) );
  AND2_X1 U6070 ( .A1(n4835), .A2(n6004), .ZN(n4838) );
  AND4_X1 U6071 ( .A1(n5440), .A2(n5439), .A3(n5438), .A4(n5437), .ZN(n9397)
         );
  INV_X1 U6072 ( .A(n9962), .ZN(n5499) );
  INV_X1 U6073 ( .A(n4936), .ZN(n5042) );
  XNOR2_X1 U6074 ( .A(n6751), .B(n8689), .ZN(n6865) );
  AND2_X1 U6075 ( .A1(n6014), .A2(n9847), .ZN(n4842) );
  INV_X1 U6076 ( .A(n8640), .ZN(n5893) );
  INV_X1 U6077 ( .A(n6028), .ZN(n8232) );
  OR2_X1 U6078 ( .A1(n9130), .A2(n10070), .ZN(n4843) );
  INV_X1 U6079 ( .A(n7895), .ZN(n5978) );
  OR2_X1 U6080 ( .A1(n8720), .A2(n9228), .ZN(n4844) );
  INV_X1 U6081 ( .A(n9228), .ZN(n5500) );
  AND2_X1 U6082 ( .A1(n9326), .A2(n7007), .ZN(n4845) );
  XOR2_X1 U6083 ( .A(n9154), .B(n8631), .Z(n4846) );
  NOR2_X1 U6084 ( .A1(n7640), .A2(n7639), .ZN(n4847) );
  AND2_X1 U6085 ( .A1(n7784), .A2(n8337), .ZN(n9835) );
  NAND2_X1 U6086 ( .A1(n5738), .A2(n7260), .ZN(n4848) );
  AND2_X1 U6087 ( .A1(n6878), .A2(n7145), .ZN(n4850) );
  AOI21_X1 U6088 ( .B1(n8386), .B2(n8385), .A(n8384), .ZN(n8388) );
  INV_X1 U6089 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n4855) );
  AND2_X1 U6090 ( .A1(n8570), .A2(n9414), .ZN(n8525) );
  INV_X1 U6091 ( .A(n8766), .ZN(n8611) );
  INV_X1 U6092 ( .A(n8110), .ZN(n5961) );
  NAND2_X1 U6093 ( .A1(n5423), .A2(n5422), .ZN(n9503) );
  INV_X1 U6094 ( .A(n6469), .ZN(n6466) );
  NAND2_X1 U6095 ( .A1(n8613), .A2(n8767), .ZN(n8614) );
  INV_X1 U6096 ( .A(n5829), .ZN(n5538) );
  INV_X1 U6097 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5572) );
  XNOR2_X1 U6098 ( .A(n6426), .B(n8689), .ZN(n6429) );
  AND2_X1 U6099 ( .A1(n9536), .A2(n4386), .ZN(n5253) );
  INV_X1 U6100 ( .A(n9752), .ZN(n5444) );
  INV_X1 U6101 ( .A(n8436), .ZN(n5027) );
  INV_X1 U6102 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5136) );
  INV_X1 U6103 ( .A(n5004), .ZN(n5005) );
  INV_X1 U6104 ( .A(n5670), .ZN(n5530) );
  NAND2_X1 U6105 ( .A1(n5538), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5839) );
  OR2_X1 U6106 ( .A1(n5745), .A2(n6781), .ZN(n5747) );
  AND2_X1 U6107 ( .A1(n5583), .A2(n5582), .ZN(n5586) );
  AOI22_X1 U6108 ( .A1(n8952), .A2(n10045), .B1(n8923), .B2(n8814), .ZN(n5975)
         );
  INV_X1 U6109 ( .A(n8220), .ZN(n7323) );
  OR2_X1 U6110 ( .A1(n6735), .A2(n6902), .ZN(n7011) );
  NOR2_X1 U6111 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5541) );
  INV_X2 U6112 ( .A(n6066), .ZN(n5527) );
  INV_X1 U6113 ( .A(n5367), .ZN(n5365) );
  INV_X1 U6114 ( .A(n6506), .ZN(n6503) );
  INV_X1 U6115 ( .A(n8658), .ZN(n8659) );
  NAND2_X1 U6116 ( .A1(n5266), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5280) );
  OR2_X1 U6117 ( .A1(n5124), .A2(n5123), .ZN(n5141) );
  INV_X1 U6118 ( .A(n9902), .ZN(n6240) );
  INV_X1 U6119 ( .A(n9543), .ZN(n5424) );
  NOR2_X1 U6120 ( .A1(n5141), .A2(n5140), .ZN(n5163) );
  NAND2_X1 U6121 ( .A1(n5080), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5103) );
  INV_X1 U6122 ( .A(n5355), .ZN(n9651) );
  INV_X1 U6123 ( .A(n6638), .ZN(n8433) );
  NAND2_X1 U6124 ( .A1(n5530), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5681) );
  INV_X1 U6125 ( .A(n8827), .ZN(n6985) );
  INV_X1 U6126 ( .A(n10047), .ZN(n6709) );
  NAND2_X1 U6127 ( .A1(n5860), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5884) );
  INV_X1 U6128 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8878) );
  AND2_X1 U6129 ( .A1(n8151), .A2(n8150), .ZN(n8225) );
  INV_X1 U6130 ( .A(n6970), .ZN(n10098) );
  INV_X1 U6131 ( .A(n5952), .ZN(n10133) );
  AND2_X1 U6132 ( .A1(n8712), .A2(n8711), .ZN(n8713) );
  AND2_X1 U6133 ( .A1(n9226), .A2(n9224), .ZN(n8717) );
  NAND2_X1 U6134 ( .A1(n8536), .A2(n9408), .ZN(n8537) );
  NAND2_X1 U6135 ( .A1(n5312), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5327) );
  INV_X1 U6136 ( .A(n4989), .ZN(n5328) );
  NAND2_X1 U6137 ( .A1(n9414), .A2(n8567), .ZN(n9437) );
  NAND2_X1 U6138 ( .A1(n8511), .A2(n8364), .ZN(n9504) );
  AND2_X1 U6139 ( .A1(n8344), .A2(n8336), .ZN(n8443) );
  OR2_X1 U6140 ( .A1(n9785), .A2(n7339), .ZN(n8329) );
  NAND2_X1 U6141 ( .A1(n10005), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6004) );
  OR2_X1 U6142 ( .A1(n9995), .A2(n6051), .ZN(n6052) );
  NAND2_X1 U6143 ( .A1(n8042), .A2(n8041), .ZN(n8046) );
  AND2_X1 U6144 ( .A1(n5195), .A2(n5176), .ZN(n5193) );
  AND2_X1 U6145 ( .A1(n5134), .A2(n5117), .ZN(n5132) );
  AND2_X1 U6146 ( .A1(n5054), .A2(n5035), .ZN(n5052) );
  OR3_X1 U6147 ( .A1(n5884), .A2(n8736), .A3(n5883), .ZN(n5981) );
  AND2_X1 U6148 ( .A1(n6295), .A2(n6294), .ZN(n10029) );
  OAI21_X1 U6149 ( .B1(n6730), .B2(n5652), .A(n5651), .ZN(n6896) );
  AND2_X1 U6150 ( .A1(n10039), .A2(n9814), .ZN(n10146) );
  NOR2_X1 U6151 ( .A1(n7920), .A2(n5929), .ZN(n10071) );
  OR2_X1 U6152 ( .A1(n8397), .A2(n6068), .ZN(n4889) );
  INV_X1 U6153 ( .A(n7647), .ZN(n7649) );
  AND2_X1 U6154 ( .A1(n8692), .A2(n8691), .ZN(n9290) );
  AND4_X1 U6155 ( .A1(n5286), .A2(n5285), .A3(n5284), .A4(n5283), .ZN(n9528)
         );
  AND2_X1 U6156 ( .A1(n8357), .A2(n8509), .ZN(n9547) );
  AND2_X1 U6157 ( .A1(n4833), .A2(n9552), .ZN(n9583) );
  OAI22_X1 U6158 ( .A1(n7301), .A2(n5051), .B1(n7311), .B2(n9975), .ZN(n7383)
         );
  INV_X1 U6159 ( .A(n9728), .ZN(n5490) );
  INV_X1 U6160 ( .A(n9767), .ZN(n5507) );
  OR2_X1 U6161 ( .A1(n9954), .A2(n9860), .ZN(n9992) );
  XNOR2_X1 U6162 ( .A(n4945), .B(n4929), .ZN(n4943) );
  INV_X1 U6163 ( .A(P2_U3966), .ZN(n8816) );
  AOI21_X1 U6164 ( .B1(n9128), .B2(n9088), .A(n5984), .ZN(n5985) );
  NAND2_X1 U6165 ( .A1(n6042), .A2(n6041), .ZN(n9132) );
  OR2_X1 U6166 ( .A1(n6393), .A2(n6459), .ZN(n10174) );
  OR2_X1 U6167 ( .A1(n6393), .A2(n6480), .ZN(n10156) );
  OR2_X1 U6168 ( .A1(n10072), .A2(n10071), .ZN(n10075) );
  AND4_X1 U6169 ( .A1(n5401), .A2(n5400), .A3(n5399), .A4(n5398), .ZN(n9228)
         );
  OR2_X1 U6170 ( .A1(n9939), .A2(n6838), .ZN(n9628) );
  OR2_X1 U6171 ( .A1(n9939), .A2(n6826), .ZN(n9589) );
  AOI21_X1 U6172 ( .B1(n9401), .B2(n5490), .A(n5489), .ZN(n5491) );
  INV_X1 U6173 ( .A(n10007), .ZN(n10005) );
  INV_X1 U6174 ( .A(n9533), .ZN(n9749) );
  INV_X1 U6175 ( .A(n9995), .ZN(n9994) );
  NAND2_X1 U6176 ( .A1(n6050), .A2(n6049), .ZN(P2_U3516) );
  NOR2_X1 U6177 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4859) );
  NOR2_X1 U6178 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n4858) );
  NOR2_X1 U6179 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n4857) );
  INV_X1 U6180 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4861) );
  INV_X1 U6181 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4862) );
  INV_X1 U6182 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4873) );
  INV_X1 U6183 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9770) );
  XNOR2_X2 U6184 ( .A(n4863), .B(n9770), .ZN(n4866) );
  NAND2_X1 U6185 ( .A1(n4933), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4872) );
  INV_X1 U6186 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n4865) );
  INV_X1 U6187 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6131) );
  INV_X1 U6188 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6835) );
  NOR2_X1 U6189 ( .A1(n4877), .A2(n4876), .ZN(n4878) );
  INV_X1 U6190 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6068) );
  AND2_X1 U6191 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4882) );
  AND2_X1 U6192 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4883) );
  NAND2_X1 U6193 ( .A1(n4928), .A2(n4883), .ZN(n4897) );
  NAND2_X1 U6194 ( .A1(n5595), .A2(n4897), .ZN(n4908) );
  INV_X1 U6195 ( .A(SI_1_), .ZN(n4884) );
  XNOR2_X1 U6196 ( .A(n4908), .B(n4884), .ZN(n4907) );
  XNOR2_X1 U6197 ( .A(n4907), .B(n4906), .ZN(n6067) );
  NOR2_X1 U6198 ( .A1(n4982), .A2(n6067), .ZN(n4887) );
  INV_X1 U6199 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4886) );
  NOR2_X1 U6200 ( .A1(n4887), .A2(n4350), .ZN(n4888) );
  AND2_X2 U6201 ( .A1(n4889), .A2(n4888), .ZN(n9943) );
  XNOR2_X2 U6202 ( .A(n6423), .B(n9943), .ZN(n6827) );
  INV_X1 U6203 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6123) );
  INV_X1 U6204 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n4890) );
  NAND2_X1 U6205 ( .A1(n6066), .A2(SI_0_), .ZN(n4896) );
  INV_X1 U6206 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n4895) );
  NAND2_X1 U6207 ( .A1(n4896), .A2(n4895), .ZN(n4898) );
  AND2_X1 U6208 ( .A1(n4898), .A2(n4897), .ZN(n9782) );
  MUX2_X1 U6209 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9782), .S(n4999), .Z(n9932) );
  NAND2_X1 U6210 ( .A1(n6423), .A2(n6839), .ZN(n4899) );
  NAND2_X1 U6211 ( .A1(n4933), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4904) );
  INV_X1 U6212 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6401) );
  OR2_X1 U6213 ( .A1(n4989), .A2(n6401), .ZN(n4903) );
  INV_X1 U6214 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6130) );
  OR2_X1 U6215 ( .A1(n4936), .A2(n6130), .ZN(n4902) );
  INV_X1 U6216 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n4900) );
  OR2_X1 U6217 ( .A1(n4932), .A2(n4900), .ZN(n4901) );
  INV_X1 U6218 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4920) );
  XNOR2_X1 U6219 ( .A(n4921), .B(n4920), .ZN(n6403) );
  INV_X1 U6220 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6079) );
  OR2_X1 U6221 ( .A1(n8397), .A2(n6079), .ZN(n4913) );
  NAND2_X1 U6222 ( .A1(n4907), .A2(n4906), .ZN(n4910) );
  NAND2_X1 U6223 ( .A1(n4908), .A2(SI_1_), .ZN(n4909) );
  NAND2_X1 U6224 ( .A1(n4910), .A2(n4909), .ZN(n4924) );
  INV_X1 U6225 ( .A(SI_2_), .ZN(n4911) );
  XNOR2_X1 U6226 ( .A(n4924), .B(n4923), .ZN(n6078) );
  OR2_X1 U6227 ( .A1(n4982), .A2(n6078), .ZN(n4912) );
  OAI211_X1 U6228 ( .C1(n4999), .C2(n6403), .A(n4913), .B(n4912), .ZN(n6494)
         );
  INV_X1 U6229 ( .A(n9329), .ZN(n8547) );
  NAND2_X1 U6230 ( .A1(n8547), .A2(n6925), .ZN(n4914) );
  NAND2_X1 U6231 ( .A1(n6635), .A2(n4914), .ZN(n6715) );
  NAND2_X1 U6232 ( .A1(n4933), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4919) );
  INV_X1 U6233 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6134) );
  OR2_X1 U6234 ( .A1(n4936), .A2(n6134), .ZN(n4918) );
  INV_X1 U6235 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n4915) );
  OR2_X1 U6236 ( .A1(n4932), .A2(n4915), .ZN(n4917) );
  OR2_X1 U6237 ( .A1(n4989), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n4916) );
  INV_X1 U6238 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4922) );
  INV_X1 U6239 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U6240 ( .A1(n4924), .A2(n4923), .ZN(n4927) );
  NAND2_X1 U6241 ( .A1(n4925), .A2(SI_2_), .ZN(n4926) );
  NAND2_X1 U6242 ( .A1(n4927), .A2(n4926), .ZN(n4944) );
  MUX2_X1 U6243 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n4928), .Z(n4945) );
  INV_X1 U6244 ( .A(SI_3_), .ZN(n4929) );
  XNOR2_X1 U6245 ( .A(n4944), .B(n4943), .ZN(n6076) );
  OR2_X1 U6246 ( .A1(n4982), .A2(n6076), .ZN(n4930) );
  NAND2_X1 U6247 ( .A1(n7095), .A2(n7124), .ZN(n8477) );
  NAND2_X1 U6248 ( .A1(n9328), .A2(n6726), .ZN(n8485) );
  NAND2_X1 U6249 ( .A1(n7095), .A2(n6726), .ZN(n4931) );
  NAND2_X1 U6250 ( .A1(n6714), .A2(n4931), .ZN(n6788) );
  NAND2_X1 U6251 ( .A1(n5993), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n4940) );
  INV_X1 U6252 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6155) );
  OR2_X1 U6253 ( .A1(n5997), .A2(n6155), .ZN(n4939) );
  INV_X1 U6254 ( .A(n4951), .ZN(n4935) );
  INV_X1 U6255 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6632) );
  INV_X1 U6256 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6343) );
  NAND2_X1 U6257 ( .A1(n6632), .A2(n6343), .ZN(n4934) );
  NAND2_X1 U6258 ( .A1(n4935), .A2(n4934), .ZN(n7094) );
  OR2_X1 U6259 ( .A1(n4989), .A2(n7094), .ZN(n4938) );
  INV_X1 U6260 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6138) );
  OR2_X1 U6261 ( .A1(n4936), .A2(n6138), .ZN(n4937) );
  OR2_X1 U6262 ( .A1(n4941), .A2(n5181), .ZN(n4942) );
  INV_X1 U6263 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4957) );
  XNOR2_X1 U6264 ( .A(n4942), .B(n4957), .ZN(n6347) );
  INV_X1 U6265 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6085) );
  OR2_X1 U6266 ( .A1(n8397), .A2(n6085), .ZN(n4949) );
  NAND2_X1 U6267 ( .A1(n4944), .A2(n4943), .ZN(n4947) );
  NAND2_X1 U6268 ( .A1(n4945), .A2(SI_3_), .ZN(n4946) );
  NAND2_X1 U6269 ( .A1(n4947), .A2(n4946), .ZN(n4962) );
  MUX2_X1 U6270 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n6066), .Z(n4963) );
  INV_X1 U6271 ( .A(SI_4_), .ZN(n7511) );
  XNOR2_X1 U6272 ( .A(n4962), .B(n4961), .ZN(n6084) );
  OR2_X1 U6273 ( .A1(n4982), .A2(n6084), .ZN(n4948) );
  OAI211_X1 U6274 ( .C1(n4999), .C2(n6347), .A(n4949), .B(n4948), .ZN(n7098)
         );
  NAND2_X1 U6275 ( .A1(n6855), .A2(n7098), .ZN(n8298) );
  NAND2_X1 U6276 ( .A1(n9327), .A2(n6798), .ZN(n8486) );
  NAND2_X1 U6277 ( .A1(n8298), .A2(n8486), .ZN(n6792) );
  NAND2_X1 U6278 ( .A1(n6788), .A2(n6792), .ZN(n6787) );
  NAND2_X1 U6279 ( .A1(n6855), .A2(n6798), .ZN(n4950) );
  NAND2_X1 U6280 ( .A1(n4933), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n4956) );
  INV_X1 U6281 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6201) );
  OR2_X1 U6282 ( .A1(n4936), .A2(n6201), .ZN(n4955) );
  OAI21_X1 U6283 ( .B1(n4951), .B2(P1_REG3_REG_5__SCAN_IN), .A(n4970), .ZN(
        n7005) );
  OR2_X1 U6284 ( .A1(n4989), .A2(n7005), .ZN(n4954) );
  INV_X1 U6285 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n4952) );
  OR2_X1 U6286 ( .A1(n4932), .A2(n4952), .ZN(n4953) );
  NAND2_X1 U6287 ( .A1(n4941), .A2(n4957), .ZN(n4959) );
  NAND2_X1 U6288 ( .A1(n4959), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4958) );
  MUX2_X1 U6289 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4958), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n4960) );
  NAND2_X1 U6290 ( .A1(n4960), .A2(n5098), .ZN(n6202) );
  INV_X1 U6291 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6087) );
  OR2_X1 U6292 ( .A1(n8397), .A2(n6087), .ZN(n4968) );
  NAND2_X1 U6293 ( .A1(n4962), .A2(n4961), .ZN(n4965) );
  NAND2_X1 U6294 ( .A1(n4963), .A2(SI_4_), .ZN(n4964) );
  NAND2_X1 U6295 ( .A1(n4965), .A2(n4964), .ZN(n4979) );
  MUX2_X1 U6296 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6066), .Z(n4980) );
  INV_X1 U6297 ( .A(SI_5_), .ZN(n4966) );
  XNOR2_X1 U6298 ( .A(n4979), .B(n4978), .ZN(n6086) );
  OR2_X1 U6299 ( .A1(n4982), .A2(n6086), .ZN(n4967) );
  OAI211_X1 U6300 ( .C1(n4999), .C2(n6202), .A(n4968), .B(n4967), .ZN(n7007)
         );
  NAND2_X1 U6301 ( .A1(n7293), .A2(n7007), .ZN(n8479) );
  INV_X1 U6302 ( .A(n7007), .ZN(n9949) );
  NAND2_X1 U6303 ( .A1(n9326), .A2(n9949), .ZN(n8307) );
  NAND2_X1 U6304 ( .A1(n5993), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n4975) );
  INV_X1 U6305 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6212) );
  OR2_X1 U6306 ( .A1(n5997), .A2(n6212), .ZN(n4974) );
  AND2_X1 U6307 ( .A1(n4970), .A2(n4969), .ZN(n4971) );
  OR2_X1 U6308 ( .A1(n4971), .A2(n4987), .ZN(n7286) );
  OR2_X1 U6309 ( .A1(n4989), .A2(n7286), .ZN(n4973) );
  INV_X1 U6310 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6217) );
  OR2_X1 U6311 ( .A1(n4936), .A2(n6217), .ZN(n4972) );
  NAND2_X1 U6312 ( .A1(n5098), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4977) );
  INV_X1 U6313 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4976) );
  XNOR2_X1 U6314 ( .A(n4977), .B(n4976), .ZN(n6218) );
  NAND2_X1 U6315 ( .A1(n4980), .A2(SI_5_), .ZN(n4981) );
  MUX2_X1 U6316 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6066), .Z(n4997) );
  XNOR2_X1 U6317 ( .A(n4996), .B(n4994), .ZN(n6080) );
  INV_X2 U6318 ( .A(n4982), .ZN(n4998) );
  NAND2_X1 U6319 ( .A1(n6080), .A2(n4998), .ZN(n4984) );
  INV_X1 U6320 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6083) );
  OR2_X1 U6321 ( .A1(n8397), .A2(n6083), .ZN(n4983) );
  OAI211_X1 U6322 ( .C1(n4999), .C2(n6218), .A(n4984), .B(n4983), .ZN(n7288)
         );
  NAND2_X1 U6323 ( .A1(n9965), .A2(n7288), .ZN(n8480) );
  INV_X1 U6324 ( .A(n9965), .ZN(n9325) );
  INV_X1 U6325 ( .A(n7288), .ZN(n9958) );
  NAND2_X1 U6326 ( .A1(n9325), .A2(n9958), .ZN(n8312) );
  NAND2_X1 U6327 ( .A1(n8480), .A2(n8312), .ZN(n8306) );
  NAND2_X1 U6328 ( .A1(n9965), .A2(n9958), .ZN(n4985) );
  NAND2_X1 U6329 ( .A1(n7281), .A2(n4985), .ZN(n7108) );
  NAND2_X1 U6330 ( .A1(n4933), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n4993) );
  INV_X1 U6331 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n4986) );
  OR2_X1 U6332 ( .A1(n4932), .A2(n4986), .ZN(n4992) );
  NAND2_X1 U6333 ( .A1(n4987), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5020) );
  OR2_X1 U6334 ( .A1(n4987), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n4988) );
  NAND2_X1 U6335 ( .A1(n5020), .A2(n4988), .ZN(n7109) );
  OR2_X1 U6336 ( .A1(n4989), .A2(n7109), .ZN(n4991) );
  INV_X1 U6337 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7110) );
  OR2_X1 U6338 ( .A1(n4936), .A2(n7110), .ZN(n4990) );
  INV_X1 U6339 ( .A(n4994), .ZN(n4995) );
  INV_X8 U6340 ( .A(n5527), .ZN(n5376) );
  MUX2_X1 U6341 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5376), .Z(n5007) );
  XNOR2_X1 U6342 ( .A(n5006), .B(n5004), .ZN(n6088) );
  NAND2_X1 U6343 ( .A1(n6088), .A2(n4998), .ZN(n5002) );
  NOR2_X1 U6344 ( .A1(n5098), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5014) );
  OR2_X1 U6345 ( .A1(n5014), .A2(n5181), .ZN(n5000) );
  XNOR2_X1 U6346 ( .A(n5000), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6235) );
  AOI22_X1 U6347 ( .A1(n5244), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6058), .B2(
        n6235), .ZN(n5001) );
  NAND2_X1 U6348 ( .A1(n5002), .A2(n5001), .ZN(n9968) );
  NAND2_X1 U6349 ( .A1(n7292), .A2(n9968), .ZN(n8435) );
  INV_X1 U6350 ( .A(n9968), .ZN(n7114) );
  INV_X1 U6351 ( .A(n7292), .ZN(n9976) );
  NAND2_X1 U6352 ( .A1(n7114), .A2(n9976), .ZN(n8313) );
  NAND2_X1 U6353 ( .A1(n8435), .A2(n8313), .ZN(n7107) );
  NAND2_X1 U6354 ( .A1(n7108), .A2(n7107), .ZN(n7106) );
  NAND2_X1 U6355 ( .A1(n7292), .A2(n7114), .ZN(n5003) );
  NAND2_X1 U6356 ( .A1(n5007), .A2(SI_7_), .ZN(n5008) );
  INV_X1 U6357 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5009) );
  INV_X1 U6358 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6095) );
  MUX2_X1 U6359 ( .A(n5009), .B(n6095), .S(n5376), .Z(n5010) );
  INV_X1 U6360 ( .A(SI_8_), .ZN(n7569) );
  NAND2_X1 U6361 ( .A1(n5010), .A2(n7569), .ZN(n5029) );
  INV_X1 U6362 ( .A(n5010), .ZN(n5011) );
  NAND2_X1 U6363 ( .A1(n5011), .A2(SI_8_), .ZN(n5012) );
  XNOR2_X1 U6364 ( .A(n5031), .B(n5030), .ZN(n6092) );
  NAND2_X1 U6365 ( .A1(n6092), .A2(n4998), .ZN(n5017) );
  INV_X1 U6366 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5013) );
  NAND2_X1 U6367 ( .A1(n5014), .A2(n5013), .ZN(n5036) );
  NAND2_X1 U6368 ( .A1(n5036), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5015) );
  XNOR2_X1 U6369 ( .A(n5015), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6238) );
  AOI22_X1 U6370 ( .A1(n5244), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6058), .B2(
        n6238), .ZN(n5016) );
  NAND2_X1 U6371 ( .A1(n5017), .A2(n5016), .ZN(n7177) );
  NAND2_X1 U6372 ( .A1(n5993), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5026) );
  INV_X1 U6373 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5018) );
  OR2_X1 U6374 ( .A1(n5997), .A2(n5018), .ZN(n5025) );
  INV_X1 U6375 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5019) );
  NAND2_X1 U6376 ( .A1(n5020), .A2(n5019), .ZN(n5021) );
  NAND2_X1 U6377 ( .A1(n5043), .A2(n5021), .ZN(n7173) );
  OR2_X1 U6378 ( .A1(n4989), .A2(n7173), .ZN(n5024) );
  INV_X1 U6379 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5022) );
  OR2_X1 U6380 ( .A1(n4936), .A2(n5022), .ZN(n5023) );
  NAND2_X1 U6381 ( .A1(n7177), .A2(n9963), .ZN(n8319) );
  INV_X1 U6382 ( .A(n9963), .ZN(n9984) );
  NAND2_X1 U6383 ( .A1(n7177), .A2(n9984), .ZN(n5028) );
  INV_X1 U6384 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6105) );
  INV_X1 U6385 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6103) );
  MUX2_X1 U6386 ( .A(n6105), .B(n6103), .S(n5376), .Z(n5033) );
  INV_X1 U6387 ( .A(SI_9_), .ZN(n5032) );
  NAND2_X1 U6388 ( .A1(n5033), .A2(n5032), .ZN(n5054) );
  INV_X1 U6389 ( .A(n5033), .ZN(n5034) );
  NAND2_X1 U6390 ( .A1(n5034), .A2(SI_9_), .ZN(n5035) );
  XNOR2_X1 U6391 ( .A(n5053), .B(n5052), .ZN(n6102) );
  NAND2_X1 U6392 ( .A1(n6102), .A2(n4998), .ZN(n5041) );
  NAND2_X1 U6393 ( .A1(n5038), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5037) );
  MUX2_X1 U6394 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5037), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n5039) );
  NAND2_X1 U6395 ( .A1(n5039), .A2(n5075), .ZN(n9902) );
  AOI22_X1 U6396 ( .A1(n5244), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6058), .B2(
        n6240), .ZN(n5040) );
  NAND2_X1 U6397 ( .A1(n5041), .A2(n5040), .ZN(n7311) );
  NAND2_X1 U6398 ( .A1(n5042), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5050) );
  INV_X1 U6399 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7242) );
  AND2_X1 U6400 ( .A1(n5043), .A2(n7242), .ZN(n5044) );
  OR2_X1 U6401 ( .A1(n5044), .A2(n5064), .ZN(n7306) );
  OR2_X1 U6402 ( .A1(n4989), .A2(n7306), .ZN(n5049) );
  INV_X1 U6403 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5045) );
  OR2_X1 U6404 ( .A1(n5997), .A2(n5045), .ZN(n5048) );
  INV_X1 U6405 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5046) );
  OR2_X1 U6406 ( .A1(n4932), .A2(n5046), .ZN(n5047) );
  NAND4_X1 U6407 ( .A1(n5050), .A2(n5049), .A3(n5048), .A4(n5047), .ZN(n9975)
         );
  AND2_X1 U6408 ( .A1(n7311), .A2(n9975), .ZN(n5051) );
  INV_X1 U6409 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6114) );
  INV_X1 U6410 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6112) );
  MUX2_X1 U6411 ( .A(n6114), .B(n6112), .S(n5376), .Z(n5057) );
  INV_X1 U6412 ( .A(SI_10_), .ZN(n5056) );
  NAND2_X1 U6413 ( .A1(n5057), .A2(n5056), .ZN(n5073) );
  INV_X1 U6414 ( .A(n5057), .ZN(n5058) );
  NAND2_X1 U6415 ( .A1(n5058), .A2(SI_10_), .ZN(n5059) );
  XNOR2_X1 U6416 ( .A(n5072), .B(n5071), .ZN(n6111) );
  NAND2_X1 U6417 ( .A1(n6111), .A2(n4998), .ZN(n5062) );
  NAND2_X1 U6418 ( .A1(n5075), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5060) );
  XNOR2_X1 U6419 ( .A(n5060), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6450) );
  AOI22_X1 U6420 ( .A1(n5244), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6058), .B2(
        n6450), .ZN(n5061) );
  NAND2_X1 U6421 ( .A1(n5993), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5069) );
  INV_X1 U6422 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5063) );
  OR2_X1 U6423 ( .A1(n5997), .A2(n5063), .ZN(n5068) );
  INV_X1 U6424 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7388) );
  OR2_X1 U6425 ( .A1(n4936), .A2(n7388), .ZN(n5067) );
  NOR2_X1 U6426 ( .A1(n5064), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5065) );
  OR2_X1 U6427 ( .A1(n5080), .A2(n5065), .ZN(n7387) );
  OR2_X1 U6428 ( .A1(n4989), .A2(n7387), .ZN(n5066) );
  NAND2_X1 U6429 ( .A1(n9785), .A2(n7339), .ZN(n8322) );
  NAND2_X1 U6430 ( .A1(n8329), .A2(n8322), .ZN(n8439) );
  INV_X1 U6431 ( .A(n7339), .ZN(n9983) );
  OR2_X1 U6432 ( .A1(n9785), .A2(n9983), .ZN(n5070) );
  INV_X1 U6433 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5074) );
  INV_X1 U6434 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6117) );
  MUX2_X1 U6435 ( .A(n5074), .B(n6117), .S(n5376), .Z(n5089) );
  NAND2_X1 U6436 ( .A1(n6115), .A2(n4998), .ZN(n5078) );
  OAI21_X1 U6437 ( .B1(n5075), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5076) );
  XNOR2_X1 U6438 ( .A(n5076), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6451) );
  AOI22_X1 U6439 ( .A1(n5244), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6058), .B2(
        n6451), .ZN(n5077) );
  NAND2_X1 U6440 ( .A1(n5993), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5086) );
  INV_X1 U6441 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5079) );
  OR2_X1 U6442 ( .A1(n5997), .A2(n5079), .ZN(n5085) );
  OR2_X1 U6443 ( .A1(n5080), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5081) );
  NAND2_X1 U6444 ( .A1(n5103), .A2(n5081), .ZN(n9842) );
  OR2_X1 U6445 ( .A1(n4989), .A2(n9842), .ZN(n5084) );
  INV_X1 U6446 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5082) );
  OR2_X1 U6447 ( .A1(n4936), .A2(n5082), .ZN(n5083) );
  OR2_X1 U6448 ( .A1(n9845), .A2(n7794), .ZN(n7784) );
  NAND2_X1 U6449 ( .A1(n9845), .A2(n7794), .ZN(n8337) );
  INV_X1 U6450 ( .A(n7794), .ZN(n9855) );
  NAND2_X1 U6451 ( .A1(n9845), .A2(n9855), .ZN(n5087) );
  NAND2_X1 U6452 ( .A1(n9833), .A2(n5087), .ZN(n7789) );
  INV_X1 U6453 ( .A(n5089), .ZN(n5090) );
  INV_X1 U6454 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5092) );
  INV_X1 U6455 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6193) );
  MUX2_X1 U6456 ( .A(n5092), .B(n6193), .S(n5376), .Z(n5093) );
  INV_X1 U6457 ( .A(n5093), .ZN(n5094) );
  NAND2_X1 U6458 ( .A1(n5094), .A2(SI_12_), .ZN(n5095) );
  NAND2_X1 U6459 ( .A1(n5111), .A2(n5095), .ZN(n5112) );
  XNOR2_X1 U6460 ( .A(n5113), .B(n5112), .ZN(n6166) );
  NAND2_X1 U6461 ( .A1(n6166), .A2(n4998), .ZN(n5101) );
  INV_X1 U6462 ( .A(n5096), .ZN(n5097) );
  OAI21_X1 U6463 ( .B1(n5098), .B2(n5097), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5099) );
  XNOR2_X1 U6464 ( .A(n5099), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6655) );
  AOI22_X1 U6465 ( .A1(n5244), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6058), .B2(
        n6655), .ZN(n5100) );
  NAND2_X1 U6466 ( .A1(n5042), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5109) );
  INV_X1 U6467 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6443) );
  OR2_X1 U6468 ( .A1(n5997), .A2(n6443), .ZN(n5108) );
  INV_X1 U6469 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5102) );
  OR2_X2 U6470 ( .A1(n5103), .A2(n5102), .ZN(n5124) );
  NAND2_X1 U6471 ( .A1(n5103), .A2(n5102), .ZN(n5104) );
  NAND2_X1 U6472 ( .A1(n5124), .A2(n5104), .ZN(n7790) );
  OR2_X1 U6473 ( .A1(n4989), .A2(n7790), .ZN(n5107) );
  INV_X1 U6474 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5105) );
  OR2_X1 U6475 ( .A1(n4932), .A2(n5105), .ZN(n5106) );
  OR2_X1 U6476 ( .A1(n7799), .A2(n7688), .ZN(n8339) );
  NAND2_X1 U6477 ( .A1(n7799), .A2(n7688), .ZN(n8338) );
  NAND2_X1 U6478 ( .A1(n8339), .A2(n8338), .ZN(n8426) );
  NAND2_X1 U6479 ( .A1(n7789), .A2(n8426), .ZN(n7788) );
  INV_X1 U6480 ( .A(n7688), .ZN(n9838) );
  NAND2_X1 U6481 ( .A1(n7799), .A2(n9838), .ZN(n5110) );
  INV_X1 U6482 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6314) );
  INV_X1 U6483 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5114) );
  MUX2_X1 U6484 ( .A(n6314), .B(n5114), .S(n5376), .Z(n5115) );
  INV_X1 U6485 ( .A(SI_13_), .ZN(n7582) );
  NAND2_X1 U6486 ( .A1(n5115), .A2(n7582), .ZN(n5134) );
  INV_X1 U6487 ( .A(n5115), .ZN(n5116) );
  NAND2_X1 U6488 ( .A1(n5116), .A2(SI_13_), .ZN(n5117) );
  XNOR2_X1 U6489 ( .A(n5133), .B(n5132), .ZN(n6249) );
  NAND2_X1 U6490 ( .A1(n6249), .A2(n4998), .ZN(n5121) );
  NAND2_X1 U6491 ( .A1(n5118), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5119) );
  XNOR2_X1 U6492 ( .A(n5119), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7073) );
  AOI22_X1 U6493 ( .A1(n5244), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6058), .B2(
        n7073), .ZN(n5120) );
  NAND2_X1 U6494 ( .A1(n5042), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5130) );
  INV_X1 U6495 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n5122) );
  OR2_X1 U6496 ( .A1(n5997), .A2(n5122), .ZN(n5129) );
  INV_X1 U6497 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5123) );
  NAND2_X1 U6498 ( .A1(n5124), .A2(n5123), .ZN(n5125) );
  NAND2_X1 U6499 ( .A1(n5141), .A2(n5125), .ZN(n7851) );
  OR2_X1 U6500 ( .A1(n4989), .A2(n7851), .ZN(n5128) );
  INV_X1 U6501 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5126) );
  OR2_X1 U6502 ( .A1(n4932), .A2(n5126), .ZN(n5127) );
  NAND4_X1 U6503 ( .A1(n5130), .A2(n5129), .A3(n5128), .A4(n5127), .ZN(n9854)
         );
  OR2_X1 U6504 ( .A1(n7859), .A2(n9854), .ZN(n5131) );
  NAND2_X1 U6505 ( .A1(n5133), .A2(n5132), .ZN(n5135) );
  INV_X1 U6506 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6318) );
  INV_X1 U6507 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6316) );
  MUX2_X1 U6508 ( .A(n6318), .B(n6316), .S(n5376), .Z(n5149) );
  XNOR2_X1 U6509 ( .A(n5149), .B(SI_14_), .ZN(n5148) );
  XNOR2_X1 U6510 ( .A(n5153), .B(n5148), .ZN(n6315) );
  NAND2_X1 U6511 ( .A1(n6315), .A2(n4998), .ZN(n5138) );
  NAND2_X1 U6512 ( .A1(n5180), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5158) );
  XNOR2_X1 U6513 ( .A(n5158), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7220) );
  AOI22_X1 U6514 ( .A1(n5244), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6058), .B2(
        n7220), .ZN(n5137) );
  NAND2_X1 U6515 ( .A1(n5993), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5146) );
  INV_X1 U6516 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n5139) );
  OR2_X1 U6517 ( .A1(n5997), .A2(n5139), .ZN(n5145) );
  INV_X1 U6518 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5140) );
  AND2_X1 U6519 ( .A1(n5141), .A2(n5140), .ZN(n5142) );
  OR2_X1 U6520 ( .A1(n5142), .A2(n5163), .ZN(n7933) );
  OR2_X1 U6521 ( .A1(n4989), .A2(n7933), .ZN(n5144) );
  INV_X1 U6522 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7934) );
  OR2_X1 U6523 ( .A1(n4936), .A2(n7934), .ZN(n5143) );
  NAND4_X1 U6524 ( .A1(n5146), .A2(n5145), .A3(n5144), .A4(n5143), .ZN(n9615)
         );
  AND2_X1 U6525 ( .A1(n7932), .A2(n9615), .ZN(n5147) );
  INV_X1 U6526 ( .A(n5148), .ZN(n5152) );
  INV_X1 U6527 ( .A(n5149), .ZN(n5150) );
  NAND2_X1 U6528 ( .A1(n5150), .A2(SI_14_), .ZN(n5151) );
  INV_X1 U6529 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6558) );
  INV_X1 U6530 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6556) );
  MUX2_X1 U6531 ( .A(n6558), .B(n6556), .S(n5376), .Z(n5155) );
  INV_X1 U6532 ( .A(SI_15_), .ZN(n5154) );
  NAND2_X1 U6533 ( .A1(n5155), .A2(n5154), .ZN(n5171) );
  INV_X1 U6534 ( .A(n5155), .ZN(n5156) );
  NAND2_X1 U6535 ( .A1(n5156), .A2(SI_15_), .ZN(n5157) );
  NAND2_X1 U6536 ( .A1(n5171), .A2(n5157), .ZN(n5172) );
  XNOR2_X1 U6537 ( .A(n5173), .B(n5172), .ZN(n6555) );
  NAND2_X1 U6538 ( .A1(n6555), .A2(n4998), .ZN(n5162) );
  INV_X1 U6539 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5178) );
  NAND2_X1 U6540 ( .A1(n5158), .A2(n5178), .ZN(n5159) );
  NAND2_X1 U6541 ( .A1(n5159), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5160) );
  XNOR2_X1 U6542 ( .A(n5160), .B(n5177), .ZN(n7668) );
  INV_X1 U6543 ( .A(n7668), .ZN(n7224) );
  AOI22_X1 U6544 ( .A1(n5244), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6058), .B2(
        n7224), .ZN(n5161) );
  NAND2_X1 U6545 ( .A1(n5993), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5168) );
  INV_X1 U6546 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9722) );
  OR2_X1 U6547 ( .A1(n5997), .A2(n9722), .ZN(n5167) );
  NAND2_X1 U6548 ( .A1(n5163), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5187) );
  OR2_X1 U6549 ( .A1(n5163), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5164) );
  NAND2_X1 U6550 ( .A1(n5187), .A2(n5164), .ZN(n9625) );
  OR2_X1 U6551 ( .A1(n4989), .A2(n9625), .ZN(n5166) );
  INV_X1 U6552 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7217) );
  OR2_X1 U6553 ( .A1(n4936), .A2(n7217), .ZN(n5165) );
  NAND4_X1 U6554 ( .A1(n5168), .A2(n5167), .A3(n5166), .A4(n5165), .ZN(n9324)
         );
  NAND2_X1 U6555 ( .A1(n9624), .A2(n9324), .ZN(n5170) );
  NOR2_X1 U6556 ( .A1(n9624), .A2(n9324), .ZN(n5169) );
  INV_X1 U6557 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6747) );
  INV_X1 U6558 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6767) );
  MUX2_X1 U6559 ( .A(n6747), .B(n6767), .S(n5376), .Z(n5174) );
  INV_X1 U6560 ( .A(SI_16_), .ZN(n7525) );
  NAND2_X1 U6561 ( .A1(n5174), .A2(n7525), .ZN(n5195) );
  INV_X1 U6562 ( .A(n5174), .ZN(n5175) );
  NAND2_X1 U6563 ( .A1(n5175), .A2(SI_16_), .ZN(n5176) );
  XNOR2_X1 U6564 ( .A(n5194), .B(n5193), .ZN(n6746) );
  NAND2_X1 U6565 ( .A1(n6746), .A2(n4998), .ZN(n5184) );
  NAND2_X1 U6566 ( .A1(n5178), .A2(n5177), .ZN(n5179) );
  NOR2_X2 U6567 ( .A1(n5180), .A2(n5179), .ZN(n5197) );
  OR2_X1 U6568 ( .A1(n5197), .A2(n5181), .ZN(n5182) );
  XNOR2_X1 U6569 ( .A(n5182), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9355) );
  AOI22_X1 U6570 ( .A1(n5244), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6058), .B2(
        n9355), .ZN(n5183) );
  NAND2_X1 U6571 ( .A1(n4933), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5192) );
  INV_X1 U6572 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n5185) );
  OR2_X1 U6573 ( .A1(n4932), .A2(n5185), .ZN(n5191) );
  INV_X1 U6574 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6575 ( .A1(n5187), .A2(n5186), .ZN(n5188) );
  NAND2_X1 U6576 ( .A1(n5204), .A2(n5188), .ZN(n9599) );
  OR2_X1 U6577 ( .A1(n4989), .A2(n9599), .ZN(n5190) );
  INV_X1 U6578 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9600) );
  OR2_X1 U6579 ( .A1(n4936), .A2(n9600), .ZN(n5189) );
  OR2_X1 U6580 ( .A1(n9715), .A2(n9586), .ZN(n8351) );
  NAND2_X1 U6581 ( .A1(n9715), .A2(n9586), .ZN(n8502) );
  NAND2_X1 U6582 ( .A1(n8351), .A2(n8502), .ZN(n9593) );
  MUX2_X1 U6583 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n5376), .Z(n5212) );
  INV_X1 U6584 ( .A(SI_17_), .ZN(n7479) );
  XNOR2_X1 U6585 ( .A(n5212), .B(n7479), .ZN(n5211) );
  XNOR2_X1 U6586 ( .A(n5214), .B(n5211), .ZN(n6743) );
  NAND2_X1 U6587 ( .A1(n6743), .A2(n4998), .ZN(n5202) );
  INV_X1 U6588 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U6589 ( .A1(n5240), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5199) );
  NAND2_X1 U6590 ( .A1(n5199), .A2(n5198), .ZN(n5215) );
  OR2_X1 U6591 ( .A1(n5199), .A2(n5198), .ZN(n5200) );
  AND2_X1 U6592 ( .A1(n5215), .A2(n5200), .ZN(n9367) );
  AOI22_X1 U6593 ( .A1(n5244), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6058), .B2(
        n9367), .ZN(n5201) );
  INV_X1 U6594 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5203) );
  AND2_X1 U6595 ( .A1(n5204), .A2(n5203), .ZN(n5205) );
  OR2_X1 U6596 ( .A1(n5205), .A2(n5219), .ZN(n9579) );
  INV_X1 U6597 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n5206) );
  OR2_X1 U6598 ( .A1(n5997), .A2(n5206), .ZN(n5208) );
  INV_X1 U6599 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9580) );
  OR2_X1 U6600 ( .A1(n4936), .A2(n9580), .ZN(n5207) );
  AND2_X1 U6601 ( .A1(n5208), .A2(n5207), .ZN(n5210) );
  NAND2_X1 U6602 ( .A1(n5993), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5209) );
  OAI211_X1 U6603 ( .C1(n9579), .C2(n4989), .A(n5210), .B(n5209), .ZN(n9604)
         );
  OR2_X1 U6604 ( .A1(n9706), .A2(n9604), .ZN(n5225) );
  AND2_X1 U6605 ( .A1(n9593), .A2(n5225), .ZN(n9558) );
  INV_X1 U6606 ( .A(n5211), .ZN(n5213) );
  MUX2_X1 U6607 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5376), .Z(n5234) );
  XNOR2_X1 U6608 ( .A(n5234), .B(SI_18_), .ZN(n5231) );
  NAND2_X1 U6609 ( .A1(n6974), .A2(n4998), .ZN(n5218) );
  NAND2_X1 U6610 ( .A1(n5215), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5216) );
  XNOR2_X1 U6611 ( .A(n5216), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9368) );
  AOI22_X1 U6612 ( .A1(n5244), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6058), .B2(
        n9368), .ZN(n5217) );
  OR2_X1 U6613 ( .A1(n5219), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5220) );
  NAND2_X1 U6614 ( .A1(n5219), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5247) );
  AND2_X1 U6615 ( .A1(n5220), .A2(n5247), .ZN(n9557) );
  NAND2_X1 U6616 ( .A1(n9557), .A2(n5328), .ZN(n5223) );
  AOI22_X1 U6617 ( .A1(n4933), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n5993), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5222) );
  INV_X1 U6618 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9567) );
  OR2_X1 U6619 ( .A1(n4936), .A2(n9567), .ZN(n5221) );
  AND3_X1 U6620 ( .A1(n5223), .A2(n5222), .A3(n5221), .ZN(n9690) );
  OR2_X1 U6621 ( .A1(n9566), .A2(n9690), .ZN(n8356) );
  NAND2_X1 U6622 ( .A1(n9566), .A2(n9690), .ZN(n8359) );
  NAND2_X1 U6623 ( .A1(n8356), .A2(n8359), .ZN(n8425) );
  AND2_X1 U6624 ( .A1(n9558), .A2(n8425), .ZN(n5224) );
  NAND2_X1 U6625 ( .A1(n9594), .A2(n5224), .ZN(n9537) );
  INV_X1 U6626 ( .A(n8425), .ZN(n5228) );
  INV_X1 U6627 ( .A(n5225), .ZN(n5226) );
  INV_X1 U6628 ( .A(n9586), .ZN(n9616) );
  NAND2_X1 U6629 ( .A1(n9715), .A2(n9616), .ZN(n9572) );
  OR2_X1 U6630 ( .A1(n5226), .A2(n9572), .ZN(n9559) );
  NAND2_X1 U6631 ( .A1(n9706), .A2(n9604), .ZN(n9561) );
  AND2_X1 U6632 ( .A1(n9559), .A2(n9561), .ZN(n5227) );
  OR2_X1 U6633 ( .A1(n5228), .A2(n5227), .ZN(n5230) );
  INV_X1 U6634 ( .A(n9690), .ZN(n9323) );
  NAND2_X1 U6635 ( .A1(n9566), .A2(n9323), .ZN(n5229) );
  INV_X1 U6636 ( .A(n5231), .ZN(n5232) );
  NAND2_X1 U6637 ( .A1(n5233), .A2(n5232), .ZN(n5236) );
  NAND2_X1 U6638 ( .A1(n5234), .A2(SI_18_), .ZN(n5235) );
  INV_X1 U6639 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7121) );
  INV_X1 U6640 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7119) );
  MUX2_X1 U6641 ( .A(n7121), .B(n7119), .S(n5376), .Z(n5237) );
  NAND2_X1 U6642 ( .A1(n5237), .A2(n7596), .ZN(n5258) );
  INV_X1 U6643 ( .A(n5237), .ZN(n5238) );
  NAND2_X1 U6644 ( .A1(n5238), .A2(SI_19_), .ZN(n5239) );
  NAND2_X1 U6645 ( .A1(n5258), .A2(n5239), .ZN(n5257) );
  XNOR2_X1 U6646 ( .A(n5256), .B(n5257), .ZN(n7118) );
  NAND2_X1 U6647 ( .A1(n7118), .A2(n4998), .ZN(n5246) );
  NAND2_X1 U6648 ( .A1(n4364), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5241) );
  MUX2_X1 U6649 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5241), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n5243) );
  INV_X1 U6650 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5242) );
  NAND2_X1 U6651 ( .A1(n5243), .A2(n5404), .ZN(n9408) );
  AOI22_X1 U6652 ( .A1(n5244), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9513), .B2(
        n6058), .ZN(n5245) );
  NAND2_X1 U6653 ( .A1(n5993), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5252) );
  INV_X1 U6654 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9369) );
  OR2_X1 U6655 ( .A1(n5997), .A2(n9369), .ZN(n5251) );
  OAI21_X1 U6656 ( .B1(P1_REG3_REG_19__SCAN_IN), .B2(n5248), .A(n5265), .ZN(
        n9540) );
  OR2_X1 U6657 ( .A1(n4989), .A2(n9540), .ZN(n5250) );
  INV_X1 U6658 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9541) );
  OR2_X1 U6659 ( .A1(n4936), .A2(n9541), .ZN(n5249) );
  NAND4_X1 U6660 ( .A1(n5252), .A2(n5251), .A3(n5250), .A4(n5249), .ZN(n9681)
         );
  NAND2_X1 U6661 ( .A1(n9537), .A2(n5253), .ZN(n5255) );
  OR2_X1 U6662 ( .A1(n9752), .A2(n9681), .ZN(n5254) );
  INV_X1 U6663 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7163) );
  INV_X1 U6664 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7160) );
  MUX2_X1 U6665 ( .A(n7163), .B(n7160), .S(n5376), .Z(n5260) );
  INV_X1 U6666 ( .A(SI_20_), .ZN(n5259) );
  NAND2_X1 U6667 ( .A1(n5260), .A2(n5259), .ZN(n5275) );
  INV_X1 U6668 ( .A(n5260), .ZN(n5261) );
  NAND2_X1 U6669 ( .A1(n5261), .A2(SI_20_), .ZN(n5262) );
  AND2_X1 U6670 ( .A1(n5275), .A2(n5262), .ZN(n5273) );
  XNOR2_X1 U6671 ( .A(n5274), .B(n5273), .ZN(n7159) );
  NAND2_X1 U6672 ( .A1(n7159), .A2(n4998), .ZN(n5264) );
  OR2_X1 U6673 ( .A1(n8397), .A2(n7160), .ZN(n5263) );
  NAND2_X1 U6674 ( .A1(n5993), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5270) );
  INV_X1 U6675 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9688) );
  OR2_X1 U6676 ( .A1(n5997), .A2(n9688), .ZN(n5269) );
  OAI21_X1 U6677 ( .B1(P1_REG3_REG_20__SCAN_IN), .B2(n5266), .A(n5280), .ZN(
        n9522) );
  OR2_X1 U6678 ( .A1(n4989), .A2(n9522), .ZN(n5268) );
  INV_X1 U6679 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9523) );
  OR2_X1 U6680 ( .A1(n4936), .A2(n9523), .ZN(n5267) );
  NAND4_X1 U6681 ( .A1(n5270), .A2(n5269), .A3(n5268), .A4(n5267), .ZN(n9543)
         );
  NOR2_X1 U6682 ( .A1(n9533), .A2(n9543), .ZN(n5272) );
  NAND2_X1 U6683 ( .A1(n9533), .A2(n9543), .ZN(n5271) );
  NAND2_X1 U6684 ( .A1(n5274), .A2(n5273), .ZN(n5276) );
  MUX2_X1 U6685 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n5376), .Z(n5288) );
  INV_X1 U6686 ( .A(SI_21_), .ZN(n5277) );
  XNOR2_X1 U6687 ( .A(n5288), .B(n5277), .ZN(n5287) );
  XNOR2_X1 U6688 ( .A(n5291), .B(n5287), .ZN(n7164) );
  NAND2_X1 U6689 ( .A1(n7164), .A2(n4998), .ZN(n5279) );
  INV_X1 U6690 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7165) );
  OR2_X1 U6691 ( .A1(n8397), .A2(n7165), .ZN(n5278) );
  NAND2_X1 U6692 ( .A1(n4933), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5286) );
  INV_X1 U6693 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9743) );
  OR2_X1 U6694 ( .A1(n4932), .A2(n9743), .ZN(n5285) );
  INV_X1 U6695 ( .A(n5280), .ZN(n5282) );
  INV_X1 U6696 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9252) );
  INV_X1 U6697 ( .A(n5297), .ZN(n5281) );
  OAI21_X1 U6698 ( .B1(P1_REG3_REG_21__SCAN_IN), .B2(n5282), .A(n5281), .ZN(
        n9512) );
  OR2_X1 U6699 ( .A1(n4989), .A2(n9512), .ZN(n5284) );
  INV_X1 U6700 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9500) );
  OR2_X1 U6701 ( .A1(n4936), .A2(n9500), .ZN(n5283) );
  NAND2_X1 U6702 ( .A1(n9502), .A2(n9528), .ZN(n8364) );
  INV_X1 U6703 ( .A(n9528), .ZN(n9682) );
  INV_X1 U6704 ( .A(n5287), .ZN(n5290) );
  NAND2_X1 U6705 ( .A1(n5288), .A2(SI_21_), .ZN(n5289) );
  INV_X1 U6706 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8018) );
  INV_X1 U6707 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7400) );
  MUX2_X1 U6708 ( .A(n8018), .B(n7400), .S(n5376), .Z(n5292) );
  INV_X1 U6709 ( .A(SI_22_), .ZN(n7581) );
  NAND2_X1 U6710 ( .A1(n5292), .A2(n7581), .ZN(n5302) );
  INV_X1 U6711 ( .A(n5292), .ZN(n5293) );
  NAND2_X1 U6712 ( .A1(n5293), .A2(SI_22_), .ZN(n5294) );
  NAND2_X1 U6713 ( .A1(n5302), .A2(n5294), .ZN(n5303) );
  XNOR2_X1 U6714 ( .A(n5304), .B(n5303), .ZN(n7398) );
  NAND2_X1 U6715 ( .A1(n7398), .A2(n4998), .ZN(n5296) );
  OR2_X1 U6716 ( .A1(n8397), .A2(n7400), .ZN(n5295) );
  NAND2_X1 U6717 ( .A1(n5993), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5301) );
  INV_X1 U6718 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9673) );
  OR2_X1 U6719 ( .A1(n5997), .A2(n9673), .ZN(n5300) );
  NAND2_X1 U6720 ( .A1(n5297), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5311) );
  OAI21_X1 U6721 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n5297), .A(n5311), .ZN(
        n9492) );
  OR2_X1 U6722 ( .A1(n4989), .A2(n9492), .ZN(n5299) );
  INV_X1 U6723 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9493) );
  OR2_X1 U6724 ( .A1(n4936), .A2(n9493), .ZN(n5298) );
  NAND4_X1 U6725 ( .A1(n5301), .A2(n5300), .A3(n5299), .A4(n5298), .ZN(n9510)
         );
  INV_X1 U6726 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5305) );
  INV_X1 U6727 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7662) );
  MUX2_X1 U6728 ( .A(n5305), .B(n7662), .S(n5376), .Z(n5306) );
  INV_X1 U6729 ( .A(SI_23_), .ZN(n7579) );
  NAND2_X1 U6730 ( .A1(n5306), .A2(n7579), .ZN(n5322) );
  INV_X1 U6731 ( .A(n5306), .ZN(n5307) );
  NAND2_X1 U6732 ( .A1(n5307), .A2(SI_23_), .ZN(n5308) );
  AND2_X1 U6733 ( .A1(n5322), .A2(n5308), .ZN(n5320) );
  NAND2_X1 U6734 ( .A1(n7659), .A2(n4998), .ZN(n5310) );
  OR2_X1 U6735 ( .A1(n8397), .A2(n7662), .ZN(n5309) );
  OAI21_X1 U6736 ( .B1(n5312), .B2(P1_REG3_REG_23__SCAN_IN), .A(n5327), .ZN(
        n9476) );
  INV_X1 U6737 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U6738 ( .A1(n5993), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U6739 ( .A1(n5042), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5313) );
  OAI211_X1 U6740 ( .C1(n5997), .C2(n5315), .A(n5314), .B(n5313), .ZN(n5316)
         );
  INV_X1 U6741 ( .A(n5316), .ZN(n5317) );
  OAI21_X1 U6742 ( .B1(n9476), .B2(n4989), .A(n5317), .ZN(n9657) );
  NOR2_X1 U6743 ( .A1(n9667), .A2(n9657), .ZN(n5319) );
  NAND2_X1 U6744 ( .A1(n9667), .A2(n9657), .ZN(n5318) );
  NAND2_X1 U6745 ( .A1(n5321), .A2(n5320), .ZN(n5323) );
  NAND2_X1 U6746 ( .A1(n5323), .A2(n5322), .ZN(n5341) );
  INV_X1 U6747 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7741) );
  INV_X1 U6748 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7739) );
  MUX2_X1 U6749 ( .A(n7741), .B(n7739), .S(n5376), .Z(n5337) );
  XNOR2_X1 U6750 ( .A(n5337), .B(SI_24_), .ZN(n5336) );
  XNOR2_X1 U6751 ( .A(n5341), .B(n5336), .ZN(n7738) );
  NAND2_X1 U6752 ( .A1(n7738), .A2(n4998), .ZN(n5325) );
  OR2_X1 U6753 ( .A1(n8397), .A2(n7739), .ZN(n5324) );
  INV_X1 U6754 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9269) );
  INV_X1 U6755 ( .A(n5327), .ZN(n5326) );
  NAND2_X1 U6756 ( .A1(n5326), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5348) );
  INV_X1 U6757 ( .A(n5348), .ZN(n5349) );
  AOI21_X1 U6758 ( .B1(n5327), .B2(n9269), .A(n5349), .ZN(n9462) );
  NAND2_X1 U6759 ( .A1(n9462), .A2(n5328), .ZN(n5334) );
  INV_X1 U6760 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5331) );
  NAND2_X1 U6761 ( .A1(n5993), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5330) );
  NAND2_X1 U6762 ( .A1(n5042), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5329) );
  OAI211_X1 U6763 ( .C1(n5997), .C2(n5331), .A(n5330), .B(n5329), .ZN(n5332)
         );
  INV_X1 U6764 ( .A(n5332), .ZN(n5333) );
  NAND2_X1 U6765 ( .A1(n5334), .A2(n5333), .ZN(n9648) );
  OR2_X1 U6766 ( .A1(n9454), .A2(n9648), .ZN(n5335) );
  INV_X1 U6767 ( .A(n5336), .ZN(n5340) );
  INV_X1 U6768 ( .A(n5337), .ZN(n5338) );
  NAND2_X1 U6769 ( .A1(n5338), .A2(SI_24_), .ZN(n5339) );
  INV_X1 U6770 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7843) );
  INV_X1 U6771 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7847) );
  MUX2_X1 U6772 ( .A(n7843), .B(n7847), .S(n5376), .Z(n5342) );
  INV_X1 U6773 ( .A(SI_25_), .ZN(n7564) );
  NAND2_X1 U6774 ( .A1(n5342), .A2(n7564), .ZN(n5356) );
  INV_X1 U6775 ( .A(n5342), .ZN(n5343) );
  NAND2_X1 U6776 ( .A1(n5343), .A2(SI_25_), .ZN(n5344) );
  NAND2_X1 U6777 ( .A1(n5356), .A2(n5344), .ZN(n5357) );
  XNOR2_X1 U6778 ( .A(n5358), .B(n5357), .ZN(n7841) );
  NAND2_X1 U6779 ( .A1(n7841), .A2(n4998), .ZN(n5346) );
  OR2_X1 U6780 ( .A1(n8397), .A2(n7847), .ZN(n5345) );
  NAND2_X1 U6781 ( .A1(n4933), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5354) );
  INV_X1 U6782 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9442) );
  OR2_X1 U6783 ( .A1(n4936), .A2(n9442), .ZN(n5353) );
  INV_X1 U6784 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5347) );
  NOR2_X2 U6785 ( .A1(n5348), .A2(n5347), .ZN(n5367) );
  OAI21_X1 U6786 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n5349), .A(n5365), .ZN(
        n9441) );
  OR2_X1 U6787 ( .A1(n4989), .A2(n9441), .ZN(n5352) );
  INV_X1 U6788 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n5350) );
  OR2_X1 U6789 ( .A1(n4932), .A2(n5350), .ZN(n5351) );
  INV_X1 U6790 ( .A(n9419), .ZN(n9656) );
  INV_X1 U6791 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7918) );
  INV_X1 U6792 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7902) );
  MUX2_X1 U6793 ( .A(n7918), .B(n7902), .S(n5376), .Z(n5359) );
  NAND2_X1 U6794 ( .A1(n5359), .A2(n7554), .ZN(n5374) );
  INV_X1 U6795 ( .A(n5359), .ZN(n5360) );
  NAND2_X1 U6796 ( .A1(n5360), .A2(SI_26_), .ZN(n5361) );
  AND2_X1 U6797 ( .A1(n5374), .A2(n5361), .ZN(n5372) );
  OR2_X1 U6798 ( .A1(n8397), .A2(n7902), .ZN(n5362) );
  NAND2_X1 U6799 ( .A1(n5993), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5371) );
  INV_X1 U6800 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9645) );
  OR2_X1 U6801 ( .A1(n5997), .A2(n9645), .ZN(n5370) );
  INV_X1 U6802 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5364) );
  INV_X1 U6803 ( .A(n5384), .ZN(n5366) );
  OAI21_X1 U6804 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n5367), .A(n5366), .ZN(
        n9428) );
  OR2_X1 U6805 ( .A1(n4989), .A2(n9428), .ZN(n5369) );
  INV_X1 U6806 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9429) );
  OR2_X1 U6807 ( .A1(n4936), .A2(n9429), .ZN(n5368) );
  NAND4_X1 U6808 ( .A1(n5371), .A2(n5370), .A3(n5369), .A4(n5368), .ZN(n9647)
         );
  NAND2_X1 U6809 ( .A1(n5373), .A2(n5372), .ZN(n5375) );
  INV_X1 U6810 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5377) );
  INV_X1 U6811 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7943) );
  MUX2_X1 U6812 ( .A(n5377), .B(n7943), .S(n5376), .Z(n5379) );
  INV_X1 U6813 ( .A(SI_27_), .ZN(n5378) );
  NAND2_X1 U6814 ( .A1(n5379), .A2(n5378), .ZN(n5393) );
  INV_X1 U6815 ( .A(n5379), .ZN(n5380) );
  NAND2_X1 U6816 ( .A1(n5380), .A2(SI_27_), .ZN(n5381) );
  AND2_X1 U6817 ( .A1(n5393), .A2(n5381), .ZN(n5391) );
  OR2_X1 U6818 ( .A1(n8397), .A2(n7943), .ZN(n5382) );
  NAND2_X1 U6819 ( .A1(n4933), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5389) );
  INV_X1 U6820 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n5506) );
  OR2_X1 U6821 ( .A1(n4932), .A2(n5506), .ZN(n5388) );
  NAND2_X1 U6822 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n5384), .ZN(n5435) );
  OAI21_X1 U6823 ( .B1(P1_REG3_REG_27__SCAN_IN), .B2(n5384), .A(n5435), .ZN(
        n9405) );
  OR2_X1 U6824 ( .A1(n4989), .A2(n9405), .ZN(n5387) );
  INV_X1 U6825 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5385) );
  OR2_X1 U6826 ( .A1(n4936), .A2(n5385), .ZN(n5386) );
  OAI22_X1 U6827 ( .A1(n5493), .A2(n8571), .B1(n9395), .B2(n5390), .ZN(n5402)
         );
  MUX2_X1 U6828 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n5376), .Z(n5897) );
  INV_X1 U6829 ( .A(SI_28_), .ZN(n5898) );
  XNOR2_X1 U6830 ( .A(n5897), .B(n5898), .ZN(n5895) );
  INV_X1 U6831 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8016) );
  OR2_X1 U6832 ( .A1(n8397), .A2(n8016), .ZN(n5395) );
  NAND2_X1 U6833 ( .A1(n5993), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5401) );
  INV_X1 U6834 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5488) );
  OR2_X1 U6835 ( .A1(n5997), .A2(n5488), .ZN(n5400) );
  INV_X1 U6836 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5397) );
  XNOR2_X1 U6837 ( .A(n5435), .B(n5397), .ZN(n9392) );
  OR2_X1 U6838 ( .A1(n4989), .A2(n9392), .ZN(n5399) );
  INV_X1 U6839 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9393) );
  OR2_X1 U6840 ( .A1(n4936), .A2(n9393), .ZN(n5398) );
  NAND2_X1 U6841 ( .A1(n5402), .A2(n8395), .ZN(n5403) );
  INV_X1 U6842 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5407) );
  NAND2_X1 U6843 ( .A1(n5408), .A2(n5407), .ZN(n5405) );
  INV_X1 U6844 ( .A(n8591), .ZN(n7399) );
  NAND2_X2 U6845 ( .A1(n7399), .A2(n9513), .ZN(n8415) );
  XNOR2_X1 U6846 ( .A(n5408), .B(n5407), .ZN(n8583) );
  INV_X1 U6847 ( .A(n8583), .ZN(n6837) );
  INV_X1 U6848 ( .A(n9787), .ZN(n9954) );
  XNOR2_X2 U6849 ( .A(n5409), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5410) );
  AND2_X2 U6850 ( .A1(n5410), .A2(n8583), .ZN(n7279) );
  OR2_X1 U6851 ( .A1(n6419), .A2(n7279), .ZN(n5412) );
  NAND3_X1 U6852 ( .A1(n7399), .A2(n5410), .A3(n5477), .ZN(n5411) );
  NAND2_X1 U6853 ( .A1(n5412), .A2(n5411), .ZN(n9860) );
  INV_X1 U6854 ( .A(n9932), .ZN(n8427) );
  INV_X1 U6855 ( .A(n8428), .ZN(n6830) );
  INV_X1 U6856 ( .A(n6423), .ZN(n6508) );
  NAND2_X1 U6857 ( .A1(n6508), .A2(n6839), .ZN(n5413) );
  OAI21_X2 U6858 ( .B1(n6827), .B2(n6830), .A(n5413), .ZN(n8549) );
  NAND2_X1 U6859 ( .A1(n8549), .A2(n6638), .ZN(n5414) );
  NAND2_X1 U6860 ( .A1(n8547), .A2(n6494), .ZN(n8546) );
  NAND2_X1 U6861 ( .A1(n5414), .A2(n8546), .ZN(n6720) );
  NAND2_X1 U6862 ( .A1(n6720), .A2(n8430), .ZN(n5415) );
  AND2_X1 U6863 ( .A1(n8479), .A2(n8298), .ZN(n8303) );
  AND2_X1 U6864 ( .A1(n8303), .A2(n8480), .ZN(n8551) );
  INV_X1 U6865 ( .A(n8307), .ZN(n5416) );
  NAND2_X1 U6866 ( .A1(n8480), .A2(n5416), .ZN(n8483) );
  AND2_X1 U6867 ( .A1(n8483), .A2(n8312), .ZN(n5417) );
  INV_X1 U6868 ( .A(n9975), .ZN(n7087) );
  OR2_X1 U6869 ( .A1(n7311), .A2(n7087), .ZN(n8324) );
  NAND2_X1 U6870 ( .A1(n8329), .A2(n8324), .ZN(n8491) );
  NAND2_X1 U6871 ( .A1(n7311), .A2(n7087), .ZN(n8320) );
  NAND2_X1 U6872 ( .A1(n8322), .A2(n8320), .ZN(n8325) );
  NAND2_X1 U6873 ( .A1(n8325), .A2(n8329), .ZN(n8471) );
  NAND2_X1 U6874 ( .A1(n5418), .A2(n8337), .ZN(n7785) );
  AND2_X1 U6875 ( .A1(n8339), .A2(n7784), .ZN(n8334) );
  INV_X1 U6876 ( .A(n9854), .ZN(n7778) );
  OR2_X1 U6877 ( .A1(n7859), .A2(n7778), .ZN(n8344) );
  NAND2_X1 U6878 ( .A1(n7859), .A2(n7778), .ZN(n8336) );
  INV_X1 U6879 ( .A(n9615), .ZN(n7855) );
  NAND2_X1 U6880 ( .A1(n7932), .A2(n7855), .ZN(n8345) );
  NAND2_X1 U6881 ( .A1(n8495), .A2(n8345), .ZN(n8445) );
  INV_X1 U6882 ( .A(n8336), .ZN(n5419) );
  NOR2_X1 U6883 ( .A1(n8445), .A2(n5419), .ZN(n5420) );
  NAND2_X1 U6884 ( .A1(n7924), .A2(n8495), .ZN(n9614) );
  INV_X1 U6885 ( .A(n9324), .ZN(n9711) );
  NAND2_X1 U6886 ( .A1(n9624), .A2(n9711), .ZN(n8498) );
  OR2_X1 U6887 ( .A1(n9624), .A2(n9711), .ZN(n9590) );
  AND2_X1 U6888 ( .A1(n8351), .A2(n9590), .ZN(n8501) );
  INV_X1 U6889 ( .A(n9604), .ZN(n9712) );
  NAND2_X1 U6890 ( .A1(n5421), .A2(n4833), .ZN(n9553) );
  OR2_X1 U6891 ( .A1(n9706), .A2(n9712), .ZN(n9552) );
  AND2_X1 U6892 ( .A1(n8356), .A2(n9552), .ZN(n8514) );
  INV_X1 U6893 ( .A(n9681), .ZN(n9556) );
  OR2_X1 U6894 ( .A1(n9752), .A2(n9556), .ZN(n8357) );
  NAND2_X1 U6895 ( .A1(n9752), .A2(n9556), .ZN(n8509) );
  INV_X1 U6896 ( .A(n9519), .ZN(n5423) );
  NOR2_X1 U6897 ( .A1(n9504), .A2(n9505), .ZN(n5425) );
  INV_X1 U6898 ( .A(n9510), .ZN(n9253) );
  OR2_X1 U6899 ( .A1(n9491), .A2(n9253), .ZN(n8518) );
  NAND2_X1 U6900 ( .A1(n9491), .A2(n9253), .ZN(n8423) );
  INV_X1 U6901 ( .A(n9657), .ZN(n9452) );
  NAND2_X1 U6902 ( .A1(n9667), .A2(n9452), .ZN(n8370) );
  NAND2_X1 U6903 ( .A1(n8519), .A2(n8370), .ZN(n8422) );
  NAND2_X1 U6904 ( .A1(n9470), .A2(n8519), .ZN(n9457) );
  INV_X1 U6905 ( .A(n9648), .ZN(n8643) );
  XNOR2_X1 U6906 ( .A(n9454), .B(n8643), .ZN(n9456) );
  NOR2_X1 U6907 ( .A1(n9457), .A2(n9456), .ZN(n9455) );
  NAND2_X1 U6908 ( .A1(n9454), .A2(n8643), .ZN(n8372) );
  INV_X1 U6909 ( .A(n8372), .ZN(n5426) );
  NAND2_X1 U6910 ( .A1(n9438), .A2(n8567), .ZN(n9415) );
  INV_X1 U6911 ( .A(n9647), .ZN(n9440) );
  NAND2_X1 U6912 ( .A1(n9415), .A2(n8525), .ZN(n5427) );
  NAND2_X1 U6913 ( .A1(n9427), .A2(n9440), .ZN(n8421) );
  NAND2_X1 U6914 ( .A1(n5427), .A2(n8421), .ZN(n5496) );
  NAND2_X1 U6915 ( .A1(n5497), .A2(n8526), .ZN(n5428) );
  NAND2_X1 U6916 ( .A1(n5428), .A2(n8450), .ZN(n5430) );
  INV_X1 U6917 ( .A(n8526), .ZN(n8380) );
  NOR2_X1 U6918 ( .A1(n8450), .A2(n8380), .ZN(n5429) );
  NAND2_X1 U6919 ( .A1(n5430), .A2(n5990), .ZN(n9390) );
  NAND2_X1 U6920 ( .A1(n8591), .A2(n9513), .ZN(n5432) );
  NAND2_X1 U6921 ( .A1(n5410), .A2(n6837), .ZN(n5431) );
  NAND2_X1 U6922 ( .A1(n5432), .A2(n5431), .ZN(n9693) );
  NAND2_X1 U6923 ( .A1(n9390), .A2(n9693), .ZN(n5446) );
  NAND2_X1 U6924 ( .A1(n8591), .A2(n5410), .ZN(n8460) );
  OR2_X1 U6925 ( .A1(n8460), .A2(n5433), .ZN(n9964) );
  NAND2_X1 U6926 ( .A1(n4933), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5440) );
  INV_X1 U6927 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n5434) );
  OR2_X1 U6928 ( .A1(n4936), .A2(n5434), .ZN(n5439) );
  INV_X1 U6929 ( .A(n5435), .ZN(n5436) );
  NAND2_X1 U6930 ( .A1(n5436), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8021) );
  OR2_X1 U6931 ( .A1(n4989), .A2(n8021), .ZN(n5438) );
  INV_X1 U6932 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6051) );
  OR2_X1 U6933 ( .A1(n4932), .A2(n6051), .ZN(n5437) );
  INV_X1 U6934 ( .A(n5433), .ZN(n6147) );
  OR2_X1 U6935 ( .A1(n8460), .A2(n6147), .ZN(n9962) );
  OAI22_X1 U6936 ( .A1(n9418), .A2(n9964), .B1(n9397), .B2(n9962), .ZN(n5441)
         );
  INV_X1 U6937 ( .A(n5441), .ZN(n5445) );
  NAND2_X1 U6938 ( .A1(n6858), .A2(n9949), .ZN(n7283) );
  INV_X1 U6939 ( .A(n7311), .ZN(n9989) );
  NAND2_X1 U6940 ( .A1(n7305), .A2(n9989), .ZN(n7385) );
  INV_X1 U6941 ( .A(n5443), .ZN(n7384) );
  INV_X1 U6942 ( .A(n7799), .ZN(n7795) );
  INV_X1 U6943 ( .A(n7859), .ZN(n7952) );
  INV_X1 U6944 ( .A(n9715), .ZN(n9607) );
  INV_X1 U6945 ( .A(n9706), .ZN(n9578) );
  NAND2_X1 U6946 ( .A1(n9574), .A2(n9578), .ZN(n9575) );
  INV_X1 U6947 ( .A(n9502), .ZN(n9745) );
  INV_X1 U6948 ( .A(n5410), .ZN(n8458) );
  AND2_X1 U6949 ( .A1(n7399), .A2(n8458), .ZN(n9931) );
  AND2_X1 U6950 ( .A1(n9931), .A2(n8583), .ZN(n9847) );
  OAI211_X1 U6951 ( .C1(n8720), .C2(n4340), .A(n9847), .B(n6000), .ZN(n9398)
         );
  NAND3_X1 U6952 ( .A1(n5446), .A2(n5445), .A3(n9398), .ZN(n5447) );
  AOI21_X1 U6953 ( .B1(n9391), .B2(n9992), .A(n5447), .ZN(n5487) );
  OR2_X1 U6954 ( .A1(n8460), .A2(n5477), .ZN(n6625) );
  NAND2_X1 U6955 ( .A1(n4351), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5448) );
  MUX2_X1 U6956 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5448), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n5449) );
  INV_X1 U6957 ( .A(n7903), .ZN(n5461) );
  NAND2_X1 U6958 ( .A1(n5450), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5451) );
  MUX2_X1 U6959 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5451), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5452) );
  NAND2_X1 U6960 ( .A1(n5452), .A2(n4351), .ZN(n7844) );
  NAND2_X1 U6961 ( .A1(n4363), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5454) );
  XNOR2_X1 U6962 ( .A(n5454), .B(n5453), .ZN(n7740) );
  NOR2_X1 U6963 ( .A1(n7844), .A2(n7740), .ZN(n5455) );
  NAND2_X1 U6964 ( .A1(n5456), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5457) );
  XNOR2_X1 U6965 ( .A(n5457), .B(n4735), .ZN(n7660) );
  AND2_X1 U6966 ( .A1(n7660), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6074) );
  AND2_X1 U6967 ( .A1(n6624), .A2(n6074), .ZN(n6355) );
  OR2_X1 U6968 ( .A1(n9787), .A2(n5410), .ZN(n5458) );
  NAND2_X1 U6969 ( .A1(n7844), .A2(P1_B_REG_SCAN_IN), .ZN(n5460) );
  INV_X1 U6970 ( .A(n7740), .ZN(n5459) );
  MUX2_X1 U6971 ( .A(n5460), .B(P1_B_REG_SCAN_IN), .S(n5459), .Z(n5462) );
  NAND2_X1 U6972 ( .A1(n5462), .A2(n5461), .ZN(n6069) );
  INV_X1 U6973 ( .A(n6069), .ZN(n5485) );
  NOR4_X1 U6974 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5466) );
  NOR4_X1 U6975 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5465) );
  NOR4_X1 U6976 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5464) );
  NOR4_X1 U6977 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5463) );
  NAND4_X1 U6978 ( .A1(n5466), .A2(n5465), .A3(n5464), .A4(n5463), .ZN(n5472)
         );
  NOR2_X1 U6979 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n5470) );
  NOR4_X1 U6980 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5469) );
  NOR4_X1 U6981 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5468) );
  NOR4_X1 U6982 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5467) );
  NAND4_X1 U6983 ( .A1(n5470), .A2(n5469), .A3(n5468), .A4(n5467), .ZN(n5471)
         );
  NOR2_X1 U6984 ( .A1(n5472), .A2(n5471), .ZN(n5482) );
  INV_X1 U6985 ( .A(n5482), .ZN(n5473) );
  NAND2_X1 U6986 ( .A1(n5485), .A2(n5473), .ZN(n5475) );
  NAND2_X1 U6987 ( .A1(n7903), .A2(n7740), .ZN(n5483) );
  OAI21_X1 U6988 ( .B1(n6069), .B2(P1_D_REG_0__SCAN_IN), .A(n5483), .ZN(n5474)
         );
  AND2_X1 U6989 ( .A1(n5475), .A2(n5474), .ZN(n6822) );
  NAND2_X1 U6990 ( .A1(n7903), .A2(n7844), .ZN(n6070) );
  OAI21_X1 U6991 ( .B1(n6069), .B2(P1_D_REG_1__SCAN_IN), .A(n6070), .ZN(n6350)
         );
  AND2_X1 U6992 ( .A1(n6822), .A2(n6350), .ZN(n5476) );
  AND2_X2 U6993 ( .A1(n6352), .A2(n5476), .ZN(n9995) );
  INV_X1 U6994 ( .A(n5477), .ZN(n8586) );
  NAND2_X1 U6995 ( .A1(n9995), .A2(n9969), .ZN(n9767) );
  INV_X1 U6996 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n5478) );
  NOR2_X1 U6997 ( .A1(n9995), .A2(n5478), .ZN(n5479) );
  NAND2_X1 U6998 ( .A1(n5481), .A2(n5480), .ZN(P1_U3519) );
  NAND2_X1 U6999 ( .A1(n5482), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5484) );
  INV_X1 U7000 ( .A(n5483), .ZN(n6073) );
  AOI21_X1 U7001 ( .B1(n5485), .B2(n5484), .A(n6073), .ZN(n6351) );
  AND2_X1 U7002 ( .A1(n6351), .A2(n6350), .ZN(n5486) );
  AND2_X2 U7003 ( .A1(n6352), .A2(n5486), .ZN(n10007) );
  NAND2_X1 U7004 ( .A1(n10007), .A2(n9969), .ZN(n9728) );
  NOR2_X1 U7005 ( .A1(n10007), .A2(n5488), .ZN(n5489) );
  NAND2_X1 U7006 ( .A1(n5492), .A2(n5491), .ZN(P1_U3551) );
  INV_X1 U7007 ( .A(n9847), .ZN(n9622) );
  AOI211_X1 U7008 ( .C1(n5390), .C2(n9425), .A(n9622), .B(n4340), .ZN(n9409)
         );
  INV_X1 U7009 ( .A(n5496), .ZN(n5498) );
  OAI211_X1 U7010 ( .C1(n5498), .C2(n8571), .A(n5497), .B(n9693), .ZN(n5504)
         );
  INV_X1 U7011 ( .A(n9964), .ZN(n9985) );
  NAND2_X1 U7012 ( .A1(n9647), .A2(n9985), .ZN(n5502) );
  NAND2_X1 U7013 ( .A1(n5500), .A2(n5499), .ZN(n5501) );
  MUX2_X1 U7014 ( .A(n5506), .B(n9638), .S(n9995), .Z(n5509) );
  INV_X1 U7015 ( .A(n5390), .ZN(n9641) );
  NAND2_X1 U7016 ( .A1(n5390), .A2(n5507), .ZN(n5508) );
  NAND2_X1 U7017 ( .A1(n5509), .A2(n5508), .ZN(P1_U3518) );
  NOR2_X1 U7018 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5513) );
  INV_X1 U7019 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5514) );
  NOR2_X1 U7020 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5521) );
  NOR2_X1 U7021 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5520) );
  NOR2_X1 U7022 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5519) );
  INV_X1 U7023 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5917) );
  INV_X1 U7024 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5523) );
  NAND2_X1 U7025 ( .A1(n4323), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5524) );
  INV_X2 U7026 ( .A(n5642), .ZN(n8047) );
  NAND2_X1 U7027 ( .A1(n7659), .A2(n8047), .ZN(n5529) );
  NAND2_X1 U7028 ( .A1(n5630), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5528) );
  INV_X1 U7029 ( .A(n9154), .ZN(n9023) );
  INV_X1 U7030 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8271) );
  INV_X1 U7031 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7059) );
  INV_X1 U7032 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6781) );
  INV_X1 U7033 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7566) );
  INV_X1 U7034 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5795) );
  INV_X1 U7035 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8004) );
  INV_X1 U7036 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8780) );
  INV_X1 U7037 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U7038 ( .A1(n5829), .A2(n8743), .ZN(n5539) );
  NAND2_X1 U7039 ( .A1(n5839), .A2(n5539), .ZN(n9020) );
  INV_X1 U7040 ( .A(n5543), .ZN(n9211) );
  INV_X1 U7041 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5542) );
  INV_X1 U7042 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5544) );
  OR2_X1 U7043 ( .A1(n9020), .A2(n5911), .ZN(n5553) );
  INV_X1 U7044 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n5550) );
  INV_X1 U7045 ( .A(n4318), .ZN(n5908) );
  NAND2_X1 U7046 ( .A1(n4320), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U7047 ( .A1(n5904), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5548) );
  OAI211_X1 U7048 ( .C1(n5550), .C2(n5908), .A(n5549), .B(n5548), .ZN(n5551)
         );
  INV_X1 U7049 ( .A(n5551), .ZN(n5552) );
  NAND2_X1 U7050 ( .A1(n5553), .A2(n5552), .ZN(n9039) );
  INV_X1 U7051 ( .A(n9039), .ZN(n9009) );
  INV_X1 U7052 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7487) );
  NAND2_X1 U7053 ( .A1(n5798), .A2(n7487), .ZN(n5554) );
  NAND2_X1 U7054 ( .A1(n5806), .A2(n5554), .ZN(n9096) );
  OR2_X1 U7055 ( .A1(n9096), .A2(n5911), .ZN(n5559) );
  INV_X1 U7056 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8904) );
  NAND2_X1 U7057 ( .A1(n4317), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U7058 ( .A1(n4318), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5555) );
  OAI211_X1 U7059 ( .C1(n4312), .C2(n8904), .A(n5556), .B(n5555), .ZN(n5557)
         );
  INV_X1 U7060 ( .A(n5557), .ZN(n5558) );
  NAND2_X1 U7061 ( .A1(n5559), .A2(n5558), .ZN(n9120) );
  INV_X1 U7062 ( .A(n9120), .ZN(n9075) );
  NAND2_X1 U7063 ( .A1(n7118), .A2(n8047), .ZN(n5565) );
  INV_X1 U7064 ( .A(n5630), .ZN(n5647) );
  INV_X1 U7065 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5561) );
  NOR2_X2 U7066 ( .A1(n5778), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n5780) );
  INV_X1 U7067 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5562) );
  INV_X1 U7068 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5946) );
  OAI22_X1 U7069 ( .A1(n5647), .A2(n7121), .B1(n4315), .B2(n4739), .ZN(n5563)
         );
  INV_X1 U7070 ( .A(n5563), .ZN(n5564) );
  INV_X1 U7071 ( .A(n9177), .ZN(n9099) );
  NAND2_X1 U7072 ( .A1(n5904), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U7073 ( .A1(n4317), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5569) );
  INV_X1 U7074 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7556) );
  NAND2_X1 U7075 ( .A1(n5747), .A2(n7556), .ZN(n5566) );
  AND2_X1 U7076 ( .A1(n5759), .A2(n5566), .ZN(n7726) );
  NAND2_X1 U7077 ( .A1(n5872), .A2(n7726), .ZN(n5568) );
  NAND2_X1 U7078 ( .A1(n4318), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5567) );
  NAND4_X1 U7079 ( .A1(n5570), .A2(n5569), .A3(n5568), .A4(n5567), .ZN(n8820)
         );
  INV_X1 U7080 ( .A(n8820), .ZN(n7891) );
  NAND2_X1 U7081 ( .A1(n6315), .A2(n8047), .ZN(n5578) );
  NAND2_X1 U7082 ( .A1(n5614), .A2(n5572), .ZN(n5631) );
  NOR2_X1 U7083 ( .A1(n5631), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5643) );
  NAND2_X1 U7084 ( .A1(n5643), .A2(n5644), .ZN(n5654) );
  NOR2_X1 U7085 ( .A1(n5677), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5690) );
  INV_X1 U7086 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U7087 ( .A1(n5690), .A2(n5573), .ZN(n5702) );
  OAI21_X1 U7088 ( .B1(n5726), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5742) );
  INV_X1 U7089 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5574) );
  NAND2_X1 U7090 ( .A1(n5742), .A2(n5574), .ZN(n5575) );
  NAND2_X1 U7091 ( .A1(n5575), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5753) );
  XNOR2_X1 U7092 ( .A(n5753), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7267) );
  AOI22_X1 U7093 ( .A1(n7267), .A2(n5653), .B1(n5630), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5577) );
  INV_X1 U7094 ( .A(n7727), .ZN(n9808) );
  NAND2_X1 U7095 ( .A1(n5630), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U7096 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5579) );
  XNOR2_X1 U7097 ( .A(n5579), .B(P2_IR_REG_1__SCAN_IN), .ZN(n8830) );
  NAND2_X1 U7098 ( .A1(n5653), .A2(n8830), .ZN(n5580) );
  NAND2_X1 U7099 ( .A1(n5598), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U7100 ( .A1(n4321), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U7101 ( .A1(n5872), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U7102 ( .A1(n4318), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U7103 ( .A1(n5872), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5591) );
  NAND2_X1 U7104 ( .A1(n5598), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7105 ( .A1(n4321), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5587) );
  AND2_X1 U7106 ( .A1(n5588), .A2(n5587), .ZN(n5590) );
  NAND2_X1 U7107 ( .A1(n4318), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5589) );
  INV_X1 U7108 ( .A(SI_0_), .ZN(n5593) );
  INV_X1 U7109 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5592) );
  OAI21_X1 U7110 ( .B1(n5376), .B2(n5593), .A(n5592), .ZN(n5594) );
  AND2_X1 U7111 ( .A1(n5595), .A2(n5594), .ZN(n9222) );
  OAI21_X1 U7112 ( .B1(n6910), .B2(n6463), .A(n6376), .ZN(n5597) );
  NAND2_X1 U7113 ( .A1(n6463), .A2(n6910), .ZN(n5596) );
  AND2_X1 U7114 ( .A1(n5597), .A2(n5596), .ZN(n6947) );
  NAND2_X1 U7115 ( .A1(n5598), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U7116 ( .A1(n4321), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U7117 ( .A1(n5630), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5607) );
  XNOR2_X1 U7118 ( .A(n5605), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6368) );
  NAND2_X1 U7119 ( .A1(n5653), .A2(n6368), .ZN(n5606) );
  NAND2_X1 U7120 ( .A1(n5608), .A2(n6949), .ZN(n5958) );
  NAND2_X1 U7121 ( .A1(n6947), .A2(n8207), .ZN(n6948) );
  NAND2_X1 U7122 ( .A1(n5608), .A2(n10086), .ZN(n5609) );
  NAND2_X1 U7123 ( .A1(n6948), .A2(n5609), .ZN(n10040) );
  NAND2_X1 U7124 ( .A1(n5904), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U7125 ( .A1(n4320), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5612) );
  INV_X1 U7126 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10061) );
  NAND2_X1 U7127 ( .A1(n5872), .A2(n10061), .ZN(n5611) );
  NAND2_X1 U7128 ( .A1(n4318), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5610) );
  NAND2_X1 U7129 ( .A1(n5630), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5619) );
  INV_X1 U7130 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5765) );
  NOR2_X1 U7131 ( .A1(n5614), .A2(n5765), .ZN(n5615) );
  MUX2_X1 U7132 ( .A(n5765), .B(n5615), .S(P2_IR_REG_3__SCAN_IN), .Z(n5617) );
  INV_X1 U7133 ( .A(n5631), .ZN(n5616) );
  NOR2_X1 U7134 ( .A1(n5617), .A2(n5616), .ZN(n8843) );
  NAND2_X1 U7135 ( .A1(n5653), .A2(n8843), .ZN(n5618) );
  NAND2_X1 U7136 ( .A1(n6961), .A2(n10056), .ZN(n8078) );
  INV_X1 U7137 ( .A(n10056), .ZN(n10094) );
  NAND2_X1 U7138 ( .A1(n5620), .A2(n10094), .ZN(n8097) );
  NAND2_X1 U7139 ( .A1(n8078), .A2(n8097), .ZN(n10042) );
  NAND2_X1 U7140 ( .A1(n10040), .A2(n10042), .ZN(n5622) );
  NAND2_X1 U7141 ( .A1(n6961), .A2(n10094), .ZN(n5621) );
  NAND2_X1 U7142 ( .A1(n5622), .A2(n5621), .ZN(n6969) );
  NAND2_X1 U7143 ( .A1(n4316), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U7144 ( .A1(n5904), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5628) );
  INV_X1 U7145 ( .A(n5636), .ZN(n5624) );
  INV_X1 U7146 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7571) );
  NAND2_X1 U7147 ( .A1(n7571), .A2(n10061), .ZN(n5623) );
  NAND2_X1 U7148 ( .A1(n5624), .A2(n5623), .ZN(n6965) );
  INV_X1 U7149 ( .A(n6965), .ZN(n5625) );
  NAND2_X1 U7150 ( .A1(n5872), .A2(n5625), .ZN(n5627) );
  NAND2_X1 U7151 ( .A1(n4318), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5626) );
  NAND4_X1 U7152 ( .A1(n5629), .A2(n5628), .A3(n5627), .A4(n5626), .ZN(n10047)
         );
  NAND2_X1 U7153 ( .A1(n5630), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U7154 ( .A1(n5631), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5632) );
  XNOR2_X1 U7155 ( .A(n5632), .B(P2_IR_REG_4__SCAN_IN), .ZN(n8860) );
  NAND2_X1 U7156 ( .A1(n5653), .A2(n8860), .ZN(n5633) );
  OAI211_X1 U7157 ( .C1(n6084), .C2(n5642), .A(n5634), .B(n5633), .ZN(n6970)
         );
  NAND2_X1 U7158 ( .A1(n6709), .A2(n6970), .ZN(n8079) );
  NAND2_X1 U7159 ( .A1(n10047), .A2(n10098), .ZN(n8098) );
  NAND2_X1 U7160 ( .A1(n8079), .A2(n8098), .ZN(n8208) );
  NAND2_X1 U7161 ( .A1(n6969), .A2(n8208), .ZN(n6968) );
  NAND2_X1 U7162 ( .A1(n6709), .A2(n10098), .ZN(n5635) );
  NAND2_X1 U7163 ( .A1(n6968), .A2(n5635), .ZN(n6730) );
  NAND2_X1 U7164 ( .A1(n5904), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U7165 ( .A1(n4318), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5640) );
  NOR2_X1 U7166 ( .A1(n5636), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5637) );
  NOR2_X1 U7167 ( .A1(n5656), .A2(n5637), .ZN(n6843) );
  NAND2_X1 U7168 ( .A1(n5872), .A2(n6843), .ZN(n5639) );
  NAND2_X1 U7169 ( .A1(n4317), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5638) );
  NAND4_X1 U7170 ( .A1(n5641), .A2(n5640), .A3(n5639), .A4(n5638), .ZN(n8829)
         );
  OR2_X1 U7171 ( .A1(n5642), .A2(n6086), .ZN(n5650) );
  INV_X1 U7172 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6065) );
  OR2_X1 U7173 ( .A1(n5643), .A2(n5765), .ZN(n5645) );
  MUX2_X1 U7174 ( .A(n5645), .B(P2_IR_REG_31__SCAN_IN), .S(n5644), .Z(n5646)
         );
  AND2_X1 U7175 ( .A1(n5646), .A2(n5654), .ZN(n6518) );
  INV_X1 U7176 ( .A(n6518), .ZN(n6064) );
  OAI22_X1 U7177 ( .A1(n5647), .A2(n6065), .B1(n4739), .B2(n6064), .ZN(n5648)
         );
  INV_X1 U7178 ( .A(n5648), .ZN(n5649) );
  NOR2_X1 U7179 ( .A1(n8829), .A2(n6736), .ZN(n5652) );
  INV_X1 U7180 ( .A(n8829), .ZN(n6962) );
  INV_X1 U7181 ( .A(n6736), .ZN(n6845) );
  NAND2_X1 U7182 ( .A1(n8829), .A2(n6845), .ZN(n8100) );
  NAND2_X1 U7183 ( .A1(n6731), .A2(n8829), .ZN(n5651) );
  NAND2_X1 U7184 ( .A1(n5654), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5655) );
  XNOR2_X1 U7185 ( .A(n5655), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6277) );
  NAND2_X1 U7186 ( .A1(n5904), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U7187 ( .A1(n4318), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5662) );
  INV_X1 U7188 ( .A(n5656), .ZN(n5657) );
  INV_X1 U7189 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7572) );
  NAND2_X1 U7190 ( .A1(n5657), .A2(n7572), .ZN(n5658) );
  NAND2_X1 U7191 ( .A1(n5670), .A2(n5658), .ZN(n10025) );
  INV_X1 U7192 ( .A(n10025), .ZN(n5659) );
  NAND2_X1 U7193 ( .A1(n5872), .A2(n5659), .ZN(n5661) );
  NAND2_X1 U7194 ( .A1(n4316), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5660) );
  AND2_X1 U7195 ( .A1(n6902), .A2(n8828), .ZN(n5664) );
  NAND2_X1 U7196 ( .A1(n6088), .A2(n8047), .ZN(n5668) );
  NAND2_X1 U7197 ( .A1(n5665), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5666) );
  XNOR2_X1 U7198 ( .A(n5666), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6541) );
  AOI22_X1 U7199 ( .A1(n5630), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5653), .B2(
        n6541), .ZN(n5667) );
  NAND2_X1 U7200 ( .A1(n5668), .A2(n5667), .ZN(n7013) );
  NAND2_X1 U7201 ( .A1(n4316), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5675) );
  NAND2_X1 U7202 ( .A1(n5904), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5674) );
  INV_X1 U7203 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U7204 ( .A1(n5670), .A2(n5669), .ZN(n5671) );
  AND2_X1 U7205 ( .A1(n5681), .A2(n5671), .ZN(n7012) );
  NAND2_X1 U7206 ( .A1(n5872), .A2(n7012), .ZN(n5673) );
  NAND2_X1 U7207 ( .A1(n4318), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5672) );
  NAND4_X1 U7208 ( .A1(n5675), .A2(n5674), .A3(n5673), .A4(n5672), .ZN(n8827)
         );
  OR2_X1 U7209 ( .A1(n7013), .A2(n6985), .ZN(n8110) );
  NAND2_X1 U7210 ( .A1(n7013), .A2(n6985), .ZN(n8109) );
  NAND2_X1 U7211 ( .A1(n8110), .A2(n8109), .ZN(n8211) );
  OR2_X1 U7212 ( .A1(n7013), .A2(n8827), .ZN(n5676) );
  NAND2_X1 U7213 ( .A1(n6092), .A2(n8047), .ZN(n5680) );
  NAND2_X1 U7214 ( .A1(n5677), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5678) );
  XNOR2_X1 U7215 ( .A(n5678), .B(P2_IR_REG_8__SCAN_IN), .ZN(n8874) );
  AOI22_X1 U7216 ( .A1(n5630), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5653), .B2(
        n8874), .ZN(n5679) );
  NAND2_X1 U7217 ( .A1(n5680), .A2(n5679), .ZN(n6684) );
  NAND2_X1 U7218 ( .A1(n4316), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U7219 ( .A1(n5904), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7220 ( .A1(n5681), .A2(n8878), .ZN(n5682) );
  AND2_X1 U7221 ( .A1(n5695), .A2(n5682), .ZN(n6991) );
  NAND2_X1 U7222 ( .A1(n5872), .A2(n6991), .ZN(n5684) );
  NAND2_X1 U7223 ( .A1(n4318), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5683) );
  NAND4_X1 U7224 ( .A1(n5686), .A2(n5685), .A3(n5684), .A4(n5683), .ZN(n8826)
         );
  INV_X1 U7225 ( .A(n8826), .ZN(n5687) );
  OR2_X1 U7226 ( .A1(n6684), .A2(n5687), .ZN(n8114) );
  NAND2_X1 U7227 ( .A1(n6684), .A2(n5687), .ZN(n8113) );
  NAND2_X1 U7228 ( .A1(n6684), .A2(n8826), .ZN(n5689) );
  NAND2_X1 U7229 ( .A1(n6980), .A2(n5689), .ZN(n7132) );
  INV_X1 U7230 ( .A(n7132), .ZN(n5701) );
  NAND2_X1 U7231 ( .A1(n6102), .A2(n8047), .ZN(n5693) );
  OR2_X1 U7232 ( .A1(n5690), .A2(n5765), .ZN(n5691) );
  XNOR2_X1 U7233 ( .A(n5691), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6545) );
  AOI22_X1 U7234 ( .A1(n5630), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5653), .B2(
        n6545), .ZN(n5692) );
  NAND2_X1 U7235 ( .A1(n5693), .A2(n5692), .ZN(n6807) );
  NAND2_X1 U7236 ( .A1(n4321), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7237 ( .A1(n4318), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5699) );
  INV_X1 U7238 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5694) );
  NAND2_X1 U7239 ( .A1(n5695), .A2(n5694), .ZN(n5696) );
  AND2_X1 U7240 ( .A1(n5708), .A2(n5696), .ZN(n7139) );
  NAND2_X1 U7241 ( .A1(n5872), .A2(n7139), .ZN(n5698) );
  NAND2_X1 U7242 ( .A1(n4317), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5697) );
  NAND4_X1 U7243 ( .A1(n5700), .A2(n5699), .A3(n5698), .A4(n5697), .ZN(n8825)
         );
  INV_X1 U7244 ( .A(n8825), .ZN(n8254) );
  OR2_X1 U7245 ( .A1(n6807), .A2(n8254), .ZN(n8118) );
  NAND2_X1 U7246 ( .A1(n6807), .A2(n8254), .ZN(n8116) );
  AOI21_X1 U7247 ( .B1(n5701), .B2(n8121), .A(n4332), .ZN(n7184) );
  NAND2_X1 U7248 ( .A1(n6111), .A2(n8047), .ZN(n5707) );
  NAND2_X1 U7249 ( .A1(n5702), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5704) );
  INV_X1 U7250 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U7251 ( .A1(n5704), .A2(n5703), .ZN(n5715) );
  OR2_X1 U7252 ( .A1(n5704), .A2(n5703), .ZN(n5705) );
  AOI22_X1 U7253 ( .A1(n5630), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6547), .B2(
        n5653), .ZN(n5706) );
  NAND2_X1 U7254 ( .A1(n4321), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5713) );
  NAND2_X1 U7255 ( .A1(n4318), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U7256 ( .A1(n5708), .A2(n8271), .ZN(n5709) );
  AND2_X1 U7257 ( .A1(n5720), .A2(n5709), .ZN(n7189) );
  NAND2_X1 U7258 ( .A1(n5872), .A2(n7189), .ZN(n5711) );
  NAND2_X1 U7259 ( .A1(n4317), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5710) );
  NAND4_X1 U7260 ( .A1(n5713), .A2(n5712), .A3(n5711), .A4(n5710), .ZN(n8824)
         );
  INV_X1 U7261 ( .A(n8824), .ZN(n5714) );
  NAND2_X1 U7262 ( .A1(n10132), .A2(n5714), .ZN(n8071) );
  NAND2_X1 U7263 ( .A1(n8119), .A2(n8071), .ZN(n8122) );
  NAND2_X1 U7264 ( .A1(n6115), .A2(n8047), .ZN(n5718) );
  NAND2_X1 U7265 ( .A1(n5715), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5716) );
  XNOR2_X1 U7266 ( .A(n5716), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6606) );
  AOI22_X1 U7267 ( .A1(n6606), .A2(n5653), .B1(n5630), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n5717) );
  NAND2_X1 U7268 ( .A1(n4321), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U7269 ( .A1(n4316), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5724) );
  INV_X1 U7270 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5719) );
  NAND2_X1 U7271 ( .A1(n5720), .A2(n5719), .ZN(n5721) );
  AND2_X1 U7272 ( .A1(n5730), .A2(n5721), .ZN(n8796) );
  NAND2_X1 U7273 ( .A1(n5872), .A2(n8796), .ZN(n5723) );
  NAND2_X1 U7274 ( .A1(n4318), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5722) );
  NAND4_X1 U7275 ( .A1(n5725), .A2(n5724), .A3(n5723), .A4(n5722), .ZN(n8823)
         );
  INV_X1 U7276 ( .A(n8823), .ZN(n8252) );
  OR2_X1 U7277 ( .A1(n10141), .A2(n8252), .ZN(n8130) );
  NAND2_X1 U7278 ( .A1(n10141), .A2(n8252), .ZN(n8070) );
  AND2_X1 U7279 ( .A1(n8122), .A2(n8219), .ZN(n7259) );
  NAND2_X1 U7280 ( .A1(n6166), .A2(n8047), .ZN(n5729) );
  NAND2_X1 U7281 ( .A1(n5726), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5727) );
  XNOR2_X1 U7282 ( .A(n5727), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6777) );
  AOI22_X1 U7283 ( .A1(n6777), .A2(n5653), .B1(n5630), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n5728) );
  NAND2_X1 U7284 ( .A1(n5904), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U7285 ( .A1(n4318), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5734) );
  NAND2_X1 U7286 ( .A1(n5730), .A2(n7059), .ZN(n5731) );
  AND2_X1 U7287 ( .A1(n5745), .A2(n5731), .ZN(n7329) );
  NAND2_X1 U7288 ( .A1(n5872), .A2(n7329), .ZN(n5733) );
  NAND2_X1 U7289 ( .A1(n4317), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5732) );
  NAND4_X1 U7290 ( .A1(n5735), .A2(n5734), .A3(n5733), .A4(n5732), .ZN(n8822)
         );
  OR2_X1 U7291 ( .A1(n7330), .A2(n8822), .ZN(n5739) );
  AND2_X1 U7292 ( .A1(n7259), .A2(n5739), .ZN(n5736) );
  NAND2_X1 U7293 ( .A1(n7184), .A2(n5736), .ZN(n5741) );
  NAND2_X1 U7294 ( .A1(n10141), .A2(n8823), .ZN(n7321) );
  INV_X1 U7295 ( .A(n8822), .ZN(n7623) );
  OR2_X1 U7296 ( .A1(n7330), .A2(n7623), .ZN(n8134) );
  NAND2_X1 U7297 ( .A1(n7330), .A2(n7623), .ZN(n8132) );
  AND2_X1 U7298 ( .A1(n7321), .A2(n8220), .ZN(n5738) );
  INV_X1 U7299 ( .A(n8219), .ZN(n5737) );
  NAND2_X1 U7300 ( .A1(n10132), .A2(n8824), .ZN(n7257) );
  OR2_X1 U7301 ( .A1(n5737), .A2(n7257), .ZN(n7260) );
  NAND2_X1 U7302 ( .A1(n4848), .A2(n5739), .ZN(n5740) );
  NAND2_X1 U7303 ( .A1(n5741), .A2(n5740), .ZN(n7621) );
  NAND2_X1 U7304 ( .A1(n6249), .A2(n8047), .ZN(n5744) );
  XNOR2_X1 U7305 ( .A(n5742), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6937) );
  AOI22_X1 U7306 ( .A1(n6937), .A2(n5653), .B1(n5630), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U7307 ( .A1(n5744), .A2(n5743), .ZN(n7048) );
  NAND2_X1 U7308 ( .A1(n4321), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5751) );
  NAND2_X1 U7309 ( .A1(n4318), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U7310 ( .A1(n5745), .A2(n6781), .ZN(n5746) );
  AND2_X1 U7311 ( .A1(n5747), .A2(n5746), .ZN(n7629) );
  NAND2_X1 U7312 ( .A1(n5872), .A2(n7629), .ZN(n5749) );
  NAND2_X1 U7313 ( .A1(n4317), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5748) );
  NAND4_X1 U7314 ( .A1(n5751), .A2(n5750), .A3(n5749), .A4(n5748), .ZN(n8821)
         );
  INV_X1 U7315 ( .A(n8821), .ZN(n7720) );
  OR2_X1 U7316 ( .A1(n7048), .A2(n7720), .ZN(n8138) );
  NAND2_X1 U7317 ( .A1(n7048), .A2(n7720), .ZN(n8139) );
  NAND2_X1 U7318 ( .A1(n8138), .A2(n8139), .ZN(n8221) );
  NAND2_X1 U7319 ( .A1(n7621), .A2(n8221), .ZN(n7620) );
  INV_X1 U7320 ( .A(n7048), .ZN(n9816) );
  NAND2_X1 U7321 ( .A1(n7727), .A2(n7891), .ZN(n8143) );
  NAND2_X1 U7322 ( .A1(n6555), .A2(n8047), .ZN(n5757) );
  INV_X1 U7323 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5752) );
  NAND2_X1 U7324 ( .A1(n5753), .A2(n5752), .ZN(n5754) );
  NAND2_X1 U7325 ( .A1(n5754), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5755) );
  XNOR2_X1 U7326 ( .A(n5755), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7866) );
  AOI22_X1 U7327 ( .A1(n7866), .A2(n5653), .B1(n5630), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5756) );
  INV_X1 U7328 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U7329 ( .A1(n5759), .A2(n5758), .ZN(n5760) );
  AND2_X1 U7330 ( .A1(n5771), .A2(n5760), .ZN(n7894) );
  NAND2_X1 U7331 ( .A1(n7894), .A2(n5872), .ZN(n5764) );
  NAND2_X1 U7332 ( .A1(n4320), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5763) );
  NAND2_X1 U7333 ( .A1(n4321), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U7334 ( .A1(n4318), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5761) );
  NAND4_X1 U7335 ( .A1(n5764), .A2(n5763), .A3(n5762), .A4(n5761), .ZN(n8819)
         );
  INV_X1 U7336 ( .A(n8819), .ZN(n7906) );
  NAND2_X1 U7337 ( .A1(n7895), .A2(n7906), .ZN(n8146) );
  NAND2_X1 U7338 ( .A1(n6746), .A2(n8047), .ZN(n5770) );
  NOR2_X1 U7339 ( .A1(n5560), .A2(n5765), .ZN(n5766) );
  MUX2_X1 U7340 ( .A(n5765), .B(n5766), .S(P2_IR_REG_16__SCAN_IN), .Z(n5767)
         );
  INV_X1 U7341 ( .A(n5767), .ZN(n5768) );
  AND2_X1 U7342 ( .A1(n5768), .A2(n5778), .ZN(n8895) );
  AOI22_X1 U7343 ( .A1(n5630), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5653), .B2(
        n8895), .ZN(n5769) );
  NAND2_X1 U7344 ( .A1(n5771), .A2(n7566), .ZN(n5772) );
  NAND2_X1 U7345 ( .A1(n5784), .A2(n5772), .ZN(n7912) );
  NAND2_X1 U7346 ( .A1(n4321), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5774) );
  NAND2_X1 U7347 ( .A1(n4318), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5773) );
  AND2_X1 U7348 ( .A1(n5774), .A2(n5773), .ZN(n5776) );
  NAND2_X1 U7349 ( .A1(n4317), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5775) );
  OAI211_X1 U7350 ( .C1(n7912), .C2(n5911), .A(n5776), .B(n5775), .ZN(n8818)
         );
  INV_X1 U7351 ( .A(n8818), .ZN(n7955) );
  NAND2_X1 U7352 ( .A1(n9191), .A2(n7955), .ZN(n8150) );
  NOR2_X1 U7353 ( .A1(n7908), .A2(n5777), .ZN(n7958) );
  NAND2_X1 U7354 ( .A1(n6743), .A2(n8047), .ZN(n5783) );
  NAND2_X1 U7355 ( .A1(n5778), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5779) );
  MUX2_X1 U7356 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5779), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5781) );
  INV_X1 U7357 ( .A(n5780), .ZN(n5790) );
  AND2_X1 U7358 ( .A1(n5781), .A2(n5790), .ZN(n7876) );
  AOI22_X1 U7359 ( .A1(n5630), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5653), .B2(
        n7876), .ZN(n5782) );
  INV_X1 U7360 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n5788) );
  INV_X1 U7361 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8262) );
  NAND2_X1 U7362 ( .A1(n5784), .A2(n8262), .ZN(n5785) );
  NAND2_X1 U7363 ( .A1(n5796), .A2(n5785), .ZN(n7960) );
  OR2_X1 U7364 ( .A1(n7960), .A2(n5911), .ZN(n5787) );
  AOI22_X1 U7365 ( .A1(n4318), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n4321), .B2(
        P2_REG1_REG_17__SCAN_IN), .ZN(n5786) );
  OAI211_X1 U7366 ( .C1(n4319), .C2(n5788), .A(n5787), .B(n5786), .ZN(n9119)
         );
  INV_X1 U7367 ( .A(n9119), .ZN(n7907) );
  NAND2_X1 U7368 ( .A1(n9188), .A2(n7907), .ZN(n8065) );
  NAND2_X1 U7369 ( .A1(n8066), .A2(n8065), .ZN(n8228) );
  NAND2_X1 U7370 ( .A1(n7958), .A2(n8228), .ZN(n7957) );
  NAND2_X1 U7371 ( .A1(n7957), .A2(n5789), .ZN(n9108) );
  NAND2_X1 U7372 ( .A1(n6974), .A2(n8047), .ZN(n5794) );
  INV_X1 U7373 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6975) );
  NAND2_X1 U7374 ( .A1(n5790), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5791) );
  XNOR2_X1 U7375 ( .A(n5791), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8907) );
  INV_X1 U7376 ( .A(n8907), .ZN(n7882) );
  OAI22_X1 U7377 ( .A1(n5647), .A2(n6975), .B1(n4739), .B2(n7882), .ZN(n5792)
         );
  INV_X1 U7378 ( .A(n5792), .ZN(n5793) );
  NAND2_X1 U7379 ( .A1(n5796), .A2(n5795), .ZN(n5797) );
  NAND2_X1 U7380 ( .A1(n5798), .A2(n5797), .ZN(n9112) );
  AOI22_X1 U7381 ( .A1(n4320), .A2(P2_REG0_REG_18__SCAN_IN), .B1(n5904), .B2(
        P2_REG1_REG_18__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U7382 ( .A1(n4318), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5799) );
  OAI211_X1 U7383 ( .C1(n9112), .C2(n5911), .A(n5800), .B(n5799), .ZN(n8817)
         );
  NOR2_X1 U7384 ( .A1(n9182), .A2(n8817), .ZN(n5801) );
  INV_X1 U7385 ( .A(n9182), .ZN(n9115) );
  INV_X1 U7386 ( .A(n8817), .ZN(n7956) );
  NOR2_X1 U7387 ( .A1(n9092), .A2(n5802), .ZN(n5803) );
  NAND2_X1 U7388 ( .A1(n7159), .A2(n8047), .ZN(n5805) );
  NAND2_X1 U7389 ( .A1(n5630), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U7390 ( .A1(n5806), .A2(n8004), .ZN(n5807) );
  AND2_X1 U7391 ( .A1(n5816), .A2(n5807), .ZN(n9084) );
  NAND2_X1 U7392 ( .A1(n9084), .A2(n5872), .ZN(n5813) );
  INV_X1 U7393 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U7394 ( .A1(n4320), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5809) );
  NAND2_X1 U7395 ( .A1(n4321), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5808) );
  OAI211_X1 U7396 ( .C1(n5810), .C2(n5908), .A(n5809), .B(n5808), .ZN(n5811)
         );
  INV_X1 U7397 ( .A(n5811), .ZN(n5812) );
  NAND2_X1 U7398 ( .A1(n5813), .A2(n5812), .ZN(n9062) );
  INV_X1 U7399 ( .A(n9062), .ZN(n8752) );
  NAND2_X1 U7400 ( .A1(n9171), .A2(n8752), .ZN(n8162) );
  NAND2_X1 U7401 ( .A1(n9059), .A2(n8162), .ZN(n9080) );
  INV_X1 U7402 ( .A(n9171), .ZN(n9086) );
  NAND2_X1 U7403 ( .A1(n7164), .A2(n8047), .ZN(n5815) );
  NAND2_X1 U7404 ( .A1(n5630), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5814) );
  INV_X1 U7405 ( .A(n9164), .ZN(n9057) );
  INV_X1 U7406 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8750) );
  NAND2_X1 U7407 ( .A1(n5816), .A2(n8750), .ZN(n5817) );
  NAND2_X1 U7408 ( .A1(n5827), .A2(n5817), .ZN(n9054) );
  OR2_X1 U7409 ( .A1(n9054), .A2(n5911), .ZN(n5823) );
  INV_X1 U7410 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n5820) );
  NAND2_X1 U7411 ( .A1(n5904), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5819) );
  NAND2_X1 U7412 ( .A1(n4317), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5818) );
  OAI211_X1 U7413 ( .C1(n5820), .C2(n5908), .A(n5819), .B(n5818), .ZN(n5821)
         );
  INV_X1 U7414 ( .A(n5821), .ZN(n5822) );
  NAND2_X1 U7415 ( .A1(n5823), .A2(n5822), .ZN(n9038) );
  INV_X1 U7416 ( .A(n9038), .ZN(n9077) );
  NAND2_X1 U7417 ( .A1(n9057), .A2(n9077), .ZN(n5824) );
  NAND2_X1 U7418 ( .A1(n7398), .A2(n8047), .ZN(n5826) );
  NAND2_X1 U7419 ( .A1(n5630), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5825) );
  NAND2_X1 U7420 ( .A1(n5827), .A2(n8780), .ZN(n5828) );
  AND2_X1 U7421 ( .A1(n5829), .A2(n5828), .ZN(n9045) );
  NAND2_X1 U7422 ( .A1(n9045), .A2(n5872), .ZN(n5835) );
  INV_X1 U7423 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n5832) );
  NAND2_X1 U7424 ( .A1(n4316), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5831) );
  NAND2_X1 U7425 ( .A1(n4321), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5830) );
  OAI211_X1 U7426 ( .C1(n5832), .C2(n5908), .A(n5831), .B(n5830), .ZN(n5833)
         );
  INV_X1 U7427 ( .A(n5833), .ZN(n5834) );
  NAND2_X1 U7428 ( .A1(n5835), .A2(n5834), .ZN(n9063) );
  INV_X1 U7429 ( .A(n9063), .ZN(n8751) );
  NAND2_X1 U7430 ( .A1(n9161), .A2(n8751), .ZN(n8169) );
  NAND2_X1 U7431 ( .A1(n9024), .A2(n8169), .ZN(n5966) );
  AOI21_X2 U7432 ( .B1(n9033), .B2(n5966), .A(n5836), .ZN(n9018) );
  OR2_X1 U7433 ( .A1(n9154), .A2(n9009), .ZN(n8062) );
  NAND2_X1 U7434 ( .A1(n7738), .A2(n8047), .ZN(n5838) );
  NAND2_X1 U7435 ( .A1(n5630), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5837) );
  INV_X1 U7436 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8771) );
  NAND2_X1 U7437 ( .A1(n5839), .A2(n8771), .ZN(n5840) );
  NAND2_X1 U7438 ( .A1(n5849), .A2(n5840), .ZN(n9002) );
  OR2_X1 U7439 ( .A1(n9002), .A2(n5911), .ZN(n5846) );
  INV_X1 U7440 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n5843) );
  NAND2_X1 U7441 ( .A1(n4321), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5842) );
  NAND2_X1 U7442 ( .A1(n4316), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5841) );
  OAI211_X1 U7443 ( .C1(n5908), .C2(n5843), .A(n5842), .B(n5841), .ZN(n5844)
         );
  INV_X1 U7444 ( .A(n5844), .ZN(n5845) );
  NAND2_X1 U7445 ( .A1(n9149), .A2(n8988), .ZN(n8173) );
  INV_X1 U7446 ( .A(n8988), .ZN(n9028) );
  NAND2_X1 U7447 ( .A1(n7841), .A2(n8047), .ZN(n5848) );
  NAND2_X1 U7448 ( .A1(n5630), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5847) );
  INV_X1 U7449 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8759) );
  NAND2_X1 U7450 ( .A1(n5849), .A2(n8759), .ZN(n5850) );
  AND2_X1 U7451 ( .A1(n5861), .A2(n5850), .ZN(n8991) );
  NAND2_X1 U7452 ( .A1(n8991), .A2(n5872), .ZN(n5856) );
  INV_X1 U7453 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n5853) );
  NAND2_X1 U7454 ( .A1(n4321), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5852) );
  NAND2_X1 U7455 ( .A1(n4317), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5851) );
  OAI211_X1 U7456 ( .C1(n5853), .C2(n5908), .A(n5852), .B(n5851), .ZN(n5854)
         );
  INV_X1 U7457 ( .A(n5854), .ZN(n5855) );
  NAND2_X1 U7458 ( .A1(n5856), .A2(n5855), .ZN(n8965) );
  INV_X1 U7459 ( .A(n8965), .ZN(n9010) );
  NAND2_X1 U7460 ( .A1(n9146), .A2(n9010), .ZN(n8176) );
  NAND2_X1 U7461 ( .A1(n8981), .A2(n5857), .ZN(n8970) );
  NAND2_X1 U7462 ( .A1(n7901), .A2(n8047), .ZN(n5859) );
  NAND2_X1 U7463 ( .A1(n5630), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5858) );
  INV_X1 U7464 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8804) );
  NAND2_X1 U7465 ( .A1(n5861), .A2(n8804), .ZN(n5862) );
  NAND2_X1 U7466 ( .A1(n5884), .A2(n5862), .ZN(n8976) );
  OR2_X1 U7467 ( .A1(n8976), .A2(n5911), .ZN(n5867) );
  INV_X1 U7468 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8974) );
  NAND2_X1 U7469 ( .A1(n5904), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U7470 ( .A1(n4320), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5863) );
  OAI211_X1 U7471 ( .C1(n5908), .C2(n8974), .A(n5864), .B(n5863), .ZN(n5865)
         );
  INV_X1 U7472 ( .A(n5865), .ZN(n5866) );
  NAND2_X1 U7473 ( .A1(n5867), .A2(n5866), .ZN(n8951) );
  INV_X1 U7474 ( .A(n8951), .ZN(n8989) );
  OR2_X1 U7475 ( .A1(n9140), .A2(n8989), .ZN(n8182) );
  NAND2_X1 U7476 ( .A1(n9140), .A2(n8989), .ZN(n8177) );
  NAND2_X1 U7477 ( .A1(n8182), .A2(n8177), .ZN(n8969) );
  NAND2_X1 U7478 ( .A1(n8970), .A2(n8969), .ZN(n8968) );
  NAND2_X1 U7479 ( .A1(n8968), .A2(n5869), .ZN(n8946) );
  NAND2_X1 U7480 ( .A1(n5630), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5870) );
  XNOR2_X1 U7481 ( .A(n5884), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8956) );
  NAND2_X1 U7482 ( .A1(n8956), .A2(n5872), .ZN(n5878) );
  INV_X1 U7483 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U7484 ( .A1(n4320), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U7485 ( .A1(n5904), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5873) );
  OAI211_X1 U7486 ( .C1(n5875), .C2(n5908), .A(n5874), .B(n5873), .ZN(n5876)
         );
  INV_X1 U7487 ( .A(n5876), .ZN(n5877) );
  NAND2_X1 U7488 ( .A1(n5878), .A2(n5877), .ZN(n8966) );
  INV_X1 U7489 ( .A(n8966), .ZN(n8057) );
  NAND2_X1 U7490 ( .A1(n8946), .A2(n8945), .ZN(n8944) );
  NAND2_X1 U7491 ( .A1(n5880), .A2(n8047), .ZN(n5882) );
  NAND2_X1 U7492 ( .A1(n5630), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5881) );
  INV_X1 U7493 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8736) );
  INV_X1 U7494 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5883) );
  OAI21_X1 U7495 ( .B1(n5884), .B2(n8736), .A(n5883), .ZN(n5885) );
  NAND2_X1 U7496 ( .A1(n5885), .A2(n5981), .ZN(n8635) );
  INV_X1 U7497 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U7498 ( .A1(n4317), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5887) );
  NAND2_X1 U7499 ( .A1(n5904), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5886) );
  OAI211_X1 U7500 ( .C1(n5888), .C2(n5908), .A(n5887), .B(n5886), .ZN(n5889)
         );
  INV_X1 U7501 ( .A(n5889), .ZN(n5890) );
  NAND2_X1 U7502 ( .A1(n5891), .A2(n5890), .ZN(n8952) );
  NAND2_X1 U7503 ( .A1(n8640), .A2(n5892), .ZN(n8188) );
  NAND2_X1 U7504 ( .A1(n5893), .A2(n5892), .ZN(n5894) );
  INV_X1 U7505 ( .A(n5897), .ZN(n5899) );
  NAND2_X1 U7506 ( .A1(n5899), .A2(n5898), .ZN(n5900) );
  MUX2_X1 U7507 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n5376), .Z(n6007) );
  INV_X1 U7508 ( .A(SI_29_), .ZN(n7589) );
  XNOR2_X1 U7509 ( .A(n6007), .B(n7589), .ZN(n6005) );
  NAND2_X1 U7510 ( .A1(n9217), .A2(n8047), .ZN(n5903) );
  NAND2_X1 U7511 ( .A1(n5630), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5902) );
  INV_X1 U7512 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U7513 ( .A1(n5904), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U7514 ( .A1(n4316), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5905) );
  OAI211_X1 U7515 ( .C1(n5908), .C2(n5907), .A(n5906), .B(n5905), .ZN(n5909)
         );
  INV_X1 U7516 ( .A(n5909), .ZN(n5910) );
  OAI21_X1 U7517 ( .B1(n5981), .B2(n5911), .A(n5910), .ZN(n8815) );
  INV_X1 U7518 ( .A(n8815), .ZN(n5912) );
  NAND2_X1 U7519 ( .A1(n5913), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5914) );
  MUX2_X1 U7520 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5914), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5915) );
  NAND2_X1 U7521 ( .A1(n5915), .A2(n5526), .ZN(n7920) );
  NAND2_X1 U7522 ( .A1(n5916), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5918) );
  MUX2_X1 U7523 ( .A(n5918), .B(P2_IR_REG_31__SCAN_IN), .S(n5917), .Z(n5919)
         );
  NAND2_X1 U7524 ( .A1(n5919), .A2(n5913), .ZN(n7842) );
  INV_X1 U7525 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5921) );
  INV_X1 U7526 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5942) );
  NAND2_X1 U7527 ( .A1(n5943), .A2(n5942), .ZN(n5922) );
  NAND2_X1 U7528 ( .A1(n5922), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5941) );
  INV_X1 U7529 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U7530 ( .A1(n5941), .A2(n5923), .ZN(n5924) );
  NAND2_X1 U7531 ( .A1(n5924), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5926) );
  INV_X1 U7532 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5925) );
  XNOR2_X1 U7533 ( .A(n5926), .B(n5925), .ZN(n7743) );
  INV_X1 U7534 ( .A(P2_B_REG_SCAN_IN), .ZN(n5927) );
  XOR2_X1 U7535 ( .A(n7743), .B(n5927), .Z(n5928) );
  AND2_X1 U7536 ( .A1(n7842), .A2(n5928), .ZN(n5929) );
  INV_X1 U7537 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10076) );
  AND2_X1 U7538 ( .A1(n7842), .A2(n7920), .ZN(n10078) );
  AOI21_X1 U7539 ( .B1(n10071), .B2(n10076), .A(n10078), .ZN(n6047) );
  NOR4_X1 U7540 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5933) );
  NOR4_X1 U7541 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5932) );
  NOR4_X1 U7542 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5931) );
  NOR4_X1 U7543 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5930) );
  NAND4_X1 U7544 ( .A1(n5933), .A2(n5932), .A3(n5931), .A4(n5930), .ZN(n5939)
         );
  NOR2_X1 U7545 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n5937) );
  NOR4_X1 U7546 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5936) );
  NOR4_X1 U7547 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5935) );
  NOR4_X1 U7548 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5934) );
  NAND4_X1 U7549 ( .A1(n5937), .A2(n5936), .A3(n5935), .A4(n5934), .ZN(n5938)
         );
  OAI21_X1 U7550 ( .B1(n5939), .B2(n5938), .A(n10071), .ZN(n6045) );
  AND2_X1 U7551 ( .A1(n6047), .A2(n6045), .ZN(n6481) );
  AND2_X1 U7552 ( .A1(n7743), .A2(n7920), .ZN(n10074) );
  INV_X1 U7553 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10073) );
  AND2_X1 U7554 ( .A1(n10071), .A2(n10073), .ZN(n5940) );
  NOR2_X1 U7555 ( .A1(n10074), .A2(n5940), .ZN(n6480) );
  OR3_X1 U7556 ( .A1(n7743), .A2(n7920), .A3(n7842), .ZN(n6580) );
  XNOR2_X1 U7557 ( .A(n5941), .B(P2_IR_REG_23__SCAN_IN), .ZN(n6096) );
  NOR2_X1 U7558 ( .A1(n6096), .A2(P2_U3152), .ZN(n10077) );
  NAND2_X1 U7559 ( .A1(n6580), .A2(n10077), .ZN(n10072) );
  INV_X1 U7560 ( .A(n5953), .ZN(n8248) );
  NAND2_X1 U7561 ( .A1(n5944), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5945) );
  INV_X1 U7562 ( .A(n8242), .ZN(n8083) );
  NAND2_X1 U7563 ( .A1(n8248), .A2(n8083), .ZN(n6461) );
  NAND2_X1 U7564 ( .A1(n5947), .A2(n5946), .ZN(n5948) );
  INV_X1 U7565 ( .A(n8238), .ZN(n7161) );
  AND2_X1 U7566 ( .A1(n7161), .A2(n4315), .ZN(n6474) );
  OR2_X1 U7567 ( .A1(n6461), .A2(n6474), .ZN(n6578) );
  INV_X1 U7568 ( .A(n6578), .ZN(n5950) );
  OR2_X1 U7569 ( .A1(n10072), .A2(n5950), .ZN(n8247) );
  NOR2_X1 U7570 ( .A1(n6480), .A2(n8247), .ZN(n5951) );
  NAND2_X1 U7571 ( .A1(n6481), .A2(n5951), .ZN(n5980) );
  INV_X1 U7572 ( .A(n7025), .ZN(n5952) );
  OR2_X1 U7573 ( .A1(n10055), .A2(n4315), .ZN(n6482) );
  NAND2_X2 U7574 ( .A1(n5980), .A2(n8975), .ZN(n9049) );
  NAND2_X1 U7575 ( .A1(n7161), .A2(n8083), .ZN(n6464) );
  XNOR2_X1 U7576 ( .A(n5953), .B(n6464), .ZN(n5954) );
  OR2_X1 U7577 ( .A1(n5954), .A2(n5979), .ZN(n10039) );
  OR2_X1 U7578 ( .A1(n6464), .A2(n4315), .ZN(n6981) );
  NAND2_X1 U7579 ( .A1(n10039), .A2(n6981), .ZN(n5955) );
  NAND2_X1 U7580 ( .A1(n9049), .A2(n5955), .ZN(n9126) );
  NAND2_X1 U7581 ( .A1(n8092), .A2(n6691), .ZN(n6380) );
  INV_X1 U7582 ( .A(n6951), .ZN(n5957) );
  NAND2_X1 U7583 ( .A1(n6950), .A2(n5958), .ZN(n5959) );
  NAND2_X1 U7584 ( .A1(n6732), .A2(n8080), .ZN(n5960) );
  NAND2_X1 U7585 ( .A1(n5960), .A2(n8100), .ZN(n6897) );
  INV_X1 U7586 ( .A(n8828), .ZN(n6592) );
  XNOR2_X1 U7587 ( .A(n6592), .B(n6902), .ZN(n8212) );
  NAND2_X1 U7588 ( .A1(n6592), .A2(n6902), .ZN(n8108) );
  INV_X1 U7589 ( .A(n8116), .ZN(n5962) );
  INV_X1 U7590 ( .A(n8122), .ZN(n8217) );
  INV_X1 U7591 ( .A(n8119), .ZN(n7248) );
  NAND2_X1 U7592 ( .A1(n8132), .A2(n8070), .ZN(n8127) );
  INV_X1 U7593 ( .A(n8224), .ZN(n7719) );
  INV_X1 U7594 ( .A(n8142), .ZN(n5963) );
  INV_X1 U7595 ( .A(n8147), .ZN(n5964) );
  INV_X1 U7596 ( .A(n8228), .ZN(n8154) );
  OR2_X1 U7597 ( .A1(n9182), .A2(n7956), .ZN(n8159) );
  NAND2_X1 U7598 ( .A1(n9182), .A2(n7956), .ZN(n8156) );
  NAND2_X1 U7599 ( .A1(n9117), .A2(n9118), .ZN(n9116) );
  NAND2_X1 U7600 ( .A1(n9116), .A2(n8156), .ZN(n9100) );
  NOR2_X1 U7601 ( .A1(n9177), .A2(n9075), .ZN(n8161) );
  NOR2_X1 U7602 ( .A1(n8161), .A2(n8158), .ZN(n9101) );
  INV_X1 U7603 ( .A(n9080), .ZN(n9069) );
  INV_X1 U7604 ( .A(n8158), .ZN(n9070) );
  OR2_X1 U7605 ( .A1(n9164), .A2(n9077), .ZN(n8166) );
  NAND2_X1 U7606 ( .A1(n9164), .A2(n9077), .ZN(n9037) );
  NAND2_X1 U7607 ( .A1(n9058), .A2(n4831), .ZN(n9035) );
  NAND2_X2 U7608 ( .A1(n9034), .A2(n4836), .ZN(n9025) );
  INV_X1 U7609 ( .A(n8969), .ZN(n8964) );
  AND2_X2 U7610 ( .A1(n8962), .A2(n8177), .ZN(n8950) );
  OR2_X1 U7611 ( .A1(n9135), .A2(n8057), .ZN(n8058) );
  NAND2_X1 U7612 ( .A1(n8948), .A2(n8058), .ZN(n6032) );
  INV_X1 U7613 ( .A(n8059), .ZN(n5969) );
  OAI21_X1 U7614 ( .B1(n8205), .B2(n5970), .A(n8035), .ZN(n5977) );
  NAND2_X1 U7615 ( .A1(n8083), .A2(n8238), .ZN(n8054) );
  NAND2_X1 U7616 ( .A1(n8239), .A2(n8054), .ZN(n10049) );
  INV_X1 U7617 ( .A(n6461), .ZN(n6253) );
  INV_X1 U7618 ( .A(n6293), .ZN(n8010) );
  AND2_X1 U7619 ( .A1(n6253), .A2(n8010), .ZN(n10045) );
  AND2_X1 U7620 ( .A1(n6253), .A2(n6293), .ZN(n10046) );
  INV_X1 U7621 ( .A(n8246), .ZN(n7921) );
  NAND2_X1 U7622 ( .A1(n7921), .A2(P2_B_REG_SCAN_IN), .ZN(n5971) );
  AND2_X1 U7623 ( .A1(n10046), .A2(n5971), .ZN(n8923) );
  NAND2_X1 U7624 ( .A1(n5598), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U7625 ( .A1(n4321), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U7626 ( .A1(n4318), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5972) );
  NAND3_X1 U7627 ( .A1(n5974), .A2(n5973), .A3(n5972), .ZN(n8814) );
  NOR2_X1 U7628 ( .A1(n10058), .A2(n6970), .ZN(n6734) );
  NAND2_X1 U7629 ( .A1(n6734), .A2(n6845), .ZN(n6735) );
  INV_X1 U7630 ( .A(n6684), .ZN(n10118) );
  INV_X1 U7631 ( .A(n6807), .ZN(n10125) );
  INV_X1 U7632 ( .A(n7330), .ZN(n10151) );
  INV_X1 U7633 ( .A(n9188), .ZN(n7963) );
  NAND2_X1 U7634 ( .A1(n4802), .A2(n9019), .ZN(n8999) );
  AOI21_X1 U7635 ( .B1(n9127), .B2(n6035), .A(n8930), .ZN(n9128) );
  OR2_X1 U7636 ( .A1(n5980), .A2(n5979), .ZN(n10065) );
  NOR2_X1 U7637 ( .A1(n10065), .A2(n10055), .ZN(n9088) );
  NOR2_X1 U7638 ( .A1(n10081), .A2(n7161), .ZN(n6477) );
  NAND2_X1 U7639 ( .A1(n9049), .A2(n6477), .ZN(n10054) );
  INV_X1 U7640 ( .A(n5981), .ZN(n5982) );
  INV_X1 U7641 ( .A(n8975), .ZN(n10062) );
  AOI22_X1 U7642 ( .A1(n5982), .A2(n10062), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n10070), .ZN(n5983) );
  OAI21_X1 U7643 ( .B1(n4486), .B2(n10054), .A(n5983), .ZN(n5984) );
  OAI211_X1 U7644 ( .C1(n9131), .C2(n9126), .A(n4843), .B(n5985), .ZN(P2_U3267) );
  NAND2_X1 U7645 ( .A1(n5986), .A2(n4844), .ZN(n5989) );
  NAND2_X1 U7646 ( .A1(n9217), .A2(n4998), .ZN(n5988) );
  INV_X1 U7647 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9778) );
  OR2_X1 U7648 ( .A1(n8397), .A2(n9778), .ZN(n5987) );
  XNOR2_X1 U7649 ( .A(n5989), .B(n8453), .ZN(n8020) );
  INV_X1 U7650 ( .A(P1_B_REG_SCAN_IN), .ZN(n5991) );
  NOR2_X1 U7651 ( .A1(n8588), .A2(n5991), .ZN(n5992) );
  NOR2_X1 U7652 ( .A1(n9962), .A2(n5992), .ZN(n6020) );
  INV_X1 U7653 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U7654 ( .A1(n5042), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U7655 ( .A1(n5993), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5994) );
  OAI211_X1 U7656 ( .C1(n5997), .C2(n5996), .A(n5995), .B(n5994), .ZN(n9322)
         );
  INV_X1 U7657 ( .A(n6000), .ZN(n6001) );
  OAI211_X1 U7658 ( .C1(n4438), .C2(n6001), .A(n9847), .B(n6013), .ZN(n8024)
         );
  NAND2_X1 U7659 ( .A1(n5500), .A2(n9985), .ZN(n6002) );
  NAND3_X1 U7660 ( .A1(n8029), .A2(n8024), .A3(n6002), .ZN(n6003) );
  OAI21_X1 U7661 ( .B1(n6055), .B2(n10005), .A(n4838), .ZN(P1_U3552) );
  INV_X1 U7662 ( .A(n6007), .ZN(n6008) );
  NAND2_X1 U7663 ( .A1(n6008), .A2(n7589), .ZN(n6009) );
  MUX2_X1 U7664 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n5376), .Z(n8038) );
  INV_X1 U7665 ( .A(SI_30_), .ZN(n8039) );
  XNOR2_X1 U7666 ( .A(n8038), .B(n8039), .ZN(n8036) );
  NAND2_X1 U7667 ( .A1(n8732), .A2(n4998), .ZN(n6012) );
  INV_X1 U7668 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8733) );
  OR2_X1 U7669 ( .A1(n8397), .A2(n8733), .ZN(n6011) );
  INV_X1 U7670 ( .A(n9380), .ZN(n6015) );
  NAND2_X1 U7671 ( .A1(n8452), .A2(n6013), .ZN(n6014) );
  NAND2_X1 U7672 ( .A1(n6015), .A2(n4842), .ZN(n9389) );
  INV_X1 U7673 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7674 ( .A1(n4933), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6018) );
  INV_X1 U7675 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6016) );
  OR2_X1 U7676 ( .A1(n4932), .A2(n6016), .ZN(n6017) );
  OAI211_X1 U7677 ( .C1(n4936), .C2(n6019), .A(n6018), .B(n6017), .ZN(n8411)
         );
  AND2_X1 U7678 ( .A1(n6020), .A2(n8411), .ZN(n9634) );
  INV_X1 U7679 ( .A(n9634), .ZN(n9382) );
  MUX2_X1 U7680 ( .A(n6024), .B(n5996), .S(n10005), .Z(n6022) );
  INV_X1 U7681 ( .A(n8452), .ZN(n9385) );
  NAND2_X1 U7682 ( .A1(n6022), .A2(n6021), .ZN(P1_U3553) );
  INV_X1 U7683 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n6023) );
  MUX2_X1 U7684 ( .A(n6024), .B(n6023), .S(n9994), .Z(n6026) );
  NAND2_X1 U7685 ( .A1(n6026), .A2(n6025), .ZN(P1_U3521) );
  OAI21_X1 U7686 ( .B1(n6029), .B2(n6028), .A(n6027), .ZN(n6030) );
  INV_X1 U7687 ( .A(n6030), .ZN(n8943) );
  NOR2_X1 U7688 ( .A1(n8238), .A2(n4315), .ZN(n6031) );
  NAND2_X1 U7689 ( .A1(n6031), .A2(n5953), .ZN(n9814) );
  XNOR2_X1 U7690 ( .A(n6032), .B(n6028), .ZN(n6033) );
  INV_X1 U7691 ( .A(n10049), .ZN(n9071) );
  NAND2_X1 U7692 ( .A1(n6033), .A2(n10049), .ZN(n6034) );
  AOI22_X1 U7693 ( .A1(n8966), .A2(n10045), .B1(n8815), .B2(n10046), .ZN(n8638) );
  NAND2_X1 U7694 ( .A1(n6034), .A2(n8638), .ZN(n8941) );
  INV_X1 U7695 ( .A(n8955), .ZN(n6037) );
  INV_X1 U7696 ( .A(n6035), .ZN(n6036) );
  AOI211_X1 U7697 ( .C1(n8640), .C2(n6037), .A(n10055), .B(n6036), .ZN(n8936)
         );
  OR2_X1 U7698 ( .A1(n10081), .A2(n6474), .ZN(n10150) );
  INV_X1 U7699 ( .A(n10150), .ZN(n10142) );
  INV_X1 U7700 ( .A(n6482), .ZN(n6043) );
  NOR2_X1 U7701 ( .A1(n8247), .A2(n6043), .ZN(n6044) );
  NAND2_X1 U7702 ( .A1(n6045), .A2(n6044), .ZN(n6046) );
  OR2_X1 U7703 ( .A1(n6047), .A2(n6046), .ZN(n6393) );
  INV_X2 U7704 ( .A(n10156), .ZN(n10158) );
  NAND2_X1 U7705 ( .A1(n9132), .A2(n10158), .ZN(n6050) );
  INV_X1 U7706 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6048) );
  OR2_X1 U7707 ( .A1(n10158), .A2(n6048), .ZN(n6049) );
  OAI21_X1 U7708 ( .B1(n6055), .B2(n9994), .A(n6054), .ZN(P1_U3520) );
  INV_X1 U7709 ( .A(n7660), .ZN(n6056) );
  OR2_X1 U7710 ( .A1(n8460), .A2(n6056), .ZN(n6057) );
  INV_X1 U7711 ( .A(n6624), .ZN(n6323) );
  NAND2_X1 U7712 ( .A1(n6323), .A2(n7660), .ZN(n6119) );
  NAND2_X1 U7713 ( .A1(n6057), .A2(n6119), .ZN(n6145) );
  OR2_X1 U7714 ( .A1(n6145), .A2(n6058), .ZN(n6125) );
  NAND2_X1 U7715 ( .A1(n6125), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NOR2_X1 U7716 ( .A1(n6580), .A2(P2_U3152), .ZN(n6251) );
  INV_X1 U7717 ( .A(n6096), .ZN(n6579) );
  AND2_X2 U7718 ( .A1(n6251), .A2(n6579), .ZN(P2_U3966) );
  INV_X1 U7719 ( .A(n6074), .ZN(n6059) );
  OR2_X1 U7720 ( .A1(n6624), .A2(n6059), .ZN(n9330) );
  INV_X2 U7721 ( .A(n9330), .ZN(P1_U4006) );
  XNOR2_X1 U7722 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AND2_X1 U7723 ( .A1(n6066), .A2(P2_U3152), .ZN(n9218) );
  AOI22_X1 U7724 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n9218), .B1(n6368), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6060) );
  OAI21_X1 U7725 ( .B1(n6078), .B2(n9221), .A(n6060), .ZN(P2_U3356) );
  INV_X1 U7726 ( .A(n9218), .ZN(n8019) );
  INV_X1 U7727 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6061) );
  INV_X1 U7728 ( .A(n8843), .ZN(n6282) );
  OAI222_X1 U7729 ( .A1(n8019), .A2(n6061), .B1(n9221), .B2(n6076), .C1(
        P2_U3152), .C2(n6282), .ZN(P2_U3355) );
  INV_X1 U7730 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6062) );
  INV_X1 U7731 ( .A(n8830), .ZN(n6279) );
  OAI222_X1 U7732 ( .A1(n8019), .A2(n6062), .B1(n9221), .B2(n6067), .C1(
        P2_U3152), .C2(n6279), .ZN(P2_U3357) );
  INV_X1 U7733 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6063) );
  INV_X1 U7734 ( .A(n8860), .ZN(n6284) );
  OAI222_X1 U7735 ( .A1(n8019), .A2(n6063), .B1(n9221), .B2(n6084), .C1(
        P2_U3152), .C2(n6284), .ZN(P2_U3354) );
  OAI222_X1 U7736 ( .A1(n8019), .A2(n6065), .B1(n9221), .B2(n6086), .C1(
        P2_U3152), .C2(n6064), .ZN(P2_U3353) );
  OR2_X1 U7737 ( .A1(n6066), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9777) );
  NAND2_X1 U7738 ( .A1(n5376), .A2(P1_U3084), .ZN(n7846) );
  OAI222_X1 U7739 ( .A1(n9777), .A2(n6068), .B1(n7846), .B2(n6067), .C1(
        P1_U3084), .C2(n6150), .ZN(P1_U3352) );
  NAND2_X1 U7740 ( .A1(n6355), .A2(n6069), .ZN(n9940) );
  INV_X1 U7741 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6072) );
  INV_X1 U7742 ( .A(n6070), .ZN(n6071) );
  AOI22_X1 U7743 ( .A1(n9940), .A2(n6072), .B1(n6074), .B2(n6071), .ZN(
        P1_U3441) );
  INV_X1 U7744 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6075) );
  AOI22_X1 U7745 ( .A1(n9940), .A2(n6075), .B1(n6074), .B2(n6073), .ZN(
        P1_U3440) );
  INV_X1 U7746 ( .A(n9777), .ZN(n6744) );
  INV_X1 U7747 ( .A(n6744), .ZN(n9771) );
  OAI222_X1 U7748 ( .A1(n9771), .A2(n6077), .B1(n7846), .B2(n6076), .C1(
        P1_U3084), .C2(n6173), .ZN(P1_U3350) );
  OAI222_X1 U7749 ( .A1(n9771), .A2(n6079), .B1(n7846), .B2(n6078), .C1(
        P1_U3084), .C2(n6403), .ZN(P1_U3351) );
  INV_X1 U7750 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6081) );
  INV_X1 U7751 ( .A(n6080), .ZN(n6082) );
  OAI222_X1 U7752 ( .A1(n8019), .A2(n6081), .B1(n9221), .B2(n6082), .C1(
        P2_U3152), .C2(n4740), .ZN(P2_U3352) );
  INV_X1 U7753 ( .A(n7846), .ZN(n8013) );
  INV_X1 U7754 ( .A(n8013), .ZN(n9781) );
  OAI222_X1 U7755 ( .A1(n9771), .A2(n6083), .B1(n9781), .B2(n6082), .C1(
        P1_U3084), .C2(n6218), .ZN(P1_U3347) );
  OAI222_X1 U7756 ( .A1(n9771), .A2(n6085), .B1(n9781), .B2(n6084), .C1(
        P1_U3084), .C2(n6347), .ZN(P1_U3349) );
  OAI222_X1 U7757 ( .A1(n9771), .A2(n6087), .B1(n9781), .B2(n6086), .C1(
        P1_U3084), .C2(n6202), .ZN(P1_U3348) );
  INV_X1 U7758 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6089) );
  INV_X1 U7759 ( .A(n6088), .ZN(n6090) );
  INV_X1 U7760 ( .A(n6235), .ZN(n6224) );
  OAI222_X1 U7761 ( .A1(n9771), .A2(n6089), .B1(n7846), .B2(n6090), .C1(
        P1_U3084), .C2(n6224), .ZN(P1_U3346) );
  INV_X1 U7762 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6091) );
  INV_X1 U7763 ( .A(n6541), .ZN(n6273) );
  OAI222_X1 U7764 ( .A1(n8019), .A2(n6091), .B1(n9221), .B2(n6090), .C1(
        P2_U3152), .C2(n6273), .ZN(P2_U3351) );
  INV_X1 U7765 ( .A(n6092), .ZN(n6094) );
  AOI22_X1 U7766 ( .A1(n8874), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n9218), .ZN(n6093) );
  OAI21_X1 U7767 ( .B1(n6094), .B2(n9221), .A(n6093), .ZN(P2_U3350) );
  INV_X1 U7768 ( .A(n6238), .ZN(n9883) );
  OAI222_X1 U7769 ( .A1(n9771), .A2(n6095), .B1(n7846), .B2(n6094), .C1(
        P1_U3084), .C2(n9883), .ZN(P1_U3345) );
  NAND2_X1 U7770 ( .A1(n6096), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8251) );
  NAND2_X1 U7771 ( .A1(n10072), .A2(n8251), .ZN(n6097) );
  NAND2_X1 U7772 ( .A1(n6097), .A2(n5653), .ZN(n6099) );
  OR2_X1 U7773 ( .A1(n10072), .A2(n6461), .ZN(n6098) );
  AND2_X1 U7774 ( .A1(n6099), .A2(n6098), .ZN(n8922) );
  INV_X1 U7775 ( .A(n8922), .ZN(n10034) );
  NOR2_X1 U7776 ( .A1(n10034), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7777 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7778 ( .A1(n8411), .A2(P1_U4006), .ZN(n6100) );
  OAI21_X1 U7779 ( .B1(P1_U4006), .B2(n6101), .A(n6100), .ZN(P1_U3586) );
  INV_X1 U7780 ( .A(n6102), .ZN(n6104) );
  OAI222_X1 U7781 ( .A1(n9781), .A2(n6104), .B1(n9902), .B2(P1_U3084), .C1(
        n6103), .C2(n9777), .ZN(P1_U3344) );
  INV_X1 U7782 ( .A(n6545), .ZN(n8293) );
  OAI222_X1 U7783 ( .A1(n8019), .A2(n6105), .B1(n9221), .B2(n6104), .C1(n8293), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U7784 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6110) );
  NAND2_X1 U7785 ( .A1(n5904), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7786 ( .A1(n4318), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U7787 ( .A1(n4317), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6106) );
  NAND3_X1 U7788 ( .A1(n6108), .A2(n6107), .A3(n6106), .ZN(n8924) );
  NAND2_X1 U7789 ( .A1(P2_U3966), .A2(n8924), .ZN(n6109) );
  OAI21_X1 U7790 ( .B1(P2_U3966), .B2(n6110), .A(n6109), .ZN(P2_U3583) );
  INV_X1 U7791 ( .A(n6111), .ZN(n6113) );
  INV_X1 U7792 ( .A(n6450), .ZN(n6231) );
  OAI222_X1 U7793 ( .A1(n9781), .A2(n6113), .B1(n6231), .B2(P1_U3084), .C1(
        n6112), .C2(n9777), .ZN(P1_U3343) );
  INV_X1 U7794 ( .A(n6547), .ZN(n8282) );
  OAI222_X1 U7795 ( .A1(n8019), .A2(n6114), .B1(n9221), .B2(n6113), .C1(n8282), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U7796 ( .A(n6115), .ZN(n6118) );
  AOI22_X1 U7797 ( .A1(n6606), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n9218), .ZN(n6116) );
  OAI21_X1 U7798 ( .B1(n6118), .B2(n9221), .A(n6116), .ZN(P2_U3347) );
  INV_X1 U7799 ( .A(n6451), .ZN(n9337) );
  OAI222_X1 U7800 ( .A1(n7846), .A2(n6118), .B1(n9337), .B2(P1_U3084), .C1(
        n6117), .C2(n9777), .ZN(P1_U3342) );
  INV_X1 U7801 ( .A(n6119), .ZN(n6329) );
  OR2_X1 U7802 ( .A1(P1_U3083), .A2(n6329), .ZN(n9924) );
  INV_X1 U7803 ( .A(n9924), .ZN(n9882) );
  OR2_X1 U7804 ( .A1(n5433), .A2(P1_U3084), .ZN(n8014) );
  NOR2_X1 U7805 ( .A1(n8588), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6120) );
  INV_X1 U7806 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6126) );
  OAI22_X1 U7807 ( .A1(n8014), .A2(n6120), .B1(P1_U3084), .B2(n6126), .ZN(
        n6328) );
  AND2_X1 U7808 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6319) );
  NAND2_X1 U7809 ( .A1(n6126), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6121) );
  OAI211_X1 U7810 ( .C1(n6319), .C2(n8588), .A(n6147), .B(n6121), .ZN(n6122)
         );
  NAND2_X1 U7811 ( .A1(n6328), .A2(n6122), .ZN(n6124) );
  OAI22_X1 U7812 ( .A1(n6125), .A2(n6124), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6123), .ZN(n6128) );
  INV_X1 U7813 ( .A(n8588), .ZN(n6144) );
  OR3_X1 U7814 ( .A1(n6145), .A2(n8014), .A3(n6144), .ZN(n9876) );
  NOR3_X1 U7815 ( .A1(n9876), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n6126), .ZN(
        n6127) );
  AOI211_X1 U7816 ( .C1(P1_ADDR_REG_0__SCAN_IN), .C2(n9882), .A(n6128), .B(
        n6127), .ZN(n6129) );
  INV_X1 U7817 ( .A(n6129), .ZN(P1_U3241) );
  INV_X1 U7818 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7413) );
  MUX2_X1 U7819 ( .A(n6130), .B(P1_REG2_REG_2__SCAN_IN), .S(n6403), .Z(n6133)
         );
  OR2_X1 U7820 ( .A1(n6150), .A2(n6131), .ZN(n6132) );
  NAND2_X1 U7821 ( .A1(n6187), .A2(n6132), .ZN(n6402) );
  NAND2_X1 U7822 ( .A1(n6133), .A2(n6402), .ZN(n6404) );
  INV_X1 U7823 ( .A(n6403), .ZN(n6410) );
  NAND2_X1 U7824 ( .A1(n6410), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U7825 ( .A1(n6404), .A2(n6174), .ZN(n6136) );
  MUX2_X1 U7826 ( .A(n6134), .B(P1_REG2_REG_3__SCAN_IN), .S(n6173), .Z(n6135)
         );
  NAND2_X1 U7827 ( .A1(n6136), .A2(n6135), .ZN(n6177) );
  INV_X1 U7828 ( .A(n6173), .ZN(n6153) );
  NAND2_X1 U7829 ( .A1(n6153), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7830 ( .A1(n6347), .A2(n6138), .ZN(n6143) );
  OAI21_X1 U7831 ( .B1(n6347), .B2(n6138), .A(n6143), .ZN(n6332) );
  INV_X1 U7832 ( .A(n6332), .ZN(n6139) );
  NAND2_X1 U7833 ( .A1(n6331), .A2(n6139), .ZN(n6335) );
  NAND2_X1 U7834 ( .A1(n6335), .A2(n6143), .ZN(n6140) );
  MUX2_X1 U7835 ( .A(n6201), .B(P1_REG2_REG_5__SCAN_IN), .S(n6202), .Z(n6141)
         );
  NAND2_X1 U7836 ( .A1(n6140), .A2(n6141), .ZN(n6204) );
  INV_X1 U7837 ( .A(n6141), .ZN(n6142) );
  NAND3_X1 U7838 ( .A1(n6335), .A2(n6143), .A3(n6142), .ZN(n6146) );
  NAND2_X1 U7839 ( .A1(n6144), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7941) );
  OR2_X1 U7840 ( .A1(n6145), .A2(n7941), .ZN(n9365) );
  OR2_X1 U7841 ( .A1(n9365), .A2(n5433), .ZN(n9895) );
  AOI21_X1 U7842 ( .B1(n6204), .B2(n6146), .A(n9895), .ZN(n6164) );
  OR2_X1 U7843 ( .A1(n9365), .A2(n6147), .ZN(n9914) );
  INV_X1 U7844 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6148) );
  NOR2_X1 U7845 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6148), .ZN(n7003) );
  INV_X1 U7846 ( .A(n7003), .ZN(n6162) );
  INV_X1 U7847 ( .A(n9876), .ZN(n9920) );
  INV_X1 U7848 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6149) );
  MUX2_X1 U7849 ( .A(n6149), .B(P1_REG1_REG_2__SCAN_IN), .S(n6403), .Z(n6399)
         );
  INV_X1 U7850 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9998) );
  MUX2_X1 U7851 ( .A(n9998), .B(P1_REG1_REG_1__SCAN_IN), .S(n6150), .Z(n6183)
         );
  AND2_X1 U7852 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6182) );
  NAND2_X1 U7853 ( .A1(n6183), .A2(n6182), .ZN(n6181) );
  INV_X1 U7854 ( .A(n6150), .ZN(n6186) );
  NAND2_X1 U7855 ( .A1(n6186), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7856 ( .A1(n6181), .A2(n6151), .ZN(n6398) );
  NAND2_X1 U7857 ( .A1(n6399), .A2(n6398), .ZN(n6397) );
  NAND2_X1 U7858 ( .A1(n6410), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6152) );
  NAND2_X1 U7859 ( .A1(n6397), .A2(n6152), .ZN(n6169) );
  XNOR2_X1 U7860 ( .A(n6173), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n6170) );
  NAND2_X1 U7861 ( .A1(n6169), .A2(n6170), .ZN(n6168) );
  NAND2_X1 U7862 ( .A1(n6153), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6154) );
  AND2_X1 U7863 ( .A1(n6168), .A2(n6154), .ZN(n6337) );
  XNOR2_X1 U7864 ( .A(n6347), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n6338) );
  NAND2_X1 U7865 ( .A1(n6337), .A2(n6338), .ZN(n6342) );
  NAND2_X1 U7866 ( .A1(n6347), .A2(n6155), .ZN(n6156) );
  NAND2_X1 U7867 ( .A1(n6342), .A2(n6156), .ZN(n6159) );
  INV_X1 U7868 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6157) );
  XNOR2_X1 U7869 ( .A(n6202), .B(n6157), .ZN(n6158) );
  OR2_X1 U7870 ( .A1(n6159), .A2(n6158), .ZN(n6196) );
  NAND2_X1 U7871 ( .A1(n6159), .A2(n6158), .ZN(n6160) );
  NAND3_X1 U7872 ( .A1(n9920), .A2(n6196), .A3(n6160), .ZN(n6161) );
  OAI211_X1 U7873 ( .C1(n9914), .C2(n6202), .A(n6162), .B(n6161), .ZN(n6163)
         );
  NOR2_X1 U7874 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  OAI21_X1 U7875 ( .B1(n7413), .B2(n9924), .A(n6165), .ZN(P1_U3246) );
  INV_X1 U7876 ( .A(n6166), .ZN(n6192) );
  AOI22_X1 U7877 ( .A1(n6777), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n9218), .ZN(n6167) );
  OAI21_X1 U7878 ( .B1(n6192), .B2(n9221), .A(n6167), .ZN(P2_U3346) );
  INV_X1 U7879 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6180) );
  OAI211_X1 U7880 ( .C1(n6170), .C2(n6169), .A(n9920), .B(n6168), .ZN(n6171)
         );
  NAND2_X1 U7881 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6628) );
  OAI211_X1 U7882 ( .C1(n9914), .C2(n6173), .A(n6171), .B(n6628), .ZN(n6172)
         );
  INV_X1 U7883 ( .A(n6172), .ZN(n6179) );
  INV_X1 U7884 ( .A(n9895), .ZN(n9911) );
  MUX2_X1 U7885 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6134), .S(n6173), .Z(n6175)
         );
  NAND3_X1 U7886 ( .A1(n6175), .A2(n6404), .A3(n6174), .ZN(n6176) );
  NAND3_X1 U7887 ( .A1(n9911), .A2(n6177), .A3(n6176), .ZN(n6178) );
  OAI211_X1 U7888 ( .C1(n6180), .C2(n9924), .A(n6179), .B(n6178), .ZN(P1_U3244) );
  INV_X1 U7889 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6191) );
  INV_X1 U7890 ( .A(n9914), .ZN(n7225) );
  OAI211_X1 U7891 ( .C1(n6183), .C2(n6182), .A(n9920), .B(n6181), .ZN(n6184)
         );
  OAI21_X1 U7892 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6835), .A(n6184), .ZN(n6185) );
  AOI21_X1 U7893 ( .B1(n6186), .B2(n7225), .A(n6185), .ZN(n6190) );
  OAI211_X1 U7894 ( .C1(n6319), .C2(n6188), .A(n9911), .B(n6187), .ZN(n6189)
         );
  OAI211_X1 U7895 ( .C1(n6191), .C2(n9924), .A(n6190), .B(n6189), .ZN(P1_U3242) );
  INV_X1 U7896 ( .A(n6655), .ZN(n6448) );
  OAI222_X1 U7897 ( .A1(n9771), .A2(n6193), .B1(n9781), .B2(n6192), .C1(
        P1_U3084), .C2(n6448), .ZN(P1_U3341) );
  NAND2_X1 U7898 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7152) );
  XNOR2_X1 U7899 ( .A(n6218), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n6198) );
  INV_X1 U7900 ( .A(n6202), .ZN(n6194) );
  NAND2_X1 U7901 ( .A1(n6194), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6195) );
  AND2_X1 U7902 ( .A1(n6196), .A2(n6195), .ZN(n6197) );
  NAND2_X1 U7903 ( .A1(n6197), .A2(n6198), .ZN(n6214) );
  OAI21_X1 U7904 ( .B1(n6198), .B2(n6197), .A(n6214), .ZN(n6199) );
  NAND2_X1 U7905 ( .A1(n9920), .A2(n6199), .ZN(n6200) );
  OAI211_X1 U7906 ( .C1(n9914), .C2(n6218), .A(n7152), .B(n6200), .ZN(n6209)
         );
  NAND2_X1 U7907 ( .A1(n6202), .A2(n6201), .ZN(n6203) );
  NAND2_X1 U7908 ( .A1(n6204), .A2(n6203), .ZN(n6207) );
  MUX2_X1 U7909 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6217), .S(n6218), .Z(n6206)
         );
  INV_X1 U7910 ( .A(n6220), .ZN(n6205) );
  AOI211_X1 U7911 ( .C1(n6207), .C2(n6206), .A(n6205), .B(n9895), .ZN(n6208)
         );
  AOI211_X1 U7912 ( .C1(P1_ADDR_REG_6__SCAN_IN), .C2(n9882), .A(n6209), .B(
        n6208), .ZN(n6210) );
  INV_X1 U7913 ( .A(n6210), .ZN(P1_U3247) );
  INV_X1 U7914 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7418) );
  NOR2_X1 U7915 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6235), .ZN(n6211) );
  AOI21_X1 U7916 ( .B1(n6235), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6211), .ZN(
        n6216) );
  NAND2_X1 U7917 ( .A1(n6218), .A2(n6212), .ZN(n6213) );
  NAND2_X1 U7918 ( .A1(n6214), .A2(n6213), .ZN(n6215) );
  NAND2_X1 U7919 ( .A1(n6215), .A2(n6216), .ZN(n6230) );
  OAI21_X1 U7920 ( .B1(n6216), .B2(n6215), .A(n6230), .ZN(n6227) );
  OR2_X1 U7921 ( .A1(n6218), .A2(n6217), .ZN(n6219) );
  NAND2_X1 U7922 ( .A1(n6220), .A2(n6219), .ZN(n6222) );
  AOI22_X1 U7923 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6224), .B1(n6235), .B2(
        n7110), .ZN(n6221) );
  NOR2_X1 U7924 ( .A1(n6221), .A2(n6222), .ZN(n6236) );
  AOI21_X1 U7925 ( .B1(n6222), .B2(n6221), .A(n6236), .ZN(n6223) );
  NOR2_X1 U7926 ( .A1(n9895), .A2(n6223), .ZN(n6226) );
  NAND2_X1 U7927 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3084), .ZN(n6890) );
  OAI21_X1 U7928 ( .B1(n9914), .B2(n6224), .A(n6890), .ZN(n6225) );
  AOI211_X1 U7929 ( .C1(n9920), .C2(n6227), .A(n6226), .B(n6225), .ZN(n6228)
         );
  OAI21_X1 U7930 ( .B1(n7418), .B2(n9924), .A(n6228), .ZN(P1_U3248) );
  INV_X1 U7931 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U7932 ( .A1(n6238), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6229) );
  OAI21_X1 U7933 ( .B1(n6238), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6229), .ZN(
        n9878) );
  OAI21_X1 U7934 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n6235), .A(n6230), .ZN(
        n9879) );
  NOR2_X1 U7935 ( .A1(n9878), .A2(n9879), .ZN(n9877) );
  AOI21_X1 U7936 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6238), .A(n9877), .ZN(
        n9894) );
  AOI22_X1 U7937 ( .A1(n6240), .A2(P1_REG1_REG_9__SCAN_IN), .B1(n5045), .B2(
        n9902), .ZN(n9893) );
  NAND2_X1 U7938 ( .A1(n9894), .A2(n9893), .ZN(n9892) );
  OAI21_X1 U7939 ( .B1(n6240), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9892), .ZN(
        n6233) );
  AOI22_X1 U7940 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n6450), .B1(n6231), .B2(
        n5063), .ZN(n6232) );
  NAND2_X1 U7941 ( .A1(n6232), .A2(n6233), .ZN(n6442) );
  OAI21_X1 U7942 ( .B1(n6233), .B2(n6232), .A(n6442), .ZN(n6234) );
  NAND2_X1 U7943 ( .A1(n6234), .A2(n9920), .ZN(n6247) );
  NAND2_X1 U7944 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3084), .ZN(n7371) );
  INV_X1 U7945 ( .A(n7371), .ZN(n6245) );
  NOR2_X1 U7946 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6235), .ZN(n6237) );
  NOR2_X1 U7947 ( .A1(n6237), .A2(n6236), .ZN(n9887) );
  NOR2_X1 U7948 ( .A1(n9883), .A2(n5022), .ZN(n9885) );
  OAI22_X1 U7949 ( .A1(n9887), .A2(n9885), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n6238), .ZN(n9898) );
  NAND2_X1 U7950 ( .A1(n6240), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6239) );
  OAI21_X1 U7951 ( .B1(n6240), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6239), .ZN(
        n9897) );
  NOR2_X1 U7952 ( .A1(n9898), .A2(n9897), .ZN(n9896) );
  NAND2_X1 U7953 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n6450), .ZN(n6241) );
  OAI21_X1 U7954 ( .B1(n6450), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6241), .ZN(
        n6242) );
  AOI211_X1 U7955 ( .C1(n6243), .C2(n6242), .A(n6449), .B(n9895), .ZN(n6244)
         );
  AOI211_X1 U7956 ( .C1(n7225), .C2(n6450), .A(n6245), .B(n6244), .ZN(n6246)
         );
  OAI211_X1 U7957 ( .C1(n9924), .C2(n6248), .A(n6247), .B(n6246), .ZN(P1_U3251) );
  INV_X1 U7958 ( .A(n6249), .ZN(n6313) );
  AOI22_X1 U7959 ( .A1(n7073), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n6744), .ZN(n6250) );
  OAI21_X1 U7960 ( .B1(n6313), .B2(n7846), .A(n6250), .ZN(P1_U3340) );
  INV_X1 U7961 ( .A(n6251), .ZN(n6252) );
  OAI211_X1 U7962 ( .C1(n10072), .C2(n6253), .A(n8251), .B(n6252), .ZN(n6271)
         );
  AND2_X1 U7963 ( .A1(n4739), .A2(n8246), .ZN(n6254) );
  NAND2_X1 U7964 ( .A1(n6271), .A2(n6254), .ZN(n10032) );
  INV_X1 U7965 ( .A(n10032), .ZN(n10027) );
  OR2_X1 U7966 ( .A1(n6541), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U7967 ( .A1(n6541), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U7968 ( .A1(n6256), .A2(n6255), .ZN(n6268) );
  INV_X1 U7969 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6257) );
  XNOR2_X1 U7970 ( .A(n8843), .B(n6257), .ZN(n8852) );
  INV_X1 U7971 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10161) );
  INV_X1 U7972 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6396) );
  MUX2_X1 U7973 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6396), .S(n8830), .Z(n8838)
         );
  AND2_X1 U7974 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n8837) );
  NAND2_X1 U7975 ( .A1(n8838), .A2(n8837), .ZN(n8836) );
  NAND2_X1 U7976 ( .A1(n8830), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6258) );
  NAND2_X1 U7977 ( .A1(n8836), .A2(n6258), .ZN(n6363) );
  NAND2_X1 U7978 ( .A1(n6368), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U7979 ( .A1(n8843), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U7980 ( .A1(n8850), .A2(n6260), .ZN(n8867) );
  INV_X1 U7981 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6261) );
  XNOR2_X1 U7982 ( .A(n8860), .B(n6261), .ZN(n8868) );
  NAND2_X1 U7983 ( .A1(n8867), .A2(n8868), .ZN(n8866) );
  NAND2_X1 U7984 ( .A1(n8860), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6262) );
  NAND2_X1 U7985 ( .A1(n6518), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6264) );
  OAI21_X1 U7986 ( .B1(n6518), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6264), .ZN(
        n6263) );
  INV_X1 U7987 ( .A(n6263), .ZN(n6517) );
  OR2_X1 U7988 ( .A1(n6277), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6266) );
  NAND2_X1 U7989 ( .A1(n6277), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6265) );
  NAND2_X1 U7990 ( .A1(n6266), .A2(n6265), .ZN(n6301) );
  AOI21_X1 U7991 ( .B1(n6277), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6300), .ZN(
        n6267) );
  NOR2_X1 U7992 ( .A1(n6267), .A2(n6268), .ZN(n6540) );
  AOI21_X1 U7993 ( .B1(n6268), .B2(n6267), .A(n6540), .ZN(n6276) );
  INV_X1 U7994 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6270) );
  NOR2_X1 U7995 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5669), .ZN(n6703) );
  INV_X1 U7996 ( .A(n6703), .ZN(n6269) );
  OAI21_X1 U7997 ( .B1(n8922), .B2(n6270), .A(n6269), .ZN(n6275) );
  NAND2_X1 U7998 ( .A1(n6271), .A2(n4739), .ZN(n6272) );
  NAND2_X1 U7999 ( .A1(n8816), .A2(n6272), .ZN(n6295) );
  NAND2_X1 U8000 ( .A1(n6295), .A2(n6293), .ZN(n10030) );
  NOR2_X1 U8001 ( .A1(n10030), .A2(n6273), .ZN(n6274) );
  AOI211_X1 U8002 ( .C1(n10027), .C2(n6276), .A(n6275), .B(n6274), .ZN(n6299)
         );
  NAND2_X1 U8003 ( .A1(n6277), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6290) );
  MUX2_X1 U8004 ( .A(n6899), .B(P2_REG2_REG_6__SCAN_IN), .S(n6277), .Z(n6278)
         );
  INV_X1 U8005 ( .A(n6278), .ZN(n6309) );
  NAND2_X1 U8006 ( .A1(n6518), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6289) );
  INV_X1 U8007 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6285) );
  INV_X1 U8008 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6905) );
  MUX2_X1 U8009 ( .A(n6905), .B(P2_REG2_REG_1__SCAN_IN), .S(n8830), .Z(n8831)
         );
  INV_X1 U8010 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10028) );
  INV_X1 U8011 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10037) );
  NOR3_X1 U8012 ( .A1(n8831), .A2(n10028), .A3(n10037), .ZN(n8832) );
  NOR2_X1 U8013 ( .A1(n6279), .A2(n6905), .ZN(n6369) );
  INV_X1 U8014 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6280) );
  MUX2_X1 U8015 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6280), .S(n6368), .Z(n6281)
         );
  OAI21_X1 U8016 ( .B1(n8832), .B2(n6369), .A(n6281), .ZN(n8848) );
  NAND2_X1 U8017 ( .A1(n6368), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8847) );
  INV_X1 U8018 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10060) );
  MUX2_X1 U8019 ( .A(n10060), .B(P2_REG2_REG_3__SCAN_IN), .S(n8843), .Z(n8846)
         );
  AOI21_X1 U8020 ( .B1(n8848), .B2(n8847), .A(n8846), .ZN(n8845) );
  NOR2_X1 U8021 ( .A1(n6282), .A2(n10060), .ZN(n8859) );
  MUX2_X1 U8022 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6285), .S(n8860), .Z(n6283)
         );
  OAI21_X1 U8023 ( .B1(n8845), .B2(n8859), .A(n6283), .ZN(n8865) );
  OAI21_X1 U8024 ( .B1(n6285), .B2(n6284), .A(n8865), .ZN(n6514) );
  INV_X1 U8025 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6286) );
  MUX2_X1 U8026 ( .A(n6286), .B(P2_REG2_REG_5__SCAN_IN), .S(n6518), .Z(n6513)
         );
  INV_X1 U8027 ( .A(n6513), .ZN(n6287) );
  NAND2_X1 U8028 ( .A1(n6514), .A2(n6287), .ZN(n6288) );
  NAND2_X1 U8029 ( .A1(n6289), .A2(n6288), .ZN(n6310) );
  NAND2_X1 U8030 ( .A1(n6309), .A2(n6310), .ZN(n6308) );
  NAND2_X1 U8031 ( .A1(n6290), .A2(n6308), .ZN(n6297) );
  INV_X1 U8032 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6291) );
  MUX2_X1 U8033 ( .A(n6291), .B(P2_REG2_REG_7__SCAN_IN), .S(n6541), .Z(n6292)
         );
  INV_X1 U8034 ( .A(n6292), .ZN(n6296) );
  NOR2_X1 U8035 ( .A1(n6293), .A2(n8246), .ZN(n6294) );
  NAND2_X1 U8036 ( .A1(n6296), .A2(n6297), .ZN(n6532) );
  OAI211_X1 U8037 ( .C1(n6297), .C2(n6296), .A(n10029), .B(n6532), .ZN(n6298)
         );
  NAND2_X1 U8038 ( .A1(n6299), .A2(n6298), .ZN(P2_U3252) );
  AOI21_X1 U8039 ( .B1(n6302), .B2(n6301), .A(n6300), .ZN(n6307) );
  INV_X1 U8040 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6304) );
  NOR2_X1 U8041 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7572), .ZN(n10016) );
  INV_X1 U8042 ( .A(n10016), .ZN(n6303) );
  OAI21_X1 U8043 ( .B1(n8922), .B2(n6304), .A(n6303), .ZN(n6306) );
  NOR2_X1 U8044 ( .A1(n10030), .A2(n4740), .ZN(n6305) );
  AOI211_X1 U8045 ( .C1(n10027), .C2(n6307), .A(n6306), .B(n6305), .ZN(n6312)
         );
  OAI211_X1 U8046 ( .C1(n6310), .C2(n6309), .A(n10029), .B(n6308), .ZN(n6311)
         );
  NAND2_X1 U8047 ( .A1(n6312), .A2(n6311), .ZN(P2_U3251) );
  INV_X1 U8048 ( .A(n6937), .ZN(n6775) );
  OAI222_X1 U8049 ( .A1(n8019), .A2(n6314), .B1(n9221), .B2(n6313), .C1(n6775), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8050 ( .A(n6315), .ZN(n6317) );
  INV_X1 U8051 ( .A(n7220), .ZN(n7212) );
  OAI222_X1 U8052 ( .A1(n7846), .A2(n6317), .B1(n7212), .B2(P1_U3084), .C1(
        n6316), .C2(n9777), .ZN(P1_U3339) );
  INV_X1 U8053 ( .A(n7267), .ZN(n7271) );
  OAI222_X1 U8054 ( .A1(n8019), .A2(n6318), .B1(n9221), .B2(n6317), .C1(n7271), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8055 ( .A(n6319), .ZN(n6327) );
  OR2_X2 U8056 ( .A1(n7279), .A2(n6323), .ZN(n8718) );
  OR2_X4 U8057 ( .A1(n8718), .A2(n6320), .ZN(n8719) );
  INV_X2 U8058 ( .A(n8719), .ZN(n6414) );
  NAND2_X1 U8059 ( .A1(n9331), .A2(n6414), .ZN(n6322) );
  AND2_X1 U8060 ( .A1(n7279), .A2(n6624), .ZN(n6615) );
  AOI22_X1 U8061 ( .A1(n9932), .A2(n8706), .B1(n6323), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n6321) );
  NAND2_X1 U8062 ( .A1(n9331), .A2(n6884), .ZN(n6325) );
  INV_X2 U8063 ( .A(n8718), .ZN(n8714) );
  AOI22_X1 U8064 ( .A1(n9932), .A2(n8714), .B1(n6323), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n6324) );
  NAND2_X1 U8065 ( .A1(n6325), .A2(n6324), .ZN(n6417) );
  NAND2_X1 U8066 ( .A1(n6326), .A2(n6417), .ZN(n6421) );
  OAI21_X1 U8067 ( .B1(n6326), .B2(n6417), .A(n6421), .ZN(n6358) );
  MUX2_X1 U8068 ( .A(n6327), .B(n6358), .S(n8588), .Z(n6330) );
  OAI211_X1 U8069 ( .C1(n6330), .C2(n5433), .A(n6329), .B(n6328), .ZN(n6411)
         );
  INV_X1 U8070 ( .A(n6331), .ZN(n6333) );
  NAND2_X1 U8071 ( .A1(n6333), .A2(n6332), .ZN(n6334) );
  NAND2_X1 U8072 ( .A1(n6335), .A2(n6334), .ZN(n6336) );
  NAND2_X1 U8073 ( .A1(n9911), .A2(n6336), .ZN(n6346) );
  INV_X1 U8074 ( .A(n6337), .ZN(n6340) );
  INV_X1 U8075 ( .A(n6338), .ZN(n6339) );
  NAND2_X1 U8076 ( .A1(n6340), .A2(n6339), .ZN(n6341) );
  NAND2_X1 U8077 ( .A1(n6342), .A2(n6341), .ZN(n6344) );
  NOR2_X1 U8078 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6343), .ZN(n6760) );
  AOI21_X1 U8079 ( .B1(n9920), .B2(n6344), .A(n6760), .ZN(n6345) );
  OAI211_X1 U8080 ( .C1(n9914), .C2(n6347), .A(n6346), .B(n6345), .ZN(n6348)
         );
  AOI21_X1 U8081 ( .B1(n9882), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6348), .ZN(
        n6349) );
  NAND2_X1 U8082 ( .A1(n6411), .A2(n6349), .ZN(P1_U3245) );
  INV_X1 U8083 ( .A(n6350), .ZN(n6823) );
  NAND2_X1 U8084 ( .A1(n6823), .A2(n6351), .ZN(n6357) );
  AND2_X1 U8085 ( .A1(n6352), .A2(n6357), .ZN(n6626) );
  INV_X1 U8086 ( .A(n6626), .ZN(n6353) );
  NAND2_X1 U8087 ( .A1(n6353), .A2(n6825), .ZN(n7653) );
  INV_X1 U8088 ( .A(n9969), .ZN(n9988) );
  INV_X1 U8089 ( .A(n9320), .ZN(n7364) );
  INV_X1 U8090 ( .A(n7279), .ZN(n6418) );
  OR2_X1 U8091 ( .A1(n6419), .A2(n6418), .ZN(n9925) );
  INV_X1 U8092 ( .A(n6355), .ZN(n8589) );
  OR3_X1 U8093 ( .A1(n9925), .A2(n6357), .A3(n8589), .ZN(n6437) );
  INV_X1 U8094 ( .A(n6437), .ZN(n6354) );
  NAND2_X1 U8095 ( .A1(n6354), .A2(n5433), .ZN(n9304) );
  INV_X1 U8096 ( .A(n9304), .ZN(n9311) );
  AOI22_X1 U8097 ( .A1(n7653), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n9311), .B2(
        n6423), .ZN(n6360) );
  NAND2_X1 U8098 ( .A1(n8460), .A2(n6355), .ZN(n6356) );
  INV_X1 U8099 ( .A(n9315), .ZN(n6757) );
  NAND2_X1 U8100 ( .A1(n6358), .A2(n6757), .ZN(n6359) );
  OAI211_X1 U8101 ( .C1(n7364), .C2(n8427), .A(n6360), .B(n6359), .ZN(P1_U3230) );
  INV_X1 U8102 ( .A(n10030), .ZN(n8896) );
  INV_X1 U8103 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6361) );
  INV_X1 U8104 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7490) );
  OAI22_X1 U8105 ( .A1(n8922), .A2(n6361), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7490), .ZN(n6367) );
  OAI21_X1 U8106 ( .B1(n6364), .B2(n6363), .A(n6362), .ZN(n6365) );
  NOR2_X1 U8107 ( .A1(n10032), .A2(n6365), .ZN(n6366) );
  AOI211_X1 U8108 ( .C1(n8896), .C2(n6368), .A(n6367), .B(n6366), .ZN(n6374)
         );
  MUX2_X1 U8109 ( .A(n6280), .B(P2_REG2_REG_2__SCAN_IN), .S(n6368), .Z(n6371)
         );
  INV_X1 U8110 ( .A(n6369), .ZN(n6370) );
  NAND2_X1 U8111 ( .A1(n6371), .A2(n6370), .ZN(n6372) );
  OAI211_X1 U8112 ( .C1(n8832), .C2(n6372), .A(n10029), .B(n8848), .ZN(n6373)
         );
  NAND2_X1 U8113 ( .A1(n6374), .A2(n6373), .ZN(P2_U3247) );
  INV_X1 U8114 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6392) );
  INV_X1 U8115 ( .A(n10146), .ZN(n10155) );
  NAND2_X1 U8116 ( .A1(n8092), .A2(n6375), .ZN(n8206) );
  INV_X1 U8117 ( .A(n6376), .ZN(n6916) );
  XNOR2_X1 U8118 ( .A(n8206), .B(n6916), .ZN(n6911) );
  INV_X1 U8119 ( .A(n6946), .ZN(n6378) );
  AOI21_X1 U8120 ( .B1(n6910), .B2(n6919), .A(n10055), .ZN(n6377) );
  NAND2_X1 U8121 ( .A1(n6378), .A2(n6377), .ZN(n6906) );
  OAI21_X1 U8122 ( .B1(n6379), .B2(n10150), .A(n6906), .ZN(n6390) );
  INV_X1 U8123 ( .A(n6375), .ZN(n6383) );
  INV_X1 U8124 ( .A(n6691), .ZN(n6381) );
  NAND2_X1 U8125 ( .A1(n8206), .A2(n6381), .ZN(n6382) );
  OAI211_X1 U8126 ( .C1(n6380), .C2(n6383), .A(n10049), .B(n6382), .ZN(n6389)
         );
  NAND2_X1 U8127 ( .A1(n6384), .A2(n10045), .ZN(n6387) );
  NAND2_X1 U8128 ( .A1(n6385), .A2(n10046), .ZN(n6386) );
  NAND2_X1 U8129 ( .A1(n6387), .A2(n6386), .ZN(n6475) );
  INV_X1 U8130 ( .A(n6475), .ZN(n6388) );
  NAND2_X1 U8131 ( .A1(n6389), .A2(n6388), .ZN(n6909) );
  AOI211_X1 U8132 ( .C1(n10155), .C2(n6911), .A(n6390), .B(n6909), .ZN(n6394)
         );
  OR2_X1 U8133 ( .A1(n6394), .A2(n10156), .ZN(n6391) );
  OAI21_X1 U8134 ( .B1(n10158), .B2(n6392), .A(n6391), .ZN(P2_U3454) );
  INV_X1 U8135 ( .A(n6480), .ZN(n6459) );
  INV_X2 U8136 ( .A(n10174), .ZN(n10176) );
  OR2_X1 U8137 ( .A1(n6394), .A2(n10174), .ZN(n6395) );
  OAI21_X1 U8138 ( .B1(n10176), .B2(n6396), .A(n6395), .ZN(P2_U3521) );
  INV_X1 U8139 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6413) );
  OAI211_X1 U8140 ( .C1(n6399), .C2(n6398), .A(n9920), .B(n6397), .ZN(n6400)
         );
  OAI21_X1 U8141 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6401), .A(n6400), .ZN(n6409) );
  INV_X1 U8142 ( .A(n6402), .ZN(n6407) );
  MUX2_X1 U8143 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6130), .S(n6403), .Z(n6406)
         );
  INV_X1 U8144 ( .A(n6404), .ZN(n6405) );
  AOI211_X1 U8145 ( .C1(n6407), .C2(n6406), .A(n6405), .B(n9895), .ZN(n6408)
         );
  AOI211_X1 U8146 ( .C1(n7225), .C2(n6410), .A(n6409), .B(n6408), .ZN(n6412)
         );
  OAI211_X1 U8147 ( .C1(n9924), .C2(n6413), .A(n6412), .B(n6411), .ZN(P1_U3243) );
  NAND2_X1 U8148 ( .A1(n6423), .A2(n6414), .ZN(n6416) );
  NAND2_X1 U8149 ( .A1(n6839), .A2(n6884), .ZN(n6415) );
  NAND2_X1 U8150 ( .A1(n6416), .A2(n6415), .ZN(n6432) );
  INV_X1 U8151 ( .A(n6432), .ZN(n6435) );
  INV_X1 U8152 ( .A(n6417), .ZN(n6420) );
  NAND2_X1 U8153 ( .A1(n6420), .A2(n8721), .ZN(n6422) );
  INV_X1 U8154 ( .A(n6430), .ZN(n6427) );
  NAND2_X1 U8155 ( .A1(n6423), .A2(n6884), .ZN(n6425) );
  NAND2_X1 U8156 ( .A1(n6839), .A2(n8714), .ZN(n6424) );
  NAND2_X1 U8157 ( .A1(n6425), .A2(n6424), .ZN(n6426) );
  INV_X1 U8158 ( .A(n6429), .ZN(n6428) );
  NAND2_X1 U8159 ( .A1(n6427), .A2(n6428), .ZN(n6492) );
  XNOR2_X1 U8160 ( .A(n6430), .B(n6428), .ZN(n6433) );
  NAND2_X1 U8161 ( .A1(n6430), .A2(n6429), .ZN(n6431) );
  NAND2_X1 U8162 ( .A1(n6431), .A2(n6432), .ZN(n6493) );
  OAI21_X1 U8163 ( .B1(n6433), .B2(n6432), .A(n6493), .ZN(n6434) );
  OAI21_X1 U8164 ( .B1(n6435), .B2(n6492), .A(n6434), .ZN(n6436) );
  NAND2_X1 U8165 ( .A1(n6436), .A2(n6757), .ZN(n6441) );
  NOR2_X1 U8166 ( .A1(n6437), .A2(n5433), .ZN(n9310) );
  INV_X1 U8167 ( .A(n9310), .ZN(n9272) );
  INV_X1 U8168 ( .A(n9331), .ZN(n6438) );
  OAI22_X1 U8169 ( .A1(n9272), .A2(n6438), .B1(n8547), .B2(n9304), .ZN(n6439)
         );
  AOI21_X1 U8170 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n7653), .A(n6439), .ZN(
        n6440) );
  OAI211_X1 U8171 ( .C1(n9943), .C2(n7364), .A(n6441), .B(n6440), .ZN(P1_U3220) );
  AOI22_X1 U8172 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n6451), .B1(n9337), .B2(
        n5079), .ZN(n9334) );
  OAI21_X1 U8173 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n6450), .A(n6442), .ZN(
        n9333) );
  NAND2_X1 U8174 ( .A1(n9334), .A2(n9333), .ZN(n9332) );
  OAI21_X1 U8175 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n6451), .A(n9332), .ZN(
        n6446) );
  NOR2_X1 U8176 ( .A1(n6448), .A2(n6443), .ZN(n6444) );
  AOI21_X1 U8177 ( .B1(n6443), .B2(n6448), .A(n6444), .ZN(n6445) );
  NAND2_X1 U8178 ( .A1(n6445), .A2(n6446), .ZN(n6647) );
  OAI21_X1 U8179 ( .B1(n6446), .B2(n6445), .A(n6647), .ZN(n6457) );
  NAND2_X1 U8180 ( .A1(n9882), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6447) );
  NAND2_X1 U8181 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n7651) );
  OAI211_X1 U8182 ( .C1(n9914), .C2(n6448), .A(n6447), .B(n7651), .ZN(n6456)
         );
  AOI22_X1 U8183 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n6451), .B1(n9337), .B2(
        n5082), .ZN(n9342) );
  OAI21_X1 U8184 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6451), .A(n9340), .ZN(
        n6454) );
  NAND2_X1 U8185 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6655), .ZN(n6452) );
  OAI21_X1 U8186 ( .B1(n6655), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6452), .ZN(
        n6453) );
  NOR2_X1 U8187 ( .A1(n6453), .A2(n6454), .ZN(n6654) );
  AOI211_X1 U8188 ( .C1(n6454), .C2(n6453), .A(n6654), .B(n9895), .ZN(n6455)
         );
  AOI211_X1 U8189 ( .C1(n9920), .C2(n6457), .A(n6456), .B(n6455), .ZN(n6458)
         );
  INV_X1 U8190 ( .A(n6458), .ZN(P1_U3253) );
  NOR2_X1 U8191 ( .A1(n6459), .A2(n10072), .ZN(n6460) );
  AND2_X1 U8192 ( .A1(n6481), .A2(n6460), .ZN(n6478) );
  AND2_X1 U8193 ( .A1(n10150), .A2(n6461), .ZN(n6462) );
  NAND2_X1 U8194 ( .A1(n6478), .A2(n6462), .ZN(n8812) );
  INV_X1 U8195 ( .A(n8812), .ZN(n10022) );
  NAND3_X1 U8196 ( .A1(n8239), .A2(n10081), .A3(n8242), .ZN(n6465) );
  NAND2_X4 U8197 ( .A1(n6465), .A2(n6464), .ZN(n8631) );
  XNOR2_X1 U8198 ( .A(n6910), .B(n8631), .ZN(n6467) );
  NAND2_X1 U8199 ( .A1(n6466), .A2(n6467), .ZN(n6470) );
  INV_X1 U8200 ( .A(n6467), .ZN(n6468) );
  NAND2_X1 U8201 ( .A1(n6469), .A2(n6468), .ZN(n6487) );
  NOR2_X1 U8202 ( .A1(n8631), .A2(n6919), .ZN(n6471) );
  AOI21_X1 U8203 ( .B1(n6376), .B2(n10055), .A(n6471), .ZN(n6472) );
  NAND2_X1 U8204 ( .A1(n6472), .A2(n6473), .ZN(n6488) );
  OAI21_X1 U8205 ( .B1(n6473), .B2(n6472), .A(n6488), .ZN(n6476) );
  NAND2_X1 U8206 ( .A1(n6478), .A2(n6474), .ZN(n8637) );
  INV_X1 U8207 ( .A(n8637), .ZN(n10018) );
  AOI22_X1 U8208 ( .A1(n10022), .A2(n6476), .B1(n10018), .B2(n6475), .ZN(n6486) );
  NAND2_X1 U8209 ( .A1(n6478), .A2(n6477), .ZN(n6479) );
  NAND2_X1 U8210 ( .A1(n6479), .A2(n8975), .ZN(n8809) );
  NAND2_X1 U8211 ( .A1(n6481), .A2(n6480), .ZN(n6483) );
  NAND2_X1 U8212 ( .A1(n6483), .A2(n6482), .ZN(n6582) );
  INV_X1 U8213 ( .A(n8247), .ZN(n6484) );
  NAND2_X1 U8214 ( .A1(n6582), .A2(n6484), .ZN(n6695) );
  AOI22_X1 U8215 ( .A1(n8809), .A2(n6910), .B1(n6695), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n6485) );
  NAND2_X1 U8216 ( .A1(n6486), .A2(n6485), .ZN(P2_U3224) );
  NAND2_X1 U8217 ( .A1(n6488), .A2(n6487), .ZN(n6562) );
  NAND2_X1 U8218 ( .A1(n6385), .A2(n10055), .ZN(n6559) );
  XNOR2_X1 U8219 ( .A(n8631), .B(n10086), .ZN(n6560) );
  XNOR2_X1 U8220 ( .A(n6559), .B(n6560), .ZN(n6561) );
  XNOR2_X1 U8221 ( .A(n6562), .B(n6561), .ZN(n6491) );
  NAND2_X1 U8222 ( .A1(n10018), .A2(n10045), .ZN(n8805) );
  INV_X1 U8223 ( .A(n8805), .ZN(n7206) );
  INV_X1 U8224 ( .A(n10046), .ZN(n9076) );
  INV_X1 U8225 ( .A(n8781), .ZN(n8808) );
  AOI22_X1 U8226 ( .A1(n7206), .A2(n6463), .B1(n8808), .B2(n5620), .ZN(n6490)
         );
  AOI22_X1 U8227 ( .A1(n8809), .A2(n6949), .B1(n6695), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n6489) );
  OAI211_X1 U8228 ( .C1(n6491), .C2(n8812), .A(n6490), .B(n6489), .ZN(P2_U3239) );
  NAND2_X1 U8229 ( .A1(n6493), .A2(n6492), .ZN(n6507) );
  NAND2_X1 U8230 ( .A1(n9329), .A2(n6884), .ZN(n6496) );
  NAND2_X1 U8231 ( .A1(n6494), .A2(n8714), .ZN(n6495) );
  NAND2_X1 U8232 ( .A1(n6496), .A2(n6495), .ZN(n6497) );
  XNOR2_X1 U8233 ( .A(n6497), .B(n8689), .ZN(n6501) );
  AND2_X1 U8234 ( .A1(n6494), .A2(n8706), .ZN(n6499) );
  AOI21_X1 U8235 ( .B1(n9329), .B2(n6414), .A(n6499), .ZN(n6500) );
  OR2_X1 U8236 ( .A1(n6501), .A2(n6500), .ZN(n6502) );
  NAND2_X1 U8237 ( .A1(n6501), .A2(n6500), .ZN(n6619) );
  NAND2_X1 U8238 ( .A1(n6502), .A2(n6619), .ZN(n6506) );
  NAND2_X1 U8239 ( .A1(n6504), .A2(n6503), .ZN(n6620) );
  INV_X1 U8240 ( .A(n6620), .ZN(n6505) );
  AOI21_X1 U8241 ( .B1(n6507), .B2(n6506), .A(n6505), .ZN(n6512) );
  OAI22_X1 U8242 ( .A1(n9272), .A2(n6508), .B1(n7095), .B2(n9304), .ZN(n6510)
         );
  NOR2_X1 U8243 ( .A1(n7364), .A2(n6925), .ZN(n6509) );
  AOI211_X1 U8244 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(n7653), .A(n6510), .B(
        n6509), .ZN(n6511) );
  OAI21_X1 U8245 ( .B1(n6512), .B2(n9315), .A(n6511), .ZN(P1_U3235) );
  XNOR2_X1 U8246 ( .A(n6514), .B(n6513), .ZN(n6524) );
  OAI21_X1 U8247 ( .B1(n6517), .B2(n6516), .A(n6515), .ZN(n6522) );
  NAND2_X1 U8248 ( .A1(n8896), .A2(n6518), .ZN(n6521) );
  INV_X1 U8249 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7448) );
  NOR2_X1 U8250 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7448), .ZN(n6519) );
  AOI21_X1 U8251 ( .B1(n10034), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6519), .ZN(
        n6520) );
  OAI211_X1 U8252 ( .C1(n10032), .C2(n6522), .A(n6521), .B(n6520), .ZN(n6523)
         );
  AOI21_X1 U8253 ( .B1(n10029), .B2(n6524), .A(n6523), .ZN(n6525) );
  INV_X1 U8254 ( .A(n6525), .ZN(P2_U3250) );
  NAND2_X1 U8255 ( .A1(n6547), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6536) );
  INV_X1 U8256 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6526) );
  MUX2_X1 U8257 ( .A(n6526), .B(P2_REG2_REG_10__SCAN_IN), .S(n6547), .Z(n6527)
         );
  INV_X1 U8258 ( .A(n6527), .ZN(n8278) );
  NAND2_X1 U8259 ( .A1(n6545), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6535) );
  INV_X1 U8260 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6528) );
  MUX2_X1 U8261 ( .A(n6528), .B(P2_REG2_REG_9__SCAN_IN), .S(n6545), .Z(n6529)
         );
  INV_X1 U8262 ( .A(n6529), .ZN(n8289) );
  NAND2_X1 U8263 ( .A1(n8874), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6534) );
  INV_X1 U8264 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6530) );
  MUX2_X1 U8265 ( .A(n6530), .B(P2_REG2_REG_8__SCAN_IN), .S(n8874), .Z(n6531)
         );
  INV_X1 U8266 ( .A(n6531), .ZN(n8876) );
  NAND2_X1 U8267 ( .A1(n6541), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6533) );
  NAND2_X1 U8268 ( .A1(n6533), .A2(n6532), .ZN(n8877) );
  NAND2_X1 U8269 ( .A1(n8876), .A2(n8877), .ZN(n8875) );
  NAND2_X1 U8270 ( .A1(n6534), .A2(n8875), .ZN(n8290) );
  NAND2_X1 U8271 ( .A1(n8289), .A2(n8290), .ZN(n8288) );
  NAND2_X1 U8272 ( .A1(n6535), .A2(n8288), .ZN(n8279) );
  NAND2_X1 U8273 ( .A1(n8278), .A2(n8279), .ZN(n8277) );
  NAND2_X1 U8274 ( .A1(n6536), .A2(n8277), .ZN(n6539) );
  INV_X1 U8275 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6537) );
  MUX2_X1 U8276 ( .A(n6537), .B(P2_REG2_REG_11__SCAN_IN), .S(n6606), .Z(n6538)
         );
  NOR2_X1 U8277 ( .A1(n6539), .A2(n6538), .ZN(n6607) );
  AOI21_X1 U8278 ( .B1(n6539), .B2(n6538), .A(n6607), .ZN(n6554) );
  INV_X1 U8279 ( .A(n10029), .ZN(n7886) );
  AND2_X1 U8280 ( .A1(P2_U3152), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8794) );
  OR2_X1 U8281 ( .A1(n8874), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6543) );
  NAND2_X1 U8282 ( .A1(n8874), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6542) );
  NAND2_X1 U8283 ( .A1(n6543), .A2(n6542), .ZN(n8881) );
  INV_X1 U8284 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6544) );
  MUX2_X1 U8285 ( .A(n6544), .B(P2_REG1_REG_9__SCAN_IN), .S(n6545), .Z(n8284)
         );
  AOI21_X1 U8286 ( .B1(n6545), .B2(P2_REG1_REG_9__SCAN_IN), .A(n8283), .ZN(
        n8274) );
  INV_X1 U8287 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6546) );
  MUX2_X1 U8288 ( .A(n6546), .B(P2_REG1_REG_10__SCAN_IN), .S(n6547), .Z(n8273)
         );
  INV_X1 U8289 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6548) );
  MUX2_X1 U8290 ( .A(n6548), .B(P2_REG1_REG_11__SCAN_IN), .S(n6606), .Z(n6549)
         );
  AOI211_X1 U8291 ( .C1(n6550), .C2(n6549), .A(n6598), .B(n10032), .ZN(n6551)
         );
  AOI211_X1 U8292 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n10034), .A(n8794), .B(
        n6551), .ZN(n6553) );
  NAND2_X1 U8293 ( .A1(n8896), .A2(n6606), .ZN(n6552) );
  OAI211_X1 U8294 ( .C1(n6554), .C2(n7886), .A(n6553), .B(n6552), .ZN(P2_U3256) );
  INV_X1 U8295 ( .A(n6555), .ZN(n6557) );
  OAI222_X1 U8296 ( .A1(n9771), .A2(n6556), .B1(n7846), .B2(n6557), .C1(
        P1_U3084), .C2(n7668), .ZN(P1_U3338) );
  INV_X1 U8297 ( .A(n7866), .ZN(n7873) );
  OAI222_X1 U8298 ( .A1(n8019), .A2(n6558), .B1(n9221), .B2(n6557), .C1(
        P2_U3152), .C2(n7873), .ZN(P2_U3343) );
  OAI22_X1 U8299 ( .A1(n8805), .A2(n6961), .B1(n8781), .B2(n6962), .ZN(n6588)
         );
  NAND2_X1 U8300 ( .A1(n5620), .A2(n10055), .ZN(n6563) );
  XNOR2_X1 U8301 ( .A(n10056), .B(n8631), .ZN(n6564) );
  XNOR2_X1 U8302 ( .A(n6563), .B(n6564), .ZN(n6707) );
  NAND2_X1 U8303 ( .A1(n6708), .A2(n6707), .ZN(n6567) );
  INV_X1 U8304 ( .A(n6563), .ZN(n6565) );
  NAND2_X1 U8305 ( .A1(n6565), .A2(n6564), .ZN(n6566) );
  NAND2_X1 U8306 ( .A1(n6567), .A2(n6566), .ZN(n6576) );
  INV_X1 U8307 ( .A(n6576), .ZN(n6574) );
  AND2_X1 U8308 ( .A1(n10047), .A2(n10055), .ZN(n6568) );
  XNOR2_X1 U8309 ( .A(n6970), .B(n8631), .ZN(n6569) );
  NAND2_X1 U8310 ( .A1(n6568), .A2(n6569), .ZN(n6572) );
  INV_X1 U8311 ( .A(n6568), .ZN(n6571) );
  INV_X1 U8312 ( .A(n6569), .ZN(n6570) );
  NAND2_X1 U8313 ( .A1(n6571), .A2(n6570), .ZN(n6589) );
  NAND2_X1 U8314 ( .A1(n6572), .A2(n6589), .ZN(n6575) );
  INV_X1 U8315 ( .A(n6575), .ZN(n6573) );
  NAND2_X1 U8316 ( .A1(n6574), .A2(n6573), .ZN(n6590) );
  NAND2_X1 U8317 ( .A1(n6576), .A2(n6575), .ZN(n6577) );
  AOI21_X1 U8318 ( .B1(n6590), .B2(n6577), .A(n8812), .ZN(n6587) );
  AND3_X1 U8319 ( .A1(n6580), .A2(n6579), .A3(n6578), .ZN(n6581) );
  NAND2_X1 U8320 ( .A1(n6582), .A2(n6581), .ZN(n6583) );
  NAND2_X1 U8321 ( .A1(n6583), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10026) );
  NOR2_X1 U8322 ( .A1(n7571), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8858) );
  INV_X1 U8323 ( .A(n8858), .ZN(n6585) );
  NAND2_X1 U8324 ( .A1(n8809), .A2(n6970), .ZN(n6584) );
  OAI211_X1 U8325 ( .C1(n10026), .C2(n6965), .A(n6585), .B(n6584), .ZN(n6586)
         );
  OR3_X1 U8326 ( .A1(n6588), .A2(n6587), .A3(n6586), .ZN(P2_U3232) );
  NAND2_X1 U8327 ( .A1(n6590), .A2(n6589), .ZN(n6683) );
  XNOR2_X1 U8328 ( .A(n6736), .B(n8606), .ZN(n6669) );
  NAND2_X1 U8329 ( .A1(n8829), .A2(n10055), .ZN(n6668) );
  XNOR2_X1 U8330 ( .A(n6669), .B(n6668), .ZN(n10008) );
  XNOR2_X1 U8331 ( .A(n10009), .B(n10008), .ZN(n6596) );
  INV_X1 U8332 ( .A(n10026), .ZN(n8784) );
  NAND2_X1 U8333 ( .A1(n8809), .A2(n6736), .ZN(n6591) );
  OAI21_X1 U8334 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n7448), .A(n6591), .ZN(n6594) );
  OAI22_X1 U8335 ( .A1(n8805), .A2(n6709), .B1(n8781), .B2(n6592), .ZN(n6593)
         );
  AOI211_X1 U8336 ( .C1(n6843), .C2(n8784), .A(n6594), .B(n6593), .ZN(n6595)
         );
  OAI21_X1 U8337 ( .B1(n6596), .B2(n8812), .A(n6595), .ZN(P2_U3229) );
  INV_X1 U8338 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6597) );
  MUX2_X1 U8339 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6597), .S(n6777), .Z(n6599)
         );
  NAND2_X1 U8340 ( .A1(n4352), .A2(n6599), .ZN(n6776) );
  OAI21_X1 U8341 ( .B1(n6599), .B2(n4352), .A(n6776), .ZN(n6605) );
  INV_X1 U8342 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6601) );
  OR2_X1 U8343 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7059), .ZN(n6600) );
  OAI21_X1 U8344 ( .B1(n8922), .B2(n6601), .A(n6600), .ZN(n6604) );
  INV_X1 U8345 ( .A(n6777), .ZN(n6602) );
  NOR2_X1 U8346 ( .A1(n10030), .A2(n6602), .ZN(n6603) );
  AOI211_X1 U8347 ( .C1(n10027), .C2(n6605), .A(n6604), .B(n6603), .ZN(n6614)
         );
  INV_X1 U8348 ( .A(n6606), .ZN(n6608) );
  AOI21_X1 U8349 ( .B1(n6608), .B2(n6537), .A(n6607), .ZN(n6612) );
  INV_X1 U8350 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6609) );
  MUX2_X1 U8351 ( .A(n6609), .B(P2_REG2_REG_12__SCAN_IN), .S(n6777), .Z(n6610)
         );
  INV_X1 U8352 ( .A(n6610), .ZN(n6611) );
  NAND2_X1 U8353 ( .A1(n6611), .A2(n6612), .ZN(n6770) );
  OAI211_X1 U8354 ( .C1(n6612), .C2(n6611), .A(n10029), .B(n6770), .ZN(n6613)
         );
  NAND2_X1 U8355 ( .A1(n6614), .A2(n6613), .ZN(P2_U3257) );
  OAI22_X1 U8356 ( .A1(n7095), .A2(n6498), .B1(n6726), .B2(n8718), .ZN(n6616)
         );
  XNOR2_X1 U8357 ( .A(n6616), .B(n8689), .ZN(n6750) );
  OR2_X1 U8358 ( .A1(n7095), .A2(n8719), .ZN(n6618) );
  NAND2_X1 U8359 ( .A1(n7124), .A2(n6884), .ZN(n6617) );
  NAND2_X1 U8360 ( .A1(n6618), .A2(n6617), .ZN(n6748) );
  XNOR2_X1 U8361 ( .A(n6750), .B(n6748), .ZN(n6622) );
  NAND2_X1 U8362 ( .A1(n6620), .A2(n6619), .ZN(n6621) );
  OAI21_X1 U8363 ( .B1(n6622), .B2(n6621), .A(n6756), .ZN(n6623) );
  NAND2_X1 U8364 ( .A1(n6623), .A2(n6757), .ZN(n6634) );
  NAND3_X1 U8365 ( .A1(n6625), .A2(n6624), .A3(n7660), .ZN(n6627) );
  AOI21_X1 U8366 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6627), .A(n6626), .ZN(n9262) );
  INV_X1 U8367 ( .A(n9262), .ZN(n9306) );
  INV_X1 U8368 ( .A(n6628), .ZN(n6629) );
  AOI21_X1 U8369 ( .B1(n9302), .B2(n9329), .A(n6629), .ZN(n6630) );
  OAI21_X1 U8370 ( .B1(n6855), .B2(n9304), .A(n6630), .ZN(n6631) );
  AOI21_X1 U8371 ( .B1(n9306), .B2(n6632), .A(n6631), .ZN(n6633) );
  OAI211_X1 U8372 ( .C1(n6726), .C2(n7364), .A(n6634), .B(n6633), .ZN(P1_U3216) );
  INV_X1 U8373 ( .A(n6635), .ZN(n6636) );
  AOI21_X1 U8374 ( .B1(n6638), .B2(n6637), .A(n6636), .ZN(n6931) );
  INV_X1 U8375 ( .A(n9992), .ZN(n9947) );
  AOI22_X1 U8376 ( .A1(n9328), .A2(n5499), .B1(n9985), .B2(n6423), .ZN(n6640)
         );
  OAI21_X1 U8377 ( .B1(n6839), .B2(n9932), .A(n6494), .ZN(n6639) );
  NAND3_X1 U8378 ( .A1(n6639), .A2(n9847), .A3(n6716), .ZN(n6924) );
  OAI211_X1 U8379 ( .C1(n6931), .C2(n9947), .A(n6640), .B(n6924), .ZN(n6642)
         );
  XNOR2_X1 U8380 ( .A(n8549), .B(n8433), .ZN(n6641) );
  INV_X1 U8381 ( .A(n9693), .ZN(n9972) );
  NOR2_X1 U8382 ( .A1(n6641), .A2(n9972), .ZN(n6928) );
  NOR2_X1 U8383 ( .A1(n6642), .A2(n6928), .ZN(n6646) );
  AOI22_X1 U8384 ( .A1(n5490), .A2(n6494), .B1(n10005), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n6643) );
  OAI21_X1 U8385 ( .B1(n6646), .B2(n10005), .A(n6643), .ZN(P1_U3525) );
  OAI22_X1 U8386 ( .A1(n9767), .A2(n6925), .B1(n9995), .B2(n4900), .ZN(n6644)
         );
  INV_X1 U8387 ( .A(n6644), .ZN(n6645) );
  OAI21_X1 U8388 ( .B1(n6646), .B2(n9994), .A(n6645), .ZN(P1_U3460) );
  NAND2_X1 U8389 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3084), .ZN(n7687) );
  OR2_X1 U8390 ( .A1(n6655), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6648) );
  NAND2_X1 U8391 ( .A1(n6648), .A2(n6647), .ZN(n6651) );
  OR2_X1 U8392 ( .A1(n7073), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7067) );
  NAND2_X1 U8393 ( .A1(n7073), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6649) );
  AND2_X1 U8394 ( .A1(n7067), .A2(n6649), .ZN(n6650) );
  NAND2_X1 U8395 ( .A1(n6650), .A2(n6651), .ZN(n7066) );
  OAI21_X1 U8396 ( .B1(n6651), .B2(n6650), .A(n7066), .ZN(n6652) );
  NAND2_X1 U8397 ( .A1(n9920), .A2(n6652), .ZN(n6653) );
  OAI211_X1 U8398 ( .C1(n9914), .C2(n4420), .A(n7687), .B(n6653), .ZN(n6660)
         );
  NAND2_X1 U8399 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7073), .ZN(n6656) );
  OAI21_X1 U8400 ( .B1(n7073), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6656), .ZN(
        n6657) );
  AOI211_X1 U8401 ( .C1(n6658), .C2(n6657), .A(n7072), .B(n9895), .ZN(n6659)
         );
  AOI211_X1 U8402 ( .C1(P1_ADDR_REG_13__SCAN_IN), .C2(n9882), .A(n6660), .B(
        n6659), .ZN(n6661) );
  INV_X1 U8403 ( .A(n6661), .ZN(P1_U3254) );
  NAND2_X1 U8404 ( .A1(n8828), .A2(n10055), .ZN(n6662) );
  NAND2_X1 U8405 ( .A1(n6663), .A2(n6662), .ZN(n6666) );
  INV_X1 U8406 ( .A(n6666), .ZN(n6672) );
  OR2_X1 U8407 ( .A1(n10008), .A2(n6672), .ZN(n6697) );
  XNOR2_X1 U8408 ( .A(n7013), .B(n8606), .ZN(n6675) );
  NAND2_X1 U8409 ( .A1(n8827), .A2(n10055), .ZN(n6676) );
  XNOR2_X1 U8410 ( .A(n6675), .B(n6676), .ZN(n6700) );
  OR2_X1 U8411 ( .A1(n6697), .A2(n6700), .ZN(n6682) );
  INV_X1 U8412 ( .A(n6662), .ZN(n6665) );
  NAND2_X1 U8413 ( .A1(n6665), .A2(n6664), .ZN(n6667) );
  INV_X1 U8414 ( .A(n6668), .ZN(n6671) );
  INV_X1 U8415 ( .A(n6669), .ZN(n6670) );
  INV_X1 U8416 ( .A(n6699), .ZN(n6674) );
  INV_X1 U8417 ( .A(n6700), .ZN(n6673) );
  NAND2_X1 U8418 ( .A1(n6674), .A2(n6673), .ZN(n6680) );
  INV_X1 U8419 ( .A(n6675), .ZN(n6678) );
  INV_X1 U8420 ( .A(n6676), .ZN(n6677) );
  NAND2_X1 U8421 ( .A1(n6678), .A2(n6677), .ZN(n6679) );
  AND2_X1 U8422 ( .A1(n6680), .A2(n6679), .ZN(n6681) );
  XNOR2_X1 U8423 ( .A(n6684), .B(n8631), .ZN(n6804) );
  NAND2_X1 U8424 ( .A1(n8826), .A2(n10055), .ZN(n6802) );
  XNOR2_X1 U8425 ( .A(n6804), .B(n6802), .ZN(n6805) );
  XNOR2_X1 U8426 ( .A(n6806), .B(n6805), .ZN(n6689) );
  NAND2_X1 U8427 ( .A1(n8809), .A2(n6684), .ZN(n6685) );
  OAI21_X1 U8428 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n8878), .A(n6685), .ZN(n6687) );
  OAI22_X1 U8429 ( .A1(n8805), .A2(n6985), .B1(n8781), .B2(n8254), .ZN(n6686)
         );
  AOI211_X1 U8430 ( .C1(n6991), .C2(n8784), .A(n6687), .B(n6686), .ZN(n6688)
         );
  OAI21_X1 U8431 ( .B1(n6689), .B2(n8812), .A(n6688), .ZN(P2_U3223) );
  INV_X1 U8432 ( .A(n6919), .ZN(n10080) );
  NAND2_X1 U8433 ( .A1(n6384), .A2(n10080), .ZN(n8090) );
  MUX2_X1 U8434 ( .A(n8090), .B(n10080), .S(n5952), .Z(n6690) );
  AOI21_X1 U8435 ( .B1(n6691), .B2(n6690), .A(n8812), .ZN(n6694) );
  INV_X1 U8436 ( .A(n8809), .ZN(n10020) );
  OAI22_X1 U8437 ( .A1(n10020), .A2(n10080), .B1(n8781), .B2(n6692), .ZN(n6693) );
  AOI211_X1 U8438 ( .C1(P2_REG3_REG_0__SCAN_IN), .C2(n6695), .A(n6694), .B(
        n6693), .ZN(n6696) );
  INV_X1 U8439 ( .A(n6696), .ZN(P2_U3234) );
  OR2_X1 U8440 ( .A1(n10009), .A2(n6697), .ZN(n6698) );
  AND2_X1 U8441 ( .A1(n6699), .A2(n6698), .ZN(n6701) );
  XNOR2_X1 U8442 ( .A(n6701), .B(n6700), .ZN(n6706) );
  AOI22_X1 U8443 ( .A1(n7206), .A2(n8828), .B1(n8808), .B2(n8826), .ZN(n6705)
         );
  NOR2_X1 U8444 ( .A1(n10020), .A2(n4503), .ZN(n6702) );
  AOI211_X1 U8445 ( .C1(n8784), .C2(n7012), .A(n6703), .B(n6702), .ZN(n6704)
         );
  OAI211_X1 U8446 ( .C1(n6706), .C2(n8812), .A(n6705), .B(n6704), .ZN(P2_U3215) );
  XNOR2_X1 U8447 ( .A(n6708), .B(n6707), .ZN(n6713) );
  OAI22_X1 U8448 ( .A1(n10020), .A2(n10094), .B1(n8781), .B2(n6709), .ZN(n6710) );
  AOI21_X1 U8449 ( .B1(n7206), .B2(n6385), .A(n6710), .ZN(n6712) );
  MUX2_X1 U8450 ( .A(n10026), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n6711) );
  OAI211_X1 U8451 ( .C1(n8812), .C2(n6713), .A(n6712), .B(n6711), .ZN(P2_U3220) );
  NAND2_X1 U8452 ( .A1(n6716), .A2(n7124), .ZN(n6717) );
  NAND2_X1 U8453 ( .A1(n6717), .A2(n9847), .ZN(n6718) );
  NOR2_X1 U8454 ( .A1(n6789), .A2(n6718), .ZN(n7122) );
  OAI22_X1 U8455 ( .A1(n8547), .A2(n9964), .B1(n6855), .B2(n9962), .ZN(n6719)
         );
  AOI211_X1 U8456 ( .C1(n7129), .C2(n9992), .A(n7122), .B(n6719), .ZN(n6722)
         );
  XNOR2_X1 U8457 ( .A(n6720), .B(n8430), .ZN(n6721) );
  NAND2_X1 U8458 ( .A1(n6721), .A2(n9693), .ZN(n7131) );
  NAND2_X1 U8459 ( .A1(n6722), .A2(n7131), .ZN(n6728) );
  OAI22_X1 U8460 ( .A1(n9767), .A2(n6726), .B1(n9995), .B2(n4915), .ZN(n6723)
         );
  AOI21_X1 U8461 ( .B1(n6728), .B2(n9995), .A(n6723), .ZN(n6724) );
  INV_X1 U8462 ( .A(n6724), .ZN(P1_U3463) );
  INV_X1 U8463 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6725) );
  OAI22_X1 U8464 ( .A1(n9728), .A2(n6726), .B1(n10007), .B2(n6725), .ZN(n6727)
         );
  AOI21_X1 U8465 ( .B1(n6728), .B2(n10007), .A(n6727), .ZN(n6729) );
  INV_X1 U8466 ( .A(n6729), .ZN(P1_U3526) );
  INV_X1 U8467 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6739) );
  XNOR2_X1 U8468 ( .A(n6730), .B(n6731), .ZN(n6850) );
  INV_X1 U8469 ( .A(n6731), .ZN(n8210) );
  XNOR2_X1 U8470 ( .A(n6732), .B(n8210), .ZN(n6733) );
  AOI222_X1 U8471 ( .A1(n10049), .A2(n6733), .B1(n8828), .B2(n10046), .C1(
        n10047), .C2(n10045), .ZN(n6842) );
  INV_X1 U8472 ( .A(n6734), .ZN(n6963) );
  INV_X1 U8473 ( .A(n6735), .ZN(n6900) );
  AOI211_X1 U8474 ( .C1(n6736), .C2(n6963), .A(n10055), .B(n6900), .ZN(n6847)
         );
  AOI21_X1 U8475 ( .B1(n10142), .B2(n6736), .A(n6847), .ZN(n6737) );
  OAI211_X1 U8476 ( .C1(n10146), .C2(n6850), .A(n6842), .B(n6737), .ZN(n6740)
         );
  NAND2_X1 U8477 ( .A1(n6740), .A2(n10158), .ZN(n6738) );
  OAI21_X1 U8478 ( .B1(n10158), .B2(n6739), .A(n6738), .ZN(P2_U3466) );
  INV_X1 U8479 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6742) );
  NAND2_X1 U8480 ( .A1(n6740), .A2(n10176), .ZN(n6741) );
  OAI21_X1 U8481 ( .B1(n10176), .B2(n6742), .A(n6741), .ZN(P2_U3525) );
  INV_X1 U8482 ( .A(n6743), .ZN(n6769) );
  AOI22_X1 U8483 ( .A1(n9367), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n6744), .ZN(n6745) );
  OAI21_X1 U8484 ( .B1(n6769), .B2(n9781), .A(n6745), .ZN(P1_U3336) );
  INV_X1 U8485 ( .A(n8895), .ZN(n7863) );
  INV_X1 U8486 ( .A(n6746), .ZN(n6766) );
  OAI222_X1 U8487 ( .A1(P2_U3152), .A2(n7863), .B1(n9221), .B2(n6766), .C1(
        n6747), .C2(n8019), .ZN(P2_U3342) );
  INV_X1 U8488 ( .A(n6748), .ZN(n6749) );
  NAND2_X1 U8489 ( .A1(n6750), .A2(n6749), .ZN(n6754) );
  AND2_X1 U8490 ( .A1(n6756), .A2(n6754), .ZN(n6759) );
  OR2_X1 U8491 ( .A1(n6855), .A2(n8719), .ZN(n6753) );
  NAND2_X1 U8492 ( .A1(n7098), .A2(n6884), .ZN(n6752) );
  NAND2_X1 U8493 ( .A1(n6753), .A2(n6752), .ZN(n6866) );
  XNOR2_X1 U8494 ( .A(n6865), .B(n6866), .ZN(n6758) );
  AND2_X1 U8495 ( .A1(n6758), .A2(n6754), .ZN(n6755) );
  OAI211_X1 U8496 ( .C1(n6759), .C2(n6758), .A(n6757), .B(n6869), .ZN(n6765)
         );
  INV_X1 U8497 ( .A(n7094), .ZN(n6763) );
  AOI21_X1 U8498 ( .B1(n9326), .B2(n9311), .A(n6760), .ZN(n6761) );
  OAI21_X1 U8499 ( .B1(n7095), .B2(n9272), .A(n6761), .ZN(n6762) );
  AOI21_X1 U8500 ( .B1(n9306), .B2(n6763), .A(n6762), .ZN(n6764) );
  OAI211_X1 U8501 ( .C1(n6798), .C2(n7364), .A(n6765), .B(n6764), .ZN(P1_U3228) );
  INV_X1 U8502 ( .A(n9355), .ZN(n7674) );
  OAI222_X1 U8503 ( .A1(n9771), .A2(n6767), .B1(n7674), .B2(P1_U3084), .C1(
        n9781), .C2(n6766), .ZN(P1_U3337) );
  INV_X1 U8504 ( .A(n7876), .ZN(n8270) );
  INV_X1 U8505 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6768) );
  OAI222_X1 U8506 ( .A1(P2_U3152), .A2(n8270), .B1(n9221), .B2(n6769), .C1(
        n6768), .C2(n8019), .ZN(P2_U3341) );
  NAND2_X1 U8507 ( .A1(n6777), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6771) );
  NAND2_X1 U8508 ( .A1(n6771), .A2(n6770), .ZN(n6774) );
  INV_X1 U8509 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6772) );
  AOI22_X1 U8510 ( .A1(n6937), .A2(n6772), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n6775), .ZN(n6773) );
  NOR2_X1 U8511 ( .A1(n6774), .A2(n6773), .ZN(n6932) );
  AOI21_X1 U8512 ( .B1(n6774), .B2(n6773), .A(n6932), .ZN(n6786) );
  INV_X1 U8513 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9821) );
  AOI22_X1 U8514 ( .A1(n6937), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n9821), .B2(
        n6775), .ZN(n6779) );
  OAI21_X1 U8515 ( .B1(n6779), .B2(n6778), .A(n6936), .ZN(n6780) );
  NAND2_X1 U8516 ( .A1(n6780), .A2(n10027), .ZN(n6785) );
  INV_X1 U8517 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n6782) );
  OAI22_X1 U8518 ( .A1(n8922), .A2(n6782), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6781), .ZN(n6783) );
  AOI21_X1 U8519 ( .B1(n8896), .B2(n6937), .A(n6783), .ZN(n6784) );
  OAI211_X1 U8520 ( .C1(n6786), .C2(n7886), .A(n6785), .B(n6784), .ZN(P2_U3258) );
  OAI21_X1 U8521 ( .B1(n6788), .B2(n6792), .A(n6787), .ZN(n7102) );
  OAI22_X1 U8522 ( .A1(n7095), .A2(n9964), .B1(n7293), .B2(n9962), .ZN(n6791)
         );
  INV_X1 U8523 ( .A(n6789), .ZN(n6790) );
  AOI211_X1 U8524 ( .C1(n7098), .C2(n6790), .A(n9622), .B(n6858), .ZN(n7093)
         );
  AOI211_X1 U8525 ( .C1(n7102), .C2(n9992), .A(n6791), .B(n7093), .ZN(n6794)
         );
  INV_X1 U8526 ( .A(n6792), .ZN(n8431) );
  XNOR2_X1 U8527 ( .A(n8300), .B(n8431), .ZN(n6793) );
  NAND2_X1 U8528 ( .A1(n6793), .A2(n9693), .ZN(n7104) );
  NAND2_X1 U8529 ( .A1(n6794), .A2(n7104), .ZN(n6800) );
  OAI22_X1 U8530 ( .A1(n9728), .A2(n6798), .B1(n10007), .B2(n6155), .ZN(n6795)
         );
  AOI21_X1 U8531 ( .B1(n6800), .B2(n10007), .A(n6795), .ZN(n6796) );
  INV_X1 U8532 ( .A(n6796), .ZN(P1_U3527) );
  INV_X1 U8533 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6797) );
  OAI22_X1 U8534 ( .A1(n9767), .A2(n6798), .B1(n9995), .B2(n6797), .ZN(n6799)
         );
  AOI21_X1 U8535 ( .B1(n6800), .B2(n9995), .A(n6799), .ZN(n6801) );
  INV_X1 U8536 ( .A(n6801), .ZN(P1_U3466) );
  INV_X1 U8537 ( .A(n6802), .ZN(n6803) );
  XNOR2_X1 U8538 ( .A(n6807), .B(n8606), .ZN(n6808) );
  NAND2_X1 U8539 ( .A1(n8825), .A2(n10055), .ZN(n6809) );
  NAND2_X1 U8540 ( .A1(n6808), .A2(n6809), .ZN(n7023) );
  INV_X1 U8541 ( .A(n6808), .ZN(n6811) );
  INV_X1 U8542 ( .A(n6809), .ZN(n6810) );
  NAND2_X1 U8543 ( .A1(n6811), .A2(n6810), .ZN(n6812) );
  AND2_X1 U8544 ( .A1(n7023), .A2(n6812), .ZN(n6813) );
  OAI21_X1 U8545 ( .B1(n6814), .B2(n6813), .A(n7024), .ZN(n6820) );
  NAND2_X1 U8546 ( .A1(n8826), .A2(n10045), .ZN(n6816) );
  NAND2_X1 U8547 ( .A1(n8824), .A2(n10046), .ZN(n6815) );
  NAND2_X1 U8548 ( .A1(n6816), .A2(n6815), .ZN(n7134) );
  AOI22_X1 U8549 ( .A1(n10018), .A2(n7134), .B1(P2_REG3_REG_9__SCAN_IN), .B2(
        P2_U3152), .ZN(n6818) );
  NAND2_X1 U8550 ( .A1(n8784), .A2(n7139), .ZN(n6817) );
  OAI211_X1 U8551 ( .C1(n10125), .C2(n10020), .A(n6818), .B(n6817), .ZN(n6819)
         );
  AOI21_X1 U8552 ( .B1(n6820), .B2(n10022), .A(n6819), .ZN(n6821) );
  INV_X1 U8553 ( .A(n6821), .ZN(P2_U3233) );
  AND2_X1 U8554 ( .A1(n6823), .A2(n6822), .ZN(n6824) );
  NAND2_X1 U8555 ( .A1(n6825), .A2(n6824), .ZN(n6922) );
  NAND2_X1 U8556 ( .A1(n9925), .A2(n8721), .ZN(n6826) );
  OAI21_X1 U8557 ( .B1(n6827), .B2(n6829), .A(n6828), .ZN(n9941) );
  XNOR2_X1 U8558 ( .A(n6830), .B(n6827), .ZN(n6831) );
  NAND2_X1 U8559 ( .A1(n6831), .A2(n9693), .ZN(n6833) );
  AOI22_X1 U8560 ( .A1(n9985), .A2(n9331), .B1(n9329), .B2(n5499), .ZN(n6832)
         );
  NAND2_X1 U8561 ( .A1(n6833), .A2(n6832), .ZN(n9944) );
  XNOR2_X1 U8562 ( .A(n9943), .B(n9932), .ZN(n6834) );
  NAND2_X1 U8563 ( .A1(n6834), .A2(n9847), .ZN(n9942) );
  OAI22_X1 U8564 ( .A1(n9942), .A2(n9513), .B1(n9598), .B2(n6835), .ZN(n6836)
         );
  INV_X1 U8565 ( .A(n9939), .ZN(n9620) );
  OAI21_X1 U8566 ( .B1(n9944), .B2(n6836), .A(n9620), .ZN(n6841) );
  NAND2_X1 U8567 ( .A1(n9931), .A2(n6837), .ZN(n6838) );
  AOI22_X1 U8568 ( .A1(n9844), .A2(n6839), .B1(n9939), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6840) );
  OAI211_X1 U8569 ( .C1(n9589), .C2(n9941), .A(n6841), .B(n6840), .ZN(P1_U3290) );
  MUX2_X1 U8570 ( .A(n6286), .B(n6842), .S(n9049), .Z(n6849) );
  INV_X1 U8571 ( .A(n10065), .ZN(n9124) );
  INV_X1 U8572 ( .A(n6843), .ZN(n6844) );
  OAI22_X1 U8573 ( .A1(n10054), .A2(n6845), .B1(n8975), .B2(n6844), .ZN(n6846)
         );
  AOI21_X1 U8574 ( .B1(n6847), .B2(n9124), .A(n6846), .ZN(n6848) );
  OAI211_X1 U8575 ( .C1(n6850), .C2(n9126), .A(n6849), .B(n6848), .ZN(P2_U3291) );
  NAND2_X1 U8576 ( .A1(n9330), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6851) );
  OAI21_X1 U8577 ( .B1(n9228), .B2(n9330), .A(n6851), .ZN(P1_U3583) );
  XNOR2_X1 U8578 ( .A(n6852), .B(n8429), .ZN(n9948) );
  NAND2_X1 U8579 ( .A1(n8301), .A2(n8298), .ZN(n6853) );
  NAND2_X1 U8580 ( .A1(n6853), .A2(n8429), .ZN(n7290) );
  OAI21_X1 U8581 ( .B1(n8429), .B2(n6853), .A(n7290), .ZN(n6854) );
  NAND2_X1 U8582 ( .A1(n6854), .A2(n9693), .ZN(n6857) );
  OR2_X1 U8583 ( .A1(n6855), .A2(n9964), .ZN(n6856) );
  NAND2_X1 U8584 ( .A1(n6857), .A2(n6856), .ZN(n9952) );
  OR2_X1 U8585 ( .A1(n6858), .A2(n9949), .ZN(n6859) );
  AND3_X1 U8586 ( .A1(n7283), .A2(n6859), .A3(n9847), .ZN(n9951) );
  INV_X1 U8587 ( .A(n9951), .ZN(n6860) );
  OAI22_X1 U8588 ( .A1(n6860), .A2(n9513), .B1(n9598), .B2(n7005), .ZN(n6861)
         );
  INV_X1 U8589 ( .A(n9939), .ZN(n9601) );
  OAI21_X1 U8590 ( .B1(n9952), .B2(n6861), .A(n9601), .ZN(n6864) );
  OR2_X1 U8591 ( .A1(n9939), .A2(n9962), .ZN(n9527) );
  INV_X1 U8592 ( .A(n9527), .ZN(n9605) );
  OAI22_X1 U8593 ( .A1(n9949), .A2(n9628), .B1(n9601), .B2(n6201), .ZN(n6862)
         );
  AOI21_X1 U8594 ( .B1(n9605), .B2(n9325), .A(n6862), .ZN(n6863) );
  OAI211_X1 U8595 ( .C1(n9948), .C2(n9589), .A(n6864), .B(n6863), .ZN(P1_U3286) );
  INV_X1 U8596 ( .A(n6865), .ZN(n6867) );
  NAND2_X1 U8597 ( .A1(n6867), .A2(n6866), .ZN(n6868) );
  OAI22_X1 U8598 ( .A1(n7293), .A2(n6498), .B1(n9949), .B2(n8718), .ZN(n6870)
         );
  XNOR2_X1 U8599 ( .A(n6870), .B(n8721), .ZN(n6873) );
  OR2_X1 U8600 ( .A1(n7293), .A2(n8719), .ZN(n6872) );
  NAND2_X1 U8601 ( .A1(n7007), .A2(n6884), .ZN(n6871) );
  NAND2_X1 U8602 ( .A1(n6872), .A2(n6871), .ZN(n7001) );
  INV_X1 U8603 ( .A(n6873), .ZN(n6998) );
  INV_X1 U8604 ( .A(n7001), .ZN(n6874) );
  NAND2_X1 U8605 ( .A1(n6998), .A2(n6874), .ZN(n6878) );
  OAI22_X1 U8606 ( .A1(n9965), .A2(n6498), .B1(n9958), .B2(n8718), .ZN(n6875)
         );
  XNOR2_X1 U8607 ( .A(n6875), .B(n8689), .ZN(n6879) );
  OR2_X1 U8608 ( .A1(n9965), .A2(n8719), .ZN(n6877) );
  NAND2_X1 U8609 ( .A1(n7288), .A2(n6884), .ZN(n6876) );
  AND2_X1 U8610 ( .A1(n6877), .A2(n6876), .ZN(n6880) );
  NAND2_X1 U8611 ( .A1(n6879), .A2(n6880), .ZN(n7145) );
  INV_X1 U8612 ( .A(n6879), .ZN(n6882) );
  INV_X1 U8613 ( .A(n6880), .ZN(n6881) );
  NAND2_X1 U8614 ( .A1(n6882), .A2(n6881), .ZN(n7146) );
  NAND2_X1 U8615 ( .A1(n6883), .A2(n7146), .ZN(n7080) );
  OR2_X1 U8616 ( .A1(n7292), .A2(n8719), .ZN(n6886) );
  NAND2_X1 U8617 ( .A1(n9968), .A2(n6884), .ZN(n6885) );
  NAND2_X1 U8618 ( .A1(n6886), .A2(n6885), .ZN(n7079) );
  NAND2_X1 U8619 ( .A1(n9968), .A2(n8714), .ZN(n6887) );
  OAI21_X1 U8620 ( .B1(n7292), .B2(n6498), .A(n6887), .ZN(n6888) );
  XNOR2_X1 U8621 ( .A(n6888), .B(n8721), .ZN(n7078) );
  XOR2_X1 U8622 ( .A(n7079), .B(n7078), .Z(n6889) );
  XNOR2_X1 U8623 ( .A(n7080), .B(n6889), .ZN(n6895) );
  OAI21_X1 U8624 ( .B1(n9963), .B2(n9304), .A(n6890), .ZN(n6891) );
  AOI21_X1 U8625 ( .B1(n9310), .B2(n9325), .A(n6891), .ZN(n6892) );
  OAI21_X1 U8626 ( .B1(n9262), .B2(n7109), .A(n6892), .ZN(n6893) );
  AOI21_X1 U8627 ( .B1(n9320), .B2(n9968), .A(n6893), .ZN(n6894) );
  OAI21_X1 U8628 ( .B1(n6895), .B2(n9315), .A(n6894), .ZN(P1_U3211) );
  XNOR2_X1 U8629 ( .A(n6896), .B(n8212), .ZN(n10104) );
  INV_X1 U8630 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6899) );
  XNOR2_X1 U8631 ( .A(n6897), .B(n8212), .ZN(n6898) );
  INV_X1 U8632 ( .A(n10045), .ZN(n9074) );
  OAI22_X1 U8633 ( .A1(n6962), .A2(n9074), .B1(n6985), .B2(n9076), .ZN(n10017)
         );
  AOI21_X1 U8634 ( .B1(n6898), .B2(n10049), .A(n10017), .ZN(n10107) );
  MUX2_X1 U8635 ( .A(n6899), .B(n10107), .S(n9049), .Z(n6904) );
  INV_X1 U8636 ( .A(n9088), .ZN(n8935) );
  INV_X1 U8637 ( .A(n6902), .ZN(n10105) );
  OAI21_X1 U8638 ( .B1(n6900), .B2(n10105), .A(n7011), .ZN(n10106) );
  OAI22_X1 U8639 ( .A1(n8935), .A2(n10106), .B1(n10025), .B2(n8975), .ZN(n6901) );
  AOI21_X1 U8640 ( .B1(n8926), .B2(n6902), .A(n6901), .ZN(n6903) );
  OAI211_X1 U8641 ( .C1(n10104), .C2(n9126), .A(n6904), .B(n6903), .ZN(
        P2_U3290) );
  NOR2_X1 U8642 ( .A1(n9049), .A2(n6905), .ZN(n6908) );
  INV_X1 U8643 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7431) );
  OAI22_X1 U8644 ( .A1(n10065), .A2(n6906), .B1(n7431), .B2(n8975), .ZN(n6907)
         );
  AOI211_X1 U8645 ( .C1(n9049), .C2(n6909), .A(n6908), .B(n6907), .ZN(n6913)
         );
  INV_X1 U8646 ( .A(n9126), .ZN(n9082) );
  AOI22_X1 U8647 ( .A1(n9082), .A2(n6911), .B1(n8926), .B2(n6910), .ZN(n6912)
         );
  NAND2_X1 U8648 ( .A1(n6913), .A2(n6912), .ZN(P2_U3295) );
  NAND2_X1 U8649 ( .A1(n6914), .A2(n10080), .ZN(n6915) );
  NAND2_X1 U8650 ( .A1(n6916), .A2(n6915), .ZN(n10082) );
  INV_X1 U8651 ( .A(n10082), .ZN(n6917) );
  AOI22_X1 U8652 ( .A1(n6917), .A2(n10049), .B1(n10046), .B2(n6463), .ZN(
        n10079) );
  INV_X1 U8653 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7568) );
  OAI22_X1 U8654 ( .A1(n10070), .A2(n10079), .B1(n7568), .B2(n8975), .ZN(n6918) );
  AOI21_X1 U8655 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n10070), .A(n6918), .ZN(
        n6921) );
  OAI21_X1 U8656 ( .B1(n9088), .B2(n8926), .A(n6919), .ZN(n6920) );
  OAI211_X1 U8657 ( .C1(n9126), .C2(n10082), .A(n6921), .B(n6920), .ZN(
        P2_U3296) );
  OR2_X1 U8658 ( .A1(n9939), .A2(n9964), .ZN(n9597) );
  INV_X1 U8659 ( .A(n9597), .ZN(n9525) );
  OR2_X1 U8660 ( .A1(n6922), .A2(n9513), .ZN(n9530) );
  INV_X1 U8661 ( .A(n9598), .ZN(n9936) );
  AOI22_X1 U8662 ( .A1(n9939), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9936), .ZN(n6923) );
  OAI21_X1 U8663 ( .B1(n9530), .B2(n6924), .A(n6923), .ZN(n6927) );
  OAI22_X1 U8664 ( .A1(n7095), .A2(n9527), .B1(n9628), .B2(n6925), .ZN(n6926)
         );
  AOI211_X1 U8665 ( .C1(n9525), .C2(n6423), .A(n6927), .B(n6926), .ZN(n6930)
         );
  NAND2_X1 U8666 ( .A1(n6928), .A2(n9601), .ZN(n6929) );
  OAI211_X1 U8667 ( .C1(n6931), .C2(n9589), .A(n6930), .B(n6929), .ZN(P1_U3289) );
  NOR2_X1 U8668 ( .A1(n6937), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6933) );
  NOR2_X1 U8669 ( .A1(n6933), .A2(n6932), .ZN(n6935) );
  INV_X1 U8670 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7270) );
  AOI22_X1 U8671 ( .A1(n7267), .A2(n7270), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7271), .ZN(n6934) );
  NOR2_X1 U8672 ( .A1(n6935), .A2(n6934), .ZN(n7269) );
  AOI21_X1 U8673 ( .B1(n6935), .B2(n6934), .A(n7269), .ZN(n6945) );
  INV_X1 U8674 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9813) );
  AOI22_X1 U8675 ( .A1(n7267), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n9813), .B2(
        n7271), .ZN(n6939) );
  OAI21_X1 U8676 ( .B1(n6939), .B2(n6938), .A(n7266), .ZN(n6940) );
  NAND2_X1 U8677 ( .A1(n6940), .A2(n10027), .ZN(n6944) );
  INV_X1 U8678 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6941) );
  NAND2_X1 U8679 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7207) );
  OAI21_X1 U8680 ( .B1(n8922), .B2(n6941), .A(n7207), .ZN(n6942) );
  AOI21_X1 U8681 ( .B1(n8896), .B2(n7267), .A(n6942), .ZN(n6943) );
  OAI211_X1 U8682 ( .C1(n6945), .C2(n7886), .A(n6944), .B(n6943), .ZN(P2_U3259) );
  OAI21_X1 U8683 ( .B1(n6946), .B2(n10086), .A(n10057), .ZN(n10087) );
  OAI21_X1 U8684 ( .B1(n6947), .B2(n8207), .A(n6948), .ZN(n10090) );
  AOI22_X1 U8685 ( .A1(n9082), .A2(n10090), .B1(n8926), .B2(n6949), .ZN(n6958)
         );
  NAND2_X1 U8686 ( .A1(n6951), .A2(n8207), .ZN(n6952) );
  NAND2_X1 U8687 ( .A1(n6950), .A2(n6952), .ZN(n6953) );
  NAND2_X1 U8688 ( .A1(n6953), .A2(n10049), .ZN(n6955) );
  AOI22_X1 U8689 ( .A1(n10045), .A2(n6463), .B1(n5620), .B2(n10046), .ZN(n6954) );
  NAND2_X1 U8690 ( .A1(n6955), .A2(n6954), .ZN(n10088) );
  OAI22_X1 U8691 ( .A1(n8975), .A2(n7490), .B1(n6280), .B2(n9049), .ZN(n6956)
         );
  AOI21_X1 U8692 ( .B1(n9049), .B2(n10088), .A(n6956), .ZN(n6957) );
  OAI211_X1 U8693 ( .C1(n8935), .C2(n10087), .A(n6958), .B(n6957), .ZN(
        P2_U3294) );
  XNOR2_X1 U8694 ( .A(n6959), .B(n8208), .ZN(n6960) );
  OAI222_X1 U8695 ( .A1(n9076), .A2(n6962), .B1(n9074), .B2(n6961), .C1(n6960), 
        .C2(n9071), .ZN(n10100) );
  INV_X1 U8696 ( .A(n10100), .ZN(n6973) );
  INV_X1 U8697 ( .A(n10058), .ZN(n6964) );
  OAI21_X1 U8698 ( .B1(n10098), .B2(n6964), .A(n6963), .ZN(n10099) );
  INV_X1 U8699 ( .A(n10099), .ZN(n6967) );
  OAI22_X1 U8700 ( .A1(n8975), .A2(n6965), .B1(n6285), .B2(n9049), .ZN(n6966)
         );
  AOI21_X1 U8701 ( .B1(n9088), .B2(n6967), .A(n6966), .ZN(n6972) );
  OAI21_X1 U8702 ( .B1(n6969), .B2(n8208), .A(n6968), .ZN(n10102) );
  AOI22_X1 U8703 ( .A1(n9082), .A2(n10102), .B1(n8926), .B2(n6970), .ZN(n6971)
         );
  OAI211_X1 U8704 ( .C1(n6973), .C2(n10070), .A(n6972), .B(n6971), .ZN(
        P2_U3292) );
  INV_X1 U8705 ( .A(n6974), .ZN(n6976) );
  OAI222_X1 U8706 ( .A1(n8019), .A2(n6975), .B1(n9221), .B2(n6976), .C1(
        P2_U3152), .C2(n7882), .ZN(P2_U3340) );
  INV_X1 U8707 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6977) );
  INV_X1 U8708 ( .A(n9368), .ZN(n9915) );
  OAI222_X1 U8709 ( .A1(n9777), .A2(n6977), .B1(n7846), .B2(n6976), .C1(
        P1_U3084), .C2(n9915), .ZN(P1_U3335) );
  NAND2_X1 U8710 ( .A1(n6978), .A2(n8215), .ZN(n6979) );
  NAND2_X1 U8711 ( .A1(n6980), .A2(n6979), .ZN(n10117) );
  INV_X1 U8712 ( .A(n6981), .ZN(n6982) );
  NAND2_X1 U8713 ( .A1(n9049), .A2(n6982), .ZN(n10053) );
  OAI21_X1 U8714 ( .B1(n8215), .B2(n6984), .A(n6983), .ZN(n6987) );
  OAI22_X1 U8715 ( .A1(n6985), .A2(n9074), .B1(n8254), .B2(n9076), .ZN(n6986)
         );
  AOI21_X1 U8716 ( .B1(n6987), .B2(n10049), .A(n6986), .ZN(n6988) );
  OAI21_X1 U8717 ( .B1(n10039), .B2(n10117), .A(n6988), .ZN(n10120) );
  NAND2_X1 U8718 ( .A1(n10120), .A2(n9049), .ZN(n6996) );
  NOR2_X1 U8719 ( .A1(n6989), .A2(n10118), .ZN(n6990) );
  OR2_X1 U8720 ( .A1(n7137), .A2(n6990), .ZN(n10119) );
  INV_X1 U8721 ( .A(n10119), .ZN(n6994) );
  AOI22_X1 U8722 ( .A1(n10070), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n6991), .B2(
        n10062), .ZN(n6992) );
  OAI21_X1 U8723 ( .B1(n10118), .B2(n10054), .A(n6992), .ZN(n6993) );
  AOI21_X1 U8724 ( .B1(n9088), .B2(n6994), .A(n6993), .ZN(n6995) );
  OAI211_X1 U8725 ( .C1(n10117), .C2(n10053), .A(n6996), .B(n6995), .ZN(
        P2_U3288) );
  INV_X1 U8726 ( .A(n6997), .ZN(n6999) );
  NAND2_X1 U8727 ( .A1(n6999), .A2(n6998), .ZN(n7147) );
  OAI21_X1 U8728 ( .B1(n6999), .B2(n6998), .A(n7147), .ZN(n7000) );
  NOR2_X1 U8729 ( .A1(n7000), .A2(n7001), .ZN(n7149) );
  AOI21_X1 U8730 ( .B1(n7001), .B2(n7000), .A(n7149), .ZN(n7009) );
  NOR2_X1 U8731 ( .A1(n9965), .A2(n9304), .ZN(n7002) );
  AOI211_X1 U8732 ( .C1(n9302), .C2(n9327), .A(n7003), .B(n7002), .ZN(n7004)
         );
  OAI21_X1 U8733 ( .B1(n9262), .B2(n7005), .A(n7004), .ZN(n7006) );
  AOI21_X1 U8734 ( .B1(n9320), .B2(n7007), .A(n7006), .ZN(n7008) );
  OAI21_X1 U8735 ( .B1(n7009), .B2(n9315), .A(n7008), .ZN(P1_U3225) );
  XNOR2_X1 U8736 ( .A(n7010), .B(n8211), .ZN(n10115) );
  XNOR2_X1 U8737 ( .A(n7011), .B(n7013), .ZN(n10112) );
  AOI22_X1 U8738 ( .A1(n8926), .A2(n7013), .B1(n10062), .B2(n7012), .ZN(n7014)
         );
  OAI21_X1 U8739 ( .B1(n8935), .B2(n10112), .A(n7014), .ZN(n7021) );
  NAND2_X1 U8740 ( .A1(n7016), .A2(n8211), .ZN(n7017) );
  NAND3_X1 U8741 ( .A1(n4597), .A2(n10049), .A3(n7017), .ZN(n7019) );
  AOI22_X1 U8742 ( .A1(n10045), .A2(n8828), .B1(n8826), .B2(n10046), .ZN(n7018) );
  NAND2_X1 U8743 ( .A1(n7019), .A2(n7018), .ZN(n10113) );
  MUX2_X1 U8744 ( .A(n10113), .B(P2_REG2_REG_7__SCAN_IN), .S(n10070), .Z(n7020) );
  AOI211_X1 U8745 ( .C1(n9082), .C2(n10115), .A(n7021), .B(n7020), .ZN(n7022)
         );
  INV_X1 U8746 ( .A(n7022), .ZN(P2_U3289) );
  INV_X1 U8747 ( .A(n8788), .ZN(n7026) );
  XNOR2_X1 U8748 ( .A(n10132), .B(n8606), .ZN(n7032) );
  NAND2_X1 U8749 ( .A1(n8824), .A2(n10055), .ZN(n7033) );
  XNOR2_X1 U8750 ( .A(n7032), .B(n7033), .ZN(n8787) );
  XNOR2_X1 U8751 ( .A(n10141), .B(n8631), .ZN(n7039) );
  INV_X1 U8752 ( .A(n5952), .ZN(n8630) );
  NAND2_X1 U8753 ( .A1(n8823), .A2(n8630), .ZN(n7037) );
  XNOR2_X1 U8754 ( .A(n7039), .B(n7037), .ZN(n8792) );
  INV_X1 U8755 ( .A(n8792), .ZN(n7036) );
  NAND2_X1 U8756 ( .A1(n7026), .A2(n4348), .ZN(n7052) );
  XNOR2_X1 U8757 ( .A(n7330), .B(n8606), .ZN(n7027) );
  NAND2_X1 U8758 ( .A1(n8822), .A2(n8630), .ZN(n7028) );
  NAND2_X1 U8759 ( .A1(n7027), .A2(n7028), .ZN(n7044) );
  INV_X1 U8760 ( .A(n7027), .ZN(n7030) );
  INV_X1 U8761 ( .A(n7028), .ZN(n7029) );
  NAND2_X1 U8762 ( .A1(n7030), .A2(n7029), .ZN(n7031) );
  NAND2_X1 U8763 ( .A1(n7044), .A2(n7031), .ZN(n7055) );
  INV_X1 U8764 ( .A(n7055), .ZN(n7042) );
  INV_X1 U8765 ( .A(n7032), .ZN(n7035) );
  INV_X1 U8766 ( .A(n7033), .ZN(n7034) );
  NAND2_X1 U8767 ( .A1(n7035), .A2(n7034), .ZN(n8789) );
  OR2_X1 U8768 ( .A1(n7036), .A2(n8789), .ZN(n7041) );
  INV_X1 U8769 ( .A(n7037), .ZN(n7038) );
  NAND2_X1 U8770 ( .A1(n7039), .A2(n7038), .ZN(n7040) );
  AND2_X1 U8771 ( .A1(n7041), .A2(n7040), .ZN(n7051) );
  AND2_X1 U8772 ( .A1(n7042), .A2(n7051), .ZN(n7043) );
  NAND2_X1 U8773 ( .A1(n7052), .A2(n7043), .ZN(n7053) );
  NAND2_X1 U8774 ( .A1(n7053), .A2(n7044), .ZN(n7203) );
  XNOR2_X1 U8775 ( .A(n7048), .B(n8606), .ZN(n7201) );
  NAND2_X1 U8776 ( .A1(n8821), .A2(n8630), .ZN(n7200) );
  XNOR2_X1 U8777 ( .A(n7201), .B(n7200), .ZN(n7202) );
  XNOR2_X1 U8778 ( .A(n7203), .B(n7202), .ZN(n7050) );
  OAI22_X1 U8779 ( .A1(n8781), .A2(n7891), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6781), .ZN(n7047) );
  INV_X1 U8780 ( .A(n7629), .ZN(n7045) );
  OAI22_X1 U8781 ( .A1(n8805), .A2(n7623), .B1(n7045), .B2(n10026), .ZN(n7046)
         );
  AOI211_X1 U8782 ( .C1(n7048), .C2(n8809), .A(n7047), .B(n7046), .ZN(n7049)
         );
  OAI21_X1 U8783 ( .B1(n7050), .B2(n8812), .A(n7049), .ZN(P2_U3236) );
  NAND2_X1 U8784 ( .A1(n7052), .A2(n7051), .ZN(n7056) );
  INV_X1 U8785 ( .A(n7053), .ZN(n7054) );
  AOI21_X1 U8786 ( .B1(n7056), .B2(n7055), .A(n7054), .ZN(n7063) );
  NAND2_X1 U8787 ( .A1(n8823), .A2(n10045), .ZN(n7058) );
  NAND2_X1 U8788 ( .A1(n8821), .A2(n10046), .ZN(n7057) );
  AND2_X1 U8789 ( .A1(n7058), .A2(n7057), .ZN(n7319) );
  OAI22_X1 U8790 ( .A1(n8637), .A2(n7319), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7059), .ZN(n7060) );
  AOI21_X1 U8791 ( .B1(n7329), .B2(n8784), .A(n7060), .ZN(n7062) );
  NAND2_X1 U8792 ( .A1(n7330), .A2(n8809), .ZN(n7061) );
  OAI211_X1 U8793 ( .C1(n7063), .C2(n8812), .A(n7062), .B(n7061), .ZN(P2_U3226) );
  NAND2_X1 U8794 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3084), .ZN(n7777) );
  OR2_X1 U8795 ( .A1(n7220), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7065) );
  NAND2_X1 U8796 ( .A1(n7220), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7064) );
  AND2_X1 U8797 ( .A1(n7065), .A2(n7064), .ZN(n7069) );
  NAND2_X1 U8798 ( .A1(n7067), .A2(n7066), .ZN(n7068) );
  NAND2_X1 U8799 ( .A1(n7069), .A2(n7068), .ZN(n7219) );
  OAI21_X1 U8800 ( .B1(n7069), .B2(n7068), .A(n7219), .ZN(n7070) );
  NAND2_X1 U8801 ( .A1(n9920), .A2(n7070), .ZN(n7071) );
  OAI211_X1 U8802 ( .C1(n9914), .C2(n7212), .A(n7777), .B(n7071), .ZN(n7076)
         );
  NOR2_X1 U8803 ( .A1(n7934), .A2(n7074), .ZN(n7214) );
  AOI211_X1 U8804 ( .C1(n7074), .C2(n7934), .A(n7214), .B(n9895), .ZN(n7075)
         );
  AOI211_X1 U8805 ( .C1(P1_ADDR_REG_14__SCAN_IN), .C2(n9882), .A(n7076), .B(
        n7075), .ZN(n7077) );
  INV_X1 U8806 ( .A(n7077), .ZN(P1_U3255) );
  NAND2_X1 U8807 ( .A1(n7177), .A2(n8716), .ZN(n7082) );
  OR2_X1 U8808 ( .A1(n9963), .A2(n8719), .ZN(n7081) );
  NAND2_X1 U8809 ( .A1(n7082), .A2(n7081), .ZN(n7239) );
  NAND2_X1 U8810 ( .A1(n7177), .A2(n8714), .ZN(n7084) );
  OR2_X1 U8811 ( .A1(n9963), .A2(n6498), .ZN(n7083) );
  NAND2_X1 U8812 ( .A1(n7084), .A2(n7083), .ZN(n7085) );
  XNOR2_X1 U8813 ( .A(n7085), .B(n8721), .ZN(n7238) );
  XOR2_X1 U8814 ( .A(n7239), .B(n7238), .Z(n7086) );
  XNOR2_X1 U8815 ( .A(n7240), .B(n7086), .ZN(n7092) );
  INV_X1 U8816 ( .A(n9306), .ZN(n9282) );
  NAND2_X1 U8817 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3084), .ZN(n9890) );
  OAI21_X1 U8818 ( .B1(n7087), .B2(n9304), .A(n9890), .ZN(n7088) );
  AOI21_X1 U8819 ( .B1(n9310), .B2(n9976), .A(n7088), .ZN(n7089) );
  OAI21_X1 U8820 ( .B1(n9282), .B2(n7173), .A(n7089), .ZN(n7090) );
  AOI21_X1 U8821 ( .B1(n9320), .B2(n7177), .A(n7090), .ZN(n7091) );
  OAI21_X1 U8822 ( .B1(n7092), .B2(n9315), .A(n7091), .ZN(P1_U3219) );
  INV_X1 U8823 ( .A(n7093), .ZN(n7100) );
  OAI22_X1 U8824 ( .A1(n9620), .A2(n6138), .B1(n7094), .B2(n9598), .ZN(n7097)
         );
  OAI22_X1 U8825 ( .A1(n7095), .A2(n9597), .B1(n9527), .B2(n7293), .ZN(n7096)
         );
  AOI211_X1 U8826 ( .C1(n9844), .C2(n7098), .A(n7097), .B(n7096), .ZN(n7099)
         );
  OAI21_X1 U8827 ( .B1(n7100), .B2(n9530), .A(n7099), .ZN(n7101) );
  AOI21_X1 U8828 ( .B1(n9595), .B2(n7102), .A(n7101), .ZN(n7103) );
  OAI21_X1 U8829 ( .B1(n9939), .B2(n7104), .A(n7103), .ZN(P1_U3287) );
  XOR2_X1 U8830 ( .A(n7105), .B(n7107), .Z(n9971) );
  NAND2_X1 U8831 ( .A1(n9620), .A2(n9693), .ZN(n9611) );
  OAI21_X1 U8832 ( .B1(n7108), .B2(n7107), .A(n7106), .ZN(n9974) );
  NAND2_X1 U8833 ( .A1(n9974), .A2(n9595), .ZN(n7117) );
  AOI211_X1 U8834 ( .C1(n9968), .C2(n7284), .A(n9622), .B(n4387), .ZN(n9966)
         );
  INV_X1 U8835 ( .A(n9530), .ZN(n9850) );
  NOR2_X1 U8836 ( .A1(n9597), .A2(n9965), .ZN(n7112) );
  OAI22_X1 U8837 ( .A1(n9620), .A2(n7110), .B1(n7109), .B2(n9598), .ZN(n7111)
         );
  AOI211_X1 U8838 ( .C1(n9605), .C2(n9984), .A(n7112), .B(n7111), .ZN(n7113)
         );
  OAI21_X1 U8839 ( .B1(n7114), .B2(n9628), .A(n7113), .ZN(n7115) );
  AOI21_X1 U8840 ( .B1(n9966), .B2(n9850), .A(n7115), .ZN(n7116) );
  OAI211_X1 U8841 ( .C1(n9971), .C2(n9611), .A(n7117), .B(n7116), .ZN(P1_U3284) );
  INV_X1 U8842 ( .A(n7118), .ZN(n7120) );
  OAI222_X1 U8843 ( .A1(n9777), .A2(n7119), .B1(n7846), .B2(n7120), .C1(n9408), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  OAI222_X1 U8844 ( .A1(n8019), .A2(n7121), .B1(n9221), .B2(n7120), .C1(
        P2_U3152), .C2(n4315), .ZN(P2_U3339) );
  INV_X1 U8845 ( .A(n7122), .ZN(n7127) );
  OAI22_X1 U8846 ( .A1(n9620), .A2(n6134), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9598), .ZN(n7123) );
  AOI21_X1 U8847 ( .B1(n9844), .B2(n7124), .A(n7123), .ZN(n7126) );
  AOI22_X1 U8848 ( .A1(n9605), .A2(n9327), .B1(n9525), .B2(n9329), .ZN(n7125)
         );
  OAI211_X1 U8849 ( .C1(n9530), .C2(n7127), .A(n7126), .B(n7125), .ZN(n7128)
         );
  AOI21_X1 U8850 ( .B1(n7129), .B2(n9595), .A(n7128), .ZN(n7130) );
  OAI21_X1 U8851 ( .B1(n9939), .B2(n7131), .A(n7130), .ZN(P1_U3288) );
  INV_X1 U8852 ( .A(n8216), .ZN(n8121) );
  XNOR2_X1 U8853 ( .A(n7132), .B(n8121), .ZN(n10124) );
  XNOR2_X1 U8854 ( .A(n7133), .B(n8216), .ZN(n7135) );
  AOI21_X1 U8855 ( .B1(n7135), .B2(n10049), .A(n7134), .ZN(n7136) );
  OAI21_X1 U8856 ( .B1(n10039), .B2(n10124), .A(n7136), .ZN(n10127) );
  NAND2_X1 U8857 ( .A1(n10127), .A2(n9049), .ZN(n7144) );
  OR2_X1 U8858 ( .A1(n7137), .A2(n10125), .ZN(n7138) );
  NAND2_X1 U8859 ( .A1(n7190), .A2(n7138), .ZN(n10126) );
  INV_X1 U8860 ( .A(n10126), .ZN(n7142) );
  AOI22_X1 U8861 ( .A1(n10070), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7139), .B2(
        n10062), .ZN(n7140) );
  OAI21_X1 U8862 ( .B1(n10125), .B2(n10054), .A(n7140), .ZN(n7141) );
  AOI21_X1 U8863 ( .B1(n7142), .B2(n9088), .A(n7141), .ZN(n7143) );
  OAI211_X1 U8864 ( .C1(n10124), .C2(n10053), .A(n7144), .B(n7143), .ZN(
        P2_U3287) );
  NAND2_X1 U8865 ( .A1(n7146), .A2(n7145), .ZN(n7151) );
  INV_X1 U8866 ( .A(n7147), .ZN(n7148) );
  NOR2_X1 U8867 ( .A1(n7149), .A2(n7148), .ZN(n7150) );
  XOR2_X1 U8868 ( .A(n7151), .B(n7150), .Z(n7158) );
  INV_X1 U8869 ( .A(n7152), .ZN(n7154) );
  NOR2_X1 U8870 ( .A1(n7292), .A2(n9304), .ZN(n7153) );
  AOI211_X1 U8871 ( .C1(n9310), .C2(n9326), .A(n7154), .B(n7153), .ZN(n7155)
         );
  OAI21_X1 U8872 ( .B1(n9282), .B2(n7286), .A(n7155), .ZN(n7156) );
  AOI21_X1 U8873 ( .B1(n9320), .B2(n7288), .A(n7156), .ZN(n7157) );
  OAI21_X1 U8874 ( .B1(n7158), .B2(n9315), .A(n7157), .ZN(P1_U3237) );
  INV_X1 U8875 ( .A(n7159), .ZN(n7162) );
  OAI222_X1 U8876 ( .A1(n9781), .A2(n7162), .B1(P1_U3084), .B2(n8583), .C1(
        n7160), .C2(n9777), .ZN(P1_U3333) );
  OAI222_X1 U8877 ( .A1(n8019), .A2(n7163), .B1(n9221), .B2(n7162), .C1(n7161), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  INV_X1 U8878 ( .A(n7164), .ZN(n7182) );
  OAI222_X1 U8879 ( .A1(n9781), .A2(n7182), .B1(P1_U3084), .B2(n8458), .C1(
        n7165), .C2(n9777), .ZN(P1_U3332) );
  INV_X1 U8880 ( .A(n7166), .ZN(n7167) );
  AOI21_X1 U8881 ( .B1(n8436), .B2(n7168), .A(n7167), .ZN(n9981) );
  INV_X1 U8882 ( .A(n9981), .ZN(n7181) );
  AOI21_X1 U8883 ( .B1(n7169), .B2(n5027), .A(n9972), .ZN(n7171) );
  AND2_X1 U8884 ( .A1(n7171), .A2(n7170), .ZN(n9980) );
  INV_X1 U8885 ( .A(n7305), .ZN(n7172) );
  OAI211_X1 U8886 ( .C1(n4623), .C2(n4387), .A(n7172), .B(n9847), .ZN(n9978)
         );
  OAI22_X1 U8887 ( .A1(n9620), .A2(n5022), .B1(n7173), .B2(n9598), .ZN(n7174)
         );
  AOI21_X1 U8888 ( .B1(n9605), .B2(n9975), .A(n7174), .ZN(n7175) );
  OAI21_X1 U8889 ( .B1(n7292), .B2(n9597), .A(n7175), .ZN(n7176) );
  AOI21_X1 U8890 ( .B1(n9844), .B2(n7177), .A(n7176), .ZN(n7178) );
  OAI21_X1 U8891 ( .B1(n9978), .B2(n9530), .A(n7178), .ZN(n7179) );
  AOI21_X1 U8892 ( .B1(n9980), .B2(n9601), .A(n7179), .ZN(n7180) );
  OAI21_X1 U8893 ( .B1(n7181), .B2(n9589), .A(n7180), .ZN(P1_U3283) );
  INV_X1 U8894 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7183) );
  OAI222_X1 U8895 ( .A1(n8019), .A2(n7183), .B1(n9221), .B2(n7182), .C1(n8242), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  NAND2_X1 U8896 ( .A1(n7184), .A2(n8122), .ZN(n7258) );
  OAI21_X1 U8897 ( .B1(n7184), .B2(n8122), .A(n7258), .ZN(n10131) );
  INV_X1 U8898 ( .A(n7249), .ZN(n7185) );
  OAI211_X1 U8899 ( .C1(n8217), .C2(n7186), .A(n7185), .B(n10049), .ZN(n7188)
         );
  AOI22_X1 U8900 ( .A1(n10045), .A2(n8825), .B1(n8823), .B2(n10046), .ZN(n7187) );
  OAI211_X1 U8901 ( .C1(n10131), .C2(n10039), .A(n7188), .B(n7187), .ZN(n10135) );
  NAND2_X1 U8902 ( .A1(n10135), .A2(n9049), .ZN(n7194) );
  INV_X1 U8903 ( .A(n7189), .ZN(n8253) );
  OAI22_X1 U8904 ( .A1(n9049), .A2(n6526), .B1(n8253), .B2(n8975), .ZN(n7192)
         );
  XNOR2_X1 U8905 ( .A(n7190), .B(n10132), .ZN(n10134) );
  NOR2_X1 U8906 ( .A1(n10134), .A2(n8935), .ZN(n7191) );
  AOI211_X1 U8907 ( .C1(n8926), .C2(n10132), .A(n7192), .B(n7191), .ZN(n7193)
         );
  OAI211_X1 U8908 ( .C1(n10131), .C2(n10053), .A(n7194), .B(n7193), .ZN(
        P2_U3286) );
  XNOR2_X1 U8909 ( .A(n7727), .B(n8606), .ZN(n7195) );
  NAND2_X1 U8910 ( .A1(n8820), .A2(n8630), .ZN(n7196) );
  NAND2_X1 U8911 ( .A1(n7195), .A2(n7196), .ZN(n7377) );
  INV_X1 U8912 ( .A(n7195), .ZN(n7198) );
  INV_X1 U8913 ( .A(n7196), .ZN(n7197) );
  NAND2_X1 U8914 ( .A1(n7198), .A2(n7197), .ZN(n7199) );
  NAND2_X1 U8915 ( .A1(n7377), .A2(n7199), .ZN(n7205) );
  AOI21_X1 U8916 ( .B1(n7205), .B2(n7204), .A(n4383), .ZN(n7211) );
  AOI22_X1 U8917 ( .A1(n7206), .A2(n8821), .B1(n7726), .B2(n8784), .ZN(n7208)
         );
  OAI211_X1 U8918 ( .C1(n7906), .C2(n8781), .A(n7208), .B(n7207), .ZN(n7209)
         );
  AOI21_X1 U8919 ( .B1(n7727), .B2(n8809), .A(n7209), .ZN(n7210) );
  OAI21_X1 U8920 ( .B1(n7211), .B2(n8812), .A(n7210), .ZN(P2_U3217) );
  INV_X1 U8921 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7228) );
  NOR2_X1 U8922 ( .A1(n7213), .A2(n7212), .ZN(n7215) );
  NOR2_X1 U8923 ( .A1(n7215), .A2(n7214), .ZN(n7663) );
  INV_X1 U8924 ( .A(n7216), .ZN(n7218) );
  OAI211_X1 U8925 ( .C1(n7218), .C2(P1_REG2_REG_15__SCAN_IN), .A(n9911), .B(
        n4408), .ZN(n7227) );
  NAND2_X1 U8926 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7765) );
  INV_X1 U8927 ( .A(n7765), .ZN(n7223) );
  OAI21_X1 U8928 ( .B1(n7220), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7219), .ZN(
        n7667) );
  XNOR2_X1 U8929 ( .A(n7668), .B(n7667), .ZN(n7221) );
  NOR2_X1 U8930 ( .A1(n9722), .A2(n7221), .ZN(n7669) );
  AOI211_X1 U8931 ( .C1(n7221), .C2(n9722), .A(n7669), .B(n9876), .ZN(n7222)
         );
  AOI211_X1 U8932 ( .C1(n7225), .C2(n7224), .A(n7223), .B(n7222), .ZN(n7226)
         );
  OAI211_X1 U8933 ( .C1(n9924), .C2(n7228), .A(n7227), .B(n7226), .ZN(P1_U3256) );
  NAND2_X1 U8934 ( .A1(n7311), .A2(n8714), .ZN(n7230) );
  NAND2_X1 U8935 ( .A1(n9975), .A2(n8716), .ZN(n7229) );
  NAND2_X1 U8936 ( .A1(n7230), .A2(n7229), .ZN(n7231) );
  XNOR2_X1 U8937 ( .A(n7231), .B(n8689), .ZN(n7233) );
  AND2_X1 U8938 ( .A1(n9975), .A2(n6414), .ZN(n7232) );
  AOI21_X1 U8939 ( .B1(n7311), .B2(n8716), .A(n7232), .ZN(n7234) );
  NAND2_X1 U8940 ( .A1(n7233), .A2(n7234), .ZN(n7365) );
  INV_X1 U8941 ( .A(n7233), .ZN(n7236) );
  INV_X1 U8942 ( .A(n7234), .ZN(n7235) );
  NAND2_X1 U8943 ( .A1(n7236), .A2(n7235), .ZN(n7237) );
  NAND2_X1 U8944 ( .A1(n7365), .A2(n7237), .ZN(n7342) );
  OR2_X1 U8945 ( .A1(n7645), .A2(n7342), .ZN(n7366) );
  INV_X1 U8946 ( .A(n7366), .ZN(n7241) );
  AOI21_X1 U8947 ( .B1(n7342), .B2(n7645), .A(n7241), .ZN(n7247) );
  NOR2_X1 U8948 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7242), .ZN(n9900) );
  NOR2_X1 U8949 ( .A1(n7339), .A2(n9304), .ZN(n7243) );
  AOI211_X1 U8950 ( .C1(n9302), .C2(n9984), .A(n9900), .B(n7243), .ZN(n7244)
         );
  OAI21_X1 U8951 ( .B1(n9262), .B2(n7306), .A(n7244), .ZN(n7245) );
  AOI21_X1 U8952 ( .B1(n9320), .B2(n7311), .A(n7245), .ZN(n7246) );
  OAI21_X1 U8953 ( .B1(n7247), .B2(n9315), .A(n7246), .ZN(P1_U3229) );
  OR2_X1 U8954 ( .A1(n7249), .A2(n7248), .ZN(n7250) );
  XNOR2_X1 U8955 ( .A(n7250), .B(n8219), .ZN(n7253) );
  NAND2_X1 U8956 ( .A1(n8824), .A2(n10045), .ZN(n7252) );
  NAND2_X1 U8957 ( .A1(n8822), .A2(n10046), .ZN(n7251) );
  NAND2_X1 U8958 ( .A1(n7252), .A2(n7251), .ZN(n8795) );
  AOI21_X1 U8959 ( .B1(n7253), .B2(n10049), .A(n8795), .ZN(n10144) );
  AOI211_X1 U8960 ( .C1(n10141), .C2(n7254), .A(n10055), .B(n7328), .ZN(n10140) );
  INV_X1 U8961 ( .A(n10141), .ZN(n7256) );
  AOI22_X1 U8962 ( .A1(n10070), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n8796), .B2(
        n10062), .ZN(n7255) );
  OAI21_X1 U8963 ( .B1(n7256), .B2(n10054), .A(n7255), .ZN(n7264) );
  NAND2_X1 U8964 ( .A1(n7258), .A2(n7257), .ZN(n7262) );
  NAND2_X1 U8965 ( .A1(n7184), .A2(n7259), .ZN(n7261) );
  AND2_X1 U8966 ( .A1(n7261), .A2(n7260), .ZN(n7322) );
  OAI21_X1 U8967 ( .B1(n7262), .B2(n8219), .A(n7322), .ZN(n10145) );
  NOR2_X1 U8968 ( .A1(n10145), .A2(n9126), .ZN(n7263) );
  AOI211_X1 U8969 ( .C1(n9124), .C2(n10140), .A(n7264), .B(n7263), .ZN(n7265)
         );
  OAI21_X1 U8970 ( .B1(n10070), .B2(n10144), .A(n7265), .ZN(P2_U3285) );
  OAI21_X1 U8971 ( .B1(n7267), .B2(P2_REG1_REG_14__SCAN_IN), .A(n7266), .ZN(
        n7872) );
  XNOR2_X1 U8972 ( .A(n7872), .B(n7873), .ZN(n7268) );
  INV_X1 U8973 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9806) );
  NOR2_X1 U8974 ( .A1(n9806), .A2(n7268), .ZN(n7874) );
  AOI211_X1 U8975 ( .C1(n7268), .C2(n9806), .A(n7874), .B(n10032), .ZN(n7278)
         );
  AOI21_X1 U8976 ( .B1(n7271), .B2(n7270), .A(n7269), .ZN(n7865) );
  XNOR2_X1 U8977 ( .A(n7865), .B(n7866), .ZN(n7272) );
  NOR2_X1 U8978 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7272), .ZN(n7867) );
  AOI21_X1 U8979 ( .B1(n7272), .B2(P2_REG2_REG_15__SCAN_IN), .A(n7867), .ZN(
        n7273) );
  NOR2_X1 U8980 ( .A1(n7273), .A2(n7886), .ZN(n7277) );
  NOR2_X1 U8981 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5758), .ZN(n7274) );
  AOI21_X1 U8982 ( .B1(n10034), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7274), .ZN(
        n7275) );
  OAI21_X1 U8983 ( .B1(n10030), .B2(n7873), .A(n7275), .ZN(n7276) );
  OR3_X1 U8984 ( .A1(n7278), .A2(n7277), .A3(n7276), .ZN(P2_U3260) );
  NAND2_X1 U8985 ( .A1(n7279), .A2(n9513), .ZN(n7280) );
  OR2_X1 U8986 ( .A1(n9939), .A2(n7280), .ZN(n9632) );
  INV_X1 U8987 ( .A(n9632), .ZN(n9851) );
  OAI21_X1 U8988 ( .B1(n7282), .B2(n8306), .A(n7281), .ZN(n9955) );
  AOI21_X1 U8989 ( .B1(n7283), .B2(n7288), .A(n9622), .ZN(n7285) );
  NAND2_X1 U8990 ( .A1(n7285), .A2(n7284), .ZN(n9956) );
  INV_X1 U8991 ( .A(n7286), .ZN(n7287) );
  AOI22_X1 U8992 ( .A1(n9844), .A2(n7288), .B1(n7287), .B2(n9936), .ZN(n7289)
         );
  OAI21_X1 U8993 ( .B1(n9956), .B2(n9530), .A(n7289), .ZN(n7299) );
  NAND2_X1 U8994 ( .A1(n7290), .A2(n8479), .ZN(n7291) );
  XNOR2_X1 U8995 ( .A(n7291), .B(n8306), .ZN(n7297) );
  NAND2_X1 U8996 ( .A1(n9955), .A2(n9860), .ZN(n7296) );
  OAI22_X1 U8997 ( .A1(n7293), .A2(n9964), .B1(n7292), .B2(n9962), .ZN(n7294)
         );
  INV_X1 U8998 ( .A(n7294), .ZN(n7295) );
  OAI211_X1 U8999 ( .C1(n9972), .C2(n7297), .A(n7296), .B(n7295), .ZN(n9960)
         );
  MUX2_X1 U9000 ( .A(n9960), .B(P1_REG2_REG_6__SCAN_IN), .S(n9939), .Z(n7298)
         );
  AOI211_X1 U9001 ( .C1(n9851), .C2(n9955), .A(n7299), .B(n7298), .ZN(n7300)
         );
  INV_X1 U9002 ( .A(n7300), .ZN(P1_U3285) );
  NAND2_X1 U9003 ( .A1(n8324), .A2(n8320), .ZN(n8438) );
  INV_X1 U9004 ( .A(n8438), .ZN(n7302) );
  XNOR2_X1 U9005 ( .A(n7301), .B(n7302), .ZN(n9993) );
  INV_X1 U9006 ( .A(n9993), .ZN(n7315) );
  OR2_X1 U9007 ( .A1(n7303), .A2(n7302), .ZN(n7304) );
  NAND2_X1 U9008 ( .A1(n7303), .A2(n7302), .ZN(n7391) );
  AND3_X1 U9009 ( .A1(n7304), .A2(n7391), .A3(n9693), .ZN(n9991) );
  OAI211_X1 U9010 ( .C1(n7305), .C2(n9989), .A(n7385), .B(n9847), .ZN(n9987)
         );
  INV_X1 U9011 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7307) );
  OAI22_X1 U9012 ( .A1(n9620), .A2(n7307), .B1(n7306), .B2(n9598), .ZN(n7308)
         );
  AOI21_X1 U9013 ( .B1(n9605), .B2(n9983), .A(n7308), .ZN(n7309) );
  OAI21_X1 U9014 ( .B1(n9963), .B2(n9597), .A(n7309), .ZN(n7310) );
  AOI21_X1 U9015 ( .B1(n9844), .B2(n7311), .A(n7310), .ZN(n7312) );
  OAI21_X1 U9016 ( .B1(n9987), .B2(n9530), .A(n7312), .ZN(n7313) );
  AOI21_X1 U9017 ( .B1(n9991), .B2(n9601), .A(n7313), .ZN(n7314) );
  OAI21_X1 U9018 ( .B1(n7315), .B2(n9589), .A(n7314), .ZN(P1_U3282) );
  INV_X1 U9019 ( .A(n8070), .ZN(n7316) );
  NOR2_X1 U9020 ( .A1(n7317), .A2(n7316), .ZN(n7318) );
  XNOR2_X1 U9021 ( .A(n7318), .B(n7323), .ZN(n7320) );
  OAI21_X1 U9022 ( .B1(n7320), .B2(n9071), .A(n7319), .ZN(n10152) );
  INV_X1 U9023 ( .A(n10152), .ZN(n7335) );
  NAND2_X1 U9024 ( .A1(n7322), .A2(n7321), .ZN(n7324) );
  INV_X1 U9025 ( .A(n7324), .ZN(n7326) );
  OR2_X1 U9026 ( .A1(n7324), .A2(n7323), .ZN(n7325) );
  OAI21_X1 U9027 ( .B1(n7326), .B2(n8220), .A(n7325), .ZN(n10154) );
  INV_X1 U9028 ( .A(n7627), .ZN(n7327) );
  OAI211_X1 U9029 ( .C1(n10151), .C2(n7328), .A(n7327), .B(n5952), .ZN(n10149)
         );
  AOI22_X1 U9030 ( .A1(n10070), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7329), .B2(
        n10062), .ZN(n7332) );
  NAND2_X1 U9031 ( .A1(n7330), .A2(n8926), .ZN(n7331) );
  OAI211_X1 U9032 ( .C1(n10149), .C2(n10065), .A(n7332), .B(n7331), .ZN(n7333)
         );
  AOI21_X1 U9033 ( .B1(n10154), .B2(n9082), .A(n7333), .ZN(n7334) );
  OAI21_X1 U9034 ( .B1(n7335), .B2(n10070), .A(n7334), .ZN(P2_U3284) );
  INV_X1 U9035 ( .A(n9845), .ZN(n9867) );
  NAND2_X1 U9036 ( .A1(n9785), .A2(n8714), .ZN(n7337) );
  OR2_X1 U9037 ( .A1(n7339), .A2(n6498), .ZN(n7336) );
  NAND2_X1 U9038 ( .A1(n7337), .A2(n7336), .ZN(n7338) );
  XNOR2_X1 U9039 ( .A(n7338), .B(n8721), .ZN(n7343) );
  NAND2_X1 U9040 ( .A1(n9785), .A2(n8716), .ZN(n7341) );
  OR2_X1 U9041 ( .A1(n7339), .A2(n8719), .ZN(n7340) );
  NAND2_X1 U9042 ( .A1(n7341), .A2(n7340), .ZN(n7344) );
  NAND2_X1 U9043 ( .A1(n7343), .A2(n7344), .ZN(n7368) );
  INV_X1 U9044 ( .A(n7368), .ZN(n7348) );
  OR2_X1 U9045 ( .A1(n7342), .A2(n7348), .ZN(n7641) );
  OR2_X1 U9046 ( .A1(n7645), .A2(n7641), .ZN(n7357) );
  INV_X1 U9047 ( .A(n7343), .ZN(n7346) );
  INV_X1 U9048 ( .A(n7344), .ZN(n7345) );
  NAND2_X1 U9049 ( .A1(n7346), .A2(n7345), .ZN(n7367) );
  AND2_X1 U9050 ( .A1(n7365), .A2(n7367), .ZN(n7347) );
  OR2_X1 U9051 ( .A1(n7348), .A2(n7347), .ZN(n7356) );
  NAND2_X1 U9052 ( .A1(n7357), .A2(n7356), .ZN(n7353) );
  NAND2_X1 U9053 ( .A1(n9845), .A2(n8714), .ZN(n7350) );
  OR2_X1 U9054 ( .A1(n7794), .A2(n6498), .ZN(n7349) );
  NAND2_X1 U9055 ( .A1(n7350), .A2(n7349), .ZN(n7351) );
  XNOR2_X1 U9056 ( .A(n7351), .B(n8689), .ZN(n7640) );
  NOR2_X1 U9057 ( .A1(n7794), .A2(n8719), .ZN(n7352) );
  AOI21_X1 U9058 ( .B1(n9845), .B2(n8716), .A(n7352), .ZN(n7639) );
  XNOR2_X1 U9059 ( .A(n7640), .B(n7639), .ZN(n7354) );
  AOI21_X1 U9060 ( .B1(n7353), .B2(n7354), .A(n9315), .ZN(n7359) );
  INV_X1 U9061 ( .A(n7354), .ZN(n7355) );
  AND2_X1 U9062 ( .A1(n7356), .A2(n7355), .ZN(n7642) );
  NAND2_X1 U9063 ( .A1(n7357), .A2(n7642), .ZN(n7358) );
  NAND2_X1 U9064 ( .A1(n7359), .A2(n7358), .ZN(n7363) );
  NAND2_X1 U9065 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3084), .ZN(n9336) );
  OAI21_X1 U9066 ( .B1(n7688), .B2(n9304), .A(n9336), .ZN(n7361) );
  NOR2_X1 U9067 ( .A1(n9282), .A2(n9842), .ZN(n7360) );
  AOI211_X1 U9068 ( .C1(n9302), .C2(n9983), .A(n7361), .B(n7360), .ZN(n7362)
         );
  OAI211_X1 U9069 ( .C1(n9867), .C2(n7364), .A(n7363), .B(n7362), .ZN(P1_U3234) );
  NAND2_X1 U9070 ( .A1(n7366), .A2(n7365), .ZN(n7370) );
  NAND2_X1 U9071 ( .A1(n7368), .A2(n7367), .ZN(n7369) );
  XNOR2_X1 U9072 ( .A(n7370), .B(n7369), .ZN(n7376) );
  OAI21_X1 U9073 ( .B1(n7794), .B2(n9304), .A(n7371), .ZN(n7372) );
  AOI21_X1 U9074 ( .B1(n9302), .B2(n9975), .A(n7372), .ZN(n7373) );
  OAI21_X1 U9075 ( .B1(n9282), .B2(n7387), .A(n7373), .ZN(n7374) );
  AOI21_X1 U9076 ( .B1(n9320), .B2(n9785), .A(n7374), .ZN(n7375) );
  OAI21_X1 U9077 ( .B1(n7376), .B2(n9315), .A(n7375), .ZN(P1_U3215) );
  XNOR2_X1 U9078 ( .A(n7895), .B(n8631), .ZN(n7702) );
  AND2_X1 U9079 ( .A1(n8819), .A2(n10055), .ZN(n7699) );
  XNOR2_X1 U9080 ( .A(n7700), .B(n7699), .ZN(n7382) );
  OAI22_X1 U9081 ( .A1(n8781), .A2(n7955), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5758), .ZN(n7380) );
  INV_X1 U9082 ( .A(n7894), .ZN(n7378) );
  OAI22_X1 U9083 ( .A1(n8805), .A2(n7891), .B1(n10026), .B2(n7378), .ZN(n7379)
         );
  AOI211_X1 U9084 ( .C1(n7895), .C2(n8809), .A(n7380), .B(n7379), .ZN(n7381)
         );
  OAI21_X1 U9085 ( .B1(n7382), .B2(n8812), .A(n7381), .ZN(P2_U3243) );
  XOR2_X1 U9086 ( .A(n7383), .B(n8439), .Z(n9788) );
  AOI211_X1 U9087 ( .C1(n9785), .C2(n7385), .A(n9622), .B(n5443), .ZN(n9784)
         );
  INV_X1 U9088 ( .A(n9785), .ZN(n7386) );
  NOR2_X1 U9089 ( .A1(n7386), .A2(n9628), .ZN(n7390) );
  OAI22_X1 U9090 ( .A1(n9620), .A2(n7388), .B1(n7387), .B2(n9598), .ZN(n7389)
         );
  AOI211_X1 U9091 ( .C1(n9784), .C2(n9850), .A(n7390), .B(n7389), .ZN(n7397)
         );
  NAND2_X1 U9092 ( .A1(n7391), .A2(n8324), .ZN(n7392) );
  XNOR2_X1 U9093 ( .A(n7392), .B(n8439), .ZN(n7393) );
  NAND2_X1 U9094 ( .A1(n7393), .A2(n9693), .ZN(n7395) );
  AOI22_X1 U9095 ( .A1(n9855), .A2(n5499), .B1(n9985), .B2(n9975), .ZN(n7394)
         );
  NAND2_X1 U9096 ( .A1(n7395), .A2(n7394), .ZN(n9783) );
  NAND2_X1 U9097 ( .A1(n9783), .A2(n9620), .ZN(n7396) );
  OAI211_X1 U9098 ( .C1(n9788), .C2(n9589), .A(n7397), .B(n7396), .ZN(P1_U3281) );
  INV_X1 U9099 ( .A(n7398), .ZN(n8017) );
  OAI222_X1 U9100 ( .A1(n9777), .A2(n7400), .B1(n7846), .B2(n8017), .C1(n7399), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  INV_X1 U9101 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10213) );
  NOR2_X1 U9102 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7401) );
  AOI21_X1 U9103 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7401), .ZN(n10184) );
  NOR2_X1 U9104 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7402) );
  AOI21_X1 U9105 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7402), .ZN(n10187) );
  NOR2_X1 U9106 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7403) );
  AOI21_X1 U9107 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7403), .ZN(n10190) );
  NOR2_X1 U9108 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7404) );
  AOI21_X1 U9109 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7404), .ZN(n10193) );
  NOR2_X1 U9110 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7405) );
  AOI21_X1 U9111 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7405), .ZN(n10196) );
  NOR2_X1 U9112 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7411) );
  XNOR2_X1 U9113 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10223) );
  NAND2_X1 U9114 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7409) );
  XOR2_X1 U9115 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10221) );
  NAND2_X1 U9116 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7407) );
  XOR2_X1 U9117 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10209) );
  AOI21_X1 U9118 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10177) );
  INV_X1 U9119 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10181) );
  NAND3_X1 U9120 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10179) );
  OAI21_X1 U9121 ( .B1(n10177), .B2(n10181), .A(n10179), .ZN(n10208) );
  NAND2_X1 U9122 ( .A1(n10209), .A2(n10208), .ZN(n7406) );
  NAND2_X1 U9123 ( .A1(n7407), .A2(n7406), .ZN(n10220) );
  NAND2_X1 U9124 ( .A1(n10221), .A2(n10220), .ZN(n7408) );
  NAND2_X1 U9125 ( .A1(n7409), .A2(n7408), .ZN(n10222) );
  NOR2_X1 U9126 ( .A1(n10223), .A2(n10222), .ZN(n7410) );
  NOR2_X1 U9127 ( .A1(n7411), .A2(n7410), .ZN(n10218) );
  NAND2_X1 U9128 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10218), .ZN(n7412) );
  NOR2_X1 U9129 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10218), .ZN(n10217) );
  AOI21_X1 U9130 ( .B1(n7413), .B2(n7412), .A(n10217), .ZN(n7414) );
  NAND2_X1 U9131 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n7414), .ZN(n7416) );
  XOR2_X1 U9132 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n7414), .Z(n10216) );
  NAND2_X1 U9133 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10216), .ZN(n7415) );
  NAND2_X1 U9134 ( .A1(n7416), .A2(n7415), .ZN(n7417) );
  NAND2_X1 U9135 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7417), .ZN(n7420) );
  XNOR2_X1 U9136 ( .A(n7418), .B(n7417), .ZN(n10215) );
  NAND2_X1 U9137 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10215), .ZN(n7419) );
  NAND2_X1 U9138 ( .A1(n7420), .A2(n7419), .ZN(n7421) );
  NAND2_X1 U9139 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7421), .ZN(n7423) );
  XOR2_X1 U9140 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7421), .Z(n10210) );
  NAND2_X1 U9141 ( .A1(n10210), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7422) );
  NAND2_X1 U9142 ( .A1(n7423), .A2(n7422), .ZN(n10206) );
  AOI222_X1 U9143 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .B1(P2_ADDR_REG_9__SCAN_IN), .B2(n10206), .C1(P1_ADDR_REG_9__SCAN_IN), 
        .C2(n10206), .ZN(n10205) );
  NAND2_X1 U9144 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7424) );
  OAI21_X1 U9145 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7424), .ZN(n10204) );
  NOR2_X1 U9146 ( .A1(n10205), .A2(n10204), .ZN(n10203) );
  AOI21_X1 U9147 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10203), .ZN(n10202) );
  NAND2_X1 U9148 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7425) );
  OAI21_X1 U9149 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7425), .ZN(n10201) );
  NOR2_X1 U9150 ( .A1(n10202), .A2(n10201), .ZN(n10200) );
  AOI21_X1 U9151 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10200), .ZN(n10199) );
  NOR2_X1 U9152 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7426) );
  AOI21_X1 U9153 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7426), .ZN(n10198) );
  NAND2_X1 U9154 ( .A1(n10199), .A2(n10198), .ZN(n10197) );
  OAI21_X1 U9155 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10197), .ZN(n10195) );
  NAND2_X1 U9156 ( .A1(n10196), .A2(n10195), .ZN(n10194) );
  OAI21_X1 U9157 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10194), .ZN(n10192) );
  NAND2_X1 U9158 ( .A1(n10193), .A2(n10192), .ZN(n10191) );
  OAI21_X1 U9159 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10191), .ZN(n10189) );
  NAND2_X1 U9160 ( .A1(n10190), .A2(n10189), .ZN(n10188) );
  OAI21_X1 U9161 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10188), .ZN(n10186) );
  NAND2_X1 U9162 ( .A1(n10187), .A2(n10186), .ZN(n10185) );
  OAI21_X1 U9163 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10185), .ZN(n10183) );
  NAND2_X1 U9164 ( .A1(n10184), .A2(n10183), .ZN(n10182) );
  OAI21_X1 U9165 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10182), .ZN(n10212) );
  NOR2_X1 U9166 ( .A1(n10213), .A2(n10212), .ZN(n7427) );
  NAND2_X1 U9167 ( .A1(n10213), .A2(n10212), .ZN(n10211) );
  OAI21_X1 U9168 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7427), .A(n10211), .ZN(
        n7617) );
  AOI22_X1 U9169 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_f61), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .ZN(n7428) );
  OAI221_X1 U9170 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_f58), .A(n7428), .ZN(n7436) );
  AOI22_X1 U9171 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_f43), .B1(SI_18_), 
        .B2(keyinput_f14), .ZN(n7429) );
  OAI221_X1 U9172 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .C1(SI_18_), .C2(keyinput_f14), .A(n7429), .ZN(n7435) );
  AOI22_X1 U9173 ( .A1(n7431), .A2(keyinput_f44), .B1(keyinput_f3), .B2(n7589), 
        .ZN(n7430) );
  OAI221_X1 U9174 ( .B1(n7431), .B2(keyinput_f44), .C1(n7589), .C2(keyinput_f3), .A(n7430), .ZN(n7434) );
  AOI22_X1 U9175 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput_f52), .B1(n5694), 
        .B2(keyinput_f53), .ZN(n7432) );
  OAI221_X1 U9176 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_f52), .C1(n5694), 
        .C2(keyinput_f53), .A(n7432), .ZN(n7433) );
  NOR4_X1 U9177 ( .A1(n7436), .A2(n7435), .A3(n7434), .A4(n7433), .ZN(n7507)
         );
  AOI22_X1 U9178 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_f46), .B1(SI_15_), .B2(keyinput_f17), .ZN(n7437) );
  OAI221_X1 U9179 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .C1(
        SI_15_), .C2(keyinput_f17), .A(n7437), .ZN(n7444) );
  AOI22_X1 U9180 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_f40), .B1(SI_9_), 
        .B2(keyinput_f23), .ZN(n7438) );
  OAI221_X1 U9181 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .C1(SI_9_), 
        .C2(keyinput_f23), .A(n7438), .ZN(n7443) );
  AOI22_X1 U9182 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_f54), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(keyinput_f50), .ZN(n7439) );
  OAI221_X1 U9183 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_f54), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_f50), .A(n7439), .ZN(n7442) );
  AOI22_X1 U9184 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_f60), .B1(SI_21_), .B2(keyinput_f11), .ZN(n7440) );
  OAI221_X1 U9185 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .C1(
        SI_21_), .C2(keyinput_f11), .A(n7440), .ZN(n7441) );
  NOR4_X1 U9186 ( .A1(n7444), .A2(n7443), .A3(n7442), .A4(n7441), .ZN(n7506)
         );
  AOI22_X1 U9187 ( .A1(keyinput_f0), .A2(P2_WR_REG_SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_f34), .ZN(n7445) );
  OAI221_X1 U9188 ( .B1(keyinput_f0), .B2(P2_WR_REG_SCAN_IN), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_f34), .A(n7445), .ZN(n7504) );
  AOI22_X1 U9189 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_f51), .B1(SI_2_), 
        .B2(keyinput_f30), .ZN(n7446) );
  OAI221_X1 U9190 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .C1(SI_2_), .C2(keyinput_f30), .A(n7446), .ZN(n7503) );
  AOI22_X1 U9191 ( .A1(SI_6_), .A2(keyinput_f26), .B1(n7448), .B2(keyinput_f49), .ZN(n7447) );
  OAI221_X1 U9192 ( .B1(SI_6_), .B2(keyinput_f26), .C1(n7448), .C2(
        keyinput_f49), .A(n7447), .ZN(n7458) );
  OAI22_X1 U9193 ( .A1(SI_5_), .A2(keyinput_f27), .B1(keyinput_f36), .B2(
        P2_REG3_REG_27__SCAN_IN), .ZN(n7449) );
  AOI221_X1 U9194 ( .B1(SI_5_), .B2(keyinput_f27), .C1(P2_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n7449), .ZN(n7456) );
  OAI22_X1 U9195 ( .A1(SI_22_), .A2(keyinput_f10), .B1(keyinput_f12), .B2(
        SI_20_), .ZN(n7450) );
  AOI221_X1 U9196 ( .B1(SI_22_), .B2(keyinput_f10), .C1(SI_20_), .C2(
        keyinput_f12), .A(n7450), .ZN(n7455) );
  OAI22_X1 U9197 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_f42), .B1(
        keyinput_f63), .B2(P2_REG3_REG_15__SCAN_IN), .ZN(n7451) );
  AOI221_X1 U9198 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput_f63), .A(n7451), .ZN(n7454) );
  OAI22_X1 U9199 ( .A1(SI_7_), .A2(keyinput_f25), .B1(keyinput_f29), .B2(SI_3_), .ZN(n7452) );
  AOI221_X1 U9200 ( .B1(SI_7_), .B2(keyinput_f25), .C1(SI_3_), .C2(
        keyinput_f29), .A(n7452), .ZN(n7453) );
  NAND4_X1 U9201 ( .A1(n7456), .A2(n7455), .A3(n7454), .A4(n7453), .ZN(n7457)
         );
  AOI211_X1 U9202 ( .C1(keyinput_f22), .C2(SI_10_), .A(n7458), .B(n7457), .ZN(
        n7459) );
  OAI21_X1 U9203 ( .B1(keyinput_f22), .B2(SI_10_), .A(n7459), .ZN(n7502) );
  INV_X1 U9204 ( .A(SI_11_), .ZN(n7553) );
  AOI22_X1 U9205 ( .A1(n7553), .A2(keyinput_f21), .B1(keyinput_f57), .B2(n8780), .ZN(n7460) );
  OAI221_X1 U9206 ( .B1(n7553), .B2(keyinput_f21), .C1(n8780), .C2(
        keyinput_f57), .A(n7460), .ZN(n7467) );
  INV_X1 U9207 ( .A(SI_24_), .ZN(n7591) );
  INV_X1 U9208 ( .A(SI_14_), .ZN(n7551) );
  AOI22_X1 U9209 ( .A1(n7591), .A2(keyinput_f8), .B1(keyinput_f18), .B2(n7551), 
        .ZN(n7461) );
  OAI221_X1 U9210 ( .B1(n7591), .B2(keyinput_f8), .C1(n7551), .C2(keyinput_f18), .A(n7461), .ZN(n7466) );
  AOI22_X1 U9211 ( .A1(n7569), .A2(keyinput_f24), .B1(n7579), .B2(keyinput_f9), 
        .ZN(n7462) );
  OAI221_X1 U9212 ( .B1(n7569), .B2(keyinput_f24), .C1(n7579), .C2(keyinput_f9), .A(n7462), .ZN(n7465) );
  AOI22_X1 U9213 ( .A1(n8804), .A2(keyinput_f62), .B1(keyinput_f55), .B2(n8004), .ZN(n7463) );
  OAI221_X1 U9214 ( .B1(n8804), .B2(keyinput_f62), .C1(n8004), .C2(
        keyinput_f55), .A(n7463), .ZN(n7464) );
  NOR4_X1 U9215 ( .A1(n7467), .A2(n7466), .A3(n7465), .A4(n7464), .ZN(n7500)
         );
  INV_X1 U9216 ( .A(SI_26_), .ZN(n7554) );
  AOI22_X1 U9217 ( .A1(n7554), .A2(keyinput_f6), .B1(keyinput_f35), .B2(n5669), 
        .ZN(n7468) );
  OAI221_X1 U9218 ( .B1(n7554), .B2(keyinput_f6), .C1(n5669), .C2(keyinput_f35), .A(n7468), .ZN(n7476) );
  AOI22_X1 U9219 ( .A1(n8759), .A2(keyinput_f47), .B1(keyinput_f39), .B2(n8271), .ZN(n7469) );
  OAI221_X1 U9220 ( .B1(n8759), .B2(keyinput_f47), .C1(n8271), .C2(
        keyinput_f39), .A(n7469), .ZN(n7475) );
  INV_X1 U9221 ( .A(SI_12_), .ZN(n7578) );
  XOR2_X1 U9222 ( .A(n7578), .B(keyinput_f20), .Z(n7473) );
  XNOR2_X1 U9223 ( .A(SI_27_), .B(keyinput_f5), .ZN(n7472) );
  XNOR2_X1 U9224 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_f33), .ZN(n7471) );
  XNOR2_X1 U9225 ( .A(SI_1_), .B(keyinput_f31), .ZN(n7470) );
  NAND4_X1 U9226 ( .A1(n7473), .A2(n7472), .A3(n7471), .A4(n7470), .ZN(n7474)
         );
  NOR3_X1 U9227 ( .A1(n7476), .A2(n7475), .A3(n7474), .ZN(n7499) );
  INV_X1 U9228 ( .A(SI_19_), .ZN(n7596) );
  AOI22_X1 U9229 ( .A1(n7596), .A2(keyinput_f13), .B1(keyinput_f4), .B2(n5898), 
        .ZN(n7477) );
  OAI221_X1 U9230 ( .B1(n7596), .B2(keyinput_f13), .C1(n5898), .C2(keyinput_f4), .A(n7477), .ZN(n7485) );
  AOI22_X1 U9231 ( .A1(n7566), .A2(keyinput_f48), .B1(n7479), .B2(keyinput_f15), .ZN(n7478) );
  OAI221_X1 U9232 ( .B1(n7566), .B2(keyinput_f48), .C1(n7479), .C2(
        keyinput_f15), .A(n7478), .ZN(n7484) );
  AOI22_X1 U9233 ( .A1(n7582), .A2(keyinput_f19), .B1(n7564), .B2(keyinput_f7), 
        .ZN(n7480) );
  OAI221_X1 U9234 ( .B1(n7582), .B2(keyinput_f19), .C1(n7564), .C2(keyinput_f7), .A(n7480), .ZN(n7483) );
  AOI22_X1 U9235 ( .A1(n8743), .A2(keyinput_f38), .B1(n7525), .B2(keyinput_f16), .ZN(n7481) );
  OAI221_X1 U9236 ( .B1(n8743), .B2(keyinput_f38), .C1(n7525), .C2(
        keyinput_f16), .A(n7481), .ZN(n7482) );
  NOR4_X1 U9237 ( .A1(n7485), .A2(n7484), .A3(n7483), .A4(n7482), .ZN(n7498)
         );
  AOI22_X1 U9238 ( .A1(n7487), .A2(keyinput_f41), .B1(keyinput_f56), .B2(n6781), .ZN(n7486) );
  OAI221_X1 U9239 ( .B1(n7487), .B2(keyinput_f41), .C1(n6781), .C2(
        keyinput_f56), .A(n7486), .ZN(n7496) );
  AOI22_X1 U9240 ( .A1(n8039), .A2(keyinput_f2), .B1(n8750), .B2(keyinput_f45), 
        .ZN(n7488) );
  OAI221_X1 U9241 ( .B1(n8039), .B2(keyinput_f2), .C1(n8750), .C2(keyinput_f45), .A(n7488), .ZN(n7495) );
  AOI22_X1 U9242 ( .A1(n7490), .A2(keyinput_f59), .B1(n7556), .B2(keyinput_f37), .ZN(n7489) );
  OAI221_X1 U9243 ( .B1(n7490), .B2(keyinput_f59), .C1(n7556), .C2(
        keyinput_f37), .A(n7489), .ZN(n7494) );
  XNOR2_X1 U9244 ( .A(SI_0_), .B(keyinput_f32), .ZN(n7492) );
  XNOR2_X1 U9245 ( .A(SI_31_), .B(keyinput_f1), .ZN(n7491) );
  NAND2_X1 U9246 ( .A1(n7492), .A2(n7491), .ZN(n7493) );
  NOR4_X1 U9247 ( .A1(n7496), .A2(n7495), .A3(n7494), .A4(n7493), .ZN(n7497)
         );
  NAND4_X1 U9248 ( .A1(n7500), .A2(n7499), .A3(n7498), .A4(n7497), .ZN(n7501)
         );
  NOR4_X1 U9249 ( .A1(n7504), .A2(n7503), .A3(n7502), .A4(n7501), .ZN(n7505)
         );
  NAND3_X1 U9250 ( .A1(n7507), .A2(n7506), .A3(n7505), .ZN(n7510) );
  INV_X1 U9251 ( .A(keyinput_f28), .ZN(n7509) );
  INV_X1 U9252 ( .A(keyinput_g28), .ZN(n7508) );
  AOI21_X1 U9253 ( .B1(n7510), .B2(n7509), .A(n7508), .ZN(n7513) );
  AOI21_X1 U9254 ( .B1(keyinput_f28), .B2(n7510), .A(keyinput_g28), .ZN(n7512)
         );
  MUX2_X1 U9255 ( .A(n7513), .B(n7512), .S(n7511), .Z(n7611) );
  OAI22_X1 U9256 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_g33), .B1(SI_20_), 
        .B2(keyinput_g12), .ZN(n7514) );
  AOI221_X1 U9257 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput_g33), .C1(
        keyinput_g12), .C2(SI_20_), .A(n7514), .ZN(n7521) );
  OAI22_X1 U9258 ( .A1(SI_0_), .A2(keyinput_g32), .B1(keyinput_g34), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n7515) );
  AOI221_X1 U9259 ( .B1(SI_0_), .B2(keyinput_g32), .C1(P2_STATE_REG_SCAN_IN), 
        .C2(keyinput_g34), .A(n7515), .ZN(n7520) );
  OAI22_X1 U9260 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_g43), .B1(SI_31_), 
        .B2(keyinput_g1), .ZN(n7516) );
  AOI221_X1 U9261 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_g43), .C1(
        keyinput_g1), .C2(SI_31_), .A(n7516), .ZN(n7519) );
  OAI22_X1 U9262 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_g49), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(keyinput_g40), .ZN(n7517) );
  AOI221_X1 U9263 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .C1(
        keyinput_g40), .C2(P2_REG3_REG_3__SCAN_IN), .A(n7517), .ZN(n7518) );
  NAND4_X1 U9264 ( .A1(n7521), .A2(n7520), .A3(n7519), .A4(n7518), .ZN(n7549)
         );
  OAI22_X1 U9265 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_g36), .B1(
        keyinput_g50), .B2(P2_REG3_REG_17__SCAN_IN), .ZN(n7522) );
  AOI221_X1 U9266 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_g50), .A(n7522), .ZN(n7529) );
  OAI22_X1 U9267 ( .A1(SI_18_), .A2(keyinput_g14), .B1(SI_10_), .B2(
        keyinput_g22), .ZN(n7523) );
  AOI221_X1 U9268 ( .B1(SI_18_), .B2(keyinput_g14), .C1(keyinput_g22), .C2(
        SI_10_), .A(n7523), .ZN(n7528) );
  OAI22_X1 U9269 ( .A1(SI_9_), .A2(keyinput_g23), .B1(P2_REG3_REG_11__SCAN_IN), 
        .B2(keyinput_g58), .ZN(n7524) );
  AOI221_X1 U9270 ( .B1(SI_9_), .B2(keyinput_g23), .C1(keyinput_g58), .C2(
        P2_REG3_REG_11__SCAN_IN), .A(n7524), .ZN(n7527) );
  XOR2_X1 U9271 ( .A(n7525), .B(keyinput_g16), .Z(n7526) );
  NAND4_X1 U9272 ( .A1(n7529), .A2(n7528), .A3(n7527), .A4(n7526), .ZN(n7548)
         );
  OAI22_X1 U9273 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_g60), .B1(
        keyinput_g46), .B2(P2_REG3_REG_12__SCAN_IN), .ZN(n7530) );
  AOI221_X1 U9274 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_g46), .A(n7530), .ZN(n7537) );
  OAI22_X1 U9275 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_g47), .B1(
        keyinput_g55), .B2(P2_REG3_REG_20__SCAN_IN), .ZN(n7531) );
  AOI221_X1 U9276 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput_g55), .A(n7531), .ZN(n7536) );
  OAI22_X1 U9277 ( .A1(SI_27_), .A2(keyinput_g5), .B1(P2_REG3_REG_19__SCAN_IN), 
        .B2(keyinput_g41), .ZN(n7532) );
  AOI221_X1 U9278 ( .B1(SI_27_), .B2(keyinput_g5), .C1(keyinput_g41), .C2(
        P2_REG3_REG_19__SCAN_IN), .A(n7532), .ZN(n7535) );
  OAI22_X1 U9279 ( .A1(SI_17_), .A2(keyinput_g15), .B1(keyinput_g44), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n7533) );
  AOI221_X1 U9280 ( .B1(SI_17_), .B2(keyinput_g15), .C1(P2_REG3_REG_1__SCAN_IN), .C2(keyinput_g44), .A(n7533), .ZN(n7534) );
  NAND4_X1 U9281 ( .A1(n7537), .A2(n7536), .A3(n7535), .A4(n7534), .ZN(n7547)
         );
  OAI22_X1 U9282 ( .A1(SI_21_), .A2(keyinput_g11), .B1(keyinput_g59), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n7538) );
  AOI221_X1 U9283 ( .B1(SI_21_), .B2(keyinput_g11), .C1(P2_REG3_REG_2__SCAN_IN), .C2(keyinput_g59), .A(n7538), .ZN(n7545) );
  OAI22_X1 U9284 ( .A1(SI_15_), .A2(keyinput_g17), .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .ZN(n7539) );
  AOI221_X1 U9285 ( .B1(SI_15_), .B2(keyinput_g17), .C1(keyinput_g51), .C2(
        P2_REG3_REG_24__SCAN_IN), .A(n7539), .ZN(n7544) );
  OAI22_X1 U9286 ( .A1(SI_28_), .A2(keyinput_g4), .B1(keyinput_g62), .B2(
        P2_REG3_REG_26__SCAN_IN), .ZN(n7540) );
  AOI221_X1 U9287 ( .B1(SI_28_), .B2(keyinput_g4), .C1(P2_REG3_REG_26__SCAN_IN), .C2(keyinput_g62), .A(n7540), .ZN(n7543) );
  OAI22_X1 U9288 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_g42), .B1(
        keyinput_g2), .B2(SI_30_), .ZN(n7541) );
  AOI221_X1 U9289 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .C1(
        SI_30_), .C2(keyinput_g2), .A(n7541), .ZN(n7542) );
  NAND4_X1 U9290 ( .A1(n7545), .A2(n7544), .A3(n7543), .A4(n7542), .ZN(n7546)
         );
  NOR4_X1 U9291 ( .A1(n7549), .A2(n7548), .A3(n7547), .A4(n7546), .ZN(n7609)
         );
  AOI22_X1 U9292 ( .A1(n7551), .A2(keyinput_g18), .B1(keyinput_g53), .B2(n5694), .ZN(n7550) );
  OAI221_X1 U9293 ( .B1(n7551), .B2(keyinput_g18), .C1(n5694), .C2(
        keyinput_g53), .A(n7550), .ZN(n7562) );
  AOI22_X1 U9294 ( .A1(n7554), .A2(keyinput_g6), .B1(keyinput_g21), .B2(n7553), 
        .ZN(n7552) );
  OAI221_X1 U9295 ( .B1(n7554), .B2(keyinput_g6), .C1(n7553), .C2(keyinput_g21), .A(n7552), .ZN(n7561) );
  AOI22_X1 U9296 ( .A1(n8780), .A2(keyinput_g57), .B1(keyinput_g37), .B2(n7556), .ZN(n7555) );
  OAI221_X1 U9297 ( .B1(n8780), .B2(keyinput_g57), .C1(n7556), .C2(
        keyinput_g37), .A(n7555), .ZN(n7560) );
  INV_X1 U9298 ( .A(SI_6_), .ZN(n7558) );
  AOI22_X1 U9299 ( .A1(n5669), .A2(keyinput_g35), .B1(n7558), .B2(keyinput_g26), .ZN(n7557) );
  OAI221_X1 U9300 ( .B1(n5669), .B2(keyinput_g35), .C1(n7558), .C2(
        keyinput_g26), .A(n7557), .ZN(n7559) );
  NOR4_X1 U9301 ( .A1(n7562), .A2(n7561), .A3(n7560), .A4(n7559), .ZN(n7608)
         );
  AOI22_X1 U9302 ( .A1(n7564), .A2(keyinput_g7), .B1(keyinput_g56), .B2(n6781), 
        .ZN(n7563) );
  OAI221_X1 U9303 ( .B1(n7564), .B2(keyinput_g7), .C1(n6781), .C2(keyinput_g56), .A(n7563), .ZN(n7576) );
  AOI22_X1 U9304 ( .A1(n5758), .A2(keyinput_g63), .B1(n7566), .B2(keyinput_g48), .ZN(n7565) );
  OAI221_X1 U9305 ( .B1(n5758), .B2(keyinput_g63), .C1(n7566), .C2(
        keyinput_g48), .A(n7565), .ZN(n7575) );
  AOI22_X1 U9306 ( .A1(n7569), .A2(keyinput_g24), .B1(keyinput_g54), .B2(n7568), .ZN(n7567) );
  OAI221_X1 U9307 ( .B1(n7569), .B2(keyinput_g24), .C1(n7568), .C2(
        keyinput_g54), .A(n7567), .ZN(n7574) );
  AOI22_X1 U9308 ( .A1(n7572), .A2(keyinput_g61), .B1(keyinput_g52), .B2(n7571), .ZN(n7570) );
  OAI221_X1 U9309 ( .B1(n7572), .B2(keyinput_g61), .C1(n7571), .C2(
        keyinput_g52), .A(n7570), .ZN(n7573) );
  NOR4_X1 U9310 ( .A1(n7576), .A2(n7575), .A3(n7574), .A4(n7573), .ZN(n7606)
         );
  AOI22_X1 U9311 ( .A1(n7579), .A2(keyinput_g9), .B1(keyinput_g20), .B2(n7578), 
        .ZN(n7577) );
  OAI221_X1 U9312 ( .B1(n7579), .B2(keyinput_g9), .C1(n7578), .C2(keyinput_g20), .A(n7577), .ZN(n7587) );
  AOI22_X1 U9313 ( .A1(n7582), .A2(keyinput_g19), .B1(n7581), .B2(keyinput_g10), .ZN(n7580) );
  OAI221_X1 U9314 ( .B1(n7582), .B2(keyinput_g19), .C1(n7581), .C2(
        keyinput_g10), .A(n7580), .ZN(n7586) );
  XNOR2_X1 U9315 ( .A(SI_2_), .B(keyinput_g30), .ZN(n7584) );
  XNOR2_X1 U9316 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_g38), .ZN(n7583)
         );
  NAND2_X1 U9317 ( .A1(n7584), .A2(n7583), .ZN(n7585) );
  NOR3_X1 U9318 ( .A1(n7587), .A2(n7586), .A3(n7585), .ZN(n7605) );
  INV_X1 U9319 ( .A(P2_WR_REG_SCAN_IN), .ZN(n9875) );
  AOI22_X1 U9320 ( .A1(n9875), .A2(keyinput_g0), .B1(n7589), .B2(keyinput_g3), 
        .ZN(n7588) );
  OAI221_X1 U9321 ( .B1(n9875), .B2(keyinput_g0), .C1(n7589), .C2(keyinput_g3), 
        .A(n7588), .ZN(n7593) );
  AOI22_X1 U9322 ( .A1(n7591), .A2(keyinput_g8), .B1(keyinput_g39), .B2(n8271), 
        .ZN(n7590) );
  OAI221_X1 U9323 ( .B1(n7591), .B2(keyinput_g8), .C1(n8271), .C2(keyinput_g39), .A(n7590), .ZN(n7592) );
  NOR2_X1 U9324 ( .A1(n7593), .A2(n7592), .ZN(n7604) );
  INV_X1 U9325 ( .A(SI_7_), .ZN(n7595) );
  AOI22_X1 U9326 ( .A1(n7596), .A2(keyinput_g13), .B1(keyinput_g25), .B2(n7595), .ZN(n7594) );
  OAI221_X1 U9327 ( .B1(n7596), .B2(keyinput_g13), .C1(n7595), .C2(
        keyinput_g25), .A(n7594), .ZN(n7602) );
  XNOR2_X1 U9328 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_g45), .ZN(n7600)
         );
  XNOR2_X1 U9329 ( .A(SI_1_), .B(keyinput_g31), .ZN(n7599) );
  XNOR2_X1 U9330 ( .A(SI_5_), .B(keyinput_g27), .ZN(n7598) );
  XNOR2_X1 U9331 ( .A(SI_3_), .B(keyinput_g29), .ZN(n7597) );
  NAND4_X1 U9332 ( .A1(n7600), .A2(n7599), .A3(n7598), .A4(n7597), .ZN(n7601)
         );
  NOR2_X1 U9333 ( .A1(n7602), .A2(n7601), .ZN(n7603) );
  AND4_X1 U9334 ( .A1(n7606), .A2(n7605), .A3(n7604), .A4(n7603), .ZN(n7607)
         );
  NAND3_X1 U9335 ( .A1(n7609), .A2(n7608), .A3(n7607), .ZN(n7610) );
  NAND2_X1 U9336 ( .A1(n7611), .A2(n7610), .ZN(n7615) );
  NOR2_X1 U9337 ( .A1(n7613), .A2(n7612), .ZN(n7614) );
  XNOR2_X1 U9338 ( .A(n7615), .B(n7614), .ZN(n7616) );
  XNOR2_X1 U9339 ( .A(n7617), .B(n7616), .ZN(ADD_1071_U4) );
  INV_X1 U9340 ( .A(n7659), .ZN(n7619) );
  NAND2_X1 U9341 ( .A1(n9218), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7618) );
  OAI211_X1 U9342 ( .C1(n7619), .C2(n9221), .A(n8251), .B(n7618), .ZN(P2_U3335) );
  OAI21_X1 U9343 ( .B1(n7621), .B2(n8221), .A(n7620), .ZN(n9815) );
  XNOR2_X1 U9344 ( .A(n7622), .B(n8221), .ZN(n7625) );
  OAI22_X1 U9345 ( .A1(n7623), .A2(n9074), .B1(n7891), .B2(n9076), .ZN(n7624)
         );
  AOI21_X1 U9346 ( .B1(n7625), .B2(n10049), .A(n7624), .ZN(n7626) );
  OAI21_X1 U9347 ( .B1(n10039), .B2(n9815), .A(n7626), .ZN(n9818) );
  NAND2_X1 U9348 ( .A1(n9818), .A2(n9049), .ZN(n7634) );
  OR2_X1 U9349 ( .A1(n7627), .A2(n9816), .ZN(n7628) );
  NAND2_X1 U9350 ( .A1(n7723), .A2(n7628), .ZN(n9817) );
  INV_X1 U9351 ( .A(n9817), .ZN(n7632) );
  AOI22_X1 U9352 ( .A1(n10070), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7629), .B2(
        n10062), .ZN(n7630) );
  OAI21_X1 U9353 ( .B1(n9816), .B2(n10054), .A(n7630), .ZN(n7631) );
  AOI21_X1 U9354 ( .B1(n7632), .B2(n9088), .A(n7631), .ZN(n7633) );
  OAI211_X1 U9355 ( .C1(n9815), .C2(n10053), .A(n7634), .B(n7633), .ZN(
        P2_U3283) );
  NAND2_X1 U9356 ( .A1(n7799), .A2(n8714), .ZN(n7636) );
  OR2_X1 U9357 ( .A1(n7688), .A2(n6498), .ZN(n7635) );
  NAND2_X1 U9358 ( .A1(n7636), .A2(n7635), .ZN(n7637) );
  XNOR2_X1 U9359 ( .A(n7637), .B(n8689), .ZN(n7679) );
  NOR2_X1 U9360 ( .A1(n7688), .A2(n8719), .ZN(n7638) );
  AOI21_X1 U9361 ( .B1(n7799), .B2(n8706), .A(n7638), .ZN(n7678) );
  XNOR2_X1 U9362 ( .A(n7679), .B(n7678), .ZN(n7650) );
  OR2_X1 U9363 ( .A1(n7641), .A2(n4847), .ZN(n7644) );
  OR2_X1 U9364 ( .A1(n4847), .A2(n7642), .ZN(n7643) );
  OAI21_X2 U9365 ( .B1(n7645), .B2(n7644), .A(n7643), .ZN(n7647) );
  INV_X1 U9366 ( .A(n7650), .ZN(n7646) );
  NAND2_X1 U9367 ( .A1(n7647), .A2(n7646), .ZN(n7681) );
  INV_X1 U9368 ( .A(n7681), .ZN(n7648) );
  AOI21_X1 U9369 ( .B1(n7650), .B2(n7649), .A(n7648), .ZN(n7658) );
  INV_X1 U9370 ( .A(n7790), .ZN(n7656) );
  NAND2_X1 U9371 ( .A1(n9855), .A2(n9302), .ZN(n7652) );
  OAI211_X1 U9372 ( .C1(n7778), .C2(n9304), .A(n7652), .B(n7651), .ZN(n7655)
         );
  NAND2_X1 U9373 ( .A1(n7799), .A2(n9969), .ZN(n9856) );
  NOR2_X1 U9374 ( .A1(n9856), .A2(n7653), .ZN(n7654) );
  AOI211_X1 U9375 ( .C1(n7656), .C2(n9306), .A(n7655), .B(n7654), .ZN(n7657)
         );
  OAI21_X1 U9376 ( .B1(n7658), .B2(n9315), .A(n7657), .ZN(P1_U3222) );
  NAND2_X1 U9377 ( .A1(n7659), .A2(n8013), .ZN(n7661) );
  NOR2_X1 U9378 ( .A1(n7660), .A2(P1_U3084), .ZN(n8584) );
  INV_X1 U9379 ( .A(n8584), .ZN(n8590) );
  OAI211_X1 U9380 ( .C1(n7662), .C2(n9771), .A(n7661), .B(n8590), .ZN(P1_U3330) );
  NOR2_X1 U9381 ( .A1(n7663), .A2(n7668), .ZN(n7664) );
  NAND2_X1 U9382 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9355), .ZN(n7665) );
  OAI21_X1 U9383 ( .B1(n9355), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7665), .ZN(
        n7666) );
  AOI211_X1 U9384 ( .C1(n4381), .C2(n7666), .A(n9354), .B(n9895), .ZN(n7677)
         );
  NOR2_X1 U9385 ( .A1(n7668), .A2(n7667), .ZN(n7670) );
  NOR2_X1 U9386 ( .A1(n7670), .A2(n7669), .ZN(n7672) );
  XNOR2_X1 U9387 ( .A(n9355), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7671) );
  NOR2_X1 U9388 ( .A1(n7672), .A2(n7671), .ZN(n9347) );
  AOI211_X1 U9389 ( .C1(n7672), .C2(n7671), .A(n9347), .B(n9876), .ZN(n7676)
         );
  NAND2_X1 U9390 ( .A1(n9882), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7673) );
  NAND2_X1 U9391 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7835) );
  OAI211_X1 U9392 ( .C1(n9914), .C2(n7674), .A(n7673), .B(n7835), .ZN(n7675)
         );
  OR3_X1 U9393 ( .A1(n7677), .A2(n7676), .A3(n7675), .ZN(P1_U3257) );
  NAND2_X1 U9394 ( .A1(n7679), .A2(n7678), .ZN(n7680) );
  NAND2_X1 U9395 ( .A1(n7859), .A2(n8714), .ZN(n7683) );
  NAND2_X1 U9396 ( .A1(n9854), .A2(n8716), .ZN(n7682) );
  NAND2_X1 U9397 ( .A1(n7683), .A2(n7682), .ZN(n7684) );
  XNOR2_X1 U9398 ( .A(n7684), .B(n8689), .ZN(n7749) );
  AND2_X1 U9399 ( .A1(n9854), .A2(n6414), .ZN(n7685) );
  AOI21_X1 U9400 ( .B1(n7859), .B2(n8706), .A(n7685), .ZN(n7750) );
  XNOR2_X1 U9401 ( .A(n7749), .B(n7750), .ZN(n7686) );
  XNOR2_X1 U9402 ( .A(n7815), .B(n7686), .ZN(n7693) );
  OAI21_X1 U9403 ( .B1(n9272), .B2(n7688), .A(n7687), .ZN(n7689) );
  AOI21_X1 U9404 ( .B1(n9311), .B2(n9615), .A(n7689), .ZN(n7690) );
  OAI21_X1 U9405 ( .B1(n9262), .B2(n7851), .A(n7690), .ZN(n7691) );
  AOI21_X1 U9406 ( .B1(n7859), .B2(n9320), .A(n7691), .ZN(n7692) );
  OAI21_X1 U9407 ( .B1(n7693), .B2(n9315), .A(n7692), .ZN(P1_U3232) );
  XNOR2_X1 U9408 ( .A(n9191), .B(n8606), .ZN(n7694) );
  NAND2_X1 U9409 ( .A1(n8818), .A2(n8630), .ZN(n7695) );
  NAND2_X1 U9410 ( .A1(n7694), .A2(n7695), .ZN(n7732) );
  INV_X1 U9411 ( .A(n7694), .ZN(n7697) );
  INV_X1 U9412 ( .A(n7695), .ZN(n7696) );
  NAND2_X1 U9413 ( .A1(n7697), .A2(n7696), .ZN(n7698) );
  NAND2_X1 U9414 ( .A1(n7732), .A2(n7698), .ZN(n7710) );
  NAND2_X1 U9415 ( .A1(n7700), .A2(n7699), .ZN(n7705) );
  INV_X1 U9416 ( .A(n7701), .ZN(n7703) );
  NAND2_X1 U9417 ( .A1(n7703), .A2(n7702), .ZN(n7704) );
  NAND2_X1 U9418 ( .A1(n7705), .A2(n7704), .ZN(n7709) );
  INV_X1 U9419 ( .A(n7709), .ZN(n7707) );
  INV_X1 U9420 ( .A(n7710), .ZN(n7706) );
  NAND2_X2 U9421 ( .A1(n7707), .A2(n7706), .ZN(n7733) );
  INV_X1 U9422 ( .A(n7733), .ZN(n7708) );
  AOI21_X1 U9423 ( .B1(n7710), .B2(n7709), .A(n7708), .ZN(n7714) );
  NAND2_X1 U9424 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8892) );
  OAI21_X1 U9425 ( .B1(n8781), .B2(n7907), .A(n8892), .ZN(n7712) );
  OAI22_X1 U9426 ( .A1(n8805), .A2(n7906), .B1(n7912), .B2(n10026), .ZN(n7711)
         );
  AOI211_X1 U9427 ( .C1(n9191), .C2(n8809), .A(n7712), .B(n7711), .ZN(n7713)
         );
  OAI21_X1 U9428 ( .B1(n7714), .B2(n8812), .A(n7713), .ZN(P2_U3228) );
  AOI21_X1 U9429 ( .B1(n8224), .B2(n7716), .A(n7715), .ZN(n9807) );
  AOI211_X1 U9430 ( .C1(n7719), .C2(n7718), .A(n9071), .B(n7717), .ZN(n7722)
         );
  OAI22_X1 U9431 ( .A1(n7906), .A2(n9076), .B1(n7720), .B2(n9074), .ZN(n7721)
         );
  OR2_X1 U9432 ( .A1(n7722), .A2(n7721), .ZN(n9810) );
  INV_X1 U9433 ( .A(n7723), .ZN(n7725) );
  OAI21_X1 U9434 ( .B1(n7725), .B2(n9808), .A(n4500), .ZN(n9809) );
  AOI22_X1 U9435 ( .A1(n10070), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7726), .B2(
        n10062), .ZN(n7729) );
  NAND2_X1 U9436 ( .A1(n7727), .A2(n8926), .ZN(n7728) );
  OAI211_X1 U9437 ( .C1(n9809), .C2(n8935), .A(n7729), .B(n7728), .ZN(n7730)
         );
  AOI21_X1 U9438 ( .B1(n9810), .B2(n9049), .A(n7730), .ZN(n7731) );
  OAI21_X1 U9439 ( .B1(n9807), .B2(n9126), .A(n7731), .ZN(P2_U3282) );
  XNOR2_X1 U9440 ( .A(n9188), .B(n8606), .ZN(n7803) );
  NAND2_X1 U9441 ( .A1(n9119), .A2(n8630), .ZN(n7802) );
  XNOR2_X1 U9442 ( .A(n7803), .B(n7802), .ZN(n7804) );
  XNOR2_X1 U9443 ( .A(n7805), .B(n7804), .ZN(n7737) );
  OAI22_X1 U9444 ( .A1(n8781), .A2(n7956), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8262), .ZN(n7735) );
  OAI22_X1 U9445 ( .A1(n8805), .A2(n7955), .B1(n7960), .B2(n10026), .ZN(n7734)
         );
  AOI211_X1 U9446 ( .C1(n9188), .C2(n8809), .A(n7735), .B(n7734), .ZN(n7736)
         );
  OAI21_X1 U9447 ( .B1(n7737), .B2(n8812), .A(n7736), .ZN(P2_U3230) );
  INV_X1 U9448 ( .A(n7738), .ZN(n7742) );
  OAI222_X1 U9449 ( .A1(n9781), .A2(n7742), .B1(P1_U3084), .B2(n7740), .C1(
        n7739), .C2(n9777), .ZN(P1_U3329) );
  OAI222_X1 U9450 ( .A1(P2_U3152), .A2(n7743), .B1(n9221), .B2(n7742), .C1(
        n7741), .C2(n8019), .ZN(P2_U3334) );
  AND2_X1 U9451 ( .A1(n7749), .A2(n7750), .ZN(n7813) );
  NAND2_X1 U9452 ( .A1(n7932), .A2(n8714), .ZN(n7745) );
  NAND2_X1 U9453 ( .A1(n9615), .A2(n8716), .ZN(n7744) );
  NAND2_X1 U9454 ( .A1(n7745), .A2(n7744), .ZN(n7746) );
  XNOR2_X1 U9455 ( .A(n7746), .B(n8689), .ZN(n7774) );
  AND2_X1 U9456 ( .A1(n9615), .A2(n6414), .ZN(n7747) );
  AOI21_X1 U9457 ( .B1(n7932), .B2(n8706), .A(n7747), .ZN(n7753) );
  NAND2_X1 U9458 ( .A1(n7774), .A2(n7753), .ZN(n7811) );
  INV_X1 U9459 ( .A(n7811), .ZN(n7756) );
  OR2_X1 U9460 ( .A1(n7813), .A2(n7756), .ZN(n7748) );
  OR2_X1 U9461 ( .A1(n7815), .A2(n7748), .ZN(n7758) );
  INV_X1 U9462 ( .A(n7749), .ZN(n7752) );
  INV_X1 U9463 ( .A(n7750), .ZN(n7751) );
  NAND2_X1 U9464 ( .A1(n7752), .A2(n7751), .ZN(n7771) );
  INV_X1 U9465 ( .A(n7774), .ZN(n7754) );
  INV_X1 U9466 ( .A(n7753), .ZN(n7773) );
  NAND2_X1 U9467 ( .A1(n7754), .A2(n7773), .ZN(n7755) );
  AND2_X1 U9468 ( .A1(n7771), .A2(n7755), .ZN(n7816) );
  OR2_X1 U9469 ( .A1(n7756), .A2(n7816), .ZN(n7757) );
  NAND2_X1 U9470 ( .A1(n7758), .A2(n7757), .ZN(n7764) );
  NAND2_X1 U9471 ( .A1(n9624), .A2(n8714), .ZN(n7760) );
  NAND2_X1 U9472 ( .A1(n9324), .A2(n8716), .ZN(n7759) );
  NAND2_X1 U9473 ( .A1(n7760), .A2(n7759), .ZN(n7761) );
  XNOR2_X1 U9474 ( .A(n7761), .B(n8689), .ZN(n7818) );
  AND2_X1 U9475 ( .A1(n9324), .A2(n6414), .ZN(n7762) );
  AOI21_X1 U9476 ( .B1(n9624), .B2(n8706), .A(n7762), .ZN(n7810) );
  INV_X1 U9477 ( .A(n7810), .ZN(n7819) );
  XNOR2_X1 U9478 ( .A(n7818), .B(n7819), .ZN(n7763) );
  XNOR2_X1 U9479 ( .A(n7764), .B(n7763), .ZN(n7770) );
  OAI21_X1 U9480 ( .B1(n9586), .B2(n9304), .A(n7765), .ZN(n7766) );
  AOI21_X1 U9481 ( .B1(n9302), .B2(n9615), .A(n7766), .ZN(n7767) );
  OAI21_X1 U9482 ( .B1(n9262), .B2(n9625), .A(n7767), .ZN(n7768) );
  AOI21_X1 U9483 ( .B1(n9624), .B2(n9320), .A(n7768), .ZN(n7769) );
  OAI21_X1 U9484 ( .B1(n7770), .B2(n9315), .A(n7769), .ZN(P1_U3239) );
  OR2_X1 U9485 ( .A1(n7815), .A2(n7813), .ZN(n7772) );
  NAND2_X1 U9486 ( .A1(n7772), .A2(n7771), .ZN(n7776) );
  XNOR2_X1 U9487 ( .A(n7774), .B(n7773), .ZN(n7775) );
  XNOR2_X1 U9488 ( .A(n7776), .B(n7775), .ZN(n7783) );
  OAI21_X1 U9489 ( .B1(n9272), .B2(n7778), .A(n7777), .ZN(n7779) );
  AOI21_X1 U9490 ( .B1(n9311), .B2(n9324), .A(n7779), .ZN(n7780) );
  OAI21_X1 U9491 ( .B1(n9282), .B2(n7933), .A(n7780), .ZN(n7781) );
  AOI21_X1 U9492 ( .B1(n7932), .B2(n9320), .A(n7781), .ZN(n7782) );
  OAI21_X1 U9493 ( .B1(n7783), .B2(n9315), .A(n7782), .ZN(P1_U3213) );
  NAND2_X1 U9494 ( .A1(n7785), .A2(n7784), .ZN(n7786) );
  XNOR2_X1 U9495 ( .A(n7786), .B(n8426), .ZN(n7787) );
  NAND2_X1 U9496 ( .A1(n7787), .A2(n9693), .ZN(n9859) );
  OAI21_X1 U9497 ( .B1(n7789), .B2(n8426), .A(n7788), .ZN(n9862) );
  INV_X1 U9498 ( .A(n9862), .ZN(n9865) );
  NAND2_X1 U9499 ( .A1(n9865), .A2(n9595), .ZN(n7801) );
  INV_X1 U9500 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7791) );
  OAI22_X1 U9501 ( .A1(n9601), .A2(n7791), .B1(n7790), .B2(n9598), .ZN(n7792)
         );
  AOI21_X1 U9502 ( .B1(n9605), .B2(n9854), .A(n7792), .ZN(n7793) );
  OAI21_X1 U9503 ( .B1(n7794), .B2(n9597), .A(n7793), .ZN(n7798) );
  OAI21_X1 U9504 ( .B1(n9846), .B2(n7795), .A(n9847), .ZN(n7796) );
  OR2_X1 U9505 ( .A1(n7796), .A2(n7856), .ZN(n9857) );
  NOR2_X1 U9506 ( .A1(n9857), .A2(n9530), .ZN(n7797) );
  AOI211_X1 U9507 ( .C1(n9844), .C2(n7799), .A(n7798), .B(n7797), .ZN(n7800)
         );
  OAI211_X1 U9508 ( .C1(n9939), .C2(n9859), .A(n7801), .B(n7800), .ZN(P1_U3279) );
  XNOR2_X1 U9509 ( .A(n9182), .B(n8631), .ZN(n7974) );
  NAND2_X1 U9510 ( .A1(n8817), .A2(n10133), .ZN(n7972) );
  XNOR2_X1 U9511 ( .A(n7974), .B(n7972), .ZN(n7970) );
  XNOR2_X1 U9512 ( .A(n7971), .B(n7970), .ZN(n7809) );
  NAND2_X1 U9513 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7881) );
  OAI21_X1 U9514 ( .B1(n8781), .B2(n9075), .A(n7881), .ZN(n7807) );
  OAI22_X1 U9515 ( .A1(n8805), .A2(n7907), .B1(n9112), .B2(n10026), .ZN(n7806)
         );
  AOI211_X1 U9516 ( .C1(n9182), .C2(n8809), .A(n7807), .B(n7806), .ZN(n7808)
         );
  OAI21_X1 U9517 ( .B1(n7809), .B2(n8812), .A(n7808), .ZN(P2_U3240) );
  NAND2_X1 U9518 ( .A1(n7818), .A2(n7810), .ZN(n7812) );
  NAND2_X1 U9519 ( .A1(n7812), .A2(n7811), .ZN(n7817) );
  OR2_X1 U9520 ( .A1(n7813), .A2(n7817), .ZN(n7814) );
  OR2_X1 U9521 ( .A1(n7817), .A2(n7816), .ZN(n7822) );
  INV_X1 U9522 ( .A(n7818), .ZN(n7820) );
  NAND2_X1 U9523 ( .A1(n7820), .A2(n7819), .ZN(n7821) );
  AND2_X1 U9524 ( .A1(n7822), .A2(n7821), .ZN(n7823) );
  NAND2_X1 U9525 ( .A1(n9715), .A2(n8714), .ZN(n7825) );
  NAND2_X1 U9526 ( .A1(n9616), .A2(n8716), .ZN(n7824) );
  NAND2_X1 U9527 ( .A1(n7825), .A2(n7824), .ZN(n7826) );
  XNOR2_X1 U9528 ( .A(n7826), .B(n8721), .ZN(n7832) );
  INV_X1 U9529 ( .A(n7832), .ZN(n7830) );
  NAND2_X1 U9530 ( .A1(n9715), .A2(n8716), .ZN(n7828) );
  NAND2_X1 U9531 ( .A1(n9616), .A2(n6414), .ZN(n7827) );
  NAND2_X1 U9532 ( .A1(n7828), .A2(n7827), .ZN(n7831) );
  INV_X1 U9533 ( .A(n7831), .ZN(n7829) );
  NAND2_X1 U9534 ( .A1(n7830), .A2(n7829), .ZN(n7990) );
  INV_X1 U9535 ( .A(n7990), .ZN(n7833) );
  AND2_X1 U9536 ( .A1(n7832), .A2(n7831), .ZN(n7991) );
  NOR2_X1 U9537 ( .A1(n7833), .A2(n7991), .ZN(n7834) );
  XNOR2_X1 U9538 ( .A(n7992), .B(n7834), .ZN(n7840) );
  OAI21_X1 U9539 ( .B1(n9712), .B2(n9304), .A(n7835), .ZN(n7836) );
  AOI21_X1 U9540 ( .B1(n9310), .B2(n9324), .A(n7836), .ZN(n7837) );
  OAI21_X1 U9541 ( .B1(n9262), .B2(n9599), .A(n7837), .ZN(n7838) );
  AOI21_X1 U9542 ( .B1(n9715), .B2(n9320), .A(n7838), .ZN(n7839) );
  OAI21_X1 U9543 ( .B1(n7840), .B2(n9315), .A(n7839), .ZN(P1_U3224) );
  INV_X1 U9544 ( .A(n7841), .ZN(n7845) );
  OAI222_X1 U9545 ( .A1(n8019), .A2(n7843), .B1(n9221), .B2(n7845), .C1(
        P2_U3152), .C2(n7842), .ZN(P2_U3333) );
  OAI222_X1 U9546 ( .A1(n9777), .A2(n7847), .B1(n7846), .B2(n7845), .C1(n7844), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  OAI21_X1 U9547 ( .B1(n7848), .B2(n8443), .A(n7926), .ZN(n7849) );
  INV_X1 U9548 ( .A(n7849), .ZN(n7946) );
  XNOR2_X1 U9549 ( .A(n7850), .B(n8443), .ZN(n7948) );
  NAND2_X1 U9550 ( .A1(n7948), .A2(n9595), .ZN(n7861) );
  NAND2_X1 U9551 ( .A1(n9525), .A2(n9838), .ZN(n7854) );
  INV_X1 U9552 ( .A(n7851), .ZN(n7852) );
  AOI22_X1 U9553 ( .A1(n9939), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7852), .B2(
        n9936), .ZN(n7853) );
  OAI211_X1 U9554 ( .C1(n7855), .C2(n9527), .A(n7854), .B(n7853), .ZN(n7858)
         );
  OAI211_X1 U9555 ( .C1(n7856), .C2(n7952), .A(n9847), .B(n4388), .ZN(n7944)
         );
  NOR2_X1 U9556 ( .A1(n7944), .A2(n9530), .ZN(n7857) );
  AOI211_X1 U9557 ( .C1(n9844), .C2(n7859), .A(n7858), .B(n7857), .ZN(n7860)
         );
  OAI211_X1 U9558 ( .C1(n7946), .C2(n9611), .A(n7861), .B(n7860), .ZN(P1_U3278) );
  NAND2_X1 U9559 ( .A1(n7876), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7870) );
  INV_X1 U9560 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7961) );
  XNOR2_X1 U9561 ( .A(n7876), .B(n7961), .ZN(n8260) );
  NAND2_X1 U9562 ( .A1(n8895), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7869) );
  INV_X1 U9563 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7864) );
  INV_X1 U9564 ( .A(n7869), .ZN(n7862) );
  AOI21_X1 U9565 ( .B1(n7864), .B2(n7863), .A(n7862), .ZN(n8898) );
  NOR2_X1 U9566 ( .A1(n7866), .A2(n7865), .ZN(n7868) );
  NOR2_X1 U9567 ( .A1(n7868), .A2(n7867), .ZN(n8899) );
  NAND2_X1 U9568 ( .A1(n8898), .A2(n8899), .ZN(n8897) );
  NAND2_X1 U9569 ( .A1(n7869), .A2(n8897), .ZN(n8261) );
  NAND2_X1 U9570 ( .A1(n8260), .A2(n8261), .ZN(n8259) );
  NAND2_X1 U9571 ( .A1(n7870), .A2(n8259), .ZN(n8906) );
  XNOR2_X1 U9572 ( .A(n8907), .B(n8906), .ZN(n7871) );
  NOR2_X1 U9573 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n7871), .ZN(n8908) );
  AOI21_X1 U9574 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n7871), .A(n8908), .ZN(
        n7887) );
  XNOR2_X1 U9575 ( .A(n7876), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8264) );
  XOR2_X1 U9576 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8895), .Z(n8889) );
  NOR2_X1 U9577 ( .A1(n7873), .A2(n7872), .ZN(n7875) );
  AOI21_X1 U9578 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n7876), .A(n8263), .ZN(
        n7879) );
  INV_X1 U9579 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7877) );
  AOI22_X1 U9580 ( .A1(n8907), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n7877), .B2(
        n7882), .ZN(n7878) );
  NAND2_X1 U9581 ( .A1(n7879), .A2(n7878), .ZN(n8903) );
  OAI21_X1 U9582 ( .B1(n7879), .B2(n7878), .A(n8903), .ZN(n7884) );
  NAND2_X1 U9583 ( .A1(n10034), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n7880) );
  OAI211_X1 U9584 ( .C1(n10030), .C2(n7882), .A(n7881), .B(n7880), .ZN(n7883)
         );
  AOI21_X1 U9585 ( .B1(n7884), .B2(n10027), .A(n7883), .ZN(n7885) );
  OAI21_X1 U9586 ( .B1(n7887), .B2(n7886), .A(n7885), .ZN(P2_U3263) );
  XNOR2_X1 U9587 ( .A(n7888), .B(n8223), .ZN(n9805) );
  INV_X1 U9588 ( .A(n9805), .ZN(n7900) );
  AOI211_X1 U9589 ( .C1(n7890), .C2(n4814), .A(n9071), .B(n7889), .ZN(n7893)
         );
  OAI22_X1 U9590 ( .A1(n7955), .A2(n9076), .B1(n7891), .B2(n9074), .ZN(n7892)
         );
  OR2_X1 U9591 ( .A1(n7893), .A2(n7892), .ZN(n9803) );
  OAI21_X1 U9592 ( .B1(n7724), .B2(n5978), .A(n7910), .ZN(n9802) );
  AOI22_X1 U9593 ( .A1(n10070), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7894), .B2(
        n10062), .ZN(n7897) );
  NAND2_X1 U9594 ( .A1(n7895), .A2(n8926), .ZN(n7896) );
  OAI211_X1 U9595 ( .C1(n9802), .C2(n8935), .A(n7897), .B(n7896), .ZN(n7898)
         );
  AOI21_X1 U9596 ( .B1(n9803), .B2(n9049), .A(n7898), .ZN(n7899) );
  OAI21_X1 U9597 ( .B1(n7900), .B2(n9126), .A(n7899), .ZN(P2_U3281) );
  INV_X1 U9598 ( .A(n7901), .ZN(n7919) );
  OAI222_X1 U9599 ( .A1(n9781), .A2(n7919), .B1(P1_U3084), .B2(n7903), .C1(
        n7902), .C2(n9777), .ZN(P1_U3327) );
  XOR2_X1 U9600 ( .A(n8225), .B(n7904), .Z(n7905) );
  OAI222_X1 U9601 ( .A1(n9076), .A2(n7907), .B1(n9074), .B2(n7906), .C1(n9071), 
        .C2(n7905), .ZN(n9193) );
  INV_X1 U9602 ( .A(n9193), .ZN(n7917) );
  AOI21_X1 U9603 ( .B1(n8225), .B2(n7909), .A(n7908), .ZN(n9195) );
  AND2_X1 U9604 ( .A1(n7910), .A2(n9191), .ZN(n7911) );
  OR2_X1 U9605 ( .A1(n7911), .A2(n7964), .ZN(n9192) );
  OAI22_X1 U9606 ( .A1(n9049), .A2(n7864), .B1(n7912), .B2(n8975), .ZN(n7913)
         );
  AOI21_X1 U9607 ( .B1(n9191), .B2(n8926), .A(n7913), .ZN(n7914) );
  OAI21_X1 U9608 ( .B1(n9192), .B2(n8935), .A(n7914), .ZN(n7915) );
  AOI21_X1 U9609 ( .B1(n9195), .B2(n9082), .A(n7915), .ZN(n7916) );
  OAI21_X1 U9610 ( .B1(n7917), .B2(n10070), .A(n7916), .ZN(P2_U3280) );
  OAI222_X1 U9611 ( .A1(P2_U3152), .A2(n7920), .B1(n9221), .B2(n7919), .C1(
        n7918), .C2(n8019), .ZN(P2_U3332) );
  INV_X1 U9612 ( .A(n7940), .ZN(n7923) );
  AOI22_X1 U9613 ( .A1(n7921), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n9218), .ZN(n7922) );
  OAI21_X1 U9614 ( .B1(n7923), .B2(n9221), .A(n7922), .ZN(P2_U3331) );
  NAND2_X1 U9615 ( .A1(n7924), .A2(n9693), .ZN(n7929) );
  INV_X1 U9616 ( .A(n8445), .ZN(n7925) );
  AOI21_X1 U9617 ( .B1(n7926), .B2(n8336), .A(n7925), .ZN(n7928) );
  AOI22_X1 U9618 ( .A1(n9985), .A2(n9854), .B1(n9324), .B2(n5499), .ZN(n7927)
         );
  OAI21_X1 U9619 ( .B1(n7929), .B2(n7928), .A(n7927), .ZN(n9724) );
  INV_X1 U9620 ( .A(n9724), .ZN(n7939) );
  XOR2_X1 U9621 ( .A(n8445), .B(n7930), .Z(n9726) );
  NAND2_X1 U9622 ( .A1(n9726), .A2(n9595), .ZN(n7938) );
  INV_X1 U9623 ( .A(n9623), .ZN(n7931) );
  AOI211_X1 U9624 ( .C1(n7932), .C2(n4388), .A(n9622), .B(n7931), .ZN(n9725)
         );
  INV_X1 U9625 ( .A(n7932), .ZN(n9768) );
  NOR2_X1 U9626 ( .A1(n9768), .A2(n9628), .ZN(n7936) );
  OAI22_X1 U9627 ( .A1(n9601), .A2(n7934), .B1(n7933), .B2(n9598), .ZN(n7935)
         );
  AOI211_X1 U9628 ( .C1(n9725), .C2(n9850), .A(n7936), .B(n7935), .ZN(n7937)
         );
  OAI211_X1 U9629 ( .C1(n9939), .C2(n7939), .A(n7938), .B(n7937), .ZN(P1_U3277) );
  NAND2_X1 U9630 ( .A1(n7940), .A2(n8013), .ZN(n7942) );
  OAI211_X1 U9631 ( .C1(n9771), .C2(n7943), .A(n7942), .B(n7941), .ZN(P1_U3326) );
  AOI22_X1 U9632 ( .A1(n9838), .A2(n9985), .B1(n5499), .B2(n9615), .ZN(n7945)
         );
  OAI211_X1 U9633 ( .C1(n7946), .C2(n9972), .A(n7945), .B(n7944), .ZN(n7947)
         );
  AOI21_X1 U9634 ( .B1(n7948), .B2(n9992), .A(n7947), .ZN(n7950) );
  MUX2_X1 U9635 ( .A(n5126), .B(n7950), .S(n9995), .Z(n7949) );
  OAI21_X1 U9636 ( .B1(n7952), .B2(n9767), .A(n7949), .ZN(P1_U3493) );
  MUX2_X1 U9637 ( .A(n5122), .B(n7950), .S(n10007), .Z(n7951) );
  OAI21_X1 U9638 ( .B1(n7952), .B2(n9728), .A(n7951), .ZN(P1_U3536) );
  XNOR2_X1 U9639 ( .A(n7953), .B(n8154), .ZN(n7954) );
  OAI222_X1 U9640 ( .A1(n9076), .A2(n7956), .B1(n9074), .B2(n7955), .C1(n7954), 
        .C2(n9071), .ZN(n9186) );
  OAI21_X1 U9641 ( .B1(n7958), .B2(n8228), .A(n7957), .ZN(n7959) );
  INV_X1 U9642 ( .A(n7959), .ZN(n9190) );
  OAI22_X1 U9643 ( .A1(n9049), .A2(n7961), .B1(n7960), .B2(n8975), .ZN(n7962)
         );
  AOI21_X1 U9644 ( .B1(n9188), .B2(n8926), .A(n7962), .ZN(n7967) );
  OAI21_X1 U9645 ( .B1(n7964), .B2(n7963), .A(n5952), .ZN(n7965) );
  NOR2_X1 U9646 ( .A1(n7965), .A2(n9109), .ZN(n9187) );
  NAND2_X1 U9647 ( .A1(n9187), .A2(n9124), .ZN(n7966) );
  OAI211_X1 U9648 ( .C1(n9190), .C2(n9126), .A(n7967), .B(n7966), .ZN(n7968)
         );
  AOI21_X1 U9649 ( .B1(n9049), .B2(n9186), .A(n7968), .ZN(n7969) );
  INV_X1 U9650 ( .A(n7969), .ZN(P2_U3279) );
  INV_X1 U9651 ( .A(n7972), .ZN(n7973) );
  XNOR2_X1 U9652 ( .A(n9177), .B(n8606), .ZN(n7975) );
  NAND2_X1 U9653 ( .A1(n9120), .A2(n8630), .ZN(n7976) );
  NAND2_X1 U9654 ( .A1(n7975), .A2(n7976), .ZN(n8002) );
  INV_X1 U9655 ( .A(n7975), .ZN(n7978) );
  INV_X1 U9656 ( .A(n7976), .ZN(n7977) );
  NAND2_X1 U9657 ( .A1(n7978), .A2(n7977), .ZN(n7979) );
  NAND2_X1 U9658 ( .A1(n8002), .A2(n7979), .ZN(n7983) );
  INV_X1 U9659 ( .A(n7984), .ZN(n7981) );
  INV_X1 U9660 ( .A(n7983), .ZN(n7980) );
  NAND2_X2 U9661 ( .A1(n7981), .A2(n7980), .ZN(n8003) );
  INV_X1 U9662 ( .A(n8003), .ZN(n7982) );
  AOI21_X1 U9663 ( .B1(n7984), .B2(n7983), .A(n7982), .ZN(n7989) );
  NOR2_X1 U9664 ( .A1(n10026), .A2(n9096), .ZN(n7987) );
  AND2_X1 U9665 ( .A1(n8817), .A2(n10045), .ZN(n7985) );
  AOI21_X1 U9666 ( .B1(n9062), .B2(n10046), .A(n7985), .ZN(n9102) );
  NAND2_X1 U9667 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8919) );
  OAI21_X1 U9668 ( .B1(n8637), .B2(n9102), .A(n8919), .ZN(n7986) );
  AOI211_X1 U9669 ( .C1(n9177), .C2(n8809), .A(n7987), .B(n7986), .ZN(n7988)
         );
  OAI21_X1 U9670 ( .B1(n7989), .B2(n8812), .A(n7988), .ZN(P2_U3221) );
  NAND2_X1 U9671 ( .A1(n9706), .A2(n8714), .ZN(n7994) );
  NAND2_X1 U9672 ( .A1(n9604), .A2(n8716), .ZN(n7993) );
  NAND2_X1 U9673 ( .A1(n7994), .A2(n7993), .ZN(n7995) );
  XNOR2_X1 U9674 ( .A(n7995), .B(n8721), .ZN(n8647) );
  AND2_X1 U9675 ( .A1(n9604), .A2(n6414), .ZN(n7996) );
  AOI21_X1 U9676 ( .B1(n9706), .B2(n8706), .A(n7996), .ZN(n8648) );
  XNOR2_X1 U9677 ( .A(n8647), .B(n8648), .ZN(n8645) );
  XOR2_X1 U9678 ( .A(n8646), .B(n8645), .Z(n8001) );
  NAND2_X1 U9679 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9352) );
  OAI21_X1 U9680 ( .B1(n9690), .B2(n9304), .A(n9352), .ZN(n7997) );
  AOI21_X1 U9681 ( .B1(n9310), .B2(n9616), .A(n7997), .ZN(n7998) );
  OAI21_X1 U9682 ( .B1(n9262), .B2(n9579), .A(n7998), .ZN(n7999) );
  AOI21_X1 U9683 ( .B1(n9706), .B2(n9320), .A(n7999), .ZN(n8000) );
  OAI21_X1 U9684 ( .B1(n8001), .B2(n9315), .A(n8000), .ZN(P1_U3226) );
  XNOR2_X1 U9685 ( .A(n9171), .B(n8606), .ZN(n8596) );
  NAND2_X1 U9686 ( .A1(n9062), .A2(n8630), .ZN(n8597) );
  XNOR2_X1 U9687 ( .A(n8596), .B(n8597), .ZN(n8601) );
  XNOR2_X1 U9688 ( .A(n8602), .B(n8601), .ZN(n8009) );
  OAI22_X1 U9689 ( .A1(n8781), .A2(n9077), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8004), .ZN(n8007) );
  INV_X1 U9690 ( .A(n9084), .ZN(n8005) );
  OAI22_X1 U9691 ( .A1(n8805), .A2(n9075), .B1(n8005), .B2(n10026), .ZN(n8006)
         );
  AOI211_X1 U9692 ( .C1(n9171), .C2(n8809), .A(n8007), .B(n8006), .ZN(n8008)
         );
  OAI21_X1 U9693 ( .B1(n8009), .B2(n8812), .A(n8008), .ZN(P2_U3235) );
  INV_X1 U9694 ( .A(n5880), .ZN(n8012) );
  AOI22_X1 U9695 ( .A1(n8010), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n9218), .ZN(n8011) );
  OAI21_X1 U9696 ( .B1(n8012), .B2(n9221), .A(n8011), .ZN(P2_U3330) );
  NAND2_X1 U9697 ( .A1(n5880), .A2(n8013), .ZN(n8015) );
  OAI211_X1 U9698 ( .C1(n9771), .C2(n8016), .A(n8015), .B(n8014), .ZN(P1_U3325) );
  OAI222_X1 U9699 ( .A1(n8019), .A2(n8018), .B1(n9221), .B2(n8017), .C1(
        P2_U3152), .C2(n5953), .ZN(P2_U3336) );
  NAND2_X1 U9700 ( .A1(n8020), .A2(n9595), .ZN(n8028) );
  INV_X1 U9701 ( .A(n8021), .ZN(n8022) );
  AOI22_X1 U9702 ( .A1(n9939), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n8022), .B2(
        n9936), .ZN(n8023) );
  OAI21_X1 U9703 ( .B1(n9597), .B2(n9228), .A(n8023), .ZN(n8026) );
  NOR2_X1 U9704 ( .A1(n8024), .A2(n9530), .ZN(n8025) );
  AOI211_X1 U9705 ( .C1(n9844), .C2(n8409), .A(n8026), .B(n8025), .ZN(n8027)
         );
  OAI211_X1 U9706 ( .C1(n8029), .C2(n9939), .A(n8028), .B(n8027), .ZN(P1_U3355) );
  NOR2_X1 U9707 ( .A1(n8924), .A2(n8242), .ZN(n8032) );
  NAND2_X1 U9708 ( .A1(n8732), .A2(n8047), .ZN(n8031) );
  NAND2_X1 U9709 ( .A1(n5630), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8030) );
  AOI21_X1 U9710 ( .B1(n8032), .B2(n9800), .A(n8186), .ZN(n8034) );
  INV_X1 U9711 ( .A(n8814), .ZN(n8050) );
  NOR2_X1 U9712 ( .A1(n9800), .A2(n8050), .ZN(n8191) );
  INV_X1 U9713 ( .A(n8032), .ZN(n8033) );
  INV_X1 U9714 ( .A(n8038), .ZN(n8040) );
  NAND2_X1 U9715 ( .A1(n8040), .A2(n8039), .ZN(n8041) );
  MUX2_X1 U9716 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n5376), .Z(n8044) );
  INV_X1 U9717 ( .A(SI_31_), .ZN(n8043) );
  XNOR2_X1 U9718 ( .A(n8044), .B(n8043), .ZN(n8045) );
  NAND2_X1 U9719 ( .A1(n9210), .A2(n8047), .ZN(n8049) );
  NAND2_X1 U9720 ( .A1(n5630), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8048) );
  INV_X1 U9721 ( .A(n8924), .ZN(n8051) );
  NAND2_X1 U9722 ( .A1(n9800), .A2(n8050), .ZN(n8192) );
  NAND2_X1 U9723 ( .A1(n8200), .A2(n8192), .ZN(n8236) );
  NAND2_X1 U9724 ( .A1(n9795), .A2(n8051), .ZN(n8199) );
  INV_X1 U9725 ( .A(n8054), .ZN(n8055) );
  NOR2_X1 U9726 ( .A1(n8242), .A2(n4315), .ZN(n8056) );
  NAND2_X1 U9727 ( .A1(n9135), .A2(n8057), .ZN(n8061) );
  AND2_X1 U9728 ( .A1(n8059), .A2(n8058), .ZN(n8060) );
  MUX2_X1 U9729 ( .A(n8061), .B(n8060), .S(n8198), .Z(n8184) );
  NAND2_X1 U9730 ( .A1(n8172), .A2(n8062), .ZN(n8064) );
  INV_X1 U9731 ( .A(n9006), .ZN(n8063) );
  NAND2_X1 U9732 ( .A1(n8156), .A2(n8065), .ZN(n8068) );
  NAND2_X1 U9733 ( .A1(n8159), .A2(n8066), .ZN(n8067) );
  MUX2_X1 U9734 ( .A(n8068), .B(n8067), .S(n8201), .Z(n8069) );
  INV_X1 U9735 ( .A(n8069), .ZN(n8155) );
  NAND2_X1 U9736 ( .A1(n8070), .A2(n8071), .ZN(n8074) );
  INV_X1 U9737 ( .A(n8071), .ZN(n8072) );
  OAI211_X1 U9738 ( .C1(n8072), .C2(n8118), .A(n8130), .B(n8119), .ZN(n8073)
         );
  MUX2_X1 U9739 ( .A(n8074), .B(n8073), .S(n8201), .Z(n8075) );
  INV_X1 U9740 ( .A(n8075), .ZN(n8126) );
  NAND2_X1 U9741 ( .A1(n8080), .A2(n8079), .ZN(n8077) );
  NAND2_X1 U9742 ( .A1(n8100), .A2(n8098), .ZN(n8076) );
  AND2_X1 U9743 ( .A1(n8079), .A2(n8078), .ZN(n8081) );
  NAND2_X1 U9744 ( .A1(n8082), .A2(n8201), .ZN(n8089) );
  INV_X1 U9745 ( .A(n8102), .ZN(n8087) );
  AND2_X1 U9746 ( .A1(n8090), .A2(n8083), .ZN(n8084) );
  OAI211_X1 U9747 ( .C1(n6380), .C2(n8084), .A(n8093), .B(n6375), .ZN(n8085)
         );
  NAND3_X1 U9748 ( .A1(n8085), .A2(n8201), .A3(n5958), .ZN(n8086) );
  NAND3_X1 U9749 ( .A1(n8087), .A2(n10041), .A3(n8086), .ZN(n8088) );
  NAND2_X1 U9750 ( .A1(n8089), .A2(n8088), .ZN(n8096) );
  NAND2_X1 U9751 ( .A1(n6375), .A2(n8090), .ZN(n8091) );
  NAND3_X1 U9752 ( .A1(n5958), .A2(n8092), .A3(n8091), .ZN(n8094) );
  NAND3_X1 U9753 ( .A1(n8094), .A2(n8198), .A3(n8093), .ZN(n8095) );
  NAND2_X1 U9754 ( .A1(n10105), .A2(n8828), .ZN(n8099) );
  NAND3_X1 U9755 ( .A1(n8096), .A2(n8095), .A3(n8099), .ZN(n8105) );
  AND2_X1 U9756 ( .A1(n8098), .A2(n8097), .ZN(n8101) );
  OAI211_X1 U9757 ( .C1(n8102), .C2(n8101), .A(n8100), .B(n8099), .ZN(n8103)
         );
  NAND2_X1 U9758 ( .A1(n8103), .A2(n8198), .ZN(n8104) );
  NAND2_X1 U9759 ( .A1(n8105), .A2(n8104), .ZN(n8107) );
  INV_X1 U9760 ( .A(n8211), .ZN(n8106) );
  OAI211_X1 U9761 ( .C1(n8108), .C2(n8201), .A(n8107), .B(n8106), .ZN(n8112)
         );
  MUX2_X1 U9762 ( .A(n8110), .B(n8109), .S(n8201), .Z(n8111) );
  NAND3_X1 U9763 ( .A1(n8112), .A2(n8215), .A3(n8111), .ZN(n8117) );
  MUX2_X1 U9764 ( .A(n8114), .B(n8113), .S(n8198), .Z(n8115) );
  NAND3_X1 U9765 ( .A1(n8117), .A2(n8116), .A3(n8115), .ZN(n8124) );
  NAND3_X1 U9766 ( .A1(n8119), .A2(n8198), .A3(n8118), .ZN(n8120) );
  OAI21_X1 U9767 ( .B1(n8122), .B2(n8121), .A(n8120), .ZN(n8123) );
  NAND2_X1 U9768 ( .A1(n8124), .A2(n8123), .ZN(n8125) );
  NAND2_X1 U9769 ( .A1(n8126), .A2(n8125), .ZN(n8131) );
  INV_X1 U9770 ( .A(n8127), .ZN(n8129) );
  INV_X1 U9771 ( .A(n8134), .ZN(n8128) );
  AOI21_X1 U9772 ( .B1(n8131), .B2(n8129), .A(n8128), .ZN(n8137) );
  NAND2_X1 U9773 ( .A1(n8131), .A2(n8130), .ZN(n8133) );
  NAND2_X1 U9774 ( .A1(n8133), .A2(n8132), .ZN(n8135) );
  NAND2_X1 U9775 ( .A1(n8135), .A2(n8134), .ZN(n8136) );
  MUX2_X1 U9776 ( .A(n8137), .B(n8136), .S(n8198), .Z(n8141) );
  MUX2_X1 U9777 ( .A(n8139), .B(n8138), .S(n8201), .Z(n8140) );
  OAI211_X1 U9778 ( .C1(n8141), .C2(n8221), .A(n8224), .B(n8140), .ZN(n8145)
         );
  MUX2_X1 U9779 ( .A(n8143), .B(n8142), .S(n8198), .Z(n8144) );
  NAND3_X1 U9780 ( .A1(n8145), .A2(n8223), .A3(n8144), .ZN(n8149) );
  MUX2_X1 U9781 ( .A(n8147), .B(n8146), .S(n8198), .Z(n8148) );
  NAND3_X1 U9782 ( .A1(n8225), .A2(n8149), .A3(n8148), .ZN(n8153) );
  MUX2_X1 U9783 ( .A(n8151), .B(n8150), .S(n8201), .Z(n8152) );
  NAND3_X1 U9784 ( .A1(n8169), .A2(n8157), .A3(n9037), .ZN(n8168) );
  AOI21_X1 U9785 ( .B1(n8160), .B2(n8159), .A(n8158), .ZN(n8164) );
  NAND2_X1 U9786 ( .A1(n9059), .A2(n4521), .ZN(n8163) );
  OAI211_X1 U9787 ( .C1(n8164), .C2(n8163), .A(n8162), .B(n9037), .ZN(n8165)
         );
  NAND3_X1 U9788 ( .A1(n9024), .A2(n8166), .A3(n8165), .ZN(n8167) );
  MUX2_X1 U9789 ( .A(n8168), .B(n8167), .S(n8198), .Z(n8171) );
  MUX2_X1 U9790 ( .A(n8169), .B(n9024), .S(n8201), .Z(n8170) );
  MUX2_X1 U9791 ( .A(n8173), .B(n8172), .S(n8201), .Z(n8174) );
  NAND2_X1 U9792 ( .A1(n8177), .A2(n8176), .ZN(n8178) );
  NAND2_X1 U9793 ( .A1(n8178), .A2(n8201), .ZN(n8179) );
  NAND2_X1 U9794 ( .A1(n8180), .A2(n8179), .ZN(n8181) );
  OAI211_X1 U9795 ( .C1(n8198), .C2(n8182), .A(n8949), .B(n8181), .ZN(n8183)
         );
  NAND2_X1 U9796 ( .A1(n8184), .A2(n8183), .ZN(n8185) );
  OAI211_X1 U9797 ( .C1(n8198), .C2(n8640), .A(n8185), .B(n8188), .ZN(n8194)
         );
  NAND2_X1 U9798 ( .A1(n8185), .A2(n5892), .ZN(n8187) );
  INV_X1 U9799 ( .A(n8186), .ZN(n8195) );
  NAND4_X1 U9800 ( .A1(n8194), .A2(n8188), .A3(n8187), .A4(n8195), .ZN(n8190)
         );
  INV_X1 U9801 ( .A(n8189), .ZN(n8193) );
  INV_X1 U9802 ( .A(n8191), .ZN(n8197) );
  NAND2_X1 U9803 ( .A1(n8199), .A2(n8197), .ZN(n8234) );
  NAND2_X1 U9804 ( .A1(n8194), .A2(n8193), .ZN(n8196) );
  INV_X1 U9805 ( .A(n8199), .ZN(n8203) );
  INV_X1 U9806 ( .A(n8200), .ZN(n8202) );
  MUX2_X1 U9807 ( .A(n8203), .B(n8202), .S(n8201), .Z(n8204) );
  INV_X1 U9808 ( .A(n8240), .ZN(n8245) );
  OAI21_X1 U9809 ( .B1(n8238), .B2(n8239), .A(n10055), .ZN(n8244) );
  INV_X1 U9810 ( .A(n8205), .ZN(n8235) );
  INV_X1 U9811 ( .A(n9005), .ZN(n8997) );
  INV_X1 U9812 ( .A(n9101), .ZN(n9091) );
  INV_X1 U9813 ( .A(n9118), .ZN(n8227) );
  NOR3_X1 U9814 ( .A1(n8208), .A2(n8207), .A3(n8206), .ZN(n8209) );
  NAND4_X1 U9815 ( .A1(n10082), .A2(n8209), .A3(n10041), .A4(n8238), .ZN(n8213) );
  NOR4_X1 U9816 ( .A1(n8213), .A2(n8212), .A3(n8211), .A4(n8210), .ZN(n8214)
         );
  NAND4_X1 U9817 ( .A1(n8217), .A2(n8216), .A3(n8215), .A4(n8214), .ZN(n8218)
         );
  NOR4_X1 U9818 ( .A1(n8221), .A2(n8220), .A3(n8219), .A4(n8218), .ZN(n8222)
         );
  NAND4_X1 U9819 ( .A1(n8225), .A2(n8224), .A3(n8223), .A4(n8222), .ZN(n8226)
         );
  NOR4_X1 U9820 ( .A1(n9091), .A2(n8228), .A3(n8227), .A4(n8226), .ZN(n8229)
         );
  NAND4_X1 U9821 ( .A1(n9036), .A2(n9060), .A3(n9069), .A4(n8229), .ZN(n8230)
         );
  NOR4_X1 U9822 ( .A1(n8982), .A2(n8997), .A3(n9017), .A4(n8230), .ZN(n8231)
         );
  NAND4_X1 U9823 ( .A1(n8232), .A2(n8964), .A3(n8231), .A4(n8949), .ZN(n8233)
         );
  NOR4_X1 U9824 ( .A1(n8236), .A2(n8235), .A3(n8234), .A4(n8233), .ZN(n8237)
         );
  XNOR2_X1 U9825 ( .A(n8237), .B(n4315), .ZN(n8243) );
  AOI21_X1 U9826 ( .B1(n8240), .B2(n8239), .A(n8238), .ZN(n8241) );
  NOR3_X1 U9827 ( .A1(n8247), .A2(n8246), .A3(n9074), .ZN(n8250) );
  OAI21_X1 U9828 ( .B1(n8251), .B2(n8248), .A(P2_B_REG_SCAN_IN), .ZN(n8249) );
  XNOR2_X1 U9829 ( .A(n8788), .B(n8787), .ZN(n8258) );
  OAI22_X1 U9830 ( .A1(n8781), .A2(n8252), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8271), .ZN(n8256) );
  OAI22_X1 U9831 ( .A1(n8805), .A2(n8254), .B1(n8253), .B2(n10026), .ZN(n8255)
         );
  AOI211_X1 U9832 ( .C1(n10132), .C2(n8809), .A(n8256), .B(n8255), .ZN(n8257)
         );
  OAI21_X1 U9833 ( .B1(n8258), .B2(n8812), .A(n8257), .ZN(P2_U3219) );
  OAI211_X1 U9834 ( .C1(n8261), .C2(n8260), .A(n10029), .B(n8259), .ZN(n8269)
         );
  NOR2_X1 U9835 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8262), .ZN(n8267) );
  AOI211_X1 U9836 ( .C1(n8265), .C2(n8264), .A(n8263), .B(n10032), .ZN(n8266)
         );
  AOI211_X1 U9837 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n10034), .A(n8267), .B(
        n8266), .ZN(n8268) );
  OAI211_X1 U9838 ( .C1(n10030), .C2(n8270), .A(n8269), .B(n8268), .ZN(
        P2_U3262) );
  NOR2_X1 U9839 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8271), .ZN(n8276) );
  AOI211_X1 U9840 ( .C1(n8274), .C2(n8273), .A(n8272), .B(n10032), .ZN(n8275)
         );
  AOI211_X1 U9841 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n10034), .A(n8276), .B(
        n8275), .ZN(n8281) );
  OAI211_X1 U9842 ( .C1(n8279), .C2(n8278), .A(n10029), .B(n8277), .ZN(n8280)
         );
  OAI211_X1 U9843 ( .C1(n10030), .C2(n8282), .A(n8281), .B(n8280), .ZN(
        P2_U3255) );
  NOR2_X1 U9844 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5694), .ZN(n8287) );
  AOI211_X1 U9845 ( .C1(n8285), .C2(n8284), .A(n8283), .B(n10032), .ZN(n8286)
         );
  AOI211_X1 U9846 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n10034), .A(n8287), .B(
        n8286), .ZN(n8292) );
  OAI211_X1 U9847 ( .C1(n8290), .C2(n8289), .A(n8288), .B(n10029), .ZN(n8291)
         );
  OAI211_X1 U9848 ( .C1(n10030), .C2(n8293), .A(n8292), .B(n8291), .ZN(
        P2_U3254) );
  NAND2_X1 U9849 ( .A1(n9427), .A2(n9414), .ZN(n8294) );
  NAND2_X1 U9850 ( .A1(n8466), .A2(n8294), .ZN(n8297) );
  NAND2_X1 U9851 ( .A1(n8567), .A2(n9647), .ZN(n8295) );
  NAND2_X1 U9852 ( .A1(n8526), .A2(n8295), .ZN(n8296) );
  MUX2_X1 U9853 ( .A(n8297), .B(n8296), .S(n8415), .Z(n8378) );
  AND2_X1 U9854 ( .A1(n8359), .A2(n4833), .ZN(n8469) );
  MUX2_X1 U9855 ( .A(n8469), .B(n8514), .S(n8415), .Z(n8355) );
  INV_X1 U9856 ( .A(n8298), .ZN(n8299) );
  OR2_X1 U9857 ( .A1(n8300), .A2(n8299), .ZN(n8302) );
  MUX2_X1 U9858 ( .A(n8302), .B(n8301), .S(n8415), .Z(n8305) );
  AND2_X1 U9859 ( .A1(n8307), .A2(n8486), .ZN(n8478) );
  MUX2_X1 U9860 ( .A(n8478), .B(n8303), .S(n8415), .Z(n8304) );
  NAND2_X1 U9861 ( .A1(n8305), .A2(n8304), .ZN(n8311) );
  INV_X1 U9862 ( .A(n8306), .ZN(n8309) );
  MUX2_X1 U9863 ( .A(n8479), .B(n8307), .S(n8415), .Z(n8308) );
  AND2_X1 U9864 ( .A1(n8309), .A2(n8308), .ZN(n8310) );
  NAND2_X1 U9865 ( .A1(n8311), .A2(n8310), .ZN(n8316) );
  AND2_X1 U9866 ( .A1(n8313), .A2(n8312), .ZN(n8484) );
  NAND2_X1 U9867 ( .A1(n8319), .A2(n8435), .ZN(n8474) );
  AOI21_X1 U9868 ( .B1(n8316), .B2(n8484), .A(n8474), .ZN(n8318) );
  AND2_X1 U9869 ( .A1(n8435), .A2(n8480), .ZN(n8315) );
  INV_X1 U9870 ( .A(n8313), .ZN(n8314) );
  AOI21_X1 U9871 ( .B1(n8316), .B2(n8315), .A(n8314), .ZN(n8317) );
  NAND2_X1 U9872 ( .A1(n8320), .A2(n8319), .ZN(n8321) );
  AOI21_X1 U9873 ( .B1(n8328), .B2(n8490), .A(n8321), .ZN(n8323) );
  OAI211_X1 U9874 ( .C1(n8323), .C2(n8491), .A(n8338), .B(n8322), .ZN(n8332)
         );
  NAND2_X1 U9875 ( .A1(n8324), .A2(n8490), .ZN(n8327) );
  INV_X1 U9876 ( .A(n8325), .ZN(n8326) );
  OAI21_X1 U9877 ( .B1(n8328), .B2(n8327), .A(n8326), .ZN(n8330) );
  NAND3_X1 U9878 ( .A1(n8330), .A2(n8339), .A3(n8329), .ZN(n8331) );
  INV_X1 U9879 ( .A(n8415), .ZN(n8402) );
  INV_X1 U9880 ( .A(n9835), .ZN(n9836) );
  INV_X1 U9881 ( .A(n8338), .ZN(n8333) );
  OR2_X1 U9882 ( .A1(n8334), .A2(n8333), .ZN(n8335) );
  AND2_X1 U9883 ( .A1(n8335), .A2(n8344), .ZN(n8492) );
  AND2_X1 U9884 ( .A1(n8492), .A2(n8495), .ZN(n8342) );
  NAND2_X1 U9885 ( .A1(n8345), .A2(n8336), .ZN(n8493) );
  NAND2_X1 U9886 ( .A1(n8338), .A2(n8337), .ZN(n8472) );
  AND2_X1 U9887 ( .A1(n8472), .A2(n8339), .ZN(n8340) );
  NOR2_X1 U9888 ( .A1(n8493), .A2(n8340), .ZN(n8341) );
  MUX2_X1 U9889 ( .A(n8342), .B(n8341), .S(n8402), .Z(n8343) );
  AND2_X1 U9890 ( .A1(n9590), .A2(n8498), .ZN(n9613) );
  NAND2_X1 U9891 ( .A1(n8495), .A2(n8344), .ZN(n8346) );
  NAND2_X1 U9892 ( .A1(n8346), .A2(n8345), .ZN(n8348) );
  NAND2_X1 U9893 ( .A1(n8493), .A2(n8495), .ZN(n8347) );
  MUX2_X1 U9894 ( .A(n8348), .B(n8347), .S(n8415), .Z(n8349) );
  AND2_X1 U9895 ( .A1(n8502), .A2(n8498), .ZN(n8470) );
  MUX2_X1 U9896 ( .A(n8470), .B(n8501), .S(n8415), .Z(n8350) );
  MUX2_X1 U9897 ( .A(n8351), .B(n8502), .S(n8415), .Z(n8352) );
  NAND3_X1 U9898 ( .A1(n8353), .A2(n9583), .A3(n8352), .ZN(n8354) );
  INV_X1 U9899 ( .A(n8357), .ZN(n8358) );
  NOR2_X1 U9900 ( .A1(n9505), .A2(n8358), .ZN(n8512) );
  AND2_X1 U9901 ( .A1(n8509), .A2(n8359), .ZN(n8510) );
  INV_X1 U9902 ( .A(n9505), .ZN(n8360) );
  AND2_X1 U9903 ( .A1(n8360), .A2(n8511), .ZN(n8362) );
  INV_X1 U9904 ( .A(n8364), .ZN(n8361) );
  AOI21_X1 U9905 ( .B1(n8368), .B2(n8362), .A(n8361), .ZN(n8363) );
  OAI21_X1 U9906 ( .B1(n8363), .B2(n4556), .A(n8423), .ZN(n8369) );
  INV_X1 U9907 ( .A(n8511), .ZN(n8367) );
  NAND2_X1 U9908 ( .A1(n8511), .A2(n8424), .ZN(n8365) );
  AND2_X1 U9909 ( .A1(n8365), .A2(n8364), .ZN(n8366) );
  AND2_X1 U9910 ( .A1(n8366), .A2(n8423), .ZN(n8508) );
  OR2_X1 U9911 ( .A1(n9454), .A2(n8643), .ZN(n8564) );
  NAND2_X1 U9912 ( .A1(n8564), .A2(n8519), .ZN(n8373) );
  NAND2_X1 U9913 ( .A1(n8372), .A2(n8370), .ZN(n8565) );
  NOR2_X1 U9914 ( .A1(n8373), .A2(n8565), .ZN(n8371) );
  NAND2_X1 U9915 ( .A1(n8373), .A2(n8372), .ZN(n8374) );
  NAND2_X1 U9916 ( .A1(n9414), .A2(n8374), .ZN(n8376) );
  NAND2_X1 U9917 ( .A1(n8565), .A2(n8564), .ZN(n8375) );
  NAND2_X1 U9918 ( .A1(n8567), .A2(n8375), .ZN(n8468) );
  MUX2_X1 U9919 ( .A(n8376), .B(n8468), .S(n8402), .Z(n8377) );
  AND2_X1 U9920 ( .A1(n9414), .A2(n9440), .ZN(n8379) );
  INV_X1 U9921 ( .A(n8421), .ZN(n8464) );
  AOI21_X1 U9922 ( .B1(n8386), .B2(n8379), .A(n8464), .ZN(n8381) );
  AOI21_X1 U9923 ( .B1(n8389), .B2(n8381), .A(n8380), .ZN(n8382) );
  NAND2_X1 U9924 ( .A1(n8382), .A2(n8402), .ZN(n8392) );
  INV_X1 U9925 ( .A(n8567), .ZN(n8383) );
  NOR2_X1 U9926 ( .A1(n8383), .A2(n9427), .ZN(n8385) );
  INV_X1 U9927 ( .A(n8570), .ZN(n8384) );
  INV_X1 U9928 ( .A(n8466), .ZN(n8387) );
  AOI21_X1 U9929 ( .B1(n8389), .B2(n8388), .A(n8387), .ZN(n8390) );
  NAND2_X1 U9930 ( .A1(n8390), .A2(n8415), .ZN(n8391) );
  MUX2_X1 U9931 ( .A(n8467), .B(n8461), .S(n8415), .Z(n8393) );
  INV_X1 U9932 ( .A(n8393), .ZN(n8394) );
  INV_X1 U9933 ( .A(n9397), .ZN(n8396) );
  INV_X1 U9934 ( .A(n9322), .ZN(n8451) );
  NAND2_X1 U9935 ( .A1(n8456), .A2(n8411), .ZN(n8400) );
  NAND2_X1 U9936 ( .A1(n9210), .A2(n4998), .ZN(n8399) );
  OR2_X1 U9937 ( .A1(n8397), .A2(n6110), .ZN(n8398) );
  NAND2_X1 U9938 ( .A1(n8400), .A2(n8413), .ZN(n8531) );
  NAND2_X1 U9939 ( .A1(n9322), .A2(n8411), .ZN(n8401) );
  NAND2_X1 U9940 ( .A1(n8452), .A2(n8401), .ZN(n8528) );
  OAI211_X1 U9941 ( .C1(n9397), .C2(n8402), .A(n8531), .B(n8528), .ZN(n8403)
         );
  INV_X1 U9942 ( .A(n8403), .ZN(n8404) );
  NAND2_X1 U9943 ( .A1(n8405), .A2(n8404), .ZN(n8407) );
  NAND2_X1 U9944 ( .A1(n8407), .A2(n8406), .ZN(n8419) );
  NAND3_X1 U9945 ( .A1(n8410), .A2(n8396), .A3(n8528), .ZN(n8408) );
  NAND2_X1 U9946 ( .A1(n8408), .A2(n8531), .ZN(n8417) );
  NAND3_X1 U9947 ( .A1(n8410), .A2(n8409), .A3(n8531), .ZN(n8414) );
  INV_X1 U9948 ( .A(n8411), .ZN(n8412) );
  AND2_X1 U9949 ( .A1(n8413), .A2(n8412), .ZN(n8455) );
  AOI21_X1 U9950 ( .B1(n8414), .B2(n8528), .A(n8455), .ZN(n8416) );
  MUX2_X1 U9951 ( .A(n8417), .B(n8416), .S(n8415), .Z(n8418) );
  NAND2_X1 U9952 ( .A1(n8570), .A2(n8421), .ZN(n9423) );
  INV_X1 U9953 ( .A(n9437), .ZN(n9435) );
  INV_X1 U9954 ( .A(n8422), .ZN(n9471) );
  NAND2_X1 U9955 ( .A1(n8518), .A2(n8423), .ZN(n9488) );
  INV_X1 U9956 ( .A(n8426), .ZN(n8442) );
  AND2_X1 U9957 ( .A1(n9331), .A2(n8427), .ZN(n8542) );
  NOR2_X1 U9958 ( .A1(n8428), .A2(n8542), .ZN(n9927) );
  NAND4_X1 U9959 ( .A1(n8431), .A2(n9927), .A3(n8430), .A4(n8429), .ZN(n8434)
         );
  INV_X1 U9960 ( .A(n8480), .ZN(n8432) );
  NOR4_X1 U9961 ( .A1(n8434), .A2(n8433), .A3(n8432), .A4(n6827), .ZN(n8437)
         );
  NAND4_X1 U9962 ( .A1(n8437), .A2(n8484), .A3(n8436), .A4(n8435), .ZN(n8440)
         );
  NOR3_X1 U9963 ( .A1(n8440), .A2(n8439), .A3(n8438), .ZN(n8441) );
  NAND4_X1 U9964 ( .A1(n8443), .A2(n8442), .A3(n9835), .A4(n8441), .ZN(n8444)
         );
  NOR4_X1 U9965 ( .A1(n9593), .A2(n4427), .A3(n8445), .A4(n8444), .ZN(n8446)
         );
  NAND4_X1 U9966 ( .A1(n9547), .A2(n5228), .A3(n9583), .A4(n8446), .ZN(n8447)
         );
  NOR4_X1 U9967 ( .A1(n9488), .A2(n9504), .A3(n9520), .A4(n8447), .ZN(n8448)
         );
  INV_X1 U9968 ( .A(n9456), .ZN(n9449) );
  NAND4_X1 U9969 ( .A1(n9435), .A2(n9471), .A3(n8448), .A4(n9449), .ZN(n8449)
         );
  NOR4_X1 U9970 ( .A1(n8450), .A2(n4440), .A3(n9423), .A4(n8449), .ZN(n8454)
         );
  NAND2_X1 U9971 ( .A1(n8452), .A2(n8451), .ZN(n8577) );
  NAND4_X1 U9972 ( .A1(n8406), .A2(n8454), .A3(n8453), .A4(n8577), .ZN(n8459)
         );
  INV_X1 U9973 ( .A(n8455), .ZN(n8457) );
  NAND2_X1 U9974 ( .A1(n8457), .A2(n8456), .ZN(n8538) );
  OAI21_X1 U9975 ( .B1(n8459), .B2(n8538), .A(n8458), .ZN(n8534) );
  INV_X1 U9976 ( .A(n8461), .ZN(n8462) );
  NOR2_X1 U9977 ( .A1(n8463), .A2(n8462), .ZN(n8539) );
  NAND2_X1 U9978 ( .A1(n8526), .A2(n8464), .ZN(n8465) );
  AND3_X1 U9979 ( .A1(n8467), .A2(n8466), .A3(n8465), .ZN(n8572) );
  INV_X1 U9980 ( .A(n8468), .ZN(n8523) );
  INV_X1 U9981 ( .A(n8469), .ZN(n8505) );
  INV_X1 U9982 ( .A(n8470), .ZN(n8475) );
  INV_X1 U9983 ( .A(n8471), .ZN(n8473) );
  OR3_X1 U9984 ( .A1(n8493), .A2(n8473), .A3(n8472), .ZN(n8497) );
  OR3_X1 U9985 ( .A1(n8475), .A2(n8497), .A3(n8474), .ZN(n8476) );
  OR2_X1 U9986 ( .A1(n8505), .A2(n8476), .ZN(n8559) );
  NAND2_X1 U9987 ( .A1(n8551), .A2(n8477), .ZN(n8541) );
  INV_X1 U9988 ( .A(n8478), .ZN(n8481) );
  NAND3_X1 U9989 ( .A1(n8481), .A2(n8480), .A3(n8479), .ZN(n8482) );
  NAND3_X1 U9990 ( .A1(n8541), .A2(n8484), .A3(n8482), .ZN(n8489) );
  NAND2_X1 U9991 ( .A1(n8484), .A2(n8483), .ZN(n8550) );
  NAND2_X1 U9992 ( .A1(n8486), .A2(n8485), .ZN(n8487) );
  NOR2_X1 U9993 ( .A1(n8550), .A2(n8487), .ZN(n8552) );
  NAND2_X1 U9994 ( .A1(n8552), .A2(n6720), .ZN(n8488) );
  NAND2_X1 U9995 ( .A1(n8489), .A2(n8488), .ZN(n8506) );
  NOR2_X1 U9996 ( .A1(n8491), .A2(n4574), .ZN(n8496) );
  OR2_X1 U9997 ( .A1(n8493), .A2(n8492), .ZN(n8494) );
  OAI211_X1 U9998 ( .C1(n8497), .C2(n8496), .A(n8495), .B(n8494), .ZN(n8499)
         );
  NAND2_X1 U9999 ( .A1(n8499), .A2(n8498), .ZN(n8500) );
  NAND2_X1 U10000 ( .A1(n8501), .A2(n8500), .ZN(n8503) );
  NAND2_X1 U10001 ( .A1(n8503), .A2(n8502), .ZN(n8504) );
  OR2_X1 U10002 ( .A1(n8505), .A2(n8504), .ZN(n8557) );
  OAI21_X1 U10003 ( .B1(n8559), .B2(n8506), .A(n8557), .ZN(n8507) );
  INV_X1 U10004 ( .A(n8507), .ZN(n8521) );
  INV_X1 U10005 ( .A(n8508), .ZN(n8516) );
  OR2_X1 U10006 ( .A1(n8516), .A2(n4461), .ZN(n8540) );
  INV_X1 U10007 ( .A(n8510), .ZN(n8513) );
  OAI211_X1 U10008 ( .C1(n8514), .C2(n8513), .A(n8512), .B(n8511), .ZN(n8515)
         );
  INV_X1 U10009 ( .A(n8515), .ZN(n8517) );
  OR2_X1 U10010 ( .A1(n8517), .A2(n8516), .ZN(n8520) );
  AND3_X1 U10011 ( .A1(n8520), .A2(n8519), .A3(n8518), .ZN(n8560) );
  OAI211_X1 U10012 ( .C1(n8521), .C2(n8540), .A(n8560), .B(n8564), .ZN(n8522)
         );
  NAND2_X1 U10013 ( .A1(n8523), .A2(n8522), .ZN(n8524) );
  NAND3_X1 U10014 ( .A1(n8526), .A2(n8525), .A3(n8524), .ZN(n8527) );
  NAND2_X1 U10015 ( .A1(n8572), .A2(n8527), .ZN(n8530) );
  INV_X1 U10016 ( .A(n8528), .ZN(n8529) );
  AOI211_X1 U10017 ( .C1(n8539), .C2(n8530), .A(n8575), .B(n8529), .ZN(n8533)
         );
  INV_X1 U10018 ( .A(n8531), .ZN(n8532) );
  OAI211_X1 U10019 ( .C1(n8533), .C2(n8532), .A(n5410), .B(n8406), .ZN(n8535)
         );
  AND2_X1 U10020 ( .A1(n8535), .A2(n8534), .ZN(n8536) );
  INV_X1 U10021 ( .A(n8538), .ZN(n8581) );
  INV_X1 U10022 ( .A(n8539), .ZN(n8579) );
  INV_X1 U10023 ( .A(n8540), .ZN(n8563) );
  INV_X1 U10024 ( .A(n8541), .ZN(n8556) );
  INV_X1 U10025 ( .A(n8542), .ZN(n8544) );
  NAND2_X1 U10026 ( .A1(n6423), .A2(n9943), .ZN(n8543) );
  NAND3_X1 U10027 ( .A1(n8544), .A2(n5410), .A3(n8543), .ZN(n8545) );
  NAND2_X1 U10028 ( .A1(n8546), .A2(n8545), .ZN(n8548) );
  OAI22_X1 U10029 ( .A1(n8549), .A2(n8548), .B1(n8547), .B2(n6494), .ZN(n8555)
         );
  OR2_X1 U10030 ( .A1(n8551), .A2(n8550), .ZN(n8554) );
  INV_X1 U10031 ( .A(n8552), .ZN(n8553) );
  AOI22_X1 U10032 ( .A1(n8556), .A2(n8555), .B1(n8554), .B2(n8553), .ZN(n8558)
         );
  OAI21_X1 U10033 ( .B1(n8559), .B2(n8558), .A(n8557), .ZN(n8562) );
  INV_X1 U10034 ( .A(n8560), .ZN(n8561) );
  AOI21_X1 U10035 ( .B1(n8563), .B2(n8562), .A(n8561), .ZN(n8566) );
  OAI211_X1 U10036 ( .C1(n8566), .C2(n8565), .A(n9414), .B(n8564), .ZN(n8568)
         );
  NAND2_X1 U10037 ( .A1(n8568), .A2(n8567), .ZN(n8569) );
  AND3_X1 U10038 ( .A1(n8571), .A2(n8570), .A3(n8569), .ZN(n8574) );
  INV_X1 U10039 ( .A(n8572), .ZN(n8573) );
  NOR2_X1 U10040 ( .A1(n8574), .A2(n8573), .ZN(n8578) );
  INV_X1 U10041 ( .A(n8575), .ZN(n8576) );
  OAI211_X1 U10042 ( .C1(n8579), .C2(n8578), .A(n8577), .B(n8576), .ZN(n8580)
         );
  NAND2_X1 U10043 ( .A1(n8581), .A2(n8580), .ZN(n8582) );
  NAND2_X1 U10044 ( .A1(n8582), .A2(n8406), .ZN(n8587) );
  AND2_X1 U10045 ( .A1(n8583), .A2(n9513), .ZN(n9930) );
  NAND2_X1 U10046 ( .A1(n8587), .A2(n9930), .ZN(n8585) );
  OAI211_X1 U10047 ( .C1(n8587), .C2(n8586), .A(n8585), .B(n8584), .ZN(n8594)
         );
  NOR4_X1 U10048 ( .A1(n9925), .A2(n8589), .A3(n5433), .A4(n8588), .ZN(n8593)
         );
  OAI21_X1 U10049 ( .B1(n8591), .B2(n8590), .A(P1_B_REG_SCAN_IN), .ZN(n8592)
         );
  OAI22_X1 U10050 ( .A1(n8595), .A2(n8594), .B1(n8593), .B2(n8592), .ZN(
        P1_U3240) );
  INV_X1 U10051 ( .A(n8596), .ZN(n8599) );
  INV_X1 U10052 ( .A(n8597), .ZN(n8598) );
  NAND2_X1 U10053 ( .A1(n8599), .A2(n8598), .ZN(n8600) );
  XNOR2_X1 U10054 ( .A(n9164), .B(n8631), .ZN(n8605) );
  NAND2_X1 U10055 ( .A1(n9038), .A2(n10133), .ZN(n8603) );
  XNOR2_X1 U10056 ( .A(n8605), .B(n8603), .ZN(n8749) );
  INV_X1 U10057 ( .A(n8603), .ZN(n8604) );
  XNOR2_X1 U10058 ( .A(n9161), .B(n8606), .ZN(n8608) );
  XNOR2_X1 U10059 ( .A(n8607), .B(n8608), .ZN(n8778) );
  NAND2_X1 U10060 ( .A1(n9063), .A2(n10133), .ZN(n8777) );
  INV_X1 U10061 ( .A(n8607), .ZN(n8609) );
  NAND2_X1 U10062 ( .A1(n8609), .A2(n8608), .ZN(n8610) );
  NAND2_X1 U10063 ( .A1(n9039), .A2(n10133), .ZN(n8766) );
  INV_X1 U10064 ( .A(n8768), .ZN(n8613) );
  NAND2_X1 U10065 ( .A1(n9028), .A2(n10055), .ZN(n8617) );
  INV_X1 U10066 ( .A(n8617), .ZN(n8767) );
  NOR2_X2 U10067 ( .A1(n8620), .A2(n8619), .ZN(n8757) );
  NAND2_X1 U10068 ( .A1(n8965), .A2(n10133), .ZN(n8622) );
  XNOR2_X1 U10069 ( .A(n9146), .B(n8631), .ZN(n8621) );
  XOR2_X1 U10070 ( .A(n8622), .B(n8621), .Z(n8758) );
  XNOR2_X1 U10071 ( .A(n9140), .B(n8631), .ZN(n8625) );
  NAND2_X1 U10072 ( .A1(n8951), .A2(n10133), .ZN(n8623) );
  XNOR2_X1 U10073 ( .A(n8625), .B(n8623), .ZN(n8802) );
  INV_X1 U10074 ( .A(n8623), .ZN(n8624) );
  NAND2_X1 U10075 ( .A1(n8966), .A2(n10133), .ZN(n8628) );
  XNOR2_X1 U10076 ( .A(n9135), .B(n8631), .ZN(n8627) );
  XOR2_X1 U10077 ( .A(n8628), .B(n8627), .Z(n8734) );
  INV_X1 U10078 ( .A(n8627), .ZN(n8629) );
  NAND2_X1 U10079 ( .A1(n8952), .A2(n8630), .ZN(n8632) );
  XNOR2_X1 U10080 ( .A(n8632), .B(n8631), .ZN(n8633) );
  XNOR2_X1 U10081 ( .A(n8640), .B(n8633), .ZN(n8634) );
  INV_X1 U10082 ( .A(n8635), .ZN(n8937) );
  AOI22_X1 U10083 ( .A1(n8937), .A2(n8784), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8636) );
  OAI21_X1 U10084 ( .B1(n8638), .B2(n8637), .A(n8636), .ZN(n8639) );
  AOI21_X1 U10085 ( .B1(n8640), .B2(n8809), .A(n8639), .ZN(n8641) );
  OAI21_X1 U10086 ( .B1(n8642), .B2(n8812), .A(n8641), .ZN(P2_U3222) );
  OAI22_X1 U10087 ( .A1(n9660), .A2(n6498), .B1(n8643), .B2(n8719), .ZN(n8697)
         );
  INV_X1 U10088 ( .A(n8697), .ZN(n8700) );
  OAI22_X1 U10089 ( .A1(n9660), .A2(n8718), .B1(n8643), .B2(n6498), .ZN(n8644)
         );
  XNOR2_X1 U10090 ( .A(n8644), .B(n8721), .ZN(n8698) );
  INV_X1 U10091 ( .A(n8698), .ZN(n8699) );
  NAND2_X1 U10092 ( .A1(n8646), .A2(n8645), .ZN(n8651) );
  INV_X1 U10093 ( .A(n8647), .ZN(n8649) );
  NAND2_X1 U10094 ( .A1(n8649), .A2(n8648), .ZN(n8650) );
  NAND2_X1 U10095 ( .A1(n8651), .A2(n8650), .ZN(n8657) );
  NAND2_X1 U10096 ( .A1(n9566), .A2(n8714), .ZN(n8653) );
  OR2_X1 U10097 ( .A1(n9690), .A2(n6498), .ZN(n8652) );
  NAND2_X1 U10098 ( .A1(n8653), .A2(n8652), .ZN(n8654) );
  XNOR2_X1 U10099 ( .A(n8654), .B(n8689), .ZN(n8658) );
  NAND2_X1 U10100 ( .A1(n8657), .A2(n8658), .ZN(n9298) );
  NAND2_X1 U10101 ( .A1(n9566), .A2(n8716), .ZN(n8656) );
  OR2_X1 U10102 ( .A1(n9690), .A2(n8719), .ZN(n8655) );
  NAND2_X1 U10103 ( .A1(n8656), .A2(n8655), .ZN(n9301) );
  NAND2_X1 U10104 ( .A1(n9298), .A2(n9301), .ZN(n8661) );
  NAND2_X1 U10105 ( .A1(n9752), .A2(n8714), .ZN(n8663) );
  NAND2_X1 U10106 ( .A1(n9681), .A2(n8716), .ZN(n8662) );
  NAND2_X1 U10107 ( .A1(n8663), .A2(n8662), .ZN(n8664) );
  XNOR2_X1 U10108 ( .A(n8664), .B(n8689), .ZN(n8667) );
  AND2_X1 U10109 ( .A1(n9681), .A2(n6414), .ZN(n8665) );
  AOI21_X1 U10110 ( .B1(n9752), .B2(n8706), .A(n8665), .ZN(n8666) );
  XNOR2_X1 U10111 ( .A(n8667), .B(n8666), .ZN(n9243) );
  NAND2_X1 U10112 ( .A1(n8667), .A2(n8666), .ZN(n9276) );
  NAND2_X1 U10113 ( .A1(n9533), .A2(n8714), .ZN(n8669) );
  NAND2_X1 U10114 ( .A1(n9543), .A2(n8716), .ZN(n8668) );
  NAND2_X1 U10115 ( .A1(n8669), .A2(n8668), .ZN(n8670) );
  XNOR2_X1 U10116 ( .A(n8670), .B(n8721), .ZN(n8675) );
  INV_X1 U10117 ( .A(n8675), .ZN(n8672) );
  AND2_X1 U10118 ( .A1(n9543), .A2(n6414), .ZN(n8671) );
  AOI21_X1 U10119 ( .B1(n9533), .B2(n8706), .A(n8671), .ZN(n8674) );
  NAND2_X1 U10120 ( .A1(n8672), .A2(n8674), .ZN(n8673) );
  INV_X1 U10121 ( .A(n8673), .ZN(n8676) );
  XNOR2_X1 U10122 ( .A(n8675), .B(n8674), .ZN(n9279) );
  NAND2_X1 U10123 ( .A1(n9502), .A2(n8714), .ZN(n8678) );
  OR2_X1 U10124 ( .A1(n9528), .A2(n6498), .ZN(n8677) );
  NAND2_X1 U10125 ( .A1(n8678), .A2(n8677), .ZN(n8679) );
  XNOR2_X1 U10126 ( .A(n8679), .B(n8721), .ZN(n8681) );
  NOR2_X1 U10127 ( .A1(n9528), .A2(n8719), .ZN(n8680) );
  AOI21_X1 U10128 ( .B1(n9502), .B2(n8716), .A(n8680), .ZN(n8682) );
  XNOR2_X1 U10129 ( .A(n8681), .B(n8682), .ZN(n9250) );
  INV_X1 U10130 ( .A(n8681), .ZN(n8683) );
  AND2_X1 U10131 ( .A1(n8683), .A2(n8682), .ZN(n8684) );
  AOI21_X1 U10132 ( .B1(n9251), .B2(n9250), .A(n8684), .ZN(n8692) );
  NAND2_X1 U10133 ( .A1(n9491), .A2(n8716), .ZN(n8686) );
  NAND2_X1 U10134 ( .A1(n9510), .A2(n6414), .ZN(n8685) );
  NAND2_X1 U10135 ( .A1(n8686), .A2(n8685), .ZN(n8691) );
  NOR2_X2 U10136 ( .A1(n8692), .A2(n8691), .ZN(n9287) );
  NAND2_X1 U10137 ( .A1(n9491), .A2(n8714), .ZN(n8688) );
  NAND2_X1 U10138 ( .A1(n9510), .A2(n8716), .ZN(n8687) );
  NAND2_X1 U10139 ( .A1(n8688), .A2(n8687), .ZN(n8690) );
  XNOR2_X1 U10140 ( .A(n8690), .B(n8689), .ZN(n9288) );
  NOR2_X1 U10141 ( .A1(n9287), .A2(n9288), .ZN(n9286) );
  NAND2_X1 U10142 ( .A1(n9667), .A2(n8714), .ZN(n8694) );
  NAND2_X1 U10143 ( .A1(n9657), .A2(n8706), .ZN(n8693) );
  NAND2_X1 U10144 ( .A1(n8694), .A2(n8693), .ZN(n8695) );
  XNOR2_X1 U10145 ( .A(n8695), .B(n8721), .ZN(n8696) );
  NOR3_X2 U10146 ( .A1(n9286), .A2(n9290), .A3(n8696), .ZN(n9233) );
  AOI22_X1 U10147 ( .A1(n9667), .A2(n8716), .B1(n6414), .B2(n9657), .ZN(n9236)
         );
  OAI21_X1 U10148 ( .B1(n9286), .B2(n9290), .A(n8696), .ZN(n9234) );
  OAI21_X1 U10149 ( .B1(n9233), .B2(n9236), .A(n9234), .ZN(n9267) );
  XNOR2_X1 U10150 ( .A(n8698), .B(n8697), .ZN(n9268) );
  NOR2_X1 U10151 ( .A1(n9267), .A2(n9268), .ZN(n9266) );
  NAND2_X1 U10152 ( .A1(n5355), .A2(n8714), .ZN(n8702) );
  OR2_X1 U10153 ( .A1(n9419), .A2(n6498), .ZN(n8701) );
  NAND2_X1 U10154 ( .A1(n8702), .A2(n8701), .ZN(n8703) );
  XNOR2_X1 U10155 ( .A(n8703), .B(n8721), .ZN(n8705) );
  OAI22_X1 U10156 ( .A1(n9651), .A2(n6498), .B1(n9419), .B2(n8719), .ZN(n8704)
         );
  XNOR2_X1 U10157 ( .A(n8705), .B(n8704), .ZN(n9259) );
  AOI22_X1 U10158 ( .A1(n9427), .A2(n8706), .B1(n6414), .B2(n9647), .ZN(n8710)
         );
  NAND2_X1 U10159 ( .A1(n9427), .A2(n8714), .ZN(n8708) );
  NAND2_X1 U10160 ( .A1(n9647), .A2(n8706), .ZN(n8707) );
  NAND2_X1 U10161 ( .A1(n8708), .A2(n8707), .ZN(n8709) );
  XOR2_X1 U10162 ( .A(n8710), .B(n8712), .Z(n9317) );
  INV_X1 U10163 ( .A(n8710), .ZN(n8711) );
  AOI22_X1 U10164 ( .A1(n5390), .A2(n8714), .B1(n8716), .B2(n9395), .ZN(n8715)
         );
  XNOR2_X1 U10165 ( .A(n8721), .B(n8715), .ZN(n9224) );
  AOI22_X1 U10166 ( .A1(n5390), .A2(n8716), .B1(n6414), .B2(n9395), .ZN(n9223)
         );
  OAI22_X1 U10167 ( .A1(n8717), .A2(n9223), .B1(n9226), .B2(n9224), .ZN(n8726)
         );
  OAI22_X1 U10168 ( .A1(n8720), .A2(n8718), .B1(n9228), .B2(n6498), .ZN(n8724)
         );
  OAI22_X1 U10169 ( .A1(n8720), .A2(n6498), .B1(n9228), .B2(n8719), .ZN(n8722)
         );
  XNOR2_X1 U10170 ( .A(n8722), .B(n8721), .ZN(n8723) );
  XOR2_X1 U10171 ( .A(n8724), .B(n8723), .Z(n8725) );
  XNOR2_X1 U10172 ( .A(n8726), .B(n8725), .ZN(n8731) );
  NOR2_X1 U10173 ( .A1(n9282), .A2(n9392), .ZN(n8729) );
  AOI22_X1 U10174 ( .A1(n9395), .A2(n9302), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8727) );
  OAI21_X1 U10175 ( .B1(n9397), .B2(n9304), .A(n8727), .ZN(n8728) );
  AOI211_X1 U10176 ( .C1(n9401), .C2(n9320), .A(n8729), .B(n8728), .ZN(n8730)
         );
  OAI21_X1 U10177 ( .B1(n8731), .B2(n9315), .A(n8730), .ZN(P1_U3218) );
  INV_X1 U10178 ( .A(n8732), .ZN(n9216) );
  OAI222_X1 U10179 ( .A1(n9781), .A2(n9216), .B1(n4866), .B2(P1_U3084), .C1(
        n8733), .C2(n9777), .ZN(P1_U3323) );
  XNOR2_X1 U10180 ( .A(n8735), .B(n8734), .ZN(n8741) );
  OAI22_X1 U10181 ( .A1(n8989), .A2(n8805), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8736), .ZN(n8739) );
  INV_X1 U10182 ( .A(n8956), .ZN(n8737) );
  OAI22_X1 U10183 ( .A1(n5892), .A2(n8781), .B1(n8737), .B2(n10026), .ZN(n8738) );
  AOI211_X1 U10184 ( .C1(n9135), .C2(n8809), .A(n8739), .B(n8738), .ZN(n8740)
         );
  OAI21_X1 U10185 ( .B1(n8741), .B2(n8812), .A(n8740), .ZN(P2_U3216) );
  XNOR2_X1 U10186 ( .A(n8742), .B(n8766), .ZN(n8747) );
  OAI22_X1 U10187 ( .A1(n8988), .A2(n8781), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8743), .ZN(n8745) );
  OAI22_X1 U10188 ( .A1(n8805), .A2(n8751), .B1(n10026), .B2(n9020), .ZN(n8744) );
  AOI211_X1 U10189 ( .C1(n9154), .C2(n8809), .A(n8745), .B(n8744), .ZN(n8746)
         );
  OAI21_X1 U10190 ( .B1(n8747), .B2(n8812), .A(n8746), .ZN(P2_U3218) );
  XNOR2_X1 U10191 ( .A(n8748), .B(n8749), .ZN(n8756) );
  OAI22_X1 U10192 ( .A1(n8781), .A2(n8751), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8750), .ZN(n8754) );
  OAI22_X1 U10193 ( .A1(n8805), .A2(n8752), .B1(n9054), .B2(n10026), .ZN(n8753) );
  AOI211_X1 U10194 ( .C1(n9164), .C2(n8809), .A(n8754), .B(n8753), .ZN(n8755)
         );
  OAI21_X1 U10195 ( .B1(n8756), .B2(n8812), .A(n8755), .ZN(P2_U3225) );
  XNOR2_X1 U10196 ( .A(n8757), .B(n8758), .ZN(n8764) );
  OAI22_X1 U10197 ( .A1(n8989), .A2(n8781), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8759), .ZN(n8762) );
  INV_X1 U10198 ( .A(n8991), .ZN(n8760) );
  OAI22_X1 U10199 ( .A1(n8760), .A2(n10026), .B1(n8988), .B2(n8805), .ZN(n8761) );
  AOI211_X1 U10200 ( .C1(n9146), .C2(n8809), .A(n8762), .B(n8761), .ZN(n8763)
         );
  OAI21_X1 U10201 ( .B1(n8764), .B2(n8812), .A(n8763), .ZN(P2_U3227) );
  OAI21_X1 U10202 ( .B1(n8742), .B2(n8766), .A(n8765), .ZN(n8770) );
  XNOR2_X1 U10203 ( .A(n8768), .B(n8767), .ZN(n8769) );
  XNOR2_X1 U10204 ( .A(n8770), .B(n8769), .ZN(n8775) );
  OAI22_X1 U10205 ( .A1(n9010), .A2(n8781), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8771), .ZN(n8773) );
  OAI22_X1 U10206 ( .A1(n9009), .A2(n8805), .B1(n10026), .B2(n9002), .ZN(n8772) );
  AOI211_X1 U10207 ( .C1(n9149), .C2(n8809), .A(n8773), .B(n8772), .ZN(n8774)
         );
  OAI21_X1 U10208 ( .B1(n8775), .B2(n8812), .A(n8774), .ZN(P2_U3231) );
  OAI21_X1 U10209 ( .B1(n8778), .B2(n8777), .A(n8776), .ZN(n8779) );
  NAND2_X1 U10210 ( .A1(n8779), .A2(n10022), .ZN(n8786) );
  NOR2_X1 U10211 ( .A1(n8805), .A2(n9077), .ZN(n8783) );
  OAI22_X1 U10212 ( .A1(n9009), .A2(n8781), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8780), .ZN(n8782) );
  AOI211_X1 U10213 ( .C1(n8784), .C2(n9045), .A(n8783), .B(n8782), .ZN(n8785)
         );
  OAI211_X1 U10214 ( .C1(n4490), .C2(n10020), .A(n8786), .B(n8785), .ZN(
        P2_U3237) );
  OR2_X1 U10215 ( .A1(n8788), .A2(n8787), .ZN(n8790) );
  NAND2_X1 U10216 ( .A1(n8790), .A2(n8789), .ZN(n8791) );
  XOR2_X1 U10217 ( .A(n8792), .B(n8791), .Z(n8793) );
  NAND2_X1 U10218 ( .A1(n8793), .A2(n10022), .ZN(n8801) );
  AOI21_X1 U10219 ( .B1(n10018), .B2(n8795), .A(n8794), .ZN(n8800) );
  NAND2_X1 U10220 ( .A1(n8809), .A2(n10141), .ZN(n8799) );
  INV_X1 U10221 ( .A(n8796), .ZN(n8797) );
  OR2_X1 U10222 ( .A1(n10026), .A2(n8797), .ZN(n8798) );
  NAND4_X1 U10223 ( .A1(n8801), .A2(n8800), .A3(n8799), .A4(n8798), .ZN(
        P2_U3238) );
  XNOR2_X1 U10224 ( .A(n8803), .B(n8802), .ZN(n8813) );
  NOR2_X1 U10225 ( .A1(n8976), .A2(n10026), .ZN(n8807) );
  OAI22_X1 U10226 ( .A1(n9010), .A2(n8805), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8804), .ZN(n8806) );
  AOI211_X1 U10227 ( .C1(n8808), .C2(n8966), .A(n8807), .B(n8806), .ZN(n8811)
         );
  NAND2_X1 U10228 ( .A1(n9140), .A2(n8809), .ZN(n8810) );
  OAI211_X1 U10229 ( .C1(n8813), .C2(n8812), .A(n8811), .B(n8810), .ZN(
        P2_U3242) );
  MUX2_X1 U10230 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8814), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U10231 ( .A(n8815), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8816), .Z(
        P2_U3581) );
  MUX2_X1 U10232 ( .A(n8952), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8816), .Z(
        P2_U3580) );
  MUX2_X1 U10233 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8966), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U10234 ( .A(n8951), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8816), .Z(
        P2_U3578) );
  MUX2_X1 U10235 ( .A(n8965), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8816), .Z(
        P2_U3577) );
  MUX2_X1 U10236 ( .A(n9028), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8816), .Z(
        P2_U3576) );
  MUX2_X1 U10237 ( .A(n9039), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8816), .Z(
        P2_U3575) );
  MUX2_X1 U10238 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9063), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10239 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9038), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U10240 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9062), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U10241 ( .A(n9120), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8816), .Z(
        P2_U3571) );
  MUX2_X1 U10242 ( .A(n8817), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8816), .Z(
        P2_U3570) );
  MUX2_X1 U10243 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9119), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U10244 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8818), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10245 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8819), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10246 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8820), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U10247 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8821), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U10248 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8822), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U10249 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8823), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U10250 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8824), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U10251 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8825), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U10252 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8826), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U10253 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8827), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U10254 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8828), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U10255 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8829), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U10256 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n10047), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U10257 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n5620), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U10258 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n6385), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U10259 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6463), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U10260 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n6384), .S(P2_U3966), .Z(
        P2_U3552) );
  NAND2_X1 U10261 ( .A1(n8896), .A2(n8830), .ZN(n8842) );
  AND2_X1 U10262 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n8835) );
  INV_X1 U10263 ( .A(n8831), .ZN(n8834) );
  INV_X1 U10264 ( .A(n8832), .ZN(n8833) );
  OAI211_X1 U10265 ( .C1(n8835), .C2(n8834), .A(n10029), .B(n8833), .ZN(n8841)
         );
  AOI22_X1 U10266 ( .A1(n10034), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n8840) );
  OAI211_X1 U10267 ( .C1(n8838), .C2(n8837), .A(n10027), .B(n8836), .ZN(n8839)
         );
  NAND4_X1 U10268 ( .A1(n8842), .A2(n8841), .A3(n8840), .A4(n8839), .ZN(
        P2_U3246) );
  NAND2_X1 U10269 ( .A1(n8896), .A2(n8843), .ZN(n8857) );
  NOR2_X1 U10270 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10061), .ZN(n8844) );
  AOI21_X1 U10271 ( .B1(n10034), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n8844), .ZN(
        n8856) );
  INV_X1 U10272 ( .A(n8845), .ZN(n8863) );
  NAND3_X1 U10273 ( .A1(n8848), .A2(n8847), .A3(n8846), .ZN(n8849) );
  NAND3_X1 U10274 ( .A1(n10029), .A2(n8863), .A3(n8849), .ZN(n8855) );
  OAI21_X1 U10275 ( .B1(n8852), .B2(n8851), .A(n8850), .ZN(n8853) );
  OR2_X1 U10276 ( .A1(n10032), .A2(n8853), .ZN(n8854) );
  NAND4_X1 U10277 ( .A1(n8857), .A2(n8856), .A3(n8855), .A4(n8854), .ZN(
        P2_U3248) );
  NAND2_X1 U10278 ( .A1(n8896), .A2(n8860), .ZN(n8873) );
  AOI21_X1 U10279 ( .B1(n10034), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n8858), .ZN(
        n8872) );
  INV_X1 U10280 ( .A(n8859), .ZN(n8862) );
  MUX2_X1 U10281 ( .A(n6285), .B(P2_REG2_REG_4__SCAN_IN), .S(n8860), .Z(n8861)
         );
  NAND3_X1 U10282 ( .A1(n8863), .A2(n8862), .A3(n8861), .ZN(n8864) );
  NAND3_X1 U10283 ( .A1(n10029), .A2(n8865), .A3(n8864), .ZN(n8871) );
  OAI21_X1 U10284 ( .B1(n8868), .B2(n8867), .A(n8866), .ZN(n8869) );
  OR2_X1 U10285 ( .A1(n10032), .A2(n8869), .ZN(n8870) );
  NAND4_X1 U10286 ( .A1(n8873), .A2(n8872), .A3(n8871), .A4(n8870), .ZN(
        P2_U3249) );
  NAND2_X1 U10287 ( .A1(n8896), .A2(n8874), .ZN(n8887) );
  OAI211_X1 U10288 ( .C1(n8877), .C2(n8876), .A(n10029), .B(n8875), .ZN(n8886)
         );
  NOR2_X1 U10289 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8878), .ZN(n8879) );
  AOI21_X1 U10290 ( .B1(n10034), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8879), .ZN(
        n8885) );
  AND2_X1 U10291 ( .A1(n8881), .A2(n8880), .ZN(n8882) );
  OR3_X1 U10292 ( .A1(n10032), .A2(n8883), .A3(n8882), .ZN(n8884) );
  NAND4_X1 U10293 ( .A1(n8887), .A2(n8886), .A3(n8885), .A4(n8884), .ZN(
        P2_U3253) );
  OAI21_X1 U10294 ( .B1(n8890), .B2(n8889), .A(n8888), .ZN(n8891) );
  NAND2_X1 U10295 ( .A1(n8891), .A2(n10027), .ZN(n8902) );
  INV_X1 U10296 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8893) );
  OAI21_X1 U10297 ( .B1(n8922), .B2(n8893), .A(n8892), .ZN(n8894) );
  AOI21_X1 U10298 ( .B1(n8896), .B2(n8895), .A(n8894), .ZN(n8901) );
  OAI211_X1 U10299 ( .C1(n8899), .C2(n8898), .A(n10029), .B(n8897), .ZN(n8900)
         );
  NAND3_X1 U10300 ( .A1(n8902), .A2(n8901), .A3(n8900), .ZN(P2_U3261) );
  INV_X1 U10301 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8921) );
  OAI21_X1 U10302 ( .B1(n8907), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8903), .ZN(
        n8905) );
  XOR2_X1 U10303 ( .A(n8905), .B(n8904), .Z(n8915) );
  NOR2_X1 U10304 ( .A1(n8907), .A2(n8906), .ZN(n8909) );
  NOR2_X1 U10305 ( .A1(n8909), .A2(n8908), .ZN(n8910) );
  XNOR2_X1 U10306 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8910), .ZN(n8913) );
  NAND2_X1 U10307 ( .A1(n8913), .A2(n10029), .ZN(n8911) );
  OAI211_X1 U10308 ( .C1(n8915), .C2(n10032), .A(n8911), .B(n10030), .ZN(n8912) );
  INV_X1 U10309 ( .A(n8912), .ZN(n8918) );
  INV_X1 U10310 ( .A(n8913), .ZN(n8914) );
  AOI22_X1 U10311 ( .A1(n8915), .A2(n10027), .B1(n10029), .B2(n8914), .ZN(
        n8917) );
  MUX2_X1 U10312 ( .A(n8918), .B(n8917), .S(n4315), .Z(n8920) );
  OAI211_X1 U10313 ( .C1(n8922), .C2(n8921), .A(n8920), .B(n8919), .ZN(
        P2_U3264) );
  INV_X1 U10314 ( .A(n9800), .ZN(n8931) );
  NAND2_X1 U10315 ( .A1(n8931), .A2(n8930), .ZN(n8929) );
  XNOR2_X1 U10316 ( .A(n8929), .B(n9795), .ZN(n9793) );
  AND2_X1 U10317 ( .A1(n8924), .A2(n8923), .ZN(n9799) );
  INV_X1 U10318 ( .A(n9799), .ZN(n8925) );
  NOR2_X1 U10319 ( .A1(n10070), .A2(n8925), .ZN(n8933) );
  AOI21_X1 U10320 ( .B1(n10070), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8933), .ZN(
        n8928) );
  NAND2_X1 U10321 ( .A1(n9795), .A2(n8926), .ZN(n8927) );
  OAI211_X1 U10322 ( .C1(n9793), .C2(n8935), .A(n8928), .B(n8927), .ZN(
        P2_U3265) );
  OAI21_X1 U10323 ( .B1(n8931), .B2(n8930), .A(n8929), .ZN(n9797) );
  NOR2_X1 U10324 ( .A1(n8931), .A2(n10054), .ZN(n8932) );
  AOI211_X1 U10325 ( .C1(n10070), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8933), .B(
        n8932), .ZN(n8934) );
  OAI21_X1 U10326 ( .B1(n8935), .B2(n9797), .A(n8934), .ZN(P2_U3266) );
  NAND2_X1 U10327 ( .A1(n8936), .A2(n9124), .ZN(n8939) );
  AOI22_X1 U10328 ( .A1(n8937), .A2(n10062), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n10070), .ZN(n8938) );
  OAI211_X1 U10329 ( .C1(n5893), .C2(n10054), .A(n8939), .B(n8938), .ZN(n8940)
         );
  AOI21_X1 U10330 ( .B1(n8941), .B2(n9049), .A(n8940), .ZN(n8942) );
  OAI21_X1 U10331 ( .B1(n8943), .B2(n9126), .A(n8942), .ZN(P2_U3268) );
  OAI21_X1 U10332 ( .B1(n8946), .B2(n8945), .A(n8944), .ZN(n8947) );
  INV_X1 U10333 ( .A(n8947), .ZN(n9137) );
  OAI211_X1 U10334 ( .C1(n8950), .C2(n8949), .A(n8948), .B(n10049), .ZN(n8954)
         );
  AOI22_X1 U10335 ( .A1(n8952), .A2(n10046), .B1(n10045), .B2(n8951), .ZN(
        n8953) );
  NAND2_X1 U10336 ( .A1(n8954), .A2(n8953), .ZN(n9133) );
  INV_X1 U10337 ( .A(n9135), .ZN(n8959) );
  AOI211_X1 U10338 ( .C1(n9135), .C2(n8971), .A(n10055), .B(n8955), .ZN(n9134)
         );
  NAND2_X1 U10339 ( .A1(n9134), .A2(n9124), .ZN(n8958) );
  AOI22_X1 U10340 ( .A1(n8956), .A2(n10062), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n10070), .ZN(n8957) );
  OAI211_X1 U10341 ( .C1(n8959), .C2(n10054), .A(n8958), .B(n8957), .ZN(n8960)
         );
  AOI21_X1 U10342 ( .B1(n9133), .B2(n9049), .A(n8960), .ZN(n8961) );
  OAI21_X1 U10343 ( .B1(n9137), .B2(n9126), .A(n8961), .ZN(P2_U3269) );
  OAI21_X1 U10344 ( .B1(n8964), .B2(n8963), .A(n8962), .ZN(n8967) );
  AOI222_X1 U10345 ( .A1(n10049), .A2(n8967), .B1(n8966), .B2(n10046), .C1(
        n8965), .C2(n10045), .ZN(n9142) );
  OAI21_X1 U10346 ( .B1(n8970), .B2(n8969), .A(n8968), .ZN(n9138) );
  NAND2_X1 U10347 ( .A1(n9138), .A2(n9082), .ZN(n8980) );
  INV_X1 U10348 ( .A(n8990), .ZN(n8973) );
  INV_X1 U10349 ( .A(n8971), .ZN(n8972) );
  AOI211_X1 U10350 ( .C1(n9140), .C2(n8973), .A(n10055), .B(n8972), .ZN(n9139)
         );
  NOR2_X1 U10351 ( .A1(n5868), .A2(n10054), .ZN(n8978) );
  OAI22_X1 U10352 ( .A1(n8976), .A2(n8975), .B1(n8974), .B2(n9049), .ZN(n8977)
         );
  AOI211_X1 U10353 ( .C1(n9139), .C2(n9124), .A(n8978), .B(n8977), .ZN(n8979)
         );
  OAI211_X1 U10354 ( .C1(n10070), .C2(n9142), .A(n8980), .B(n8979), .ZN(
        P2_U3270) );
  OAI21_X1 U10355 ( .B1(n8983), .B2(n8982), .A(n8981), .ZN(n8984) );
  INV_X1 U10356 ( .A(n8984), .ZN(n9148) );
  XNOR2_X1 U10357 ( .A(n8985), .B(n8986), .ZN(n8987) );
  OAI222_X1 U10358 ( .A1(n9076), .A2(n8989), .B1(n9074), .B2(n8988), .C1(n9071), .C2(n8987), .ZN(n9144) );
  INV_X1 U10359 ( .A(n9146), .ZN(n8994) );
  AOI211_X1 U10360 ( .C1(n9146), .C2(n8999), .A(n10055), .B(n8990), .ZN(n9145)
         );
  NAND2_X1 U10361 ( .A1(n9145), .A2(n9124), .ZN(n8993) );
  AOI22_X1 U10362 ( .A1(n8991), .A2(n10062), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n10070), .ZN(n8992) );
  OAI211_X1 U10363 ( .C1(n8994), .C2(n10054), .A(n8993), .B(n8992), .ZN(n8995)
         );
  AOI21_X1 U10364 ( .B1(n9144), .B2(n9049), .A(n8995), .ZN(n8996) );
  OAI21_X1 U10365 ( .B1(n9148), .B2(n9126), .A(n8996), .ZN(P2_U3271) );
  XNOR2_X1 U10366 ( .A(n8998), .B(n8997), .ZN(n9153) );
  INV_X1 U10367 ( .A(n9019), .ZN(n9001) );
  INV_X1 U10368 ( .A(n8999), .ZN(n9000) );
  AOI21_X1 U10369 ( .B1(n9149), .B2(n9001), .A(n9000), .ZN(n9150) );
  INV_X1 U10370 ( .A(n9002), .ZN(n9003) );
  AOI22_X1 U10371 ( .A1(n9003), .A2(n10062), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n10070), .ZN(n9004) );
  OAI21_X1 U10372 ( .B1(n4802), .B2(n10054), .A(n9004), .ZN(n9014) );
  AOI21_X1 U10373 ( .B1(n9025), .B2(n9006), .A(n9005), .ZN(n9007) );
  NOR2_X1 U10374 ( .A1(n9007), .A2(n9071), .ZN(n9012) );
  OAI22_X1 U10375 ( .A1(n9010), .A2(n9076), .B1(n9009), .B2(n9074), .ZN(n9011)
         );
  AOI21_X1 U10376 ( .B1(n9012), .B2(n9008), .A(n9011), .ZN(n9152) );
  NOR2_X1 U10377 ( .A1(n9152), .A2(n10070), .ZN(n9013) );
  AOI211_X1 U10378 ( .C1(n9150), .C2(n9088), .A(n9014), .B(n9013), .ZN(n9015)
         );
  OAI21_X1 U10379 ( .B1(n9153), .B2(n9126), .A(n9015), .ZN(P2_U3272) );
  OAI21_X1 U10380 ( .B1(n9018), .B2(n9017), .A(n9016), .ZN(n9158) );
  AOI21_X1 U10381 ( .B1(n9154), .B2(n9043), .A(n9019), .ZN(n9155) );
  INV_X1 U10382 ( .A(n9020), .ZN(n9021) );
  AOI22_X1 U10383 ( .A1(P2_REG2_REG_23__SCAN_IN), .A2(n10070), .B1(n9021), 
        .B2(n10062), .ZN(n9022) );
  OAI21_X1 U10384 ( .B1(n9023), .B2(n10054), .A(n9022), .ZN(n9031) );
  AND2_X1 U10385 ( .A1(n9034), .A2(n9024), .ZN(n9027) );
  OAI21_X1 U10386 ( .B1(n9027), .B2(n9026), .A(n9025), .ZN(n9029) );
  AOI222_X1 U10387 ( .A1(n10049), .A2(n9029), .B1(n9063), .B2(n10045), .C1(
        n9028), .C2(n10046), .ZN(n9157) );
  NOR2_X1 U10388 ( .A1(n9157), .A2(n10070), .ZN(n9030) );
  AOI211_X1 U10389 ( .C1(n9155), .C2(n9088), .A(n9031), .B(n9030), .ZN(n9032)
         );
  OAI21_X1 U10390 ( .B1(n9126), .B2(n9158), .A(n9032), .ZN(P2_U3273) );
  XNOR2_X1 U10391 ( .A(n9033), .B(n9036), .ZN(n9163) );
  NAND2_X1 U10392 ( .A1(n9034), .A2(n10049), .ZN(n9042) );
  AOI21_X1 U10393 ( .B1(n9035), .B2(n9037), .A(n9036), .ZN(n9041) );
  AOI22_X1 U10394 ( .A1(n9039), .A2(n10046), .B1(n10045), .B2(n9038), .ZN(
        n9040) );
  OAI21_X1 U10395 ( .B1(n9042), .B2(n9041), .A(n9040), .ZN(n9159) );
  INV_X1 U10396 ( .A(n9043), .ZN(n9044) );
  AOI211_X1 U10397 ( .C1(n9161), .C2(n9052), .A(n10055), .B(n9044), .ZN(n9160)
         );
  NAND2_X1 U10398 ( .A1(n9160), .A2(n9124), .ZN(n9047) );
  AOI22_X1 U10399 ( .A1(n10070), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9045), 
        .B2(n10062), .ZN(n9046) );
  OAI211_X1 U10400 ( .C1(n4490), .C2(n10054), .A(n9047), .B(n9046), .ZN(n9048)
         );
  AOI21_X1 U10401 ( .B1(n9159), .B2(n9049), .A(n9048), .ZN(n9050) );
  OAI21_X1 U10402 ( .B1(n9163), .B2(n9126), .A(n9050), .ZN(P2_U3274) );
  XOR2_X1 U10403 ( .A(n9060), .B(n9051), .Z(n9168) );
  INV_X1 U10404 ( .A(n9052), .ZN(n9053) );
  AOI21_X1 U10405 ( .B1(n9164), .B2(n4494), .A(n9053), .ZN(n9165) );
  INV_X1 U10406 ( .A(n9054), .ZN(n9055) );
  AOI22_X1 U10407 ( .A1(n10070), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9055), 
        .B2(n10062), .ZN(n9056) );
  OAI21_X1 U10408 ( .B1(n9057), .B2(n10054), .A(n9056), .ZN(n9066) );
  AND2_X1 U10409 ( .A1(n9058), .A2(n9059), .ZN(n9061) );
  OAI21_X1 U10410 ( .B1(n9061), .B2(n9060), .A(n9035), .ZN(n9064) );
  AOI222_X1 U10411 ( .A1(n10049), .A2(n9064), .B1(n9063), .B2(n10046), .C1(
        n9062), .C2(n10045), .ZN(n9167) );
  NOR2_X1 U10412 ( .A1(n9167), .A2(n10070), .ZN(n9065) );
  AOI211_X1 U10413 ( .C1(n9165), .C2(n9088), .A(n9066), .B(n9065), .ZN(n9067)
         );
  OAI21_X1 U10414 ( .B1(n9126), .B2(n9168), .A(n9067), .ZN(P2_U3275) );
  INV_X1 U10415 ( .A(n9058), .ZN(n9073) );
  AOI21_X1 U10416 ( .B1(n9068), .B2(n9070), .A(n9069), .ZN(n9072) );
  NOR3_X1 U10417 ( .A1(n9073), .A2(n9072), .A3(n9071), .ZN(n9079) );
  OAI22_X1 U10418 ( .A1(n9077), .A2(n9076), .B1(n9075), .B2(n9074), .ZN(n9078)
         );
  NOR2_X1 U10419 ( .A1(n9079), .A2(n9078), .ZN(n9174) );
  OR2_X1 U10420 ( .A1(n9081), .A2(n9080), .ZN(n9170) );
  NAND3_X1 U10421 ( .A1(n9170), .A2(n9169), .A3(n9082), .ZN(n9090) );
  AOI21_X1 U10422 ( .B1(n9171), .B2(n9093), .A(n9083), .ZN(n9172) );
  AOI22_X1 U10423 ( .A1(n10070), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9084), 
        .B2(n10062), .ZN(n9085) );
  OAI21_X1 U10424 ( .B1(n9086), .B2(n10054), .A(n9085), .ZN(n9087) );
  AOI21_X1 U10425 ( .B1(n9172), .B2(n9088), .A(n9087), .ZN(n9089) );
  OAI211_X1 U10426 ( .C1(n9174), .C2(n10070), .A(n9090), .B(n9089), .ZN(
        P2_U3276) );
  XNOR2_X1 U10427 ( .A(n9092), .B(n9091), .ZN(n9180) );
  INV_X1 U10428 ( .A(n9110), .ZN(n9095) );
  INV_X1 U10429 ( .A(n9093), .ZN(n9094) );
  AOI211_X1 U10430 ( .C1(n9177), .C2(n9095), .A(n10055), .B(n9094), .ZN(n9176)
         );
  INV_X1 U10431 ( .A(n9096), .ZN(n9097) );
  AOI22_X1 U10432 ( .A1(n10070), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n9097), 
        .B2(n10062), .ZN(n9098) );
  OAI21_X1 U10433 ( .B1(n9099), .B2(n10054), .A(n9098), .ZN(n9106) );
  OAI21_X1 U10434 ( .B1(n9101), .B2(n9100), .A(n9068), .ZN(n9104) );
  INV_X1 U10435 ( .A(n9102), .ZN(n9103) );
  AOI21_X1 U10436 ( .B1(n9104), .B2(n10049), .A(n9103), .ZN(n9179) );
  NOR2_X1 U10437 ( .A1(n9179), .A2(n10070), .ZN(n9105) );
  AOI211_X1 U10438 ( .C1(n9176), .C2(n9124), .A(n9106), .B(n9105), .ZN(n9107)
         );
  OAI21_X1 U10439 ( .B1(n9126), .B2(n9180), .A(n9107), .ZN(P2_U3277) );
  XNOR2_X1 U10440 ( .A(n9108), .B(n9118), .ZN(n9185) );
  INV_X1 U10441 ( .A(n9109), .ZN(n9111) );
  AOI211_X1 U10442 ( .C1(n9182), .C2(n9111), .A(n10055), .B(n9110), .ZN(n9181)
         );
  INV_X1 U10443 ( .A(n9112), .ZN(n9113) );
  AOI22_X1 U10444 ( .A1(n10070), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9113), 
        .B2(n10062), .ZN(n9114) );
  OAI21_X1 U10445 ( .B1(n9115), .B2(n10054), .A(n9114), .ZN(n9123) );
  OAI21_X1 U10446 ( .B1(n9118), .B2(n9117), .A(n9116), .ZN(n9121) );
  AOI222_X1 U10447 ( .A1(n10049), .A2(n9121), .B1(n9120), .B2(n10046), .C1(
        n9119), .C2(n10045), .ZN(n9184) );
  NOR2_X1 U10448 ( .A1(n9184), .A2(n10070), .ZN(n9122) );
  AOI211_X1 U10449 ( .C1(n9181), .C2(n9124), .A(n9123), .B(n9122), .ZN(n9125)
         );
  OAI21_X1 U10450 ( .B1(n9185), .B2(n9126), .A(n9125), .ZN(P2_U3278) );
  AOI22_X1 U10451 ( .A1(n9128), .A2(n5952), .B1(n10142), .B2(n9127), .ZN(n9129) );
  OAI211_X1 U10452 ( .C1(n9131), .C2(n10146), .A(n9130), .B(n9129), .ZN(n9197)
         );
  MUX2_X1 U10453 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9197), .S(n10176), .Z(
        P2_U3549) );
  MUX2_X1 U10454 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9132), .S(n10176), .Z(
        P2_U3548) );
  AOI211_X1 U10455 ( .C1(n10142), .C2(n9135), .A(n9134), .B(n9133), .ZN(n9136)
         );
  OAI21_X1 U10456 ( .B1(n9137), .B2(n10146), .A(n9136), .ZN(n9198) );
  MUX2_X1 U10457 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9198), .S(n10176), .Z(
        P2_U3547) );
  INV_X1 U10458 ( .A(n9138), .ZN(n9143) );
  AOI21_X1 U10459 ( .B1(n10142), .B2(n9140), .A(n9139), .ZN(n9141) );
  OAI211_X1 U10460 ( .C1(n9143), .C2(n10146), .A(n9142), .B(n9141), .ZN(n9199)
         );
  MUX2_X1 U10461 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9199), .S(n10176), .Z(
        P2_U3546) );
  AOI211_X1 U10462 ( .C1(n10142), .C2(n9146), .A(n9145), .B(n9144), .ZN(n9147)
         );
  OAI21_X1 U10463 ( .B1(n9148), .B2(n10146), .A(n9147), .ZN(n9200) );
  MUX2_X1 U10464 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9200), .S(n10176), .Z(
        P2_U3545) );
  AOI22_X1 U10465 ( .A1(n9150), .A2(n5952), .B1(n10142), .B2(n9149), .ZN(n9151) );
  OAI211_X1 U10466 ( .C1(n9153), .C2(n10146), .A(n9152), .B(n9151), .ZN(n9201)
         );
  MUX2_X1 U10467 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9201), .S(n10176), .Z(
        P2_U3544) );
  AOI22_X1 U10468 ( .A1(n9155), .A2(n5952), .B1(n10142), .B2(n9154), .ZN(n9156) );
  OAI211_X1 U10469 ( .C1(n9158), .C2(n10146), .A(n9157), .B(n9156), .ZN(n9202)
         );
  MUX2_X1 U10470 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9202), .S(n10176), .Z(
        P2_U3543) );
  AOI211_X1 U10471 ( .C1(n10142), .C2(n9161), .A(n9160), .B(n9159), .ZN(n9162)
         );
  OAI21_X1 U10472 ( .B1(n9163), .B2(n10146), .A(n9162), .ZN(n9203) );
  MUX2_X1 U10473 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9203), .S(n10176), .Z(
        P2_U3542) );
  AOI22_X1 U10474 ( .A1(n9165), .A2(n5952), .B1(n10142), .B2(n9164), .ZN(n9166) );
  OAI211_X1 U10475 ( .C1(n9168), .C2(n10146), .A(n9167), .B(n9166), .ZN(n9204)
         );
  MUX2_X1 U10476 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9204), .S(n10176), .Z(
        P2_U3541) );
  NAND3_X1 U10477 ( .A1(n9170), .A2(n9169), .A3(n10155), .ZN(n9175) );
  AOI22_X1 U10478 ( .A1(n9172), .A2(n5952), .B1(n10142), .B2(n9171), .ZN(n9173) );
  NAND3_X1 U10479 ( .A1(n9175), .A2(n9174), .A3(n9173), .ZN(n9205) );
  MUX2_X1 U10480 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9205), .S(n10176), .Z(
        P2_U3540) );
  AOI21_X1 U10481 ( .B1(n10142), .B2(n9177), .A(n9176), .ZN(n9178) );
  OAI211_X1 U10482 ( .C1(n9180), .C2(n10146), .A(n9179), .B(n9178), .ZN(n9206)
         );
  MUX2_X1 U10483 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9206), .S(n10176), .Z(
        P2_U3539) );
  AOI21_X1 U10484 ( .B1(n10142), .B2(n9182), .A(n9181), .ZN(n9183) );
  OAI211_X1 U10485 ( .C1(n10146), .C2(n9185), .A(n9184), .B(n9183), .ZN(n9207)
         );
  MUX2_X1 U10486 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9207), .S(n10176), .Z(
        P2_U3538) );
  AOI211_X1 U10487 ( .C1(n10142), .C2(n9188), .A(n9187), .B(n9186), .ZN(n9189)
         );
  OAI21_X1 U10488 ( .B1(n10146), .B2(n9190), .A(n9189), .ZN(n9208) );
  MUX2_X1 U10489 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9208), .S(n10176), .Z(
        P2_U3537) );
  OAI22_X1 U10490 ( .A1(n9192), .A2(n10133), .B1(n4496), .B2(n10150), .ZN(
        n9194) );
  AOI211_X1 U10491 ( .C1(n9195), .C2(n10155), .A(n9194), .B(n9193), .ZN(n9196)
         );
  INV_X1 U10492 ( .A(n9196), .ZN(n9209) );
  MUX2_X1 U10493 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9209), .S(n10176), .Z(
        P2_U3536) );
  MUX2_X1 U10494 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9197), .S(n10158), .Z(
        P2_U3517) );
  MUX2_X1 U10495 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9198), .S(n10158), .Z(
        P2_U3515) );
  MUX2_X1 U10496 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9199), .S(n10158), .Z(
        P2_U3514) );
  MUX2_X1 U10497 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9200), .S(n10158), .Z(
        P2_U3513) );
  MUX2_X1 U10498 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9201), .S(n10158), .Z(
        P2_U3512) );
  MUX2_X1 U10499 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9202), .S(n10158), .Z(
        P2_U3511) );
  MUX2_X1 U10500 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9203), .S(n10158), .Z(
        P2_U3510) );
  MUX2_X1 U10501 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9204), .S(n10158), .Z(
        P2_U3509) );
  MUX2_X1 U10502 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9205), .S(n10158), .Z(
        P2_U3508) );
  MUX2_X1 U10503 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9206), .S(n10158), .Z(
        P2_U3507) );
  MUX2_X1 U10504 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9207), .S(n10158), .Z(
        P2_U3505) );
  MUX2_X1 U10505 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9208), .S(n10158), .Z(
        P2_U3502) );
  MUX2_X1 U10506 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9209), .S(n10158), .Z(
        P2_U3499) );
  INV_X1 U10507 ( .A(n9210), .ZN(n9776) );
  NOR4_X1 U10508 ( .A1(n9211), .A2(P2_IR_REG_30__SCAN_IN), .A3(n5765), .A4(
        P2_U3152), .ZN(n9212) );
  AOI21_X1 U10509 ( .B1(n9218), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9212), .ZN(
        n9213) );
  OAI21_X1 U10510 ( .B1(n9776), .B2(n9221), .A(n9213), .ZN(P2_U3327) );
  AOI22_X1 U10511 ( .A1(n9214), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9218), .ZN(n9215) );
  OAI21_X1 U10512 ( .B1(n9216), .B2(n9221), .A(n9215), .ZN(P2_U3328) );
  INV_X1 U10513 ( .A(n9217), .ZN(n9780) );
  AOI22_X1 U10514 ( .A1(n9219), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9218), .ZN(n9220) );
  OAI21_X1 U10515 ( .B1(n9780), .B2(n9221), .A(n9220), .ZN(P2_U3329) );
  MUX2_X1 U10516 ( .A(n9222), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10517 ( .A(n9224), .B(n9223), .ZN(n9225) );
  XNOR2_X1 U10518 ( .A(n9226), .B(n9225), .ZN(n9232) );
  NOR2_X1 U10519 ( .A1(n9282), .A2(n9405), .ZN(n9230) );
  AOI22_X1 U10520 ( .A1(n9310), .A2(n9647), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n9227) );
  OAI21_X1 U10521 ( .B1(n9228), .B2(n9304), .A(n9227), .ZN(n9229) );
  AOI211_X1 U10522 ( .C1(n5390), .C2(n9320), .A(n9230), .B(n9229), .ZN(n9231)
         );
  OAI21_X1 U10523 ( .B1(n9232), .B2(n9315), .A(n9231), .ZN(P1_U3212) );
  INV_X1 U10524 ( .A(n9233), .ZN(n9235) );
  NAND2_X1 U10525 ( .A1(n9235), .A2(n9234), .ZN(n9237) );
  XNOR2_X1 U10526 ( .A(n9237), .B(n9236), .ZN(n9242) );
  NAND2_X1 U10527 ( .A1(n9648), .A2(n9311), .ZN(n9239) );
  AOI22_X1 U10528 ( .A1(n9310), .A2(n9510), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9238) );
  OAI211_X1 U10529 ( .C1(n9476), .C2(n9282), .A(n9239), .B(n9238), .ZN(n9240)
         );
  AOI21_X1 U10530 ( .B1(n9667), .B2(n9320), .A(n9240), .ZN(n9241) );
  OAI21_X1 U10531 ( .B1(n9242), .B2(n9315), .A(n9241), .ZN(P1_U3214) );
  XOR2_X1 U10532 ( .A(n9244), .B(n9243), .Z(n9249) );
  NAND2_X1 U10533 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9377) );
  OAI21_X1 U10534 ( .B1(n5424), .B2(n9304), .A(n9377), .ZN(n9245) );
  AOI21_X1 U10535 ( .B1(n9323), .B2(n9310), .A(n9245), .ZN(n9246) );
  OAI21_X1 U10536 ( .B1(n9282), .B2(n9540), .A(n9246), .ZN(n9247) );
  AOI21_X1 U10537 ( .B1(n9752), .B2(n9320), .A(n9247), .ZN(n9248) );
  OAI21_X1 U10538 ( .B1(n9249), .B2(n9315), .A(n9248), .ZN(P1_U3217) );
  XOR2_X1 U10539 ( .A(n9251), .B(n9250), .Z(n9258) );
  OAI22_X1 U10540 ( .A1(n9253), .A2(n9304), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9252), .ZN(n9254) );
  AOI21_X1 U10541 ( .B1(n9310), .B2(n9543), .A(n9254), .ZN(n9255) );
  OAI21_X1 U10542 ( .B1(n9282), .B2(n9512), .A(n9255), .ZN(n9256) );
  AOI21_X1 U10543 ( .B1(n9502), .B2(n9320), .A(n9256), .ZN(n9257) );
  OAI21_X1 U10544 ( .B1(n9258), .B2(n9315), .A(n9257), .ZN(P1_U3221) );
  XOR2_X1 U10545 ( .A(n9259), .B(n4344), .Z(n9265) );
  NAND2_X1 U10546 ( .A1(n9648), .A2(n9302), .ZN(n9261) );
  AOI22_X1 U10547 ( .A1(n9311), .A2(n9647), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9260) );
  OAI211_X1 U10548 ( .C1(n9262), .C2(n9441), .A(n9261), .B(n9260), .ZN(n9263)
         );
  AOI21_X1 U10549 ( .B1(n5355), .B2(n9320), .A(n9263), .ZN(n9264) );
  OAI21_X1 U10550 ( .B1(n9265), .B2(n9315), .A(n9264), .ZN(P1_U3223) );
  AOI21_X1 U10551 ( .B1(n9268), .B2(n9267), .A(n9266), .ZN(n9275) );
  OAI22_X1 U10552 ( .A1(n9419), .A2(n9304), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9269), .ZN(n9270) );
  AOI21_X1 U10553 ( .B1(n9306), .B2(n9462), .A(n9270), .ZN(n9271) );
  OAI21_X1 U10554 ( .B1(n9452), .B2(n9272), .A(n9271), .ZN(n9273) );
  AOI21_X1 U10555 ( .B1(n9454), .B2(n9320), .A(n9273), .ZN(n9274) );
  OAI21_X1 U10556 ( .B1(n9275), .B2(n9315), .A(n9274), .ZN(P1_U3227) );
  NAND2_X1 U10557 ( .A1(n9277), .A2(n9276), .ZN(n9278) );
  XOR2_X1 U10558 ( .A(n9279), .B(n9278), .Z(n9285) );
  AOI22_X1 U10559 ( .A1(n9682), .A2(n9311), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9281) );
  NAND2_X1 U10560 ( .A1(n9302), .A2(n9681), .ZN(n9280) );
  OAI211_X1 U10561 ( .C1(n9282), .C2(n9522), .A(n9281), .B(n9280), .ZN(n9283)
         );
  AOI21_X1 U10562 ( .B1(n9533), .B2(n9320), .A(n9283), .ZN(n9284) );
  OAI21_X1 U10563 ( .B1(n9285), .B2(n9315), .A(n9284), .ZN(P1_U3231) );
  INV_X1 U10564 ( .A(n9286), .ZN(n9292) );
  OAI21_X1 U10565 ( .B1(n9287), .B2(n9290), .A(n9288), .ZN(n9291) );
  INV_X1 U10566 ( .A(n9288), .ZN(n9289) );
  AOI22_X1 U10567 ( .A1(n9292), .A2(n9291), .B1(n9290), .B2(n9289), .ZN(n9297)
         );
  NAND2_X1 U10568 ( .A1(n9657), .A2(n9311), .ZN(n9294) );
  AOI22_X1 U10569 ( .A1(n9682), .A2(n9302), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9293) );
  OAI211_X1 U10570 ( .C1(n9262), .C2(n9492), .A(n9294), .B(n9293), .ZN(n9295)
         );
  AOI21_X1 U10571 ( .B1(n9491), .B2(n9320), .A(n9295), .ZN(n9296) );
  OAI21_X1 U10572 ( .B1(n9297), .B2(n9315), .A(n9296), .ZN(P1_U3233) );
  NAND2_X1 U10573 ( .A1(n9299), .A2(n9298), .ZN(n9300) );
  XOR2_X1 U10574 ( .A(n9301), .B(n9300), .Z(n9309) );
  NAND2_X1 U10575 ( .A1(n9302), .A2(n9604), .ZN(n9303) );
  NAND2_X1 U10576 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9912) );
  OAI211_X1 U10577 ( .C1(n9556), .C2(n9304), .A(n9303), .B(n9912), .ZN(n9305)
         );
  AOI21_X1 U10578 ( .B1(n9306), .B2(n9557), .A(n9305), .ZN(n9308) );
  NAND2_X1 U10579 ( .A1(n9566), .A2(n9320), .ZN(n9307) );
  OAI211_X1 U10580 ( .C1(n9309), .C2(n9315), .A(n9308), .B(n9307), .ZN(
        P1_U3236) );
  AOI22_X1 U10581 ( .A1(n9656), .A2(n9310), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9313) );
  NAND2_X1 U10582 ( .A1(n9395), .A2(n9311), .ZN(n9312) );
  OAI211_X1 U10583 ( .C1(n9262), .C2(n9428), .A(n9313), .B(n9312), .ZN(n9319)
         );
  AOI211_X1 U10584 ( .C1(n9317), .C2(n9316), .A(n9315), .B(n9314), .ZN(n9318)
         );
  AOI211_X1 U10585 ( .C1(n9320), .C2(n9427), .A(n9319), .B(n9318), .ZN(n9321)
         );
  INV_X1 U10586 ( .A(n9321), .ZN(P1_U3238) );
  MUX2_X1 U10587 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9322), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10588 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n8396), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10589 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9395), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10590 ( .A(n9647), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9330), .Z(
        P1_U3581) );
  MUX2_X1 U10591 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9656), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10592 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9648), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10593 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9657), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10594 ( .A(n9510), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9330), .Z(
        P1_U3577) );
  MUX2_X1 U10595 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9682), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10596 ( .A(n9543), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9330), .Z(
        P1_U3575) );
  MUX2_X1 U10597 ( .A(n9681), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9330), .Z(
        P1_U3574) );
  MUX2_X1 U10598 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9323), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10599 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9604), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10600 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9616), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10601 ( .A(n9324), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9330), .Z(
        P1_U3570) );
  MUX2_X1 U10602 ( .A(n9615), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9330), .Z(
        P1_U3569) );
  MUX2_X1 U10603 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9854), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10604 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9838), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10605 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9855), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10606 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9983), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10607 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9975), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10608 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9984), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10609 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9976), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10610 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9325), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10611 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9326), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10612 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9327), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10613 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9328), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10614 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9329), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10615 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6423), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10616 ( .A(n9331), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9330), .Z(
        P1_U3555) );
  OAI21_X1 U10617 ( .B1(n9334), .B2(n9333), .A(n9332), .ZN(n9335) );
  NAND2_X1 U10618 ( .A1(n9335), .A2(n9920), .ZN(n9346) );
  INV_X1 U10619 ( .A(n9336), .ZN(n9339) );
  NOR2_X1 U10620 ( .A1(n9914), .A2(n9337), .ZN(n9338) );
  AOI211_X1 U10621 ( .C1(P1_ADDR_REG_11__SCAN_IN), .C2(n9882), .A(n9339), .B(
        n9338), .ZN(n9345) );
  OAI21_X1 U10622 ( .B1(n9342), .B2(n9341), .A(n9340), .ZN(n9343) );
  NAND2_X1 U10623 ( .A1(n9343), .A2(n9911), .ZN(n9344) );
  NAND3_X1 U10624 ( .A1(n9346), .A2(n9345), .A3(n9344), .ZN(P1_U3252) );
  INV_X1 U10625 ( .A(n9367), .ZN(n9353) );
  XNOR2_X1 U10626 ( .A(n9367), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9349) );
  AOI21_X1 U10627 ( .B1(n9355), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9347), .ZN(
        n9348) );
  NOR2_X1 U10628 ( .A1(n9348), .A2(n9349), .ZN(n9366) );
  AOI21_X1 U10629 ( .B1(n9349), .B2(n9348), .A(n9366), .ZN(n9350) );
  NAND2_X1 U10630 ( .A1(n9920), .A2(n9350), .ZN(n9351) );
  OAI211_X1 U10631 ( .C1(n9914), .C2(n9353), .A(n9352), .B(n9351), .ZN(n9360)
         );
  AOI21_X1 U10632 ( .B1(n9355), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9354), .ZN(
        n9358) );
  NAND2_X1 U10633 ( .A1(n9367), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9356) );
  OAI21_X1 U10634 ( .B1(n9367), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9356), .ZN(
        n9357) );
  NOR2_X1 U10635 ( .A1(n9358), .A2(n9357), .ZN(n9362) );
  AOI211_X1 U10636 ( .C1(n9358), .C2(n9357), .A(n9362), .B(n9895), .ZN(n9359)
         );
  AOI211_X1 U10637 ( .C1(P1_ADDR_REG_17__SCAN_IN), .C2(n9882), .A(n9360), .B(
        n9359), .ZN(n9361) );
  INV_X1 U10638 ( .A(n9361), .ZN(P1_U3258) );
  INV_X1 U10639 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9379) );
  OR2_X1 U10640 ( .A1(n9368), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9364) );
  NAND2_X1 U10641 ( .A1(n9368), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9363) );
  NAND2_X1 U10642 ( .A1(n9364), .A2(n9363), .ZN(n9909) );
  INV_X1 U10643 ( .A(n9374), .ZN(n9372) );
  INV_X1 U10644 ( .A(n9365), .ZN(n9886) );
  INV_X1 U10645 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9702) );
  AOI22_X1 U10646 ( .A1(n9368), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n9702), .B2(
        n9915), .ZN(n9918) );
  AOI21_X1 U10647 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9367), .A(n9366), .ZN(
        n9919) );
  NAND2_X1 U10648 ( .A1(n9918), .A2(n9919), .ZN(n9917) );
  OAI21_X1 U10649 ( .B1(n9368), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9917), .ZN(
        n9370) );
  XOR2_X1 U10650 ( .A(n9370), .B(n9369), .Z(n9373) );
  OAI21_X1 U10651 ( .B1(n9373), .B2(n9876), .A(n9914), .ZN(n9371) );
  AOI21_X1 U10652 ( .B1(n9372), .B2(n9886), .A(n9371), .ZN(n9376) );
  AOI22_X1 U10653 ( .A1(n9374), .A2(n9911), .B1(n9920), .B2(n9373), .ZN(n9375)
         );
  MUX2_X1 U10654 ( .A(n9376), .B(n9375), .S(n9408), .Z(n9378) );
  OAI211_X1 U10655 ( .C1(n9379), .C2(n9924), .A(n9378), .B(n9377), .ZN(
        P1_U3260) );
  XNOR2_X1 U10656 ( .A(n9731), .B(n9380), .ZN(n9381) );
  NAND2_X1 U10657 ( .A1(n9635), .A2(n9850), .ZN(n9384) );
  NOR2_X1 U10658 ( .A1(n9382), .A2(n9939), .ZN(n9387) );
  AOI21_X1 U10659 ( .B1(n9939), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9387), .ZN(
        n9383) );
  OAI211_X1 U10660 ( .C1(n9731), .C2(n9628), .A(n9384), .B(n9383), .ZN(
        P1_U3261) );
  NOR2_X1 U10661 ( .A1(n9385), .A2(n9628), .ZN(n9386) );
  AOI211_X1 U10662 ( .C1(n9939), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9387), .B(
        n9386), .ZN(n9388) );
  OAI21_X1 U10663 ( .B1(n9530), .B2(n9389), .A(n9388), .ZN(P1_U3262) );
  INV_X1 U10664 ( .A(n9390), .ZN(n9404) );
  NAND2_X1 U10665 ( .A1(n9391), .A2(n9595), .ZN(n9403) );
  OAI22_X1 U10666 ( .A1(n9620), .A2(n9393), .B1(n9392), .B2(n9598), .ZN(n9394)
         );
  AOI21_X1 U10667 ( .B1(n9525), .B2(n9395), .A(n9394), .ZN(n9396) );
  OAI21_X1 U10668 ( .B1(n9397), .B2(n9527), .A(n9396), .ZN(n9400) );
  NOR2_X1 U10669 ( .A1(n9398), .A2(n9530), .ZN(n9399) );
  AOI211_X1 U10670 ( .C1(n9844), .C2(n9401), .A(n9400), .B(n9399), .ZN(n9402)
         );
  OAI211_X1 U10671 ( .C1(n9404), .C2(n9611), .A(n9403), .B(n9402), .ZN(
        P1_U3263) );
  NOR2_X1 U10672 ( .A1(n9598), .A2(n9405), .ZN(n9407) );
  AOI211_X1 U10673 ( .C1(n9409), .C2(n9408), .A(n9407), .B(n9406), .ZN(n9413)
         );
  NAND2_X1 U10674 ( .A1(n9410), .A2(n9595), .ZN(n9412) );
  AOI22_X1 U10675 ( .A1(n5390), .A2(n9844), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9939), .ZN(n9411) );
  OAI211_X1 U10676 ( .C1(n9939), .C2(n9413), .A(n9412), .B(n9411), .ZN(
        P1_U3264) );
  NAND2_X1 U10677 ( .A1(n9415), .A2(n9414), .ZN(n9416) );
  XNOR2_X1 U10678 ( .A(n9416), .B(n9423), .ZN(n9417) );
  NAND2_X1 U10679 ( .A1(n9417), .A2(n9693), .ZN(n9422) );
  OAI22_X1 U10680 ( .A1(n9419), .A2(n9964), .B1(n9418), .B2(n9962), .ZN(n9420)
         );
  INV_X1 U10681 ( .A(n9420), .ZN(n9421) );
  NAND2_X1 U10682 ( .A1(n9422), .A2(n9421), .ZN(n9642) );
  INV_X1 U10683 ( .A(n9642), .ZN(n9434) );
  XNOR2_X1 U10684 ( .A(n9424), .B(n9423), .ZN(n9644) );
  NAND2_X1 U10685 ( .A1(n9644), .A2(n9595), .ZN(n9433) );
  INV_X1 U10686 ( .A(n9425), .ZN(n9426) );
  AOI211_X1 U10687 ( .C1(n9427), .C2(n9439), .A(n9622), .B(n9426), .ZN(n9643)
         );
  INV_X1 U10688 ( .A(n9427), .ZN(n9735) );
  NOR2_X1 U10689 ( .A1(n9735), .A2(n9628), .ZN(n9431) );
  OAI22_X1 U10690 ( .A1(n9601), .A2(n9429), .B1(n9428), .B2(n9598), .ZN(n9430)
         );
  AOI211_X1 U10691 ( .C1(n9643), .C2(n9850), .A(n9431), .B(n9430), .ZN(n9432)
         );
  OAI211_X1 U10692 ( .C1(n9939), .C2(n9434), .A(n9433), .B(n9432), .ZN(
        P1_U3265) );
  XNOR2_X1 U10693 ( .A(n9436), .B(n9435), .ZN(n9655) );
  XNOR2_X1 U10694 ( .A(n9438), .B(n9437), .ZN(n9653) );
  INV_X1 U10695 ( .A(n9611), .ZN(n9549) );
  OAI211_X1 U10696 ( .C1(n9651), .C2(n9460), .A(n9847), .B(n9439), .ZN(n9650)
         );
  NOR2_X1 U10697 ( .A1(n9527), .A2(n9440), .ZN(n9444) );
  OAI22_X1 U10698 ( .A1(n9601), .A2(n9442), .B1(n9441), .B2(n9598), .ZN(n9443)
         );
  AOI211_X1 U10699 ( .C1(n9648), .C2(n9525), .A(n9444), .B(n9443), .ZN(n9446)
         );
  NAND2_X1 U10700 ( .A1(n5355), .A2(n9844), .ZN(n9445) );
  OAI211_X1 U10701 ( .C1(n9650), .C2(n9530), .A(n9446), .B(n9445), .ZN(n9447)
         );
  AOI21_X1 U10702 ( .B1(n9653), .B2(n9549), .A(n9447), .ZN(n9448) );
  OAI21_X1 U10703 ( .B1(n9655), .B2(n9589), .A(n9448), .ZN(P1_U3266) );
  XNOR2_X1 U10704 ( .A(n9450), .B(n9449), .ZN(n9663) );
  INV_X1 U10705 ( .A(n9663), .ZN(n9467) );
  AOI22_X1 U10706 ( .A1(n9605), .A2(n9656), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9939), .ZN(n9451) );
  OAI21_X1 U10707 ( .B1(n9452), .B2(n9597), .A(n9451), .ZN(n9453) );
  AOI21_X1 U10708 ( .B1(n9454), .B2(n9844), .A(n9453), .ZN(n9466) );
  INV_X1 U10709 ( .A(n9455), .ZN(n9459) );
  NAND2_X1 U10710 ( .A1(n9457), .A2(n9456), .ZN(n9458) );
  AOI21_X1 U10711 ( .B1(n9459), .B2(n9458), .A(n9972), .ZN(n9662) );
  OAI21_X1 U10712 ( .B1(n9660), .B2(n9475), .A(n9847), .ZN(n9461) );
  OR2_X1 U10713 ( .A1(n9461), .A2(n9460), .ZN(n9659) );
  INV_X1 U10714 ( .A(n9462), .ZN(n9463) );
  OAI22_X1 U10715 ( .A1(n9659), .A2(n9513), .B1(n9598), .B2(n9463), .ZN(n9464)
         );
  OAI21_X1 U10716 ( .B1(n9662), .B2(n9464), .A(n9620), .ZN(n9465) );
  OAI211_X1 U10717 ( .C1(n9467), .C2(n9589), .A(n9466), .B(n9465), .ZN(
        P1_U3267) );
  XNOR2_X1 U10718 ( .A(n9468), .B(n9471), .ZN(n9669) );
  INV_X1 U10719 ( .A(n9469), .ZN(n9472) );
  OAI211_X1 U10720 ( .C1(n9472), .C2(n9471), .A(n9470), .B(n9693), .ZN(n9474)
         );
  AOI22_X1 U10721 ( .A1(n9648), .A2(n5499), .B1(n9985), .B2(n9510), .ZN(n9473)
         );
  NAND2_X1 U10722 ( .A1(n9474), .A2(n9473), .ZN(n9665) );
  INV_X1 U10723 ( .A(n9667), .ZN(n9480) );
  AOI211_X1 U10724 ( .C1(n9667), .C2(n4849), .A(n9622), .B(n9475), .ZN(n9666)
         );
  NAND2_X1 U10725 ( .A1(n9666), .A2(n9850), .ZN(n9479) );
  INV_X1 U10726 ( .A(n9476), .ZN(n9477) );
  AOI22_X1 U10727 ( .A1(n9477), .A2(n9936), .B1(n9939), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9478) );
  OAI211_X1 U10728 ( .C1(n9480), .C2(n9628), .A(n9479), .B(n9478), .ZN(n9481)
         );
  AOI21_X1 U10729 ( .B1(n9601), .B2(n9665), .A(n9481), .ZN(n9482) );
  OAI21_X1 U10730 ( .B1(n9669), .B2(n9589), .A(n9482), .ZN(P1_U3268) );
  INV_X1 U10731 ( .A(n9488), .ZN(n9483) );
  XNOR2_X1 U10732 ( .A(n9484), .B(n9483), .ZN(n9485) );
  NAND2_X1 U10733 ( .A1(n9485), .A2(n9693), .ZN(n9487) );
  AOI22_X1 U10734 ( .A1(n9657), .A2(n5499), .B1(n9985), .B2(n9682), .ZN(n9486)
         );
  NAND2_X1 U10735 ( .A1(n9487), .A2(n9486), .ZN(n9670) );
  INV_X1 U10736 ( .A(n9670), .ZN(n9498) );
  XOR2_X1 U10737 ( .A(n9489), .B(n9488), .Z(n9672) );
  NAND2_X1 U10738 ( .A1(n9672), .A2(n9595), .ZN(n9497) );
  INV_X1 U10739 ( .A(n4849), .ZN(n9490) );
  AOI211_X1 U10740 ( .C1(n9491), .C2(n9511), .A(n9622), .B(n9490), .ZN(n9671)
         );
  NOR2_X1 U10741 ( .A1(n4621), .A2(n9628), .ZN(n9495) );
  OAI22_X1 U10742 ( .A1(n9601), .A2(n9493), .B1(n9492), .B2(n9598), .ZN(n9494)
         );
  AOI211_X1 U10743 ( .C1(n9671), .C2(n9850), .A(n9495), .B(n9494), .ZN(n9496)
         );
  OAI211_X1 U10744 ( .C1(n9939), .C2(n9498), .A(n9497), .B(n9496), .ZN(
        P1_U3269) );
  XOR2_X1 U10745 ( .A(n9499), .B(n9504), .Z(n9678) );
  INV_X1 U10746 ( .A(n9678), .ZN(n9518) );
  OAI22_X1 U10747 ( .A1(n5424), .A2(n9597), .B1(n9601), .B2(n9500), .ZN(n9501)
         );
  AOI21_X1 U10748 ( .B1(n9502), .B2(n9844), .A(n9501), .ZN(n9517) );
  INV_X1 U10749 ( .A(n9503), .ZN(n9506) );
  OAI21_X1 U10750 ( .B1(n9506), .B2(n9505), .A(n9504), .ZN(n9508) );
  AOI21_X1 U10751 ( .B1(n9508), .B2(n9507), .A(n9972), .ZN(n9509) );
  AOI21_X1 U10752 ( .B1(n5499), .B2(n9510), .A(n9509), .ZN(n9676) );
  INV_X1 U10753 ( .A(n9676), .ZN(n9515) );
  OAI211_X1 U10754 ( .C1(n9745), .C2(n9529), .A(n9511), .B(n9847), .ZN(n9675)
         );
  OAI22_X1 U10755 ( .A1(n9675), .A2(n9513), .B1(n9598), .B2(n9512), .ZN(n9514)
         );
  OAI21_X1 U10756 ( .B1(n9515), .B2(n9514), .A(n9620), .ZN(n9516) );
  OAI211_X1 U10757 ( .C1(n9518), .C2(n9589), .A(n9517), .B(n9516), .ZN(
        P1_U3270) );
  XNOR2_X1 U10758 ( .A(n9519), .B(n9520), .ZN(n9685) );
  XNOR2_X1 U10759 ( .A(n9521), .B(n9520), .ZN(n9687) );
  NAND2_X1 U10760 ( .A1(n9687), .A2(n9595), .ZN(n9535) );
  OAI22_X1 U10761 ( .A1(n9601), .A2(n9523), .B1(n9522), .B2(n9598), .ZN(n9524)
         );
  AOI21_X1 U10762 ( .B1(n9525), .B2(n9681), .A(n9524), .ZN(n9526) );
  OAI21_X1 U10763 ( .B1(n9528), .B2(n9527), .A(n9526), .ZN(n9532) );
  OAI211_X1 U10764 ( .C1(n9749), .C2(n4325), .A(n4622), .B(n9847), .ZN(n9683)
         );
  NOR2_X1 U10765 ( .A1(n9683), .A2(n9530), .ZN(n9531) );
  AOI211_X1 U10766 ( .C1(n9844), .C2(n9533), .A(n9532), .B(n9531), .ZN(n9534)
         );
  OAI211_X1 U10767 ( .C1(n9685), .C2(n9611), .A(n9535), .B(n9534), .ZN(
        P1_U3271) );
  NAND2_X1 U10768 ( .A1(n9537), .A2(n9536), .ZN(n9538) );
  XOR2_X1 U10769 ( .A(n9547), .B(n9538), .Z(n9696) );
  INV_X1 U10770 ( .A(n9539), .ZN(n9564) );
  AOI211_X1 U10771 ( .C1(n9752), .C2(n9564), .A(n9622), .B(n4325), .ZN(n9691)
         );
  NAND2_X1 U10772 ( .A1(n9752), .A2(n9844), .ZN(n9545) );
  OAI22_X1 U10773 ( .A1(n9601), .A2(n9541), .B1(n9540), .B2(n9598), .ZN(n9542)
         );
  AOI21_X1 U10774 ( .B1(n9605), .B2(n9543), .A(n9542), .ZN(n9544) );
  OAI211_X1 U10775 ( .C1(n9690), .C2(n9597), .A(n9545), .B(n9544), .ZN(n9546)
         );
  AOI21_X1 U10776 ( .B1(n9691), .B2(n9850), .A(n9546), .ZN(n9551) );
  XNOR2_X1 U10777 ( .A(n9548), .B(n9547), .ZN(n9694) );
  NAND2_X1 U10778 ( .A1(n9694), .A2(n9549), .ZN(n9550) );
  OAI211_X1 U10779 ( .C1(n9696), .C2(n9589), .A(n9551), .B(n9550), .ZN(
        P1_U3272) );
  NAND2_X1 U10780 ( .A1(n9553), .A2(n9552), .ZN(n9554) );
  XNOR2_X1 U10781 ( .A(n9554), .B(n5228), .ZN(n9555) );
  OAI222_X1 U10782 ( .A1(n9962), .A2(n9556), .B1(n9964), .B2(n9712), .C1(n9972), .C2(n9555), .ZN(n9699) );
  AOI21_X1 U10783 ( .B1(n9557), .B2(n9936), .A(n9699), .ZN(n9571) );
  NAND2_X1 U10784 ( .A1(n9594), .A2(n9558), .ZN(n9560) );
  AND2_X1 U10785 ( .A1(n9560), .A2(n9559), .ZN(n9562) );
  NAND2_X1 U10786 ( .A1(n9562), .A2(n9561), .ZN(n9563) );
  XNOR2_X1 U10787 ( .A(n9563), .B(n5228), .ZN(n9701) );
  NAND2_X1 U10788 ( .A1(n9701), .A2(n9595), .ZN(n9570) );
  AOI21_X1 U10789 ( .B1(n9575), .B2(n9566), .A(n9622), .ZN(n9565) );
  AND2_X1 U10790 ( .A1(n9565), .A2(n9564), .ZN(n9700) );
  INV_X1 U10791 ( .A(n9566), .ZN(n9757) );
  OAI22_X1 U10792 ( .A1(n9757), .A2(n9628), .B1(n9567), .B2(n9601), .ZN(n9568)
         );
  AOI21_X1 U10793 ( .B1(n9700), .B2(n9850), .A(n9568), .ZN(n9569) );
  OAI211_X1 U10794 ( .C1(n9939), .C2(n9571), .A(n9570), .B(n9569), .ZN(
        P1_U3273) );
  NAND2_X1 U10795 ( .A1(n9594), .A2(n9593), .ZN(n9709) );
  NAND2_X1 U10796 ( .A1(n9709), .A2(n9572), .ZN(n9573) );
  XOR2_X1 U10797 ( .A(n9583), .B(n9573), .Z(n9708) );
  INV_X1 U10798 ( .A(n9574), .ZN(n9577) );
  INV_X1 U10799 ( .A(n9575), .ZN(n9576) );
  AOI211_X1 U10800 ( .C1(n9706), .C2(n9577), .A(n9622), .B(n9576), .ZN(n9705)
         );
  NOR2_X1 U10801 ( .A1(n9578), .A2(n9628), .ZN(n9582) );
  OAI22_X1 U10802 ( .A1(n9601), .A2(n9580), .B1(n9579), .B2(n9598), .ZN(n9581)
         );
  AOI211_X1 U10803 ( .C1(n9705), .C2(n9850), .A(n9582), .B(n9581), .ZN(n9588)
         );
  XOR2_X1 U10804 ( .A(n9584), .B(n9583), .Z(n9585) );
  OAI222_X1 U10805 ( .A1(n9962), .A2(n9690), .B1(n9964), .B2(n9586), .C1(n9585), .C2(n9972), .ZN(n9704) );
  NAND2_X1 U10806 ( .A1(n9704), .A2(n9601), .ZN(n9587) );
  OAI211_X1 U10807 ( .C1(n9708), .C2(n9589), .A(n9588), .B(n9587), .ZN(
        P1_U3274) );
  NAND2_X1 U10808 ( .A1(n9591), .A2(n9590), .ZN(n9592) );
  XOR2_X1 U10809 ( .A(n9593), .B(n9592), .Z(n9718) );
  OR2_X1 U10810 ( .A1(n9594), .A2(n9593), .ZN(n9710) );
  NAND3_X1 U10811 ( .A1(n9710), .A2(n9709), .A3(n9595), .ZN(n9610) );
  INV_X1 U10812 ( .A(n9621), .ZN(n9596) );
  AOI211_X1 U10813 ( .C1(n9715), .C2(n9596), .A(n9622), .B(n9574), .ZN(n9713)
         );
  NOR2_X1 U10814 ( .A1(n9597), .A2(n9711), .ZN(n9603) );
  OAI22_X1 U10815 ( .A1(n9601), .A2(n9600), .B1(n9599), .B2(n9598), .ZN(n9602)
         );
  AOI211_X1 U10816 ( .C1(n9605), .C2(n9604), .A(n9603), .B(n9602), .ZN(n9606)
         );
  OAI21_X1 U10817 ( .B1(n9607), .B2(n9628), .A(n9606), .ZN(n9608) );
  AOI21_X1 U10818 ( .B1(n9713), .B2(n9850), .A(n9608), .ZN(n9609) );
  OAI211_X1 U10819 ( .C1(n9718), .C2(n9611), .A(n9610), .B(n9609), .ZN(
        P1_U3275) );
  XNOR2_X1 U10820 ( .A(n9612), .B(n4427), .ZN(n9721) );
  INV_X1 U10821 ( .A(n9721), .ZN(n9633) );
  XNOR2_X1 U10822 ( .A(n9614), .B(n9613), .ZN(n9619) );
  NAND2_X1 U10823 ( .A1(n9721), .A2(n9860), .ZN(n9618) );
  AOI22_X1 U10824 ( .A1(n9616), .A2(n5499), .B1(n9985), .B2(n9615), .ZN(n9617)
         );
  OAI211_X1 U10825 ( .C1(n9972), .C2(n9619), .A(n9618), .B(n9617), .ZN(n9719)
         );
  NAND2_X1 U10826 ( .A1(n9719), .A2(n9620), .ZN(n9631) );
  AOI211_X1 U10827 ( .C1(n9624), .C2(n9623), .A(n9622), .B(n9621), .ZN(n9720)
         );
  INV_X1 U10828 ( .A(n9624), .ZN(n9763) );
  INV_X1 U10829 ( .A(n9625), .ZN(n9626) );
  AOI22_X1 U10830 ( .A1(n9939), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9626), .B2(
        n9936), .ZN(n9627) );
  OAI21_X1 U10831 ( .B1(n9763), .B2(n9628), .A(n9627), .ZN(n9629) );
  AOI21_X1 U10832 ( .B1(n9720), .B2(n9850), .A(n9629), .ZN(n9630) );
  OAI211_X1 U10833 ( .C1(n9633), .C2(n9632), .A(n9631), .B(n9630), .ZN(
        P1_U3276) );
  INV_X1 U10834 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9636) );
  NOR2_X1 U10835 ( .A1(n9635), .A2(n9634), .ZN(n9729) );
  MUX2_X1 U10836 ( .A(n9636), .B(n9729), .S(n10007), .Z(n9637) );
  OAI21_X1 U10837 ( .B1(n9731), .B2(n9728), .A(n9637), .ZN(P1_U3554) );
  INV_X1 U10838 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9639) );
  OAI21_X1 U10839 ( .B1(n9641), .B2(n9728), .A(n9640), .ZN(P1_U3550) );
  MUX2_X1 U10840 ( .A(n9645), .B(n9732), .S(n10007), .Z(n9646) );
  OAI21_X1 U10841 ( .B1(n9735), .B2(n9728), .A(n9646), .ZN(P1_U3549) );
  AOI22_X1 U10842 ( .A1(n9648), .A2(n9985), .B1(n5499), .B2(n9647), .ZN(n9649)
         );
  OAI211_X1 U10843 ( .C1(n9651), .C2(n9988), .A(n9650), .B(n9649), .ZN(n9652)
         );
  AOI21_X1 U10844 ( .B1(n9653), .B2(n9693), .A(n9652), .ZN(n9654) );
  OAI21_X1 U10845 ( .B1(n9655), .B2(n9947), .A(n9654), .ZN(n9736) );
  MUX2_X1 U10846 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9736), .S(n10007), .Z(
        P1_U3548) );
  AOI22_X1 U10847 ( .A1(n9657), .A2(n9985), .B1(n5499), .B2(n9656), .ZN(n9658)
         );
  OAI211_X1 U10848 ( .C1(n9660), .C2(n9988), .A(n9659), .B(n9658), .ZN(n9661)
         );
  AOI211_X1 U10849 ( .C1(n9663), .C2(n9992), .A(n9662), .B(n9661), .ZN(n9664)
         );
  INV_X1 U10850 ( .A(n9664), .ZN(n9737) );
  MUX2_X1 U10851 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9737), .S(n10007), .Z(
        P1_U3547) );
  AOI211_X1 U10852 ( .C1(n9969), .C2(n9667), .A(n9666), .B(n9665), .ZN(n9668)
         );
  OAI21_X1 U10853 ( .B1(n9669), .B2(n9947), .A(n9668), .ZN(n9738) );
  MUX2_X1 U10854 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9738), .S(n10007), .Z(
        P1_U3546) );
  AOI211_X1 U10855 ( .C1(n9672), .C2(n9992), .A(n9671), .B(n9670), .ZN(n9739)
         );
  MUX2_X1 U10856 ( .A(n9673), .B(n9739), .S(n10007), .Z(n9674) );
  OAI21_X1 U10857 ( .B1(n4621), .B2(n9728), .A(n9674), .ZN(P1_U3545) );
  INV_X1 U10858 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9679) );
  OAI211_X1 U10859 ( .C1(n5424), .C2(n9964), .A(n9676), .B(n9675), .ZN(n9677)
         );
  AOI21_X1 U10860 ( .B1(n9678), .B2(n9992), .A(n9677), .ZN(n9742) );
  MUX2_X1 U10861 ( .A(n9679), .B(n9742), .S(n10007), .Z(n9680) );
  OAI21_X1 U10862 ( .B1(n9745), .B2(n9728), .A(n9680), .ZN(P1_U3544) );
  AOI22_X1 U10863 ( .A1(n9682), .A2(n5499), .B1(n9985), .B2(n9681), .ZN(n9684)
         );
  OAI211_X1 U10864 ( .C1(n9685), .C2(n9972), .A(n9684), .B(n9683), .ZN(n9686)
         );
  AOI21_X1 U10865 ( .B1(n9687), .B2(n9992), .A(n9686), .ZN(n9746) );
  MUX2_X1 U10866 ( .A(n9688), .B(n9746), .S(n10007), .Z(n9689) );
  OAI21_X1 U10867 ( .B1(n9749), .B2(n9728), .A(n9689), .ZN(P1_U3543) );
  OAI22_X1 U10868 ( .A1(n9690), .A2(n9964), .B1(n5424), .B2(n9962), .ZN(n9692)
         );
  AOI211_X1 U10869 ( .C1(n9694), .C2(n9693), .A(n9692), .B(n9691), .ZN(n9695)
         );
  OAI21_X1 U10870 ( .B1(n9696), .B2(n9947), .A(n9695), .ZN(n9750) );
  MUX2_X1 U10871 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9750), .S(n10007), .Z(
        n9697) );
  AOI21_X1 U10872 ( .B1(n5490), .B2(n9752), .A(n9697), .ZN(n9698) );
  INV_X1 U10873 ( .A(n9698), .ZN(P1_U3542) );
  AOI211_X1 U10874 ( .C1(n9701), .C2(n9992), .A(n9700), .B(n9699), .ZN(n9754)
         );
  MUX2_X1 U10875 ( .A(n9702), .B(n9754), .S(n10007), .Z(n9703) );
  OAI21_X1 U10876 ( .B1(n9757), .B2(n9728), .A(n9703), .ZN(P1_U3541) );
  AOI211_X1 U10877 ( .C1(n9969), .C2(n9706), .A(n9705), .B(n9704), .ZN(n9707)
         );
  OAI21_X1 U10878 ( .B1(n9708), .B2(n9947), .A(n9707), .ZN(n9758) );
  MUX2_X1 U10879 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9758), .S(n10007), .Z(
        P1_U3540) );
  NAND3_X1 U10880 ( .A1(n9710), .A2(n9992), .A3(n9709), .ZN(n9717) );
  OAI22_X1 U10881 ( .A1(n9712), .A2(n9962), .B1(n9711), .B2(n9964), .ZN(n9714)
         );
  AOI211_X1 U10882 ( .C1(n9969), .C2(n9715), .A(n9714), .B(n9713), .ZN(n9716)
         );
  OAI211_X1 U10883 ( .C1(n9972), .C2(n9718), .A(n9717), .B(n9716), .ZN(n9759)
         );
  MUX2_X1 U10884 ( .A(n9759), .B(P1_REG1_REG_16__SCAN_IN), .S(n10005), .Z(
        P1_U3539) );
  AOI211_X1 U10885 ( .C1(n9954), .C2(n9721), .A(n9720), .B(n9719), .ZN(n9760)
         );
  MUX2_X1 U10886 ( .A(n9722), .B(n9760), .S(n10007), .Z(n9723) );
  OAI21_X1 U10887 ( .B1(n9763), .B2(n9728), .A(n9723), .ZN(P1_U3538) );
  AOI211_X1 U10888 ( .C1(n9726), .C2(n9992), .A(n9725), .B(n9724), .ZN(n9764)
         );
  MUX2_X1 U10889 ( .A(n5139), .B(n9764), .S(n10007), .Z(n9727) );
  OAI21_X1 U10890 ( .B1(n9768), .B2(n9728), .A(n9727), .ZN(P1_U3537) );
  MUX2_X1 U10891 ( .A(n6016), .B(n9729), .S(n9995), .Z(n9730) );
  OAI21_X1 U10892 ( .B1(n9731), .B2(n9767), .A(n9730), .ZN(P1_U3522) );
  INV_X1 U10893 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9733) );
  MUX2_X1 U10894 ( .A(n9733), .B(n9732), .S(n9995), .Z(n9734) );
  OAI21_X1 U10895 ( .B1(n9735), .B2(n9767), .A(n9734), .ZN(P1_U3517) );
  MUX2_X1 U10896 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9736), .S(n9995), .Z(
        P1_U3516) );
  MUX2_X1 U10897 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9737), .S(n9995), .Z(
        P1_U3515) );
  MUX2_X1 U10898 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9738), .S(n9995), .Z(
        P1_U3514) );
  INV_X1 U10899 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9740) );
  MUX2_X1 U10900 ( .A(n9740), .B(n9739), .S(n9995), .Z(n9741) );
  OAI21_X1 U10901 ( .B1(n4621), .B2(n9767), .A(n9741), .ZN(P1_U3513) );
  MUX2_X1 U10902 ( .A(n9743), .B(n9742), .S(n9995), .Z(n9744) );
  OAI21_X1 U10903 ( .B1(n9745), .B2(n9767), .A(n9744), .ZN(P1_U3512) );
  INV_X1 U10904 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9747) );
  MUX2_X1 U10905 ( .A(n9747), .B(n9746), .S(n9995), .Z(n9748) );
  OAI21_X1 U10906 ( .B1(n9749), .B2(n9767), .A(n9748), .ZN(P1_U3511) );
  MUX2_X1 U10907 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9750), .S(n9995), .Z(n9751) );
  AOI21_X1 U10908 ( .B1(n5507), .B2(n9752), .A(n9751), .ZN(n9753) );
  INV_X1 U10909 ( .A(n9753), .ZN(P1_U3510) );
  INV_X1 U10910 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9755) );
  MUX2_X1 U10911 ( .A(n9755), .B(n9754), .S(n9995), .Z(n9756) );
  OAI21_X1 U10912 ( .B1(n9757), .B2(n9767), .A(n9756), .ZN(P1_U3508) );
  MUX2_X1 U10913 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9758), .S(n9995), .Z(
        P1_U3505) );
  MUX2_X1 U10914 ( .A(n9759), .B(P1_REG0_REG_16__SCAN_IN), .S(n9994), .Z(
        P1_U3502) );
  INV_X1 U10915 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9761) );
  MUX2_X1 U10916 ( .A(n9761), .B(n9760), .S(n9995), .Z(n9762) );
  OAI21_X1 U10917 ( .B1(n9763), .B2(n9767), .A(n9762), .ZN(P1_U3499) );
  INV_X1 U10918 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9765) );
  MUX2_X1 U10919 ( .A(n9765), .B(n9764), .S(n9995), .Z(n9766) );
  OAI21_X1 U10920 ( .B1(n9768), .B2(n9767), .A(n9766), .ZN(P1_U3496) );
  INV_X1 U10921 ( .A(n9769), .ZN(n9773) );
  NAND3_X1 U10922 ( .A1(n9770), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n9772) );
  OAI22_X1 U10923 ( .A1(n9773), .A2(n9772), .B1(n6110), .B2(n9771), .ZN(n9774)
         );
  INV_X1 U10924 ( .A(n9774), .ZN(n9775) );
  OAI21_X1 U10925 ( .B1(n9776), .B2(n9781), .A(n9775), .ZN(P1_U3322) );
  OAI222_X1 U10926 ( .A1(n9781), .A2(n9780), .B1(n9779), .B2(P1_U3084), .C1(
        n9778), .C2(n9777), .ZN(P1_U3324) );
  MUX2_X1 U10927 ( .A(n9782), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U10928 ( .A(n9788), .ZN(n9790) );
  AOI211_X1 U10929 ( .C1(n9969), .C2(n9785), .A(n9784), .B(n9783), .ZN(n9786)
         );
  OAI21_X1 U10930 ( .B1(n9788), .B2(n9787), .A(n9786), .ZN(n9789) );
  AOI21_X1 U10931 ( .B1(n9860), .B2(n9790), .A(n9789), .ZN(n9792) );
  INV_X1 U10932 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9791) );
  AOI22_X1 U10933 ( .A1(n9995), .A2(n9792), .B1(n9791), .B2(n9994), .ZN(
        P1_U3484) );
  AOI22_X1 U10934 ( .A1(n10007), .A2(n9792), .B1(n5063), .B2(n10005), .ZN(
        P1_U3533) );
  NOR2_X1 U10935 ( .A1(n9793), .A2(n10055), .ZN(n9794) );
  INV_X1 U10936 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9796) );
  AOI22_X1 U10937 ( .A1(n10176), .A2(n9823), .B1(n9796), .B2(n10174), .ZN(
        P2_U3551) );
  NOR2_X1 U10938 ( .A1(n9797), .A2(n10055), .ZN(n9798) );
  AOI211_X1 U10939 ( .C1(n10142), .C2(n9800), .A(n9799), .B(n9798), .ZN(n9825)
         );
  INV_X1 U10940 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9801) );
  AOI22_X1 U10941 ( .A1(n10176), .A2(n9825), .B1(n9801), .B2(n10174), .ZN(
        P2_U3550) );
  OAI22_X1 U10942 ( .A1(n9802), .A2(n10133), .B1(n5978), .B2(n10150), .ZN(
        n9804) );
  AOI211_X1 U10943 ( .C1(n10155), .C2(n9805), .A(n9804), .B(n9803), .ZN(n9827)
         );
  AOI22_X1 U10944 ( .A1(n10176), .A2(n9827), .B1(n9806), .B2(n10174), .ZN(
        P2_U3535) );
  INV_X1 U10945 ( .A(n9807), .ZN(n9812) );
  OAI22_X1 U10946 ( .A1(n9809), .A2(n10133), .B1(n9808), .B2(n10150), .ZN(
        n9811) );
  AOI211_X1 U10947 ( .C1(n10155), .C2(n9812), .A(n9811), .B(n9810), .ZN(n9829)
         );
  AOI22_X1 U10948 ( .A1(n10176), .A2(n9829), .B1(n9813), .B2(n10174), .ZN(
        P2_U3534) );
  INV_X1 U10949 ( .A(n9814), .ZN(n10138) );
  INV_X1 U10950 ( .A(n9815), .ZN(n9820) );
  OAI22_X1 U10951 ( .A1(n9817), .A2(n10133), .B1(n9816), .B2(n10150), .ZN(
        n9819) );
  AOI211_X1 U10952 ( .C1(n10138), .C2(n9820), .A(n9819), .B(n9818), .ZN(n9831)
         );
  AOI22_X1 U10953 ( .A1(n10176), .A2(n9831), .B1(n9821), .B2(n10174), .ZN(
        P2_U3533) );
  INV_X1 U10954 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9822) );
  AOI22_X1 U10955 ( .A1(n10158), .A2(n9823), .B1(n9822), .B2(n10156), .ZN(
        P2_U3519) );
  INV_X1 U10956 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9824) );
  AOI22_X1 U10957 ( .A1(n10158), .A2(n9825), .B1(n9824), .B2(n10156), .ZN(
        P2_U3518) );
  INV_X1 U10958 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9826) );
  AOI22_X1 U10959 ( .A1(n10158), .A2(n9827), .B1(n9826), .B2(n10156), .ZN(
        P2_U3496) );
  INV_X1 U10960 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9828) );
  AOI22_X1 U10961 ( .A1(n10158), .A2(n9829), .B1(n9828), .B2(n10156), .ZN(
        P2_U3493) );
  INV_X1 U10962 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9830) );
  AOI22_X1 U10963 ( .A1(n10158), .A2(n9831), .B1(n9830), .B2(n10156), .ZN(
        P2_U3490) );
  INV_X1 U10964 ( .A(n9833), .ZN(n9834) );
  AOI21_X1 U10965 ( .B1(n9835), .B2(n9832), .A(n9834), .ZN(n9871) );
  XNOR2_X1 U10966 ( .A(n9837), .B(n9836), .ZN(n9840) );
  AOI22_X1 U10967 ( .A1(n9985), .A2(n9983), .B1(n9838), .B2(n5499), .ZN(n9839)
         );
  OAI21_X1 U10968 ( .B1(n9840), .B2(n9972), .A(n9839), .ZN(n9841) );
  AOI21_X1 U10969 ( .B1(n9871), .B2(n9860), .A(n9841), .ZN(n9868) );
  INV_X1 U10970 ( .A(n9842), .ZN(n9843) );
  AOI222_X1 U10971 ( .A1(n9845), .A2(n9844), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n9939), .C1(n9843), .C2(n9936), .ZN(n9853) );
  INV_X1 U10972 ( .A(n9846), .ZN(n9848) );
  OAI211_X1 U10973 ( .C1(n9867), .C2(n5443), .A(n9848), .B(n9847), .ZN(n9866)
         );
  INV_X1 U10974 ( .A(n9866), .ZN(n9849) );
  AOI22_X1 U10975 ( .A1(n9871), .A2(n9851), .B1(n9850), .B2(n9849), .ZN(n9852)
         );
  OAI211_X1 U10976 ( .C1(n9939), .C2(n9868), .A(n9853), .B(n9852), .ZN(
        P1_U3280) );
  AOI22_X1 U10977 ( .A1(n9855), .A2(n9985), .B1(n5499), .B2(n9854), .ZN(n9858)
         );
  NAND4_X1 U10978 ( .A1(n9859), .A2(n9858), .A3(n9857), .A4(n9856), .ZN(n9864)
         );
  INV_X1 U10979 ( .A(n9860), .ZN(n9861) );
  NOR2_X1 U10980 ( .A1(n9862), .A2(n9861), .ZN(n9863) );
  AOI211_X1 U10981 ( .C1(n9865), .C2(n9954), .A(n9864), .B(n9863), .ZN(n9872)
         );
  AOI22_X1 U10982 ( .A1(n10007), .A2(n9872), .B1(n6443), .B2(n10005), .ZN(
        P1_U3535) );
  OAI21_X1 U10983 ( .B1(n9867), .B2(n9988), .A(n9866), .ZN(n9870) );
  INV_X1 U10984 ( .A(n9868), .ZN(n9869) );
  AOI211_X1 U10985 ( .C1(n9954), .C2(n9871), .A(n9870), .B(n9869), .ZN(n9874)
         );
  AOI22_X1 U10986 ( .A1(n10007), .A2(n9874), .B1(n5079), .B2(n10005), .ZN(
        P1_U3534) );
  AOI22_X1 U10987 ( .A1(n9995), .A2(n9872), .B1(n5105), .B2(n9994), .ZN(
        P1_U3490) );
  INV_X1 U10988 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9873) );
  AOI22_X1 U10989 ( .A1(n9995), .A2(n9874), .B1(n9873), .B2(n9994), .ZN(
        P1_U3487) );
  XOR2_X1 U10990 ( .A(n9875), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  NOR2_X1 U10991 ( .A1(n9914), .A2(n9883), .ZN(n9881) );
  AOI211_X1 U10992 ( .C1(n9879), .C2(n9878), .A(n9877), .B(n9876), .ZN(n9880)
         );
  AOI211_X1 U10993 ( .C1(P1_ADDR_REG_8__SCAN_IN), .C2(n9882), .A(n9881), .B(
        n9880), .ZN(n9891) );
  NAND2_X1 U10994 ( .A1(n9883), .A2(n5022), .ZN(n9884) );
  OAI211_X1 U10995 ( .C1(n9887), .C2(n9884), .A(n9898), .B(n9911), .ZN(n9889)
         );
  NAND3_X1 U10996 ( .A1(n9887), .A2(n9886), .A3(n9885), .ZN(n9888) );
  NAND4_X1 U10997 ( .A1(n9891), .A2(n9890), .A3(n9889), .A4(n9888), .ZN(
        P1_U3249) );
  OAI21_X1 U10998 ( .B1(n9894), .B2(n9893), .A(n9892), .ZN(n9901) );
  AOI211_X1 U10999 ( .C1(n9898), .C2(n9897), .A(n9896), .B(n9895), .ZN(n9899)
         );
  AOI211_X1 U11000 ( .C1(n9920), .C2(n9901), .A(n9900), .B(n9899), .ZN(n9906)
         );
  INV_X1 U11001 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9903) );
  OAI22_X1 U11002 ( .A1(n9924), .A2(n9903), .B1(n9902), .B2(n9914), .ZN(n9904)
         );
  INV_X1 U11003 ( .A(n9904), .ZN(n9905) );
  NAND2_X1 U11004 ( .A1(n9906), .A2(n9905), .ZN(P1_U3250) );
  AOI21_X1 U11005 ( .B1(n9909), .B2(n9908), .A(n9907), .ZN(n9910) );
  NAND2_X1 U11006 ( .A1(n9911), .A2(n9910), .ZN(n9913) );
  OAI211_X1 U11007 ( .C1(n9915), .C2(n9914), .A(n9913), .B(n9912), .ZN(n9916)
         );
  INV_X1 U11008 ( .A(n9916), .ZN(n9923) );
  OAI21_X1 U11009 ( .B1(n9919), .B2(n9918), .A(n9917), .ZN(n9921) );
  NAND2_X1 U11010 ( .A1(n9921), .A2(n9920), .ZN(n9922) );
  OAI211_X1 U11011 ( .C1(n10213), .C2(n9924), .A(n9923), .B(n9922), .ZN(
        P1_U3259) );
  INV_X1 U11012 ( .A(n9925), .ZN(n9926) );
  OR3_X1 U11013 ( .A1(n9927), .A2(n9926), .A3(n9931), .ZN(n9929) );
  NAND2_X1 U11014 ( .A1(n6423), .A2(n5499), .ZN(n9928) );
  NAND2_X1 U11015 ( .A1(n9929), .A2(n9928), .ZN(n9935) );
  INV_X1 U11016 ( .A(n9930), .ZN(n9934) );
  AOI21_X1 U11017 ( .B1(n9932), .B2(n9931), .A(n9935), .ZN(n9997) );
  INV_X1 U11018 ( .A(n9997), .ZN(n9933) );
  OAI21_X1 U11019 ( .B1(n9935), .B2(n9934), .A(n9933), .ZN(n9938) );
  AOI22_X1 U11020 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(n9939), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n9936), .ZN(n9937) );
  OAI21_X1 U11021 ( .B1(n9939), .B2(n9938), .A(n9937), .ZN(P1_U3291) );
  AND2_X1 U11022 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9940), .ZN(P1_U3292) );
  AND2_X1 U11023 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9940), .ZN(P1_U3293) );
  AND2_X1 U11024 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9940), .ZN(P1_U3294) );
  AND2_X1 U11025 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9940), .ZN(P1_U3295) );
  AND2_X1 U11026 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9940), .ZN(P1_U3296) );
  AND2_X1 U11027 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9940), .ZN(P1_U3297) );
  AND2_X1 U11028 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9940), .ZN(P1_U3298) );
  AND2_X1 U11029 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9940), .ZN(P1_U3299) );
  AND2_X1 U11030 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9940), .ZN(P1_U3300) );
  AND2_X1 U11031 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9940), .ZN(P1_U3301) );
  AND2_X1 U11032 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9940), .ZN(P1_U3302) );
  AND2_X1 U11033 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9940), .ZN(P1_U3303) );
  AND2_X1 U11034 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9940), .ZN(P1_U3304) );
  AND2_X1 U11035 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9940), .ZN(P1_U3305) );
  AND2_X1 U11036 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9940), .ZN(P1_U3306) );
  AND2_X1 U11037 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9940), .ZN(P1_U3307) );
  AND2_X1 U11038 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9940), .ZN(P1_U3308) );
  AND2_X1 U11039 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9940), .ZN(P1_U3309) );
  AND2_X1 U11040 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9940), .ZN(P1_U3310) );
  AND2_X1 U11041 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9940), .ZN(P1_U3311) );
  AND2_X1 U11042 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9940), .ZN(P1_U3312) );
  AND2_X1 U11043 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9940), .ZN(P1_U3313) );
  AND2_X1 U11044 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9940), .ZN(P1_U3314) );
  AND2_X1 U11045 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9940), .ZN(P1_U3315) );
  AND2_X1 U11046 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9940), .ZN(P1_U3316) );
  AND2_X1 U11047 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9940), .ZN(P1_U3317) );
  AND2_X1 U11048 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9940), .ZN(P1_U3318) );
  AND2_X1 U11049 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9940), .ZN(P1_U3319) );
  AND2_X1 U11050 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9940), .ZN(P1_U3320) );
  AND2_X1 U11051 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9940), .ZN(P1_U3321) );
  AOI22_X1 U11052 ( .A1(n9995), .A2(n9997), .B1(n4890), .B2(n9994), .ZN(
        P1_U3454) );
  INV_X1 U11053 ( .A(n9941), .ZN(n9946) );
  OAI21_X1 U11054 ( .B1(n9943), .B2(n9988), .A(n9942), .ZN(n9945) );
  AOI211_X1 U11055 ( .C1(n9946), .C2(n9992), .A(n9945), .B(n9944), .ZN(n9999)
         );
  AOI22_X1 U11056 ( .A1(n9995), .A2(n9999), .B1(n4865), .B2(n9994), .ZN(
        P1_U3457) );
  NOR2_X1 U11057 ( .A1(n9948), .A2(n9947), .ZN(n9953) );
  OAI22_X1 U11058 ( .A1(n9965), .A2(n9962), .B1(n9949), .B2(n9988), .ZN(n9950)
         );
  NOR4_X1 U11059 ( .A1(n9953), .A2(n9952), .A3(n9951), .A4(n9950), .ZN(n10000)
         );
  AOI22_X1 U11060 ( .A1(n9995), .A2(n10000), .B1(n4952), .B2(n9994), .ZN(
        P1_U3469) );
  NAND2_X1 U11061 ( .A1(n9955), .A2(n9954), .ZN(n9957) );
  OAI211_X1 U11062 ( .C1(n9958), .C2(n9988), .A(n9957), .B(n9956), .ZN(n9959)
         );
  NOR2_X1 U11063 ( .A1(n9960), .A2(n9959), .ZN(n10001) );
  INV_X1 U11064 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9961) );
  AOI22_X1 U11065 ( .A1(n9995), .A2(n10001), .B1(n9961), .B2(n9994), .ZN(
        P1_U3472) );
  OAI22_X1 U11066 ( .A1(n9965), .A2(n9964), .B1(n9963), .B2(n9962), .ZN(n9967)
         );
  AOI211_X1 U11067 ( .C1(n9969), .C2(n9968), .A(n9967), .B(n9966), .ZN(n9970)
         );
  OAI21_X1 U11068 ( .B1(n9972), .B2(n9971), .A(n9970), .ZN(n9973) );
  AOI21_X1 U11069 ( .B1(n9992), .B2(n9974), .A(n9973), .ZN(n10003) );
  AOI22_X1 U11070 ( .A1(n9995), .A2(n10003), .B1(n4986), .B2(n9994), .ZN(
        P1_U3475) );
  AOI22_X1 U11071 ( .A1(n9976), .A2(n9985), .B1(n5499), .B2(n9975), .ZN(n9977)
         );
  OAI211_X1 U11072 ( .C1(n4623), .C2(n9988), .A(n9978), .B(n9977), .ZN(n9979)
         );
  AOI211_X1 U11073 ( .C1(n9981), .C2(n9992), .A(n9980), .B(n9979), .ZN(n10004)
         );
  INV_X1 U11074 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9982) );
  AOI22_X1 U11075 ( .A1(n9995), .A2(n10004), .B1(n9982), .B2(n9994), .ZN(
        P1_U3478) );
  AOI22_X1 U11076 ( .A1(n9985), .A2(n9984), .B1(n9983), .B2(n5499), .ZN(n9986)
         );
  OAI211_X1 U11077 ( .C1(n9989), .C2(n9988), .A(n9987), .B(n9986), .ZN(n9990)
         );
  AOI211_X1 U11078 ( .C1(n9993), .C2(n9992), .A(n9991), .B(n9990), .ZN(n10006)
         );
  AOI22_X1 U11079 ( .A1(n9995), .A2(n10006), .B1(n5046), .B2(n9994), .ZN(
        P1_U3481) );
  INV_X1 U11080 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9996) );
  AOI22_X1 U11081 ( .A1(n10007), .A2(n9997), .B1(n9996), .B2(n10005), .ZN(
        P1_U3523) );
  AOI22_X1 U11082 ( .A1(n10007), .A2(n9999), .B1(n9998), .B2(n10005), .ZN(
        P1_U3524) );
  AOI22_X1 U11083 ( .A1(n10007), .A2(n10000), .B1(n6157), .B2(n10005), .ZN(
        P1_U3528) );
  AOI22_X1 U11084 ( .A1(n10007), .A2(n10001), .B1(n6212), .B2(n10005), .ZN(
        P1_U3529) );
  INV_X1 U11085 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10002) );
  AOI22_X1 U11086 ( .A1(n10007), .A2(n10003), .B1(n10002), .B2(n10005), .ZN(
        P1_U3530) );
  AOI22_X1 U11087 ( .A1(n10007), .A2(n10004), .B1(n5018), .B2(n10005), .ZN(
        P1_U3531) );
  AOI22_X1 U11088 ( .A1(n10007), .A2(n10006), .B1(n5045), .B2(n10005), .ZN(
        P1_U3532) );
  OR2_X1 U11089 ( .A1(n10009), .A2(n10008), .ZN(n10012) );
  AND2_X1 U11090 ( .A1(n10012), .A2(n10010), .ZN(n10014) );
  NAND2_X1 U11091 ( .A1(n10012), .A2(n10011), .ZN(n10013) );
  OAI21_X1 U11092 ( .B1(n10015), .B2(n10014), .A(n10013), .ZN(n10023) );
  AOI21_X1 U11093 ( .B1(n10018), .B2(n10017), .A(n10016), .ZN(n10019) );
  OAI21_X1 U11094 ( .B1(n10020), .B2(n10105), .A(n10019), .ZN(n10021) );
  AOI21_X1 U11095 ( .B1(n10023), .B2(n10022), .A(n10021), .ZN(n10024) );
  OAI21_X1 U11096 ( .B1(n10026), .B2(n10025), .A(n10024), .ZN(P2_U3241) );
  AOI22_X1 U11097 ( .A1(n10029), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10027), .ZN(n10038) );
  NAND2_X1 U11098 ( .A1(n10029), .A2(n10028), .ZN(n10031) );
  OAI211_X1 U11099 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n10032), .A(n10031), .B(
        n10030), .ZN(n10033) );
  INV_X1 U11100 ( .A(n10033), .ZN(n10036) );
  AOI22_X1 U11101 ( .A1(n10034), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10035) );
  OAI221_X1 U11102 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n10038), .C1(n10037), .C2(
        n10036), .A(n10035), .ZN(P2_U3245) );
  INV_X1 U11103 ( .A(n10039), .ZN(n10051) );
  XNOR2_X1 U11104 ( .A(n10040), .B(n10041), .ZN(n10052) );
  INV_X1 U11105 ( .A(n10052), .ZN(n10096) );
  NAND3_X1 U11106 ( .A1(n6950), .A2(n10042), .A3(n5958), .ZN(n10043) );
  NAND2_X1 U11107 ( .A1(n10044), .A2(n10043), .ZN(n10048) );
  AOI222_X1 U11108 ( .A1(n10049), .A2(n10048), .B1(n10047), .B2(n10046), .C1(
        n6385), .C2(n10045), .ZN(n10093) );
  INV_X1 U11109 ( .A(n10093), .ZN(n10050) );
  AOI21_X1 U11110 ( .B1(n10051), .B2(n10096), .A(n10050), .ZN(n10069) );
  OAI22_X1 U11111 ( .A1(n10094), .A2(n10054), .B1(n10053), .B2(n10052), .ZN(
        n10067) );
  AOI21_X1 U11112 ( .B1(n10057), .B2(n10056), .A(n10055), .ZN(n10059) );
  NAND2_X1 U11113 ( .A1(n10059), .A2(n10058), .ZN(n10092) );
  OR2_X1 U11114 ( .A1(n9049), .A2(n10060), .ZN(n10064) );
  NAND2_X1 U11115 ( .A1(n10062), .A2(n10061), .ZN(n10063) );
  OAI211_X1 U11116 ( .C1(n10065), .C2(n10092), .A(n10064), .B(n10063), .ZN(
        n10066) );
  NOR2_X1 U11117 ( .A1(n10067), .A2(n10066), .ZN(n10068) );
  OAI21_X1 U11118 ( .B1(n10070), .B2(n10069), .A(n10068), .ZN(P2_U3293) );
  AND2_X1 U11119 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10075), .ZN(P2_U3297) );
  AND2_X1 U11120 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10075), .ZN(P2_U3298) );
  AND2_X1 U11121 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10075), .ZN(P2_U3299) );
  AND2_X1 U11122 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10075), .ZN(P2_U3300) );
  AND2_X1 U11123 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10075), .ZN(P2_U3301) );
  AND2_X1 U11124 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10075), .ZN(P2_U3302) );
  AND2_X1 U11125 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10075), .ZN(P2_U3303) );
  AND2_X1 U11126 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10075), .ZN(P2_U3304) );
  AND2_X1 U11127 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10075), .ZN(P2_U3305) );
  AND2_X1 U11128 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10075), .ZN(P2_U3306) );
  AND2_X1 U11129 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10075), .ZN(P2_U3307) );
  AND2_X1 U11130 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10075), .ZN(P2_U3308) );
  AND2_X1 U11131 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10075), .ZN(P2_U3309) );
  AND2_X1 U11132 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10075), .ZN(P2_U3310) );
  AND2_X1 U11133 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10075), .ZN(P2_U3311) );
  AND2_X1 U11134 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10075), .ZN(P2_U3312) );
  AND2_X1 U11135 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10075), .ZN(P2_U3313) );
  AND2_X1 U11136 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10075), .ZN(P2_U3314) );
  AND2_X1 U11137 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10075), .ZN(P2_U3315) );
  AND2_X1 U11138 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10075), .ZN(P2_U3316) );
  AND2_X1 U11139 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10075), .ZN(P2_U3317) );
  AND2_X1 U11140 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10075), .ZN(P2_U3318) );
  AND2_X1 U11141 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10075), .ZN(P2_U3319) );
  AND2_X1 U11142 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10075), .ZN(P2_U3320) );
  AND2_X1 U11143 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10075), .ZN(P2_U3321) );
  AND2_X1 U11144 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10075), .ZN(P2_U3322) );
  AND2_X1 U11145 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10075), .ZN(P2_U3323) );
  AND2_X1 U11146 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10075), .ZN(P2_U3324) );
  AND2_X1 U11147 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10075), .ZN(P2_U3325) );
  AND2_X1 U11148 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10075), .ZN(P2_U3326) );
  AOI22_X1 U11149 ( .A1(n10074), .A2(n10077), .B1(n10073), .B2(n10075), .ZN(
        P2_U3437) );
  AOI22_X1 U11150 ( .A1(n10078), .A2(n10077), .B1(n10076), .B2(n10075), .ZN(
        P2_U3438) );
  INV_X1 U11151 ( .A(n10079), .ZN(n10084) );
  OAI22_X1 U11152 ( .A1(n10082), .A2(n10146), .B1(n10081), .B2(n10080), .ZN(
        n10083) );
  NOR2_X1 U11153 ( .A1(n10084), .A2(n10083), .ZN(n10160) );
  INV_X1 U11154 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10085) );
  AOI22_X1 U11155 ( .A1(n10158), .A2(n10160), .B1(n10085), .B2(n10156), .ZN(
        P2_U3451) );
  OAI22_X1 U11156 ( .A1(n10087), .A2(n10133), .B1(n10086), .B2(n10150), .ZN(
        n10089) );
  AOI211_X1 U11157 ( .C1(n10155), .C2(n10090), .A(n10089), .B(n10088), .ZN(
        n10162) );
  INV_X1 U11158 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10091) );
  AOI22_X1 U11159 ( .A1(n10158), .A2(n10162), .B1(n10091), .B2(n10156), .ZN(
        P2_U3457) );
  OAI211_X1 U11160 ( .C1(n10094), .C2(n10150), .A(n10093), .B(n10092), .ZN(
        n10095) );
  AOI21_X1 U11161 ( .B1(n10155), .B2(n10096), .A(n10095), .ZN(n10163) );
  INV_X1 U11162 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10097) );
  AOI22_X1 U11163 ( .A1(n10158), .A2(n10163), .B1(n10097), .B2(n10156), .ZN(
        P2_U3460) );
  OAI22_X1 U11164 ( .A1(n10099), .A2(n10133), .B1(n10098), .B2(n10150), .ZN(
        n10101) );
  AOI211_X1 U11165 ( .C1(n10155), .C2(n10102), .A(n10101), .B(n10100), .ZN(
        n10164) );
  INV_X1 U11166 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10103) );
  AOI22_X1 U11167 ( .A1(n10158), .A2(n10164), .B1(n10103), .B2(n10156), .ZN(
        P2_U3463) );
  INV_X1 U11168 ( .A(n10104), .ZN(n10110) );
  OAI22_X1 U11169 ( .A1(n10106), .A2(n10133), .B1(n10105), .B2(n10150), .ZN(
        n10109) );
  INV_X1 U11170 ( .A(n10107), .ZN(n10108) );
  AOI211_X1 U11171 ( .C1(n10155), .C2(n10110), .A(n10109), .B(n10108), .ZN(
        n10166) );
  INV_X1 U11172 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10111) );
  AOI22_X1 U11173 ( .A1(n10158), .A2(n10166), .B1(n10111), .B2(n10156), .ZN(
        P2_U3469) );
  OAI22_X1 U11174 ( .A1(n10112), .A2(n10133), .B1(n4503), .B2(n10150), .ZN(
        n10114) );
  AOI211_X1 U11175 ( .C1(n10155), .C2(n10115), .A(n10114), .B(n10113), .ZN(
        n10168) );
  INV_X1 U11176 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10116) );
  AOI22_X1 U11177 ( .A1(n10158), .A2(n10168), .B1(n10116), .B2(n10156), .ZN(
        P2_U3472) );
  INV_X1 U11178 ( .A(n10117), .ZN(n10122) );
  OAI22_X1 U11179 ( .A1(n10119), .A2(n10133), .B1(n10118), .B2(n10150), .ZN(
        n10121) );
  AOI211_X1 U11180 ( .C1(n10138), .C2(n10122), .A(n10121), .B(n10120), .ZN(
        n10170) );
  INV_X1 U11181 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10123) );
  AOI22_X1 U11182 ( .A1(n10158), .A2(n10170), .B1(n10123), .B2(n10156), .ZN(
        P2_U3475) );
  INV_X1 U11183 ( .A(n10124), .ZN(n10129) );
  OAI22_X1 U11184 ( .A1(n10126), .A2(n10133), .B1(n10125), .B2(n10150), .ZN(
        n10128) );
  AOI211_X1 U11185 ( .C1(n10138), .C2(n10129), .A(n10128), .B(n10127), .ZN(
        n10171) );
  INV_X1 U11186 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10130) );
  AOI22_X1 U11187 ( .A1(n10158), .A2(n10171), .B1(n10130), .B2(n10156), .ZN(
        P2_U3478) );
  INV_X1 U11188 ( .A(n10131), .ZN(n10137) );
  OAI22_X1 U11189 ( .A1(n10134), .A2(n10133), .B1(n4506), .B2(n10150), .ZN(
        n10136) );
  AOI211_X1 U11190 ( .C1(n10138), .C2(n10137), .A(n10136), .B(n10135), .ZN(
        n10172) );
  INV_X1 U11191 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10139) );
  AOI22_X1 U11192 ( .A1(n10158), .A2(n10172), .B1(n10139), .B2(n10156), .ZN(
        P2_U3481) );
  AOI21_X1 U11193 ( .B1(n10142), .B2(n10141), .A(n10140), .ZN(n10143) );
  OAI211_X1 U11194 ( .C1(n10146), .C2(n10145), .A(n10144), .B(n10143), .ZN(
        n10147) );
  INV_X1 U11195 ( .A(n10147), .ZN(n10173) );
  INV_X1 U11196 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10148) );
  AOI22_X1 U11197 ( .A1(n10158), .A2(n10173), .B1(n10148), .B2(n10156), .ZN(
        P2_U3484) );
  OAI21_X1 U11198 ( .B1(n10151), .B2(n10150), .A(n10149), .ZN(n10153) );
  AOI211_X1 U11199 ( .C1(n10155), .C2(n10154), .A(n10153), .B(n10152), .ZN(
        n10175) );
  INV_X1 U11200 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10157) );
  AOI22_X1 U11201 ( .A1(n10158), .A2(n10175), .B1(n10157), .B2(n10156), .ZN(
        P2_U3487) );
  INV_X1 U11202 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10159) );
  AOI22_X1 U11203 ( .A1(n10176), .A2(n10160), .B1(n10159), .B2(n10174), .ZN(
        P2_U3520) );
  AOI22_X1 U11204 ( .A1(n10176), .A2(n10162), .B1(n10161), .B2(n10174), .ZN(
        P2_U3522) );
  AOI22_X1 U11205 ( .A1(n10176), .A2(n10163), .B1(n6257), .B2(n10174), .ZN(
        P2_U3523) );
  AOI22_X1 U11206 ( .A1(n10176), .A2(n10164), .B1(n6261), .B2(n10174), .ZN(
        P2_U3524) );
  INV_X1 U11207 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10165) );
  AOI22_X1 U11208 ( .A1(n10176), .A2(n10166), .B1(n10165), .B2(n10174), .ZN(
        P2_U3526) );
  INV_X1 U11209 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10167) );
  AOI22_X1 U11210 ( .A1(n10176), .A2(n10168), .B1(n10167), .B2(n10174), .ZN(
        P2_U3527) );
  INV_X1 U11211 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10169) );
  AOI22_X1 U11212 ( .A1(n10176), .A2(n10170), .B1(n10169), .B2(n10174), .ZN(
        P2_U3528) );
  AOI22_X1 U11213 ( .A1(n10176), .A2(n10171), .B1(n6544), .B2(n10174), .ZN(
        P2_U3529) );
  AOI22_X1 U11214 ( .A1(n10176), .A2(n10172), .B1(n6546), .B2(n10174), .ZN(
        P2_U3530) );
  AOI22_X1 U11215 ( .A1(n10176), .A2(n10173), .B1(n6548), .B2(n10174), .ZN(
        P2_U3531) );
  AOI22_X1 U11216 ( .A1(n10176), .A2(n10175), .B1(n6597), .B2(n10174), .ZN(
        P2_U3532) );
  INV_X1 U11217 ( .A(n10177), .ZN(n10178) );
  NAND2_X1 U11218 ( .A1(n10179), .A2(n10178), .ZN(n10180) );
  XOR2_X1 U11219 ( .A(n10181), .B(n10180), .Z(ADD_1071_U5) );
  XOR2_X1 U11220 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11221 ( .B1(n10184), .B2(n10183), .A(n10182), .ZN(ADD_1071_U56) );
  OAI21_X1 U11222 ( .B1(n10187), .B2(n10186), .A(n10185), .ZN(ADD_1071_U57) );
  OAI21_X1 U11223 ( .B1(n10190), .B2(n10189), .A(n10188), .ZN(ADD_1071_U58) );
  OAI21_X1 U11224 ( .B1(n10193), .B2(n10192), .A(n10191), .ZN(ADD_1071_U59) );
  OAI21_X1 U11225 ( .B1(n10196), .B2(n10195), .A(n10194), .ZN(ADD_1071_U60) );
  OAI21_X1 U11226 ( .B1(n10199), .B2(n10198), .A(n10197), .ZN(ADD_1071_U61) );
  AOI21_X1 U11227 ( .B1(n10202), .B2(n10201), .A(n10200), .ZN(ADD_1071_U62) );
  AOI21_X1 U11228 ( .B1(n10205), .B2(n10204), .A(n10203), .ZN(ADD_1071_U63) );
  XNOR2_X1 U11229 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10207) );
  XNOR2_X1 U11230 ( .A(n10207), .B(n10206), .ZN(ADD_1071_U47) );
  XOR2_X1 U11231 ( .A(n10209), .B(n10208), .Z(ADD_1071_U54) );
  XOR2_X1 U11232 ( .A(n10210), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  OAI21_X1 U11233 ( .B1(n10213), .B2(n10212), .A(n10211), .ZN(n10214) );
  XNOR2_X1 U11234 ( .A(n10214), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11235 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10215), .Z(ADD_1071_U49) );
  XOR2_X1 U11236 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10216), .Z(ADD_1071_U50) );
  AOI21_X1 U11237 ( .B1(n10218), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n10217), .ZN(
        n10219) );
  XOR2_X1 U11238 ( .A(n10219), .B(P1_ADDR_REG_5__SCAN_IN), .Z(ADD_1071_U51) );
  XOR2_X1 U11239 ( .A(n10221), .B(n10220), .Z(ADD_1071_U53) );
  XNOR2_X1 U11240 ( .A(n10223), .B(n10222), .ZN(ADD_1071_U52) );
  XNOR2_X1 U4860 ( .A(n5945), .B(n4527), .ZN(n8242) );
  CLKBUF_X1 U4818 ( .A(n8916), .Z(n4314) );
  AND3_X1 U4842 ( .A1(n5560), .A2(n4839), .A3(n4612), .ZN(n5543) );
  INV_X1 U4851 ( .A(n5546), .ZN(n9219) );
  NAND2_X1 U5955 ( .A1(n5062), .A2(n5061), .ZN(n9785) );
  NAND2_X1 U5973 ( .A1(n4558), .A2(n4557), .ZN(n4874) );
  CLKBUF_X1 U6049 ( .A(n8916), .Z(n4315) );
endmodule

