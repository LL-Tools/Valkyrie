

module b15_C_SARLock_k_128_5 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3445, 
        U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, 
        U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, 
        U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, 
        U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, 
        U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, 
        U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, 
        U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, 
        U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, 
        U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, 
        U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, 
        U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, 
        U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, 
        U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, 
        U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, 
        U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, 
        U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, 
        U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, 
        U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, 
        U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, 
        U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, 
        U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, 
        U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, 
        U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, 
        U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, 
        U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, 
        U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, 
        U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, 
        U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, 
        U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, 
        U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, 
        U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, 
        U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, 
        U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, 
        U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, 
        U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, 
        U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, 
        U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, 
        U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, 
        U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, 
        U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, 
        U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, 
        U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, 
        U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, 
        U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, 
        U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5358, n5359,
         n5360, n5361, n5362, n5363, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983;

  AND2_X1 U3548 ( .A1(n5553), .A2(n5552), .ZN(n5904) );
  OR2_X1 U3549 ( .A1(n5553), .A2(n5500), .ZN(n5505) );
  AND2_X1 U3551 ( .A1(n5356), .A2(n5496), .ZN(n5470) );
  NAND2_X1 U3552 ( .A1(n5373), .A2(n5355), .ZN(n5553) );
  AND2_X2 U3553 ( .A1(n5593), .A2(n5594), .ZN(n5373) );
  NAND2_X1 U3554 ( .A1(n5593), .A2(n4134), .ZN(n5569) );
  OR2_X1 U3555 ( .A1(n5261), .A2(n3979), .ZN(n5332) );
  NAND2_X1 U3556 ( .A1(n5225), .A2(n5226), .ZN(n5224) );
  INV_X1 U3557 ( .A(n4382), .ZN(n5485) );
  CLKBUF_X1 U3559 ( .A(n3346), .Z(n5435) );
  AND2_X1 U3560 ( .A1(n3244), .A2(n4404), .ZN(n3268) );
  CLKBUF_X2 U3561 ( .A(n3327), .Z(n4315) );
  CLKBUF_X2 U3562 ( .A(n3345), .Z(n5438) );
  CLKBUF_X2 U3563 ( .A(n3328), .Z(n4320) );
  CLKBUF_X2 U3564 ( .A(n3329), .Z(n3101) );
  CLKBUF_X2 U3565 ( .A(n3293), .Z(n5427) );
  CLKBUF_X2 U3566 ( .A(n3351), .Z(n5433) );
  CLKBUF_X2 U3567 ( .A(n3294), .Z(n5437) );
  CLKBUF_X2 U3568 ( .A(n4296), .Z(n4218) );
  NAND2_X1 U3569 ( .A1(n3770), .A2(n3241), .ZN(n3563) );
  AND4_X2 U3570 ( .A1(n3197), .A2(n3196), .A3(n3195), .A4(n3194), .ZN(n3658)
         );
  CLKBUF_X2 U3571 ( .A(n3292), .Z(n5428) );
  AND4_X1 U3572 ( .A1(n3189), .A2(n3188), .A3(n3187), .A4(n3186), .ZN(n3195)
         );
  INV_X1 U3573 ( .A(n4025), .ZN(n5502) );
  XNOR2_X1 U3574 ( .A(n4517), .B(n4722), .ZN(n4489) );
  AND2_X1 U3575 ( .A1(n3824), .A2(n3825), .ZN(n5483) );
  OR2_X1 U3576 ( .A1(n5569), .A2(n5586), .ZN(n5584) );
  BUF_X1 U3578 ( .A(n3852), .Z(n5800) );
  AND2_X1 U3579 ( .A1(n6148), .A2(n4258), .ZN(n6133) );
  NAND2_X1 U3581 ( .A1(n5259), .A2(n5260), .ZN(n5310) );
  AOI21_X1 U3582 ( .B1(n5498), .B2(n5553), .A(n5356), .ZN(n5901) );
  INV_X1 U3583 ( .A(n6133), .ZN(n6128) );
  OR2_X1 U3584 ( .A1(n5470), .A2(n4338), .ZN(n5424) );
  OAI21_X1 U3585 ( .B1(n5373), .B2(n5372), .A(n5569), .ZN(n5862) );
  NAND2_X1 U3587 ( .A1(n5167), .A2(n5166), .ZN(n5169) );
  NOR2_X2 U3588 ( .A1(n4355), .A2(n4710), .ZN(n4712) );
  NAND2_X2 U3589 ( .A1(n3382), .A2(n3381), .ZN(n3386) );
  OAI21_X2 U3590 ( .B1(n5313), .B2(n3542), .A(n3541), .ZN(n5290) );
  OAI21_X2 U3591 ( .B1(n5280), .B2(n3536), .A(n3535), .ZN(n5313) );
  AOI21_X1 U3592 ( .B1(n5523), .B2(n3099), .A(n5509), .ZN(n5510) );
  CLKBUF_X2 U3593 ( .A(n6254), .Z(n6259) );
  CLKBUF_X2 U3594 ( .A(n3251), .Z(n4558) );
  INV_X1 U3595 ( .A(n3330), .ZN(n3100) );
  INV_X2 U3597 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3560) );
  OR2_X1 U3598 ( .A1(n5653), .A2(n5477), .ZN(n3814) );
  NAND2_X1 U3599 ( .A1(n5367), .A2(n3548), .ZN(n5774) );
  AOI21_X1 U3600 ( .B1(n5586), .B2(n5569), .A(n5585), .ZN(n5913) );
  NAND2_X1 U3601 ( .A1(n5691), .A2(n3546), .ZN(n5367) );
  AND2_X2 U3603 ( .A1(n5602), .A2(n5603), .ZN(n5593) );
  CLKBUF_X1 U3604 ( .A(n5313), .Z(n5322) );
  NAND2_X1 U3605 ( .A1(n5263), .A2(n5262), .ZN(n5261) );
  AND2_X1 U3606 ( .A1(n5056), .A2(n3930), .ZN(n5210) );
  NAND2_X1 U3607 ( .A1(n3520), .A2(n3519), .ZN(n3521) );
  AND2_X2 U3608 ( .A1(n3525), .A2(n3524), .ZN(n3556) );
  OR2_X2 U3609 ( .A1(n6288), .A2(n4563), .ZN(n6296) );
  XNOR2_X1 U3610 ( .A(n3492), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6283)
         );
  XNOR2_X1 U3611 ( .A(n3412), .B(n3420), .ZN(n3874) );
  NAND2_X1 U3612 ( .A1(n3489), .A2(n3488), .ZN(n3492) );
  CLKBUF_X1 U3613 ( .A(n4526), .Z(n4797) );
  XNOR2_X1 U3614 ( .A(n3449), .B(n3452), .ZN(n4526) );
  NAND2_X1 U3615 ( .A1(n3286), .A2(n3368), .ZN(n4517) );
  CLKBUF_X1 U3616 ( .A(n3840), .Z(n5252) );
  AND2_X1 U3617 ( .A1(n4401), .A2(n4586), .ZN(n4234) );
  NAND2_X2 U3618 ( .A1(n4374), .A2(n4586), .ZN(n3755) );
  AND2_X1 U3619 ( .A1(n3413), .A2(n3658), .ZN(n3783) );
  BUF_X2 U3620 ( .A(n3654), .Z(n4580) );
  NAND2_X1 U3621 ( .A1(n3228), .A2(n3454), .ZN(n3624) );
  CLKBUF_X1 U3622 ( .A(n3454), .Z(n4594) );
  INV_X2 U3623 ( .A(n3654), .ZN(n3241) );
  NAND2_X1 U3624 ( .A1(n4598), .A2(n3227), .ZN(n3245) );
  AND4_X2 U3625 ( .A1(n3113), .A2(n3140), .A3(n3139), .A4(n3138), .ZN(n4373)
         );
  INV_X2 U3626 ( .A(n4586), .ZN(n3770) );
  OR2_X2 U3627 ( .A1(n3150), .A2(n3149), .ZN(n4541) );
  INV_X1 U3628 ( .A(n3227), .ZN(n3454) );
  AND4_X1 U3629 ( .A1(n3181), .A2(n3180), .A3(n3179), .A4(n3178), .ZN(n3197)
         );
  AND4_X1 U3630 ( .A1(n3137), .A2(n3136), .A3(n3135), .A4(n3134), .ZN(n3138)
         );
  AND4_X1 U3631 ( .A1(n3193), .A2(n3192), .A3(n3191), .A4(n3190), .ZN(n3194)
         );
  AND4_X1 U3632 ( .A1(n3185), .A2(n3184), .A3(n3183), .A4(n3182), .ZN(n3196)
         );
  AND4_X1 U3633 ( .A1(n3131), .A2(n3130), .A3(n3129), .A4(n3128), .ZN(n3139)
         );
  INV_X2 U3634 ( .A(n6645), .ZN(n6194) );
  INV_X2 U3635 ( .A(n6266), .ZN(n3099) );
  BUF_X2 U3636 ( .A(n3370), .Z(n3322) );
  CLKBUF_X3 U3637 ( .A(n3169), .Z(n4145) );
  NOR2_X2 U3638 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4490) );
  XNOR2_X2 U3639 ( .A(n3483), .B(n4538), .ZN(n3852) );
  AND3_X2 U3640 ( .A1(n3214), .A2(n3213), .A3(n3212), .ZN(n3219) );
  NOR2_X4 U3641 ( .A1(n5310), .A2(n5311), .ZN(n5309) );
  NAND2_X2 U3642 ( .A1(n3307), .A2(n3306), .ZN(n4538) );
  NAND2_X1 U3643 ( .A1(n3448), .A2(n3447), .ZN(n6291) );
  AOI211_X1 U3645 ( .C1(n6648), .C2(n6735), .A(n6647), .B(n6646), .ZN(n6649)
         );
  INV_X1 U3646 ( .A(n4381), .ZN(n5522) );
  NOR2_X4 U3647 ( .A1(n5384), .A2(n5385), .ZN(n5631) );
  NAND2_X2 U3648 ( .A1(n5309), .A2(n5301), .ZN(n5384) );
  AOI21_X2 U3649 ( .B1(n3545), .B2(n3107), .A(n3106), .ZN(n5691) );
  AOI21_X2 U3650 ( .B1(n4479), .B2(n4478), .A(n3475), .ZN(n6289) );
  AND2_X1 U3651 ( .A1(n3133), .A2(n4407), .ZN(n3102) );
  AND2_X4 U3652 ( .A1(n3132), .A2(n4407), .ZN(n3346) );
  BUF_X4 U3653 ( .A(n3209), .Z(n4314) );
  OR2_X1 U3654 ( .A1(n6532), .A2(n6539), .ZN(n4611) );
  AND2_X1 U3655 ( .A1(n3494), .A2(n3420), .ZN(n3421) );
  NAND3_X1 U3656 ( .A1(n3272), .A2(n3276), .A3(n3275), .ZN(n3309) );
  OR2_X1 U3657 ( .A1(n4586), .A2(n6910), .ZN(n3383) );
  NOR2_X2 U3658 ( .A1(n5609), .A2(n5610), .ZN(n5602) );
  XNOR2_X1 U3659 ( .A(n3496), .B(n3495), .ZN(n3860) );
  NAND2_X1 U3660 ( .A1(n6148), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5513) );
  AND2_X1 U3661 ( .A1(n4116), .A2(n4115), .ZN(n5594) );
  OR2_X1 U3662 ( .A1(n4611), .A2(n5539), .ZN(n6198) );
  NAND2_X1 U3663 ( .A1(n3651), .A2(n3650), .ZN(n3794) );
  AND2_X2 U3664 ( .A1(n3228), .A2(n4381), .ZN(n3261) );
  AND2_X2 U3665 ( .A1(n4399), .A2(n3132), .ZN(n3209) );
  AND2_X1 U3666 ( .A1(n4232), .A2(n5372), .ZN(n4287) );
  INV_X1 U3667 ( .A(n5447), .ZN(n4330) );
  NAND2_X1 U3668 ( .A1(n4472), .A2(n3111), .ZN(n4355) );
  INV_X1 U3669 ( .A(n3833), .ZN(n4025) );
  AND2_X1 U3670 ( .A1(n3755), .A2(n3764), .ZN(n3771) );
  AND2_X1 U3671 ( .A1(n5279), .A2(n3534), .ZN(n3535) );
  XNOR2_X1 U3672 ( .A(n3344), .B(n3310), .ZN(n4400) );
  INV_X1 U3673 ( .A(n3617), .ZN(n3609) );
  INV_X1 U3674 ( .A(n3636), .ZN(n3608) );
  CLKBUF_X1 U3675 ( .A(n3413), .Z(n3567) );
  AND2_X1 U3676 ( .A1(n3615), .A2(n3614), .ZN(n3619) );
  NAND2_X1 U3677 ( .A1(n3337), .A2(n3383), .ZN(n3616) );
  OR2_X1 U3678 ( .A1(n5513), .A2(n4251), .ZN(n6131) );
  INV_X1 U3680 ( .A(n4191), .ZN(n5501) );
  AND2_X1 U3681 ( .A1(n5594), .A2(n5372), .ZN(n4134) );
  XNOR2_X1 U3682 ( .A(n5261), .B(n3979), .ZN(n5307) );
  NAND2_X1 U3683 ( .A1(n4712), .A2(n4960), .ZN(n5058) );
  NOR2_X1 U3684 ( .A1(n6929), .A2(n3875), .ZN(n3882) );
  NAND2_X1 U3685 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n3882), .ZN(n3886)
         );
  NOR2_X1 U3686 ( .A1(n3864), .A2(n6103), .ZN(n3869) );
  NAND2_X1 U3687 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n3869), .ZN(n3875)
         );
  INV_X1 U3689 ( .A(n3556), .ZN(n5406) );
  OR2_X1 U3690 ( .A1(n3653), .A2(n3652), .ZN(n6516) );
  OR3_X1 U3691 ( .A1(n4397), .A2(n4396), .A3(n4395), .ZN(n6499) );
  INV_X1 U3692 ( .A(n3619), .ZN(n3641) );
  NAND2_X1 U3693 ( .A1(n3583), .A2(n3567), .ZN(n3617) );
  AND2_X1 U3694 ( .A1(n3616), .A2(n3619), .ZN(n3618) );
  AND2_X1 U3695 ( .A1(n6198), .A2(n4235), .ZN(n6644) );
  NAND2_X1 U3696 ( .A1(n6133), .A2(n5656), .ZN(n4259) );
  NAND2_X1 U3697 ( .A1(n4380), .A2(n4379), .ZN(n6159) );
  AND2_X1 U3698 ( .A1(n5640), .A2(n5378), .ZN(n6167) );
  AND2_X1 U3699 ( .A1(n5640), .A2(n4613), .ZN(n6168) );
  INV_X1 U3700 ( .A(n5640), .ZN(n6170) );
  XNOR2_X1 U3701 ( .A(n5470), .B(n5469), .ZN(n5894) );
  INV_X1 U3702 ( .A(n5497), .ZN(n5469) );
  XNOR2_X1 U3703 ( .A(n3558), .B(n3557), .ZN(n5476) );
  AOI21_X1 U3704 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5479), .A(n3811), 
        .ZN(n3558) );
  OR2_X1 U3705 ( .A1(n5739), .A2(n3804), .ZN(n5941) );
  INV_X1 U3706 ( .A(n6532), .ZN(n4398) );
  INV_X1 U3707 ( .A(n4598), .ZN(n3228) );
  OR2_X1 U3708 ( .A1(n3336), .A2(n3335), .ZN(n3527) );
  OR2_X1 U3709 ( .A1(n3397), .A2(n3396), .ZN(n3497) );
  OR2_X1 U3710 ( .A1(n3380), .A2(n3379), .ZN(n3414) );
  OR2_X1 U3712 ( .A1(n4558), .A2(n6910), .ZN(n3337) );
  OR3_X1 U3713 ( .A1(n3613), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(n6387), 
        .ZN(n3636) );
  INV_X1 U3714 ( .A(n4287), .ZN(n4288) );
  NOR2_X1 U3715 ( .A1(n4413), .A2(n6910), .ZN(n5447) );
  NAND2_X1 U3716 ( .A1(n3900), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3915)
         );
  INV_X1 U3717 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6929) );
  AND2_X1 U3718 ( .A1(n5378), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3841) );
  NAND2_X1 U3719 ( .A1(n3442), .A2(n3441), .ZN(n3507) );
  OR2_X1 U3720 ( .A1(n3358), .A2(n3357), .ZN(n3466) );
  NAND2_X1 U3721 ( .A1(n3344), .A2(n3343), .ZN(n3840) );
  NAND2_X1 U3722 ( .A1(n3277), .A2(n3309), .ZN(n3369) );
  INV_X1 U3723 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4719) );
  AND4_X1 U3724 ( .A1(n3127), .A2(n3126), .A3(n3125), .A4(n3124), .ZN(n3140)
         );
  OAI21_X1 U3725 ( .B1(n6651), .B2(n4530), .A(n6626), .ZN(n4540) );
  INV_X1 U3726 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6505) );
  INV_X1 U3727 ( .A(n3583), .ZN(n3605) );
  NOR2_X1 U3728 ( .A1(n6110), .A2(n4244), .ZN(n6015) );
  AND2_X1 U3729 ( .A1(n4337), .A2(n4336), .ZN(n5496) );
  OR2_X1 U3730 ( .A1(n5816), .A2(n5449), .ZN(n4336) );
  OR2_X2 U3731 ( .A1(n3168), .A2(n3167), .ZN(n4381) );
  BUF_X1 U3732 ( .A(n5609), .Z(n5628) );
  OR2_X1 U3733 ( .A1(n4282), .A2(n4281), .ZN(n4307) );
  NAND2_X1 U3734 ( .A1(n4204), .A2(n4183), .ZN(n4238) );
  AND2_X1 U3735 ( .A1(n4133), .A2(n4132), .ZN(n5372) );
  NOR2_X1 U3736 ( .A1(n4113), .A2(n5875), .ZN(n4114) );
  CLKBUF_X1 U3737 ( .A(n5602), .Z(n5611) );
  NOR2_X1 U3738 ( .A1(n4079), .A2(n5698), .ZN(n4080) );
  NOR2_X1 U3739 ( .A1(n4045), .A2(n6019), .ZN(n4046) );
  INV_X1 U3740 ( .A(n4044), .ZN(n4045) );
  NAND2_X1 U3742 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n3995), .ZN(n3996)
         );
  BUF_X1 U3743 ( .A(n5395), .Z(n5634) );
  AND3_X1 U3744 ( .A1(n3994), .A2(n3993), .A3(n3992), .ZN(n5333) );
  CLKBUF_X1 U3745 ( .A(n5331), .Z(n5394) );
  NAND2_X1 U3746 ( .A1(n3964), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3991)
         );
  INV_X1 U3747 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6037) );
  INV_X1 U3748 ( .A(n5307), .ZN(n3978) );
  NOR2_X1 U3749 ( .A1(n3949), .A2(n3948), .ZN(n3964) );
  NAND2_X1 U3750 ( .A1(n3931), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3949)
         );
  INV_X1 U3751 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3948) );
  CLKBUF_X1 U3752 ( .A(n5210), .Z(n5215) );
  AOI21_X1 U3753 ( .B1(n3881), .B2(n3988), .A(n3885), .ZN(n4710) );
  CLKBUF_X1 U3754 ( .A(n4712), .Z(n4959) );
  AOI21_X1 U3755 ( .B1(n3874), .B2(n3988), .A(n3873), .ZN(n4616) );
  NAND2_X1 U3756 ( .A1(n3868), .A2(n3867), .ZN(n4469) );
  NAND2_X1 U3757 ( .A1(n3854), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3864)
         );
  NAND2_X1 U3758 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3853) );
  INV_X1 U3759 ( .A(n3771), .ZN(n5486) );
  BUF_X1 U3761 ( .A(n3664), .Z(n5616) );
  NAND2_X1 U3762 ( .A1(n5950), .A2(n5618), .ZN(n5606) );
  CLKBUF_X1 U3763 ( .A(n5691), .Z(n5692) );
  AND2_X1 U3764 ( .A1(n5323), .A2(n3540), .ZN(n3541) );
  OR2_X1 U3765 ( .A1(n5406), .A2(n5388), .ZN(n5288) );
  NAND2_X1 U3766 ( .A1(n4618), .A2(n4357), .ZN(n4714) );
  AND2_X1 U3767 ( .A1(n6395), .A2(n6537), .ZN(n4364) );
  OR2_X1 U3768 ( .A1(n5297), .A2(n5299), .ZN(n6330) );
  CLKBUF_X1 U3769 ( .A(n4400), .Z(n6136) );
  OR2_X1 U3770 ( .A1(n3780), .A2(n4590), .ZN(n4413) );
  AND2_X2 U3771 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4513) );
  NAND2_X1 U3772 ( .A1(n3291), .A2(n3290), .ZN(n4722) );
  NAND2_X1 U3773 ( .A1(n3222), .A2(n3770), .ZN(n3223) );
  AND2_X1 U3774 ( .A1(n4924), .A2(n4865), .ZN(n5109) );
  AND2_X1 U3775 ( .A1(n4718), .A2(n4717), .ZN(n5019) );
  OR2_X1 U3776 ( .A1(n4861), .A2(n4797), .ZN(n4690) );
  INV_X1 U3777 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6647) );
  INV_X1 U3778 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6917) );
  OR2_X1 U3779 ( .A1(n4842), .A2(n5018), .ZN(n4804) );
  NAND2_X1 U3780 ( .A1(n6910), .A2(n4540), .ZN(n4764) );
  OR2_X1 U3781 ( .A1(n4798), .A2(n4797), .ZN(n4842) );
  INV_X1 U3782 ( .A(n5522), .ZN(n4554) );
  AND2_X1 U3783 ( .A1(n6621), .A2(n4540), .ZN(n4599) );
  INV_X1 U3784 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6537) );
  AOI22_X1 U3785 ( .A1(n5910), .A2(n6079), .B1(n5840), .B2(n6083), .ZN(n5843)
         );
  INV_X1 U3786 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U3787 ( .A1(n6644), .A2(n4237), .ZN(n6148) );
  OR2_X1 U3788 ( .A1(n6340), .A2(n6541), .ZN(n4236) );
  INV_X1 U3789 ( .A(n6138), .ZN(n6115) );
  NOR2_X1 U3790 ( .A1(n5483), .A2(n3827), .ZN(n5812) );
  INV_X1 U3791 ( .A(n5904), .ZN(n5567) );
  INV_X1 U3792 ( .A(n5573), .ZN(n5574) );
  OR2_X1 U3793 ( .A1(n5572), .A2(n5571), .ZN(n5575) );
  OR2_X1 U3794 ( .A1(n5596), .A2(n5595), .ZN(n5870) );
  INV_X1 U3795 ( .A(n5601), .ZN(n6156) );
  NAND2_X1 U3796 ( .A1(n6159), .A2(n5522), .ZN(n6150) );
  INV_X2 U3797 ( .A(n6175), .ZN(n6980) );
  OR2_X2 U3798 ( .A1(n4611), .A2(n4605), .ZN(n6261) );
  INV_X1 U3799 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5204) );
  OR2_X1 U3800 ( .A1(n5754), .A2(n3802), .ZN(n5739) );
  NOR2_X1 U3801 ( .A1(n5298), .A2(n6299), .ZN(n5965) );
  OR2_X1 U3802 ( .A1(n5297), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4485)
         );
  NAND2_X1 U3803 ( .A1(n3794), .A2(n3661), .ZN(n6378) );
  INV_X1 U3804 ( .A(n6378), .ZN(n6342) );
  INV_X1 U3805 ( .A(n4797), .ZN(n4717) );
  CLKBUF_X1 U3806 ( .A(n4533), .Z(n4875) );
  CLKBUF_X1 U3807 ( .A(n4501), .Z(n6116) );
  CLKBUF_X1 U3808 ( .A(n4489), .Z(n6107) );
  AND2_X2 U3809 ( .A1(n3117), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4399)
         );
  INV_X1 U3810 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3117) );
  AND2_X1 U3811 ( .A1(n5019), .A2(n5018), .ZN(n6434) );
  OR2_X1 U3812 ( .A1(n4861), .A2(n4874), .ZN(n6495) );
  NAND2_X1 U3813 ( .A1(n4582), .A2(n4581), .ZN(n4835) );
  INV_X1 U3814 ( .A(n5140), .ZN(n6447) );
  INV_X1 U3815 ( .A(n5118), .ZN(n6453) );
  INV_X1 U3816 ( .A(n5145), .ZN(n6481) );
  INV_X1 U3817 ( .A(n5153), .ZN(n6461) );
  INV_X1 U3818 ( .A(n4804), .ZN(n4913) );
  INV_X1 U3819 ( .A(n5130), .ZN(n6489) );
  AND2_X1 U3820 ( .A1(n3644), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6525) );
  NAND2_X1 U3821 ( .A1(n3622), .A2(n3621), .ZN(n6532) );
  OAI21_X1 U3822 ( .B1(n3620), .B2(n3618), .A(n3617), .ZN(n3622) );
  INV_X1 U3823 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6910) );
  INV_X1 U3824 ( .A(n6525), .ZN(n6539) );
  NAND2_X1 U3825 ( .A1(n4260), .A2(n4259), .ZN(n4261) );
  AND2_X1 U3826 ( .A1(n6167), .A2(DATAI_29_), .ZN(n5897) );
  AOI21_X1 U3827 ( .B1(n5894), .B2(n3099), .A(n5474), .ZN(n5475) );
  AND2_X2 U3828 ( .A1(n3132), .A2(n5528), .ZN(n3329) );
  INV_X1 U3829 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3116) );
  NAND2_X1 U3830 ( .A1(n3859), .A2(n3858), .ZN(n4440) );
  OR2_X1 U3831 ( .A1(n4611), .A2(n6516), .ZN(n5984) );
  INV_X1 U3832 ( .A(n6340), .ZN(n6376) );
  AND2_X2 U3833 ( .A1(n5984), .A2(n4341), .ZN(n6288) );
  NAND2_X1 U3834 ( .A1(n3671), .A2(n3670), .ZN(n3103) );
  INV_X1 U3835 ( .A(n5726), .ZN(n4262) );
  AND2_X1 U3836 ( .A1(n3794), .A2(n3657), .ZN(n6381) );
  AND2_X2 U3837 ( .A1(n4490), .A2(n5528), .ZN(n3293) );
  AND2_X2 U3838 ( .A1(n5528), .A2(n4513), .ZN(n3294) );
  INV_X1 U3839 ( .A(n4170), .ZN(n3330) );
  AND4_X1 U3840 ( .A1(n3158), .A2(n3157), .A3(n3156), .A4(n3155), .ZN(n3104)
         );
  NAND2_X1 U3841 ( .A1(n5406), .A2(n5388), .ZN(n3105) );
  AND2_X1 U3842 ( .A1(n5406), .A2(n5790), .ZN(n3106) );
  OR2_X1 U3843 ( .A1(n5693), .A2(n5790), .ZN(n3107) );
  AND3_X1 U3844 ( .A1(n3227), .A2(n4374), .A3(n4373), .ZN(n3108) );
  AND4_X1 U3845 ( .A1(n3154), .A2(n3153), .A3(n3152), .A4(n3151), .ZN(n3109)
         );
  AND4_X1 U3846 ( .A1(n3218), .A2(n3217), .A3(n3216), .A4(n3215), .ZN(n3110)
         );
  NAND2_X1 U3847 ( .A1(n3245), .A2(n3658), .ZN(n3242) );
  AND2_X1 U3848 ( .A1(n3880), .A2(n3879), .ZN(n3111) );
  AND4_X1 U3849 ( .A1(n3173), .A2(n3172), .A3(n3171), .A4(n3170), .ZN(n3112)
         );
  AND4_X1 U3850 ( .A1(n3121), .A2(n3120), .A3(n3119), .A4(n3118), .ZN(n3113)
         );
  NAND2_X1 U3851 ( .A1(n3285), .A2(n3284), .ZN(n3368) );
  AND4_X1 U3852 ( .A1(n3177), .A2(n3176), .A3(n3175), .A4(n3174), .ZN(n3114)
         );
  INV_X1 U3853 ( .A(n6083), .ZN(n6120) );
  AND2_X1 U3854 ( .A1(n5812), .A2(n6083), .ZN(n3115) );
  OR2_X1 U3855 ( .A1(n3565), .A2(n3586), .ZN(n3570) );
  INV_X1 U3856 ( .A(n3242), .ZN(n3243) );
  INV_X1 U3857 ( .A(n3567), .ZN(n3434) );
  NAND2_X1 U3858 ( .A1(n3243), .A2(n4554), .ZN(n3627) );
  OR2_X1 U3860 ( .A1(n3409), .A2(n3408), .ZN(n3438) );
  INV_X1 U3861 ( .A(n3494), .ZN(n3495) );
  OR2_X1 U3862 ( .A1(n3431), .A2(n3430), .ZN(n3516) );
  OR2_X1 U3863 ( .A1(n3305), .A2(n3304), .ZN(n3484) );
  INV_X1 U3864 ( .A(n4354), .ZN(n3879) );
  INV_X1 U3865 ( .A(n4616), .ZN(n3880) );
  OR2_X1 U3866 ( .A1(n3514), .A2(n3434), .ZN(n3520) );
  OR2_X1 U3867 ( .A1(n3320), .A2(n3319), .ZN(n3453) );
  NAND2_X1 U3868 ( .A1(n3464), .A2(n3523), .ZN(n3451) );
  NAND2_X1 U3869 ( .A1(n4489), .A2(n6910), .ZN(n3307) );
  INV_X1 U3870 ( .A(n5630), .ZN(n4064) );
  INV_X1 U3871 ( .A(n4541), .ZN(n4374) );
  NOR2_X1 U3872 ( .A1(n4307), .A2(n4303), .ZN(n4332) );
  NOR2_X2 U3873 ( .A1(n5935), .A2(n5934), .ZN(n5626) );
  NOR2_X1 U3874 ( .A1(n3915), .A2(n5204), .ZN(n3931) );
  AND2_X1 U3875 ( .A1(n3433), .A2(n3432), .ZN(n3435) );
  INV_X1 U3876 ( .A(n3841), .ZN(n3863) );
  OR2_X1 U3877 ( .A1(n3362), .A2(n6910), .ZN(n3523) );
  OR2_X1 U3878 ( .A1(n5406), .A2(n6312), .ZN(n3534) );
  INV_X1 U3879 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3477) );
  AND2_X1 U3880 ( .A1(n3654), .A2(n3454), .ZN(n3413) );
  XNOR2_X1 U3881 ( .A(n3451), .B(n3450), .ZN(n3452) );
  AND3_X2 U3882 ( .A1(n4558), .A2(n4586), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3583) );
  OR2_X1 U3883 ( .A1(n4238), .A2(n4256), .ZN(n4282) );
  NOR2_X1 U3884 ( .A1(n6786), .A2(n5855), .ZN(n5860) );
  NAND2_X1 U3885 ( .A1(n5626), .A2(n4064), .ZN(n5609) );
  OR2_X1 U3886 ( .A1(n5451), .A2(n5459), .ZN(n4239) );
  NOR2_X1 U3887 ( .A1(n5550), .A2(n4288), .ZN(n5355) );
  NOR2_X1 U3888 ( .A1(n3991), .A2(n6037), .ZN(n3995) );
  INV_X1 U3889 ( .A(n5212), .ZN(n3930) );
  NAND2_X1 U3890 ( .A1(n5558), .A2(n5362), .ZN(n3762) );
  OR2_X1 U3891 ( .A1(n5406), .A2(n3547), .ZN(n3548) );
  NAND2_X1 U3892 ( .A1(n4382), .A2(n3764), .ZN(n3752) );
  CLKBUF_X1 U3893 ( .A(n5265), .Z(n6274) );
  OR2_X1 U3894 ( .A1(n4611), .A2(n3649), .ZN(n3650) );
  XNOR2_X1 U3895 ( .A(n3443), .B(n3482), .ZN(n4533) );
  INV_X1 U3896 ( .A(n4373), .ZN(n4590) );
  NAND2_X1 U3897 ( .A1(n3611), .A2(n3610), .ZN(n3620) );
  NOR2_X1 U3898 ( .A1(n4180), .A2(n5371), .ZN(n4202) );
  NOR2_X1 U3899 ( .A1(n3996), .A2(n6834), .ZN(n4044) );
  INV_X1 U3900 ( .A(n3886), .ZN(n3900) );
  AND2_X1 U3901 ( .A1(n5508), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4258) );
  OR2_X1 U3902 ( .A1(n5513), .A2(n4242), .ZN(n6110) );
  NAND2_X1 U3903 ( .A1(n3745), .A2(n3705), .ZN(n3748) );
  INV_X1 U3904 ( .A(n5452), .ZN(n5449) );
  XNOR2_X1 U3905 ( .A(n4239), .B(n5517), .ZN(n5508) );
  INV_X1 U3906 ( .A(n5411), .ZN(n5412) );
  INV_X1 U3907 ( .A(n5627), .ZN(n5937) );
  AOI21_X1 U3908 ( .B1(n3878), .B2(n3988), .A(n3877), .ZN(n4354) );
  AND2_X1 U3909 ( .A1(n5406), .A2(n5728), .ZN(n3555) );
  NAND2_X1 U3910 ( .A1(n5409), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5408) );
  OR2_X1 U3911 ( .A1(n5965), .A2(n3798), .ZN(n5948) );
  INV_X2 U3912 ( .A(n3556), .ZN(n5693) );
  OR2_X1 U3913 ( .A1(n5406), .A2(n3533), .ZN(n5279) );
  NAND2_X1 U3915 ( .A1(n6330), .A2(n4485), .ZN(n6369) );
  AND2_X2 U3916 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5528) );
  OR3_X1 U3917 ( .A1(n4875), .A2(n5800), .A3(n4721), .ZN(n4899) );
  INV_X1 U3918 ( .A(n4764), .ZN(n4918) );
  OR2_X1 U3919 ( .A1(n4690), .A2(n3838), .ZN(n5064) );
  INV_X1 U3920 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6734) );
  NAND2_X1 U3921 ( .A1(n3620), .A2(n3641), .ZN(n3621) );
  AND2_X1 U3922 ( .A1(n6537), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3644) );
  AND2_X1 U3923 ( .A1(n4202), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4204)
         );
  NAND2_X1 U3924 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n4114), .ZN(n4180)
         );
  NAND2_X1 U3925 ( .A1(n4046), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4079)
         );
  INV_X1 U3926 ( .A(n5890), .ZN(n6079) );
  INV_X1 U3927 ( .A(n6085), .ZN(n6094) );
  AND2_X1 U3928 ( .A1(n6148), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6130) );
  AND2_X1 U3929 ( .A1(n5381), .A2(n3736), .ZN(n5590) );
  INV_X1 U3930 ( .A(n6159), .ZN(n5620) );
  INV_X1 U3931 ( .A(n6150), .ZN(n6155) );
  AND2_X1 U3932 ( .A1(n4209), .A2(n4231), .ZN(n5573) );
  AND2_X1 U3933 ( .A1(n4448), .A2(n4447), .ZN(n6981) );
  INV_X1 U3934 ( .A(n6256), .ZN(n6258) );
  INV_X1 U3935 ( .A(n5666), .ZN(n5907) );
  NAND2_X1 U3936 ( .A1(n4080), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4113)
         );
  NAND2_X1 U3937 ( .A1(n3978), .A2(n3977), .ZN(n5334) );
  INV_X1 U3938 ( .A(n5056), .ZN(n5211) );
  CLKBUF_X1 U3939 ( .A(n4355), .Z(n4711) );
  INV_X1 U3940 ( .A(n3853), .ZN(n3854) );
  INV_X1 U3941 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5480) );
  AND2_X1 U3942 ( .A1(n3762), .A2(n5363), .ZN(n5823) );
  OAI21_X1 U3943 ( .B1(n3556), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5679), 
        .ZN(n5409) );
  CLKBUF_X1 U3944 ( .A(n5221), .Z(n5222) );
  NAND2_X1 U3945 ( .A1(n3794), .A2(n4386), .ZN(n6329) );
  AND2_X1 U3946 ( .A1(n3794), .A2(n6498), .ZN(n5297) );
  NAND2_X1 U3947 ( .A1(n4398), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6626) );
  NOR2_X1 U3948 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5972) );
  INV_X1 U3949 ( .A(n5158), .ZN(n5120) );
  NOR3_X1 U3950 ( .A1(n5800), .A2(n4875), .A3(n4797), .ZN(n4665) );
  INV_X1 U3951 ( .A(n5117), .ZN(n5155) );
  INV_X1 U3952 ( .A(n4899), .ZN(n4754) );
  OAI21_X1 U3953 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n5105), .A(n4918), 
        .ZN(n5012) );
  AND2_X1 U3954 ( .A1(n4875), .A2(n4630), .ZN(n4718) );
  OR2_X1 U3955 ( .A1(n4767), .A2(n4766), .ZN(n4793) );
  INV_X1 U3956 ( .A(n3838), .ZN(n5018) );
  INV_X1 U3957 ( .A(n5064), .ZN(n5096) );
  INV_X1 U3958 ( .A(n5125), .ZN(n6441) );
  INV_X1 U3959 ( .A(n5135), .ZN(n6475) );
  INV_X1 U3960 ( .A(n5111), .ZN(n6427) );
  NOR2_X1 U3961 ( .A1(n4798), .A2(n4874), .ZN(n4948) );
  INV_X1 U3962 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6565) );
  AOI21_X1 U3963 ( .B1(n4262), .B2(n6083), .A(n4261), .ZN(n4263) );
  INV_X1 U3964 ( .A(n4248), .ZN(n4264) );
  OR2_X1 U3965 ( .A1(n5513), .A2(n4255), .ZN(n6138) );
  NAND2_X1 U3966 ( .A1(n6148), .A2(n4240), .ZN(n5890) );
  INV_X1 U3967 ( .A(n6130), .ZN(n6105) );
  NAND2_X1 U3968 ( .A1(n5575), .A2(n5574), .ZN(n5666) );
  INV_X1 U3969 ( .A(n6156), .ZN(n5636) );
  OAI21_X1 U3970 ( .B1(n5573), .B2(n4233), .A(n5551), .ZN(n5655) );
  OAI211_X2 U3971 ( .C1(n4611), .C2(n5540), .A(n6261), .B(n4610), .ZN(n5640)
         );
  INV_X1 U3972 ( .A(n6168), .ZN(n5639) );
  NAND2_X1 U3973 ( .A1(n6645), .A2(n6196), .ZN(n6175) );
  INV_X1 U3974 ( .A(n6981), .ZN(n6196) );
  OR2_X1 U3975 ( .A1(n4611), .A2(n6529), .ZN(n6256) );
  OR2_X1 U3976 ( .A1(n5736), .A2(n3792), .ZN(n5947) );
  INV_X1 U3977 ( .A(n6381), .ZN(n6354) );
  INV_X1 U3978 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U3979 ( .A1(n4665), .A2(n3838), .ZN(n4999) );
  NAND2_X1 U3980 ( .A1(n4718), .A2(n4631), .ZN(n6472) );
  OR2_X1 U3981 ( .A1(n4690), .A2(n5018), .ZN(n4796) );
  INV_X1 U3982 ( .A(n6448), .ZN(n5139) );
  INV_X1 U3983 ( .A(n6426), .ZN(n5110) );
  NOR2_X1 U3984 ( .A1(n4803), .A2(n4802), .ZN(n4841) );
  OR2_X1 U3985 ( .A1(n4842), .A2(n3838), .ZN(n4958) );
  INV_X1 U3986 ( .A(n4948), .ZN(n4952) );
  NAND2_X1 U3987 ( .A1(n4264), .A2(n4263), .ZN(U2801) );
  AND2_X2 U3988 ( .A1(n3116), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3132)
         );
  AND2_X4 U3989 ( .A1(n3132), .A2(n3123), .ZN(n3391) );
  NAND2_X1 U3990 ( .A1(n3391), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3121) );
  AND2_X4 U3991 ( .A1(n3123), .A2(n4513), .ZN(n3352) );
  NAND2_X1 U3992 ( .A1(n3299), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3120)
         );
  AND2_X2 U3993 ( .A1(n4399), .A2(n4513), .ZN(n3370) );
  NAND2_X1 U3994 ( .A1(n3370), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3119)
         );
  NOR2_X4 U3995 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4407) );
  NAND2_X1 U3996 ( .A1(n3346), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3118) );
  AND2_X2 U3997 ( .A1(n3123), .A2(n4490), .ZN(n3292) );
  NAND2_X1 U3998 ( .A1(n3292), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3127) );
  INV_X1 U3999 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3122) );
  NOR2_X2 U4000 ( .A1(n3122), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3133)
         );
  AND2_X2 U4001 ( .A1(n3123), .A2(n3133), .ZN(n3345) );
  NAND2_X1 U4002 ( .A1(n3345), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3126)
         );
  AND2_X2 U4003 ( .A1(n4399), .A2(n4490), .ZN(n3351) );
  NAND2_X1 U4004 ( .A1(n3351), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3125) );
  NAND2_X1 U4005 ( .A1(n3293), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3124) );
  AND2_X2 U4006 ( .A1(n3133), .A2(n5528), .ZN(n3328) );
  NAND2_X1 U4007 ( .A1(n3328), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3131)
         );
  AND2_X2 U4008 ( .A1(n3133), .A2(n4399), .ZN(n3327) );
  NAND2_X1 U4009 ( .A1(n3327), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3130) );
  NAND2_X1 U4010 ( .A1(n3329), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3129) );
  AND2_X2 U4011 ( .A1(n4407), .A2(n4490), .ZN(n3169) );
  NAND2_X1 U4012 ( .A1(n4145), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3128) );
  NAND2_X1 U4013 ( .A1(n4314), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3137) );
  AND2_X2 U4014 ( .A1(n3133), .A2(n4407), .ZN(n4170) );
  NAND2_X1 U4015 ( .A1(n4170), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3136) );
  AND2_X2 U4016 ( .A1(n4407), .A2(n4513), .ZN(n4087) );
  NAND2_X1 U4017 ( .A1(n4087), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3135)
         );
  NAND2_X1 U4018 ( .A1(n3294), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3134)
         );
  AOI22_X1 U4019 ( .A1(n3292), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3144) );
  AOI22_X1 U4020 ( .A1(n3345), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3143) );
  AOI22_X1 U4021 ( .A1(n4170), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3142) );
  AOI22_X1 U4022 ( .A1(n3293), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3141) );
  NAND4_X1 U4023 ( .A1(n3144), .A2(n3143), .A3(n3142), .A4(n3141), .ZN(n3150)
         );
  AOI22_X1 U4024 ( .A1(n3391), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3329), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3148) );
  AOI22_X1 U4025 ( .A1(n3352), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3147) );
  BUF_X4 U4026 ( .A(n3169), .Z(n5436) );
  AOI22_X1 U4027 ( .A1(n3327), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3146) );
  AOI22_X1 U4028 ( .A1(n3328), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3145) );
  NAND4_X1 U4029 ( .A1(n3148), .A2(n3147), .A3(n3146), .A4(n3145), .ZN(n3149)
         );
  NAND2_X1 U4030 ( .A1(n4373), .A2(n4541), .ZN(n3772) );
  AOI22_X1 U4031 ( .A1(n3391), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3154) );
  AOI22_X1 U4032 ( .A1(n3328), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3153) );
  AOI22_X1 U4033 ( .A1(n4170), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3152) );
  AOI22_X1 U4034 ( .A1(n3209), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3151) );
  AOI22_X1 U4035 ( .A1(n3329), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3158) );
  AOI22_X1 U4036 ( .A1(n3327), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3157) );
  AOI22_X1 U4037 ( .A1(n3345), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3156) );
  AOI22_X1 U4038 ( .A1(n3292), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3155) );
  AND2_X2 U4039 ( .A1(n3109), .A2(n3104), .ZN(n3227) );
  AOI22_X1 U4040 ( .A1(n3327), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3162) );
  AOI22_X1 U4041 ( .A1(n3292), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3161) );
  AOI22_X1 U4042 ( .A1(n3391), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3329), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3160) );
  AOI22_X1 U4043 ( .A1(n3209), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3159) );
  NAND4_X1 U4044 ( .A1(n3162), .A2(n3161), .A3(n3160), .A4(n3159), .ZN(n3168)
         );
  AOI22_X1 U4045 ( .A1(n3352), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3166) );
  AOI22_X1 U4046 ( .A1(n3370), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3165) );
  AOI22_X1 U4047 ( .A1(n3351), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3164) );
  AOI22_X1 U4048 ( .A1(n3345), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3163) );
  NAND4_X1 U4049 ( .A1(n3166), .A2(n3165), .A3(n3164), .A4(n3163), .ZN(n3167)
         );
  NAND2_X1 U4050 ( .A1(n3227), .A2(n4381), .ZN(n5377) );
  NOR2_X1 U4051 ( .A1(n3772), .A2(n5377), .ZN(n3198) );
  AOI22_X1 U4052 ( .A1(n3391), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3329), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3173) );
  AOI22_X1 U4053 ( .A1(n3352), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3172) );
  AOI22_X1 U4054 ( .A1(n3327), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3171) );
  AOI22_X1 U4055 ( .A1(n3328), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3170) );
  AOI22_X1 U4056 ( .A1(n3345), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3177) );
  AOI22_X1 U4057 ( .A1(n3102), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3176) );
  AOI22_X1 U4058 ( .A1(n3293), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3175) );
  AOI22_X1 U4059 ( .A1(n3292), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3209), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3174) );
  NAND2_X2 U4060 ( .A1(n3112), .A2(n3114), .ZN(n4598) );
  NAND2_X1 U4061 ( .A1(n3345), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3181)
         );
  NAND2_X1 U4062 ( .A1(n3370), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3180)
         );
  NAND2_X1 U4063 ( .A1(n4314), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3179) );
  NAND2_X1 U4064 ( .A1(n3292), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3178) );
  NAND2_X1 U4065 ( .A1(n3329), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3185) );
  NAND2_X1 U4066 ( .A1(n3391), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3184) );
  NAND2_X1 U4067 ( .A1(n3352), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3183)
         );
  NAND2_X1 U4068 ( .A1(n3346), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3182) );
  NAND2_X1 U4069 ( .A1(n3327), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3189) );
  NAND2_X1 U4070 ( .A1(n3328), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3188)
         );
  NAND2_X1 U4071 ( .A1(n4145), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3187) );
  BUF_X2 U4072 ( .A(n4087), .Z(n4296) );
  NAND2_X1 U4073 ( .A1(n4296), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3186)
         );
  NAND2_X1 U4074 ( .A1(n4170), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3193) );
  NAND2_X1 U4075 ( .A1(n3351), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3192) );
  NAND2_X1 U4076 ( .A1(n3293), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3191) );
  NAND2_X1 U4077 ( .A1(n3294), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3190)
         );
  AND2_X2 U4078 ( .A1(n3198), .A2(n3243), .ZN(n4401) );
  AOI22_X1 U4079 ( .A1(n3345), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3202) );
  AOI22_X1 U4080 ( .A1(n4170), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3201) );
  AOI22_X1 U4081 ( .A1(n3391), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3329), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3200) );
  AOI22_X1 U4082 ( .A1(n3292), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3199) );
  NAND4_X1 U4083 ( .A1(n3202), .A2(n3201), .A3(n3200), .A4(n3199), .ZN(n3208)
         );
  AOI22_X1 U4084 ( .A1(n3327), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3206) );
  AOI22_X1 U4085 ( .A1(n3346), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3205) );
  AOI22_X1 U4086 ( .A1(n3370), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3204) );
  AOI22_X1 U4087 ( .A1(n3209), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3203) );
  NAND4_X1 U4088 ( .A1(n3206), .A2(n3205), .A3(n3204), .A4(n3203), .ZN(n3207)
         );
  OR2_X4 U4089 ( .A1(n3208), .A2(n3207), .ZN(n4586) );
  AOI22_X1 U4090 ( .A1(n3346), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3214) );
  AOI22_X1 U4091 ( .A1(n3370), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3209), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3213) );
  AOI22_X1 U4092 ( .A1(n3351), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3211) );
  AOI22_X1 U4093 ( .A1(n3391), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3210) );
  AND2_X1 U4094 ( .A1(n3211), .A2(n3210), .ZN(n3212) );
  AOI22_X1 U4095 ( .A1(n3345), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3292), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3218) );
  AOI22_X1 U4096 ( .A1(n3327), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3329), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3217) );
  AOI22_X1 U4097 ( .A1(n3328), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3216) );
  AOI22_X1 U4098 ( .A1(n4170), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3215) );
  NAND2_X2 U4099 ( .A1(n3219), .A2(n3110), .ZN(n3654) );
  INV_X1 U4100 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6555) );
  NOR2_X1 U4101 ( .A1(n6555), .A2(n6565), .ZN(n6550) );
  NOR2_X1 U4102 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n3220) );
  OR2_X1 U4103 ( .A1(n6550), .A2(n3220), .ZN(n3633) );
  NAND2_X1 U4104 ( .A1(n3241), .A2(n3633), .ZN(n3248) );
  INV_X1 U4105 ( .A(n3563), .ZN(n3221) );
  NAND2_X1 U4106 ( .A1(n3221), .A2(n3108), .ZN(n4402) );
  NAND2_X1 U4107 ( .A1(n4598), .A2(n4554), .ZN(n4612) );
  NOR2_X2 U4108 ( .A1(n4402), .A2(n4612), .ZN(n3659) );
  AOI21_X1 U4109 ( .B1(n4234), .B2(n3248), .A(n3659), .ZN(n3232) );
  INV_X1 U4110 ( .A(n3261), .ZN(n3222) );
  NOR2_X1 U4111 ( .A1(n3223), .A2(n3242), .ZN(n3231) );
  NAND2_X1 U4112 ( .A1(n3245), .A2(n4373), .ZN(n3224) );
  NAND2_X1 U4113 ( .A1(n3224), .A2(n4381), .ZN(n3226) );
  NAND2_X1 U4115 ( .A1(n3251), .A2(n3261), .ZN(n3225) );
  NAND2_X1 U4116 ( .A1(n3226), .A2(n3225), .ZN(n3229) );
  NAND2_X1 U4117 ( .A1(n3624), .A2(n4541), .ZN(n3264) );
  NAND2_X1 U4118 ( .A1(n3229), .A2(n3264), .ZN(n3240) );
  INV_X1 U4119 ( .A(n3240), .ZN(n3230) );
  AND2_X2 U4120 ( .A1(n3231), .A2(n3230), .ZN(n5546) );
  NAND2_X2 U4121 ( .A1(n5546), .A2(n3241), .ZN(n3655) );
  NAND2_X1 U4122 ( .A1(n3232), .A2(n3655), .ZN(n3233) );
  NAND2_X1 U4123 ( .A1(n3233), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3272) );
  NAND2_X1 U4124 ( .A1(n5972), .A2(n6910), .ZN(n4340) );
  INV_X1 U4125 ( .A(n4340), .ZN(n3283) );
  XNOR2_X1 U4126 ( .A(n6917), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6389)
         );
  NAND2_X1 U4127 ( .A1(n3283), .A2(n6389), .ZN(n3235) );
  INV_X1 U4128 ( .A(n3644), .ZN(n3282) );
  NAND2_X1 U4129 ( .A1(n3282), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3234) );
  NAND2_X1 U4130 ( .A1(n3235), .A2(n3234), .ZN(n3273) );
  NOR2_X1 U4131 ( .A1(n3273), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3236)
         );
  OR2_X2 U4132 ( .A1(n3272), .A2(n3236), .ZN(n3308) );
  NAND2_X1 U4133 ( .A1(n3261), .A2(n4590), .ZN(n3238) );
  NAND2_X1 U4134 ( .A1(n3242), .A2(n4590), .ZN(n3237) );
  NAND3_X1 U4135 ( .A1(n3238), .A2(n3237), .A3(n3241), .ZN(n3239) );
  OAI21_X2 U4136 ( .B1(n3240), .B2(n3239), .A(n3770), .ZN(n3256) );
  AND2_X4 U4137 ( .A1(n3241), .A2(n4586), .ZN(n6648) );
  NAND2_X1 U4138 ( .A1(n6648), .A2(n3627), .ZN(n3244) );
  NAND2_X1 U4139 ( .A1(n3783), .A2(n4541), .ZN(n4404) );
  AND2_X1 U4141 ( .A1(n3245), .A2(n4381), .ZN(n3246) );
  NOR2_X2 U4143 ( .A1(n3769), .A2(n3772), .ZN(n3629) );
  NAND2_X1 U4144 ( .A1(n3248), .A2(n3227), .ZN(n3249) );
  NAND4_X1 U4145 ( .A1(n3256), .A2(n3268), .A3(n3629), .A4(n3249), .ZN(n3250)
         );
  NAND2_X1 U4146 ( .A1(n3250), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3253) );
  NAND2_X1 U4147 ( .A1(n3624), .A2(n3583), .ZN(n3252) );
  NAND2_X1 U4148 ( .A1(n3253), .A2(n3252), .ZN(n3274) );
  NAND2_X1 U4149 ( .A1(n3274), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3255) );
  MUX2_X1 U4150 ( .A(n3644), .B(n4340), .S(n6917), .Z(n3254) );
  NAND2_X1 U4151 ( .A1(n3255), .A2(n3254), .ZN(n3342) );
  INV_X1 U4152 ( .A(n3256), .ZN(n3258) );
  INV_X1 U4153 ( .A(n3783), .ZN(n3257) );
  NAND2_X1 U4154 ( .A1(n3258), .A2(n3257), .ZN(n3778) );
  NAND2_X1 U4155 ( .A1(n3624), .A2(n4558), .ZN(n3259) );
  NAND2_X1 U4156 ( .A1(n3259), .A2(n4541), .ZN(n3260) );
  OAI21_X1 U4157 ( .B1(n3769), .B2(n3260), .A(n4580), .ZN(n3267) );
  AND3_X1 U4158 ( .A1(n4374), .A2(n3770), .A3(n4373), .ZN(n3779) );
  NAND2_X1 U4159 ( .A1(n5972), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6538) );
  INV_X1 U4160 ( .A(n6538), .ZN(n3262) );
  OAI21_X1 U4161 ( .B1(n3770), .B2(n4373), .A(n3262), .ZN(n3263) );
  AOI21_X1 U4162 ( .B1(n3261), .B2(n3779), .A(n3263), .ZN(n3266) );
  NAND2_X1 U4163 ( .A1(n3264), .A2(n6648), .ZN(n3265) );
  NAND3_X1 U4164 ( .A1(n3267), .A2(n3266), .A3(n3265), .ZN(n3270) );
  INV_X1 U4165 ( .A(n3268), .ZN(n3269) );
  NOR2_X1 U4166 ( .A1(n3270), .A2(n3269), .ZN(n3271) );
  NAND2_X1 U4167 ( .A1(n3778), .A2(n3271), .ZN(n3341) );
  NAND2_X2 U4168 ( .A1(n3342), .A2(n3341), .ZN(n3344) );
  NAND2_X1 U4169 ( .A1(n3308), .A2(n3344), .ZN(n3277) );
  INV_X1 U4170 ( .A(n3273), .ZN(n3276) );
  NAND2_X1 U4171 ( .A1(n3278), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3275) );
  INV_X1 U4172 ( .A(n3369), .ZN(n3286) );
  NAND2_X1 U4173 ( .A1(n3278), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3285) );
  AND2_X1 U4174 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3279) );
  NAND2_X1 U4175 ( .A1(n3279), .A2(n6505), .ZN(n4866) );
  INV_X1 U4176 ( .A(n3279), .ZN(n3280) );
  NAND2_X1 U4177 ( .A1(n3280), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3281) );
  NAND2_X1 U4178 ( .A1(n4866), .A2(n3281), .ZN(n4726) );
  AOI22_X1 U4179 ( .A1(n3283), .A2(n4726), .B1(n3282), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3284) );
  NAND2_X1 U4180 ( .A1(n3278), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3291) );
  NAND3_X1 U4181 ( .A1(n6734), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6388) );
  INV_X1 U4182 ( .A(n6388), .ZN(n3287) );
  NAND2_X1 U4183 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3287), .ZN(n4632) );
  NAND2_X1 U4184 ( .A1(n6734), .A2(n4632), .ZN(n3288) );
  NAND3_X1 U4185 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4917) );
  INV_X1 U4186 ( .A(n4917), .ZN(n4544) );
  NAND2_X1 U4187 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4544), .ZN(n4654) );
  NAND2_X1 U4188 ( .A1(n3288), .A2(n4654), .ZN(n4759) );
  OAI22_X1 U4189 ( .A1(n4340), .A2(n4759), .B1(n3644), .B2(n6734), .ZN(n3289)
         );
  INV_X1 U4190 ( .A(n3289), .ZN(n3290) );
  AOI22_X1 U4191 ( .A1(n5438), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4192 ( .A1(n5428), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3297) );
  INV_X1 U4193 ( .A(n3330), .ZN(n5434) );
  AOI22_X1 U4194 ( .A1(n5434), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5433), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4195 ( .A1(n5427), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3295) );
  NAND4_X1 U4196 ( .A1(n3298), .A2(n3297), .A3(n3296), .A4(n3295), .ZN(n3305)
         );
  AOI22_X1 U4198 ( .A1(n4122), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3303) );
  AOI22_X1 U4199 ( .A1(n4295), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5435), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4201 ( .A1(n4315), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4202 ( .A1(n4320), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3300) );
  NAND4_X1 U4203 ( .A1(n3303), .A2(n3302), .A3(n3301), .A4(n3300), .ZN(n3304)
         );
  AOI22_X1 U4204 ( .A1(n3616), .A2(n3484), .B1(n3583), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3306) );
  NAND2_X1 U4205 ( .A1(n3309), .A2(n3308), .ZN(n3310) );
  INV_X1 U4206 ( .A(n3337), .ZN(n4376) );
  AOI22_X1 U4207 ( .A1(n4320), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4208 ( .A1(n5438), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4209 ( .A1(n3101), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5435), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3312) );
  AOI22_X1 U4210 ( .A1(n5428), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3311) );
  NAND4_X1 U4211 ( .A1(n3314), .A2(n3313), .A3(n3312), .A4(n3311), .ZN(n3320)
         );
  AOI22_X1 U4212 ( .A1(n3391), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3299), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U4213 ( .A1(n5434), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5433), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3317) );
  AOI22_X1 U4214 ( .A1(n4315), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4215 ( .A1(n4218), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3315) );
  NAND4_X1 U4216 ( .A1(n3318), .A2(n3317), .A3(n3316), .A4(n3315), .ZN(n3319)
         );
  NAND2_X1 U4217 ( .A1(n4376), .A2(n3453), .ZN(n3321) );
  OAI21_X2 U4218 ( .B1(n4400), .B2(STATE2_REG_0__SCAN_IN), .A(n3321), .ZN(
        n3449) );
  INV_X1 U4219 ( .A(n3453), .ZN(n3340) );
  AOI22_X1 U4220 ( .A1(n3299), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4221 ( .A1(n5438), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3325) );
  AOI22_X1 U4222 ( .A1(n5428), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3324) );
  AOI22_X1 U4223 ( .A1(n5433), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3323) );
  NAND4_X1 U4224 ( .A1(n3326), .A2(n3325), .A3(n3324), .A4(n3323), .ZN(n3336)
         );
  AOI22_X1 U4225 ( .A1(n4315), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4320), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4226 ( .A1(n3391), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3333) );
  AOI22_X1 U4227 ( .A1(n5435), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3332) );
  AOI22_X1 U4228 ( .A1(n3100), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3331) );
  NAND4_X1 U4229 ( .A1(n3334), .A2(n3333), .A3(n3332), .A4(n3331), .ZN(n3335)
         );
  NOR2_X1 U4230 ( .A1(n3337), .A2(n3527), .ZN(n3359) );
  INV_X1 U4231 ( .A(n3359), .ZN(n3339) );
  NAND2_X1 U4232 ( .A1(n3583), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3338) );
  OAI211_X1 U4233 ( .C1(n3340), .C2(n3383), .A(n3339), .B(n3338), .ZN(n3450)
         );
  OR2_X2 U4234 ( .A1(n3342), .A2(n3341), .ZN(n3343) );
  AOI22_X1 U4235 ( .A1(n3391), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3350) );
  AOI22_X1 U4236 ( .A1(n5438), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3349) );
  AOI22_X1 U4237 ( .A1(n4315), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5435), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3348) );
  AOI22_X1 U4238 ( .A1(n4320), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3347) );
  NAND4_X1 U4239 ( .A1(n3350), .A2(n3349), .A3(n3348), .A4(n3347), .ZN(n3358)
         );
  AOI22_X1 U4240 ( .A1(n5428), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3356) );
  AOI22_X1 U4241 ( .A1(n3100), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5433), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3355) );
  AOI22_X1 U4242 ( .A1(n3299), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3354) );
  AOI22_X1 U4243 ( .A1(n5427), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3353) );
  NAND4_X1 U4244 ( .A1(n3356), .A2(n3355), .A3(n3354), .A4(n3353), .ZN(n3357)
         );
  NAND2_X1 U4245 ( .A1(n3658), .A2(n3527), .ZN(n3362) );
  NAND2_X1 U4246 ( .A1(n3359), .A2(n3466), .ZN(n3461) );
  OAI21_X1 U4247 ( .B1(n3466), .B2(n3523), .A(n3461), .ZN(n3360) );
  INV_X1 U4248 ( .A(n3360), .ZN(n3361) );
  OAI21_X1 U4249 ( .B1(n3840), .B2(STATE2_REG_0__SCAN_IN), .A(n3361), .ZN(
        n3365) );
  NAND2_X1 U4250 ( .A1(n3583), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3364) );
  AOI21_X1 U4251 ( .B1(n3770), .B2(n3466), .A(n6910), .ZN(n3363) );
  NAND3_X1 U4252 ( .A1(n3364), .A2(n3363), .A3(n3362), .ZN(n3460) );
  NAND2_X1 U4253 ( .A1(n3365), .A2(n3460), .ZN(n3464) );
  OAI21_X1 U4254 ( .B1(n3449), .B2(n3450), .A(n3451), .ZN(n3367) );
  NAND2_X1 U4255 ( .A1(n3449), .A2(n3450), .ZN(n3366) );
  NAND2_X1 U4256 ( .A1(n3367), .A2(n3366), .ZN(n3481) );
  XNOR2_X2 U4257 ( .A(n3369), .B(n3368), .ZN(n4501) );
  NAND2_X1 U4258 ( .A1(n4501), .A2(n6910), .ZN(n3382) );
  AOI22_X1 U4259 ( .A1(n5438), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4260 ( .A1(n5428), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4261 ( .A1(n5434), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5433), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3372) );
  AOI22_X1 U4262 ( .A1(n5427), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3371) );
  NAND4_X1 U4263 ( .A1(n3374), .A2(n3373), .A3(n3372), .A4(n3371), .ZN(n3380)
         );
  AOI22_X1 U4264 ( .A1(n3391), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4265 ( .A1(n3352), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5435), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3377) );
  AOI22_X1 U4266 ( .A1(n4315), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U4267 ( .A1(n4320), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3375) );
  NAND4_X1 U4268 ( .A1(n3378), .A2(n3377), .A3(n3376), .A4(n3375), .ZN(n3379)
         );
  NAND2_X1 U4269 ( .A1(n4376), .A2(n3414), .ZN(n3381) );
  INV_X1 U4270 ( .A(n3383), .ZN(n3384) );
  AOI22_X1 U4271 ( .A1(n3583), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3384), 
        .B2(n3414), .ZN(n3385) );
  XNOR2_X2 U4272 ( .A(n3386), .B(n3385), .ZN(n3482) );
  AND3_X2 U4273 ( .A1(n4538), .A2(n3481), .A3(n3482), .ZN(n3496) );
  AOI22_X1 U4274 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n5438), .B1(n3322), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3390) );
  AOI22_X1 U4275 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4117), .B1(n5428), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3389) );
  AOI22_X1 U4276 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5434), .B1(n5433), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3388) );
  AOI22_X1 U4277 ( .A1(n5427), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3387) );
  NAND4_X1 U4278 ( .A1(n3390), .A2(n3389), .A3(n3388), .A4(n3387), .ZN(n3397)
         );
  AOI22_X1 U4279 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n4122), .B1(n3101), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3395) );
  AOI22_X1 U4280 ( .A1(n4295), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n5435), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4281 ( .A1(n4315), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3393) );
  AOI22_X1 U4282 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4320), .B1(n4218), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3392) );
  NAND4_X1 U4283 ( .A1(n3395), .A2(n3394), .A3(n3393), .A4(n3392), .ZN(n3396)
         );
  NAND2_X1 U4284 ( .A1(n3616), .A2(n3497), .ZN(n3399) );
  NAND2_X1 U4285 ( .A1(n3583), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3398) );
  NAND2_X1 U4286 ( .A1(n3399), .A2(n3398), .ZN(n3494) );
  NAND2_X1 U4287 ( .A1(n3496), .A2(n3494), .ZN(n3412) );
  AOI22_X1 U4288 ( .A1(n5438), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3403) );
  INV_X1 U4289 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n6791) );
  AOI22_X1 U4290 ( .A1(n5428), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3402) );
  AOI22_X1 U4291 ( .A1(n5434), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5433), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3401) );
  AOI22_X1 U4292 ( .A1(n5427), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3400) );
  NAND4_X1 U4293 ( .A1(n3403), .A2(n3402), .A3(n3401), .A4(n3400), .ZN(n3409)
         );
  AOI22_X1 U4294 ( .A1(n4122), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3407) );
  AOI22_X1 U4295 ( .A1(n4295), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5435), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3406) );
  AOI22_X1 U4296 ( .A1(n4315), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3405) );
  AOI22_X1 U4297 ( .A1(n4320), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3404) );
  NAND4_X1 U4298 ( .A1(n3407), .A2(n3406), .A3(n3405), .A4(n3404), .ZN(n3408)
         );
  NAND2_X1 U4299 ( .A1(n3616), .A2(n3438), .ZN(n3411) );
  NAND2_X1 U4300 ( .A1(n3583), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3410) );
  NAND2_X1 U4301 ( .A1(n3411), .A2(n3410), .ZN(n3420) );
  NAND2_X1 U4302 ( .A1(n3874), .A2(n3567), .ZN(n3419) );
  NAND2_X1 U4303 ( .A1(n3466), .A2(n3453), .ZN(n3445) );
  INV_X1 U4304 ( .A(n3414), .ZN(n3444) );
  NAND2_X1 U4305 ( .A1(n3445), .A2(n3444), .ZN(n3486) );
  NAND2_X1 U4306 ( .A1(n3486), .A2(n3484), .ZN(n3498) );
  INV_X1 U4307 ( .A(n3497), .ZN(n3415) );
  OR2_X1 U4308 ( .A1(n3498), .A2(n3415), .ZN(n3416) );
  XNOR2_X1 U4309 ( .A(n3416), .B(n3438), .ZN(n3417) );
  NAND2_X1 U4310 ( .A1(n3417), .A2(n6648), .ZN(n3418) );
  NAND2_X1 U4311 ( .A1(n3419), .A2(n3418), .ZN(n3505) );
  INV_X1 U4312 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5187) );
  XNOR2_X1 U4313 ( .A(n3505), .B(n5187), .ZN(n6273) );
  NAND2_X1 U4314 ( .A1(n3496), .A2(n3421), .ZN(n3436) );
  AOI22_X1 U4315 ( .A1(n5438), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3425) );
  AOI22_X1 U4316 ( .A1(n5428), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3424) );
  AOI22_X1 U4317 ( .A1(n5434), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5433), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3423) );
  AOI22_X1 U4318 ( .A1(n5427), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3422) );
  NAND4_X1 U4319 ( .A1(n3425), .A2(n3424), .A3(n3423), .A4(n3422), .ZN(n3431)
         );
  AOI22_X1 U4320 ( .A1(n4122), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4321 ( .A1(n4295), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n5435), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3428) );
  AOI22_X1 U4322 ( .A1(n4315), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3427) );
  AOI22_X1 U4323 ( .A1(n4320), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3426) );
  NAND4_X1 U4324 ( .A1(n3429), .A2(n3428), .A3(n3427), .A4(n3426), .ZN(n3430)
         );
  NAND2_X1 U4325 ( .A1(n3616), .A2(n3516), .ZN(n3433) );
  NAND2_X1 U4326 ( .A1(n3583), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3432) );
  NOR2_X2 U4327 ( .A1(n3436), .A2(n3435), .ZN(n3510) );
  NOR2_X1 U4328 ( .A1(n3510), .A2(n3434), .ZN(n3437) );
  NAND2_X1 U4329 ( .A1(n3436), .A2(n3435), .ZN(n3878) );
  NAND2_X1 U4330 ( .A1(n3437), .A2(n3878), .ZN(n3442) );
  NAND2_X1 U4331 ( .A1(n3497), .A2(n3438), .ZN(n3439) );
  OR2_X1 U4332 ( .A1(n3498), .A2(n3439), .ZN(n3515) );
  XNOR2_X1 U4333 ( .A(n3515), .B(n3516), .ZN(n3440) );
  NAND2_X1 U4334 ( .A1(n3440), .A2(n6648), .ZN(n3441) );
  INV_X1 U4335 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6752) );
  XNOR2_X1 U4336 ( .A(n3507), .B(n6752), .ZN(n5270) );
  AND2_X1 U4337 ( .A1(n6273), .A2(n5270), .ZN(n3504) );
  INV_X1 U4338 ( .A(n3481), .ZN(n3443) );
  NAND2_X1 U4339 ( .A1(n4533), .A2(n3567), .ZN(n3448) );
  XNOR2_X1 U4340 ( .A(n3445), .B(n3444), .ZN(n3446) );
  AND2_X1 U4341 ( .A1(n3770), .A2(n4541), .ZN(n3782) );
  AOI21_X1 U4342 ( .B1(n3446), .B2(n6648), .A(n3782), .ZN(n3447) );
  NAND2_X1 U4343 ( .A1(n6291), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3476)
         );
  NAND2_X1 U4344 ( .A1(n4526), .A2(n3567), .ZN(n3459) );
  XNOR2_X1 U4345 ( .A(n3466), .B(n3453), .ZN(n3456) );
  INV_X1 U4346 ( .A(n6648), .ZN(n3467) );
  INV_X1 U4347 ( .A(n3772), .ZN(n3455) );
  OAI211_X1 U4348 ( .C1(n3456), .C2(n3467), .A(n3455), .B(n4594), .ZN(n3457)
         );
  INV_X1 U4349 ( .A(n3457), .ZN(n3458) );
  NAND2_X1 U4350 ( .A1(n3459), .A2(n3458), .ZN(n4479) );
  INV_X1 U4351 ( .A(n3460), .ZN(n3462) );
  NAND2_X1 U4352 ( .A1(n3462), .A2(n3461), .ZN(n3463) );
  NAND2_X2 U4353 ( .A1(n3464), .A2(n3463), .ZN(n3838) );
  OR2_X1 U4354 ( .A1(n3838), .A2(n3434), .ZN(n3470) );
  INV_X1 U4355 ( .A(n3782), .ZN(n3465) );
  OAI21_X1 U4356 ( .B1(n3467), .B2(n3466), .A(n3465), .ZN(n3468) );
  INV_X1 U4357 ( .A(n3468), .ZN(n3469) );
  NAND2_X1 U4358 ( .A1(n3470), .A2(n3469), .ZN(n4425) );
  NAND2_X1 U4359 ( .A1(n4425), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3471)
         );
  INV_X1 U4360 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4486) );
  NAND2_X1 U4361 ( .A1(n3471), .A2(n4486), .ZN(n3473) );
  AND2_X1 U4362 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3472) );
  NAND2_X1 U4363 ( .A1(n4425), .A2(n3472), .ZN(n3474) );
  AND2_X1 U4364 ( .A1(n3473), .A2(n3474), .ZN(n4478) );
  INV_X1 U4365 ( .A(n3474), .ZN(n3475) );
  NAND2_X1 U4366 ( .A1(n3476), .A2(n6289), .ZN(n3480) );
  INV_X1 U4367 ( .A(n6291), .ZN(n3478) );
  NAND2_X1 U4368 ( .A1(n3478), .A2(n3477), .ZN(n3479) );
  NAND2_X1 U4369 ( .A1(n3480), .A2(n3479), .ZN(n6282) );
  INV_X1 U4370 ( .A(n6282), .ZN(n3491) );
  NAND2_X1 U4371 ( .A1(n3482), .A2(n3481), .ZN(n3483) );
  NAND2_X1 U4372 ( .A1(n3852), .A2(n3567), .ZN(n3489) );
  INV_X1 U4373 ( .A(n3484), .ZN(n3485) );
  XNOR2_X1 U4374 ( .A(n3486), .B(n3485), .ZN(n3487) );
  NAND2_X1 U4375 ( .A1(n3487), .A2(n6648), .ZN(n3488) );
  INV_X1 U4376 ( .A(n6283), .ZN(n3490) );
  NAND2_X1 U4377 ( .A1(n3491), .A2(n3490), .ZN(n6280) );
  NAND2_X1 U4378 ( .A1(n3492), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3493)
         );
  NAND2_X1 U4379 ( .A1(n6280), .A2(n3493), .ZN(n5167) );
  NAND2_X1 U4380 ( .A1(n3860), .A2(n3567), .ZN(n3501) );
  XNOR2_X1 U4381 ( .A(n3498), .B(n3497), .ZN(n3499) );
  NAND2_X1 U4382 ( .A1(n3499), .A2(n6648), .ZN(n3500) );
  NAND2_X1 U4383 ( .A1(n3501), .A2(n3500), .ZN(n3502) );
  INV_X1 U4384 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6361) );
  XNOR2_X1 U4385 ( .A(n3502), .B(n6361), .ZN(n5166) );
  NAND2_X1 U4386 ( .A1(n3502), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3503)
         );
  NAND2_X1 U4387 ( .A1(n5169), .A2(n3503), .ZN(n5265) );
  NAND2_X1 U4388 ( .A1(n3504), .A2(n5265), .ZN(n5268) );
  XNOR2_X1 U4389 ( .A(n3507), .B(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3506)
         );
  NAND2_X1 U4390 ( .A1(n3505), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5266)
         );
  OR2_X1 U4391 ( .A1(n3506), .A2(n5266), .ZN(n5267) );
  NAND2_X1 U4392 ( .A1(n3507), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3508)
         );
  AND2_X1 U4393 ( .A1(n5267), .A2(n3508), .ZN(n3509) );
  NAND2_X1 U4394 ( .A1(n5268), .A2(n3509), .ZN(n6263) );
  INV_X1 U4395 ( .A(n3510), .ZN(n3525) );
  NAND2_X1 U4396 ( .A1(n3616), .A2(n3527), .ZN(n3512) );
  NAND2_X1 U4397 ( .A1(n3583), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3511) );
  NAND2_X1 U4398 ( .A1(n3512), .A2(n3511), .ZN(n3513) );
  XNOR2_X2 U4399 ( .A(n3525), .B(n3513), .ZN(n3881) );
  INV_X1 U4400 ( .A(n3881), .ZN(n3514) );
  INV_X1 U4401 ( .A(n3515), .ZN(n3517) );
  NAND2_X1 U4402 ( .A1(n3517), .A2(n3516), .ZN(n3526) );
  XNOR2_X1 U4403 ( .A(n3526), .B(n3527), .ZN(n3518) );
  NAND2_X1 U4404 ( .A1(n3518), .A2(n6648), .ZN(n3519) );
  INV_X1 U4405 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n5189) );
  XNOR2_X1 U4406 ( .A(n3521), .B(n5189), .ZN(n6262) );
  NAND2_X1 U4407 ( .A1(n6263), .A2(n6262), .ZN(n6265) );
  NAND2_X1 U4408 ( .A1(n3521), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3522)
         );
  NAND2_X1 U4409 ( .A1(n6265), .A2(n3522), .ZN(n5181) );
  NOR2_X1 U4410 ( .A1(n3523), .A2(n3434), .ZN(n3524) );
  INV_X1 U4411 ( .A(n3526), .ZN(n3528) );
  NAND3_X1 U4412 ( .A1(n3528), .A2(n6648), .A3(n3527), .ZN(n3529) );
  NAND2_X1 U4413 ( .A1(n5693), .A2(n3529), .ZN(n3530) );
  INV_X1 U4414 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6799) );
  XNOR2_X1 U4415 ( .A(n3530), .B(n6799), .ZN(n5183) );
  NAND2_X1 U4416 ( .A1(n5181), .A2(n5183), .ZN(n5182) );
  NAND2_X1 U4417 ( .A1(n3530), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3531)
         );
  NAND2_X1 U4418 ( .A1(n5182), .A2(n3531), .ZN(n5200) );
  INV_X1 U4419 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6801) );
  NAND2_X1 U4420 ( .A1(n5406), .A2(n6801), .ZN(n5201) );
  NAND2_X1 U4421 ( .A1(n5200), .A2(n5201), .ZN(n3532) );
  OR2_X1 U4422 ( .A1(n5406), .A2(n6801), .ZN(n5202) );
  NAND2_X1 U4423 ( .A1(n3532), .A2(n5202), .ZN(n5221) );
  INV_X1 U4424 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3533) );
  NAND2_X1 U4425 ( .A1(n5406), .A2(n3533), .ZN(n5220) );
  NAND2_X1 U4426 ( .A1(n5221), .A2(n5220), .ZN(n5280) );
  INV_X1 U4427 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6312) );
  AND2_X1 U4428 ( .A1(n5406), .A2(n6312), .ZN(n3536) );
  INV_X1 U4429 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3538) );
  NOR2_X1 U4430 ( .A1(n5693), .A2(n3538), .ZN(n5321) );
  XNOR2_X1 U4431 ( .A(n5693), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5325)
         );
  INV_X1 U4432 ( .A(n5325), .ZN(n3537) );
  OR2_X1 U4433 ( .A1(n5321), .A2(n3537), .ZN(n3542) );
  NAND2_X1 U4434 ( .A1(n5406), .A2(n3538), .ZN(n5323) );
  INV_X1 U4435 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3539) );
  NAND2_X1 U4436 ( .A1(n5406), .A2(n3539), .ZN(n3540) );
  INV_X1 U4437 ( .A(n5290), .ZN(n3543) );
  INV_X1 U4438 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5388) );
  NAND2_X1 U4439 ( .A1(n3543), .A2(n3105), .ZN(n3544) );
  NAND2_X1 U4440 ( .A1(n3544), .A2(n5288), .ZN(n5382) );
  INV_X1 U4441 ( .A(n5382), .ZN(n3545) );
  INV_X1 U4442 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5790) );
  INV_X1 U4443 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5791) );
  NAND2_X1 U4444 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5763) );
  OAI21_X1 U4445 ( .B1(n5791), .B2(n5763), .A(n5693), .ZN(n3546) );
  INV_X1 U4446 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5762) );
  INV_X1 U4447 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5959) );
  AND3_X1 U4448 ( .A1(n5791), .A2(n5762), .A3(n5959), .ZN(n3547) );
  AND2_X1 U4449 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3803) );
  AND2_X1 U4450 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5764) );
  AND2_X1 U4451 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3800) );
  NAND3_X1 U4452 ( .A1(n3803), .A2(n5764), .A3(n3800), .ZN(n3549) );
  NAND2_X1 U4453 ( .A1(n5693), .A2(n3549), .ZN(n3554) );
  INV_X1 U4454 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5417) );
  INV_X1 U4455 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6785) );
  INV_X1 U4456 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5744) );
  INV_X1 U4457 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3550) );
  NAND4_X1 U4458 ( .A1(n5417), .A2(n6785), .A3(n5744), .A4(n3550), .ZN(n3551)
         );
  INV_X1 U4459 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3722) );
  INV_X1 U4460 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U4461 ( .A1(n3722), .A2(n5780), .ZN(n5765) );
  NOR2_X1 U4462 ( .A1(n3551), .A2(n5765), .ZN(n3552) );
  NOR2_X1 U4463 ( .A1(n5693), .A2(n3552), .ZN(n3553) );
  AOI21_X1 U4464 ( .B1(n5774), .B2(n3554), .A(n3553), .ZN(n5663) );
  XNOR2_X1 U4465 ( .A(n5693), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5662)
         );
  AND2_X2 U4466 ( .A1(n5663), .A2(n5662), .ZN(n5664) );
  INV_X1 U4467 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5728) );
  NOR2_X2 U4468 ( .A1(n5664), .A2(n3555), .ZN(n5653) );
  INV_X1 U4469 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5729) );
  NOR2_X1 U4470 ( .A1(n3556), .A2(n5729), .ZN(n5652) );
  NAND2_X1 U4472 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5712) );
  NOR2_X4 U4473 ( .A1(n5643), .A2(n5712), .ZN(n5479) );
  NOR2_X1 U4474 ( .A1(n5693), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5651)
         );
  NOR2_X1 U4475 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U4476 ( .A1(n5651), .A2(n5711), .ZN(n5477) );
  NOR2_X1 U4477 ( .A1(n3814), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3811)
         );
  INV_X1 U4478 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3557) );
  NAND2_X1 U4479 ( .A1(n3616), .A2(n4580), .ZN(n3559) );
  NAND2_X1 U4480 ( .A1(n3559), .A2(n4594), .ZN(n3571) );
  XNOR2_X1 U4481 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3578) );
  NAND2_X1 U4482 ( .A1(n6917), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3577) );
  XNOR2_X1 U4483 ( .A(n3578), .B(n3577), .ZN(n3638) );
  NAND2_X1 U4484 ( .A1(n3560), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3561) );
  AND2_X1 U4485 ( .A1(n3577), .A2(n3561), .ZN(n3562) );
  AND2_X1 U4486 ( .A1(n3616), .A2(n3562), .ZN(n3566) );
  NAND2_X1 U4487 ( .A1(n3658), .A2(n4594), .ZN(n3652) );
  AOI21_X1 U4488 ( .B1(n3652), .B2(n3562), .A(n3770), .ZN(n3565) );
  NAND2_X1 U4489 ( .A1(n3241), .A2(n4594), .ZN(n3564) );
  NAND2_X1 U4490 ( .A1(n3563), .A2(n3564), .ZN(n3586) );
  OAI211_X1 U4491 ( .C1(n3571), .C2(n3638), .A(n3566), .B(n3570), .ZN(n3569)
         );
  NAND3_X1 U4492 ( .A1(n3571), .A2(STATE2_REG_0__SCAN_IN), .A3(n3638), .ZN(
        n3568) );
  NAND3_X1 U4493 ( .A1(n3569), .A2(n3617), .A3(n3568), .ZN(n3575) );
  INV_X1 U4494 ( .A(n3570), .ZN(n3573) );
  INV_X1 U4495 ( .A(n3571), .ZN(n3572) );
  NAND3_X1 U4496 ( .A1(n3573), .A2(n3572), .A3(n3638), .ZN(n3574) );
  NAND2_X1 U4497 ( .A1(n3575), .A2(n3574), .ZN(n3584) );
  INV_X1 U4498 ( .A(n3586), .ZN(n3576) );
  NAND2_X1 U4499 ( .A1(n3584), .A2(n3576), .ZN(n3582) );
  INV_X1 U4500 ( .A(n3577), .ZN(n3579) );
  NAND2_X1 U4501 ( .A1(n3579), .A2(n3578), .ZN(n3581) );
  NAND2_X1 U4502 ( .A1(n4719), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3580) );
  NAND2_X1 U4503 ( .A1(n3581), .A2(n3580), .ZN(n3592) );
  XNOR2_X1 U4504 ( .A(n5537), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3590)
         );
  XNOR2_X1 U4505 ( .A(n3592), .B(n3590), .ZN(n3637) );
  NAND3_X1 U4506 ( .A1(n3582), .A2(n3637), .A3(n3616), .ZN(n3589) );
  NOR2_X1 U4507 ( .A1(n3605), .A2(n3637), .ZN(n3587) );
  INV_X1 U4508 ( .A(n3584), .ZN(n3585) );
  OAI21_X1 U4509 ( .B1(n3587), .B2(n3586), .A(n3585), .ZN(n3588) );
  NAND2_X1 U4510 ( .A1(n3589), .A2(n3588), .ZN(n3596) );
  INV_X1 U4511 ( .A(n3590), .ZN(n3591) );
  NAND2_X1 U4512 ( .A1(n3592), .A2(n3591), .ZN(n3594) );
  NAND2_X1 U4513 ( .A1(n6505), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3593) );
  NAND2_X1 U4514 ( .A1(n3594), .A2(n3593), .ZN(n3602) );
  XNOR2_X1 U4515 ( .A(n3122), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3600)
         );
  XNOR2_X1 U4516 ( .A(n3602), .B(n3600), .ZN(n3639) );
  INV_X1 U4517 ( .A(n3639), .ZN(n3597) );
  NAND2_X1 U4518 ( .A1(n3605), .A2(n3597), .ZN(n3595) );
  NAND2_X1 U4519 ( .A1(n3596), .A2(n3595), .ZN(n3599) );
  NAND2_X1 U4520 ( .A1(n3609), .A2(n3597), .ZN(n3598) );
  NAND2_X1 U4521 ( .A1(n3599), .A2(n3598), .ZN(n3607) );
  INV_X1 U4522 ( .A(n3600), .ZN(n3601) );
  NAND2_X1 U4523 ( .A1(n3602), .A2(n3601), .ZN(n3604) );
  NAND2_X1 U4524 ( .A1(n6734), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3603) );
  NAND2_X1 U4525 ( .A1(n3604), .A2(n3603), .ZN(n3613) );
  INV_X1 U4526 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6387) );
  NAND2_X1 U4527 ( .A1(n3605), .A2(n3608), .ZN(n3606) );
  NAND2_X1 U4528 ( .A1(n3607), .A2(n3606), .ZN(n3611) );
  AOI22_X1 U4529 ( .A1(n3609), .A2(n3608), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6910), .ZN(n3610) );
  AND2_X1 U4530 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6387), .ZN(n3612)
         );
  OR2_X1 U4531 ( .A1(n3613), .A2(n3612), .ZN(n3615) );
  INV_X1 U4532 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U4533 ( .A1(n5974), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3614) );
  NOR2_X1 U4534 ( .A1(n3227), .A2(n3658), .ZN(n3623) );
  NAND2_X1 U4535 ( .A1(n3261), .A2(n3623), .ZN(n3780) );
  NOR2_X1 U4536 ( .A1(n4413), .A2(n3241), .ZN(n3786) );
  NAND2_X1 U4537 ( .A1(n6532), .A2(n3786), .ZN(n3643) );
  INV_X1 U4538 ( .A(n3624), .ZN(n3626) );
  AND2_X1 U4539 ( .A1(n3624), .A2(n4586), .ZN(n3625) );
  OAI22_X1 U4540 ( .A1(n3627), .A2(n3626), .B1(n6648), .B2(n3625), .ZN(n3776)
         );
  INV_X1 U4541 ( .A(n3776), .ZN(n3630) );
  NAND2_X1 U4542 ( .A1(n3780), .A2(n3770), .ZN(n3628) );
  NAND2_X1 U4543 ( .A1(n3629), .A2(n3628), .ZN(n3653) );
  OR2_X1 U4544 ( .A1(n3630), .A2(n3653), .ZN(n3632) );
  INV_X1 U4545 ( .A(n5546), .ZN(n3631) );
  NAND2_X1 U4546 ( .A1(n3632), .A2(n3631), .ZN(n4393) );
  INV_X1 U4547 ( .A(n3633), .ZN(n3635) );
  INV_X1 U4548 ( .A(STATE_REG_0__SCAN_IN), .ZN(n3634) );
  NAND2_X1 U4549 ( .A1(n3635), .A2(n3634), .ZN(n6554) );
  INV_X1 U4550 ( .A(n6554), .ZN(n4447) );
  NAND4_X1 U4551 ( .A1(n3639), .A2(n3638), .A3(n3637), .A4(n3636), .ZN(n3640)
         );
  NAND2_X1 U4552 ( .A1(n3641), .A2(n3640), .ZN(n5541) );
  NOR2_X1 U4553 ( .A1(READY_N), .A2(n5541), .ZN(n4606) );
  OAI211_X1 U4554 ( .C1(n3241), .C2(n4447), .A(n4590), .B(n4606), .ZN(n3642)
         );
  NAND3_X1 U4555 ( .A1(n3643), .A2(n4393), .A3(n3642), .ZN(n3645) );
  NAND2_X1 U4556 ( .A1(n3645), .A2(n6525), .ZN(n3651) );
  NAND2_X1 U4557 ( .A1(n3241), .A2(n6554), .ZN(n4241) );
  INV_X1 U4558 ( .A(READY_N), .ZN(n3646) );
  NAND3_X1 U4559 ( .A1(n4401), .A2(n4241), .A3(n3646), .ZN(n3647) );
  NAND3_X1 U4560 ( .A1(n3647), .A2(n4586), .A3(n4612), .ZN(n3648) );
  NAND2_X1 U4561 ( .A1(n3648), .A2(n4373), .ZN(n3649) );
  OR2_X1 U4562 ( .A1(n3653), .A2(n3563), .ZN(n5540) );
  NAND2_X1 U4563 ( .A1(n4586), .A2(n3654), .ZN(n3665) );
  INV_X2 U4564 ( .A(n3665), .ZN(n4382) );
  AOI22_X1 U4565 ( .A1(n3659), .A2(n4558), .B1(n4401), .B2(n4382), .ZN(n3656)
         );
  NAND4_X1 U4566 ( .A1(n6516), .A2(n5540), .A3(n3656), .A4(n3655), .ZN(n3657)
         );
  NAND2_X1 U4567 ( .A1(n4401), .A2(n6648), .ZN(n6529) );
  NAND2_X1 U4568 ( .A1(n3659), .A2(n3658), .ZN(n3660) );
  NAND2_X1 U4569 ( .A1(n6529), .A2(n3660), .ZN(n3661) );
  NAND2_X4 U4570 ( .A1(n4541), .A2(n4580), .ZN(n3764) );
  INV_X2 U4571 ( .A(n3764), .ZN(n3664) );
  NOR2_X1 U4572 ( .A1(n3752), .A2(EBX_REG_5__SCAN_IN), .ZN(n3662) );
  AOI21_X1 U4573 ( .B1(EBX_REG_5__SCAN_IN), .B2(n5616), .A(n3662), .ZN(n3663)
         );
  OAI21_X1 U4574 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n5486), .A(n3663), 
        .ZN(n4620) );
  AND2_X4 U4575 ( .A1(n3664), .A2(n4382), .ZN(n3753) );
  INV_X1 U4576 ( .A(EBX_REG_1__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U4577 ( .A1(n3753), .A2(n6139), .ZN(n3668) );
  NAND2_X1 U4578 ( .A1(n3755), .A2(n4486), .ZN(n3666) );
  OAI211_X1 U4579 ( .C1(n5485), .C2(EBX_REG_1__SCAN_IN), .A(n3666), .B(n3764), 
        .ZN(n3667) );
  INV_X1 U4581 ( .A(n3672), .ZN(n3673) );
  NAND2_X1 U4582 ( .A1(n3755), .A2(EBX_REG_0__SCAN_IN), .ZN(n3671) );
  INV_X1 U4583 ( .A(EBX_REG_0__SCAN_IN), .ZN(n3669) );
  NAND2_X1 U4584 ( .A1(n3764), .A2(n3669), .ZN(n3670) );
  XNOR2_X1 U4585 ( .A(n3103), .B(n3672), .ZN(n4383) );
  AND2_X2 U4586 ( .A1(n4383), .A2(n4382), .ZN(n6134) );
  NOR2_X2 U4587 ( .A1(n3673), .A2(n6134), .ZN(n4434) );
  INV_X1 U4588 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4439) );
  NAND2_X1 U4589 ( .A1(n3753), .A2(n4439), .ZN(n3676) );
  INV_X1 U4590 ( .A(n3755), .ZN(n3745) );
  INV_X1 U4591 ( .A(n4382), .ZN(n3705) );
  OR2_X1 U4592 ( .A1(n3755), .A2(n4439), .ZN(n3675) );
  NAND2_X1 U4593 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n3705), .ZN(n3674)
         );
  NAND4_X1 U4594 ( .A1(n3676), .A2(n3748), .A3(n3675), .A4(n3674), .ZN(n4433)
         );
  NAND2_X1 U4595 ( .A1(n4434), .A2(n4433), .ZN(n4441) );
  NAND2_X1 U4596 ( .A1(n3764), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3677)
         );
  OAI211_X1 U4597 ( .C1(n3705), .C2(EBX_REG_3__SCAN_IN), .A(n3755), .B(n3677), 
        .ZN(n3678) );
  OAI21_X1 U4598 ( .B1(n3752), .B2(EBX_REG_3__SCAN_IN), .A(n3678), .ZN(n4442)
         );
  NOR2_X2 U4599 ( .A1(n4441), .A2(n4442), .ZN(n4473) );
  INV_X1 U4600 ( .A(EBX_REG_4__SCAN_IN), .ZN(n3679) );
  NAND2_X1 U4601 ( .A1(n3753), .A2(n3679), .ZN(n3682) );
  NAND2_X1 U4602 ( .A1(n3755), .A2(n6361), .ZN(n3680) );
  OAI211_X1 U4603 ( .C1(n3705), .C2(EBX_REG_4__SCAN_IN), .A(n3680), .B(n3764), 
        .ZN(n3681) );
  NAND2_X1 U4604 ( .A1(n3682), .A2(n3681), .ZN(n4474) );
  INV_X1 U4606 ( .A(EBX_REG_6__SCAN_IN), .ZN(n3683) );
  NAND2_X1 U4607 ( .A1(n3753), .A2(n3683), .ZN(n3686) );
  NAND2_X1 U4608 ( .A1(n3755), .A2(n6752), .ZN(n3684) );
  OAI211_X1 U4609 ( .C1(n3705), .C2(EBX_REG_6__SCAN_IN), .A(n3684), .B(n3764), 
        .ZN(n3685) );
  NAND2_X1 U4610 ( .A1(n3686), .A2(n3685), .ZN(n4357) );
  NOR2_X1 U4611 ( .A1(n3752), .A2(EBX_REG_7__SCAN_IN), .ZN(n3687) );
  AOI21_X1 U4612 ( .B1(EBX_REG_7__SCAN_IN), .B2(n5616), .A(n3687), .ZN(n3688)
         );
  OAI21_X1 U4613 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n5486), .A(n3688), 
        .ZN(n4715) );
  INV_X1 U4615 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U4616 ( .A1(n3753), .A2(n6066), .ZN(n3691) );
  NAND2_X1 U4617 ( .A1(n3755), .A2(n6799), .ZN(n3689) );
  OAI211_X1 U4618 ( .C1(n3705), .C2(EBX_REG_8__SCAN_IN), .A(n3689), .B(n3764), 
        .ZN(n3690) );
  NAND2_X1 U4619 ( .A1(n3691), .A2(n3690), .ZN(n4962) );
  NOR2_X1 U4620 ( .A1(n3752), .A2(EBX_REG_9__SCAN_IN), .ZN(n3692) );
  AOI21_X1 U4621 ( .B1(n5616), .B2(EBX_REG_9__SCAN_IN), .A(n3692), .ZN(n3693)
         );
  OAI21_X1 U4622 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n5486), .A(n3693), 
        .ZN(n5062) );
  NOR2_X4 U4623 ( .A1(n5061), .A2(n5062), .ZN(n5225) );
  INV_X1 U4624 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5244) );
  NAND2_X1 U4625 ( .A1(n3753), .A2(n5244), .ZN(n3696) );
  OR2_X1 U4626 ( .A1(n3755), .A2(n5244), .ZN(n3695) );
  NAND2_X1 U4627 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n3705), .ZN(n3694) );
  NAND4_X1 U4628 ( .A1(n3696), .A2(n3748), .A3(n3695), .A4(n3694), .ZN(n5226)
         );
  INV_X1 U4629 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5238) );
  NAND2_X1 U4630 ( .A1(n4382), .A2(n5238), .ZN(n3697) );
  OAI211_X1 U4631 ( .C1(n5616), .C2(n6312), .A(n3697), .B(n3755), .ZN(n3698)
         );
  OAI21_X1 U4632 ( .B1(n3752), .B2(EBX_REG_11__SCAN_IN), .A(n3698), .ZN(n5218)
         );
  NOR2_X2 U4633 ( .A1(n5224), .A2(n5218), .ZN(n5259) );
  INV_X1 U4634 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5264) );
  NAND2_X1 U4635 ( .A1(n3753), .A2(n5264), .ZN(n3701) );
  OR2_X1 U4636 ( .A1(n3755), .A2(n5264), .ZN(n3700) );
  NAND2_X1 U4637 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n3705), .ZN(n3699) );
  NAND4_X1 U4638 ( .A1(n3701), .A2(n3748), .A3(n3700), .A4(n3699), .ZN(n5260)
         );
  OAI21_X1 U4639 ( .B1(n5616), .B2(n3539), .A(n3755), .ZN(n3703) );
  NOR2_X1 U4640 ( .A1(n3705), .A2(EBX_REG_13__SCAN_IN), .ZN(n3702) );
  OAI22_X1 U4641 ( .A1(n3703), .A2(n3702), .B1(EBX_REG_13__SCAN_IN), .B2(n3752), .ZN(n5311) );
  INV_X1 U4642 ( .A(EBX_REG_14__SCAN_IN), .ZN(n3704) );
  NAND2_X1 U4643 ( .A1(n3753), .A2(n3704), .ZN(n3708) );
  OR2_X1 U4644 ( .A1(n3755), .A2(n3704), .ZN(n3707) );
  NAND2_X1 U4645 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n3705), .ZN(n3706) );
  NAND4_X1 U4646 ( .A1(n3708), .A2(n3748), .A3(n3707), .A4(n3706), .ZN(n5301)
         );
  INV_X1 U4647 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U4648 ( .A1(n4382), .A2(n6160), .ZN(n3709) );
  OAI211_X1 U4649 ( .C1(n5616), .C2(n5790), .A(n3709), .B(n3755), .ZN(n3710)
         );
  OAI21_X1 U4650 ( .B1(n3752), .B2(EBX_REG_15__SCAN_IN), .A(n3710), .ZN(n5385)
         );
  INV_X1 U4651 ( .A(EBX_REG_16__SCAN_IN), .ZN(n3711) );
  NAND2_X1 U4652 ( .A1(n3753), .A2(n3711), .ZN(n3714) );
  OR2_X1 U4653 ( .A1(n3755), .A2(n3711), .ZN(n3713) );
  NAND2_X1 U4654 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n3705), .ZN(n3712) );
  NAND4_X1 U4655 ( .A1(n3714), .A2(n3748), .A3(n3713), .A4(n3712), .ZN(n5632)
         );
  NAND2_X2 U4656 ( .A1(n5631), .A2(n5632), .ZN(n5951) );
  NAND2_X1 U4657 ( .A1(n3764), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3715) );
  OAI211_X1 U4658 ( .C1(n3705), .C2(EBX_REG_17__SCAN_IN), .A(n3755), .B(n3715), 
        .ZN(n3716) );
  OAI21_X1 U4659 ( .B1(n3752), .B2(EBX_REG_17__SCAN_IN), .A(n3716), .ZN(n5952)
         );
  NOR2_X4 U4660 ( .A1(n5951), .A2(n5952), .ZN(n5950) );
  INV_X1 U4661 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6897) );
  NAND2_X1 U4662 ( .A1(n3753), .A2(n6897), .ZN(n3720) );
  NAND2_X1 U4663 ( .A1(n3755), .A2(n5780), .ZN(n3718) );
  NAND2_X1 U4664 ( .A1(n4382), .A2(n6897), .ZN(n3717) );
  NAND3_X1 U4665 ( .A1(n3718), .A2(n3764), .A3(n3717), .ZN(n3719) );
  NAND2_X1 U4666 ( .A1(n3720), .A2(n3719), .ZN(n5618) );
  NOR2_X1 U4667 ( .A1(n3705), .A2(EBX_REG_20__SCAN_IN), .ZN(n3721) );
  AOI21_X1 U4668 ( .B1(n3771), .B2(n3722), .A(n3721), .ZN(n5607) );
  OR2_X1 U4669 ( .A1(n5486), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3724)
         );
  INV_X1 U4670 ( .A(EBX_REG_18__SCAN_IN), .ZN(n3723) );
  NAND2_X1 U4671 ( .A1(n4382), .A2(n3723), .ZN(n5613) );
  NAND2_X1 U4672 ( .A1(n3724), .A2(n5613), .ZN(n5617) );
  NAND2_X1 U4673 ( .A1(n5616), .A2(EBX_REG_20__SCAN_IN), .ZN(n3726) );
  NAND2_X1 U4674 ( .A1(n5617), .A2(n3764), .ZN(n3725) );
  OAI211_X1 U4675 ( .C1(n5607), .C2(n5617), .A(n3726), .B(n3725), .ZN(n3727)
         );
  OR2_X1 U4676 ( .A1(n5486), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3729)
         );
  NAND2_X1 U4677 ( .A1(n5616), .A2(EBX_REG_21__SCAN_IN), .ZN(n3728) );
  OAI211_X1 U4678 ( .C1(n3752), .C2(EBX_REG_21__SCAN_IN), .A(n3729), .B(n3728), 
        .ZN(n5597) );
  OR2_X1 U4679 ( .A1(n5486), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3732)
         );
  INV_X1 U4680 ( .A(n3752), .ZN(n3821) );
  INV_X1 U4681 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5591) );
  NAND2_X1 U4682 ( .A1(n3821), .A2(n5591), .ZN(n3731) );
  NAND2_X1 U4683 ( .A1(n5616), .A2(EBX_REG_23__SCAN_IN), .ZN(n3730) );
  AND3_X1 U4684 ( .A1(n3732), .A2(n3731), .A3(n3730), .ZN(n5587) );
  INV_X1 U4685 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5858) );
  NAND2_X1 U4686 ( .A1(n3753), .A2(n5858), .ZN(n3735) );
  NAND2_X1 U4687 ( .A1(n3745), .A2(EBX_REG_22__SCAN_IN), .ZN(n3734) );
  NAND2_X1 U4688 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n5485), .ZN(n3733) );
  NAND4_X1 U4689 ( .A1(n3735), .A2(n3748), .A3(n3734), .A4(n3733), .ZN(n5588)
         );
  AND2_X1 U4690 ( .A1(n5587), .A2(n5588), .ZN(n3736) );
  INV_X1 U4691 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U4692 ( .A1(n3753), .A2(n5583), .ZN(n3739) );
  OR2_X1 U4693 ( .A1(n3755), .A2(n5583), .ZN(n3738) );
  NAND2_X1 U4694 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n5485), .ZN(n3737) );
  NAND4_X1 U4695 ( .A1(n3739), .A2(n3748), .A3(n3738), .A4(n3737), .ZN(n5577)
         );
  INV_X1 U4696 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U4697 ( .A1(n3753), .A2(n5581), .ZN(n3742) );
  NAND2_X1 U4698 ( .A1(n3755), .A2(n5728), .ZN(n3740) );
  OAI211_X1 U4699 ( .C1(EBX_REG_25__SCAN_IN), .C2(n3705), .A(n3740), .B(n3764), 
        .ZN(n3741) );
  NAND2_X1 U4700 ( .A1(n3742), .A2(n3741), .ZN(n5576) );
  AND2_X1 U4701 ( .A1(n5577), .A2(n5576), .ZN(n3743) );
  AND2_X2 U4702 ( .A1(n5590), .A2(n3743), .ZN(n5579) );
  INV_X1 U4703 ( .A(EBX_REG_26__SCAN_IN), .ZN(n3744) );
  NAND2_X1 U4704 ( .A1(n3753), .A2(n3744), .ZN(n3749) );
  NAND2_X1 U4705 ( .A1(n3745), .A2(EBX_REG_26__SCAN_IN), .ZN(n3747) );
  NAND2_X1 U4706 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n5485), .ZN(n3746) );
  NAND4_X1 U4707 ( .A1(n3749), .A2(n3748), .A3(n3747), .A4(n3746), .ZN(n4249)
         );
  NAND2_X1 U4708 ( .A1(n5579), .A2(n4249), .ZN(n5556) );
  OR2_X1 U4709 ( .A1(n5486), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3751)
         );
  NAND2_X1 U4710 ( .A1(n5616), .A2(EBX_REG_27__SCAN_IN), .ZN(n3750) );
  OAI211_X1 U4711 ( .C1(n3752), .C2(EBX_REG_27__SCAN_IN), .A(n3751), .B(n3750), 
        .ZN(n5555) );
  NOR2_X2 U4712 ( .A1(n5556), .A2(n5555), .ZN(n5558) );
  INV_X1 U4713 ( .A(EBX_REG_28__SCAN_IN), .ZN(n3756) );
  NAND2_X1 U4714 ( .A1(n3753), .A2(n3756), .ZN(n3760) );
  INV_X1 U4715 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3754) );
  NAND2_X1 U4716 ( .A1(n3755), .A2(n3754), .ZN(n3758) );
  NAND2_X1 U4717 ( .A1(n4382), .A2(n3756), .ZN(n3757) );
  NAND3_X1 U4718 ( .A1(n3758), .A2(n3764), .A3(n3757), .ZN(n3759) );
  NAND2_X1 U4719 ( .A1(n3760), .A2(n3759), .ZN(n5362) );
  INV_X1 U4720 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3815) );
  AND2_X1 U4721 ( .A1(n3771), .A2(n3815), .ZN(n3820) );
  INV_X1 U4722 ( .A(EBX_REG_29__SCAN_IN), .ZN(n6789) );
  AND2_X1 U4723 ( .A1(n4382), .A2(n6789), .ZN(n3761) );
  NOR3_X2 U4724 ( .A1(n3762), .A2(n3820), .A3(n3761), .ZN(n3766) );
  NOR2_X1 U4725 ( .A1(n3766), .A2(n5616), .ZN(n5482) );
  AOI22_X1 U4726 ( .A1(n5486), .A2(EBX_REG_30__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5485), .ZN(n5484) );
  OAI21_X1 U4727 ( .B1(n3766), .B2(n3762), .A(n5484), .ZN(n3767) );
  INV_X1 U4728 ( .A(n3762), .ZN(n3824) );
  INV_X1 U4729 ( .A(n5484), .ZN(n3763) );
  OAI21_X1 U4730 ( .B1(n3824), .B2(n3764), .A(n3763), .ZN(n3765) );
  OAI22_X1 U4731 ( .A1(n5482), .A2(n3767), .B1(n3766), .B2(n3765), .ZN(n5466)
         );
  NOR2_X2 U4732 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6395) );
  AND2_X2 U4733 ( .A1(n4364), .A2(n6910), .ZN(n6340) );
  AND2_X1 U4734 ( .A1(n6340), .A2(REIP_REG_30__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U4735 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U4736 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5229) );
  NOR2_X1 U4737 ( .A1(n5228), .A2(n5229), .ZN(n3787) );
  INV_X1 U4738 ( .A(n4612), .ZN(n5378) );
  AOI21_X1 U4739 ( .B1(n5378), .B2(n3770), .A(n4373), .ZN(n3768) );
  AOI21_X1 U4740 ( .B1(n3769), .B2(n5616), .A(n3768), .ZN(n3775) );
  NAND2_X1 U4741 ( .A1(n3770), .A2(n4580), .ZN(n5251) );
  OR2_X1 U4742 ( .A1(n5251), .A2(n4590), .ZN(n4392) );
  NAND2_X1 U4743 ( .A1(n3771), .A2(n4392), .ZN(n3773) );
  NAND2_X1 U4744 ( .A1(n3773), .A2(n3772), .ZN(n3774) );
  AND3_X1 U4745 ( .A1(n3776), .A2(n3775), .A3(n3774), .ZN(n3777) );
  NAND2_X1 U4746 ( .A1(n3778), .A2(n3777), .ZN(n4406) );
  INV_X1 U4747 ( .A(n3779), .ZN(n3781) );
  OR2_X1 U4748 ( .A1(n3781), .A2(n3780), .ZN(n4505) );
  NAND2_X1 U4749 ( .A1(n3783), .A2(n3782), .ZN(n3784) );
  OAI211_X1 U4750 ( .C1(n4402), .C2(n3222), .A(n4505), .B(n3784), .ZN(n3785)
         );
  NOR2_X1 U4751 ( .A1(n4406), .A2(n3785), .ZN(n3788) );
  NAND2_X1 U4752 ( .A1(n3788), .A2(n3786), .ZN(n5544) );
  INV_X1 U4753 ( .A(n5544), .ZN(n4386) );
  INV_X1 U4754 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6372) );
  OAI21_X1 U4755 ( .B1(n4486), .B2(n6372), .A(n3477), .ZN(n6371) );
  INV_X1 U4756 ( .A(n6371), .ZN(n6352) );
  INV_X1 U4757 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6367) );
  NOR2_X1 U4758 ( .A1(n6367), .A2(n6361), .ZN(n6353) );
  INV_X1 U4759 ( .A(n6353), .ZN(n6343) );
  NOR2_X1 U4760 ( .A1(n6352), .A2(n6343), .ZN(n6339) );
  NAND2_X1 U4761 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6339), .ZN(n6332)
         );
  NOR3_X1 U4762 ( .A1(n6752), .A2(n6329), .A3(n6332), .ZN(n5184) );
  NAND2_X1 U4763 ( .A1(n3787), .A2(n5184), .ZN(n5291) );
  INV_X1 U4764 ( .A(n5291), .ZN(n5298) );
  NAND2_X1 U4765 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6373) );
  NOR4_X1 U4766 ( .A1(n5187), .A2(n6752), .A3(n6373), .A4(n6343), .ZN(n5185)
         );
  NAND2_X1 U4767 ( .A1(n5185), .A2(n3787), .ZN(n5293) );
  AND2_X1 U4768 ( .A1(n5546), .A2(n4580), .ZN(n6498) );
  INV_X1 U4769 ( .A(n3788), .ZN(n3789) );
  AND2_X1 U4770 ( .A1(n3794), .A2(n3789), .ZN(n5299) );
  NOR2_X1 U4771 ( .A1(n5293), .A2(n6369), .ZN(n6299) );
  NAND2_X1 U4772 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6298) );
  INV_X1 U4773 ( .A(n6298), .ZN(n5295) );
  NAND2_X1 U4774 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5295), .ZN(n5389) );
  NOR2_X1 U4775 ( .A1(n5388), .A2(n5389), .ZN(n5386) );
  NAND3_X1 U4776 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5386), .ZN(n3798) );
  INV_X1 U4777 ( .A(n5763), .ZN(n3790) );
  AND2_X1 U4778 ( .A1(n3790), .A2(n5764), .ZN(n5746) );
  NAND2_X1 U4779 ( .A1(n5746), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3791) );
  NOR2_X1 U4780 ( .A1(n5948), .A2(n3791), .ZN(n5745) );
  NAND2_X1 U4781 ( .A1(n5745), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5736) );
  INV_X1 U4782 ( .A(n3803), .ZN(n3792) );
  AND2_X1 U4783 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5727) );
  INV_X1 U4784 ( .A(n5727), .ZN(n3805) );
  NOR2_X1 U4785 ( .A1(n5947), .A2(n3805), .ZN(n5718) );
  INV_X1 U4786 ( .A(n5712), .ZN(n3793) );
  NAND2_X1 U4787 ( .A1(n5718), .A2(n3793), .ZN(n5491) );
  NOR2_X1 U4788 ( .A1(n5491), .A2(n3815), .ZN(n3808) );
  INV_X1 U4789 ( .A(n6330), .ZN(n5186) );
  NAND2_X1 U4790 ( .A1(n5186), .A2(n6329), .ZN(n6331) );
  INV_X1 U4791 ( .A(n6331), .ZN(n5387) );
  AND2_X1 U4792 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5489) );
  NOR2_X1 U4793 ( .A1(n3798), .A2(n5291), .ZN(n5759) );
  OR2_X1 U4794 ( .A1(n3794), .A2(n6340), .ZN(n4429) );
  INV_X1 U4795 ( .A(n6329), .ZN(n6375) );
  NOR2_X1 U4796 ( .A1(n6375), .A2(n5299), .ZN(n5294) );
  OR2_X1 U4797 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5294), .ZN(n4426)
         );
  NAND2_X1 U4798 ( .A1(n4429), .A2(n4426), .ZN(n6328) );
  INV_X1 U4799 ( .A(n6328), .ZN(n3795) );
  NAND2_X1 U4800 ( .A1(n6329), .A2(n3795), .ZN(n5292) );
  INV_X1 U4801 ( .A(n5292), .ZN(n5758) );
  OAI21_X1 U4802 ( .B1(n5759), .B2(n5758), .A(n5746), .ZN(n3797) );
  NAND2_X1 U4803 ( .A1(n5186), .A2(n5758), .ZN(n3796) );
  NAND2_X1 U4804 ( .A1(n3797), .A2(n3796), .ZN(n3799) );
  OAI21_X1 U4805 ( .B1(n5293), .B2(n3798), .A(n6330), .ZN(n5757) );
  NAND2_X1 U4806 ( .A1(n3799), .A2(n5757), .ZN(n5754) );
  INV_X1 U4807 ( .A(n3800), .ZN(n3801) );
  AND2_X1 U4808 ( .A1(n6331), .A2(n3801), .ZN(n3802) );
  AOI21_X1 U4809 ( .B1(n6369), .B2(n6329), .A(n3803), .ZN(n3804) );
  INV_X1 U4810 ( .A(n5941), .ZN(n3807) );
  NAND2_X1 U4811 ( .A1(n6331), .A2(n3805), .ZN(n3806) );
  NAND2_X1 U4812 ( .A1(n3807), .A2(n3806), .ZN(n5723) );
  AOI21_X1 U4813 ( .B1(n6331), .B2(n5712), .A(n5723), .ZN(n3819) );
  OAI21_X1 U4814 ( .B1(n5387), .B2(n5489), .A(n3819), .ZN(n5492) );
  MUX2_X1 U4815 ( .A(n3808), .B(n5492), .S(INSTADDRPOINTER_REG_30__SCAN_IN), 
        .Z(n3809) );
  AOI211_X1 U4816 ( .C1(n6342), .C2(n5466), .A(n5471), .B(n3809), .ZN(n3810)
         );
  OAI21_X1 U4817 ( .B1(n5476), .B2(n6354), .A(n3810), .ZN(U2988) );
  NAND2_X1 U4818 ( .A1(n5479), .A2(n3815), .ZN(n3813) );
  INV_X1 U4819 ( .A(n3811), .ZN(n3812) );
  NAND2_X1 U4820 ( .A1(n3813), .A2(n3812), .ZN(n3818) );
  INV_X1 U4821 ( .A(n3814), .ZN(n3816) );
  NOR3_X1 U4822 ( .A1(n5479), .A2(n3816), .A3(n3815), .ZN(n3817) );
  OR2_X2 U4823 ( .A1(n3818), .A2(n3817), .ZN(n4265) );
  NAND2_X1 U4824 ( .A1(n4265), .A2(n6381), .ZN(n3832) );
  INV_X1 U4825 ( .A(n3819), .ZN(n3830) );
  INV_X1 U4826 ( .A(n3820), .ZN(n3823) );
  AOI22_X1 U4827 ( .A1(n3821), .A2(n6789), .B1(n5616), .B2(EBX_REG_29__SCAN_IN), .ZN(n3822) );
  AND2_X1 U4828 ( .A1(n3823), .A2(n3822), .ZN(n3825) );
  INV_X1 U4829 ( .A(n3825), .ZN(n3826) );
  AND2_X1 U4830 ( .A1(n3762), .A2(n3826), .ZN(n3827) );
  AND2_X1 U4831 ( .A1(n6340), .A2(REIP_REG_29__SCAN_IN), .ZN(n4344) );
  AOI21_X1 U4832 ( .B1(n5812), .B2(n6342), .A(n4344), .ZN(n3828) );
  OAI21_X1 U4833 ( .B1(n5491), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n3828), 
        .ZN(n3829) );
  AOI21_X1 U4834 ( .B1(n3830), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n3829), 
        .ZN(n3831) );
  NAND2_X1 U4835 ( .A1(n3832), .A2(n3831), .ZN(U2989) );
  NOR2_X2 U4836 ( .A1(n4598), .A2(n6647), .ZN(n3988) );
  NAND2_X1 U4837 ( .A1(n4526), .A2(n3988), .ZN(n3837) );
  NOR2_X1 U4838 ( .A1(n4381), .A2(n6647), .ZN(n3833) );
  AOI22_X1 U4839 ( .A1(n5502), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6647), .ZN(n3835) );
  NAND2_X1 U4840 ( .A1(n3841), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3834) );
  AND2_X1 U4841 ( .A1(n3835), .A2(n3834), .ZN(n3836) );
  NAND2_X1 U4842 ( .A1(n3837), .A2(n3836), .ZN(n4369) );
  NAND2_X1 U4843 ( .A1(n3838), .A2(n3261), .ZN(n3839) );
  NAND2_X1 U4844 ( .A1(n3839), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4420) );
  INV_X1 U4845 ( .A(n5252), .ZN(n4867) );
  NAND2_X1 U4846 ( .A1(n5502), .A2(EAX_REG_0__SCAN_IN), .ZN(n3843) );
  NAND2_X1 U4847 ( .A1(n6647), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3842)
         );
  OAI211_X1 U4848 ( .C1(n3863), .C2(n3560), .A(n3843), .B(n3842), .ZN(n3844)
         );
  AOI21_X1 U4849 ( .B1(n4867), .B2(n3988), .A(n3844), .ZN(n4421) );
  OR2_X1 U4850 ( .A1(n4420), .A2(n4421), .ZN(n4422) );
  NOR2_X2 U4851 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n5452) );
  NAND2_X1 U4852 ( .A1(n4421), .A2(n5452), .ZN(n3845) );
  NAND2_X1 U4853 ( .A1(n4422), .A2(n3845), .ZN(n4368) );
  AND2_X2 U4854 ( .A1(n4369), .A2(n4368), .ZN(n4371) );
  NAND2_X1 U4855 ( .A1(n4533), .A2(n3988), .ZN(n3846) );
  NAND2_X1 U4856 ( .A1(n6647), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4191) );
  NAND2_X1 U4857 ( .A1(n3846), .A2(n4191), .ZN(n3849) );
  OR2_X2 U4858 ( .A1(n4371), .A2(n3849), .ZN(n4437) );
  OAI21_X1 U4859 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3853), .ZN(n6297) );
  AOI22_X1 U4860 ( .A1(n5452), .A2(n6297), .B1(n5501), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3848) );
  NAND2_X1 U4861 ( .A1(n5502), .A2(EAX_REG_2__SCAN_IN), .ZN(n3847) );
  OAI211_X1 U4862 ( .C1(n3863), .C2(n5537), .A(n3848), .B(n3847), .ZN(n4436)
         );
  NAND2_X1 U4863 ( .A1(n4437), .A2(n4436), .ZN(n3851) );
  NAND2_X1 U4864 ( .A1(n3849), .A2(n4371), .ZN(n3850) );
  NAND2_X2 U4865 ( .A1(n3851), .A2(n3850), .ZN(n4470) );
  NAND2_X1 U4866 ( .A1(n5800), .A2(n3988), .ZN(n3859) );
  OAI21_X1 U4867 ( .B1(n3854), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n3864), 
        .ZN(n6287) );
  AOI22_X1 U4868 ( .A1(n6287), .A2(n5452), .B1(n5501), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3856) );
  NAND2_X1 U4869 ( .A1(n5502), .A2(EAX_REG_3__SCAN_IN), .ZN(n3855) );
  OAI211_X1 U4870 ( .C1(n3863), .C2(n3116), .A(n3856), .B(n3855), .ZN(n3857)
         );
  INV_X1 U4871 ( .A(n3857), .ZN(n3858) );
  NAND2_X1 U4872 ( .A1(n3860), .A2(n3988), .ZN(n3868) );
  NAND2_X1 U4873 ( .A1(n6647), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3862)
         );
  NAND2_X1 U4874 ( .A1(n5502), .A2(EAX_REG_4__SCAN_IN), .ZN(n3861) );
  OAI211_X1 U4875 ( .C1(n3863), .C2(n5974), .A(n3862), .B(n3861), .ZN(n3866)
         );
  AOI21_X1 U4876 ( .B1(n3864), .B2(n6103), .A(n3869), .ZN(n5170) );
  NOR2_X1 U4877 ( .A1(n5170), .A2(n5449), .ZN(n3865) );
  AOI21_X1 U4878 ( .B1(n3866), .B2(n5449), .A(n3865), .ZN(n3867) );
  NAND3_X2 U4879 ( .A1(n4470), .A2(n4440), .A3(n4469), .ZN(n4617) );
  INV_X1 U4880 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3872) );
  NAND2_X1 U4881 ( .A1(n5501), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3871)
         );
  OAI21_X1 U4882 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n3869), .A(n3875), 
        .ZN(n6279) );
  NAND2_X1 U4883 ( .A1(n6279), .A2(n5452), .ZN(n3870) );
  OAI211_X1 U4884 ( .C1(n4025), .C2(n3872), .A(n3871), .B(n3870), .ZN(n3873)
         );
  AOI21_X1 U4885 ( .B1(n6929), .B2(n3875), .A(n3882), .ZN(n5273) );
  AOI22_X1 U4886 ( .A1(n5502), .A2(EAX_REG_6__SCAN_IN), .B1(n5501), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3876) );
  OAI21_X1 U4887 ( .B1(n5273), .B2(n5449), .A(n3876), .ZN(n3877) );
  OAI21_X1 U4888 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n3882), .A(n3886), 
        .ZN(n6271) );
  NAND2_X1 U4889 ( .A1(n6271), .A2(n5452), .ZN(n3884) );
  AOI22_X1 U4890 ( .A1(n5502), .A2(EAX_REG_7__SCAN_IN), .B1(n5501), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3883) );
  NAND2_X1 U4891 ( .A1(n3884), .A2(n3883), .ZN(n3885) );
  XOR2_X1 U4892 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3900), .Z(n6068) );
  AOI22_X1 U4893 ( .A1(n4315), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4894 ( .A1(n3322), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n5428), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4895 ( .A1(n4320), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4896 ( .A1(n5433), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3887) );
  NAND4_X1 U4897 ( .A1(n3890), .A2(n3889), .A3(n3888), .A4(n3887), .ZN(n3896)
         );
  AOI22_X1 U4898 ( .A1(n5438), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4899 ( .A1(n4295), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4900 ( .A1(n5435), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4901 ( .A1(n5434), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3891) );
  NAND4_X1 U4902 ( .A1(n3894), .A2(n3893), .A3(n3892), .A4(n3891), .ZN(n3895)
         );
  OR2_X1 U4903 ( .A1(n3896), .A2(n3895), .ZN(n3897) );
  AOI22_X1 U4904 ( .A1(n3988), .A2(n3897), .B1(n5501), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3899) );
  NAND2_X1 U4905 ( .A1(n5502), .A2(EAX_REG_8__SCAN_IN), .ZN(n3898) );
  OAI211_X1 U4906 ( .C1(n6068), .C2(n5449), .A(n3899), .B(n3898), .ZN(n4960)
         );
  XNOR2_X1 U4907 ( .A(n3915), .B(n5204), .ZN(n5161) );
  INV_X1 U4908 ( .A(n3988), .ZN(n4010) );
  AOI22_X1 U4909 ( .A1(n3322), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4910 ( .A1(n5428), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5433), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4911 ( .A1(n4295), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4912 ( .A1(n4315), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3901) );
  NAND4_X1 U4913 ( .A1(n3904), .A2(n3903), .A3(n3902), .A4(n3901), .ZN(n3910)
         );
  AOI22_X1 U4914 ( .A1(n4122), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4915 ( .A1(n4320), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5435), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4916 ( .A1(n5438), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4917 ( .A1(n5434), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3905) );
  NAND4_X1 U4918 ( .A1(n3908), .A2(n3907), .A3(n3906), .A4(n3905), .ZN(n3909)
         );
  NOR2_X1 U4919 ( .A1(n3910), .A2(n3909), .ZN(n3913) );
  NAND2_X1 U4920 ( .A1(n5502), .A2(EAX_REG_9__SCAN_IN), .ZN(n3912) );
  NAND2_X1 U4921 ( .A1(n5501), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3911)
         );
  OAI211_X1 U4922 ( .C1(n4010), .C2(n3913), .A(n3912), .B(n3911), .ZN(n3914)
         );
  AOI21_X1 U4923 ( .B1(n5161), .B2(n5452), .A(n3914), .ZN(n5057) );
  NOR2_X2 U4924 ( .A1(n5058), .A2(n5057), .ZN(n5056) );
  XOR2_X1 U4925 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3931), .Z(n6055) );
  INV_X1 U4926 ( .A(n6055), .ZN(n5246) );
  AOI22_X1 U4927 ( .A1(n4315), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4320), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4928 ( .A1(n5434), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5433), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4929 ( .A1(n4295), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4930 ( .A1(n5428), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3916) );
  NAND4_X1 U4931 ( .A1(n3919), .A2(n3918), .A3(n3917), .A4(n3916), .ZN(n3925)
         );
  AOI22_X1 U4932 ( .A1(n5438), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4933 ( .A1(n4122), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4934 ( .A1(n5435), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3921) );
  AOI22_X1 U4935 ( .A1(n4117), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3920) );
  NAND4_X1 U4936 ( .A1(n3923), .A2(n3922), .A3(n3921), .A4(n3920), .ZN(n3924)
         );
  NOR2_X1 U4937 ( .A1(n3925), .A2(n3924), .ZN(n3928) );
  NAND2_X1 U4938 ( .A1(n5502), .A2(EAX_REG_10__SCAN_IN), .ZN(n3927) );
  NAND2_X1 U4939 ( .A1(n5501), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3926)
         );
  OAI211_X1 U4940 ( .C1(n4010), .C2(n3928), .A(n3927), .B(n3926), .ZN(n3929)
         );
  AOI21_X1 U4941 ( .B1(n5246), .B2(n5452), .A(n3929), .ZN(n5212) );
  XNOR2_X1 U4942 ( .A(n3949), .B(n3948), .ZN(n5283) );
  NAND2_X1 U4943 ( .A1(n5283), .A2(n5452), .ZN(n3947) );
  AOI22_X1 U4944 ( .A1(n4320), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4945 ( .A1(n5428), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4946 ( .A1(n4122), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4947 ( .A1(n5433), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3932) );
  NAND4_X1 U4948 ( .A1(n3935), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(n3941)
         );
  AOI22_X1 U4949 ( .A1(n4295), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n5435), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4950 ( .A1(n4315), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3938) );
  AOI22_X1 U4951 ( .A1(n5438), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4952 ( .A1(n5434), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3936) );
  NAND4_X1 U4953 ( .A1(n3939), .A2(n3938), .A3(n3937), .A4(n3936), .ZN(n3940)
         );
  NOR2_X1 U4954 ( .A1(n3941), .A2(n3940), .ZN(n3944) );
  NAND2_X1 U4955 ( .A1(n5502), .A2(EAX_REG_11__SCAN_IN), .ZN(n3943) );
  NAND2_X1 U4956 ( .A1(n5501), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3942)
         );
  OAI211_X1 U4957 ( .C1(n4010), .C2(n3944), .A(n3943), .B(n3942), .ZN(n3945)
         );
  INV_X1 U4958 ( .A(n3945), .ZN(n3946) );
  NAND2_X1 U4959 ( .A1(n3947), .A2(n3946), .ZN(n5214) );
  AND2_X2 U4960 ( .A1(n5210), .A2(n5214), .ZN(n5263) );
  XOR2_X1 U4961 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3964), .Z(n6050) );
  INV_X1 U4962 ( .A(EAX_REG_12__SCAN_IN), .ZN(n3950) );
  INV_X1 U4963 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5317) );
  OAI22_X1 U4964 ( .A1(n4025), .A2(n3950), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5317), .ZN(n3962) );
  AOI22_X1 U4965 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n5428), .B1(n4320), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4966 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n5434), .B1(n5433), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3953) );
  AOI22_X1 U4967 ( .A1(n3101), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5435), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3952) );
  AOI22_X1 U4968 ( .A1(n4315), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3951) );
  NAND4_X1 U4969 ( .A1(n3954), .A2(n3953), .A3(n3952), .A4(n3951), .ZN(n3960)
         );
  AOI22_X1 U4970 ( .A1(n4122), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4295), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4971 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n5438), .B1(n4117), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4972 ( .A1(n3322), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4973 ( .A1(n5427), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3955) );
  NAND4_X1 U4974 ( .A1(n3958), .A2(n3957), .A3(n3956), .A4(n3955), .ZN(n3959)
         );
  OR2_X1 U4975 ( .A1(n3960), .A2(n3959), .ZN(n3961) );
  AOI22_X1 U4976 ( .A1(n3962), .A2(n5449), .B1(n3988), .B2(n3961), .ZN(n3963)
         );
  OAI21_X1 U4977 ( .B1(n6050), .B2(n5449), .A(n3963), .ZN(n5262) );
  XNOR2_X1 U4978 ( .A(n3991), .B(n6037), .ZN(n6040) );
  INV_X1 U4979 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6178) );
  OAI22_X1 U4980 ( .A1(n4025), .A2(n6178), .B1(n4191), .B2(n6037), .ZN(n3965)
         );
  AOI21_X1 U4981 ( .B1(n6040), .B2(n5452), .A(n3965), .ZN(n3979) );
  AOI22_X1 U4982 ( .A1(n5434), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5433), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3969) );
  AOI22_X1 U4983 ( .A1(n4117), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n5435), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4984 ( .A1(n4320), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4985 ( .A1(n5438), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3966) );
  NAND4_X1 U4986 ( .A1(n3969), .A2(n3968), .A3(n3967), .A4(n3966), .ZN(n3975)
         );
  AOI22_X1 U4987 ( .A1(n3322), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5428), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4988 ( .A1(n4315), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4989 ( .A1(n4122), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3971) );
  AOI22_X1 U4990 ( .A1(n4295), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3970) );
  NAND4_X1 U4991 ( .A1(n3973), .A2(n3972), .A3(n3971), .A4(n3970), .ZN(n3974)
         );
  OR2_X1 U4992 ( .A1(n3975), .A2(n3974), .ZN(n3976) );
  NAND2_X1 U4993 ( .A1(n3988), .A2(n3976), .ZN(n5306) );
  INV_X1 U4994 ( .A(n5306), .ZN(n3977) );
  AOI22_X1 U4995 ( .A1(n3322), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n5433), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4996 ( .A1(n4122), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4997 ( .A1(n3346), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4998 ( .A1(n4320), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3980) );
  NAND4_X1 U4999 ( .A1(n3983), .A2(n3982), .A3(n3981), .A4(n3980), .ZN(n3990)
         );
  AOI22_X1 U5000 ( .A1(n4315), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4295), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U5001 ( .A1(n5438), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3986) );
  AOI22_X1 U5002 ( .A1(n5428), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U5003 ( .A1(n3100), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3984) );
  NAND4_X1 U5004 ( .A1(n3987), .A2(n3986), .A3(n3985), .A4(n3984), .ZN(n3989)
         );
  OAI21_X1 U5005 ( .B1(n3990), .B2(n3989), .A(n3988), .ZN(n3994) );
  XNOR2_X1 U5006 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3995), .ZN(n5348)
         );
  AOI22_X1 U5007 ( .A1(n5452), .A2(n5348), .B1(n5501), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3993) );
  NAND2_X1 U5008 ( .A1(n5502), .A2(EAX_REG_14__SCAN_IN), .ZN(n3992) );
  AOI21_X2 U5009 ( .B1(n5334), .B2(n5332), .A(n5333), .ZN(n5331) );
  INV_X1 U5010 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6834) );
  AOI21_X1 U5011 ( .B1(n3996), .B2(n6834), .A(n4044), .ZN(n6031) );
  OR2_X1 U5012 ( .A1(n6031), .A2(n5449), .ZN(n4013) );
  AOI22_X1 U5013 ( .A1(n4122), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U5014 ( .A1(n5438), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5428), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U5015 ( .A1(n4320), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U5016 ( .A1(n3100), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3997) );
  NAND4_X1 U5017 ( .A1(n4000), .A2(n3999), .A3(n3998), .A4(n3997), .ZN(n4006)
         );
  AOI22_X1 U5018 ( .A1(n3322), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U5019 ( .A1(n4295), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U5020 ( .A1(n4315), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U5021 ( .A1(n5433), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4001) );
  NAND4_X1 U5022 ( .A1(n4004), .A2(n4003), .A3(n4002), .A4(n4001), .ZN(n4005)
         );
  NOR2_X1 U5023 ( .A1(n4006), .A2(n4005), .ZN(n4009) );
  NAND2_X1 U5024 ( .A1(n3833), .A2(EAX_REG_15__SCAN_IN), .ZN(n4008) );
  NAND2_X1 U5025 ( .A1(n5501), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4007)
         );
  OAI211_X1 U5026 ( .C1(n4010), .C2(n4009), .A(n4008), .B(n4007), .ZN(n4011)
         );
  INV_X1 U5027 ( .A(n4011), .ZN(n4012) );
  NAND2_X1 U5028 ( .A1(n4013), .A2(n4012), .ZN(n5393) );
  AND2_X2 U5029 ( .A1(n5331), .A2(n5393), .ZN(n5395) );
  XNOR2_X1 U5030 ( .A(n4044), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6021)
         );
  NAND2_X1 U5031 ( .A1(n6021), .A2(n5452), .ZN(n4029) );
  AOI22_X1 U5032 ( .A1(n4320), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U5033 ( .A1(n5434), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5433), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U5034 ( .A1(n4295), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U5035 ( .A1(n5428), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4014) );
  NAND4_X1 U5036 ( .A1(n4017), .A2(n4016), .A3(n4015), .A4(n4014), .ZN(n4023)
         );
  AOI22_X1 U5037 ( .A1(n4122), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U5038 ( .A1(n4315), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U5039 ( .A1(n3322), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U5040 ( .A1(n5438), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4018) );
  NAND4_X1 U5041 ( .A1(n4021), .A2(n4020), .A3(n4019), .A4(n4018), .ZN(n4022)
         );
  OR2_X1 U5042 ( .A1(n4023), .A2(n4022), .ZN(n4027) );
  INV_X1 U5043 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4024) );
  INV_X1 U5044 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6019) );
  OAI22_X1 U5045 ( .A1(n4025), .A2(n4024), .B1(n4191), .B2(n6019), .ZN(n4026)
         );
  AOI21_X1 U5046 ( .B1(n5447), .B2(n4027), .A(n4026), .ZN(n4028) );
  NAND2_X1 U5047 ( .A1(n4029), .A2(n4028), .ZN(n5633) );
  AOI22_X1 U5049 ( .A1(n5438), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U5050 ( .A1(n5428), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3100), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U5051 ( .A1(n4295), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U5052 ( .A1(n3322), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4030) );
  NAND4_X1 U5053 ( .A1(n4033), .A2(n4032), .A3(n4031), .A4(n4030), .ZN(n4039)
         );
  AOI22_X1 U5054 ( .A1(n4315), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4320), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U5055 ( .A1(n4122), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U5056 ( .A1(n4218), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U5057 ( .A1(n5433), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4034) );
  NAND4_X1 U5058 ( .A1(n4037), .A2(n4036), .A3(n4035), .A4(n4034), .ZN(n4038)
         );
  NOR2_X1 U5059 ( .A1(n4039), .A2(n4038), .ZN(n4043) );
  NAND2_X1 U5060 ( .A1(n6647), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4040)
         );
  NAND2_X1 U5061 ( .A1(n5449), .A2(n4040), .ZN(n4041) );
  AOI21_X1 U5062 ( .B1(n3833), .B2(EAX_REG_17__SCAN_IN), .A(n4041), .ZN(n4042)
         );
  OAI21_X1 U5063 ( .B1(n4330), .B2(n4043), .A(n4042), .ZN(n4048) );
  OAI21_X1 U5064 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n4046), .A(n4079), 
        .ZN(n6014) );
  OR2_X1 U5065 ( .A1(n5449), .A2(n6014), .ZN(n4047) );
  NAND2_X1 U5066 ( .A1(n4048), .A2(n4047), .ZN(n5934) );
  AOI22_X1 U5067 ( .A1(n4295), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4320), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4052) );
  AOI22_X1 U5068 ( .A1(n5428), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n5434), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U5069 ( .A1(n4122), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4050) );
  AOI22_X1 U5070 ( .A1(n4314), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4049) );
  NAND4_X1 U5071 ( .A1(n4052), .A2(n4051), .A3(n4050), .A4(n4049), .ZN(n4058)
         );
  AOI22_X1 U5072 ( .A1(n4315), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U5073 ( .A1(n5435), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4055) );
  AOI22_X1 U5074 ( .A1(n5433), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4054) );
  AOI22_X1 U5075 ( .A1(n5438), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4053) );
  NAND4_X1 U5076 ( .A1(n4056), .A2(n4055), .A3(n4054), .A4(n4053), .ZN(n4057)
         );
  NOR2_X1 U5077 ( .A1(n4058), .A2(n4057), .ZN(n4061) );
  INV_X1 U5078 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5698) );
  OAI21_X1 U5079 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5698), .A(n5449), .ZN(
        n4059) );
  AOI21_X1 U5080 ( .B1(n3833), .B2(EAX_REG_18__SCAN_IN), .A(n4059), .ZN(n4060)
         );
  OAI21_X1 U5081 ( .B1(n4330), .B2(n4061), .A(n4060), .ZN(n4063) );
  XNOR2_X1 U5082 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n4079), .ZN(n6003)
         );
  NAND2_X1 U5083 ( .A1(n5452), .A2(n6003), .ZN(n4062) );
  NAND2_X1 U5084 ( .A1(n4063), .A2(n4062), .ZN(n5630) );
  AOI22_X1 U5085 ( .A1(n4315), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U5086 ( .A1(n5438), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U5087 ( .A1(n5428), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3100), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U5088 ( .A1(n3101), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4065) );
  NAND4_X1 U5089 ( .A1(n4068), .A2(n4067), .A3(n4066), .A4(n4065), .ZN(n4074)
         );
  AOI22_X1 U5090 ( .A1(n4122), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4295), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U5091 ( .A1(n4320), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U5092 ( .A1(n5433), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4070) );
  AOI22_X1 U5093 ( .A1(n4218), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4069) );
  NAND4_X1 U5094 ( .A1(n4072), .A2(n4071), .A3(n4070), .A4(n4069), .ZN(n4073)
         );
  NOR2_X1 U5095 ( .A1(n4074), .A2(n4073), .ZN(n4078) );
  INV_X1 U5096 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4075) );
  OAI21_X1 U5097 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4075), .A(n5449), .ZN(
        n4076) );
  AOI21_X1 U5098 ( .B1(n3833), .B2(EAX_REG_19__SCAN_IN), .A(n4076), .ZN(n4077)
         );
  OAI21_X1 U5099 ( .B1(n4330), .B2(n4078), .A(n4077), .ZN(n4082) );
  OAI21_X1 U5100 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n4080), .A(n4113), 
        .ZN(n5930) );
  OR2_X1 U5101 ( .A1(n5449), .A2(n5930), .ZN(n4081) );
  NAND2_X1 U5102 ( .A1(n4082), .A2(n4081), .ZN(n5610) );
  AOI22_X1 U5103 ( .A1(n5438), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4086) );
  AOI22_X1 U5104 ( .A1(n5428), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U5105 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n5433), .B1(n5434), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U5106 ( .A1(n5427), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4083) );
  NAND4_X1 U5107 ( .A1(n4086), .A2(n4085), .A3(n4084), .A4(n4083), .ZN(n4093)
         );
  AOI22_X1 U5108 ( .A1(n4122), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U5109 ( .A1(n4295), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n5435), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U5110 ( .A1(n4315), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U5111 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n4320), .B1(n4087), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4088) );
  NAND4_X1 U5112 ( .A1(n4091), .A2(n4090), .A3(n4089), .A4(n4088), .ZN(n4092)
         );
  NOR2_X1 U5113 ( .A1(n4093), .A2(n4092), .ZN(n4096) );
  INV_X1 U5114 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5875) );
  AOI21_X1 U5115 ( .B1(n5875), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4094) );
  AOI21_X1 U5116 ( .B1(n3833), .B2(EAX_REG_20__SCAN_IN), .A(n4094), .ZN(n4095)
         );
  OAI21_X1 U5117 ( .B1(n4330), .B2(n4096), .A(n4095), .ZN(n4098) );
  XNOR2_X1 U5118 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n4113), .ZN(n5880)
         );
  NAND2_X1 U5119 ( .A1(n5452), .A2(n5880), .ZN(n4097) );
  AND2_X1 U5120 ( .A1(n4098), .A2(n4097), .ZN(n5603) );
  AOI22_X1 U5121 ( .A1(n5438), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5122 ( .A1(n5428), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5433), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4101) );
  AOI22_X1 U5123 ( .A1(n3299), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n5435), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4100) );
  AOI22_X1 U5124 ( .A1(n4320), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4099) );
  NAND4_X1 U5125 ( .A1(n4102), .A2(n4101), .A3(n4100), .A4(n4099), .ZN(n4108)
         );
  AOI22_X1 U5126 ( .A1(n4122), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U5127 ( .A1(n4315), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4105) );
  AOI22_X1 U5128 ( .A1(n3100), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U5129 ( .A1(n4117), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4103) );
  NAND4_X1 U5130 ( .A1(n4106), .A2(n4105), .A3(n4104), .A4(n4103), .ZN(n4107)
         );
  NOR2_X1 U5131 ( .A1(n4108), .A2(n4107), .ZN(n4112) );
  INV_X1 U5132 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6735) );
  OAI21_X1 U5133 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6735), .A(n6647), 
        .ZN(n4109) );
  INV_X1 U5134 ( .A(n4109), .ZN(n4110) );
  AOI21_X1 U5135 ( .B1(n3833), .B2(EAX_REG_21__SCAN_IN), .A(n4110), .ZN(n4111)
         );
  OAI21_X1 U5136 ( .B1(n4330), .B2(n4112), .A(n4111), .ZN(n4116) );
  OAI21_X1 U5137 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n4114), .A(n4180), 
        .ZN(n5874) );
  OR2_X1 U5138 ( .A1(n5874), .A2(n5449), .ZN(n4115) );
  AOI22_X1 U5139 ( .A1(n5438), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4121) );
  AOI22_X1 U5140 ( .A1(n5428), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4120) );
  AOI22_X1 U5141 ( .A1(n3100), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5433), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4119) );
  AOI22_X1 U5142 ( .A1(n5427), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4118) );
  NAND4_X1 U5143 ( .A1(n4121), .A2(n4120), .A3(n4119), .A4(n4118), .ZN(n4128)
         );
  AOI22_X1 U5144 ( .A1(n4122), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U5145 ( .A1(n3299), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5146 ( .A1(n4315), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5147 ( .A1(n4320), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4123) );
  NAND4_X1 U5148 ( .A1(n4126), .A2(n4125), .A3(n4124), .A4(n4123), .ZN(n4127)
         );
  NOR2_X1 U5149 ( .A1(n4128), .A2(n4127), .ZN(n4131) );
  INV_X1 U5150 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5371) );
  AOI21_X1 U5151 ( .B1(n5371), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4129) );
  AOI21_X1 U5152 ( .B1(n3833), .B2(EAX_REG_22__SCAN_IN), .A(n4129), .ZN(n4130)
         );
  OAI21_X1 U5153 ( .B1(n4330), .B2(n4131), .A(n4130), .ZN(n4133) );
  XNOR2_X1 U5154 ( .A(n4180), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5856)
         );
  NAND2_X1 U5155 ( .A1(n5856), .A2(n5452), .ZN(n4132) );
  INV_X1 U5156 ( .A(n5569), .ZN(n4209) );
  AOI22_X1 U5157 ( .A1(n4315), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4320), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4138) );
  AOI22_X1 U5158 ( .A1(n3322), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n5428), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4137) );
  AOI22_X1 U5159 ( .A1(n4295), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U5160 ( .A1(n5434), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4135) );
  NAND4_X1 U5161 ( .A1(n4138), .A2(n4137), .A3(n4136), .A4(n4135), .ZN(n4144)
         );
  AOI22_X1 U5162 ( .A1(n5438), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4142) );
  AOI22_X1 U5163 ( .A1(n4122), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4141) );
  AOI22_X1 U5164 ( .A1(n5435), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4140) );
  AOI22_X1 U5165 ( .A1(n5433), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4139) );
  NAND4_X1 U5166 ( .A1(n4142), .A2(n4141), .A3(n4140), .A4(n4139), .ZN(n4143)
         );
  NOR2_X1 U5167 ( .A1(n4144), .A2(n4143), .ZN(n4196) );
  AOI22_X1 U5168 ( .A1(n4122), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U5169 ( .A1(n4295), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n5435), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U5170 ( .A1(n4315), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4147) );
  AOI22_X1 U5171 ( .A1(n4320), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4146) );
  NAND4_X1 U5172 ( .A1(n4149), .A2(n4148), .A3(n4147), .A4(n4146), .ZN(n4155)
         );
  AOI22_X1 U5173 ( .A1(n5438), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4153) );
  AOI22_X1 U5174 ( .A1(n4117), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5428), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4152) );
  AOI22_X1 U5175 ( .A1(n5434), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5433), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4151) );
  AOI22_X1 U5176 ( .A1(n5427), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4150) );
  NAND4_X1 U5177 ( .A1(n4153), .A2(n4152), .A3(n4151), .A4(n4150), .ZN(n4154)
         );
  NOR2_X1 U5178 ( .A1(n4155), .A2(n4154), .ZN(n4197) );
  OR2_X1 U5179 ( .A1(n4196), .A2(n4197), .ZN(n4210) );
  AOI22_X1 U5180 ( .A1(n4320), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4159) );
  AOI22_X1 U5181 ( .A1(n5428), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n5433), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4158) );
  AOI22_X1 U5182 ( .A1(n4295), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4157) );
  AOI22_X1 U5183 ( .A1(n5435), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4156) );
  NAND4_X1 U5184 ( .A1(n4159), .A2(n4158), .A3(n4157), .A4(n4156), .ZN(n4165)
         );
  AOI22_X1 U5185 ( .A1(n4315), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4163) );
  AOI22_X1 U5186 ( .A1(n5438), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4162) );
  AOI22_X1 U5187 ( .A1(n5434), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4161) );
  AOI22_X1 U5188 ( .A1(n4117), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4160) );
  NAND4_X1 U5189 ( .A1(n4163), .A2(n4162), .A3(n4161), .A4(n4160), .ZN(n4164)
         );
  NOR2_X1 U5190 ( .A1(n4165), .A2(n4164), .ZN(n4212) );
  NOR2_X1 U5191 ( .A1(n4210), .A2(n4212), .ZN(n4188) );
  AOI22_X1 U5192 ( .A1(n4315), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4320), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U5193 ( .A1(n4295), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U5194 ( .A1(n5428), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4167) );
  AOI22_X1 U5195 ( .A1(n5433), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4166) );
  NAND4_X1 U5196 ( .A1(n4169), .A2(n4168), .A3(n4167), .A4(n4166), .ZN(n4176)
         );
  AOI22_X1 U5197 ( .A1(n4122), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4174) );
  AOI22_X1 U5198 ( .A1(n5438), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4173) );
  AOI22_X1 U5199 ( .A1(n3322), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n5435), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4172) );
  AOI22_X1 U5200 ( .A1(n5434), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4171) );
  NAND4_X1 U5201 ( .A1(n4174), .A2(n4173), .A3(n4172), .A4(n4171), .ZN(n4175)
         );
  NOR2_X1 U5202 ( .A1(n4176), .A2(n4175), .ZN(n4211) );
  XNOR2_X1 U5203 ( .A(n4188), .B(n4211), .ZN(n4177) );
  NAND2_X1 U5204 ( .A1(n4177), .A2(n5447), .ZN(n4187) );
  NAND2_X1 U5205 ( .A1(n6647), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4178)
         );
  NAND2_X1 U5206 ( .A1(n5449), .A2(n4178), .ZN(n4179) );
  AOI21_X1 U5207 ( .B1(n3833), .B2(EAX_REG_25__SCAN_IN), .A(n4179), .ZN(n4186)
         );
  NAND2_X1 U5208 ( .A1(n4204), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4182)
         );
  INV_X1 U5209 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4181) );
  NAND2_X1 U5210 ( .A1(n4182), .A2(n4181), .ZN(n4184) );
  AND2_X1 U5211 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4183) );
  AND2_X1 U5212 ( .A1(n4184), .A2(n4238), .ZN(n5830) );
  AND2_X1 U5213 ( .A1(n5830), .A2(n5452), .ZN(n4185) );
  AOI21_X1 U5214 ( .B1(n4187), .B2(n4186), .A(n4185), .ZN(n5571) );
  INV_X1 U5215 ( .A(n5571), .ZN(n4208) );
  NAND2_X1 U5216 ( .A1(n4212), .A2(n4210), .ZN(n4190) );
  INV_X1 U5217 ( .A(n4188), .ZN(n4189) );
  NAND3_X1 U5218 ( .A1(n5447), .A2(n4190), .A3(n4189), .ZN(n4195) );
  INV_X1 U5219 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5414) );
  XNOR2_X1 U5220 ( .A(n4204), .B(n5414), .ZN(n5837) );
  NOR2_X1 U5221 ( .A1(n5837), .A2(n5449), .ZN(n4193) );
  NOR2_X1 U5222 ( .A1(n4191), .A2(n5414), .ZN(n4192) );
  AOI211_X1 U5223 ( .C1(n5502), .C2(EAX_REG_24__SCAN_IN), .A(n4193), .B(n4192), 
        .ZN(n4194) );
  AND2_X1 U5224 ( .A1(n4195), .A2(n4194), .ZN(n5411) );
  XNOR2_X1 U5225 ( .A(n4197), .B(n4196), .ZN(n4201) );
  NAND2_X1 U5226 ( .A1(n6647), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4198)
         );
  NAND2_X1 U5227 ( .A1(n5449), .A2(n4198), .ZN(n4199) );
  AOI21_X1 U5228 ( .B1(n5502), .B2(EAX_REG_23__SCAN_IN), .A(n4199), .ZN(n4200)
         );
  OAI21_X1 U5229 ( .B1(n4330), .B2(n4201), .A(n4200), .ZN(n4207) );
  NOR2_X1 U5230 ( .A1(n4202), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4203)
         );
  OR2_X1 U5231 ( .A1(n4204), .A2(n4203), .ZN(n5852) );
  INV_X1 U5232 ( .A(n5852), .ZN(n4205) );
  NAND2_X1 U5233 ( .A1(n4205), .A2(n5452), .ZN(n4206) );
  NAND2_X1 U5234 ( .A1(n4207), .A2(n4206), .ZN(n5586) );
  OR2_X1 U5235 ( .A1(n5411), .A2(n5586), .ZN(n5570) );
  NOR2_X1 U5236 ( .A1(n4208), .A2(n5570), .ZN(n4231) );
  NOR3_X1 U5237 ( .A1(n4212), .A2(n4211), .A3(n4210), .ZN(n4267) );
  AOI22_X1 U5238 ( .A1(n5438), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3322), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4216) );
  AOI22_X1 U5239 ( .A1(n5428), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4215) );
  AOI22_X1 U5240 ( .A1(n3100), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5433), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4214) );
  AOI22_X1 U5241 ( .A1(n5427), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4213) );
  NAND4_X1 U5242 ( .A1(n4216), .A2(n4215), .A3(n4214), .A4(n4213), .ZN(n4224)
         );
  AOI22_X1 U5243 ( .A1(n3391), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4222) );
  AOI22_X1 U5244 ( .A1(n4295), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4221) );
  AOI22_X1 U5245 ( .A1(n4315), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4220) );
  AOI22_X1 U5246 ( .A1(n4320), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4219) );
  NAND4_X1 U5247 ( .A1(n4222), .A2(n4221), .A3(n4220), .A4(n4219), .ZN(n4223)
         );
  OR2_X1 U5248 ( .A1(n4224), .A2(n4223), .ZN(n4266) );
  INV_X1 U5249 ( .A(n4266), .ZN(n4225) );
  XNOR2_X1 U5250 ( .A(n4267), .B(n4225), .ZN(n4226) );
  NAND2_X1 U5251 ( .A1(n4226), .A2(n5447), .ZN(n4230) );
  INV_X1 U5252 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4256) );
  AOI21_X1 U5253 ( .B1(n4256), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4227) );
  AOI21_X1 U5254 ( .B1(n3833), .B2(EAX_REG_26__SCAN_IN), .A(n4227), .ZN(n4229)
         );
  XNOR2_X1 U5255 ( .A(n4238), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5656)
         );
  AND2_X1 U5256 ( .A1(n5656), .A2(n5452), .ZN(n4228) );
  AOI21_X1 U5257 ( .B1(n4230), .B2(n4229), .A(n4228), .ZN(n4233) );
  AND2_X1 U5258 ( .A1(n4233), .A2(n4231), .ZN(n4232) );
  NAND2_X1 U5259 ( .A1(n5596), .A2(n4287), .ZN(n5551) );
  INV_X1 U5260 ( .A(n4234), .ZN(n5539) );
  INV_X1 U5261 ( .A(n5541), .ZN(n5545) );
  AND3_X1 U5262 ( .A1(n5546), .A2(n6525), .A3(n5545), .ZN(n5811) );
  INV_X1 U5263 ( .A(n5811), .ZN(n4235) );
  NOR2_X1 U5264 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6651) );
  NAND2_X1 U5265 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6651), .ZN(n6531) );
  NOR2_X1 U5266 ( .A1(n6910), .A2(n6531), .ZN(n6526) );
  NAND2_X1 U5267 ( .A1(n6910), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6546) );
  INV_X1 U5268 ( .A(n6546), .ZN(n4339) );
  AND2_X1 U5269 ( .A1(n4339), .A2(n5452), .ZN(n6541) );
  NOR2_X1 U5270 ( .A1(n6526), .A2(n4236), .ZN(n4237) );
  INV_X1 U5271 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4281) );
  INV_X1 U5272 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4303) );
  NAND2_X1 U5273 ( .A1(n4332), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5451)
         );
  INV_X1 U5274 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5459) );
  INV_X1 U5275 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5517) );
  NOR2_X1 U5276 ( .A1(n5508), .A2(n6537), .ZN(n4240) );
  INV_X1 U5277 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6601) );
  INV_X1 U5278 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6786) );
  NAND2_X1 U5279 ( .A1(n3646), .A2(n6735), .ZN(n4253) );
  INV_X1 U5280 ( .A(n4253), .ZN(n4252) );
  NAND3_X1 U5281 ( .A1(n4241), .A2(n4586), .A3(n4252), .ZN(n4242) );
  INV_X1 U5282 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6582) );
  INV_X1 U5283 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6725) );
  INV_X1 U5284 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6572) );
  NAND3_X1 U5285 ( .A1(REIP_REG_2__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .ZN(n6092) );
  NOR3_X1 U5286 ( .A1(n6725), .A2(n6572), .A3(n6092), .ZN(n4350) );
  NAND4_X1 U5287 ( .A1(REIP_REG_6__SCAN_IN), .A2(n4350), .A3(
        REIP_REG_8__SCAN_IN), .A4(REIP_REG_7__SCAN_IN), .ZN(n5159) );
  NAND2_X1 U5288 ( .A1(REIP_REG_9__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .ZN(
        n5235) );
  NOR3_X1 U5289 ( .A1(n6582), .A2(n5159), .A3(n5235), .ZN(n4245) );
  NAND3_X1 U5290 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        REIP_REG_12__SCAN_IN), .ZN(n4246) );
  INV_X1 U5291 ( .A(n4246), .ZN(n4243) );
  NAND2_X1 U5292 ( .A1(n4245), .A2(n4243), .ZN(n4244) );
  NAND4_X1 U5293 ( .A1(n6015), .A2(REIP_REG_17__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .A4(REIP_REG_15__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U5294 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5884) );
  NOR2_X1 U5295 ( .A1(n6001), .A2(n5884), .ZN(n5877) );
  NAND2_X1 U5296 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5877), .ZN(n5855) );
  NAND3_X1 U5297 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        n5860), .ZN(n5832) );
  NOR2_X1 U5298 ( .A1(n6601), .A2(n5832), .ZN(n5829) );
  AOI21_X1 U5299 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5829), .A(
        REIP_REG_26__SCAN_IN), .ZN(n4247) );
  INV_X1 U5300 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6896) );
  NAND2_X1 U5301 ( .A1(n4245), .A2(n6148), .ZN(n5236) );
  NOR2_X1 U5302 ( .A1(n4246), .A2(n5236), .ZN(n5345) );
  NAND4_X1 U5303 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .A4(n5345), .ZN(n5885) );
  NOR3_X1 U5304 ( .A1(n6896), .A2(n5884), .A3(n5885), .ZN(n5853) );
  NAND4_X1 U5305 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5853), .ZN(n5831) );
  NAND3_X1 U5306 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U5307 ( .A1(n6110), .A2(n6148), .ZN(n5886) );
  OAI21_X1 U5308 ( .B1(n5831), .B2(n5462), .A(n5886), .ZN(n5554) );
  OAI22_X1 U5309 ( .A1(n5655), .A2(n5890), .B1(n4247), .B2(n5554), .ZN(n4248)
         );
  OR2_X1 U5310 ( .A1(n5579), .A2(n4249), .ZN(n4250) );
  NAND2_X1 U5311 ( .A1(n5556), .A2(n4250), .ZN(n5726) );
  NAND2_X1 U5312 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4253), .ZN(n4251) );
  NOR2_X2 U5313 ( .A1(n6131), .A2(n3705), .ZN(n6083) );
  NAND2_X1 U5314 ( .A1(n4447), .A2(n4252), .ZN(n6528) );
  INV_X1 U5315 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5565) );
  AND3_X1 U5316 ( .A1(n4586), .A2(n4253), .A3(n5565), .ZN(n4254) );
  AOI21_X1 U5317 ( .B1(n6648), .B2(n6528), .A(n4254), .ZN(n4255) );
  OAI22_X1 U5318 ( .A1(n3744), .A2(n6138), .B1(n4256), .B2(n6105), .ZN(n4257)
         );
  INV_X1 U5319 ( .A(n4257), .ZN(n4260) );
  NAND2_X1 U5320 ( .A1(n4265), .A2(n6293), .ZN(n4348) );
  NAND2_X1 U5321 ( .A1(n4267), .A2(n4266), .ZN(n4289) );
  AOI22_X1 U5322 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4117), .B1(n3322), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4271) );
  AOI22_X1 U5323 ( .A1(n3391), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4270) );
  AOI22_X1 U5324 ( .A1(n5435), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4269) );
  AOI22_X1 U5325 ( .A1(n5433), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4268) );
  NAND4_X1 U5326 ( .A1(n4271), .A2(n4270), .A3(n4269), .A4(n4268), .ZN(n4277)
         );
  AOI22_X1 U5327 ( .A1(n4315), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3299), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4275) );
  AOI22_X1 U5328 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n5438), .B1(n5428), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4274) );
  AOI22_X1 U5329 ( .A1(n4320), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4273) );
  AOI22_X1 U5330 ( .A1(n3100), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4272) );
  NAND4_X1 U5331 ( .A1(n4275), .A2(n4274), .A3(n4273), .A4(n4272), .ZN(n4276)
         );
  NOR2_X1 U5332 ( .A1(n4277), .A2(n4276), .ZN(n4290) );
  XNOR2_X1 U5333 ( .A(n4289), .B(n4290), .ZN(n4280) );
  OAI21_X1 U5334 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4281), .A(n5449), .ZN(
        n4278) );
  AOI21_X1 U5335 ( .B1(n5502), .B2(EAX_REG_27__SCAN_IN), .A(n4278), .ZN(n4279)
         );
  OAI21_X1 U5336 ( .B1(n4280), .B2(n4330), .A(n4279), .ZN(n4286) );
  NAND2_X1 U5337 ( .A1(n4282), .A2(n4281), .ZN(n4283) );
  NAND2_X1 U5338 ( .A1(n4307), .A2(n4283), .ZN(n5648) );
  INV_X1 U5339 ( .A(n5648), .ZN(n4284) );
  NAND2_X1 U5340 ( .A1(n4284), .A2(n5452), .ZN(n4285) );
  NAND2_X1 U5341 ( .A1(n4286), .A2(n4285), .ZN(n5550) );
  NOR2_X1 U5342 ( .A1(n4290), .A2(n4289), .ZN(n4313) );
  AOI22_X1 U5343 ( .A1(n5438), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4294) );
  AOI22_X1 U5344 ( .A1(n5428), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4293) );
  AOI22_X1 U5345 ( .A1(n3100), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5433), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4292) );
  AOI22_X1 U5346 ( .A1(n5427), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4291) );
  NAND4_X1 U5347 ( .A1(n4294), .A2(n4293), .A3(n4292), .A4(n4291), .ZN(n4302)
         );
  AOI22_X1 U5348 ( .A1(n3391), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4300) );
  AOI22_X1 U5349 ( .A1(n4295), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n5435), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4299) );
  AOI22_X1 U5350 ( .A1(n4315), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4298) );
  AOI22_X1 U5351 ( .A1(n4320), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4297) );
  NAND4_X1 U5352 ( .A1(n4300), .A2(n4299), .A3(n4298), .A4(n4297), .ZN(n4301)
         );
  OR2_X1 U5353 ( .A1(n4302), .A2(n4301), .ZN(n4312) );
  XNOR2_X1 U5354 ( .A(n4313), .B(n4312), .ZN(n4306) );
  OAI21_X1 U5355 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4303), .A(n5449), .ZN(
        n4304) );
  AOI21_X1 U5356 ( .B1(n5502), .B2(EAX_REG_28__SCAN_IN), .A(n4304), .ZN(n4305)
         );
  OAI21_X1 U5357 ( .B1(n4306), .B2(n4330), .A(n4305), .ZN(n4309) );
  XNOR2_X1 U5358 ( .A(n4307), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5822)
         );
  NAND2_X1 U5359 ( .A1(n5822), .A2(n5452), .ZN(n4308) );
  NAND2_X1 U5360 ( .A1(n4309), .A2(n4308), .ZN(n5498) );
  INV_X1 U5361 ( .A(n5498), .ZN(n4310) );
  AND2_X1 U5362 ( .A1(n5355), .A2(n4310), .ZN(n4311) );
  AND2_X2 U5363 ( .A1(n5373), .A2(n4311), .ZN(n5356) );
  NAND2_X1 U5364 ( .A1(n4313), .A2(n4312), .ZN(n5425) );
  AOI22_X1 U5365 ( .A1(n5438), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4319) );
  AOI22_X1 U5366 ( .A1(n3100), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5433), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4318) );
  AOI22_X1 U5367 ( .A1(n4315), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4317) );
  AOI22_X1 U5368 ( .A1(n5428), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4316) );
  NAND4_X1 U5369 ( .A1(n4319), .A2(n4318), .A3(n4317), .A4(n4316), .ZN(n4326)
         );
  AOI22_X1 U5370 ( .A1(n3391), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3299), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4324) );
  AOI22_X1 U5371 ( .A1(n3346), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4323) );
  AOI22_X1 U5372 ( .A1(n4320), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4322) );
  AOI22_X1 U5373 ( .A1(n3370), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4321) );
  NAND4_X1 U5374 ( .A1(n4324), .A2(n4323), .A3(n4322), .A4(n4321), .ZN(n4325)
         );
  NOR2_X1 U5375 ( .A1(n4326), .A2(n4325), .ZN(n5426) );
  XNOR2_X1 U5376 ( .A(n5425), .B(n5426), .ZN(n4331) );
  NAND2_X1 U5377 ( .A1(n6647), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4327)
         );
  NAND2_X1 U5378 ( .A1(n5449), .A2(n4327), .ZN(n4328) );
  AOI21_X1 U5379 ( .B1(n5502), .B2(EAX_REG_29__SCAN_IN), .A(n4328), .ZN(n4329)
         );
  OAI21_X1 U5380 ( .B1(n4331), .B2(n4330), .A(n4329), .ZN(n4337) );
  INV_X1 U5381 ( .A(n4332), .ZN(n4334) );
  INV_X1 U5382 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4333) );
  NAND2_X1 U5383 ( .A1(n4334), .A2(n4333), .ZN(n4335) );
  NAND2_X1 U5384 ( .A1(n5451), .A2(n4335), .ZN(n5816) );
  NOR2_X1 U5385 ( .A1(n5356), .A2(n5496), .ZN(n4338) );
  INV_X1 U5386 ( .A(n5424), .ZN(n5898) );
  NAND3_X1 U5387 ( .A1(n4339), .A2(n6395), .A3(STATEBS16_REG_SCAN_IN), .ZN(
        n6266) );
  INV_X1 U5388 ( .A(n6395), .ZN(n6392) );
  NAND2_X1 U5389 ( .A1(n6392), .A2(n4340), .ZN(n6642) );
  NAND2_X1 U5390 ( .A1(n6642), .A2(n6910), .ZN(n4341) );
  NAND2_X1 U5391 ( .A1(n6910), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4343) );
  NAND2_X1 U5392 ( .A1(n6735), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4342) );
  AND2_X1 U5393 ( .A1(n4343), .A2(n4342), .ZN(n4563) );
  AOI21_X1 U5394 ( .B1(n6288), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n4344), 
        .ZN(n4345) );
  OAI21_X1 U5395 ( .B1(n6296), .B2(n5816), .A(n4345), .ZN(n4346) );
  AOI21_X1 U5396 ( .B1(n5898), .B2(n3099), .A(n4346), .ZN(n4347) );
  NAND2_X1 U5397 ( .A1(n4348), .A2(n4347), .ZN(U2957) );
  NOR2_X1 U5398 ( .A1(n6110), .A2(n6092), .ZN(n6095) );
  INV_X1 U5399 ( .A(n6095), .ZN(n4349) );
  NOR2_X1 U5400 ( .A1(n4349), .A2(n6725), .ZN(n6089) );
  NAND2_X1 U5401 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6089), .ZN(n6074) );
  NOR2_X1 U5402 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6074), .ZN(n4362) );
  INV_X1 U5403 ( .A(n6110), .ZN(n6121) );
  INV_X1 U5404 ( .A(n4350), .ZN(n4351) );
  NAND2_X1 U5405 ( .A1(n6121), .A2(n4351), .ZN(n4352) );
  AND2_X1 U5406 ( .A1(n4352), .A2(n6148), .ZN(n6087) );
  INV_X1 U5407 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6574) );
  AOI22_X1 U5408 ( .A1(EBX_REG_6__SCAN_IN), .A2(n6115), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6130), .ZN(n4353) );
  NAND2_X1 U5409 ( .A1(n6148), .A2(n4364), .ZN(n6085) );
  OAI211_X1 U5410 ( .C1(n6087), .C2(n6574), .A(n4353), .B(n6085), .ZN(n4361)
         );
  OAI21_X1 U5411 ( .B1(n4617), .B2(n4616), .A(n4354), .ZN(n4356) );
  NAND2_X1 U5412 ( .A1(n4356), .A2(n4711), .ZN(n5278) );
  NOR2_X1 U5413 ( .A1(n5278), .A2(n5890), .ZN(n4360) );
  XNOR2_X1 U5414 ( .A(n4357), .B(n4618), .ZN(n4622) );
  NAND2_X1 U5415 ( .A1(n5273), .A2(n6133), .ZN(n4358) );
  OAI21_X1 U5416 ( .B1(n6120), .B2(n4622), .A(n4358), .ZN(n4359) );
  OR4_X1 U5417 ( .A1(n4362), .A2(n4361), .A3(n4360), .A4(n4359), .ZN(U2821) );
  INV_X1 U5418 ( .A(n6644), .ZN(n4367) );
  INV_X1 U5419 ( .A(n5251), .ZN(n4363) );
  OR2_X1 U5420 ( .A1(n6648), .A2(n4363), .ZN(n5548) );
  INV_X1 U5421 ( .A(n4364), .ZN(n4365) );
  AND2_X1 U5422 ( .A1(n6198), .A2(n4365), .ZN(n5809) );
  NOR2_X1 U5423 ( .A1(n5811), .A2(READREQUEST_REG_SCAN_IN), .ZN(n4366) );
  AOI22_X1 U5424 ( .A1(n4367), .A2(n5548), .B1(n5809), .B2(n4366), .ZN(U3474)
         );
  NOR2_X1 U5425 ( .A1(n4369), .A2(n4368), .ZN(n4370) );
  OR2_X1 U5426 ( .A1(n4371), .A2(n4370), .ZN(n6144) );
  NOR2_X1 U5427 ( .A1(n5544), .A2(n6539), .ZN(n4372) );
  NAND2_X1 U5428 ( .A1(n6532), .A2(n4372), .ZN(n4380) );
  INV_X1 U5429 ( .A(n3245), .ZN(n4377) );
  AND3_X1 U5430 ( .A1(n4374), .A2(n4373), .A3(n6537), .ZN(n4375) );
  NAND4_X1 U5431 ( .A1(n4377), .A2(n4376), .A3(n3833), .A4(n4375), .ZN(n4607)
         );
  INV_X1 U5432 ( .A(n4607), .ZN(n4378) );
  NAND2_X1 U5433 ( .A1(n4378), .A2(n4382), .ZN(n4379) );
  NAND2_X1 U5434 ( .A1(n6159), .A2(n4381), .ZN(n5601) );
  NOR2_X1 U5435 ( .A1(n4383), .A2(n4382), .ZN(n4384) );
  OR2_X1 U5436 ( .A1(n6134), .A2(n4384), .ZN(n4480) );
  AOI22_X1 U5437 ( .A1(n6155), .A2(n4480), .B1(n5620), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4385) );
  OAI21_X1 U5438 ( .B1(n6144), .B2(n5601), .A(n4385), .ZN(U2858) );
  NAND2_X1 U5439 ( .A1(n6532), .A2(n4386), .ZN(n4387) );
  OAI21_X1 U5440 ( .B1(n6532), .B2(n5540), .A(n4387), .ZN(n4397) );
  NOR2_X1 U5441 ( .A1(n3705), .A2(READY_N), .ZN(n4388) );
  NAND2_X1 U5442 ( .A1(n4401), .A2(n4388), .ZN(n4605) );
  NAND2_X1 U5443 ( .A1(n4447), .A2(n3646), .ZN(n4389) );
  NAND2_X1 U5444 ( .A1(n4605), .A2(n4389), .ZN(n4390) );
  OAI21_X1 U5445 ( .B1(n6498), .B2(n4401), .A(n4390), .ZN(n4391) );
  NOR2_X1 U5446 ( .A1(n6532), .A2(n4391), .ZN(n4396) );
  INV_X1 U5447 ( .A(n4606), .ZN(n4394) );
  OAI211_X1 U5448 ( .C1(n3655), .C2(n4394), .A(n4393), .B(n4392), .ZN(n4395)
         );
  NOR2_X1 U5449 ( .A1(n6537), .A2(n6647), .ZN(n4530) );
  NAND2_X1 U5450 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4530), .ZN(n4524) );
  INV_X1 U5451 ( .A(n4524), .ZN(n6622) );
  AOI22_X1 U5452 ( .A1(n6525), .A2(n6499), .B1(FLUSH_REG_SCAN_IN), .B2(n6622), 
        .ZN(n5976) );
  NAND2_X1 U5453 ( .A1(n6910), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4539) );
  NAND2_X1 U5454 ( .A1(n5976), .A2(n4539), .ZN(n6630) );
  INV_X1 U5455 ( .A(n4399), .ZN(n4410) );
  NAND2_X1 U5456 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5530) );
  OAI22_X1 U5457 ( .A1(n4486), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n5480), .B2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5529) );
  INV_X1 U5458 ( .A(n5972), .ZN(n6628) );
  INV_X1 U5459 ( .A(n6136), .ZN(n4660) );
  INV_X1 U5460 ( .A(n4401), .ZN(n4403) );
  NAND4_X1 U5461 ( .A1(n3655), .A2(n4404), .A3(n4403), .A4(n4402), .ZN(n4405)
         );
  OR2_X1 U5462 ( .A1(n4406), .A2(n4405), .ZN(n4502) );
  INV_X1 U5463 ( .A(n6498), .ZN(n4445) );
  NOR2_X1 U5464 ( .A1(n4445), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4409)
         );
  NOR3_X1 U5465 ( .A1(n4413), .A2(n5528), .A3(n4407), .ZN(n4408) );
  AOI211_X1 U5466 ( .C1(n4660), .C2(n4502), .A(n4409), .B(n4408), .ZN(n6500)
         );
  OAI222_X1 U5467 ( .A1(n6626), .A2(n4410), .B1(n5530), .B2(n5529), .C1(n6628), 
        .C2(n6500), .ZN(n4411) );
  OAI21_X1 U5468 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6626), .A(n6630), 
        .ZN(n4416) );
  AOI22_X1 U5469 ( .A1(n6630), .A2(n4411), .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n4416), .ZN(n4412) );
  INV_X1 U5470 ( .A(n4412), .ZN(U3460) );
  NOR2_X1 U5471 ( .A1(n6630), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4419)
         );
  INV_X1 U5472 ( .A(n4502), .ZN(n4414) );
  OAI22_X1 U5473 ( .A1(n5252), .A2(n4414), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n4413), .ZN(n6497) );
  NOR2_X1 U5474 ( .A1(n6537), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4415)
         );
  AOI211_X1 U5475 ( .C1(n6497), .C2(n5972), .A(n4416), .B(n4415), .ZN(n4418)
         );
  NAND3_X1 U5476 ( .A1(n6498), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n5972), .ZN(n4417) );
  OAI21_X1 U5477 ( .B1(n4419), .B2(n4418), .A(n4417), .ZN(U3461) );
  OAI21_X1 U5478 ( .B1(n5486), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n3103), 
        .ZN(n5258) );
  INV_X1 U5479 ( .A(n4420), .ZN(n4424) );
  INV_X1 U5480 ( .A(n4421), .ZN(n4423) );
  OAI21_X1 U5481 ( .B1(n4424), .B2(n4423), .A(n4422), .ZN(n5253) );
  OAI222_X1 U5482 ( .A1(n5258), .A2(n6150), .B1(n6159), .B2(n3669), .C1(n5636), 
        .C2(n5253), .ZN(U2859) );
  XNOR2_X1 U5483 ( .A(n4425), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4568)
         );
  INV_X1 U5484 ( .A(n5258), .ZN(n4428) );
  INV_X1 U5485 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6638) );
  NOR2_X1 U5486 ( .A1(n6376), .A2(n6638), .ZN(n4565) );
  INV_X1 U5487 ( .A(n4426), .ZN(n4427) );
  AOI211_X1 U5488 ( .C1(n6342), .C2(n4428), .A(n4565), .B(n4427), .ZN(n4432)
         );
  INV_X1 U5489 ( .A(n4429), .ZN(n4430) );
  OAI21_X1 U5490 ( .B1(n4430), .B2(n5297), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4431) );
  OAI211_X1 U5491 ( .C1(n4568), .C2(n6354), .A(n4432), .B(n4431), .ZN(U3018)
         );
  OR2_X1 U5492 ( .A1(n4434), .A2(n4433), .ZN(n4435) );
  NAND2_X1 U5493 ( .A1(n4435), .A2(n4441), .ZN(n6377) );
  NOR2_X1 U5494 ( .A1(n4437), .A2(n4436), .ZN(n4438) );
  NOR2_X1 U5495 ( .A1(n4470), .A2(n4438), .ZN(n6292) );
  INV_X1 U5496 ( .A(n6292), .ZN(n4625) );
  OAI222_X1 U5497 ( .A1(n6377), .A2(n6150), .B1(n4439), .B2(n6159), .C1(n4625), 
        .C2(n5636), .ZN(U2857) );
  XOR2_X1 U5498 ( .A(n4440), .B(n4470), .Z(n6284) );
  INV_X1 U5499 ( .A(n6284), .ZN(n4615) );
  XNOR2_X1 U5500 ( .A(n4442), .B(n4441), .ZN(n6362) );
  INV_X1 U5501 ( .A(n6362), .ZN(n4443) );
  AOI22_X1 U5502 ( .A1(n6155), .A2(n4443), .B1(n5620), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4444) );
  OAI21_X1 U5503 ( .B1(n4615), .B2(n5601), .A(n4444), .ZN(U2856) );
  INV_X1 U5504 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6213) );
  OR2_X1 U5505 ( .A1(n4611), .A2(n4445), .ZN(n4446) );
  NAND2_X1 U5506 ( .A1(n6256), .A2(n4446), .ZN(n4448) );
  NAND2_X1 U5507 ( .A1(n6981), .A2(n4586), .ZN(n4468) );
  NAND2_X1 U5508 ( .A1(n6910), .A2(n4530), .ZN(n6645) );
  AOI22_X1 U5509 ( .A1(DATAO_REG_25__SCAN_IN), .A2(n6980), .B1(n6194), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n4449) );
  OAI21_X1 U5510 ( .B1(n6213), .B2(n4468), .A(n4449), .ZN(U2898) );
  INV_X1 U5511 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6900) );
  AOI22_X1 U5512 ( .A1(DATAO_REG_29__SCAN_IN), .A2(n6980), .B1(n6194), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n4450) );
  OAI21_X1 U5513 ( .B1(n6900), .B2(n4468), .A(n4450), .ZN(U2894) );
  INV_X1 U5514 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6221) );
  AOI22_X1 U5515 ( .A1(DATAO_REG_28__SCAN_IN), .A2(n6980), .B1(n6194), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n4451) );
  OAI21_X1 U5516 ( .B1(n6221), .B2(n4468), .A(n4451), .ZN(U2895) );
  INV_X1 U5517 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4453) );
  AOI22_X1 U5518 ( .A1(DATAO_REG_21__SCAN_IN), .A2(n6980), .B1(
        UWORD_REG_5__SCAN_IN), .B2(n6194), .ZN(n4452) );
  OAI21_X1 U5519 ( .B1(n4453), .B2(n4468), .A(n4452), .ZN(U2902) );
  INV_X1 U5520 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4455) );
  AOI22_X1 U5521 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n6194), .B1(n6980), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4454) );
  OAI21_X1 U5522 ( .B1(n4455), .B2(n4468), .A(n4454), .ZN(U2904) );
  INV_X1 U5523 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6225) );
  AOI22_X1 U5524 ( .A1(n6194), .A2(UWORD_REG_14__SCAN_IN), .B1(n6980), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4456) );
  OAI21_X1 U5525 ( .B1(n6225), .B2(n4468), .A(n4456), .ZN(U2893) );
  INV_X1 U5526 ( .A(EAX_REG_24__SCAN_IN), .ZN(n6210) );
  AOI22_X1 U5527 ( .A1(n6194), .A2(UWORD_REG_8__SCAN_IN), .B1(n6980), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4457) );
  OAI21_X1 U5528 ( .B1(n6210), .B2(n4468), .A(n4457), .ZN(U2899) );
  AOI22_X1 U5529 ( .A1(n6194), .A2(UWORD_REG_0__SCAN_IN), .B1(n6980), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4458) );
  OAI21_X1 U5530 ( .B1(n4024), .B2(n4468), .A(n4458), .ZN(U2907) );
  INV_X1 U5531 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6803) );
  AOI22_X1 U5532 ( .A1(n6194), .A2(UWORD_REG_1__SCAN_IN), .B1(n6980), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4459) );
  OAI21_X1 U5533 ( .B1(n6803), .B2(n4468), .A(n4459), .ZN(U2906) );
  INV_X1 U5534 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4461) );
  AOI22_X1 U5535 ( .A1(n6194), .A2(UWORD_REG_2__SCAN_IN), .B1(n6980), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4460) );
  OAI21_X1 U5536 ( .B1(n4461), .B2(n4468), .A(n4460), .ZN(U2905) );
  INV_X1 U5537 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4463) );
  AOI22_X1 U5538 ( .A1(n6194), .A2(UWORD_REG_4__SCAN_IN), .B1(n6980), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4462) );
  OAI21_X1 U5539 ( .B1(n4463), .B2(n4468), .A(n4462), .ZN(U2903) );
  INV_X1 U5540 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6763) );
  AOI22_X1 U5541 ( .A1(n6194), .A2(UWORD_REG_6__SCAN_IN), .B1(n6980), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4464) );
  OAI21_X1 U5542 ( .B1(n6763), .B2(n4468), .A(n4464), .ZN(U2901) );
  INV_X1 U5543 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6806) );
  AOI22_X1 U5544 ( .A1(n6194), .A2(UWORD_REG_7__SCAN_IN), .B1(n6980), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4465) );
  OAI21_X1 U5545 ( .B1(n6806), .B2(n4468), .A(n4465), .ZN(U2900) );
  INV_X1 U5546 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6792) );
  AOI22_X1 U5547 ( .A1(n6194), .A2(UWORD_REG_10__SCAN_IN), .B1(n6980), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4466) );
  OAI21_X1 U5548 ( .B1(n6792), .B2(n4468), .A(n4466), .ZN(U2897) );
  INV_X1 U5549 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6218) );
  AOI22_X1 U5550 ( .A1(n6194), .A2(UWORD_REG_11__SCAN_IN), .B1(n6980), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4467) );
  OAI21_X1 U5551 ( .B1(n6218), .B2(n4468), .A(n4467), .ZN(U2896) );
  INV_X1 U5552 ( .A(n4617), .ZN(n4472) );
  AOI21_X1 U5553 ( .B1(n4470), .B2(n4440), .A(n4469), .ZN(n4471) );
  NOR2_X1 U5554 ( .A1(n4472), .A2(n4471), .ZN(n5173) );
  INV_X1 U5555 ( .A(n5173), .ZN(n6098) );
  OR2_X1 U5556 ( .A1(n4474), .A2(n4473), .ZN(n4475) );
  NAND2_X1 U5557 ( .A1(n4475), .A2(n4619), .ZN(n6356) );
  INV_X1 U5558 ( .A(n6356), .ZN(n4476) );
  AOI22_X1 U5559 ( .A1(n6155), .A2(n4476), .B1(n5620), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4477) );
  OAI21_X1 U5560 ( .B1(n6098), .B2(n5601), .A(n4477), .ZN(U2855) );
  XNOR2_X1 U5561 ( .A(n4479), .B(n4478), .ZN(n5180) );
  INV_X1 U5562 ( .A(n4480), .ZN(n4483) );
  AND2_X1 U5563 ( .A1(n6340), .A2(REIP_REG_1__SCAN_IN), .ZN(n5175) );
  INV_X1 U5564 ( .A(n5175), .ZN(n4482) );
  NAND2_X1 U5565 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6328), .ZN(n4481)
         );
  OAI211_X1 U5566 ( .C1(n6378), .C2(n4483), .A(n4482), .B(n4481), .ZN(n4484)
         );
  INV_X1 U5567 ( .A(n4484), .ZN(n4488) );
  NAND3_X1 U5568 ( .A1(n6331), .A2(n4486), .A3(n4485), .ZN(n4487) );
  OAI211_X1 U5569 ( .C1(n5180), .C2(n6354), .A(n4488), .B(n4487), .ZN(U3017)
         );
  NAND2_X1 U5570 ( .A1(n6107), .A2(n4502), .ZN(n4500) );
  NAND2_X1 U5571 ( .A1(n5544), .A2(n5540), .ZN(n4508) );
  MUX2_X1 U5572 ( .A(n4490), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n5528), 
        .Z(n4491) );
  NOR2_X1 U5573 ( .A1(n4491), .A2(n4513), .ZN(n4498) );
  AOI21_X1 U5574 ( .B1(n5528), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3122), 
        .ZN(n4492) );
  NOR2_X1 U5575 ( .A1(n3101), .A2(n4492), .ZN(n6627) );
  AND2_X1 U5576 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4494) );
  INV_X1 U5577 ( .A(n4494), .ZN(n4493) );
  MUX2_X1 U5578 ( .A(n4494), .B(n4493), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4495) );
  NAND2_X1 U5579 ( .A1(n6498), .A2(n4495), .ZN(n4496) );
  OAI21_X1 U5580 ( .B1(n6627), .B2(n4505), .A(n4496), .ZN(n4497) );
  AOI21_X1 U5581 ( .B1(n4508), .B2(n4498), .A(n4497), .ZN(n4499) );
  NAND2_X1 U5582 ( .A1(n4500), .A2(n4499), .ZN(n6625) );
  MUX2_X1 U5583 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6625), .S(n6499), 
        .Z(n6511) );
  OR2_X1 U5584 ( .A1(n6499), .A2(n5537), .ZN(n4512) );
  NAND2_X1 U5585 ( .A1(n6116), .A2(n4502), .ZN(n4510) );
  XNOR2_X1 U5586 ( .A(n5528), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4507)
         );
  XNOR2_X1 U5587 ( .A(n5537), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4503)
         );
  NAND2_X1 U5588 ( .A1(n6498), .A2(n4503), .ZN(n4504) );
  OAI21_X1 U5589 ( .B1(n4507), .B2(n4505), .A(n4504), .ZN(n4506) );
  AOI21_X1 U5590 ( .B1(n4508), .B2(n4507), .A(n4506), .ZN(n4509) );
  NAND2_X1 U5591 ( .A1(n4510), .A2(n4509), .ZN(n5534) );
  NAND2_X1 U5592 ( .A1(n6499), .A2(n5534), .ZN(n4511) );
  NAND2_X1 U5593 ( .A1(n4512), .A2(n4511), .ZN(n6506) );
  NAND3_X1 U5594 ( .A1(n6511), .A2(n6537), .A3(n6506), .ZN(n4515) );
  NOR2_X1 U5595 ( .A1(FLUSH_REG_SCAN_IN), .A2(n6537), .ZN(n4520) );
  NAND2_X1 U5596 ( .A1(n4520), .A2(n4513), .ZN(n4514) );
  NAND2_X1 U5597 ( .A1(n4515), .A2(n4514), .ZN(n6512) );
  INV_X1 U5598 ( .A(n4407), .ZN(n4523) );
  INV_X1 U5599 ( .A(n4722), .ZN(n4516) );
  NOR2_X1 U5600 ( .A1(n4517), .A2(n4516), .ZN(n4518) );
  XNOR2_X1 U5601 ( .A(n4518), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6096)
         );
  OAI22_X1 U5602 ( .A1(n6096), .A2(n3655), .B1(n5974), .B2(n6499), .ZN(n4519)
         );
  NAND2_X1 U5603 ( .A1(n4519), .A2(n6537), .ZN(n4522) );
  NAND2_X1 U5604 ( .A1(n4520), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4521) );
  NAND2_X1 U5605 ( .A1(n4522), .A2(n4521), .ZN(n6520) );
  AOI21_X1 U5606 ( .B1(n6512), .B2(n4523), .A(n6520), .ZN(n6524) );
  INV_X1 U5607 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6515) );
  AND2_X1 U5608 ( .A1(n6524), .A2(n6515), .ZN(n4525) );
  OAI21_X1 U5609 ( .B1(n4525), .B2(n4524), .A(n4764), .ZN(n6386) );
  INV_X1 U5610 ( .A(n6386), .ZN(n4537) );
  AOI21_X1 U5611 ( .B1(n4717), .B2(n6735), .A(n6392), .ZN(n4527) );
  NAND2_X1 U5612 ( .A1(n4797), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4863) );
  INV_X1 U5613 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n5105) );
  NAND2_X1 U5614 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5105), .ZN(n5804) );
  AOI22_X1 U5615 ( .A1(n4527), .A2(n4863), .B1(n4660), .B2(n5804), .ZN(n4529)
         );
  NAND2_X1 U5616 ( .A1(n4537), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4528) );
  OAI21_X1 U5617 ( .B1(n4537), .B2(n4529), .A(n4528), .ZN(U3464) );
  AOI222_X1 U5618 ( .A1(n6524), .A2(n4530), .B1(n4867), .B2(n5804), .C1(n5018), 
        .C2(n6395), .ZN(n4532) );
  NAND2_X1 U5619 ( .A1(n4537), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4531) );
  OAI21_X1 U5620 ( .B1(n4537), .B2(n4532), .A(n4531), .ZN(U3465) );
  XNOR2_X1 U5621 ( .A(n4875), .B(n4863), .ZN(n4534) );
  AOI22_X1 U5622 ( .A1(n4534), .A2(n6395), .B1(n5804), .B2(n6116), .ZN(n4536)
         );
  NAND2_X1 U5623 ( .A1(n4537), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4535) );
  OAI21_X1 U5624 ( .B1(n4537), .B2(n4536), .A(n4535), .ZN(U3463) );
  NAND2_X1 U5625 ( .A1(n4875), .A2(n4538), .ZN(n4798) );
  NAND2_X1 U5626 ( .A1(n4797), .A2(n3838), .ZN(n4874) );
  NAND2_X1 U5627 ( .A1(n3099), .A2(DATAI_27_), .ZN(n6479) );
  NAND2_X1 U5628 ( .A1(n3099), .A2(DATAI_19_), .ZN(n6417) );
  INV_X1 U5629 ( .A(n6417), .ZN(n6474) );
  NAND2_X1 U5630 ( .A1(n4797), .A2(n5018), .ZN(n4721) );
  NOR2_X2 U5631 ( .A1(n4798), .A2(n4721), .ZN(n4996) );
  INV_X1 U5632 ( .A(n4539), .ZN(n6621) );
  NAND2_X1 U5633 ( .A1(n4599), .A2(n4541), .ZN(n5135) );
  AND2_X1 U5634 ( .A1(n6107), .A2(n4867), .ZN(n4845) );
  NAND2_X1 U5635 ( .A1(n6116), .A2(n4660), .ZN(n4925) );
  INV_X1 U5636 ( .A(n4925), .ZN(n4543) );
  INV_X1 U5637 ( .A(n4654), .ZN(n4542) );
  AOI21_X1 U5638 ( .B1(n4845), .B2(n4543), .A(n4542), .ZN(n4548) );
  INV_X1 U5639 ( .A(n4548), .ZN(n4545) );
  AOI22_X1 U5640 ( .A1(n4545), .A2(n6395), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4544), .ZN(n4653) );
  INV_X1 U5641 ( .A(DATAI_3_), .ZN(n6231) );
  NOR2_X1 U5642 ( .A1(n6231), .A2(n4764), .ZN(n6476) );
  INV_X1 U5643 ( .A(n6476), .ZN(n5134) );
  OAI22_X1 U5644 ( .A1(n5135), .A2(n4654), .B1(n4653), .B2(n5134), .ZN(n4546)
         );
  AOI21_X1 U5645 ( .B1(n6474), .B2(n4996), .A(n4546), .ZN(n4553) );
  OAI21_X1 U5646 ( .B1(n4798), .B2(n4717), .A(n3099), .ZN(n4547) );
  AND2_X1 U5647 ( .A1(n6395), .A2(n6735), .ZN(n4971) );
  INV_X1 U5648 ( .A(n4971), .ZN(n5806) );
  NAND2_X1 U5649 ( .A1(n4547), .A2(n5806), .ZN(n4549) );
  NAND2_X1 U5650 ( .A1(n4549), .A2(n4548), .ZN(n4551) );
  AOI21_X1 U5651 ( .B1(n6392), .B2(n4917), .A(n5012), .ZN(n4550) );
  NAND2_X1 U5652 ( .A1(n4551), .A2(n4550), .ZN(n4656) );
  NAND2_X1 U5653 ( .A1(n4656), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4552)
         );
  OAI211_X1 U5654 ( .C1(n4952), .C2(n6479), .A(n4553), .B(n4552), .ZN(U3143)
         );
  NAND2_X1 U5655 ( .A1(n3099), .A2(DATAI_31_), .ZN(n6496) );
  NAND2_X1 U5656 ( .A1(n3099), .A2(DATAI_23_), .ZN(n6439) );
  INV_X1 U5657 ( .A(n6439), .ZN(n6487) );
  NAND2_X1 U5658 ( .A1(n4599), .A2(n4554), .ZN(n5130) );
  INV_X1 U5659 ( .A(DATAI_7_), .ZN(n6237) );
  NOR2_X1 U5660 ( .A1(n6237), .A2(n4764), .ZN(n6491) );
  INV_X1 U5661 ( .A(n6491), .ZN(n5129) );
  OAI22_X1 U5662 ( .A1(n5130), .A2(n4654), .B1(n4653), .B2(n5129), .ZN(n4555)
         );
  AOI21_X1 U5663 ( .B1(n6487), .B2(n4996), .A(n4555), .ZN(n4557) );
  NAND2_X1 U5664 ( .A1(n4656), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4556)
         );
  OAI211_X1 U5665 ( .C1(n4952), .C2(n6496), .A(n4557), .B(n4556), .ZN(U3147)
         );
  NAND2_X1 U5666 ( .A1(n3099), .A2(DATAI_28_), .ZN(n6485) );
  NAND2_X1 U5667 ( .A1(n3099), .A2(DATAI_20_), .ZN(n6421) );
  INV_X1 U5668 ( .A(n6421), .ZN(n6480) );
  NAND2_X1 U5669 ( .A1(n4599), .A2(n4558), .ZN(n5145) );
  INV_X1 U5670 ( .A(DATAI_4_), .ZN(n6805) );
  NOR2_X1 U5671 ( .A1(n6805), .A2(n4764), .ZN(n6482) );
  INV_X1 U5672 ( .A(n6482), .ZN(n5144) );
  OAI22_X1 U5673 ( .A1(n5145), .A2(n4654), .B1(n4653), .B2(n5144), .ZN(n4559)
         );
  AOI21_X1 U5674 ( .B1(n6480), .B2(n4996), .A(n4559), .ZN(n4561) );
  NAND2_X1 U5675 ( .A1(n4656), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4560)
         );
  OAI211_X1 U5676 ( .C1(n4952), .C2(n6485), .A(n4561), .B(n4560), .ZN(U3144)
         );
  INV_X1 U5677 ( .A(n5253), .ZN(n4566) );
  INV_X1 U5678 ( .A(n6288), .ZN(n5699) );
  INV_X1 U5679 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4562) );
  AOI21_X1 U5680 ( .B1(n5699), .B2(n4563), .A(n4562), .ZN(n4564) );
  AOI211_X1 U5681 ( .C1(n4566), .C2(n3099), .A(n4565), .B(n4564), .ZN(n4567)
         );
  OAI21_X1 U5682 ( .B1(n4568), .B2(n5984), .A(n4567), .ZN(U2986) );
  INV_X1 U5683 ( .A(n4875), .ZN(n4569) );
  NAND2_X1 U5684 ( .A1(n4569), .A2(n5800), .ZN(n4861) );
  OR2_X1 U5685 ( .A1(n4861), .A2(n4863), .ZN(n4570) );
  NAND2_X1 U5686 ( .A1(n4570), .A2(n6395), .ZN(n4579) );
  NOR2_X1 U5687 ( .A1(n6116), .A2(n6136), .ZN(n4865) );
  AND2_X1 U5688 ( .A1(n4865), .A2(n6107), .ZN(n5067) );
  NAND2_X1 U5689 ( .A1(n5067), .A2(n4867), .ZN(n4572) );
  INV_X1 U5690 ( .A(n4866), .ZN(n4571) );
  NAND2_X1 U5691 ( .A1(n4571), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6473) );
  NAND2_X1 U5692 ( .A1(n4572), .A2(n6473), .ZN(n4578) );
  INV_X1 U5693 ( .A(n4578), .ZN(n4573) );
  OR2_X1 U5694 ( .A1(n4579), .A2(n4573), .ZN(n4576) );
  NAND3_X1 U5695 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6505), .ZN(n5068) );
  INV_X1 U5696 ( .A(n5068), .ZN(n4574) );
  NAND2_X1 U5697 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4574), .ZN(n4575) );
  NAND2_X1 U5698 ( .A1(n4576), .A2(n4575), .ZN(n6490) );
  INV_X1 U5699 ( .A(n6490), .ZN(n4604) );
  INV_X1 U5700 ( .A(DATAI_1_), .ZN(n6751) );
  NOR2_X1 U5701 ( .A1(n6751), .A2(n4764), .ZN(n6448) );
  AOI21_X1 U5702 ( .B1(n5068), .B2(n6392), .A(n5012), .ZN(n4577) );
  OAI21_X1 U5703 ( .B1(n4579), .B2(n4578), .A(n4577), .ZN(n6492) );
  NAND2_X1 U5704 ( .A1(n6492), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4585)
         );
  INV_X1 U5705 ( .A(n6495), .ZN(n4601) );
  NAND2_X1 U5706 ( .A1(n3099), .A2(DATAI_25_), .ZN(n6451) );
  INV_X1 U5707 ( .A(n6451), .ZN(n6406) );
  NAND2_X1 U5708 ( .A1(n4599), .A2(n4580), .ZN(n5140) );
  NAND2_X1 U5709 ( .A1(n3099), .A2(DATAI_17_), .ZN(n6409) );
  INV_X1 U5710 ( .A(n4861), .ZN(n4582) );
  INV_X1 U5711 ( .A(n4721), .ZN(n4581) );
  OAI22_X1 U5712 ( .A1(n5140), .A2(n6473), .B1(n6409), .B2(n4835), .ZN(n4583)
         );
  AOI21_X1 U5713 ( .B1(n4601), .B2(n6406), .A(n4583), .ZN(n4584) );
  OAI211_X1 U5714 ( .C1(n4604), .C2(n5139), .A(n4585), .B(n4584), .ZN(U3109)
         );
  INV_X1 U5715 ( .A(DATAI_0_), .ZN(n6227) );
  NOR2_X1 U5716 ( .A1(n6227), .A2(n4764), .ZN(n6442) );
  INV_X1 U5717 ( .A(n6442), .ZN(n5124) );
  NAND2_X1 U5718 ( .A1(n6492), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4589)
         );
  NAND2_X1 U5719 ( .A1(n3099), .A2(DATAI_24_), .ZN(n6445) );
  INV_X1 U5720 ( .A(n6445), .ZN(n6402) );
  NAND2_X1 U5721 ( .A1(n4599), .A2(n4586), .ZN(n5125) );
  NAND2_X1 U5722 ( .A1(n3099), .A2(DATAI_16_), .ZN(n6405) );
  OAI22_X1 U5723 ( .A1(n5125), .A2(n6473), .B1(n6405), .B2(n4835), .ZN(n4587)
         );
  AOI21_X1 U5724 ( .B1(n4601), .B2(n6402), .A(n4587), .ZN(n4588) );
  OAI211_X1 U5725 ( .C1(n4604), .C2(n5124), .A(n4589), .B(n4588), .ZN(U3108)
         );
  INV_X1 U5726 ( .A(DATAI_2_), .ZN(n6888) );
  NOR2_X1 U5727 ( .A1(n6888), .A2(n4764), .ZN(n6454) );
  INV_X1 U5728 ( .A(n6454), .ZN(n5123) );
  NAND2_X1 U5729 ( .A1(n6492), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4593)
         );
  NAND2_X1 U5730 ( .A1(n3099), .A2(DATAI_26_), .ZN(n6457) );
  INV_X1 U5731 ( .A(n6457), .ZN(n6410) );
  NAND2_X1 U5732 ( .A1(n4599), .A2(n4590), .ZN(n5118) );
  NAND2_X1 U5733 ( .A1(n3099), .A2(DATAI_18_), .ZN(n6413) );
  OAI22_X1 U5734 ( .A1(n5118), .A2(n6473), .B1(n6413), .B2(n4835), .ZN(n4591)
         );
  AOI21_X1 U5735 ( .B1(n4601), .B2(n6410), .A(n4591), .ZN(n4592) );
  OAI211_X1 U5736 ( .C1(n4604), .C2(n5123), .A(n4593), .B(n4592), .ZN(U3110)
         );
  INV_X1 U5737 ( .A(DATAI_5_), .ZN(n6234) );
  NOR2_X1 U5738 ( .A1(n6234), .A2(n4764), .ZN(n6462) );
  INV_X1 U5739 ( .A(n6462), .ZN(n5150) );
  NAND2_X1 U5740 ( .A1(n6492), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4597)
         );
  NAND2_X1 U5741 ( .A1(n3099), .A2(DATAI_29_), .ZN(n6465) );
  INV_X1 U5742 ( .A(n6465), .ZN(n6422) );
  NAND2_X1 U5743 ( .A1(n4599), .A2(n4594), .ZN(n5153) );
  NAND2_X1 U5744 ( .A1(n3099), .A2(DATAI_21_), .ZN(n6425) );
  OAI22_X1 U5745 ( .A1(n5153), .A2(n6473), .B1(n6425), .B2(n4835), .ZN(n4595)
         );
  AOI21_X1 U5746 ( .B1(n4601), .B2(n6422), .A(n4595), .ZN(n4596) );
  OAI211_X1 U5747 ( .C1(n4604), .C2(n5150), .A(n4597), .B(n4596), .ZN(U3113)
         );
  INV_X1 U5748 ( .A(DATAI_6_), .ZN(n6728) );
  NOR2_X1 U5749 ( .A1(n6728), .A2(n4764), .ZN(n6426) );
  NAND2_X1 U5750 ( .A1(n6492), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4603)
         );
  AND2_X1 U5751 ( .A1(n3099), .A2(DATAI_30_), .ZN(n6428) );
  NAND2_X1 U5752 ( .A1(n4599), .A2(n4598), .ZN(n5111) );
  NAND2_X1 U5753 ( .A1(n3099), .A2(DATAI_22_), .ZN(n6431) );
  OAI22_X1 U5754 ( .A1(n5111), .A2(n6473), .B1(n6431), .B2(n4835), .ZN(n4600)
         );
  AOI21_X1 U5755 ( .B1(n4601), .B2(n6428), .A(n4600), .ZN(n4602) );
  OAI211_X1 U5756 ( .C1(n4604), .C2(n5110), .A(n4603), .B(n4602), .ZN(U3114)
         );
  NAND2_X1 U5757 ( .A1(n6525), .A2(n4606), .ZN(n4608) );
  OAI22_X1 U5758 ( .A1(n3655), .A2(n4608), .B1(n3563), .B2(n4607), .ZN(n4609)
         );
  INV_X1 U5759 ( .A(n4609), .ZN(n4610) );
  AND2_X1 U5760 ( .A1(n5377), .A2(n4612), .ZN(n4613) );
  INV_X1 U5761 ( .A(n4613), .ZN(n4614) );
  NAND2_X1 U5762 ( .A1(n5640), .A2(n4614), .ZN(n5642) );
  INV_X1 U5763 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6191) );
  OAI222_X1 U5764 ( .A1(n4615), .A2(n5639), .B1(n5642), .B2(n6231), .C1(n5640), 
        .C2(n6191), .ZN(U2888) );
  INV_X1 U5765 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6197) );
  OAI222_X1 U5766 ( .A1(n5253), .A2(n5639), .B1(n5642), .B2(n6227), .C1(n5640), 
        .C2(n6197), .ZN(U2891) );
  INV_X1 U5767 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6189) );
  OAI222_X1 U5768 ( .A1(n6098), .A2(n5639), .B1(n5642), .B2(n6805), .C1(n5640), 
        .C2(n6189), .ZN(U2887) );
  INV_X1 U5769 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6193) );
  OAI222_X1 U5770 ( .A1(n6144), .A2(n5639), .B1(n5642), .B2(n6751), .C1(n5640), 
        .C2(n6193), .ZN(U2890) );
  XOR2_X1 U5771 ( .A(n4617), .B(n4616), .Z(n6276) );
  INV_X1 U5772 ( .A(n6276), .ZN(n4629) );
  AOI21_X1 U5773 ( .B1(n4620), .B2(n4619), .A(n4618), .ZN(n6341) );
  AOI22_X1 U5774 ( .A1(n6155), .A2(n6341), .B1(n5620), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n4621) );
  OAI21_X1 U5775 ( .B1(n4629), .B2(n5601), .A(n4621), .ZN(U2854) );
  INV_X1 U5776 ( .A(n4622), .ZN(n6334) );
  AOI22_X1 U5777 ( .A1(n6155), .A2(n6334), .B1(n5620), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4623) );
  OAI21_X1 U5778 ( .B1(n5278), .B2(n5601), .A(n4623), .ZN(U2853) );
  INV_X1 U5779 ( .A(n5642), .ZN(n5342) );
  AOI22_X1 U5780 ( .A1(n5342), .A2(DATAI_2_), .B1(EAX_REG_2__SCAN_IN), .B2(
        n6170), .ZN(n4624) );
  OAI21_X1 U5781 ( .B1(n4625), .B2(n5639), .A(n4624), .ZN(U2889) );
  INV_X1 U5782 ( .A(n4996), .ZN(n5001) );
  OAI22_X1 U5783 ( .A1(n5118), .A2(n4654), .B1(n6413), .B2(n5001), .ZN(n4626)
         );
  AOI21_X1 U5784 ( .B1(n6410), .B2(n4948), .A(n4626), .ZN(n4628) );
  NAND2_X1 U5785 ( .A1(n4656), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4627)
         );
  OAI211_X1 U5786 ( .C1(n5123), .C2(n4653), .A(n4628), .B(n4627), .ZN(U3142)
         );
  OAI222_X1 U5787 ( .A1(n5639), .A2(n4629), .B1(n5642), .B2(n6234), .C1(n5640), 
        .C2(n3872), .ZN(U2886) );
  INV_X1 U5788 ( .A(n4538), .ZN(n4630) );
  INV_X1 U5789 ( .A(n4874), .ZN(n4631) );
  OR2_X1 U5790 ( .A1(n6107), .A2(n4925), .ZN(n6394) );
  INV_X1 U5791 ( .A(n6394), .ZN(n4633) );
  INV_X1 U5792 ( .A(n4632), .ZN(n6467) );
  AOI21_X1 U5793 ( .B1(n4633), .B2(n4867), .A(n6467), .ZN(n4638) );
  INV_X1 U5794 ( .A(n4638), .ZN(n4636) );
  INV_X1 U5795 ( .A(n4863), .ZN(n4634) );
  NAND2_X1 U5796 ( .A1(n4718), .A2(n4634), .ZN(n5801) );
  NAND2_X1 U5797 ( .A1(n6395), .A2(n5801), .ZN(n4637) );
  AOI21_X1 U5798 ( .B1(n6392), .B2(n6388), .A(n5012), .ZN(n4635) );
  OAI21_X1 U5799 ( .B1(n4636), .B2(n4637), .A(n4635), .ZN(n6469) );
  OAI22_X1 U5800 ( .A1(n4638), .A2(n4637), .B1(n6647), .B2(n6388), .ZN(n6468)
         );
  AOI22_X1 U5801 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6469), .B1(n6476), 
        .B2(n6468), .ZN(n4641) );
  INV_X1 U5802 ( .A(n4718), .ZN(n4639) );
  NOR2_X2 U5803 ( .A1(n4639), .A2(n4721), .ZN(n6466) );
  AOI22_X1 U5804 ( .A1(n6475), .A2(n6467), .B1(n6474), .B2(n6466), .ZN(n4640)
         );
  OAI211_X1 U5805 ( .C1(n6479), .C2(n6472), .A(n4641), .B(n4640), .ZN(U3079)
         );
  INV_X1 U5806 ( .A(n6428), .ZN(n5116) );
  AOI22_X1 U5807 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6469), .B1(n6426), 
        .B2(n6468), .ZN(n4643) );
  INV_X1 U5808 ( .A(n6431), .ZN(n5113) );
  AOI22_X1 U5809 ( .A1(n6427), .A2(n6467), .B1(n5113), .B2(n6466), .ZN(n4642)
         );
  OAI211_X1 U5810 ( .C1(n5116), .C2(n6472), .A(n4643), .B(n4642), .ZN(U3082)
         );
  INV_X1 U5811 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6866) );
  OAI222_X1 U5812 ( .A1(n5278), .A2(n5639), .B1(n5642), .B2(n6728), .C1(n5640), 
        .C2(n6866), .ZN(U2885) );
  OAI22_X1 U5813 ( .A1(n5111), .A2(n4654), .B1(n4653), .B2(n5110), .ZN(n4644)
         );
  AOI21_X1 U5814 ( .B1(n5113), .B2(n4996), .A(n4644), .ZN(n4646) );
  NAND2_X1 U5815 ( .A1(n4656), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4645)
         );
  OAI211_X1 U5816 ( .C1(n4952), .C2(n5116), .A(n4646), .B(n4645), .ZN(U3146)
         );
  INV_X1 U5817 ( .A(n6409), .ZN(n6446) );
  OAI22_X1 U5818 ( .A1(n5140), .A2(n4654), .B1(n4653), .B2(n5139), .ZN(n4647)
         );
  AOI21_X1 U5819 ( .B1(n6446), .B2(n4996), .A(n4647), .ZN(n4649) );
  NAND2_X1 U5820 ( .A1(n4656), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4648)
         );
  OAI211_X1 U5821 ( .C1(n4952), .C2(n6451), .A(n4649), .B(n4648), .ZN(U3141)
         );
  INV_X1 U5822 ( .A(n6425), .ZN(n6460) );
  OAI22_X1 U5823 ( .A1(n5153), .A2(n4654), .B1(n4653), .B2(n5150), .ZN(n4650)
         );
  AOI21_X1 U5824 ( .B1(n6460), .B2(n4996), .A(n4650), .ZN(n4652) );
  NAND2_X1 U5825 ( .A1(n4656), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4651)
         );
  OAI211_X1 U5826 ( .C1(n4952), .C2(n6465), .A(n4652), .B(n4651), .ZN(U3145)
         );
  INV_X1 U5827 ( .A(n6405), .ZN(n6440) );
  OAI22_X1 U5828 ( .A1(n5125), .A2(n4654), .B1(n4653), .B2(n5124), .ZN(n4655)
         );
  AOI21_X1 U5829 ( .B1(n6440), .B2(n4996), .A(n4655), .ZN(n4658) );
  NAND2_X1 U5830 ( .A1(n4656), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4657)
         );
  OAI211_X1 U5831 ( .C1(n4952), .C2(n6445), .A(n4658), .B(n4657), .ZN(U3140)
         );
  INV_X1 U5832 ( .A(n4665), .ZN(n4659) );
  OAI21_X1 U5833 ( .B1(n4659), .B2(n6735), .A(n6395), .ZN(n4664) );
  OR2_X1 U5834 ( .A1(n6116), .A2(n4660), .ZN(n4685) );
  OR2_X1 U5835 ( .A1(n4685), .A2(n6107), .ZN(n4970) );
  INV_X1 U5836 ( .A(n4970), .ZN(n4976) );
  NAND3_X1 U5837 ( .A1(n6734), .A2(n6505), .A3(n4719), .ZN(n4968) );
  NOR2_X1 U5838 ( .A1(n6917), .A2(n4968), .ZN(n4682) );
  AOI21_X1 U5839 ( .B1(n4976), .B2(n4867), .A(n4682), .ZN(n4663) );
  INV_X1 U5840 ( .A(n4663), .ZN(n4662) );
  AOI21_X1 U5841 ( .B1(n6392), .B2(n4968), .A(n5012), .ZN(n4661) );
  OAI21_X1 U5842 ( .B1(n4664), .B2(n4662), .A(n4661), .ZN(n4681) );
  OAI22_X1 U5843 ( .A1(n4664), .A2(n4663), .B1(n6647), .B2(n4968), .ZN(n4680)
         );
  AOI22_X1 U5844 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4681), .B1(n6448), 
        .B2(n4680), .ZN(n4667) );
  NAND2_X1 U5845 ( .A1(n4665), .A2(n5018), .ZN(n5158) );
  AOI22_X1 U5846 ( .A1(n6447), .A2(n4682), .B1(n6446), .B2(n5120), .ZN(n4666)
         );
  OAI211_X1 U5847 ( .C1(n6451), .C2(n4999), .A(n4667), .B(n4666), .ZN(U3029)
         );
  AOI22_X1 U5848 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4681), .B1(n6454), 
        .B2(n4680), .ZN(n4669) );
  INV_X1 U5849 ( .A(n6413), .ZN(n6452) );
  AOI22_X1 U5850 ( .A1(n6453), .A2(n4682), .B1(n6452), .B2(n5120), .ZN(n4668)
         );
  OAI211_X1 U5851 ( .C1(n6457), .C2(n4999), .A(n4669), .B(n4668), .ZN(U3030)
         );
  AOI22_X1 U5852 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4681), .B1(n6442), 
        .B2(n4680), .ZN(n4671) );
  AOI22_X1 U5853 ( .A1(n6441), .A2(n4682), .B1(n6440), .B2(n5120), .ZN(n4670)
         );
  OAI211_X1 U5854 ( .C1(n6445), .C2(n4999), .A(n4671), .B(n4670), .ZN(U3028)
         );
  AOI22_X1 U5855 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4681), .B1(n6482), 
        .B2(n4680), .ZN(n4673) );
  AOI22_X1 U5856 ( .A1(n6481), .A2(n4682), .B1(n6480), .B2(n5120), .ZN(n4672)
         );
  OAI211_X1 U5857 ( .C1(n6485), .C2(n4999), .A(n4673), .B(n4672), .ZN(U3032)
         );
  AOI22_X1 U5858 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4681), .B1(n6426), 
        .B2(n4680), .ZN(n4675) );
  AOI22_X1 U5859 ( .A1(n6427), .A2(n4682), .B1(n5113), .B2(n5120), .ZN(n4674)
         );
  OAI211_X1 U5860 ( .C1(n5116), .C2(n4999), .A(n4675), .B(n4674), .ZN(U3034)
         );
  AOI22_X1 U5861 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4681), .B1(n6462), 
        .B2(n4680), .ZN(n4677) );
  AOI22_X1 U5862 ( .A1(n6461), .A2(n4682), .B1(n6460), .B2(n5120), .ZN(n4676)
         );
  OAI211_X1 U5863 ( .C1(n6465), .C2(n4999), .A(n4677), .B(n4676), .ZN(U3033)
         );
  AOI22_X1 U5864 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4681), .B1(n6476), 
        .B2(n4680), .ZN(n4679) );
  AOI22_X1 U5865 ( .A1(n6475), .A2(n4682), .B1(n6474), .B2(n5120), .ZN(n4678)
         );
  OAI211_X1 U5866 ( .C1(n6479), .C2(n4999), .A(n4679), .B(n4678), .ZN(U3031)
         );
  AOI22_X1 U5867 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4681), .B1(n6491), 
        .B2(n4680), .ZN(n4684) );
  AOI22_X1 U5868 ( .A1(n6489), .A2(n4682), .B1(n6487), .B2(n5120), .ZN(n4683)
         );
  OAI211_X1 U5869 ( .C1(n6496), .C2(n4999), .A(n4684), .B(n4683), .ZN(U3035)
         );
  OAI21_X1 U5870 ( .B1(n4690), .B2(n6735), .A(n6395), .ZN(n4688) );
  INV_X1 U5871 ( .A(n4685), .ZN(n4758) );
  NAND3_X1 U5872 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6505), .A3(n4719), .ZN(n4757) );
  NOR2_X1 U5873 ( .A1(n6917), .A2(n4757), .ZN(n4707) );
  AOI21_X1 U5874 ( .B1(n4845), .B2(n4758), .A(n4707), .ZN(n4689) );
  INV_X1 U5875 ( .A(n4689), .ZN(n4687) );
  AOI21_X1 U5876 ( .B1(n6392), .B2(n4757), .A(n5012), .ZN(n4686) );
  OAI21_X1 U5877 ( .B1(n4688), .B2(n4687), .A(n4686), .ZN(n4706) );
  OAI22_X1 U5878 ( .A1(n4689), .A2(n4688), .B1(n6647), .B2(n4757), .ZN(n4705)
         );
  AOI22_X1 U5879 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4706), .B1(n6491), 
        .B2(n4705), .ZN(n4692) );
  AOI22_X1 U5880 ( .A1(n6489), .A2(n4707), .B1(n5096), .B2(n6487), .ZN(n4691)
         );
  OAI211_X1 U5881 ( .C1(n6496), .C2(n4796), .A(n4692), .B(n4691), .ZN(U3099)
         );
  AOI22_X1 U5882 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4706), .B1(n6476), 
        .B2(n4705), .ZN(n4694) );
  AOI22_X1 U5883 ( .A1(n6475), .A2(n4707), .B1(n5096), .B2(n6474), .ZN(n4693)
         );
  OAI211_X1 U5884 ( .C1(n6479), .C2(n4796), .A(n4694), .B(n4693), .ZN(U3095)
         );
  AOI22_X1 U5885 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4706), .B1(n6454), 
        .B2(n4705), .ZN(n4696) );
  AOI22_X1 U5886 ( .A1(n6453), .A2(n4707), .B1(n5096), .B2(n6452), .ZN(n4695)
         );
  OAI211_X1 U5887 ( .C1(n6457), .C2(n4796), .A(n4696), .B(n4695), .ZN(U3094)
         );
  AOI22_X1 U5888 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4706), .B1(n6482), 
        .B2(n4705), .ZN(n4698) );
  AOI22_X1 U5889 ( .A1(n6481), .A2(n4707), .B1(n5096), .B2(n6480), .ZN(n4697)
         );
  OAI211_X1 U5890 ( .C1(n6485), .C2(n4796), .A(n4698), .B(n4697), .ZN(U3096)
         );
  AOI22_X1 U5891 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4706), .B1(n6462), 
        .B2(n4705), .ZN(n4700) );
  AOI22_X1 U5892 ( .A1(n6461), .A2(n4707), .B1(n5096), .B2(n6460), .ZN(n4699)
         );
  OAI211_X1 U5893 ( .C1(n6465), .C2(n4796), .A(n4700), .B(n4699), .ZN(U3097)
         );
  AOI22_X1 U5894 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4706), .B1(n6426), 
        .B2(n4705), .ZN(n4702) );
  AOI22_X1 U5895 ( .A1(n6427), .A2(n4707), .B1(n5096), .B2(n5113), .ZN(n4701)
         );
  OAI211_X1 U5896 ( .C1(n5116), .C2(n4796), .A(n4702), .B(n4701), .ZN(U3098)
         );
  AOI22_X1 U5897 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4706), .B1(n6442), 
        .B2(n4705), .ZN(n4704) );
  AOI22_X1 U5898 ( .A1(n6441), .A2(n4707), .B1(n5096), .B2(n6440), .ZN(n4703)
         );
  OAI211_X1 U5899 ( .C1(n6445), .C2(n4796), .A(n4704), .B(n4703), .ZN(U3092)
         );
  AOI22_X1 U5900 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4706), .B1(n6448), 
        .B2(n4705), .ZN(n4709) );
  AOI22_X1 U5901 ( .A1(n6447), .A2(n4707), .B1(n5096), .B2(n6446), .ZN(n4708)
         );
  OAI211_X1 U5902 ( .C1(n6451), .C2(n4796), .A(n4709), .B(n4708), .ZN(U3093)
         );
  AND2_X1 U5903 ( .A1(n4711), .A2(n4710), .ZN(n4713) );
  OR2_X1 U5904 ( .A1(n4713), .A2(n4959), .ZN(n6267) );
  AOI21_X1 U5905 ( .B1(n4715), .B2(n4714), .A(n4961), .ZN(n6322) );
  AOI22_X1 U5906 ( .A1(n6155), .A2(n6322), .B1(n5620), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n4716) );
  OAI21_X1 U5907 ( .B1(n6267), .B2(n5636), .A(n4716), .ZN(U2852) );
  NAND2_X1 U5908 ( .A1(n5019), .A2(n3838), .ZN(n5050) );
  NAND2_X1 U5909 ( .A1(n4719), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4850) );
  INV_X1 U5910 ( .A(n4850), .ZN(n4800) );
  NAND2_X1 U5911 ( .A1(n4800), .A2(n6734), .ZN(n5015) );
  OR2_X1 U5912 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5015), .ZN(n4752)
         );
  NOR2_X1 U5913 ( .A1(n4726), .A2(n6647), .ZN(n6398) );
  INV_X1 U5914 ( .A(n4759), .ZN(n4720) );
  NOR2_X1 U5915 ( .A1(n6389), .A2(n4720), .ZN(n4975) );
  OAI21_X1 U5916 ( .B1(n4975), .B2(n6647), .A(n4918), .ZN(n4969) );
  AOI211_X1 U5917 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4752), .A(n6398), .B(
        n4969), .ZN(n4724) );
  AOI21_X1 U5918 ( .B1(n5019), .B2(STATEBS16_REG_SCAN_IN), .A(n6392), .ZN(
        n5008) );
  NAND2_X1 U5919 ( .A1(n6116), .A2(n6136), .ZN(n4725) );
  OR2_X1 U5920 ( .A1(n4725), .A2(n4722), .ZN(n5009) );
  OAI211_X1 U5921 ( .C1(n4971), .C2(n4899), .A(n5008), .B(n5009), .ZN(n4723)
         );
  NAND2_X1 U5922 ( .A1(n4724), .A2(n4723), .ZN(n4750) );
  NAND2_X1 U5923 ( .A1(n4750), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4730) );
  INV_X1 U5924 ( .A(n6485), .ZN(n6418) );
  INV_X1 U5925 ( .A(n4725), .ZN(n4844) );
  NAND2_X1 U5926 ( .A1(n4844), .A2(n6395), .ZN(n4806) );
  AND2_X1 U5927 ( .A1(n4726), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6390) );
  INV_X1 U5928 ( .A(n6390), .ZN(n4926) );
  INV_X1 U5929 ( .A(n4975), .ZN(n4727) );
  OAI22_X1 U5930 ( .A1(n4806), .A2(n6107), .B1(n4926), .B2(n4727), .ZN(n4738)
         );
  INV_X1 U5931 ( .A(n4738), .ZN(n4751) );
  OAI22_X1 U5932 ( .A1(n5145), .A2(n4752), .B1(n4751), .B2(n5144), .ZN(n4728)
         );
  AOI21_X1 U5933 ( .B1(n6418), .B2(n4754), .A(n4728), .ZN(n4729) );
  OAI211_X1 U5934 ( .C1(n5050), .C2(n6421), .A(n4730), .B(n4729), .ZN(U3056)
         );
  NAND2_X1 U5935 ( .A1(n4750), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4733) );
  INV_X1 U5936 ( .A(n6496), .ZN(n6435) );
  OAI22_X1 U5937 ( .A1(n5130), .A2(n4752), .B1(n4751), .B2(n5129), .ZN(n4731)
         );
  AOI21_X1 U5938 ( .B1(n6435), .B2(n4754), .A(n4731), .ZN(n4732) );
  OAI211_X1 U5939 ( .C1(n5050), .C2(n6439), .A(n4733), .B(n4732), .ZN(U3059)
         );
  NAND2_X1 U5940 ( .A1(n4750), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4736) );
  INV_X1 U5941 ( .A(n6479), .ZN(n6414) );
  OAI22_X1 U5942 ( .A1(n5135), .A2(n4752), .B1(n4751), .B2(n5134), .ZN(n4734)
         );
  AOI21_X1 U5943 ( .B1(n6414), .B2(n4754), .A(n4734), .ZN(n4735) );
  OAI211_X1 U5944 ( .C1(n5050), .C2(n6417), .A(n4736), .B(n4735), .ZN(U3055)
         );
  NAND2_X1 U5945 ( .A1(n4750), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4740) );
  OAI22_X1 U5946 ( .A1(n5118), .A2(n4752), .B1(n6457), .B2(n4899), .ZN(n4737)
         );
  AOI21_X1 U5947 ( .B1(n6454), .B2(n4738), .A(n4737), .ZN(n4739) );
  OAI211_X1 U5948 ( .C1(n5050), .C2(n6413), .A(n4740), .B(n4739), .ZN(U3054)
         );
  NAND2_X1 U5949 ( .A1(n4750), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4743) );
  OAI22_X1 U5950 ( .A1(n5111), .A2(n4752), .B1(n4751), .B2(n5110), .ZN(n4741)
         );
  AOI21_X1 U5951 ( .B1(n6428), .B2(n4754), .A(n4741), .ZN(n4742) );
  OAI211_X1 U5952 ( .C1(n5050), .C2(n6431), .A(n4743), .B(n4742), .ZN(U3058)
         );
  NAND2_X1 U5953 ( .A1(n4750), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4746) );
  OAI22_X1 U5954 ( .A1(n5125), .A2(n4752), .B1(n4751), .B2(n5124), .ZN(n4744)
         );
  AOI21_X1 U5955 ( .B1(n6402), .B2(n4754), .A(n4744), .ZN(n4745) );
  OAI211_X1 U5956 ( .C1(n6405), .C2(n5050), .A(n4746), .B(n4745), .ZN(U3052)
         );
  NAND2_X1 U5957 ( .A1(n4750), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4749) );
  OAI22_X1 U5958 ( .A1(n5140), .A2(n4752), .B1(n4751), .B2(n5139), .ZN(n4747)
         );
  AOI21_X1 U5959 ( .B1(n6406), .B2(n4754), .A(n4747), .ZN(n4748) );
  OAI211_X1 U5960 ( .C1(n5050), .C2(n6409), .A(n4749), .B(n4748), .ZN(U3053)
         );
  NAND2_X1 U5961 ( .A1(n4750), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4756) );
  OAI22_X1 U5962 ( .A1(n5153), .A2(n4752), .B1(n4751), .B2(n5150), .ZN(n4753)
         );
  AOI21_X1 U5963 ( .B1(n6422), .B2(n4754), .A(n4753), .ZN(n4755) );
  OAI211_X1 U5964 ( .C1(n5050), .C2(n6425), .A(n4756), .B(n4755), .ZN(U3057)
         );
  NOR2_X1 U5965 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4757), .ZN(n4765)
         );
  INV_X1 U5966 ( .A(n4765), .ZN(n4791) );
  NAND2_X1 U5967 ( .A1(n4758), .A2(n6107), .ZN(n4761) );
  INV_X1 U5968 ( .A(n6398), .ZN(n5107) );
  OR2_X1 U5969 ( .A1(n6389), .A2(n4759), .ZN(n4805) );
  OAI22_X1 U5970 ( .A1(n4761), .A2(n6392), .B1(n5107), .B2(n4805), .ZN(n4781)
         );
  INV_X1 U5971 ( .A(n4781), .ZN(n4790) );
  OAI22_X1 U5972 ( .A1(n5153), .A2(n4791), .B1(n4790), .B2(n5150), .ZN(n4760)
         );
  AOI21_X1 U5973 ( .B1(n6422), .B2(n6466), .A(n4760), .ZN(n4769) );
  INV_X1 U5974 ( .A(n6466), .ZN(n4779) );
  NAND3_X1 U5975 ( .A1(n4779), .A2(n6395), .A3(n4796), .ZN(n4763) );
  INV_X1 U5976 ( .A(n4761), .ZN(n4762) );
  AOI21_X1 U5977 ( .B1(n4763), .B2(n5806), .A(n4762), .ZN(n4767) );
  AOI21_X1 U5978 ( .B1(n4805), .B2(STATE2_REG_2__SCAN_IN), .A(n4764), .ZN(
        n4801) );
  OAI211_X1 U5979 ( .C1(n5105), .C2(n4765), .A(n4926), .B(n4801), .ZN(n4766)
         );
  NAND2_X1 U5980 ( .A1(n4793), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4768) );
  OAI211_X1 U5981 ( .C1(n4796), .C2(n6425), .A(n4769), .B(n4768), .ZN(U3089)
         );
  OAI22_X1 U5982 ( .A1(n5130), .A2(n4791), .B1(n4790), .B2(n5129), .ZN(n4770)
         );
  AOI21_X1 U5983 ( .B1(n6435), .B2(n6466), .A(n4770), .ZN(n4772) );
  NAND2_X1 U5984 ( .A1(n4793), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4771) );
  OAI211_X1 U5985 ( .C1(n4796), .C2(n6439), .A(n4772), .B(n4771), .ZN(U3091)
         );
  OAI22_X1 U5986 ( .A1(n5125), .A2(n4791), .B1(n4790), .B2(n5124), .ZN(n4773)
         );
  AOI21_X1 U5987 ( .B1(n6402), .B2(n6466), .A(n4773), .ZN(n4775) );
  NAND2_X1 U5988 ( .A1(n4793), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4774) );
  OAI211_X1 U5989 ( .C1(n4796), .C2(n6405), .A(n4775), .B(n4774), .ZN(U3084)
         );
  OAI22_X1 U5990 ( .A1(n5140), .A2(n4791), .B1(n4790), .B2(n5139), .ZN(n4776)
         );
  AOI21_X1 U5991 ( .B1(n6406), .B2(n6466), .A(n4776), .ZN(n4778) );
  NAND2_X1 U5992 ( .A1(n4793), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4777) );
  OAI211_X1 U5993 ( .C1(n4796), .C2(n6409), .A(n4778), .B(n4777), .ZN(U3085)
         );
  OAI22_X1 U5994 ( .A1(n5118), .A2(n4791), .B1(n4779), .B2(n6457), .ZN(n4780)
         );
  AOI21_X1 U5995 ( .B1(n6454), .B2(n4781), .A(n4780), .ZN(n4783) );
  NAND2_X1 U5996 ( .A1(n4793), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4782) );
  OAI211_X1 U5997 ( .C1(n4796), .C2(n6413), .A(n4783), .B(n4782), .ZN(U3086)
         );
  OAI22_X1 U5998 ( .A1(n5135), .A2(n4791), .B1(n4790), .B2(n5134), .ZN(n4784)
         );
  AOI21_X1 U5999 ( .B1(n6414), .B2(n6466), .A(n4784), .ZN(n4786) );
  NAND2_X1 U6000 ( .A1(n4793), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4785) );
  OAI211_X1 U6001 ( .C1(n4796), .C2(n6417), .A(n4786), .B(n4785), .ZN(U3087)
         );
  OAI22_X1 U6002 ( .A1(n5145), .A2(n4791), .B1(n4790), .B2(n5144), .ZN(n4787)
         );
  AOI21_X1 U6003 ( .B1(n6418), .B2(n6466), .A(n4787), .ZN(n4789) );
  NAND2_X1 U6004 ( .A1(n4793), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4788) );
  OAI211_X1 U6005 ( .C1(n4796), .C2(n6421), .A(n4789), .B(n4788), .ZN(U3088)
         );
  OAI22_X1 U6006 ( .A1(n5111), .A2(n4791), .B1(n4790), .B2(n5110), .ZN(n4792)
         );
  AOI21_X1 U6007 ( .B1(n6428), .B2(n6466), .A(n4792), .ZN(n4795) );
  NAND2_X1 U6008 ( .A1(n4793), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4794) );
  OAI211_X1 U6009 ( .C1(n4796), .C2(n6431), .A(n4795), .B(n4794), .ZN(U3090)
         );
  AOI21_X1 U6010 ( .B1(n4835), .B2(n4804), .A(n6735), .ZN(n4799) );
  AOI211_X1 U6011 ( .C1(n4844), .C2(n6107), .A(n6392), .B(n4799), .ZN(n4803)
         );
  NAND2_X1 U6012 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4800), .ZN(n4846) );
  NOR2_X1 U6013 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4846), .ZN(n4836)
         );
  OAI211_X1 U6014 ( .C1(n4836), .C2(n5105), .A(n4801), .B(n5107), .ZN(n4802)
         );
  INV_X1 U6015 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4810) );
  INV_X1 U6016 ( .A(n6107), .ZN(n4924) );
  OAI22_X1 U6017 ( .A1(n4806), .A2(n4924), .B1(n4926), .B2(n4805), .ZN(n4837)
         );
  AOI22_X1 U6018 ( .A1(n6461), .A2(n4836), .B1(n6462), .B2(n4837), .ZN(n4807)
         );
  OAI21_X1 U6019 ( .B1(n6465), .B2(n4835), .A(n4807), .ZN(n4808) );
  AOI21_X1 U6020 ( .B1(n6460), .B2(n4913), .A(n4808), .ZN(n4809) );
  OAI21_X1 U6021 ( .B1(n4841), .B2(n4810), .A(n4809), .ZN(U3121) );
  INV_X1 U6022 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4814) );
  AOI22_X1 U6023 ( .A1(n6441), .A2(n4836), .B1(n6442), .B2(n4837), .ZN(n4811)
         );
  OAI21_X1 U6024 ( .B1(n6445), .B2(n4835), .A(n4811), .ZN(n4812) );
  AOI21_X1 U6025 ( .B1(n6440), .B2(n4913), .A(n4812), .ZN(n4813) );
  OAI21_X1 U6026 ( .B1(n4841), .B2(n4814), .A(n4813), .ZN(U3116) );
  INV_X1 U6027 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4818) );
  AOI22_X1 U6028 ( .A1(n6489), .A2(n4836), .B1(n6491), .B2(n4837), .ZN(n4815)
         );
  OAI21_X1 U6029 ( .B1(n6496), .B2(n4835), .A(n4815), .ZN(n4816) );
  AOI21_X1 U6030 ( .B1(n6487), .B2(n4913), .A(n4816), .ZN(n4817) );
  OAI21_X1 U6031 ( .B1(n4841), .B2(n4818), .A(n4817), .ZN(U3123) );
  INV_X1 U6032 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4822) );
  AOI22_X1 U6033 ( .A1(n6447), .A2(n4836), .B1(n6448), .B2(n4837), .ZN(n4819)
         );
  OAI21_X1 U6034 ( .B1(n6451), .B2(n4835), .A(n4819), .ZN(n4820) );
  AOI21_X1 U6035 ( .B1(n6446), .B2(n4913), .A(n4820), .ZN(n4821) );
  OAI21_X1 U6036 ( .B1(n4841), .B2(n4822), .A(n4821), .ZN(U3117) );
  INV_X1 U6037 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4826) );
  AOI22_X1 U6038 ( .A1(n6475), .A2(n4836), .B1(n6476), .B2(n4837), .ZN(n4823)
         );
  OAI21_X1 U6039 ( .B1(n6479), .B2(n4835), .A(n4823), .ZN(n4824) );
  AOI21_X1 U6040 ( .B1(n6474), .B2(n4913), .A(n4824), .ZN(n4825) );
  OAI21_X1 U6041 ( .B1(n4841), .B2(n4826), .A(n4825), .ZN(U3119) );
  INV_X1 U6042 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4830) );
  AOI22_X1 U6043 ( .A1(n6481), .A2(n4836), .B1(n6482), .B2(n4837), .ZN(n4827)
         );
  OAI21_X1 U6044 ( .B1(n6485), .B2(n4835), .A(n4827), .ZN(n4828) );
  AOI21_X1 U6045 ( .B1(n6480), .B2(n4913), .A(n4828), .ZN(n4829) );
  OAI21_X1 U6046 ( .B1(n4841), .B2(n4830), .A(n4829), .ZN(U3120) );
  INV_X1 U6047 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4834) );
  AOI22_X1 U6048 ( .A1(n6427), .A2(n4836), .B1(n6426), .B2(n4837), .ZN(n4831)
         );
  OAI21_X1 U6049 ( .B1(n5116), .B2(n4835), .A(n4831), .ZN(n4832) );
  AOI21_X1 U6050 ( .B1(n5113), .B2(n4913), .A(n4832), .ZN(n4833) );
  OAI21_X1 U6051 ( .B1(n4841), .B2(n4834), .A(n4833), .ZN(U3122) );
  INV_X1 U6052 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6185) );
  OAI222_X1 U6053 ( .A1(n6267), .A2(n5639), .B1(n5642), .B2(n6237), .C1(n5640), 
        .C2(n6185), .ZN(U2884) );
  INV_X1 U6054 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4840) );
  INV_X1 U6055 ( .A(n4835), .ZN(n6486) );
  AOI22_X1 U6056 ( .A1(n6453), .A2(n4836), .B1(n6410), .B2(n6486), .ZN(n4839)
         );
  AOI22_X1 U6057 ( .A1(n6454), .A2(n4837), .B1(n6452), .B2(n4913), .ZN(n4838)
         );
  OAI211_X1 U6058 ( .C1(n4841), .C2(n4840), .A(n4839), .B(n4838), .ZN(U3118)
         );
  INV_X1 U6059 ( .A(n4842), .ZN(n4843) );
  NAND2_X1 U6060 ( .A1(n4843), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4862) );
  NAND2_X1 U6061 ( .A1(n6395), .A2(n4862), .ZN(n4851) );
  NOR2_X1 U6062 ( .A1(n6917), .A2(n4846), .ZN(n4914) );
  AOI21_X1 U6063 ( .B1(n4845), .B2(n4844), .A(n4914), .ZN(n4852) );
  INV_X1 U6064 ( .A(n4852), .ZN(n4848) );
  AOI21_X1 U6065 ( .B1(n6392), .B2(n4846), .A(n5012), .ZN(n4847) );
  OAI21_X1 U6066 ( .B1(n4851), .B2(n4848), .A(n4847), .ZN(n4912) );
  NAND2_X1 U6067 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4849) );
  OAI22_X1 U6068 ( .A1(n4852), .A2(n4851), .B1(n4850), .B2(n4849), .ZN(n4911)
         );
  AOI22_X1 U6069 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4912), .B1(n6476), 
        .B2(n4911), .ZN(n4854) );
  AOI22_X1 U6070 ( .A1(n6475), .A2(n4914), .B1(n6414), .B2(n4913), .ZN(n4853)
         );
  OAI211_X1 U6071 ( .C1(n6417), .C2(n4958), .A(n4854), .B(n4853), .ZN(U3127)
         );
  AOI22_X1 U6072 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4912), .B1(n6491), 
        .B2(n4911), .ZN(n4856) );
  AOI22_X1 U6073 ( .A1(n6489), .A2(n4914), .B1(n6435), .B2(n4913), .ZN(n4855)
         );
  OAI211_X1 U6074 ( .C1(n6439), .C2(n4958), .A(n4856), .B(n4855), .ZN(U3131)
         );
  AOI22_X1 U6075 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4912), .B1(n6482), 
        .B2(n4911), .ZN(n4858) );
  AOI22_X1 U6076 ( .A1(n6481), .A2(n4914), .B1(n6418), .B2(n4913), .ZN(n4857)
         );
  OAI211_X1 U6077 ( .C1(n6421), .C2(n4958), .A(n4858), .B(n4857), .ZN(U3128)
         );
  AOI22_X1 U6078 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4912), .B1(n6454), 
        .B2(n4911), .ZN(n4860) );
  AOI22_X1 U6079 ( .A1(n6453), .A2(n4914), .B1(n6410), .B2(n4913), .ZN(n4859)
         );
  OAI211_X1 U6080 ( .C1(n6413), .C2(n4958), .A(n4860), .B(n4859), .ZN(U3126)
         );
  AND2_X1 U6081 ( .A1(n4862), .A2(n4861), .ZN(n5802) );
  NOR2_X1 U6082 ( .A1(n4875), .A2(n4863), .ZN(n4864) );
  AOI21_X1 U6083 ( .B1(n5802), .B2(n4864), .A(n6392), .ZN(n4870) );
  NOR2_X1 U6084 ( .A1(n4866), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4876)
         );
  AOI21_X1 U6085 ( .B1(n5109), .B2(n4867), .A(n4876), .ZN(n4869) );
  INV_X1 U6086 ( .A(n4869), .ZN(n4868) );
  NAND3_X1 U6087 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6734), .A3(n6505), .ZN(n5100) );
  INV_X1 U6088 ( .A(n5100), .ZN(n4873) );
  AOI22_X1 U6089 ( .A1(n4870), .A2(n4868), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4873), .ZN(n4904) );
  INV_X1 U6090 ( .A(n5012), .ZN(n4872) );
  NAND2_X1 U6091 ( .A1(n4870), .A2(n4869), .ZN(n4871) );
  OAI211_X1 U6092 ( .C1(n6395), .C2(n4873), .A(n4872), .B(n4871), .ZN(n4898)
         );
  NAND2_X1 U6093 ( .A1(n4898), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4879) );
  OR3_X1 U6094 ( .A1(n4875), .A2(n5800), .A3(n4874), .ZN(n5117) );
  INV_X1 U6095 ( .A(n4876), .ZN(n4900) );
  OAI22_X1 U6096 ( .A1(n5118), .A2(n4900), .B1(n6413), .B2(n4899), .ZN(n4877)
         );
  AOI21_X1 U6097 ( .B1(n6410), .B2(n5155), .A(n4877), .ZN(n4878) );
  OAI211_X1 U6098 ( .C1(n4904), .C2(n5123), .A(n4879), .B(n4878), .ZN(U3046)
         );
  NAND2_X1 U6099 ( .A1(n4898), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4882) );
  OAI22_X1 U6100 ( .A1(n5145), .A2(n4900), .B1(n6421), .B2(n4899), .ZN(n4880)
         );
  AOI21_X1 U6101 ( .B1(n6418), .B2(n5155), .A(n4880), .ZN(n4881) );
  OAI211_X1 U6102 ( .C1(n4904), .C2(n5144), .A(n4882), .B(n4881), .ZN(U3048)
         );
  NAND2_X1 U6103 ( .A1(n4898), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4885) );
  OAI22_X1 U6104 ( .A1(n5140), .A2(n4900), .B1(n6409), .B2(n4899), .ZN(n4883)
         );
  AOI21_X1 U6105 ( .B1(n6406), .B2(n5155), .A(n4883), .ZN(n4884) );
  OAI211_X1 U6106 ( .C1(n4904), .C2(n5139), .A(n4885), .B(n4884), .ZN(U3045)
         );
  NAND2_X1 U6107 ( .A1(n4898), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4888) );
  OAI22_X1 U6108 ( .A1(n5130), .A2(n4900), .B1(n6439), .B2(n4899), .ZN(n4886)
         );
  AOI21_X1 U6109 ( .B1(n6435), .B2(n5155), .A(n4886), .ZN(n4887) );
  OAI211_X1 U6110 ( .C1(n4904), .C2(n5129), .A(n4888), .B(n4887), .ZN(U3051)
         );
  NAND2_X1 U6111 ( .A1(n4898), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4891) );
  OAI22_X1 U6112 ( .A1(n5125), .A2(n4900), .B1(n6405), .B2(n4899), .ZN(n4889)
         );
  AOI21_X1 U6113 ( .B1(n6402), .B2(n5155), .A(n4889), .ZN(n4890) );
  OAI211_X1 U6114 ( .C1(n4904), .C2(n5124), .A(n4891), .B(n4890), .ZN(U3044)
         );
  NAND2_X1 U6115 ( .A1(n4898), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4894) );
  OAI22_X1 U6116 ( .A1(n5153), .A2(n4900), .B1(n6425), .B2(n4899), .ZN(n4892)
         );
  AOI21_X1 U6117 ( .B1(n6422), .B2(n5155), .A(n4892), .ZN(n4893) );
  OAI211_X1 U6118 ( .C1(n4904), .C2(n5150), .A(n4894), .B(n4893), .ZN(U3049)
         );
  NAND2_X1 U6119 ( .A1(n4898), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4897) );
  OAI22_X1 U6120 ( .A1(n5135), .A2(n4900), .B1(n6417), .B2(n4899), .ZN(n4895)
         );
  AOI21_X1 U6121 ( .B1(n6414), .B2(n5155), .A(n4895), .ZN(n4896) );
  OAI211_X1 U6122 ( .C1(n4904), .C2(n5134), .A(n4897), .B(n4896), .ZN(U3047)
         );
  NAND2_X1 U6123 ( .A1(n4898), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4903) );
  OAI22_X1 U6124 ( .A1(n5111), .A2(n4900), .B1(n6431), .B2(n4899), .ZN(n4901)
         );
  AOI21_X1 U6125 ( .B1(n6428), .B2(n5155), .A(n4901), .ZN(n4902) );
  OAI211_X1 U6126 ( .C1(n4904), .C2(n5110), .A(n4903), .B(n4902), .ZN(U3050)
         );
  AOI22_X1 U6127 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4912), .B1(n6462), 
        .B2(n4911), .ZN(n4906) );
  AOI22_X1 U6128 ( .A1(n6461), .A2(n4914), .B1(n6422), .B2(n4913), .ZN(n4905)
         );
  OAI211_X1 U6129 ( .C1(n6425), .C2(n4958), .A(n4906), .B(n4905), .ZN(U3129)
         );
  AOI22_X1 U6130 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4912), .B1(n6442), 
        .B2(n4911), .ZN(n4908) );
  AOI22_X1 U6131 ( .A1(n6441), .A2(n4914), .B1(n6402), .B2(n4913), .ZN(n4907)
         );
  OAI211_X1 U6132 ( .C1(n6405), .C2(n4958), .A(n4908), .B(n4907), .ZN(U3124)
         );
  AOI22_X1 U6133 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4912), .B1(n6426), 
        .B2(n4911), .ZN(n4910) );
  AOI22_X1 U6134 ( .A1(n6427), .A2(n4914), .B1(n6428), .B2(n4913), .ZN(n4909)
         );
  OAI211_X1 U6135 ( .C1(n6431), .C2(n4958), .A(n4910), .B(n4909), .ZN(U3130)
         );
  AOI22_X1 U6136 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4912), .B1(n6448), 
        .B2(n4911), .ZN(n4916) );
  AOI22_X1 U6137 ( .A1(n6447), .A2(n4914), .B1(n6406), .B2(n4913), .ZN(n4915)
         );
  OAI211_X1 U6138 ( .C1(n6409), .C2(n4958), .A(n4916), .B(n4915), .ZN(U3125)
         );
  NOR2_X1 U6139 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4917), .ZN(n4923)
         );
  OAI21_X1 U6140 ( .B1(n6389), .B2(n6647), .A(n4918), .ZN(n6397) );
  NOR3_X1 U6141 ( .A1(n6397), .A2(n6734), .A3(n6398), .ZN(n4922) );
  INV_X1 U6142 ( .A(n4958), .ZN(n4919) );
  OAI21_X1 U6143 ( .B1(n4919), .B2(n4948), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4920) );
  NAND3_X1 U6144 ( .A1(n4925), .A2(n6395), .A3(n4920), .ZN(n4921) );
  OAI211_X1 U6145 ( .C1(n4923), .C2(n5105), .A(n4922), .B(n4921), .ZN(n4951)
         );
  NAND2_X1 U6146 ( .A1(n4951), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4930)
         );
  INV_X1 U6147 ( .A(n4923), .ZN(n4953) );
  INV_X1 U6148 ( .A(n6389), .ZN(n4927) );
  OAI33_X1 U6149 ( .A1(n6734), .A2(n4927), .A3(n4926), .B1(n4925), .B2(n6392), 
        .B3(n4924), .ZN(n4955) );
  INV_X1 U6150 ( .A(n4955), .ZN(n4946) );
  OAI22_X1 U6151 ( .A1(n5125), .A2(n4953), .B1(n4946), .B2(n5124), .ZN(n4928)
         );
  AOI21_X1 U6152 ( .B1(n6440), .B2(n4948), .A(n4928), .ZN(n4929) );
  OAI211_X1 U6153 ( .C1(n4958), .C2(n6445), .A(n4930), .B(n4929), .ZN(U3132)
         );
  NAND2_X1 U6154 ( .A1(n4951), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4933)
         );
  OAI22_X1 U6155 ( .A1(n5111), .A2(n4953), .B1(n4946), .B2(n5110), .ZN(n4931)
         );
  AOI21_X1 U6156 ( .B1(n5113), .B2(n4948), .A(n4931), .ZN(n4932) );
  OAI211_X1 U6157 ( .C1(n4958), .C2(n5116), .A(n4933), .B(n4932), .ZN(U3138)
         );
  NAND2_X1 U6158 ( .A1(n4951), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4936)
         );
  OAI22_X1 U6159 ( .A1(n5130), .A2(n4953), .B1(n4946), .B2(n5129), .ZN(n4934)
         );
  AOI21_X1 U6160 ( .B1(n6487), .B2(n4948), .A(n4934), .ZN(n4935) );
  OAI211_X1 U6161 ( .C1(n4958), .C2(n6496), .A(n4936), .B(n4935), .ZN(U3139)
         );
  NAND2_X1 U6162 ( .A1(n4951), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4939)
         );
  OAI22_X1 U6163 ( .A1(n5135), .A2(n4953), .B1(n4946), .B2(n5134), .ZN(n4937)
         );
  AOI21_X1 U6164 ( .B1(n6474), .B2(n4948), .A(n4937), .ZN(n4938) );
  OAI211_X1 U6165 ( .C1(n4958), .C2(n6479), .A(n4939), .B(n4938), .ZN(U3135)
         );
  NAND2_X1 U6166 ( .A1(n4951), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4942)
         );
  OAI22_X1 U6167 ( .A1(n5145), .A2(n4953), .B1(n4946), .B2(n5144), .ZN(n4940)
         );
  AOI21_X1 U6168 ( .B1(n6480), .B2(n4948), .A(n4940), .ZN(n4941) );
  OAI211_X1 U6169 ( .C1(n4958), .C2(n6485), .A(n4942), .B(n4941), .ZN(U3136)
         );
  NAND2_X1 U6170 ( .A1(n4951), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4945)
         );
  OAI22_X1 U6171 ( .A1(n5153), .A2(n4953), .B1(n4946), .B2(n5150), .ZN(n4943)
         );
  AOI21_X1 U6172 ( .B1(n6460), .B2(n4948), .A(n4943), .ZN(n4944) );
  OAI211_X1 U6173 ( .C1(n4958), .C2(n6465), .A(n4945), .B(n4944), .ZN(U3137)
         );
  NAND2_X1 U6174 ( .A1(n4951), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4950)
         );
  OAI22_X1 U6175 ( .A1(n5140), .A2(n4953), .B1(n4946), .B2(n5139), .ZN(n4947)
         );
  AOI21_X1 U6176 ( .B1(n6446), .B2(n4948), .A(n4947), .ZN(n4949) );
  OAI211_X1 U6177 ( .C1(n4958), .C2(n6451), .A(n4950), .B(n4949), .ZN(U3133)
         );
  NAND2_X1 U6178 ( .A1(n4951), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4957)
         );
  OAI22_X1 U6179 ( .A1(n5118), .A2(n4953), .B1(n6413), .B2(n4952), .ZN(n4954)
         );
  AOI21_X1 U6180 ( .B1(n6454), .B2(n4955), .A(n4954), .ZN(n4956) );
  OAI211_X1 U6181 ( .C1(n4958), .C2(n6457), .A(n4957), .B(n4956), .ZN(U3134)
         );
  XOR2_X1 U6182 ( .A(n4960), .B(n4959), .Z(n6069) );
  INV_X1 U6183 ( .A(n6069), .ZN(n4967) );
  OR2_X1 U6184 ( .A1(n4962), .A2(n4961), .ZN(n4963) );
  NAND2_X1 U6185 ( .A1(n4963), .A2(n5061), .ZN(n6065) );
  INV_X1 U6186 ( .A(n6065), .ZN(n4964) );
  AOI22_X1 U6187 ( .A1(n6155), .A2(n4964), .B1(n5620), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n4965) );
  OAI21_X1 U6188 ( .B1(n4967), .B2(n5636), .A(n4965), .ZN(U2851) );
  AOI22_X1 U6189 ( .A1(n5342), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n6170), .ZN(n4966) );
  OAI21_X1 U6190 ( .B1(n4967), .B2(n5639), .A(n4966), .ZN(U2883) );
  OR2_X1 U6191 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4968), .ZN(n5002)
         );
  AOI211_X1 U6192 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5002), .A(n6390), .B(
        n4969), .ZN(n4974) );
  INV_X1 U6193 ( .A(n4999), .ZN(n5004) );
  NOR3_X1 U6194 ( .A1(n5004), .A2(n4996), .A3(n6392), .ZN(n4972) );
  OAI21_X1 U6195 ( .B1(n4972), .B2(n4971), .A(n4970), .ZN(n4973) );
  NAND2_X1 U6196 ( .A1(n4974), .A2(n4973), .ZN(n5000) );
  NAND2_X1 U6197 ( .A1(n5000), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4979) );
  AOI22_X1 U6198 ( .A1(n4976), .A2(n6395), .B1(n6398), .B2(n4975), .ZN(n5007)
         );
  OAI22_X1 U6199 ( .A1(n5140), .A2(n5002), .B1(n5007), .B2(n5139), .ZN(n4977)
         );
  AOI21_X1 U6200 ( .B1(n6406), .B2(n4996), .A(n4977), .ZN(n4978) );
  OAI211_X1 U6201 ( .C1(n4999), .C2(n6409), .A(n4979), .B(n4978), .ZN(U3021)
         );
  NAND2_X1 U6202 ( .A1(n5000), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4982) );
  OAI22_X1 U6203 ( .A1(n5130), .A2(n5002), .B1(n5007), .B2(n5129), .ZN(n4980)
         );
  AOI21_X1 U6204 ( .B1(n6435), .B2(n4996), .A(n4980), .ZN(n4981) );
  OAI211_X1 U6205 ( .C1(n4999), .C2(n6439), .A(n4982), .B(n4981), .ZN(U3027)
         );
  NAND2_X1 U6206 ( .A1(n5000), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4985) );
  OAI22_X1 U6207 ( .A1(n5125), .A2(n5002), .B1(n5007), .B2(n5124), .ZN(n4983)
         );
  AOI21_X1 U6208 ( .B1(n6402), .B2(n4996), .A(n4983), .ZN(n4984) );
  OAI211_X1 U6209 ( .C1(n4999), .C2(n6405), .A(n4985), .B(n4984), .ZN(U3020)
         );
  NAND2_X1 U6210 ( .A1(n5000), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4988) );
  OAI22_X1 U6211 ( .A1(n5135), .A2(n5002), .B1(n5007), .B2(n5134), .ZN(n4986)
         );
  AOI21_X1 U6212 ( .B1(n6414), .B2(n4996), .A(n4986), .ZN(n4987) );
  OAI211_X1 U6213 ( .C1(n4999), .C2(n6417), .A(n4988), .B(n4987), .ZN(U3023)
         );
  NAND2_X1 U6214 ( .A1(n5000), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4991) );
  OAI22_X1 U6215 ( .A1(n5145), .A2(n5002), .B1(n5007), .B2(n5144), .ZN(n4989)
         );
  AOI21_X1 U6216 ( .B1(n6418), .B2(n4996), .A(n4989), .ZN(n4990) );
  OAI211_X1 U6217 ( .C1(n4999), .C2(n6421), .A(n4991), .B(n4990), .ZN(U3024)
         );
  NAND2_X1 U6218 ( .A1(n5000), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4994) );
  OAI22_X1 U6219 ( .A1(n5153), .A2(n5002), .B1(n5007), .B2(n5150), .ZN(n4992)
         );
  AOI21_X1 U6220 ( .B1(n6422), .B2(n4996), .A(n4992), .ZN(n4993) );
  OAI211_X1 U6221 ( .C1(n4999), .C2(n6425), .A(n4994), .B(n4993), .ZN(U3025)
         );
  NAND2_X1 U6222 ( .A1(n5000), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4998) );
  OAI22_X1 U6223 ( .A1(n5111), .A2(n5002), .B1(n5007), .B2(n5110), .ZN(n4995)
         );
  AOI21_X1 U6224 ( .B1(n6428), .B2(n4996), .A(n4995), .ZN(n4997) );
  OAI211_X1 U6225 ( .C1(n4999), .C2(n6431), .A(n4998), .B(n4997), .ZN(U3026)
         );
  NAND2_X1 U6226 ( .A1(n5000), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5006) );
  OAI22_X1 U6227 ( .A1(n5118), .A2(n5002), .B1(n6457), .B2(n5001), .ZN(n5003)
         );
  AOI21_X1 U6228 ( .B1(n6452), .B2(n5004), .A(n5003), .ZN(n5005) );
  OAI211_X1 U6229 ( .C1(n5007), .C2(n5123), .A(n5006), .B(n5005), .ZN(U3022)
         );
  INV_X1 U6230 ( .A(n5008), .ZN(n5017) );
  OR2_X1 U6231 ( .A1(n5009), .A2(n5252), .ZN(n5011) );
  NOR2_X1 U6232 ( .A1(n6917), .A2(n5015), .ZN(n5048) );
  INV_X1 U6233 ( .A(n5048), .ZN(n5010) );
  NAND2_X1 U6234 ( .A1(n5011), .A2(n5010), .ZN(n5014) );
  NOR2_X1 U6235 ( .A1(n5017), .A2(n5014), .ZN(n5013) );
  INV_X1 U6236 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n5023) );
  INV_X1 U6237 ( .A(n5014), .ZN(n5016) );
  OAI22_X1 U6238 ( .A1(n5017), .A2(n5016), .B1(n5015), .B2(n6647), .ZN(n5052)
         );
  AOI22_X1 U6239 ( .A1(n6447), .A2(n5048), .B1(n6446), .B2(n6434), .ZN(n5020)
         );
  OAI21_X1 U6240 ( .B1(n6451), .B2(n5050), .A(n5020), .ZN(n5021) );
  AOI21_X1 U6241 ( .B1(n6448), .B2(n5052), .A(n5021), .ZN(n5022) );
  OAI21_X1 U6242 ( .B1(n5055), .B2(n5023), .A(n5022), .ZN(U3061) );
  INV_X1 U6243 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5027) );
  AOI22_X1 U6244 ( .A1(n6489), .A2(n5048), .B1(n6487), .B2(n6434), .ZN(n5024)
         );
  OAI21_X1 U6245 ( .B1(n6496), .B2(n5050), .A(n5024), .ZN(n5025) );
  AOI21_X1 U6246 ( .B1(n6491), .B2(n5052), .A(n5025), .ZN(n5026) );
  OAI21_X1 U6247 ( .B1(n5055), .B2(n5027), .A(n5026), .ZN(U3067) );
  INV_X1 U6248 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n5031) );
  AOI22_X1 U6249 ( .A1(n6475), .A2(n5048), .B1(n6474), .B2(n6434), .ZN(n5028)
         );
  OAI21_X1 U6250 ( .B1(n6479), .B2(n5050), .A(n5028), .ZN(n5029) );
  AOI21_X1 U6251 ( .B1(n6476), .B2(n5052), .A(n5029), .ZN(n5030) );
  OAI21_X1 U6252 ( .B1(n5055), .B2(n5031), .A(n5030), .ZN(U3063) );
  INV_X1 U6253 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n5035) );
  AOI22_X1 U6254 ( .A1(n6441), .A2(n5048), .B1(n6440), .B2(n6434), .ZN(n5032)
         );
  OAI21_X1 U6255 ( .B1(n6445), .B2(n5050), .A(n5032), .ZN(n5033) );
  AOI21_X1 U6256 ( .B1(n6442), .B2(n5052), .A(n5033), .ZN(n5034) );
  OAI21_X1 U6257 ( .B1(n5055), .B2(n5035), .A(n5034), .ZN(U3060) );
  INV_X1 U6258 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n5039) );
  AOI22_X1 U6259 ( .A1(n6461), .A2(n5048), .B1(n6460), .B2(n6434), .ZN(n5036)
         );
  OAI21_X1 U6260 ( .B1(n6465), .B2(n5050), .A(n5036), .ZN(n5037) );
  AOI21_X1 U6261 ( .B1(n6462), .B2(n5052), .A(n5037), .ZN(n5038) );
  OAI21_X1 U6262 ( .B1(n5055), .B2(n5039), .A(n5038), .ZN(U3065) );
  INV_X1 U6263 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5043) );
  AOI22_X1 U6264 ( .A1(n6481), .A2(n5048), .B1(n6480), .B2(n6434), .ZN(n5040)
         );
  OAI21_X1 U6265 ( .B1(n6485), .B2(n5050), .A(n5040), .ZN(n5041) );
  AOI21_X1 U6266 ( .B1(n6482), .B2(n5052), .A(n5041), .ZN(n5042) );
  OAI21_X1 U6267 ( .B1(n5055), .B2(n5043), .A(n5042), .ZN(U3064) );
  INV_X1 U6268 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n5047) );
  AOI22_X1 U6269 ( .A1(n6453), .A2(n5048), .B1(n6452), .B2(n6434), .ZN(n5044)
         );
  OAI21_X1 U6270 ( .B1(n6457), .B2(n5050), .A(n5044), .ZN(n5045) );
  AOI21_X1 U6271 ( .B1(n6454), .B2(n5052), .A(n5045), .ZN(n5046) );
  OAI21_X1 U6272 ( .B1(n5055), .B2(n5047), .A(n5046), .ZN(U3062) );
  INV_X1 U6273 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5054) );
  AOI22_X1 U6274 ( .A1(n6427), .A2(n5048), .B1(n5113), .B2(n6434), .ZN(n5049)
         );
  OAI21_X1 U6275 ( .B1(n5116), .B2(n5050), .A(n5049), .ZN(n5051) );
  AOI21_X1 U6276 ( .B1(n6426), .B2(n5052), .A(n5051), .ZN(n5053) );
  OAI21_X1 U6277 ( .B1(n5055), .B2(n5054), .A(n5053), .ZN(U3066) );
  NAND2_X1 U6278 ( .A1(n5058), .A2(n5057), .ZN(n5059) );
  NAND2_X1 U6279 ( .A1(n5211), .A2(n5059), .ZN(n5209) );
  AOI22_X1 U6280 ( .A1(n5342), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n6170), .ZN(n5060) );
  OAI21_X1 U6281 ( .B1(n5209), .B2(n5639), .A(n5060), .ZN(U2882) );
  AOI21_X1 U6282 ( .B1(n5062), .B2(n5061), .A(n5225), .ZN(n6316) );
  AOI22_X1 U6283 ( .A1(n6155), .A2(n6316), .B1(n5620), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n5063) );
  OAI21_X1 U6284 ( .B1(n5209), .B2(n5636), .A(n5063), .ZN(U2850) );
  NAND2_X1 U6285 ( .A1(n5064), .A2(n6495), .ZN(n5065) );
  AOI21_X1 U6286 ( .B1(n5065), .B2(STATEBS16_REG_SCAN_IN), .A(n6392), .ZN(
        n5070) );
  NOR2_X1 U6287 ( .A1(n5107), .A2(n6734), .ZN(n5066) );
  AOI22_X1 U6288 ( .A1(n5070), .A2(n5067), .B1(n6389), .B2(n5066), .ZN(n5099)
         );
  NOR2_X1 U6289 ( .A1(n6390), .A2(n6397), .ZN(n5103) );
  INV_X1 U6290 ( .A(n5067), .ZN(n5069) );
  OR2_X1 U6291 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5068), .ZN(n5094)
         );
  AOI22_X1 U6292 ( .A1(n5070), .A2(n5069), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5094), .ZN(n5071) );
  OAI211_X1 U6293 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6647), .A(n5103), .B(n5071), .ZN(n5093) );
  NAND2_X1 U6294 ( .A1(n5093), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5074)
         );
  OAI22_X1 U6295 ( .A1(n5145), .A2(n5094), .B1(n6495), .B2(n6421), .ZN(n5072)
         );
  AOI21_X1 U6296 ( .B1(n5096), .B2(n6418), .A(n5072), .ZN(n5073) );
  OAI211_X1 U6297 ( .C1(n5099), .C2(n5144), .A(n5074), .B(n5073), .ZN(U3104)
         );
  NAND2_X1 U6298 ( .A1(n5093), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5077)
         );
  OAI22_X1 U6299 ( .A1(n5153), .A2(n5094), .B1(n6495), .B2(n6425), .ZN(n5075)
         );
  AOI21_X1 U6300 ( .B1(n5096), .B2(n6422), .A(n5075), .ZN(n5076) );
  OAI211_X1 U6301 ( .C1(n5099), .C2(n5150), .A(n5077), .B(n5076), .ZN(U3105)
         );
  NAND2_X1 U6302 ( .A1(n5093), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5080)
         );
  OAI22_X1 U6303 ( .A1(n5111), .A2(n5094), .B1(n6495), .B2(n6431), .ZN(n5078)
         );
  AOI21_X1 U6304 ( .B1(n5096), .B2(n6428), .A(n5078), .ZN(n5079) );
  OAI211_X1 U6305 ( .C1(n5099), .C2(n5110), .A(n5080), .B(n5079), .ZN(U3106)
         );
  NAND2_X1 U6306 ( .A1(n5093), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5083)
         );
  OAI22_X1 U6307 ( .A1(n5135), .A2(n5094), .B1(n6495), .B2(n6417), .ZN(n5081)
         );
  AOI21_X1 U6308 ( .B1(n5096), .B2(n6414), .A(n5081), .ZN(n5082) );
  OAI211_X1 U6309 ( .C1(n5099), .C2(n5134), .A(n5083), .B(n5082), .ZN(U3103)
         );
  NAND2_X1 U6310 ( .A1(n5093), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5086)
         );
  OAI22_X1 U6311 ( .A1(n5140), .A2(n5094), .B1(n6495), .B2(n6409), .ZN(n5084)
         );
  AOI21_X1 U6312 ( .B1(n5096), .B2(n6406), .A(n5084), .ZN(n5085) );
  OAI211_X1 U6313 ( .C1(n5099), .C2(n5139), .A(n5086), .B(n5085), .ZN(U3101)
         );
  NAND2_X1 U6314 ( .A1(n5093), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5089)
         );
  OAI22_X1 U6315 ( .A1(n5118), .A2(n5094), .B1(n6495), .B2(n6413), .ZN(n5087)
         );
  AOI21_X1 U6316 ( .B1(n5096), .B2(n6410), .A(n5087), .ZN(n5088) );
  OAI211_X1 U6317 ( .C1(n5099), .C2(n5123), .A(n5089), .B(n5088), .ZN(U3102)
         );
  NAND2_X1 U6318 ( .A1(n5093), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5092)
         );
  OAI22_X1 U6319 ( .A1(n5130), .A2(n5094), .B1(n6495), .B2(n6439), .ZN(n5090)
         );
  AOI21_X1 U6320 ( .B1(n5096), .B2(n6435), .A(n5090), .ZN(n5091) );
  OAI211_X1 U6321 ( .C1(n5099), .C2(n5129), .A(n5092), .B(n5091), .ZN(U3107)
         );
  NAND2_X1 U6322 ( .A1(n5093), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5098)
         );
  OAI22_X1 U6323 ( .A1(n5125), .A2(n5094), .B1(n6495), .B2(n6405), .ZN(n5095)
         );
  AOI21_X1 U6324 ( .B1(n5096), .B2(n6402), .A(n5095), .ZN(n5097) );
  OAI211_X1 U6325 ( .C1(n5099), .C2(n5124), .A(n5098), .B(n5097), .ZN(U3100)
         );
  NOR2_X1 U6326 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5100), .ZN(n5106)
         );
  OAI21_X1 U6327 ( .B1(n5120), .B2(n5155), .A(n5806), .ZN(n5102) );
  INV_X1 U6328 ( .A(n5109), .ZN(n5101) );
  NAND2_X1 U6329 ( .A1(n5102), .A2(n5101), .ZN(n5104) );
  OAI221_X1 U6330 ( .B1(n5106), .B2(n5105), .C1(n5106), .C2(n5104), .A(n5103), 
        .ZN(n5149) );
  NAND2_X1 U6331 ( .A1(n5149), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5115) );
  INV_X1 U6332 ( .A(n5106), .ZN(n5152) );
  NOR2_X1 U6333 ( .A1(n5107), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5108)
         );
  AOI22_X1 U6334 ( .A1(n5109), .A2(n6395), .B1(n6389), .B2(n5108), .ZN(n5151)
         );
  OAI22_X1 U6335 ( .A1(n5111), .A2(n5152), .B1(n5151), .B2(n5110), .ZN(n5112)
         );
  AOI21_X1 U6336 ( .B1(n5113), .B2(n5155), .A(n5112), .ZN(n5114) );
  OAI211_X1 U6337 ( .C1(n5158), .C2(n5116), .A(n5115), .B(n5114), .ZN(U3042)
         );
  NAND2_X1 U6338 ( .A1(n5149), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5122) );
  OAI22_X1 U6339 ( .A1(n5118), .A2(n5152), .B1(n6413), .B2(n5117), .ZN(n5119)
         );
  AOI21_X1 U6340 ( .B1(n6410), .B2(n5120), .A(n5119), .ZN(n5121) );
  OAI211_X1 U6341 ( .C1(n5151), .C2(n5123), .A(n5122), .B(n5121), .ZN(U3038)
         );
  NAND2_X1 U6342 ( .A1(n5149), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5128) );
  OAI22_X1 U6343 ( .A1(n5125), .A2(n5152), .B1(n5151), .B2(n5124), .ZN(n5126)
         );
  AOI21_X1 U6344 ( .B1(n6440), .B2(n5155), .A(n5126), .ZN(n5127) );
  OAI211_X1 U6345 ( .C1(n6445), .C2(n5158), .A(n5128), .B(n5127), .ZN(U3036)
         );
  NAND2_X1 U6346 ( .A1(n5149), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5133) );
  OAI22_X1 U6347 ( .A1(n5130), .A2(n5152), .B1(n5151), .B2(n5129), .ZN(n5131)
         );
  AOI21_X1 U6348 ( .B1(n6487), .B2(n5155), .A(n5131), .ZN(n5132) );
  OAI211_X1 U6349 ( .C1(n5158), .C2(n6496), .A(n5133), .B(n5132), .ZN(U3043)
         );
  NAND2_X1 U6350 ( .A1(n5149), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5138) );
  OAI22_X1 U6351 ( .A1(n5135), .A2(n5152), .B1(n5151), .B2(n5134), .ZN(n5136)
         );
  AOI21_X1 U6352 ( .B1(n6474), .B2(n5155), .A(n5136), .ZN(n5137) );
  OAI211_X1 U6353 ( .C1(n5158), .C2(n6479), .A(n5138), .B(n5137), .ZN(U3039)
         );
  NAND2_X1 U6354 ( .A1(n5149), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5143) );
  OAI22_X1 U6355 ( .A1(n5140), .A2(n5152), .B1(n5151), .B2(n5139), .ZN(n5141)
         );
  AOI21_X1 U6356 ( .B1(n6446), .B2(n5155), .A(n5141), .ZN(n5142) );
  OAI211_X1 U6357 ( .C1(n5158), .C2(n6451), .A(n5143), .B(n5142), .ZN(U3037)
         );
  NAND2_X1 U6358 ( .A1(n5149), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5148) );
  OAI22_X1 U6359 ( .A1(n5145), .A2(n5152), .B1(n5151), .B2(n5144), .ZN(n5146)
         );
  AOI21_X1 U6360 ( .B1(n6480), .B2(n5155), .A(n5146), .ZN(n5147) );
  OAI211_X1 U6361 ( .C1(n5158), .C2(n6485), .A(n5148), .B(n5147), .ZN(U3040)
         );
  NAND2_X1 U6362 ( .A1(n5149), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5157) );
  OAI22_X1 U6363 ( .A1(n5153), .A2(n5152), .B1(n5151), .B2(n5150), .ZN(n5154)
         );
  AOI21_X1 U6364 ( .B1(n6460), .B2(n5155), .A(n5154), .ZN(n5156) );
  OAI211_X1 U6365 ( .C1(n5158), .C2(n6465), .A(n5157), .B(n5156), .ZN(U3041)
         );
  NOR2_X1 U6366 ( .A1(n6574), .A2(n6074), .ZN(n6078) );
  NAND3_X1 U6367 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        n6078), .ZN(n6064) );
  INV_X1 U6368 ( .A(n6064), .ZN(n5160) );
  INV_X1 U6369 ( .A(n6148), .ZN(n6111) );
  OAI21_X1 U6370 ( .B1(n6111), .B2(n5159), .A(n5886), .ZN(n6073) );
  OAI21_X1 U6371 ( .B1(n6064), .B2(REIP_REG_9__SCAN_IN), .A(n6073), .ZN(n6060)
         );
  OAI21_X1 U6372 ( .B1(REIP_REG_9__SCAN_IN), .B2(n5160), .A(n6060), .ZN(n5165)
         );
  INV_X1 U6373 ( .A(n5161), .ZN(n5206) );
  AOI22_X1 U6374 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6115), .B1(n6083), .B2(n6316), 
        .ZN(n5162) );
  OAI211_X1 U6375 ( .C1(n6105), .C2(n5204), .A(n5162), .B(n6085), .ZN(n5163)
         );
  AOI21_X1 U6376 ( .B1(n6133), .B2(n5206), .A(n5163), .ZN(n5164) );
  OAI211_X1 U6377 ( .C1(n5890), .C2(n5209), .A(n5165), .B(n5164), .ZN(U2818)
         );
  OR2_X1 U6378 ( .A1(n5167), .A2(n5166), .ZN(n5168) );
  NAND2_X1 U6379 ( .A1(n5169), .A2(n5168), .ZN(n6355) );
  INV_X1 U6380 ( .A(n5170), .ZN(n6097) );
  AOI22_X1 U6381 ( .A1(n6288), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n6340), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n5171) );
  OAI21_X1 U6382 ( .B1(n6296), .B2(n6097), .A(n5171), .ZN(n5172) );
  AOI21_X1 U6383 ( .B1(n5173), .B2(n3099), .A(n5172), .ZN(n5174) );
  OAI21_X1 U6384 ( .B1(n5984), .B2(n6355), .A(n5174), .ZN(U2982) );
  INV_X1 U6385 ( .A(n6144), .ZN(n5178) );
  AOI21_X1 U6386 ( .B1(n6288), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n5175), 
        .ZN(n5176) );
  OAI21_X1 U6387 ( .B1(n6296), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n5176), 
        .ZN(n5177) );
  AOI21_X1 U6388 ( .B1(n5178), .B2(n3099), .A(n5177), .ZN(n5179) );
  OAI21_X1 U6389 ( .B1(n5180), .B2(n5984), .A(n5179), .ZN(U2985) );
  OAI21_X1 U6390 ( .B1(n5181), .B2(n5183), .A(n5182), .ZN(n5199) );
  OAI22_X1 U6391 ( .A1(n5186), .A2(n5185), .B1(n5758), .B2(n5184), .ZN(n6324)
         );
  INV_X1 U6392 ( .A(n6324), .ZN(n5188) );
  NOR2_X1 U6393 ( .A1(n6369), .A2(n6373), .ZN(n6345) );
  OAI21_X1 U6394 ( .B1(n6375), .B2(n6345), .A(n6371), .ZN(n6368) );
  NOR3_X1 U6395 ( .A1(n5187), .A2(n6343), .A3(n6368), .ZN(n6336) );
  NAND2_X1 U6396 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6336), .ZN(n5227)
         );
  OR2_X1 U6397 ( .A1(n5227), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6325)
         );
  AOI21_X1 U6398 ( .B1(n5188), .B2(n6325), .A(n6799), .ZN(n5192) );
  NOR3_X1 U6399 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n5189), .A3(n5227), 
        .ZN(n5191) );
  NAND2_X1 U6400 ( .A1(n6340), .A2(REIP_REG_8__SCAN_IN), .ZN(n5195) );
  OAI21_X1 U6401 ( .B1(n6378), .B2(n6065), .A(n5195), .ZN(n5190) );
  NOR3_X1 U6402 ( .A1(n5192), .A2(n5191), .A3(n5190), .ZN(n5193) );
  OAI21_X1 U6403 ( .B1(n6354), .B2(n5199), .A(n5193), .ZN(U3010) );
  INV_X1 U6404 ( .A(n6068), .ZN(n5196) );
  NAND2_X1 U6405 ( .A1(n6288), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5194)
         );
  OAI211_X1 U6406 ( .C1(n6296), .C2(n5196), .A(n5195), .B(n5194), .ZN(n5197)
         );
  AOI21_X1 U6407 ( .B1(n6069), .B2(n3099), .A(n5197), .ZN(n5198) );
  OAI21_X1 U6408 ( .B1(n5199), .B2(n5984), .A(n5198), .ZN(U2978) );
  NAND2_X1 U6409 ( .A1(n5202), .A2(n5201), .ZN(n5203) );
  XNOR2_X1 U6410 ( .A(n5200), .B(n5203), .ZN(n6317) );
  INV_X1 U6411 ( .A(n5984), .ZN(n6293) );
  NAND2_X1 U6412 ( .A1(n6317), .A2(n6293), .ZN(n5208) );
  INV_X1 U6413 ( .A(n6296), .ZN(n5701) );
  NAND2_X1 U6414 ( .A1(n6340), .A2(REIP_REG_9__SCAN_IN), .ZN(n6314) );
  OAI21_X1 U6415 ( .B1(n5699), .B2(n5204), .A(n6314), .ZN(n5205) );
  AOI21_X1 U6416 ( .B1(n5701), .B2(n5206), .A(n5205), .ZN(n5207) );
  OAI211_X1 U6417 ( .C1(n6266), .C2(n5209), .A(n5208), .B(n5207), .ZN(U2977)
         );
  AOI21_X1 U6418 ( .B1(n5212), .B2(n5211), .A(n5215), .ZN(n6059) );
  INV_X1 U6419 ( .A(n6059), .ZN(n5243) );
  AOI22_X1 U6420 ( .A1(n5342), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n6170), .ZN(n5213) );
  OAI21_X1 U6421 ( .B1(n5243), .B2(n5639), .A(n5213), .ZN(U2881) );
  NOR2_X1 U6422 ( .A1(n5215), .A2(n5214), .ZN(n5216) );
  OR2_X1 U6423 ( .A1(n5263), .A2(n5216), .ZN(n5287) );
  AOI22_X1 U6424 ( .A1(n5342), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n6170), .ZN(n5217) );
  OAI21_X1 U6425 ( .B1(n5287), .B2(n5639), .A(n5217), .ZN(U2880) );
  AOI21_X1 U6426 ( .B1(n5218), .B2(n5224), .A(n5259), .ZN(n6307) );
  AOI22_X1 U6427 ( .A1(n6155), .A2(n6307), .B1(n5620), .B2(EBX_REG_11__SCAN_IN), .ZN(n5219) );
  OAI21_X1 U6428 ( .B1(n5287), .B2(n5636), .A(n5219), .ZN(U2848) );
  NAND2_X1 U6429 ( .A1(n5279), .A2(n5220), .ZN(n5223) );
  XOR2_X1 U6430 ( .A(n5223), .B(n5222), .Z(n5249) );
  AOI21_X1 U6431 ( .B1(n5228), .B2(n6331), .A(n6324), .ZN(n6321) );
  INV_X1 U6432 ( .A(n6321), .ZN(n5233) );
  OAI21_X1 U6433 ( .B1(n5226), .B2(n5225), .A(n5224), .ZN(n6057) );
  INV_X1 U6434 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6579) );
  OAI22_X1 U6435 ( .A1(n6378), .A2(n6057), .B1(n6579), .B2(n6376), .ZN(n5232)
         );
  NOR2_X1 U6436 ( .A1(n5228), .A2(n5227), .ZN(n6318) );
  OAI211_X1 U6437 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6318), .B(n5229), .ZN(n5230) );
  INV_X1 U6438 ( .A(n5230), .ZN(n5231) );
  AOI211_X1 U6439 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n5233), .A(n5232), .B(n5231), .ZN(n5234) );
  OAI21_X1 U6440 ( .B1(n5249), .B2(n6354), .A(n5234), .ZN(U3008) );
  NOR2_X1 U6441 ( .A1(n5235), .A2(n6064), .ZN(n5344) );
  AND2_X1 U6442 ( .A1(n5886), .A2(n5236), .ZN(n6046) );
  OAI21_X1 U6443 ( .B1(REIP_REG_11__SCAN_IN), .B2(n5344), .A(n6046), .ZN(n5242) );
  INV_X1 U6444 ( .A(n5283), .ZN(n5240) );
  AOI22_X1 U6445 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n6130), .B1(n6083), 
        .B2(n6307), .ZN(n5237) );
  OAI211_X1 U6446 ( .C1(n6138), .C2(n5238), .A(n5237), .B(n6085), .ZN(n5239)
         );
  AOI21_X1 U6447 ( .B1(n6133), .B2(n5240), .A(n5239), .ZN(n5241) );
  OAI211_X1 U6448 ( .C1(n5890), .C2(n5287), .A(n5242), .B(n5241), .ZN(U2816)
         );
  OAI222_X1 U6449 ( .A1(n6057), .A2(n6150), .B1(n5244), .B2(n6159), .C1(n5636), 
        .C2(n5243), .ZN(U2849) );
  AOI22_X1 U6450 ( .A1(n6288), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6340), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5245) );
  OAI21_X1 U6451 ( .B1(n6296), .B2(n5246), .A(n5245), .ZN(n5247) );
  AOI21_X1 U6452 ( .B1(n6059), .B2(n3099), .A(n5247), .ZN(n5248) );
  OAI21_X1 U6453 ( .B1(n5249), .B2(n5984), .A(n5248), .ZN(U2976) );
  OR2_X1 U6454 ( .A1(n5513), .A2(n3563), .ZN(n5250) );
  NAND2_X1 U6455 ( .A1(n5250), .A2(n5890), .ZN(n6126) );
  INV_X1 U6456 ( .A(n6126), .ZN(n6143) );
  OR2_X1 U6457 ( .A1(n5513), .A2(n5251), .ZN(n6137) );
  OAI22_X1 U6458 ( .A1(n6143), .A2(n5253), .B1(n5252), .B2(n6137), .ZN(n5254)
         );
  AOI21_X1 U6459 ( .B1(REIP_REG_0__SCAN_IN), .B2(n5886), .A(n5254), .ZN(n5257)
         );
  NAND2_X1 U6460 ( .A1(n6105), .A2(n6128), .ZN(n5255) );
  AOI22_X1 U6461 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n5255), .B1(n6115), 
        .B2(EBX_REG_0__SCAN_IN), .ZN(n5256) );
  OAI211_X1 U6462 ( .C1(n6120), .C2(n5258), .A(n5257), .B(n5256), .ZN(U2827)
         );
  OAI21_X1 U6463 ( .B1(n5260), .B2(n5259), .A(n5310), .ZN(n6300) );
  OAI21_X1 U6464 ( .B1(n5263), .B2(n5262), .A(n5261), .ZN(n6049) );
  OAI222_X1 U6465 ( .A1(n6300), .A2(n6150), .B1(n5264), .B2(n6159), .C1(n5636), 
        .C2(n6049), .ZN(U2847) );
  INV_X1 U6466 ( .A(DATAI_12_), .ZN(n6219) );
  OAI222_X1 U6467 ( .A1(n6219), .A2(n5642), .B1(n5640), .B2(n3950), .C1(n5639), 
        .C2(n6049), .ZN(U2879) );
  NAND2_X1 U6468 ( .A1(n6274), .A2(n6273), .ZN(n6272) );
  NAND2_X1 U6469 ( .A1(n6272), .A2(n5266), .ZN(n5271) );
  AND2_X1 U6470 ( .A1(n5268), .A2(n5267), .ZN(n5269) );
  OAI21_X1 U6471 ( .B1(n5271), .B2(n5270), .A(n5269), .ZN(n5272) );
  INV_X1 U6472 ( .A(n5272), .ZN(n6335) );
  NAND2_X1 U6473 ( .A1(n6335), .A2(n6293), .ZN(n5277) );
  NOR2_X1 U6474 ( .A1(n6376), .A2(n6574), .ZN(n6333) );
  INV_X1 U6475 ( .A(n5273), .ZN(n5274) );
  NOR2_X1 U6476 ( .A1(n6296), .A2(n5274), .ZN(n5275) );
  AOI211_X1 U6477 ( .C1(n6288), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6333), 
        .B(n5275), .ZN(n5276) );
  OAI211_X1 U6478 ( .C1(n6266), .C2(n5278), .A(n5277), .B(n5276), .ZN(U2980)
         );
  NAND2_X1 U6479 ( .A1(n5280), .A2(n5279), .ZN(n5282) );
  XNOR2_X1 U6480 ( .A(n5693), .B(n6312), .ZN(n5281) );
  XNOR2_X1 U6481 ( .A(n5282), .B(n5281), .ZN(n6309) );
  NAND2_X1 U6482 ( .A1(n6309), .A2(n6293), .ZN(n5286) );
  NOR2_X1 U6483 ( .A1(n6376), .A2(n6582), .ZN(n6306) );
  NOR2_X1 U6484 ( .A1(n6296), .A2(n5283), .ZN(n5284) );
  AOI211_X1 U6485 ( .C1(n6288), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6306), 
        .B(n5284), .ZN(n5285) );
  OAI211_X1 U6486 ( .C1(n6266), .C2(n5287), .A(n5286), .B(n5285), .ZN(U2975)
         );
  NAND2_X1 U6487 ( .A1(n3105), .A2(n5288), .ZN(n5289) );
  XNOR2_X1 U6488 ( .A(n5290), .B(n5289), .ZN(n5340) );
  AOI22_X1 U6489 ( .A1(n6330), .A2(n5293), .B1(n5292), .B2(n5291), .ZN(n6313)
         );
  OAI21_X1 U6490 ( .B1(n5295), .B2(n5294), .A(n6313), .ZN(n5296) );
  AOI21_X1 U6491 ( .B1(n5297), .B2(n5389), .A(n5296), .ZN(n5970) );
  OAI21_X1 U6492 ( .B1(n5299), .B2(n5298), .A(n3539), .ZN(n5300) );
  AOI21_X1 U6493 ( .B1(n5970), .B2(n5300), .A(n5388), .ZN(n5304) );
  NOR3_X1 U6494 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5965), .A3(n5389), 
        .ZN(n5303) );
  OAI21_X1 U6495 ( .B1(n5301), .B2(n5309), .A(n5384), .ZN(n5637) );
  NAND2_X1 U6496 ( .A1(n6340), .A2(REIP_REG_14__SCAN_IN), .ZN(n5337) );
  OAI21_X1 U6497 ( .B1(n6378), .B2(n5637), .A(n5337), .ZN(n5302) );
  NOR3_X1 U6498 ( .A1(n5304), .A2(n5303), .A3(n5302), .ZN(n5305) );
  OAI21_X1 U6499 ( .B1(n5340), .B2(n6354), .A(n5305), .ZN(U3004) );
  NAND2_X1 U6500 ( .A1(n5307), .A2(n5306), .ZN(n5308) );
  NAND2_X1 U6501 ( .A1(n5334), .A2(n5308), .ZN(n6039) );
  AOI21_X1 U6502 ( .B1(n5311), .B2(n5310), .A(n5309), .ZN(n6035) );
  AOI22_X1 U6503 ( .A1(n6155), .A2(n6035), .B1(n5620), .B2(EBX_REG_13__SCAN_IN), .ZN(n5312) );
  OAI21_X1 U6504 ( .B1(n6039), .B2(n5636), .A(n5312), .ZN(U2846) );
  INV_X1 U6505 ( .A(n5323), .ZN(n5314) );
  NOR2_X1 U6506 ( .A1(n5321), .A2(n5314), .ZN(n5315) );
  XNOR2_X1 U6507 ( .A(n5322), .B(n5315), .ZN(n6301) );
  INV_X1 U6508 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5316) );
  OAI22_X1 U6509 ( .A1(n5699), .A2(n5317), .B1(n6376), .B2(n5316), .ZN(n5319)
         );
  NOR2_X1 U6510 ( .A1(n6049), .A2(n6266), .ZN(n5318) );
  AOI211_X1 U6511 ( .C1(n5701), .C2(n6050), .A(n5319), .B(n5318), .ZN(n5320)
         );
  OAI21_X1 U6512 ( .B1(n6301), .B2(n5984), .A(n5320), .ZN(U2974) );
  INV_X1 U6513 ( .A(DATAI_13_), .ZN(n6252) );
  OAI222_X1 U6514 ( .A1(n6039), .A2(n5639), .B1(n5642), .B2(n6252), .C1(n6178), 
        .C2(n5640), .ZN(U2878) );
  OR2_X1 U6515 ( .A1(n5322), .A2(n5321), .ZN(n5324) );
  NAND2_X1 U6516 ( .A1(n5324), .A2(n5323), .ZN(n5326) );
  XNOR2_X1 U6517 ( .A(n5326), .B(n5325), .ZN(n5967) );
  NAND2_X1 U6518 ( .A1(n5967), .A2(n6293), .ZN(n5330) );
  INV_X1 U6519 ( .A(REIP_REG_13__SCAN_IN), .ZN(n5327) );
  NOR2_X1 U6520 ( .A1(n6376), .A2(n5327), .ZN(n5964) );
  NOR2_X1 U6521 ( .A1(n6296), .A2(n6040), .ZN(n5328) );
  AOI211_X1 U6522 ( .C1(n6288), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5964), 
        .B(n5328), .ZN(n5329) );
  OAI211_X1 U6523 ( .C1(n6266), .C2(n6039), .A(n5330), .B(n5329), .ZN(U2973)
         );
  AND3_X1 U6524 ( .A1(n5334), .A2(n5333), .A3(n5332), .ZN(n5335) );
  NOR2_X1 U6525 ( .A1(n5394), .A2(n5335), .ZN(n5341) );
  NAND2_X1 U6526 ( .A1(n6288), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5336)
         );
  OAI211_X1 U6527 ( .C1(n6296), .C2(n5348), .A(n5337), .B(n5336), .ZN(n5338)
         );
  AOI21_X1 U6528 ( .B1(n5341), .B2(n3099), .A(n5338), .ZN(n5339) );
  OAI21_X1 U6529 ( .B1(n5340), .B2(n5984), .A(n5339), .ZN(U2972) );
  INV_X1 U6530 ( .A(n5341), .ZN(n5635) );
  AOI22_X1 U6531 ( .A1(n5342), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n6170), .ZN(n5343) );
  OAI21_X1 U6532 ( .B1(n5635), .B2(n5639), .A(n5343), .ZN(U2877) );
  NAND2_X1 U6533 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n6034) );
  NAND2_X1 U6534 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5344), .ZN(n6054) );
  INV_X1 U6535 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6585) );
  OAI21_X1 U6536 ( .B1(n6034), .B2(n6054), .A(n6585), .ZN(n5351) );
  INV_X1 U6537 ( .A(n5886), .ZN(n5854) );
  NOR2_X1 U6538 ( .A1(n5854), .A2(n5345), .ZN(n6026) );
  INV_X1 U6539 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5346) );
  OAI22_X1 U6540 ( .A1(n5346), .A2(n6105), .B1(n6120), .B2(n5637), .ZN(n5350)
         );
  NAND2_X1 U6541 ( .A1(n6115), .A2(EBX_REG_14__SCAN_IN), .ZN(n5347) );
  OAI211_X1 U6542 ( .C1(n6128), .C2(n5348), .A(n5347), .B(n6085), .ZN(n5349)
         );
  AOI211_X1 U6543 ( .C1(n5351), .C2(n6026), .A(n5350), .B(n5349), .ZN(n5352)
         );
  OAI21_X1 U6544 ( .B1(n5890), .B2(n5635), .A(n5352), .ZN(U2813) );
  OAI222_X1 U6545 ( .A1(n5636), .A2(n5655), .B1(n6159), .B2(n3744), .C1(n5726), 
        .C2(n6150), .ZN(U2833) );
  INV_X1 U6546 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6940) );
  NAND3_X1 U6547 ( .A1(n5664), .A2(n3556), .A3(n6940), .ZN(n5353) );
  AOI22_X1 U6548 ( .A1(n5643), .A2(n5353), .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n6940), .ZN(n5354) );
  XNOR2_X1 U6549 ( .A(n5354), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5709)
         );
  INV_X1 U6550 ( .A(n5822), .ZN(n5359) );
  AND2_X1 U6551 ( .A1(n6340), .A2(REIP_REG_28__SCAN_IN), .ZN(n5710) );
  AOI21_X1 U6552 ( .B1(n6288), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5710), 
        .ZN(n5358) );
  OAI21_X1 U6553 ( .B1(n6296), .B2(n5359), .A(n5358), .ZN(n5360) );
  AOI21_X1 U6554 ( .B1(n5901), .B2(n3099), .A(n5360), .ZN(n5361) );
  OAI21_X1 U6555 ( .B1(n5984), .B2(n5709), .A(n5361), .ZN(U2958) );
  INV_X1 U6556 ( .A(n5901), .ZN(n5366) );
  OR2_X1 U6557 ( .A1(n5558), .A2(n5362), .ZN(n5363) );
  AOI22_X1 U6558 ( .A1(n5823), .A2(n6155), .B1(n5620), .B2(EBX_REG_28__SCAN_IN), .ZN(n5365) );
  OAI21_X1 U6559 ( .B1(n5366), .B2(n5636), .A(n5365), .ZN(U2831) );
  NOR2_X1 U6560 ( .A1(n5774), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5773)
         );
  INV_X1 U6561 ( .A(n5367), .ZN(n5672) );
  AOI21_X1 U6562 ( .B1(n5672), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n3556), 
        .ZN(n5368) );
  NOR2_X1 U6563 ( .A1(n5773), .A2(n5368), .ZN(n5687) );
  XNOR2_X1 U6564 ( .A(n5693), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5686)
         );
  AOI22_X1 U6565 ( .A1(n5687), .A2(n5686), .B1(n3556), .B2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5681) );
  XNOR2_X1 U6566 ( .A(n5693), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5680)
         );
  NAND2_X1 U6567 ( .A1(n5681), .A2(n5680), .ZN(n5679) );
  NOR2_X1 U6568 ( .A1(n3556), .A2(n5744), .ZN(n5671) );
  OR2_X1 U6569 ( .A1(n5406), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5674)
         );
  INV_X1 U6570 ( .A(n5674), .ZN(n5369) );
  NOR2_X1 U6571 ( .A1(n5671), .A2(n5369), .ZN(n5370) );
  XNOR2_X1 U6572 ( .A(n5409), .B(n5370), .ZN(n5750) );
  NAND2_X1 U6573 ( .A1(n6340), .A2(REIP_REG_22__SCAN_IN), .ZN(n5742) );
  OAI21_X1 U6574 ( .B1(n5699), .B2(n5371), .A(n5742), .ZN(n5375) );
  NOR2_X1 U6575 ( .A1(n5862), .A2(n6266), .ZN(n5374) );
  AOI211_X1 U6576 ( .C1(n5701), .C2(n5856), .A(n5375), .B(n5374), .ZN(n5376)
         );
  OAI21_X1 U6577 ( .B1(n5750), .B2(n5984), .A(n5376), .ZN(U2964) );
  NOR2_X2 U6578 ( .A1(n6170), .A2(n5377), .ZN(n6171) );
  AOI22_X1 U6579 ( .A1(n6171), .A2(DATAI_6_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n6170), .ZN(n5380) );
  NAND2_X1 U6580 ( .A1(n6167), .A2(DATAI_22_), .ZN(n5379) );
  OAI211_X1 U6581 ( .C1(n5862), .C2(n5639), .A(n5380), .B(n5379), .ZN(U2869)
         );
  XNOR2_X1 U6582 ( .A(n5381), .B(n5588), .ZN(n5865) );
  OAI222_X1 U6583 ( .A1(n5862), .A2(n5601), .B1(n6150), .B2(n5865), .C1(n6159), 
        .C2(n5858), .ZN(U2837) );
  XNOR2_X1 U6584 ( .A(n5693), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5383)
         );
  XNOR2_X1 U6585 ( .A(n5382), .B(n5383), .ZN(n5403) );
  AOI21_X1 U6586 ( .B1(n5385), .B2(n5384), .A(n5631), .ZN(n6154) );
  NAND2_X1 U6587 ( .A1(n6340), .A2(REIP_REG_15__SCAN_IN), .ZN(n5399) );
  OAI21_X1 U6588 ( .B1(n5387), .B2(n5386), .A(n6313), .ZN(n5797) );
  NOR3_X1 U6589 ( .A1(n5965), .A2(n5389), .A3(n5388), .ZN(n5793) );
  AOI22_X1 U6590 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n5797), .B1(n5793), .B2(n5790), .ZN(n5390) );
  NAND2_X1 U6591 ( .A1(n5399), .A2(n5390), .ZN(n5391) );
  AOI21_X1 U6592 ( .B1(n6342), .B2(n6154), .A(n5391), .ZN(n5392) );
  OAI21_X1 U6593 ( .B1(n5403), .B2(n6354), .A(n5392), .ZN(U3003) );
  INV_X1 U6594 ( .A(n5393), .ZN(n5397) );
  INV_X1 U6595 ( .A(n5394), .ZN(n5396) );
  AOI21_X1 U6596 ( .B1(n5397), .B2(n5396), .A(n5634), .ZN(n6157) );
  INV_X1 U6597 ( .A(n6031), .ZN(n5400) );
  NAND2_X1 U6598 ( .A1(n6288), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5398)
         );
  OAI211_X1 U6599 ( .C1(n6296), .C2(n5400), .A(n5399), .B(n5398), .ZN(n5401)
         );
  AOI21_X1 U6600 ( .B1(n6157), .B2(n3099), .A(n5401), .ZN(n5402) );
  OAI21_X1 U6601 ( .B1(n5403), .B2(n5984), .A(n5402), .ZN(U2971) );
  AOI22_X1 U6602 ( .A1(n6171), .A2(DATAI_10_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6170), .ZN(n5405) );
  NAND2_X1 U6603 ( .A1(n6167), .A2(DATAI_26_), .ZN(n5404) );
  OAI211_X1 U6604 ( .C1(n5655), .C2(n5639), .A(n5405), .B(n5404), .ZN(U2865)
         );
  MUX2_X1 U6605 ( .A(n5744), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .S(n5406), 
        .Z(n5407) );
  OAI211_X1 U6606 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5409), .A(n5408), .B(n5407), .ZN(n5410) );
  XNOR2_X1 U6607 ( .A(n5410), .B(n5417), .ZN(n5422) );
  XNOR2_X2 U6608 ( .A(n5584), .B(n5412), .ZN(n5910) );
  NAND2_X1 U6609 ( .A1(n5701), .A2(n5837), .ZN(n5413) );
  NAND2_X1 U6610 ( .A1(n6340), .A2(REIP_REG_24__SCAN_IN), .ZN(n5418) );
  OAI211_X1 U6611 ( .C1(n5414), .C2(n5699), .A(n5413), .B(n5418), .ZN(n5415)
         );
  AOI21_X1 U6612 ( .B1(n5910), .B2(n3099), .A(n5415), .ZN(n5416) );
  OAI21_X1 U6613 ( .B1(n5422), .B2(n5984), .A(n5416), .ZN(U2962) );
  OAI21_X1 U6614 ( .B1(n5736), .B2(n6785), .A(n5417), .ZN(n5420) );
  XNOR2_X1 U6615 ( .A(n5590), .B(n5577), .ZN(n5839) );
  OAI21_X1 U6616 ( .B1(n6378), .B2(n5839), .A(n5418), .ZN(n5419) );
  AOI21_X1 U6617 ( .B1(n5420), .B2(n5941), .A(n5419), .ZN(n5421) );
  OAI21_X1 U6618 ( .B1(n5422), .B2(n6354), .A(n5421), .ZN(U2994) );
  AOI22_X1 U6619 ( .A1(n5812), .A2(n6155), .B1(EBX_REG_29__SCAN_IN), .B2(n5620), .ZN(n5423) );
  OAI21_X1 U6620 ( .B1(n5424), .B2(n5636), .A(n5423), .ZN(U2830) );
  NOR2_X1 U6621 ( .A1(n5426), .A2(n5425), .ZN(n5446) );
  AOI22_X1 U6622 ( .A1(n3391), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3299), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5432) );
  AOI22_X1 U6623 ( .A1(n4315), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4320), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5431) );
  AOI22_X1 U6624 ( .A1(n4117), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5430) );
  AOI22_X1 U6625 ( .A1(n5428), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5427), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n5429) );
  NAND4_X1 U6626 ( .A1(n5432), .A2(n5431), .A3(n5430), .A4(n5429), .ZN(n5444)
         );
  AOI22_X1 U6627 ( .A1(n5434), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5433), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5442) );
  AOI22_X1 U6628 ( .A1(n3101), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5435), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5441) );
  AOI22_X1 U6629 ( .A1(n3370), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n5436), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5440) );
  AOI22_X1 U6630 ( .A1(n5438), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n5437), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5439) );
  NAND4_X1 U6631 ( .A1(n5442), .A2(n5441), .A3(n5440), .A4(n5439), .ZN(n5443)
         );
  NOR2_X1 U6632 ( .A1(n5444), .A2(n5443), .ZN(n5445) );
  XNOR2_X1 U6633 ( .A(n5446), .B(n5445), .ZN(n5448) );
  NAND2_X1 U6634 ( .A1(n5448), .A2(n5447), .ZN(n5455) );
  OAI21_X1 U6635 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5459), .A(n5449), .ZN(
        n5450) );
  AOI21_X1 U6636 ( .B1(n5502), .B2(EAX_REG_30__SCAN_IN), .A(n5450), .ZN(n5454)
         );
  XNOR2_X1 U6637 ( .A(n5451), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5457)
         );
  AND2_X1 U6638 ( .A1(n5457), .A2(n5452), .ZN(n5453) );
  AOI21_X1 U6639 ( .B1(n5455), .B2(n5454), .A(n5453), .ZN(n5497) );
  XNOR2_X1 U6640 ( .A(n5497), .B(n5470), .ZN(n5468) );
  INV_X1 U6641 ( .A(n5466), .ZN(n5456) );
  INV_X1 U6642 ( .A(EBX_REG_30__SCAN_IN), .ZN(n6756) );
  OAI222_X1 U6643 ( .A1(n5468), .A2(n5601), .B1(n6150), .B2(n5456), .C1(n6159), 
        .C2(n6756), .ZN(U2829) );
  INV_X1 U6644 ( .A(n5457), .ZN(n5473) );
  INV_X1 U6645 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6816) );
  INV_X1 U6646 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6606) );
  NOR2_X1 U6647 ( .A1(n6816), .A2(n6606), .ZN(n5458) );
  OAI21_X1 U6648 ( .B1(n5458), .B2(n6110), .A(n5554), .ZN(n5821) );
  INV_X1 U6649 ( .A(REIP_REG_29__SCAN_IN), .ZN(n5815) );
  NOR2_X1 U6650 ( .A1(n5821), .A2(n5815), .ZN(n5813) );
  INV_X1 U6651 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6615) );
  NOR3_X1 U6652 ( .A1(n5854), .A2(n5813), .A3(n6615), .ZN(n5461) );
  OAI22_X1 U6653 ( .A1(n6756), .A2(n6138), .B1(n5459), .B2(n6105), .ZN(n5460)
         );
  NOR2_X1 U6654 ( .A1(n5461), .A2(n5460), .ZN(n5464) );
  NOR2_X1 U6655 ( .A1(n5832), .A2(n5462), .ZN(n5824) );
  NAND3_X1 U6656 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .A3(
        n5824), .ZN(n5814) );
  INV_X1 U6657 ( .A(n5814), .ZN(n5512) );
  NAND3_X1 U6658 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6615), .A3(n5512), .ZN(
        n5463) );
  OAI211_X1 U6659 ( .C1(n6128), .C2(n5473), .A(n5464), .B(n5463), .ZN(n5465)
         );
  AOI21_X1 U6660 ( .B1(n5466), .B2(n6083), .A(n5465), .ZN(n5467) );
  OAI21_X1 U6661 ( .B1(n5468), .B2(n5890), .A(n5467), .ZN(U2797) );
  AOI21_X1 U6662 ( .B1(n6288), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5471), 
        .ZN(n5472) );
  OAI21_X1 U6663 ( .B1(n6296), .B2(n5473), .A(n5472), .ZN(n5474) );
  OAI21_X1 U6664 ( .B1(n5476), .B2(n5984), .A(n5475), .ZN(U2956) );
  NOR3_X1 U6665 ( .A1(n5477), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5478) );
  AOI22_X1 U6666 ( .A1(n5479), .A2(n5489), .B1(n5664), .B2(n5478), .ZN(n5481)
         );
  XNOR2_X1 U6667 ( .A(n5481), .B(n5480), .ZN(n5511) );
  AOI22_X1 U6668 ( .A1(n5486), .A2(EBX_REG_31__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5485), .ZN(n5487) );
  XNOR2_X1 U6669 ( .A(n5488), .B(n5487), .ZN(n5564) );
  AND2_X1 U6670 ( .A1(n6340), .A2(REIP_REG_31__SCAN_IN), .ZN(n5506) );
  INV_X1 U6671 ( .A(n5489), .ZN(n5490) );
  NOR2_X1 U6672 ( .A1(n5491), .A2(n5490), .ZN(n5493) );
  MUX2_X1 U6673 ( .A(n5493), .B(n5492), .S(INSTADDRPOINTER_REG_31__SCAN_IN), 
        .Z(n5494) );
  AOI211_X1 U6674 ( .C1(n6342), .C2(n5564), .A(n5506), .B(n5494), .ZN(n5495)
         );
  OAI21_X1 U6675 ( .B1(n5511), .B2(n6354), .A(n5495), .ZN(U2987) );
  NAND2_X1 U6676 ( .A1(n5497), .A2(n5496), .ZN(n5499) );
  OR2_X1 U6677 ( .A1(n5499), .A2(n5498), .ZN(n5500) );
  AOI22_X1 U6678 ( .A1(n5502), .A2(EAX_REG_31__SCAN_IN), .B1(n5501), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5503) );
  INV_X1 U6679 ( .A(n5503), .ZN(n5504) );
  XNOR2_X2 U6680 ( .A(n5505), .B(n5504), .ZN(n5523) );
  AOI21_X1 U6681 ( .B1(n6288), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5506), 
        .ZN(n5507) );
  OAI21_X1 U6682 ( .B1(n6296), .B2(n5508), .A(n5507), .ZN(n5509) );
  OAI21_X1 U6683 ( .B1(n5511), .B2(n5984), .A(n5510), .ZN(U2955) );
  INV_X1 U6684 ( .A(n5523), .ZN(n5521) );
  INV_X1 U6685 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6749) );
  NAND4_X1 U6686 ( .A1(n6749), .A2(REIP_REG_30__SCAN_IN), .A3(
        REIP_REG_29__SCAN_IN), .A4(n5512), .ZN(n5516) );
  INV_X1 U6687 ( .A(n5513), .ZN(n5514) );
  NAND4_X1 U6688 ( .A1(n5514), .A2(n6648), .A3(EBX_REG_31__SCAN_IN), .A4(n6528), .ZN(n5515) );
  OAI211_X1 U6689 ( .C1(n6105), .C2(n5517), .A(n5516), .B(n5515), .ZN(n5519)
         );
  AOI211_X1 U6690 ( .C1(n5813), .C2(REIP_REG_30__SCAN_IN), .A(n5854), .B(n6749), .ZN(n5518) );
  AOI211_X1 U6691 ( .C1(n6083), .C2(n5564), .A(n5519), .B(n5518), .ZN(n5520)
         );
  OAI21_X1 U6692 ( .B1(n5521), .B2(n5890), .A(n5520), .ZN(U2796) );
  NAND3_X1 U6693 ( .A1(n5523), .A2(n5522), .A3(n5640), .ZN(n5525) );
  AOI22_X1 U6694 ( .A1(n6167), .A2(DATAI_31_), .B1(n6170), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U6695 ( .A1(n5525), .A2(n5524), .ZN(U2860) );
  INV_X1 U6696 ( .A(n6626), .ZN(n5527) );
  INV_X1 U6697 ( .A(n5528), .ZN(n5526) );
  INV_X1 U6698 ( .A(n6630), .ZN(n5535) );
  AOI21_X1 U6699 ( .B1(n5527), .B2(n5526), .A(n5535), .ZN(n5538) );
  NAND2_X1 U6700 ( .A1(n5528), .A2(n5537), .ZN(n5532) );
  INV_X1 U6701 ( .A(n5529), .ZN(n5531) );
  OAI22_X1 U6702 ( .A1(n6626), .A2(n5532), .B1(n5531), .B2(n5530), .ZN(n5533)
         );
  AOI21_X1 U6703 ( .B1(n5972), .B2(n5534), .A(n5533), .ZN(n5536) );
  OAI22_X1 U6704 ( .A1(n5538), .A2(n5537), .B1(n5536), .B2(n5535), .ZN(U3459)
         );
  NAND3_X1 U6705 ( .A1(n6516), .A2(n5540), .A3(n5539), .ZN(n5542) );
  AOI22_X1 U6706 ( .A1(n6532), .A2(n5542), .B1(n5546), .B2(n5541), .ZN(n5543)
         );
  OAI21_X1 U6707 ( .B1(n6532), .B2(n5544), .A(n5543), .ZN(n6517) );
  AOI21_X1 U6708 ( .B1(n5546), .B2(n5545), .A(n4234), .ZN(n5547) );
  AOI21_X1 U6709 ( .B1(n6532), .B2(n3563), .A(n5547), .ZN(n5978) );
  NAND2_X1 U6710 ( .A1(n5548), .A2(n6554), .ZN(n5549) );
  NAND2_X1 U6711 ( .A1(n5549), .A2(n3646), .ZN(n6646) );
  NAND2_X1 U6712 ( .A1(n5978), .A2(n6646), .ZN(n6513) );
  AND2_X1 U6713 ( .A1(n6513), .A2(n6525), .ZN(n5985) );
  MUX2_X1 U6714 ( .A(MORE_REG_SCAN_IN), .B(n6517), .S(n5985), .Z(U3471) );
  NAND2_X1 U6715 ( .A1(n5551), .A2(n5550), .ZN(n5552) );
  OAI22_X1 U6716 ( .A1(n4281), .A2(n6105), .B1(n6606), .B2(n5554), .ZN(n5562)
         );
  AND2_X1 U6717 ( .A1(n5556), .A2(n5555), .ZN(n5557) );
  OR2_X1 U6718 ( .A1(n5558), .A2(n5557), .ZN(n5721) );
  NOR2_X1 U6719 ( .A1(n5648), .A2(n6128), .ZN(n5559) );
  AOI21_X1 U6720 ( .B1(n6115), .B2(EBX_REG_27__SCAN_IN), .A(n5559), .ZN(n5560)
         );
  OAI21_X1 U6721 ( .B1(n6120), .B2(n5721), .A(n5560), .ZN(n5561) );
  AOI211_X1 U6722 ( .C1(n5824), .C2(n6606), .A(n5562), .B(n5561), .ZN(n5563)
         );
  OAI21_X1 U6723 ( .B1(n5567), .B2(n5890), .A(n5563), .ZN(U2800) );
  INV_X1 U6724 ( .A(n5564), .ZN(n5566) );
  OAI22_X1 U6725 ( .A1(n5566), .A2(n6150), .B1(n5565), .B2(n6159), .ZN(U2828)
         );
  INV_X1 U6726 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5568) );
  OAI222_X1 U6727 ( .A1(n5568), .A2(n6159), .B1(n6150), .B2(n5721), .C1(n5567), 
        .C2(n5636), .ZN(U2832) );
  NOR2_X1 U6728 ( .A1(n5569), .A2(n5570), .ZN(n5572) );
  AOI21_X1 U6729 ( .B1(n5590), .B2(n5577), .A(n5576), .ZN(n5578) );
  NOR2_X1 U6730 ( .A1(n5579), .A2(n5578), .ZN(n5943) );
  INV_X1 U6731 ( .A(n5943), .ZN(n5580) );
  OAI222_X1 U6732 ( .A1(n5666), .A2(n5601), .B1(n6159), .B2(n5581), .C1(n5580), 
        .C2(n6150), .ZN(U2834) );
  INV_X1 U6733 ( .A(n5910), .ZN(n5582) );
  OAI222_X1 U6734 ( .A1(n6159), .A2(n5583), .B1(n6150), .B2(n5839), .C1(n5636), 
        .C2(n5582), .ZN(U2835) );
  INV_X1 U6735 ( .A(n5584), .ZN(n5585) );
  INV_X1 U6736 ( .A(n5913), .ZN(n5592) );
  AOI21_X1 U6737 ( .B1(n5381), .B2(n5588), .A(n5587), .ZN(n5589) );
  OR2_X1 U6738 ( .A1(n5590), .A2(n5589), .ZN(n5848) );
  OAI222_X1 U6739 ( .A1(n5636), .A2(n5592), .B1(n6159), .B2(n5591), .C1(n5848), 
        .C2(n6150), .ZN(U2836) );
  NOR2_X1 U6740 ( .A1(n5593), .A2(n5594), .ZN(n5595) );
  INV_X1 U6741 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5600) );
  AND2_X1 U6742 ( .A1(n5598), .A2(n5597), .ZN(n5599) );
  OR2_X1 U6743 ( .A1(n5599), .A2(n5381), .ZN(n5869) );
  OAI222_X1 U6744 ( .A1(n5870), .A2(n5601), .B1(n6159), .B2(n5600), .C1(n5869), 
        .C2(n6150), .ZN(U2838) );
  NOR2_X1 U6745 ( .A1(n5611), .A2(n5603), .ZN(n5604) );
  OR2_X1 U6746 ( .A1(n5593), .A2(n5604), .ZN(n5879) );
  NAND2_X1 U6747 ( .A1(n5606), .A2(n5616), .ZN(n5605) );
  OAI21_X1 U6748 ( .B1(n5606), .B2(n5617), .A(n5605), .ZN(n5608) );
  XNOR2_X1 U6749 ( .A(n5608), .B(n5607), .ZN(n5883) );
  INV_X1 U6750 ( .A(EBX_REG_20__SCAN_IN), .ZN(n6930) );
  OAI222_X1 U6751 ( .A1(n5879), .A2(n5636), .B1(n6150), .B2(n5883), .C1(n6159), 
        .C2(n6930), .ZN(U2839) );
  AND2_X1 U6752 ( .A1(n5628), .A2(n5610), .ZN(n5612) );
  OR2_X1 U6753 ( .A1(n5612), .A2(n5611), .ZN(n5922) );
  INV_X1 U6754 ( .A(n5613), .ZN(n5614) );
  NAND2_X1 U6755 ( .A1(n5614), .A2(n5616), .ZN(n5615) );
  OAI21_X1 U6756 ( .B1(n5617), .B2(n5616), .A(n5615), .ZN(n5623) );
  NAND2_X1 U6757 ( .A1(n5623), .A2(n5950), .ZN(n5625) );
  INV_X1 U6758 ( .A(n5618), .ZN(n5619) );
  XNOR2_X1 U6759 ( .A(n5625), .B(n5619), .ZN(n5889) );
  INV_X1 U6760 ( .A(n5889), .ZN(n5621) );
  AOI22_X1 U6761 ( .A1(n6155), .A2(n5621), .B1(n5620), .B2(EBX_REG_19__SCAN_IN), .ZN(n5622) );
  OAI21_X1 U6762 ( .B1(n5922), .B2(n5636), .A(n5622), .ZN(U2840) );
  OR2_X1 U6763 ( .A1(n5950), .A2(n5623), .ZN(n5624) );
  NAND2_X1 U6764 ( .A1(n5625), .A2(n5624), .ZN(n6006) );
  INV_X1 U6765 ( .A(n5628), .ZN(n5629) );
  AOI21_X1 U6766 ( .B1(n5630), .B2(n5937), .A(n5629), .ZN(n6161) );
  INV_X1 U6767 ( .A(n6161), .ZN(n5703) );
  OAI222_X1 U6768 ( .A1(n6006), .A2(n6150), .B1(n6159), .B2(n3723), .C1(n5636), 
        .C2(n5703), .ZN(U2841) );
  OAI21_X1 U6769 ( .B1(n5632), .B2(n5631), .A(n5951), .ZN(n6025) );
  OAI21_X1 U6770 ( .B1(n5634), .B2(n5633), .A(n5935), .ZN(n5705) );
  OAI222_X1 U6771 ( .A1(n6025), .A2(n6150), .B1(n6159), .B2(n3711), .C1(n5636), 
        .C2(n5705), .ZN(U2843) );
  OAI222_X1 U6772 ( .A1(n5637), .A2(n6150), .B1(n6159), .B2(n3704), .C1(n5636), 
        .C2(n5635), .ZN(U2845) );
  INV_X1 U6773 ( .A(DATAI_15_), .ZN(n5641) );
  INV_X1 U6774 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6822) );
  INV_X1 U6775 ( .A(n6157), .ZN(n5638) );
  OAI222_X1 U6776 ( .A1(n5642), .A2(n5641), .B1(n5640), .B2(n6822), .C1(n5639), 
        .C2(n5638), .ZN(U2876) );
  INV_X1 U6777 ( .A(n5643), .ZN(n5644) );
  AOI21_X1 U6778 ( .B1(n5651), .B2(n5664), .A(n5644), .ZN(n5645) );
  XNOR2_X1 U6779 ( .A(n5645), .B(n6940), .ZN(n5725) );
  NAND2_X1 U6780 ( .A1(n6340), .A2(REIP_REG_27__SCAN_IN), .ZN(n5719) );
  INV_X1 U6781 ( .A(n5719), .ZN(n5646) );
  AOI21_X1 U6782 ( .B1(n6288), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5646), 
        .ZN(n5647) );
  OAI21_X1 U6783 ( .B1(n6296), .B2(n5648), .A(n5647), .ZN(n5649) );
  AOI21_X1 U6784 ( .B1(n5904), .B2(n3099), .A(n5649), .ZN(n5650) );
  OAI21_X1 U6785 ( .B1(n5725), .B2(n5984), .A(n5650), .ZN(U2959) );
  NOR2_X1 U6786 ( .A1(n5652), .A2(n5651), .ZN(n5654) );
  XOR2_X1 U6787 ( .A(n5654), .B(n5653), .Z(n5734) );
  INV_X1 U6788 ( .A(n5655), .ZN(n5660) );
  INV_X1 U6789 ( .A(n5656), .ZN(n5658) );
  AND2_X1 U6790 ( .A1(n6340), .A2(REIP_REG_26__SCAN_IN), .ZN(n5731) );
  AOI21_X1 U6791 ( .B1(n6288), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5731), 
        .ZN(n5657) );
  OAI21_X1 U6792 ( .B1(n6296), .B2(n5658), .A(n5657), .ZN(n5659) );
  AOI21_X1 U6793 ( .B1(n5660), .B2(n3099), .A(n5659), .ZN(n5661) );
  OAI21_X1 U6794 ( .B1(n5734), .B2(n5984), .A(n5661), .ZN(U2960) );
  NOR2_X1 U6795 ( .A1(n5663), .A2(n5662), .ZN(n5665) );
  NOR2_X1 U6796 ( .A1(n5665), .A2(n5664), .ZN(n5942) );
  INV_X1 U6797 ( .A(n5830), .ZN(n5668) );
  AOI22_X1 U6798 ( .A1(n6288), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .B1(n6340), 
        .B2(REIP_REG_25__SCAN_IN), .ZN(n5667) );
  OAI21_X1 U6799 ( .B1(n6296), .B2(n5668), .A(n5667), .ZN(n5669) );
  AOI21_X1 U6800 ( .B1(n5907), .B2(n3099), .A(n5669), .ZN(n5670) );
  OAI21_X1 U6801 ( .B1(n5942), .B2(n5984), .A(n5670), .ZN(U2961) );
  NAND4_X1 U6802 ( .A1(n5672), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n5764), .A4(n5671), .ZN(n5673) );
  OAI21_X1 U6803 ( .B1(n5679), .B2(n5674), .A(n5673), .ZN(n5675) );
  XNOR2_X1 U6804 ( .A(n5675), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5741)
         );
  NAND2_X1 U6805 ( .A1(n6340), .A2(REIP_REG_23__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U6806 ( .A1(n6288), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5676)
         );
  OAI211_X1 U6807 ( .C1(n6296), .C2(n5852), .A(n5735), .B(n5676), .ZN(n5677)
         );
  AOI21_X1 U6808 ( .B1(n5913), .B2(n3099), .A(n5677), .ZN(n5678) );
  OAI21_X1 U6809 ( .B1(n5741), .B2(n5984), .A(n5678), .ZN(U2963) );
  OAI21_X1 U6810 ( .B1(n5681), .B2(n5680), .A(n5679), .ZN(n5682) );
  INV_X1 U6811 ( .A(n5682), .ZN(n5756) );
  INV_X1 U6812 ( .A(n5870), .ZN(n5916) );
  AOI22_X1 U6813 ( .A1(n6288), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .B1(n6340), 
        .B2(REIP_REG_21__SCAN_IN), .ZN(n5683) );
  OAI21_X1 U6814 ( .B1(n6296), .B2(n5874), .A(n5683), .ZN(n5684) );
  AOI21_X1 U6815 ( .B1(n5916), .B2(n3099), .A(n5684), .ZN(n5685) );
  OAI21_X1 U6816 ( .B1(n5756), .B2(n5984), .A(n5685), .ZN(U2965) );
  XNOR2_X1 U6817 ( .A(n5687), .B(n5686), .ZN(n5772) );
  NAND2_X1 U6818 ( .A1(n6340), .A2(REIP_REG_20__SCAN_IN), .ZN(n5767) );
  OAI21_X1 U6819 ( .B1(n5699), .B2(n5875), .A(n5767), .ZN(n5689) );
  NOR2_X1 U6820 ( .A1(n5879), .A2(n6266), .ZN(n5688) );
  AOI211_X1 U6821 ( .C1(n5701), .C2(n5880), .A(n5689), .B(n5688), .ZN(n5690)
         );
  OAI21_X1 U6822 ( .B1(n5772), .B2(n5984), .A(n5690), .ZN(U2966) );
  NAND2_X1 U6823 ( .A1(n6340), .A2(REIP_REG_18__SCAN_IN), .ZN(n5785) );
  NOR2_X1 U6824 ( .A1(n5693), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5932)
         );
  NAND2_X1 U6825 ( .A1(n5932), .A2(n5959), .ZN(n5695) );
  NOR2_X1 U6826 ( .A1(n3556), .A2(n5791), .ZN(n5931) );
  NAND3_X1 U6827 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5692), .A3(n5931), .ZN(n5694) );
  OAI21_X1 U6828 ( .B1(n5692), .B2(n5695), .A(n5694), .ZN(n5696) );
  XOR2_X1 U6829 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .B(n5696), .Z(n5787) );
  NAND2_X1 U6830 ( .A1(n6293), .A2(n5787), .ZN(n5697) );
  OAI211_X1 U6831 ( .C1(n5699), .C2(n5698), .A(n5785), .B(n5697), .ZN(n5700)
         );
  AOI21_X1 U6832 ( .B1(n5701), .B2(n6003), .A(n5700), .ZN(n5702) );
  OAI21_X1 U6833 ( .B1(n5703), .B2(n6266), .A(n5702), .ZN(U2968) );
  NOR2_X1 U6834 ( .A1(n5931), .A2(n5932), .ZN(n5704) );
  XOR2_X1 U6835 ( .A(n5704), .B(n5692), .Z(n5799) );
  INV_X1 U6836 ( .A(n5705), .ZN(n6169) );
  NAND2_X1 U6837 ( .A1(n6340), .A2(REIP_REG_16__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U6838 ( .A1(n6288), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5706)
         );
  OAI211_X1 U6839 ( .C1(n6296), .C2(n6021), .A(n5794), .B(n5706), .ZN(n5707)
         );
  AOI21_X1 U6840 ( .B1(n6169), .B2(n3099), .A(n5707), .ZN(n5708) );
  OAI21_X1 U6841 ( .B1(n5799), .B2(n5984), .A(n5708), .ZN(U2970) );
  OR2_X1 U6842 ( .A1(n5709), .A2(n6354), .ZN(n5717) );
  AOI21_X1 U6843 ( .B1(n6342), .B2(n5823), .A(n5710), .ZN(n5716) );
  NAND2_X1 U6844 ( .A1(n5723), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5715) );
  INV_X1 U6845 ( .A(n5711), .ZN(n5713) );
  NAND3_X1 U6846 ( .A1(n5718), .A2(n5713), .A3(n5712), .ZN(n5714) );
  NAND4_X1 U6847 ( .A1(n5717), .A2(n5716), .A3(n5715), .A4(n5714), .ZN(U2990)
         );
  NAND2_X1 U6848 ( .A1(n5718), .A2(n6940), .ZN(n5720) );
  OAI211_X1 U6849 ( .C1(n6378), .C2(n5721), .A(n5720), .B(n5719), .ZN(n5722)
         );
  AOI21_X1 U6850 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5723), .A(n5722), 
        .ZN(n5724) );
  OAI21_X1 U6851 ( .B1(n5725), .B2(n6354), .A(n5724), .ZN(U2991) );
  AOI211_X1 U6852 ( .C1(n5729), .C2(n5728), .A(n5727), .B(n5947), .ZN(n5730)
         );
  AOI211_X1 U6853 ( .C1(n6342), .C2(n4262), .A(n5731), .B(n5730), .ZN(n5733)
         );
  NAND2_X1 U6854 ( .A1(n5941), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5732) );
  OAI211_X1 U6855 ( .C1(n5734), .C2(n6354), .A(n5733), .B(n5732), .ZN(U2992)
         );
  OAI21_X1 U6856 ( .B1(n6378), .B2(n5848), .A(n5735), .ZN(n5738) );
  NOR2_X1 U6857 ( .A1(n5736), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5737)
         );
  AOI211_X1 U6858 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5739), .A(n5738), .B(n5737), .ZN(n5740) );
  OAI21_X1 U6859 ( .B1(n5741), .B2(n6354), .A(n5740), .ZN(U2995) );
  OAI21_X1 U6860 ( .B1(n6378), .B2(n5865), .A(n5742), .ZN(n5743) );
  AOI21_X1 U6861 ( .B1(n5745), .B2(n5744), .A(n5743), .ZN(n5749) );
  INV_X1 U6862 ( .A(n5746), .ZN(n5747) );
  NOR3_X1 U6863 ( .A1(n5948), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n5747), 
        .ZN(n5752) );
  OAI21_X1 U6864 ( .B1(n5752), .B2(n5754), .A(INSTADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n5748) );
  OAI211_X1 U6865 ( .C1(n5750), .C2(n6354), .A(n5749), .B(n5748), .ZN(U2996)
         );
  NAND2_X1 U6866 ( .A1(n6340), .A2(REIP_REG_21__SCAN_IN), .ZN(n5751) );
  OAI21_X1 U6867 ( .B1(n6378), .B2(n5869), .A(n5751), .ZN(n5753) );
  AOI211_X1 U6868 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5754), .A(n5753), .B(n5752), .ZN(n5755) );
  OAI21_X1 U6869 ( .B1(n5756), .B2(n6354), .A(n5755), .ZN(U2997) );
  INV_X1 U6870 ( .A(n5757), .ZN(n5761) );
  AOI21_X1 U6871 ( .B1(n5759), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5758), 
        .ZN(n5760) );
  NOR2_X1 U6872 ( .A1(n5761), .A2(n5760), .ZN(n5960) );
  OAI21_X1 U6873 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n6369), .A(n5960), 
        .ZN(n5783) );
  AOI21_X1 U6874 ( .B1(n5762), .B2(n6331), .A(n5783), .ZN(n5777) );
  INV_X1 U6875 ( .A(n5777), .ZN(n5770) );
  NOR2_X1 U6876 ( .A1(n5948), .A2(n5763), .ZN(n5781) );
  INV_X1 U6877 ( .A(n5764), .ZN(n5766) );
  NAND3_X1 U6878 ( .A1(n5781), .A2(n5766), .A3(n5765), .ZN(n5768) );
  OAI211_X1 U6879 ( .C1(n5883), .C2(n6378), .A(n5768), .B(n5767), .ZN(n5769)
         );
  AOI21_X1 U6880 ( .B1(n5770), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5769), 
        .ZN(n5771) );
  OAI21_X1 U6881 ( .B1(n5772), .B2(n6354), .A(n5771), .ZN(U2998) );
  AOI21_X1 U6882 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5774), .A(n5773), 
        .ZN(n5775) );
  XNOR2_X1 U6883 ( .A(n5775), .B(n3556), .ZN(n5925) );
  NAND2_X1 U6884 ( .A1(n6340), .A2(REIP_REG_19__SCAN_IN), .ZN(n5776) );
  OAI21_X1 U6885 ( .B1(n6378), .B2(n5889), .A(n5776), .ZN(n5779) );
  NOR2_X1 U6886 ( .A1(n5777), .A2(n5780), .ZN(n5778) );
  AOI211_X1 U6887 ( .C1(n5781), .C2(n5780), .A(n5779), .B(n5778), .ZN(n5782)
         );
  OAI21_X1 U6888 ( .B1(n5925), .B2(n6354), .A(n5782), .ZN(U2999) );
  NAND2_X1 U6889 ( .A1(n5783), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5789) );
  OR3_X1 U6890 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5959), .A3(n5948), 
        .ZN(n5784) );
  OAI211_X1 U6891 ( .C1(n6378), .C2(n6006), .A(n5785), .B(n5784), .ZN(n5786)
         );
  AOI21_X1 U6892 ( .B1(n6381), .B2(n5787), .A(n5786), .ZN(n5788) );
  NAND2_X1 U6893 ( .A1(n5789), .A2(n5788), .ZN(U3000) );
  AOI22_X1 U6894 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .B1(n5791), .B2(n5790), .ZN(n5792)
         );
  NAND2_X1 U6895 ( .A1(n5793), .A2(n5792), .ZN(n5795) );
  OAI211_X1 U6896 ( .C1(n6378), .C2(n6025), .A(n5795), .B(n5794), .ZN(n5796)
         );
  AOI21_X1 U6897 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n5797), .A(n5796), 
        .ZN(n5798) );
  OAI21_X1 U6898 ( .B1(n5799), .B2(n6354), .A(n5798), .ZN(U3002) );
  INV_X1 U6899 ( .A(n5800), .ZN(n5807) );
  AOI21_X1 U6900 ( .B1(n5802), .B2(n5801), .A(n6392), .ZN(n5803) );
  AOI21_X1 U6901 ( .B1(n6107), .B2(n5804), .A(n5803), .ZN(n5805) );
  OAI21_X1 U6902 ( .B1(n5807), .B2(n5806), .A(n5805), .ZN(n5808) );
  MUX2_X1 U6903 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n5808), .S(n6386), 
        .Z(U3462) );
  AND2_X1 U6904 ( .A1(DATAO_REG_31__SCAN_IN), .A2(n6980), .ZN(U2892) );
  INV_X1 U6905 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n5810) );
  OAI21_X1 U6906 ( .B1(n5811), .B2(n5810), .A(n5809), .ZN(U2788) );
  AOI21_X1 U6907 ( .B1(n5898), .B2(n6079), .A(n3115), .ZN(n5820) );
  AOI21_X1 U6908 ( .B1(n5815), .B2(n5814), .A(n5813), .ZN(n5818) );
  OAI22_X1 U6909 ( .A1(n4333), .A2(n6105), .B1(n5816), .B2(n6128), .ZN(n5817)
         );
  AOI211_X1 U6910 ( .C1(n6115), .C2(EBX_REG_29__SCAN_IN), .A(n5818), .B(n5817), 
        .ZN(n5819) );
  NAND2_X1 U6911 ( .A1(n5820), .A2(n5819), .ZN(U2798) );
  AOI22_X1 U6912 ( .A1(EBX_REG_28__SCAN_IN), .A2(n6115), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6130), .ZN(n5828) );
  AOI22_X1 U6913 ( .A1(n5822), .A2(n6133), .B1(REIP_REG_28__SCAN_IN), .B2(
        n5821), .ZN(n5827) );
  AOI22_X1 U6914 ( .A1(n5901), .A2(n6079), .B1(n5823), .B2(n6083), .ZN(n5826)
         );
  NAND3_X1 U6915 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5824), .A3(n6816), .ZN(
        n5825) );
  NAND4_X1 U6916 ( .A1(n5828), .A2(n5827), .A3(n5826), .A4(n5825), .ZN(U2799)
         );
  AOI22_X1 U6917 ( .A1(n5907), .A2(n6079), .B1(n6083), .B2(n5943), .ZN(n5836)
         );
  INV_X1 U6918 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6604) );
  AOI22_X1 U6919 ( .A1(n5830), .A2(n6133), .B1(n5829), .B2(n6604), .ZN(n5835)
         );
  AOI22_X1 U6920 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6115), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6130), .ZN(n5834) );
  NAND2_X1 U6921 ( .A1(n5886), .A2(n5831), .ZN(n5846) );
  INV_X1 U6922 ( .A(n5846), .ZN(n5838) );
  NOR2_X1 U6923 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5832), .ZN(n5841) );
  OAI21_X1 U6924 ( .B1(n5838), .B2(n5841), .A(REIP_REG_25__SCAN_IN), .ZN(n5833) );
  NAND4_X1 U6925 ( .A1(n5836), .A2(n5835), .A3(n5834), .A4(n5833), .ZN(U2802)
         );
  AOI22_X1 U6926 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n6130), .B1(n5837), 
        .B2(n6133), .ZN(n5845) );
  AOI22_X1 U6927 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5838), .B1(
        EBX_REG_24__SCAN_IN), .B2(n6115), .ZN(n5844) );
  INV_X1 U6928 ( .A(n5839), .ZN(n5840) );
  INV_X1 U6929 ( .A(n5841), .ZN(n5842) );
  NAND4_X1 U6930 ( .A1(n5845), .A2(n5844), .A3(n5843), .A4(n5842), .ZN(U2803)
         );
  AOI22_X1 U6931 ( .A1(EBX_REG_23__SCAN_IN), .A2(n6115), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6130), .ZN(n5851) );
  AOI21_X1 U6932 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5860), .A(
        REIP_REG_23__SCAN_IN), .ZN(n5847) );
  OAI22_X1 U6933 ( .A1(n6120), .A2(n5848), .B1(n5847), .B2(n5846), .ZN(n5849)
         );
  AOI21_X1 U6934 ( .B1(n5913), .B2(n6079), .A(n5849), .ZN(n5850) );
  OAI211_X1 U6935 ( .C1(n5852), .C2(n6128), .A(n5851), .B(n5850), .ZN(U2804)
         );
  NOR2_X1 U6936 ( .A1(n5854), .A2(n5853), .ZN(n5878) );
  NOR2_X1 U6937 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5855), .ZN(n5868) );
  INV_X1 U6938 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6599) );
  AOI22_X1 U6939 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n6130), .B1(n6133), 
        .B2(n5856), .ZN(n5857) );
  OAI21_X1 U6940 ( .B1(n5858), .B2(n6138), .A(n5857), .ZN(n5859) );
  AOI21_X1 U6941 ( .B1(n5860), .B2(n6599), .A(n5859), .ZN(n5861) );
  OAI21_X1 U6942 ( .B1(n5862), .B2(n5890), .A(n5861), .ZN(n5863) );
  AOI221_X1 U6943 ( .B1(n5878), .B2(REIP_REG_22__SCAN_IN), .C1(n5868), .C2(
        REIP_REG_22__SCAN_IN), .A(n5863), .ZN(n5864) );
  OAI21_X1 U6944 ( .B1(n5865), .B2(n6120), .A(n5864), .ZN(U2805) );
  AOI22_X1 U6945 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n6130), .B1(
        REIP_REG_21__SCAN_IN), .B2(n5878), .ZN(n5866) );
  INV_X1 U6946 ( .A(n5866), .ZN(n5867) );
  AOI211_X1 U6947 ( .C1(n6115), .C2(EBX_REG_21__SCAN_IN), .A(n5868), .B(n5867), 
        .ZN(n5873) );
  OAI22_X1 U6948 ( .A1(n5870), .A2(n5890), .B1(n6120), .B2(n5869), .ZN(n5871)
         );
  INV_X1 U6949 ( .A(n5871), .ZN(n5872) );
  OAI211_X1 U6950 ( .C1(n5874), .C2(n6128), .A(n5873), .B(n5872), .ZN(U2806)
         );
  OAI22_X1 U6951 ( .A1(n6930), .A2(n6138), .B1(n5875), .B2(n6105), .ZN(n5876)
         );
  AOI221_X1 U6952 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5878), .C1(n5877), .C2(
        n5878), .A(n5876), .ZN(n5882) );
  INV_X1 U6953 ( .A(n5879), .ZN(n5919) );
  AOI22_X1 U6954 ( .A1(n5919), .A2(n6079), .B1(n6133), .B2(n5880), .ZN(n5881)
         );
  OAI211_X1 U6955 ( .C1(n5883), .C2(n6120), .A(n5882), .B(n5881), .ZN(U2807)
         );
  OAI21_X1 U6956 ( .B1(REIP_REG_19__SCAN_IN), .B2(REIP_REG_18__SCAN_IN), .A(
        n5884), .ZN(n5887) );
  INV_X1 U6957 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U6958 ( .A1(n5886), .A2(n5885), .ZN(n6008) );
  OAI22_X1 U6959 ( .A1(n6001), .A2(n5887), .B1(n6595), .B2(n6008), .ZN(n5888)
         );
  AOI211_X1 U6960 ( .C1(n6130), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6094), 
        .B(n5888), .ZN(n5893) );
  OAI222_X1 U6961 ( .A1(n5922), .A2(n5890), .B1(n6120), .B2(n5889), .C1(n5930), 
        .C2(n6128), .ZN(n5891) );
  INV_X1 U6962 ( .A(n5891), .ZN(n5892) );
  OAI211_X1 U6963 ( .C1(n6897), .C2(n6138), .A(n5893), .B(n5892), .ZN(U2808)
         );
  AOI22_X1 U6964 ( .A1(n5894), .A2(n6168), .B1(n6167), .B2(DATAI_30_), .ZN(
        n5896) );
  AOI22_X1 U6965 ( .A1(n6171), .A2(DATAI_14_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6170), .ZN(n5895) );
  NAND2_X1 U6966 ( .A1(n5896), .A2(n5895), .ZN(U2861) );
  AOI21_X1 U6967 ( .B1(n5898), .B2(n6168), .A(n5897), .ZN(n5900) );
  AOI22_X1 U6968 ( .A1(n6171), .A2(DATAI_13_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6170), .ZN(n5899) );
  NAND2_X1 U6969 ( .A1(n5900), .A2(n5899), .ZN(U2862) );
  AOI22_X1 U6970 ( .A1(n5901), .A2(n6168), .B1(n6167), .B2(DATAI_28_), .ZN(
        n5903) );
  AOI22_X1 U6971 ( .A1(n6171), .A2(DATAI_12_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6170), .ZN(n5902) );
  NAND2_X1 U6972 ( .A1(n5903), .A2(n5902), .ZN(U2863) );
  AOI22_X1 U6973 ( .A1(n5904), .A2(n6168), .B1(n6167), .B2(DATAI_27_), .ZN(
        n5906) );
  AOI22_X1 U6974 ( .A1(n6171), .A2(DATAI_11_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6170), .ZN(n5905) );
  NAND2_X1 U6975 ( .A1(n5906), .A2(n5905), .ZN(U2864) );
  AOI22_X1 U6976 ( .A1(n5907), .A2(n6168), .B1(n6167), .B2(DATAI_25_), .ZN(
        n5909) );
  AOI22_X1 U6977 ( .A1(n6171), .A2(DATAI_9_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6170), .ZN(n5908) );
  NAND2_X1 U6978 ( .A1(n5909), .A2(n5908), .ZN(U2866) );
  AOI22_X1 U6979 ( .A1(n5910), .A2(n6168), .B1(DATAI_24_), .B2(n6167), .ZN(
        n5912) );
  AOI22_X1 U6980 ( .A1(n6171), .A2(DATAI_8_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6170), .ZN(n5911) );
  NAND2_X1 U6981 ( .A1(n5912), .A2(n5911), .ZN(U2867) );
  AOI22_X1 U6982 ( .A1(n5913), .A2(n6168), .B1(n6167), .B2(DATAI_23_), .ZN(
        n5915) );
  AOI22_X1 U6983 ( .A1(n6171), .A2(DATAI_7_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n6170), .ZN(n5914) );
  NAND2_X1 U6984 ( .A1(n5915), .A2(n5914), .ZN(U2868) );
  AOI22_X1 U6985 ( .A1(n5916), .A2(n6168), .B1(n6167), .B2(DATAI_21_), .ZN(
        n5918) );
  AOI22_X1 U6986 ( .A1(n6171), .A2(DATAI_5_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n6170), .ZN(n5917) );
  NAND2_X1 U6987 ( .A1(n5918), .A2(n5917), .ZN(U2870) );
  AOI22_X1 U6988 ( .A1(n5919), .A2(n6168), .B1(n6167), .B2(DATAI_20_), .ZN(
        n5921) );
  AOI22_X1 U6989 ( .A1(n6171), .A2(DATAI_4_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n6170), .ZN(n5920) );
  NAND2_X1 U6990 ( .A1(n5921), .A2(n5920), .ZN(U2871) );
  INV_X1 U6991 ( .A(n5922), .ZN(n5926) );
  AOI22_X1 U6992 ( .A1(n5926), .A2(n6168), .B1(n6167), .B2(DATAI_19_), .ZN(
        n5924) );
  AOI22_X1 U6993 ( .A1(n6171), .A2(DATAI_3_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n6170), .ZN(n5923) );
  NAND2_X1 U6994 ( .A1(n5924), .A2(n5923), .ZN(U2872) );
  AOI22_X1 U6995 ( .A1(n6340), .A2(REIP_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6288), .ZN(n5929) );
  INV_X1 U6996 ( .A(n5925), .ZN(n5927) );
  AOI22_X1 U6997 ( .A1(n5927), .A2(n6293), .B1(n3099), .B2(n5926), .ZN(n5928)
         );
  OAI211_X1 U6998 ( .C1(n5930), .C2(n6296), .A(n5929), .B(n5928), .ZN(U2967)
         );
  MUX2_X1 U6999 ( .A(n5932), .B(n5931), .S(n5692), .Z(n5933) );
  XNOR2_X1 U7000 ( .A(n5933), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5963)
         );
  AOI22_X1 U7001 ( .A1(n6340), .A2(REIP_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6288), .ZN(n5940) );
  NAND2_X1 U7002 ( .A1(n5935), .A2(n5934), .ZN(n5936) );
  AND2_X1 U7003 ( .A1(n5937), .A2(n5936), .ZN(n6164) );
  NOR2_X1 U7004 ( .A1(n6296), .A2(n6014), .ZN(n5938) );
  AOI21_X1 U7005 ( .B1(n6164), .B2(n3099), .A(n5938), .ZN(n5939) );
  OAI211_X1 U7006 ( .C1(n5963), .C2(n5984), .A(n5940), .B(n5939), .ZN(U2969)
         );
  AOI22_X1 U7007 ( .A1(n6340), .A2(REIP_REG_25__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5941), .ZN(n5946) );
  INV_X1 U7008 ( .A(n5942), .ZN(n5944) );
  AOI22_X1 U7009 ( .A1(n5944), .A2(n6381), .B1(n6342), .B2(n5943), .ZN(n5945)
         );
  OAI211_X1 U7010 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5947), .A(n5946), .B(n5945), .ZN(U2993) );
  INV_X1 U7011 ( .A(n5948), .ZN(n5949) );
  NAND2_X1 U7012 ( .A1(n5949), .A2(n5959), .ZN(n5958) );
  INV_X1 U7013 ( .A(n5950), .ZN(n5954) );
  NAND2_X1 U7014 ( .A1(n5952), .A2(n5951), .ZN(n5953) );
  NAND2_X1 U7015 ( .A1(n5954), .A2(n5953), .ZN(n6149) );
  NAND2_X1 U7016 ( .A1(n6340), .A2(REIP_REG_17__SCAN_IN), .ZN(n5955) );
  OAI21_X1 U7017 ( .B1(n6378), .B2(n6149), .A(n5955), .ZN(n5956) );
  INV_X1 U7018 ( .A(n5956), .ZN(n5957) );
  OAI211_X1 U7019 ( .C1(n5960), .C2(n5959), .A(n5958), .B(n5957), .ZN(n5961)
         );
  INV_X1 U7020 ( .A(n5961), .ZN(n5962) );
  OAI21_X1 U7021 ( .B1(n5963), .B2(n6354), .A(n5962), .ZN(U3001) );
  AOI21_X1 U7022 ( .B1(n6342), .B2(n6035), .A(n5964), .ZN(n5969) );
  NOR2_X1 U7023 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6298), .ZN(n5966)
         );
  INV_X1 U7024 ( .A(n5965), .ZN(n6308) );
  AOI22_X1 U7025 ( .A1(n5967), .A2(n6381), .B1(n5966), .B2(n6308), .ZN(n5968)
         );
  OAI211_X1 U7026 ( .C1(n5970), .C2(n3539), .A(n5969), .B(n5968), .ZN(U3005)
         );
  INV_X1 U7027 ( .A(n6096), .ZN(n5973) );
  INV_X1 U7028 ( .A(n3655), .ZN(n5971) );
  NAND3_X1 U7029 ( .A1(n5973), .A2(n5972), .A3(n5971), .ZN(n5975) );
  OAI22_X1 U7030 ( .A1(n5976), .A2(n5975), .B1(n5974), .B2(n6630), .ZN(U3455)
         );
  AOI21_X1 U7031 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6565), .A(n3634), .ZN(n5982) );
  INV_X1 U7032 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5977) );
  AND2_X1 U7033 ( .A1(n3634), .A2(STATE_REG_1__SCAN_IN), .ZN(n6655) );
  AOI21_X1 U7034 ( .B1(n5982), .B2(n5977), .A(n6655), .ZN(U2789) );
  INV_X1 U7035 ( .A(n5978), .ZN(n5979) );
  OAI21_X1 U7036 ( .B1(n5979), .B2(n6539), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5980) );
  OAI21_X1 U7037 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6538), .A(n5980), .ZN(
        U2790) );
  INV_X2 U7038 ( .A(n6655), .ZN(n6656) );
  NOR2_X1 U7039 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5983) );
  OAI21_X1 U7040 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5983), .A(n6656), .ZN(n5981)
         );
  OAI21_X1 U7041 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6656), .A(n5981), .ZN(
        U2791) );
  NOR2_X1 U7042 ( .A1(n6655), .A2(n5982), .ZN(n6620) );
  OAI21_X1 U7043 ( .B1(BS16_N), .B2(n5983), .A(n6620), .ZN(n6618) );
  OAI21_X1 U7044 ( .B1(n6620), .B2(n6735), .A(n6618), .ZN(U2792) );
  OAI21_X1 U7045 ( .B1(n5985), .B2(n6515), .A(n5984), .ZN(U2793) );
  NOR4_X1 U7046 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_20__SCAN_IN), .ZN(n5989) );
  NOR4_X1 U7047 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_12__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n5988) );
  NOR4_X1 U7048 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5987) );
  NOR4_X1 U7049 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_22__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n5986) );
  NAND4_X1 U7050 ( .A1(n5989), .A2(n5988), .A3(n5987), .A4(n5986), .ZN(n5995)
         );
  NOR4_X1 U7051 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(DATAWIDTH_REG_23__SCAN_IN), .ZN(n5993)
         );
  AOI211_X1 U7052 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_13__SCAN_IN), .B(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n5992) );
  NOR4_X1 U7053 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_9__SCAN_IN), .ZN(
        n5991) );
  NOR4_X1 U7054 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), .A3(DATAWIDTH_REG_4__SCAN_IN), .A4(DATAWIDTH_REG_5__SCAN_IN), .ZN(n5990) );
  NAND4_X1 U7055 ( .A1(n5993), .A2(n5992), .A3(n5991), .A4(n5990), .ZN(n5994)
         );
  NOR2_X1 U7056 ( .A1(n5995), .A2(n5994), .ZN(n6636) );
  INV_X1 U7057 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6927) );
  NOR3_X1 U7058 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5997) );
  OAI21_X1 U7059 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5997), .A(n6636), .ZN(n5996)
         );
  OAI21_X1 U7060 ( .B1(n6636), .B2(n6927), .A(n5996), .ZN(U2794) );
  INV_X1 U7061 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6632) );
  INV_X1 U7062 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6619) );
  AOI21_X1 U7063 ( .B1(n6632), .B2(n6619), .A(n5997), .ZN(n5999) );
  INV_X1 U7064 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5998) );
  INV_X1 U7065 ( .A(n6636), .ZN(n6639) );
  AOI22_X1 U7066 ( .A1(n6636), .A2(n5999), .B1(n5998), .B2(n6639), .ZN(U2795)
         );
  INV_X1 U7067 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6592) );
  AOI21_X1 U7068 ( .B1(n6130), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6094), 
        .ZN(n6000) );
  OAI221_X1 U7069 ( .B1(REIP_REG_18__SCAN_IN), .B2(n6001), .C1(n6592), .C2(
        n6008), .A(n6000), .ZN(n6002) );
  AOI21_X1 U7070 ( .B1(EBX_REG_18__SCAN_IN), .B2(n6115), .A(n6002), .ZN(n6005)
         );
  AOI22_X1 U7071 ( .A1(n6161), .A2(n6079), .B1(n6133), .B2(n6003), .ZN(n6004)
         );
  OAI211_X1 U7072 ( .C1(n6120), .C2(n6006), .A(n6005), .B(n6004), .ZN(U2809)
         );
  INV_X1 U7073 ( .A(n6015), .ZN(n6007) );
  INV_X1 U7074 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6587) );
  NOR2_X1 U7075 ( .A1(n6007), .A2(n6587), .ZN(n6016) );
  AOI21_X1 U7076 ( .B1(REIP_REG_16__SCAN_IN), .B2(n6016), .A(
        REIP_REG_17__SCAN_IN), .ZN(n6009) );
  INV_X1 U7077 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6153) );
  OAI22_X1 U7078 ( .A1(n6009), .A2(n6008), .B1(n6153), .B2(n6138), .ZN(n6010)
         );
  AOI211_X1 U7079 ( .C1(n6130), .C2(PHYADDRPOINTER_REG_17__SCAN_IN), .A(n6094), 
        .B(n6010), .ZN(n6013) );
  INV_X1 U7080 ( .A(n6149), .ZN(n6011) );
  AOI22_X1 U7081 ( .A1(n6164), .A2(n6079), .B1(n6083), .B2(n6011), .ZN(n6012)
         );
  OAI211_X1 U7082 ( .C1(n6014), .C2(n6128), .A(n6013), .B(n6012), .ZN(U2810)
         );
  INV_X1 U7084 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6590) );
  AND2_X1 U7085 ( .A1(n6015), .A2(n6587), .ZN(n6027) );
  OAI33_X1 U7086 ( .A1(1'b0), .A2(n6016), .A3(REIP_REG_16__SCAN_IN), .B1(n6590), .B2(n6026), .B3(n6027), .ZN(n6018) );
  OAI211_X1 U7087 ( .C1(n6105), .C2(n6019), .A(n6018), .B(n6085), .ZN(n6020)
         );
  AOI21_X1 U7088 ( .B1(EBX_REG_16__SCAN_IN), .B2(n6115), .A(n6020), .ZN(n6024)
         );
  INV_X1 U7089 ( .A(n6021), .ZN(n6022) );
  AOI22_X1 U7090 ( .A1(n6169), .A2(n6079), .B1(n6022), .B2(n6133), .ZN(n6023)
         );
  OAI211_X1 U7091 ( .C1(n6120), .C2(n6025), .A(n6024), .B(n6023), .ZN(U2811)
         );
  AOI22_X1 U7092 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6115), .B1(
        REIP_REG_15__SCAN_IN), .B2(n6026), .ZN(n6029) );
  AOI211_X1 U7093 ( .C1(n6130), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6094), 
        .B(n6027), .ZN(n6028) );
  NAND2_X1 U7094 ( .A1(n6029), .A2(n6028), .ZN(n6030) );
  AOI21_X1 U7095 ( .B1(n6157), .B2(n6079), .A(n6030), .ZN(n6033) );
  AOI22_X1 U7096 ( .A1(n6031), .A2(n6133), .B1(n6083), .B2(n6154), .ZN(n6032)
         );
  NAND2_X1 U7097 ( .A1(n6033), .A2(n6032), .ZN(U2812) );
  OAI21_X1 U7098 ( .B1(REIP_REG_13__SCAN_IN), .B2(REIP_REG_12__SCAN_IN), .A(
        n6034), .ZN(n6045) );
  AOI22_X1 U7099 ( .A1(n6083), .A2(n6035), .B1(REIP_REG_13__SCAN_IN), .B2(
        n6046), .ZN(n6036) );
  OAI211_X1 U7100 ( .C1(n6105), .C2(n6037), .A(n6036), .B(n6085), .ZN(n6038)
         );
  AOI21_X1 U7101 ( .B1(EBX_REG_13__SCAN_IN), .B2(n6115), .A(n6038), .ZN(n6044)
         );
  INV_X1 U7102 ( .A(n6039), .ZN(n6042) );
  INV_X1 U7103 ( .A(n6040), .ZN(n6041) );
  AOI22_X1 U7104 ( .A1(n6042), .A2(n6079), .B1(n6133), .B2(n6041), .ZN(n6043)
         );
  OAI211_X1 U7105 ( .C1(n6054), .C2(n6045), .A(n6044), .B(n6043), .ZN(U2814)
         );
  AOI22_X1 U7106 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6115), .B1(
        REIP_REG_12__SCAN_IN), .B2(n6046), .ZN(n6047) );
  OAI21_X1 U7107 ( .B1(n6120), .B2(n6300), .A(n6047), .ZN(n6048) );
  AOI211_X1 U7108 ( .C1(n6130), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6094), 
        .B(n6048), .ZN(n6053) );
  INV_X1 U7109 ( .A(n6049), .ZN(n6051) );
  AOI22_X1 U7110 ( .A1(n6051), .A2(n6079), .B1(n6050), .B2(n6133), .ZN(n6052)
         );
  OAI211_X1 U7111 ( .C1(REIP_REG_12__SCAN_IN), .C2(n6054), .A(n6053), .B(n6052), .ZN(U2815) );
  NAND2_X1 U7112 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6579), .ZN(n6063) );
  AOI22_X1 U7113 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6115), .B1(n6055), .B2(n6133), .ZN(n6056) );
  OAI21_X1 U7114 ( .B1(n6120), .B2(n6057), .A(n6056), .ZN(n6058) );
  AOI211_X1 U7115 ( .C1(n6130), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6094), 
        .B(n6058), .ZN(n6062) );
  AOI22_X1 U7116 ( .A1(n6060), .A2(REIP_REG_10__SCAN_IN), .B1(n6079), .B2(
        n6059), .ZN(n6061) );
  OAI211_X1 U7117 ( .C1(n6064), .C2(n6063), .A(n6062), .B(n6061), .ZN(U2817)
         );
  AOI21_X1 U7118 ( .B1(REIP_REG_7__SCAN_IN), .B2(n6078), .A(
        REIP_REG_8__SCAN_IN), .ZN(n6072) );
  OAI22_X1 U7119 ( .A1(n6066), .A2(n6138), .B1(n6120), .B2(n6065), .ZN(n6067)
         );
  AOI211_X1 U7120 ( .C1(n6130), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6094), 
        .B(n6067), .ZN(n6071) );
  AOI22_X1 U7121 ( .A1(n6069), .A2(n6079), .B1(n6133), .B2(n6068), .ZN(n6070)
         );
  OAI211_X1 U7122 ( .C1(n6073), .C2(n6072), .A(n6071), .B(n6070), .ZN(U2819)
         );
  INV_X1 U7123 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6576) );
  OAI21_X1 U7124 ( .B1(REIP_REG_6__SCAN_IN), .B2(n6074), .A(n6087), .ZN(n6077)
         );
  INV_X1 U7125 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6755) );
  AOI22_X1 U7126 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6115), .B1(n6083), .B2(n6322), 
        .ZN(n6075) );
  OAI211_X1 U7127 ( .C1(n6105), .C2(n6755), .A(n6075), .B(n6085), .ZN(n6076)
         );
  AOI221_X1 U7128 ( .B1(n6078), .B2(n6576), .C1(n6077), .C2(
        REIP_REG_7__SCAN_IN), .A(n6076), .ZN(n6082) );
  INV_X1 U7129 ( .A(n6267), .ZN(n6080) );
  NAND2_X1 U7130 ( .A1(n6080), .A2(n6079), .ZN(n6081) );
  OAI211_X1 U7131 ( .C1(n6128), .C2(n6271), .A(n6082), .B(n6081), .ZN(U2820)
         );
  INV_X1 U7132 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6885) );
  AOI22_X1 U7133 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6115), .B1(n6083), .B2(n6341), 
        .ZN(n6084) );
  OAI211_X1 U7134 ( .C1(n6105), .C2(n6885), .A(n6085), .B(n6084), .ZN(n6086)
         );
  AOI21_X1 U7135 ( .B1(n6276), .B2(n6126), .A(n6086), .ZN(n6091) );
  INV_X1 U7136 ( .A(n6087), .ZN(n6088) );
  OAI21_X1 U7137 ( .B1(REIP_REG_5__SCAN_IN), .B2(n6089), .A(n6088), .ZN(n6090)
         );
  OAI211_X1 U7138 ( .C1(n6128), .C2(n6279), .A(n6091), .B(n6090), .ZN(U2822)
         );
  INV_X1 U7139 ( .A(n6092), .ZN(n6093) );
  OAI21_X1 U7140 ( .B1(n6110), .B2(n6093), .A(n6148), .ZN(n6112) );
  AOI221_X1 U7141 ( .B1(n6095), .B2(n6725), .C1(n6112), .C2(
        REIP_REG_4__SCAN_IN), .A(n6094), .ZN(n6102) );
  OAI22_X1 U7142 ( .A1(n6120), .A2(n6356), .B1(n6096), .B2(n6137), .ZN(n6100)
         );
  OAI22_X1 U7143 ( .A1(n6098), .A2(n6143), .B1(n6097), .B2(n6128), .ZN(n6099)
         );
  AOI211_X1 U7144 ( .C1(EBX_REG_4__SCAN_IN), .C2(n6115), .A(n6100), .B(n6099), 
        .ZN(n6101) );
  OAI211_X1 U7145 ( .C1(n6103), .C2(n6105), .A(n6102), .B(n6101), .ZN(U2823)
         );
  INV_X1 U7146 ( .A(n6137), .ZN(n6117) );
  INV_X1 U7147 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6104) );
  INV_X1 U7148 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6963) );
  OAI22_X1 U7149 ( .A1(n6105), .A2(n6104), .B1(n6138), .B2(n6963), .ZN(n6106)
         );
  AOI21_X1 U7150 ( .B1(n6117), .B2(n6107), .A(n6106), .ZN(n6108) );
  OAI21_X1 U7151 ( .B1(n6362), .B2(n6120), .A(n6108), .ZN(n6109) );
  AOI21_X1 U7152 ( .B1(n6284), .B2(n6126), .A(n6109), .ZN(n6114) );
  NOR2_X1 U7153 ( .A1(n6110), .A2(REIP_REG_1__SCAN_IN), .ZN(n6129) );
  INV_X1 U7154 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6955) );
  NOR3_X1 U7155 ( .A1(n6129), .A2(n6111), .A3(n6955), .ZN(n6123) );
  OAI21_X1 U7156 ( .B1(REIP_REG_3__SCAN_IN), .B2(n6123), .A(n6112), .ZN(n6113)
         );
  OAI211_X1 U7157 ( .C1(n6128), .C2(n6287), .A(n6114), .B(n6113), .ZN(U2824)
         );
  AOI22_X1 U7158 ( .A1(n6115), .A2(EBX_REG_2__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n6130), .ZN(n6119) );
  NAND2_X1 U7159 ( .A1(n6117), .A2(n6116), .ZN(n6118) );
  OAI211_X1 U7160 ( .C1(n6120), .C2(n6377), .A(n6119), .B(n6118), .ZN(n6125)
         );
  AOI21_X1 U7161 ( .B1(n6121), .B2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .ZN(n6122) );
  NOR2_X1 U7162 ( .A1(n6123), .A2(n6122), .ZN(n6124) );
  AOI211_X1 U7163 ( .C1(n6292), .C2(n6126), .A(n6125), .B(n6124), .ZN(n6127)
         );
  OAI21_X1 U7164 ( .B1(n6297), .B2(n6128), .A(n6127), .ZN(U2825) );
  AOI21_X1 U7165 ( .B1(n6130), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n6129), 
        .ZN(n6147) );
  INV_X1 U7166 ( .A(n6131), .ZN(n6135) );
  INV_X1 U7167 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6132) );
  AOI22_X1 U7168 ( .A1(n6135), .A2(n6134), .B1(n6133), .B2(n6132), .ZN(n6142)
         );
  OAI22_X1 U7169 ( .A1(n6139), .A2(n6138), .B1(n6137), .B2(n6136), .ZN(n6140)
         );
  INV_X1 U7170 ( .A(n6140), .ZN(n6141) );
  OAI211_X1 U7171 ( .C1(n6144), .C2(n6143), .A(n6142), .B(n6141), .ZN(n6145)
         );
  INV_X1 U7172 ( .A(n6145), .ZN(n6146) );
  OAI211_X1 U7173 ( .C1(n6148), .C2(n6632), .A(n6147), .B(n6146), .ZN(U2826)
         );
  NOR2_X1 U7174 ( .A1(n6150), .A2(n6149), .ZN(n6151) );
  AOI21_X1 U7175 ( .B1(n6164), .B2(n6156), .A(n6151), .ZN(n6152) );
  OAI21_X1 U7176 ( .B1(n6153), .B2(n6159), .A(n6152), .ZN(U2842) );
  AOI22_X1 U7177 ( .A1(n6157), .A2(n6156), .B1(n6155), .B2(n6154), .ZN(n6158)
         );
  OAI21_X1 U7178 ( .B1(n6160), .B2(n6159), .A(n6158), .ZN(U2844) );
  AOI22_X1 U7179 ( .A1(n6161), .A2(n6168), .B1(n6167), .B2(DATAI_18_), .ZN(
        n6163) );
  AOI22_X1 U7180 ( .A1(n6171), .A2(DATAI_2_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n6170), .ZN(n6162) );
  NAND2_X1 U7181 ( .A1(n6163), .A2(n6162), .ZN(U2873) );
  AOI22_X1 U7182 ( .A1(n6164), .A2(n6168), .B1(n6167), .B2(DATAI_17_), .ZN(
        n6166) );
  AOI22_X1 U7183 ( .A1(n6171), .A2(DATAI_1_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n6170), .ZN(n6165) );
  NAND2_X1 U7184 ( .A1(n6166), .A2(n6165), .ZN(U2874) );
  AOI22_X1 U7185 ( .A1(n6169), .A2(n6168), .B1(n6167), .B2(DATAI_16_), .ZN(
        n6173) );
  AOI22_X1 U7186 ( .A1(n6171), .A2(DATAI_0_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n6170), .ZN(n6172) );
  NAND2_X1 U7187 ( .A1(n6173), .A2(n6172), .ZN(U2875) );
  INV_X1 U7188 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n6873) );
  AOI22_X1 U7189 ( .A1(EAX_REG_15__SCAN_IN), .A2(n6981), .B1(n6194), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n6174) );
  OAI21_X1 U7190 ( .B1(n6873), .B2(n6175), .A(n6174), .ZN(U2908) );
  INV_X1 U7191 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6257) );
  AOI22_X1 U7192 ( .A1(LWORD_REG_14__SCAN_IN), .A2(n6194), .B1(n6980), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6176) );
  OAI21_X1 U7193 ( .B1(n6257), .B2(n6196), .A(n6176), .ZN(U2909) );
  AOI22_X1 U7194 ( .A1(n6194), .A2(LWORD_REG_13__SCAN_IN), .B1(n6980), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6177) );
  OAI21_X1 U7195 ( .B1(n6178), .B2(n6196), .A(n6177), .ZN(U2910) );
  AOI22_X1 U7196 ( .A1(n6194), .A2(LWORD_REG_12__SCAN_IN), .B1(n6980), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6179) );
  OAI21_X1 U7197 ( .B1(n3950), .B2(n6196), .A(n6179), .ZN(U2911) );
  INV_X1 U7198 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6248) );
  AOI22_X1 U7199 ( .A1(n6194), .A2(LWORD_REG_11__SCAN_IN), .B1(n6980), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6180) );
  OAI21_X1 U7200 ( .B1(n6248), .B2(n6196), .A(n6180), .ZN(U2912) );
  INV_X1 U7201 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6245) );
  AOI22_X1 U7202 ( .A1(n6194), .A2(LWORD_REG_10__SCAN_IN), .B1(n6980), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6181) );
  OAI21_X1 U7203 ( .B1(n6245), .B2(n6196), .A(n6181), .ZN(U2913) );
  INV_X1 U7204 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6242) );
  AOI22_X1 U7205 ( .A1(n6194), .A2(LWORD_REG_9__SCAN_IN), .B1(n6980), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6182) );
  OAI21_X1 U7206 ( .B1(n6242), .B2(n6196), .A(n6182), .ZN(U2914) );
  INV_X1 U7207 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6819) );
  AOI22_X1 U7208 ( .A1(DATAO_REG_8__SCAN_IN), .A2(n6980), .B1(n6194), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n6183) );
  OAI21_X1 U7209 ( .B1(n6819), .B2(n6196), .A(n6183), .ZN(U2915) );
  AOI22_X1 U7210 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n6194), .B1(n6980), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6184) );
  OAI21_X1 U7211 ( .B1(n6185), .B2(n6196), .A(n6184), .ZN(U2916) );
  AOI22_X1 U7212 ( .A1(DATAO_REG_6__SCAN_IN), .A2(n6980), .B1(n6194), .B2(
        LWORD_REG_6__SCAN_IN), .ZN(n6186) );
  OAI21_X1 U7213 ( .B1(n6866), .B2(n6196), .A(n6186), .ZN(U2917) );
  AOI22_X1 U7214 ( .A1(n6194), .A2(LWORD_REG_5__SCAN_IN), .B1(n6980), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6187) );
  OAI21_X1 U7215 ( .B1(n3872), .B2(n6196), .A(n6187), .ZN(U2918) );
  AOI22_X1 U7216 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n6194), .B1(n6980), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6188) );
  OAI21_X1 U7217 ( .B1(n6189), .B2(n6196), .A(n6188), .ZN(U2919) );
  AOI22_X1 U7218 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n6194), .B1(n6980), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6190) );
  OAI21_X1 U7219 ( .B1(n6191), .B2(n6196), .A(n6190), .ZN(U2920) );
  AOI22_X1 U7220 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n6194), .B1(n6980), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6192) );
  OAI21_X1 U7221 ( .B1(n6193), .B2(n6196), .A(n6192), .ZN(U2922) );
  AOI22_X1 U7222 ( .A1(n6194), .A2(LWORD_REG_0__SCAN_IN), .B1(n6980), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6195) );
  OAI21_X1 U7223 ( .B1(n6197), .B2(n6196), .A(n6195), .ZN(U2923) );
  INV_X1 U7224 ( .A(n6198), .ZN(n6199) );
  OAI21_X1 U7225 ( .B1(n6648), .B2(n3646), .A(n6199), .ZN(n6254) );
  AOI22_X1 U7226 ( .A1(n6259), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n6258), .ZN(n6200) );
  OAI21_X1 U7227 ( .B1(n6261), .B2(n6227), .A(n6200), .ZN(U2924) );
  AOI22_X1 U7228 ( .A1(n6259), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n6258), .ZN(n6201) );
  OAI21_X1 U7229 ( .B1(n6261), .B2(n6751), .A(n6201), .ZN(U2925) );
  AOI22_X1 U7230 ( .A1(n6259), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6258), .ZN(n6202) );
  OAI21_X1 U7231 ( .B1(n6261), .B2(n6888), .A(n6202), .ZN(U2926) );
  AOI22_X1 U7232 ( .A1(n6259), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6258), .ZN(n6203) );
  OAI21_X1 U7233 ( .B1(n6261), .B2(n6231), .A(n6203), .ZN(U2927) );
  AOI22_X1 U7234 ( .A1(n6259), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n6258), .ZN(n6204) );
  OAI21_X1 U7235 ( .B1(n6261), .B2(n6805), .A(n6204), .ZN(U2928) );
  AOI22_X1 U7236 ( .A1(n6259), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6258), .ZN(n6205) );
  OAI21_X1 U7237 ( .B1(n6261), .B2(n6234), .A(n6205), .ZN(U2929) );
  AOI22_X1 U7238 ( .A1(n6259), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6258), .ZN(n6206) );
  OAI21_X1 U7239 ( .B1(n6261), .B2(n6728), .A(n6206), .ZN(U2930) );
  AOI22_X1 U7240 ( .A1(n6259), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6258), .ZN(n6207) );
  OAI21_X1 U7241 ( .B1(n6261), .B2(n6237), .A(n6207), .ZN(U2931) );
  INV_X1 U7242 ( .A(DATAI_8_), .ZN(n6208) );
  NOR2_X1 U7243 ( .A1(n6261), .A2(n6208), .ZN(n6238) );
  AOI21_X1 U7244 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n6254), .A(n6238), .ZN(n6209) );
  OAI21_X1 U7245 ( .B1(n6210), .B2(n6256), .A(n6209), .ZN(U2932) );
  INV_X1 U7246 ( .A(DATAI_9_), .ZN(n6211) );
  NOR2_X1 U7247 ( .A1(n6261), .A2(n6211), .ZN(n6240) );
  AOI21_X1 U7248 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6259), .A(n6240), .ZN(n6212) );
  OAI21_X1 U7249 ( .B1(n6213), .B2(n6256), .A(n6212), .ZN(U2933) );
  INV_X1 U7250 ( .A(DATAI_10_), .ZN(n6214) );
  NOR2_X1 U7251 ( .A1(n6261), .A2(n6214), .ZN(n6243) );
  AOI21_X1 U7252 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n6259), .A(n6243), .ZN(
        n6215) );
  OAI21_X1 U7253 ( .B1(n6792), .B2(n6256), .A(n6215), .ZN(U2934) );
  INV_X1 U7254 ( .A(DATAI_11_), .ZN(n6216) );
  NOR2_X1 U7255 ( .A1(n6261), .A2(n6216), .ZN(n6246) );
  AOI21_X1 U7256 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n6259), .A(n6246), .ZN(
        n6217) );
  OAI21_X1 U7257 ( .B1(n6218), .B2(n6256), .A(n6217), .ZN(U2935) );
  NOR2_X1 U7258 ( .A1(n6261), .A2(n6219), .ZN(n6249) );
  AOI21_X1 U7259 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6259), .A(n6249), .ZN(
        n6220) );
  OAI21_X1 U7260 ( .B1(n6221), .B2(n6256), .A(n6220), .ZN(U2936) );
  AOI22_X1 U7261 ( .A1(n6259), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n6258), .ZN(n6222) );
  OAI21_X1 U7262 ( .B1(n6261), .B2(n6252), .A(n6222), .ZN(U2937) );
  INV_X1 U7263 ( .A(DATAI_14_), .ZN(n6223) );
  NOR2_X1 U7264 ( .A1(n6261), .A2(n6223), .ZN(n6253) );
  AOI21_X1 U7265 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6259), .A(n6253), .ZN(
        n6224) );
  OAI21_X1 U7266 ( .B1(n6225), .B2(n6256), .A(n6224), .ZN(U2938) );
  AOI22_X1 U7267 ( .A1(n6259), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n6258), .ZN(n6226) );
  OAI21_X1 U7268 ( .B1(n6261), .B2(n6227), .A(n6226), .ZN(U2939) );
  AOI22_X1 U7269 ( .A1(n6259), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6258), .ZN(n6228) );
  OAI21_X1 U7270 ( .B1(n6261), .B2(n6751), .A(n6228), .ZN(U2940) );
  AOI22_X1 U7271 ( .A1(n6259), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6258), .ZN(n6229) );
  OAI21_X1 U7272 ( .B1(n6261), .B2(n6888), .A(n6229), .ZN(U2941) );
  AOI22_X1 U7273 ( .A1(n6259), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6258), .ZN(n6230) );
  OAI21_X1 U7274 ( .B1(n6261), .B2(n6231), .A(n6230), .ZN(U2942) );
  AOI22_X1 U7275 ( .A1(n6259), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6258), .ZN(n6232) );
  OAI21_X1 U7276 ( .B1(n6261), .B2(n6805), .A(n6232), .ZN(U2943) );
  AOI22_X1 U7277 ( .A1(n6259), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6258), .ZN(n6233) );
  OAI21_X1 U7278 ( .B1(n6261), .B2(n6234), .A(n6233), .ZN(U2944) );
  AOI22_X1 U7279 ( .A1(n6259), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6258), .ZN(n6235) );
  OAI21_X1 U7280 ( .B1(n6261), .B2(n6728), .A(n6235), .ZN(U2945) );
  AOI22_X1 U7281 ( .A1(n6259), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6258), .ZN(n6236) );
  OAI21_X1 U7282 ( .B1(n6261), .B2(n6237), .A(n6236), .ZN(U2946) );
  AOI21_X1 U7283 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n6259), .A(n6238), .ZN(n6239) );
  OAI21_X1 U7284 ( .B1(n6819), .B2(n6256), .A(n6239), .ZN(U2947) );
  AOI21_X1 U7285 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n6254), .A(n6240), .ZN(n6241) );
  OAI21_X1 U7286 ( .B1(n6242), .B2(n6256), .A(n6241), .ZN(U2948) );
  AOI21_X1 U7287 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6254), .A(n6243), .ZN(
        n6244) );
  OAI21_X1 U7288 ( .B1(n6245), .B2(n6256), .A(n6244), .ZN(U2949) );
  AOI21_X1 U7289 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n6254), .A(n6246), .ZN(
        n6247) );
  OAI21_X1 U7290 ( .B1(n6248), .B2(n6256), .A(n6247), .ZN(U2950) );
  AOI21_X1 U7291 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n6254), .A(n6249), .ZN(
        n6250) );
  OAI21_X1 U7292 ( .B1(n3950), .B2(n6256), .A(n6250), .ZN(U2951) );
  AOI22_X1 U7293 ( .A1(n6259), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n6258), .ZN(n6251) );
  OAI21_X1 U7294 ( .B1(n6261), .B2(n6252), .A(n6251), .ZN(U2952) );
  AOI21_X1 U7295 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6254), .A(n6253), .ZN(
        n6255) );
  OAI21_X1 U7296 ( .B1(n6257), .B2(n6256), .A(n6255), .ZN(U2953) );
  AOI22_X1 U7297 ( .A1(n6259), .A2(LWORD_REG_15__SCAN_IN), .B1(
        EAX_REG_15__SCAN_IN), .B2(n6258), .ZN(n6260) );
  OAI21_X1 U7298 ( .B1(n6261), .B2(n5641), .A(n6260), .ZN(U2954) );
  AOI22_X1 U7299 ( .A1(n6340), .A2(REIP_REG_7__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n6288), .ZN(n6270) );
  OR2_X1 U7300 ( .A1(n6263), .A2(n6262), .ZN(n6264) );
  AND2_X1 U7301 ( .A1(n6265), .A2(n6264), .ZN(n6323) );
  NOR2_X1 U7302 ( .A1(n6267), .A2(n6266), .ZN(n6268) );
  AOI21_X1 U7303 ( .B1(n6323), .B2(n6293), .A(n6268), .ZN(n6269) );
  OAI211_X1 U7304 ( .C1(n6271), .C2(n6296), .A(n6270), .B(n6269), .ZN(U2979)
         );
  AOI22_X1 U7305 ( .A1(n6340), .A2(REIP_REG_5__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n6288), .ZN(n6278) );
  OAI21_X1 U7306 ( .B1(n6274), .B2(n6273), .A(n6272), .ZN(n6275) );
  INV_X1 U7307 ( .A(n6275), .ZN(n6346) );
  AOI22_X1 U7308 ( .A1(n6346), .A2(n6293), .B1(n3099), .B2(n6276), .ZN(n6277)
         );
  OAI211_X1 U7309 ( .C1(n6279), .C2(n6296), .A(n6278), .B(n6277), .ZN(U2981)
         );
  AOI22_X1 U7310 ( .A1(n6340), .A2(REIP_REG_3__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n6288), .ZN(n6286) );
  INV_X1 U7311 ( .A(n6280), .ZN(n6281) );
  AOI21_X1 U7312 ( .B1(n6283), .B2(n6282), .A(n6281), .ZN(n6364) );
  AOI22_X1 U7313 ( .A1(n6364), .A2(n6293), .B1(n6284), .B2(n3099), .ZN(n6285)
         );
  OAI211_X1 U7314 ( .C1(n6287), .C2(n6296), .A(n6286), .B(n6285), .ZN(U2983)
         );
  AOI22_X1 U7315 ( .A1(n6340), .A2(REIP_REG_2__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n6288), .ZN(n6295) );
  XOR2_X1 U7316 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .B(n6289), .Z(n6290) );
  XNOR2_X1 U7317 ( .A(n6291), .B(n6290), .ZN(n6382) );
  AOI22_X1 U7318 ( .A1(n6382), .A2(n6293), .B1(n3099), .B2(n6292), .ZN(n6294)
         );
  OAI211_X1 U7319 ( .C1(n6297), .C2(n6296), .A(n6295), .B(n6294), .ZN(U2984)
         );
  AOI21_X1 U7320 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6308), .A(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6305) );
  OAI21_X1 U7321 ( .B1(n6375), .B2(n6299), .A(n6298), .ZN(n6304) );
  OAI22_X1 U7322 ( .A1(n6301), .A2(n6354), .B1(n6378), .B2(n6300), .ZN(n6302)
         );
  AOI21_X1 U7323 ( .B1(n6340), .B2(REIP_REG_12__SCAN_IN), .A(n6302), .ZN(n6303) );
  OAI221_X1 U7324 ( .B1(n6305), .B2(n6313), .C1(n6305), .C2(n6304), .A(n6303), 
        .ZN(U3006) );
  AOI21_X1 U7325 ( .B1(n6342), .B2(n6307), .A(n6306), .ZN(n6311) );
  AOI22_X1 U7326 ( .A1(n6381), .A2(n6309), .B1(n6312), .B2(n6308), .ZN(n6310)
         );
  OAI211_X1 U7327 ( .C1(n6313), .C2(n6312), .A(n6311), .B(n6310), .ZN(U3007)
         );
  INV_X1 U7328 ( .A(n6314), .ZN(n6315) );
  AOI21_X1 U7329 ( .B1(n6342), .B2(n6316), .A(n6315), .ZN(n6320) );
  AOI22_X1 U7330 ( .A1(n6318), .A2(n6801), .B1(n6381), .B2(n6317), .ZN(n6319)
         );
  OAI211_X1 U7331 ( .C1(n6321), .C2(n6801), .A(n6320), .B(n6319), .ZN(U3009)
         );
  AOI22_X1 U7332 ( .A1(n6342), .A2(n6322), .B1(n6340), .B2(REIP_REG_7__SCAN_IN), .ZN(n6327) );
  AOI22_X1 U7333 ( .A1(n6324), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .B1(n6381), 
        .B2(n6323), .ZN(n6326) );
  NAND3_X1 U7334 ( .A1(n6327), .A2(n6326), .A3(n6325), .ZN(U3011) );
  AOI22_X1 U7335 ( .A1(n6330), .A2(n6373), .B1(n6329), .B2(n6328), .ZN(n6384)
         );
  INV_X1 U7336 ( .A(n6384), .ZN(n6351) );
  AOI21_X1 U7337 ( .B1(n6332), .B2(n6331), .A(n6351), .ZN(n6350) );
  AOI21_X1 U7338 ( .B1(n6342), .B2(n6334), .A(n6333), .ZN(n6338) );
  AOI22_X1 U7339 ( .A1(n6336), .A2(n6752), .B1(n6335), .B2(n6381), .ZN(n6337)
         );
  OAI211_X1 U7340 ( .C1(n6350), .C2(n6752), .A(n6338), .B(n6337), .ZN(U3012)
         );
  AOI21_X1 U7341 ( .B1(n6375), .B2(n6339), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6349) );
  AOI22_X1 U7342 ( .A1(n6342), .A2(n6341), .B1(n6340), .B2(REIP_REG_5__SCAN_IN), .ZN(n6348) );
  NOR2_X1 U7343 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6343), .ZN(n6344)
         );
  AOI22_X1 U7344 ( .A1(n6346), .A2(n6381), .B1(n6345), .B2(n6344), .ZN(n6347)
         );
  OAI211_X1 U7345 ( .C1(n6350), .C2(n6349), .A(n6348), .B(n6347), .ZN(U3013)
         );
  AOI21_X1 U7346 ( .B1(n6375), .B2(n6352), .A(n6351), .ZN(n6366) );
  AOI211_X1 U7347 ( .C1(n6367), .C2(n6361), .A(n6353), .B(n6368), .ZN(n6359)
         );
  NOR2_X1 U7348 ( .A1(n6355), .A2(n6354), .ZN(n6358) );
  OAI22_X1 U7349 ( .A1(n6378), .A2(n6356), .B1(n6725), .B2(n6376), .ZN(n6357)
         );
  NOR3_X1 U7350 ( .A1(n6359), .A2(n6358), .A3(n6357), .ZN(n6360) );
  OAI21_X1 U7351 ( .B1(n6366), .B2(n6361), .A(n6360), .ZN(U3014) );
  INV_X1 U7352 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6569) );
  OAI22_X1 U7353 ( .A1(n6378), .A2(n6362), .B1(n6569), .B2(n6376), .ZN(n6363)
         );
  AOI21_X1 U7354 ( .B1(n6364), .B2(n6381), .A(n6363), .ZN(n6365) );
  OAI221_X1 U7355 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n6368), .C1(n6367), .C2(n6366), .A(n6365), .ZN(U3015) );
  INV_X1 U7356 ( .A(n6369), .ZN(n6370) );
  NAND2_X1 U7357 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6370), .ZN(n6385)
         );
  OAI21_X1 U7358 ( .B1(n6373), .B2(n6372), .A(n6371), .ZN(n6374) );
  AND2_X1 U7359 ( .A1(n6375), .A2(n6374), .ZN(n6380) );
  OAI22_X1 U7360 ( .A1(n6378), .A2(n6377), .B1(n6955), .B2(n6376), .ZN(n6379)
         );
  AOI211_X1 U7361 ( .C1(n6382), .C2(n6381), .A(n6380), .B(n6379), .ZN(n6383)
         );
  OAI221_X1 U7362 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6385), .C1(n3477), .C2(n6384), .A(n6383), .ZN(U3016) );
  NOR2_X1 U7363 ( .A1(n6387), .A2(n6386), .ZN(U3019) );
  NOR2_X1 U7364 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6388), .ZN(n6433)
         );
  NAND3_X1 U7365 ( .A1(n6390), .A2(n6389), .A3(n6734), .ZN(n6391) );
  OAI21_X1 U7366 ( .B1(n6394), .B2(n6392), .A(n6391), .ZN(n6432) );
  AOI22_X1 U7367 ( .A1(n6441), .A2(n6433), .B1(n6442), .B2(n6432), .ZN(n6404)
         );
  INV_X1 U7368 ( .A(n6472), .ZN(n6393) );
  OAI21_X1 U7369 ( .B1(n6434), .B2(n6393), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6396) );
  NAND3_X1 U7370 ( .A1(n6396), .A2(n6395), .A3(n6394), .ZN(n6401) );
  INV_X1 U7371 ( .A(n6433), .ZN(n6399) );
  AOI211_X1 U7372 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6399), .A(n6398), .B(
        n6397), .ZN(n6400) );
  NAND3_X1 U7373 ( .A1(n6734), .A2(n6401), .A3(n6400), .ZN(n6436) );
  AOI22_X1 U7374 ( .A1(n6436), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6402), 
        .B2(n6434), .ZN(n6403) );
  OAI211_X1 U7375 ( .C1(n6405), .C2(n6472), .A(n6404), .B(n6403), .ZN(U3068)
         );
  AOI22_X1 U7376 ( .A1(n6447), .A2(n6433), .B1(n6448), .B2(n6432), .ZN(n6408)
         );
  AOI22_X1 U7377 ( .A1(n6436), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6406), 
        .B2(n6434), .ZN(n6407) );
  OAI211_X1 U7378 ( .C1(n6409), .C2(n6472), .A(n6408), .B(n6407), .ZN(U3069)
         );
  AOI22_X1 U7379 ( .A1(n6454), .A2(n6432), .B1(n6453), .B2(n6433), .ZN(n6412)
         );
  AOI22_X1 U7380 ( .A1(n6436), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6410), 
        .B2(n6434), .ZN(n6411) );
  OAI211_X1 U7381 ( .C1(n6413), .C2(n6472), .A(n6412), .B(n6411), .ZN(U3070)
         );
  AOI22_X1 U7382 ( .A1(n6475), .A2(n6433), .B1(n6476), .B2(n6432), .ZN(n6416)
         );
  AOI22_X1 U7383 ( .A1(n6436), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6414), 
        .B2(n6434), .ZN(n6415) );
  OAI211_X1 U7384 ( .C1(n6417), .C2(n6472), .A(n6416), .B(n6415), .ZN(U3071)
         );
  AOI22_X1 U7385 ( .A1(n6481), .A2(n6433), .B1(n6482), .B2(n6432), .ZN(n6420)
         );
  AOI22_X1 U7386 ( .A1(n6436), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6418), 
        .B2(n6434), .ZN(n6419) );
  OAI211_X1 U7387 ( .C1(n6421), .C2(n6472), .A(n6420), .B(n6419), .ZN(U3072)
         );
  AOI22_X1 U7388 ( .A1(n6461), .A2(n6433), .B1(n6462), .B2(n6432), .ZN(n6424)
         );
  AOI22_X1 U7389 ( .A1(n6436), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6422), 
        .B2(n6434), .ZN(n6423) );
  OAI211_X1 U7390 ( .C1(n6425), .C2(n6472), .A(n6424), .B(n6423), .ZN(U3073)
         );
  AOI22_X1 U7391 ( .A1(n6427), .A2(n6433), .B1(n6426), .B2(n6432), .ZN(n6430)
         );
  AOI22_X1 U7392 ( .A1(n6436), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6428), 
        .B2(n6434), .ZN(n6429) );
  OAI211_X1 U7393 ( .C1(n6431), .C2(n6472), .A(n6430), .B(n6429), .ZN(U3074)
         );
  AOI22_X1 U7394 ( .A1(n6489), .A2(n6433), .B1(n6491), .B2(n6432), .ZN(n6438)
         );
  AOI22_X1 U7395 ( .A1(n6436), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6435), 
        .B2(n6434), .ZN(n6437) );
  OAI211_X1 U7396 ( .C1(n6439), .C2(n6472), .A(n6438), .B(n6437), .ZN(U3075)
         );
  AOI22_X1 U7397 ( .A1(n6441), .A2(n6467), .B1(n6440), .B2(n6466), .ZN(n6444)
         );
  AOI22_X1 U7398 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6469), .B1(n6442), 
        .B2(n6468), .ZN(n6443) );
  OAI211_X1 U7399 ( .C1(n6445), .C2(n6472), .A(n6444), .B(n6443), .ZN(U3076)
         );
  AOI22_X1 U7400 ( .A1(n6447), .A2(n6467), .B1(n6446), .B2(n6466), .ZN(n6450)
         );
  AOI22_X1 U7401 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6469), .B1(n6448), 
        .B2(n6468), .ZN(n6449) );
  OAI211_X1 U7402 ( .C1(n6451), .C2(n6472), .A(n6450), .B(n6449), .ZN(U3077)
         );
  AOI22_X1 U7403 ( .A1(n6453), .A2(n6467), .B1(n6452), .B2(n6466), .ZN(n6456)
         );
  AOI22_X1 U7404 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6469), .B1(n6454), 
        .B2(n6468), .ZN(n6455) );
  OAI211_X1 U7405 ( .C1(n6457), .C2(n6472), .A(n6456), .B(n6455), .ZN(U3078)
         );
  AOI22_X1 U7406 ( .A1(n6481), .A2(n6467), .B1(n6480), .B2(n6466), .ZN(n6459)
         );
  AOI22_X1 U7407 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6469), .B1(n6482), 
        .B2(n6468), .ZN(n6458) );
  OAI211_X1 U7408 ( .C1(n6485), .C2(n6472), .A(n6459), .B(n6458), .ZN(U3080)
         );
  AOI22_X1 U7409 ( .A1(n6461), .A2(n6467), .B1(n6460), .B2(n6466), .ZN(n6464)
         );
  AOI22_X1 U7410 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6469), .B1(n6462), 
        .B2(n6468), .ZN(n6463) );
  OAI211_X1 U7411 ( .C1(n6465), .C2(n6472), .A(n6464), .B(n6463), .ZN(U3081)
         );
  AOI22_X1 U7412 ( .A1(n6489), .A2(n6467), .B1(n6487), .B2(n6466), .ZN(n6471)
         );
  AOI22_X1 U7413 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6469), .B1(n6491), 
        .B2(n6468), .ZN(n6470) );
  OAI211_X1 U7414 ( .C1(n6496), .C2(n6472), .A(n6471), .B(n6470), .ZN(U3083)
         );
  INV_X1 U7415 ( .A(n6473), .ZN(n6488) );
  AOI22_X1 U7416 ( .A1(n6475), .A2(n6488), .B1(n6474), .B2(n6486), .ZN(n6478)
         );
  AOI22_X1 U7417 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6492), .B1(n6476), 
        .B2(n6490), .ZN(n6477) );
  OAI211_X1 U7418 ( .C1(n6479), .C2(n6495), .A(n6478), .B(n6477), .ZN(U3111)
         );
  AOI22_X1 U7419 ( .A1(n6481), .A2(n6488), .B1(n6480), .B2(n6486), .ZN(n6484)
         );
  AOI22_X1 U7420 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6492), .B1(n6482), 
        .B2(n6490), .ZN(n6483) );
  OAI211_X1 U7421 ( .C1(n6485), .C2(n6495), .A(n6484), .B(n6483), .ZN(U3112)
         );
  AOI22_X1 U7422 ( .A1(n6489), .A2(n6488), .B1(n6487), .B2(n6486), .ZN(n6494)
         );
  AOI22_X1 U7423 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6492), .B1(n6491), 
        .B2(n6490), .ZN(n6493) );
  OAI211_X1 U7424 ( .C1(n6496), .C2(n6495), .A(n6494), .B(n6493), .ZN(U3115)
         );
  AOI211_X1 U7425 ( .C1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n6498), .A(n6917), .B(n6497), .ZN(n6502) );
  INV_X1 U7426 ( .A(n6499), .ZN(n6501) );
  OAI22_X1 U7427 ( .A1(n6502), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n6501), .B2(n6500), .ZN(n6504) );
  NAND2_X1 U7428 ( .A1(n6502), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6503) );
  OAI211_X1 U7429 ( .C1(n6506), .C2(n6505), .A(n6504), .B(n6503), .ZN(n6509)
         );
  NAND2_X1 U7430 ( .A1(n6506), .A2(n6505), .ZN(n6508) );
  INV_X1 U7431 ( .A(n6511), .ZN(n6507) );
  AOI22_X1 U7432 ( .A1(n6509), .A2(n6508), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6507), .ZN(n6510) );
  AOI21_X1 U7433 ( .B1(n6511), .B2(n6734), .A(n6510), .ZN(n6523) );
  INV_X1 U7434 ( .A(n6512), .ZN(n6522) );
  INV_X1 U7435 ( .A(MORE_REG_SCAN_IN), .ZN(n6514) );
  AOI21_X1 U7436 ( .B1(n6515), .B2(n6514), .A(n6513), .ZN(n6519) );
  INV_X1 U7437 ( .A(n6516), .ZN(n6518) );
  NOR4_X1 U7438 ( .A1(n6520), .A2(n6519), .A3(n6518), .A4(n6517), .ZN(n6521)
         );
  OAI211_X1 U7439 ( .C1(n6523), .C2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(n6522), .B(n6521), .ZN(n6530) );
  AOI22_X1 U7440 ( .A1(n6530), .A2(n6525), .B1(n6524), .B2(n6622), .ZN(n6536)
         );
  INV_X1 U7441 ( .A(n6526), .ZN(n6535) );
  OAI21_X1 U7442 ( .B1(n6537), .B2(n3646), .A(n6910), .ZN(n6527) );
  OAI211_X1 U7443 ( .C1(n6529), .C2(n6528), .A(STATE2_REG_2__SCAN_IN), .B(
        n6527), .ZN(n6544) );
  NOR2_X1 U7444 ( .A1(n6544), .A2(n6530), .ZN(n6623) );
  NOR2_X1 U7445 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n3646), .ZN(n6542) );
  OAI21_X1 U7446 ( .B1(n6623), .B2(n6542), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n6534) );
  OAI211_X1 U7447 ( .C1(n6532), .C2(n6531), .A(n6910), .B(n6544), .ZN(n6533)
         );
  NAND4_X1 U7448 ( .A1(n6536), .A2(n6535), .A3(n6534), .A4(n6533), .ZN(U3148)
         );
  NOR2_X1 U7449 ( .A1(n6910), .A2(n6537), .ZN(n6545) );
  AOI221_X1 U7450 ( .B1(READY_N), .B2(n6539), .C1(n6538), .C2(n6539), .A(n6623), .ZN(n6540) );
  AOI211_X1 U7451 ( .C1(n6542), .C2(n6545), .A(n6541), .B(n6540), .ZN(n6543)
         );
  OAI21_X1 U7452 ( .B1(n6546), .B2(n6544), .A(n6543), .ZN(U3149) );
  AOI21_X1 U7453 ( .B1(n6545), .B2(n3646), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n6547) );
  OAI22_X1 U7454 ( .A1(n6622), .A2(n6547), .B1(n6735), .B2(n6546), .ZN(U3150)
         );
  INV_X1 U7455 ( .A(n6620), .ZN(n6548) );
  AND2_X1 U7456 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6548), .ZN(U3151) );
  AND2_X1 U7457 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6548), .ZN(U3152) );
  AND2_X1 U7458 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6548), .ZN(U3153) );
  AND2_X1 U7459 ( .A1(n6548), .A2(DATAWIDTH_REG_28__SCAN_IN), .ZN(U3154) );
  AND2_X1 U7460 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6548), .ZN(U3155) );
  AND2_X1 U7461 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6548), .ZN(U3156) );
  AND2_X1 U7462 ( .A1(n6548), .A2(DATAWIDTH_REG_25__SCAN_IN), .ZN(U3157) );
  AND2_X1 U7463 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6548), .ZN(U3158) );
  AND2_X1 U7464 ( .A1(n6548), .A2(DATAWIDTH_REG_23__SCAN_IN), .ZN(U3159) );
  AND2_X1 U7465 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6548), .ZN(U3160) );
  AND2_X1 U7466 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6548), .ZN(U3161) );
  AND2_X1 U7467 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6548), .ZN(U3162) );
  INV_X1 U7468 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n6933) );
  NOR2_X1 U7469 ( .A1(n6620), .A2(n6933), .ZN(U3163) );
  AND2_X1 U7470 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6548), .ZN(U3164) );
  AND2_X1 U7471 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6548), .ZN(U3165) );
  AND2_X1 U7472 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6548), .ZN(U3166) );
  AND2_X1 U7473 ( .A1(n6548), .A2(DATAWIDTH_REG_15__SCAN_IN), .ZN(U3167) );
  AND2_X1 U7474 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6548), .ZN(U3168) );
  AND2_X1 U7475 ( .A1(n6548), .A2(DATAWIDTH_REG_13__SCAN_IN), .ZN(U3169) );
  AND2_X1 U7476 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6548), .ZN(U3170) );
  AND2_X1 U7477 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6548), .ZN(U3171) );
  AND2_X1 U7478 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6548), .ZN(U3172) );
  AND2_X1 U7479 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6548), .ZN(U3173) );
  AND2_X1 U7480 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6548), .ZN(U3174) );
  AND2_X1 U7481 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6548), .ZN(U3175) );
  AND2_X1 U7482 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6548), .ZN(U3176) );
  AND2_X1 U7483 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6548), .ZN(U3177) );
  AND2_X1 U7484 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6548), .ZN(U3178) );
  AND2_X1 U7485 ( .A1(n6548), .A2(DATAWIDTH_REG_3__SCAN_IN), .ZN(U3179) );
  AND2_X1 U7486 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6548), .ZN(U3180) );
  AOI22_X1 U7487 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6564) );
  AND2_X1 U7488 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6551) );
  INV_X1 U7489 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6653) );
  OAI21_X1 U7490 ( .B1(n6551), .B2(n6653), .A(n6656), .ZN(n6549) );
  INV_X1 U7491 ( .A(n6550), .ZN(n6563) );
  OAI211_X1 U7492 ( .C1(NA_N), .C2(n6565), .A(n3634), .B(n6563), .ZN(n6560) );
  OAI211_X1 U7493 ( .C1(n6550), .C2(n6564), .A(n6549), .B(n6560), .ZN(U3181)
         );
  NOR2_X1 U7494 ( .A1(n3634), .A2(n6653), .ZN(n6552) );
  NAND2_X1 U7495 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6557) );
  OAI21_X1 U7496 ( .B1(n6552), .B2(n6551), .A(n6557), .ZN(n6553) );
  OAI211_X1 U7497 ( .C1(n6555), .C2(n3646), .A(n6554), .B(n6553), .ZN(U3182)
         );
  NOR4_X1 U7498 ( .A1(NA_N), .A2(n3634), .A3(n3646), .A4(n6653), .ZN(n6561) );
  NOR2_X1 U7499 ( .A1(NA_N), .A2(n3646), .ZN(n6556) );
  OAI211_X1 U7500 ( .C1(n6556), .C2(n6555), .A(HOLD), .B(n6653), .ZN(n6558) );
  NAND3_X1 U7501 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6558), .A3(n6557), .ZN(
        n6559) );
  AOI22_X1 U7502 ( .A1(STATE_REG_1__SCAN_IN), .A2(n6561), .B1(n6560), .B2(
        n6559), .ZN(n6562) );
  OAI21_X1 U7503 ( .B1(n6564), .B2(n6563), .A(n6562), .ZN(U3183) );
  NOR2_X2 U7504 ( .A1(n6565), .A2(n6656), .ZN(n6609) );
  INV_X1 U7505 ( .A(n6609), .ZN(n6614) );
  NAND2_X1 U7506 ( .A1(n6565), .A2(n6655), .ZN(n6611) );
  INV_X1 U7507 ( .A(n6611), .ZN(n6612) );
  AOI22_X1 U7508 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6656), .ZN(n6566) );
  OAI21_X1 U7509 ( .B1(n6632), .B2(n6614), .A(n6566), .ZN(U3184) );
  AOI22_X1 U7510 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6656), .ZN(n6567) );
  OAI21_X1 U7511 ( .B1(n6955), .B2(n6614), .A(n6567), .ZN(U3185) );
  AOI22_X1 U7512 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6656), .ZN(n6568) );
  OAI21_X1 U7513 ( .B1(n6569), .B2(n6614), .A(n6568), .ZN(U3186) );
  AOI22_X1 U7514 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6656), .ZN(n6570) );
  OAI21_X1 U7515 ( .B1(n6725), .B2(n6614), .A(n6570), .ZN(U3187) );
  AOI22_X1 U7516 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6656), .ZN(n6571) );
  OAI21_X1 U7517 ( .B1(n6572), .B2(n6614), .A(n6571), .ZN(U3188) );
  AOI22_X1 U7518 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6656), .ZN(n6573) );
  OAI21_X1 U7519 ( .B1(n6574), .B2(n6614), .A(n6573), .ZN(U3189) );
  AOI22_X1 U7520 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6656), .ZN(n6575) );
  OAI21_X1 U7521 ( .B1(n6576), .B2(n6614), .A(n6575), .ZN(U3190) );
  INV_X1 U7522 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6813) );
  AOI22_X1 U7523 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6656), .ZN(n6577) );
  OAI21_X1 U7524 ( .B1(n6813), .B2(n6611), .A(n6577), .ZN(U3191) );
  AOI22_X1 U7525 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6656), .ZN(n6578) );
  OAI21_X1 U7526 ( .B1(n6579), .B2(n6611), .A(n6578), .ZN(U3192) );
  AOI22_X1 U7527 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6656), .ZN(n6580) );
  OAI21_X1 U7528 ( .B1(n6582), .B2(n6611), .A(n6580), .ZN(U3193) );
  AOI22_X1 U7529 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6656), .ZN(n6581) );
  OAI21_X1 U7530 ( .B1(n6582), .B2(n6614), .A(n6581), .ZN(U3194) );
  AOI22_X1 U7531 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6656), .ZN(n6583) );
  OAI21_X1 U7532 ( .B1(n5316), .B2(n6614), .A(n6583), .ZN(U3195) );
  AOI22_X1 U7533 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6656), .ZN(n6584) );
  OAI21_X1 U7534 ( .B1(n6585), .B2(n6611), .A(n6584), .ZN(U3196) );
  AOI22_X1 U7535 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6656), .ZN(n6586) );
  OAI21_X1 U7536 ( .B1(n6587), .B2(n6611), .A(n6586), .ZN(U3197) );
  AOI22_X1 U7537 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6656), .ZN(n6588) );
  OAI21_X1 U7538 ( .B1(n6590), .B2(n6611), .A(n6588), .ZN(U3198) );
  AOI22_X1 U7539 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6656), .ZN(n6589) );
  OAI21_X1 U7540 ( .B1(n6590), .B2(n6614), .A(n6589), .ZN(U3199) );
  AOI22_X1 U7541 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6656), .ZN(n6591) );
  OAI21_X1 U7542 ( .B1(n6592), .B2(n6611), .A(n6591), .ZN(U3200) );
  AOI22_X1 U7543 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6656), .ZN(n6593) );
  OAI21_X1 U7544 ( .B1(n6595), .B2(n6611), .A(n6593), .ZN(U3201) );
  AOI22_X1 U7545 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6656), .ZN(n6594) );
  OAI21_X1 U7546 ( .B1(n6595), .B2(n6614), .A(n6594), .ZN(U3202) );
  AOI22_X1 U7547 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6656), .ZN(n6596) );
  OAI21_X1 U7548 ( .B1(n6786), .B2(n6611), .A(n6596), .ZN(U3203) );
  AOI22_X1 U7549 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6656), .ZN(n6597) );
  OAI21_X1 U7550 ( .B1(n6786), .B2(n6614), .A(n6597), .ZN(U3204) );
  AOI22_X1 U7551 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6656), .ZN(n6598) );
  OAI21_X1 U7552 ( .B1(n6599), .B2(n6614), .A(n6598), .ZN(U3205) );
  AOI22_X1 U7553 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6656), .ZN(n6600) );
  OAI21_X1 U7554 ( .B1(n6601), .B2(n6611), .A(n6600), .ZN(U3206) );
  AOI222_X1 U7555 ( .A1(n6612), .A2(REIP_REG_25__SCAN_IN), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6656), .C1(REIP_REG_24__SCAN_IN), .C2(
        n6609), .ZN(n6602) );
  INV_X1 U7556 ( .A(n6602), .ZN(U3207) );
  AOI22_X1 U7557 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6656), .ZN(n6603) );
  OAI21_X1 U7558 ( .B1(n6604), .B2(n6614), .A(n6603), .ZN(U3208) );
  AOI22_X1 U7559 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6656), .ZN(n6605) );
  OAI21_X1 U7560 ( .B1(n6606), .B2(n6611), .A(n6605), .ZN(U3209) );
  AOI222_X1 U7561 ( .A1(n6609), .A2(REIP_REG_27__SCAN_IN), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6656), .C1(REIP_REG_28__SCAN_IN), .C2(
        n6612), .ZN(n6607) );
  INV_X1 U7562 ( .A(n6607), .ZN(U3210) );
  AOI22_X1 U7563 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6656), .ZN(n6608) );
  OAI21_X1 U7564 ( .B1(n6816), .B2(n6614), .A(n6608), .ZN(U3211) );
  AOI22_X1 U7565 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6656), .ZN(n6610) );
  OAI21_X1 U7566 ( .B1(n6615), .B2(n6611), .A(n6610), .ZN(U3212) );
  AOI22_X1 U7567 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6656), .ZN(n6613) );
  OAI21_X1 U7568 ( .B1(n6615), .B2(n6614), .A(n6613), .ZN(U3213) );
  OAI22_X1 U7569 ( .A1(n6656), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n6655), .ZN(n6616) );
  INV_X1 U7570 ( .A(n6616), .ZN(U3445) );
  MUX2_X1 U7571 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6656), .Z(U3446) );
  MUX2_X1 U7572 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6656), .Z(U3447) );
  MUX2_X1 U7573 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6656), .Z(U3448) );
  OAI21_X1 U7574 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6620), .A(n6618), .ZN(
        n6617) );
  INV_X1 U7575 ( .A(n6617), .ZN(U3451) );
  OAI21_X1 U7576 ( .B1(n6620), .B2(n6619), .A(n6618), .ZN(U3452) );
  AOI211_X1 U7577 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6623), .A(n6622), .B(
        n6621), .ZN(n6624) );
  INV_X1 U7578 ( .A(n6624), .ZN(U3453) );
  INV_X1 U7579 ( .A(n6625), .ZN(n6629) );
  OAI22_X1 U7580 ( .A1(n6629), .A2(n6628), .B1(n6627), .B2(n6626), .ZN(n6631)
         );
  MUX2_X1 U7581 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6631), .S(n6630), 
        .Z(U3456) );
  AOI21_X1 U7582 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6633) );
  AOI22_X1 U7583 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6633), .B2(n6632), .ZN(n6635) );
  INV_X1 U7584 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6634) );
  AOI22_X1 U7585 ( .A1(n6636), .A2(n6635), .B1(n6634), .B2(n6639), .ZN(U3468)
         );
  INV_X1 U7586 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6640) );
  NOR2_X1 U7587 ( .A1(n6639), .A2(REIP_REG_1__SCAN_IN), .ZN(n6637) );
  AOI22_X1 U7588 ( .A1(n6640), .A2(n6639), .B1(n6638), .B2(n6637), .ZN(U3469)
         );
  NAND2_X1 U7589 ( .A1(n6656), .A2(W_R_N_REG_SCAN_IN), .ZN(n6641) );
  OAI21_X1 U7590 ( .B1(n6656), .B2(READREQUEST_REG_SCAN_IN), .A(n6641), .ZN(
        U3470) );
  INV_X1 U7591 ( .A(n6642), .ZN(n6643) );
  OAI211_X1 U7592 ( .C1(READY_N), .C2(n6645), .A(n6644), .B(n6643), .ZN(n6654)
         );
  NOR2_X1 U7593 ( .A1(n6649), .A2(n6910), .ZN(n6650) );
  OAI21_X1 U7594 ( .B1(n6651), .B2(n6650), .A(n6654), .ZN(n6652) );
  OAI21_X1 U7595 ( .B1(n6654), .B2(n6653), .A(n6652), .ZN(U3472) );
  OAI22_X1 U7596 ( .A1(n6656), .A2(MEMORYFETCH_REG_SCAN_IN), .B1(
        M_IO_N_REG_SCAN_IN), .B2(n6655), .ZN(n6657) );
  INV_X1 U7597 ( .A(n6657), .ZN(U3473) );
  INV_X1 U7598 ( .A(keyinput123), .ZN(n6717) );
  NAND2_X1 U7599 ( .A1(keyinput53), .A2(keyinput97), .ZN(n6658) );
  NOR3_X1 U7600 ( .A1(keyinput22), .A2(keyinput34), .A3(n6658), .ZN(n6659) );
  NAND3_X1 U7601 ( .A1(keyinput82), .A2(keyinput28), .A3(n6659), .ZN(n6672) );
  NAND2_X1 U7602 ( .A1(keyinput127), .A2(keyinput37), .ZN(n6660) );
  NOR3_X1 U7603 ( .A1(keyinput80), .A2(keyinput25), .A3(n6660), .ZN(n6670) );
  NOR4_X1 U7604 ( .A1(keyinput115), .A2(keyinput14), .A3(keyinput26), .A4(
        keyinput88), .ZN(n6669) );
  NOR2_X1 U7605 ( .A1(keyinput18), .A2(keyinput62), .ZN(n6661) );
  NAND3_X1 U7606 ( .A1(keyinput109), .A2(keyinput56), .A3(n6661), .ZN(n6667)
         );
  NOR2_X1 U7607 ( .A1(keyinput2), .A2(keyinput74), .ZN(n6662) );
  NAND3_X1 U7608 ( .A1(keyinput24), .A2(keyinput59), .A3(n6662), .ZN(n6666) );
  NOR2_X1 U7609 ( .A1(keyinput48), .A2(keyinput95), .ZN(n6663) );
  NAND3_X1 U7610 ( .A1(keyinput119), .A2(keyinput126), .A3(n6663), .ZN(n6665)
         );
  NAND4_X1 U7611 ( .A1(keyinput49), .A2(keyinput19), .A3(keyinput41), .A4(
        keyinput92), .ZN(n6664) );
  NOR4_X1 U7612 ( .A1(n6667), .A2(n6666), .A3(n6665), .A4(n6664), .ZN(n6668)
         );
  NAND3_X1 U7613 ( .A1(n6670), .A2(n6669), .A3(n6668), .ZN(n6671) );
  NOR4_X1 U7614 ( .A1(keyinput39), .A2(keyinput11), .A3(n6672), .A4(n6671), 
        .ZN(n6715) );
  INV_X1 U7615 ( .A(keyinput42), .ZN(n6673) );
  NAND4_X1 U7616 ( .A1(keyinput46), .A2(keyinput12), .A3(keyinput1), .A4(n6673), .ZN(n6679) );
  NOR2_X1 U7617 ( .A1(keyinput71), .A2(keyinput113), .ZN(n6674) );
  NAND3_X1 U7618 ( .A1(keyinput83), .A2(keyinput91), .A3(n6674), .ZN(n6678) );
  NOR2_X1 U7619 ( .A1(keyinput70), .A2(keyinput101), .ZN(n6675) );
  NAND3_X1 U7620 ( .A1(keyinput76), .A2(keyinput10), .A3(n6675), .ZN(n6677) );
  NAND4_X1 U7621 ( .A1(keyinput98), .A2(keyinput114), .A3(keyinput122), .A4(
        keyinput8), .ZN(n6676) );
  NOR4_X1 U7622 ( .A1(n6679), .A2(n6678), .A3(n6677), .A4(n6676), .ZN(n6714)
         );
  INV_X1 U7623 ( .A(keyinput31), .ZN(n6680) );
  NAND4_X1 U7624 ( .A1(keyinput69), .A2(keyinput21), .A3(keyinput124), .A4(
        n6680), .ZN(n6684) );
  OR4_X1 U7625 ( .A1(keyinput20), .A2(keyinput4), .A3(keyinput118), .A4(
        keyinput40), .ZN(n6683) );
  OR4_X1 U7626 ( .A1(keyinput65), .A2(keyinput107), .A3(keyinput60), .A4(
        keyinput106), .ZN(n6682) );
  NAND4_X1 U7627 ( .A1(keyinput67), .A2(keyinput104), .A3(keyinput64), .A4(
        keyinput79), .ZN(n6681) );
  NOR4_X1 U7628 ( .A1(n6684), .A2(n6683), .A3(n6682), .A4(n6681), .ZN(n6713)
         );
  NOR4_X1 U7629 ( .A1(keyinput35), .A2(keyinput55), .A3(keyinput27), .A4(
        keyinput103), .ZN(n6685) );
  INV_X1 U7630 ( .A(keyinput43), .ZN(n6846) );
  NAND3_X1 U7631 ( .A1(keyinput89), .A2(n6685), .A3(n6846), .ZN(n6711) );
  NOR2_X1 U7632 ( .A1(keyinput17), .A2(keyinput9), .ZN(n6686) );
  NAND3_X1 U7633 ( .A1(keyinput125), .A2(keyinput111), .A3(n6686), .ZN(n6687)
         );
  NOR3_X1 U7634 ( .A1(keyinput32), .A2(keyinput13), .A3(n6687), .ZN(n6695) );
  NOR3_X1 U7635 ( .A1(keyinput68), .A2(keyinput100), .A3(keyinput57), .ZN(
        n6688) );
  NAND2_X1 U7636 ( .A1(keyinput116), .A2(n6688), .ZN(n6693) );
  NAND4_X1 U7637 ( .A1(keyinput61), .A2(keyinput108), .A3(keyinput44), .A4(
        keyinput66), .ZN(n6692) );
  NOR2_X1 U7638 ( .A1(keyinput47), .A2(keyinput15), .ZN(n6689) );
  NAND3_X1 U7639 ( .A1(keyinput75), .A2(keyinput16), .A3(n6689), .ZN(n6691) );
  NAND4_X1 U7640 ( .A1(keyinput96), .A2(keyinput86), .A3(keyinput121), .A4(
        keyinput23), .ZN(n6690) );
  NOR4_X1 U7641 ( .A1(n6693), .A2(n6692), .A3(n6691), .A4(n6690), .ZN(n6694)
         );
  NAND4_X1 U7642 ( .A1(keyinput120), .A2(keyinput73), .A3(n6695), .A4(n6694), 
        .ZN(n6710) );
  NAND4_X1 U7643 ( .A1(keyinput93), .A2(keyinput51), .A3(keyinput90), .A4(
        keyinput33), .ZN(n6696) );
  NOR3_X1 U7644 ( .A1(keyinput110), .A2(keyinput81), .A3(n6696), .ZN(n6708) );
  INV_X1 U7645 ( .A(keyinput105), .ZN(n6815) );
  NOR4_X1 U7646 ( .A1(keyinput0), .A2(keyinput3), .A3(keyinput38), .A4(n6815), 
        .ZN(n6697) );
  NAND3_X1 U7647 ( .A1(keyinput99), .A2(keyinput77), .A3(n6697), .ZN(n6706) );
  NAND2_X1 U7648 ( .A1(keyinput85), .A2(keyinput63), .ZN(n6698) );
  NOR3_X1 U7649 ( .A1(keyinput72), .A2(keyinput102), .A3(n6698), .ZN(n6704) );
  NAND2_X1 U7650 ( .A1(keyinput7), .A2(keyinput30), .ZN(n6699) );
  NOR3_X1 U7651 ( .A1(keyinput36), .A2(keyinput94), .A3(n6699), .ZN(n6703) );
  NAND2_X1 U7652 ( .A1(keyinput54), .A2(keyinput112), .ZN(n6700) );
  NOR3_X1 U7653 ( .A1(keyinput78), .A2(keyinput29), .A3(n6700), .ZN(n6702) );
  NOR4_X1 U7654 ( .A1(keyinput84), .A2(keyinput5), .A3(keyinput6), .A4(
        keyinput58), .ZN(n6701) );
  NAND4_X1 U7655 ( .A1(n6704), .A2(n6703), .A3(n6702), .A4(n6701), .ZN(n6705)
         );
  NOR4_X1 U7656 ( .A1(keyinput45), .A2(keyinput52), .A3(n6706), .A4(n6705), 
        .ZN(n6707) );
  NAND4_X1 U7657 ( .A1(keyinput117), .A2(keyinput87), .A3(n6708), .A4(n6707), 
        .ZN(n6709) );
  NOR4_X1 U7658 ( .A1(keyinput50), .A2(n6711), .A3(n6710), .A4(n6709), .ZN(
        n6712) );
  NAND4_X1 U7659 ( .A1(n6715), .A2(n6714), .A3(n6713), .A4(n6712), .ZN(n6716)
         );
  AOI21_X1 U7660 ( .B1(n6717), .B2(n6716), .A(DATAO_REG_15__SCAN_IN), .ZN(
        n6979) );
  INV_X1 U7661 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n6719) );
  AOI22_X1 U7662 ( .A1(n6719), .A2(keyinput4), .B1(n5035), .B2(keyinput118), 
        .ZN(n6718) );
  OAI221_X1 U7663 ( .B1(n6719), .B2(keyinput4), .C1(n5035), .C2(keyinput118), 
        .A(n6718), .ZN(n6732) );
  INV_X1 U7664 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n6722) );
  INV_X1 U7665 ( .A(keyinput69), .ZN(n6721) );
  AOI22_X1 U7666 ( .A1(n6722), .A2(keyinput40), .B1(ADDRESS_REG_25__SCAN_IN), 
        .B2(n6721), .ZN(n6720) );
  OAI221_X1 U7667 ( .B1(n6722), .B2(keyinput40), .C1(n6721), .C2(
        ADDRESS_REG_25__SCAN_IN), .A(n6720), .ZN(n6731) );
  INV_X1 U7668 ( .A(keyinput21), .ZN(n6724) );
  AOI22_X1 U7669 ( .A1(n6725), .A2(keyinput31), .B1(DATAO_REG_21__SCAN_IN), 
        .B2(n6724), .ZN(n6723) );
  OAI221_X1 U7670 ( .B1(n6725), .B2(keyinput31), .C1(n6724), .C2(
        DATAO_REG_21__SCAN_IN), .A(n6723), .ZN(n6730) );
  INV_X1 U7671 ( .A(keyinput67), .ZN(n6727) );
  AOI22_X1 U7672 ( .A1(n6728), .A2(keyinput124), .B1(ADDRESS_REG_4__SCAN_IN), 
        .B2(n6727), .ZN(n6726) );
  OAI221_X1 U7673 ( .B1(n6728), .B2(keyinput124), .C1(n6727), .C2(
        ADDRESS_REG_4__SCAN_IN), .A(n6726), .ZN(n6729) );
  NOR4_X1 U7674 ( .A1(n6732), .A2(n6731), .A3(n6730), .A4(n6729), .ZN(n6780)
         );
  AOI22_X1 U7675 ( .A1(n6735), .A2(keyinput104), .B1(n6734), .B2(keyinput65), 
        .ZN(n6733) );
  OAI221_X1 U7676 ( .B1(n6735), .B2(keyinput104), .C1(n6734), .C2(keyinput65), 
        .A(n6733), .ZN(n6747) );
  INV_X1 U7677 ( .A(keyinput60), .ZN(n6737) );
  AOI22_X1 U7678 ( .A1(n3533), .A2(keyinput107), .B1(DATAWIDTH_REG_15__SCAN_IN), .B2(n6737), .ZN(n6736) );
  OAI221_X1 U7679 ( .B1(n3533), .B2(keyinput107), .C1(n6737), .C2(
        DATAWIDTH_REG_15__SCAN_IN), .A(n6736), .ZN(n6746) );
  INV_X1 U7680 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n6740) );
  INV_X1 U7681 ( .A(keyinput106), .ZN(n6739) );
  AOI22_X1 U7682 ( .A1(n6740), .A2(keyinput64), .B1(UWORD_REG_3__SCAN_IN), 
        .B2(n6739), .ZN(n6738) );
  OAI221_X1 U7683 ( .B1(n6740), .B2(keyinput64), .C1(n6739), .C2(
        UWORD_REG_3__SCAN_IN), .A(n6738), .ZN(n6745) );
  INV_X1 U7684 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n6743) );
  INV_X1 U7685 ( .A(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n6742) );
  AOI22_X1 U7686 ( .A1(n6743), .A2(keyinput79), .B1(n6742), .B2(keyinput71), 
        .ZN(n6741) );
  OAI221_X1 U7687 ( .B1(n6743), .B2(keyinput79), .C1(n6742), .C2(keyinput71), 
        .A(n6741), .ZN(n6744) );
  NOR4_X1 U7688 ( .A1(n6747), .A2(n6746), .A3(n6745), .A4(n6744), .ZN(n6779)
         );
  AOI22_X1 U7689 ( .A1(n6749), .A2(keyinput83), .B1(n3646), .B2(keyinput91), 
        .ZN(n6748) );
  OAI221_X1 U7690 ( .B1(n6749), .B2(keyinput83), .C1(n3646), .C2(keyinput91), 
        .A(n6748), .ZN(n6760) );
  AOI22_X1 U7691 ( .A1(n6752), .A2(keyinput113), .B1(keyinput46), .B2(n6751), 
        .ZN(n6750) );
  OAI221_X1 U7692 ( .B1(n6752), .B2(keyinput113), .C1(n6751), .C2(keyinput46), 
        .A(n6750), .ZN(n6759) );
  AOI22_X1 U7693 ( .A1(n4333), .A2(keyinput42), .B1(n4075), .B2(keyinput12), 
        .ZN(n6753) );
  OAI221_X1 U7694 ( .B1(n4333), .B2(keyinput42), .C1(n4075), .C2(keyinput12), 
        .A(n6753), .ZN(n6758) );
  AOI22_X1 U7695 ( .A1(n6756), .A2(keyinput1), .B1(n6755), .B2(keyinput98), 
        .ZN(n6754) );
  OAI221_X1 U7696 ( .B1(n6756), .B2(keyinput1), .C1(n6755), .C2(keyinput98), 
        .A(n6754), .ZN(n6757) );
  NOR4_X1 U7697 ( .A1(n6760), .A2(n6759), .A3(n6758), .A4(n6757), .ZN(n6778)
         );
  INV_X1 U7698 ( .A(keyinput114), .ZN(n6762) );
  AOI22_X1 U7699 ( .A1(n6763), .A2(keyinput122), .B1(DATAWIDTH_REG_3__SCAN_IN), 
        .B2(n6762), .ZN(n6761) );
  OAI221_X1 U7700 ( .B1(n6763), .B2(keyinput122), .C1(n6762), .C2(
        DATAWIDTH_REG_3__SCAN_IN), .A(n6761), .ZN(n6776) );
  INV_X1 U7701 ( .A(keyinput8), .ZN(n6766) );
  INV_X1 U7702 ( .A(keyinput70), .ZN(n6765) );
  AOI22_X1 U7703 ( .A1(n6766), .A2(ADDRESS_REG_12__SCAN_IN), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6765), .ZN(n6764) );
  OAI221_X1 U7704 ( .B1(n6766), .B2(ADDRESS_REG_12__SCAN_IN), .C1(n6765), .C2(
        ADDRESS_REG_26__SCAN_IN), .A(n6764), .ZN(n6775) );
  INV_X1 U7705 ( .A(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n6769) );
  INV_X1 U7706 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n6768) );
  AOI22_X1 U7707 ( .A1(n6769), .A2(keyinput76), .B1(n6768), .B2(keyinput101), 
        .ZN(n6767) );
  OAI221_X1 U7708 ( .B1(n6769), .B2(keyinput76), .C1(n6768), .C2(keyinput101), 
        .A(n6767), .ZN(n6774) );
  INV_X1 U7709 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n6772) );
  INV_X1 U7710 ( .A(DATAI_22_), .ZN(n6771) );
  AOI22_X1 U7711 ( .A1(n6772), .A2(keyinput10), .B1(keyinput117), .B2(n6771), 
        .ZN(n6770) );
  OAI221_X1 U7712 ( .B1(n6772), .B2(keyinput10), .C1(n6771), .C2(keyinput117), 
        .A(n6770), .ZN(n6773) );
  NOR4_X1 U7713 ( .A1(n6776), .A2(n6775), .A3(n6774), .A4(n6773), .ZN(n6777)
         );
  NAND4_X1 U7714 ( .A1(n6780), .A2(n6779), .A3(n6778), .A4(n6777), .ZN(n6978)
         );
  INV_X1 U7715 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n6783) );
  INV_X1 U7716 ( .A(keyinput87), .ZN(n6782) );
  AOI22_X1 U7717 ( .A1(n6783), .A2(keyinput93), .B1(DATAO_REG_28__SCAN_IN), 
        .B2(n6782), .ZN(n6781) );
  OAI221_X1 U7718 ( .B1(n6783), .B2(keyinput93), .C1(n6782), .C2(
        DATAO_REG_28__SCAN_IN), .A(n6781), .ZN(n6796) );
  AOI22_X1 U7719 ( .A1(n6786), .A2(keyinput51), .B1(n6785), .B2(keyinput90), 
        .ZN(n6784) );
  OAI221_X1 U7720 ( .B1(n6786), .B2(keyinput51), .C1(n6785), .C2(keyinput90), 
        .A(n6784), .ZN(n6795) );
  INV_X1 U7721 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n6788) );
  AOI22_X1 U7722 ( .A1(n6789), .A2(keyinput33), .B1(n6788), .B2(keyinput110), 
        .ZN(n6787) );
  OAI221_X1 U7723 ( .B1(n6789), .B2(keyinput33), .C1(n6788), .C2(keyinput110), 
        .A(n6787), .ZN(n6794) );
  AOI22_X1 U7724 ( .A1(n6792), .A2(keyinput81), .B1(n6791), .B2(keyinput36), 
        .ZN(n6790) );
  OAI221_X1 U7725 ( .B1(n6792), .B2(keyinput81), .C1(n6791), .C2(keyinput36), 
        .A(n6790), .ZN(n6793) );
  NOR4_X1 U7726 ( .A1(n6796), .A2(n6795), .A3(n6794), .A4(n6793), .ZN(n6844)
         );
  INV_X1 U7727 ( .A(DATAI_26_), .ZN(n6798) );
  AOI22_X1 U7728 ( .A1(n6799), .A2(keyinput30), .B1(keyinput7), .B2(n6798), 
        .ZN(n6797) );
  OAI221_X1 U7729 ( .B1(n6799), .B2(keyinput30), .C1(n6798), .C2(keyinput7), 
        .A(n6797), .ZN(n6810) );
  AOI22_X1 U7730 ( .A1(n6801), .A2(keyinput94), .B1(n5054), .B2(keyinput63), 
        .ZN(n6800) );
  OAI221_X1 U7731 ( .B1(n6801), .B2(keyinput94), .C1(n5054), .C2(keyinput63), 
        .A(n6800), .ZN(n6809) );
  AOI22_X1 U7732 ( .A1(n3950), .A2(keyinput72), .B1(keyinput85), .B2(n6803), 
        .ZN(n6802) );
  OAI221_X1 U7733 ( .B1(n3950), .B2(keyinput72), .C1(n6803), .C2(keyinput85), 
        .A(n6802), .ZN(n6808) );
  AOI22_X1 U7734 ( .A1(n6806), .A2(keyinput102), .B1(keyinput99), .B2(n6805), 
        .ZN(n6804) );
  OAI221_X1 U7735 ( .B1(n6806), .B2(keyinput102), .C1(n6805), .C2(keyinput99), 
        .A(n6804), .ZN(n6807) );
  NOR4_X1 U7736 ( .A1(n6810), .A2(n6809), .A3(n6808), .A4(n6807), .ZN(n6843)
         );
  INV_X1 U7737 ( .A(keyinput45), .ZN(n6812) );
  AOI22_X1 U7738 ( .A1(n6813), .A2(keyinput77), .B1(LWORD_REG_1__SCAN_IN), 
        .B2(n6812), .ZN(n6811) );
  OAI221_X1 U7739 ( .B1(n6813), .B2(keyinput77), .C1(n6812), .C2(
        LWORD_REG_1__SCAN_IN), .A(n6811), .ZN(n6826) );
  AOI22_X1 U7740 ( .A1(n6816), .A2(keyinput52), .B1(LWORD_REG_14__SCAN_IN), 
        .B2(n6815), .ZN(n6814) );
  OAI221_X1 U7741 ( .B1(n6816), .B2(keyinput52), .C1(n6815), .C2(
        LWORD_REG_14__SCAN_IN), .A(n6814), .ZN(n6825) );
  INV_X1 U7742 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n6818) );
  AOI22_X1 U7743 ( .A1(n6819), .A2(keyinput3), .B1(n6818), .B2(keyinput0), 
        .ZN(n6817) );
  OAI221_X1 U7744 ( .B1(n6819), .B2(keyinput3), .C1(n6818), .C2(keyinput0), 
        .A(n6817), .ZN(n6824) );
  INV_X1 U7745 ( .A(keyinput38), .ZN(n6821) );
  AOI22_X1 U7746 ( .A1(n6822), .A2(keyinput84), .B1(ADDRESS_REG_15__SCAN_IN), 
        .B2(n6821), .ZN(n6820) );
  OAI221_X1 U7747 ( .B1(n6822), .B2(keyinput84), .C1(n6821), .C2(
        ADDRESS_REG_15__SCAN_IN), .A(n6820), .ZN(n6823) );
  NOR4_X1 U7748 ( .A1(n6826), .A2(n6825), .A3(n6824), .A4(n6823), .ZN(n6842)
         );
  INV_X1 U7749 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n6829) );
  INV_X1 U7750 ( .A(DATAI_29_), .ZN(n6828) );
  AOI22_X1 U7751 ( .A1(n6829), .A2(keyinput5), .B1(keyinput6), .B2(n6828), 
        .ZN(n6827) );
  OAI221_X1 U7752 ( .B1(n6829), .B2(keyinput5), .C1(n6828), .C2(keyinput6), 
        .A(n6827), .ZN(n6840) );
  INV_X1 U7753 ( .A(keyinput58), .ZN(n6832) );
  INV_X1 U7754 ( .A(keyinput78), .ZN(n6831) );
  AOI22_X1 U7755 ( .A1(n6832), .A2(CODEFETCH_REG_SCAN_IN), .B1(
        BYTEENABLE_REG_0__SCAN_IN), .B2(n6831), .ZN(n6830) );
  OAI221_X1 U7756 ( .B1(n6832), .B2(CODEFETCH_REG_SCAN_IN), .C1(n6831), .C2(
        BYTEENABLE_REG_0__SCAN_IN), .A(n6830), .ZN(n6839) );
  AOI22_X1 U7757 ( .A1(n6834), .A2(keyinput112), .B1(n3872), .B2(keyinput54), 
        .ZN(n6833) );
  OAI221_X1 U7758 ( .B1(n6834), .B2(keyinput112), .C1(n3872), .C2(keyinput54), 
        .A(n6833), .ZN(n6838) );
  INV_X1 U7759 ( .A(keyinput29), .ZN(n6836) );
  AOI22_X1 U7760 ( .A1(n3711), .A2(keyinput50), .B1(DATAWIDTH_REG_28__SCAN_IN), 
        .B2(n6836), .ZN(n6835) );
  OAI221_X1 U7761 ( .B1(n3711), .B2(keyinput50), .C1(n6836), .C2(
        DATAWIDTH_REG_28__SCAN_IN), .A(n6835), .ZN(n6837) );
  NOR4_X1 U7762 ( .A1(n6840), .A2(n6839), .A3(n6838), .A4(n6837), .ZN(n6841)
         );
  NAND4_X1 U7763 ( .A1(n6844), .A2(n6843), .A3(n6842), .A4(n6841), .ZN(n6977)
         );
  INV_X1 U7764 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6847) );
  AOI22_X1 U7765 ( .A1(n6847), .A2(keyinput61), .B1(DATAO_REG_31__SCAN_IN), 
        .B2(n6846), .ZN(n6845) );
  OAI221_X1 U7766 ( .B1(n6847), .B2(keyinput61), .C1(n6846), .C2(
        DATAO_REG_31__SCAN_IN), .A(n6845), .ZN(n6876) );
  INV_X1 U7767 ( .A(keyinput103), .ZN(n6850) );
  INV_X1 U7768 ( .A(keyinput89), .ZN(n6849) );
  AOI22_X1 U7769 ( .A1(n6850), .A2(M_IO_N_REG_SCAN_IN), .B1(
        DATAO_REG_6__SCAN_IN), .B2(n6849), .ZN(n6848) );
  OAI221_X1 U7770 ( .B1(n6850), .B2(M_IO_N_REG_SCAN_IN), .C1(n6849), .C2(
        DATAO_REG_6__SCAN_IN), .A(n6848), .ZN(n6875) );
  INV_X1 U7771 ( .A(keyinput35), .ZN(n6855) );
  INV_X1 U7772 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n6854) );
  INV_X1 U7773 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n6852) );
  AOI22_X1 U7774 ( .A1(n4826), .A2(keyinput55), .B1(n6852), .B2(keyinput27), 
        .ZN(n6851) );
  OAI221_X1 U7775 ( .B1(n4826), .B2(keyinput55), .C1(n6852), .C2(keyinput27), 
        .A(n6851), .ZN(n6853) );
  AOI221_X1 U7776 ( .B1(INSTQUEUE_REG_15__3__SCAN_IN), .B2(n6855), .C1(n6854), 
        .C2(keyinput35), .A(n6853), .ZN(n6872) );
  INV_X1 U7777 ( .A(keyinput66), .ZN(n6857) );
  AOI22_X1 U7778 ( .A1(n3744), .A2(keyinput116), .B1(ADDRESS_REG_24__SCAN_IN), 
        .B2(n6857), .ZN(n6856) );
  OAI221_X1 U7779 ( .B1(n3744), .B2(keyinput116), .C1(n6857), .C2(
        ADDRESS_REG_24__SCAN_IN), .A(n6856), .ZN(n6870) );
  INV_X1 U7780 ( .A(DATAI_27_), .ZN(n6860) );
  INV_X1 U7781 ( .A(keyinput108), .ZN(n6859) );
  AOI22_X1 U7782 ( .A1(n6860), .A2(keyinput44), .B1(BS16_N), .B2(n6859), .ZN(
        n6858) );
  OAI221_X1 U7783 ( .B1(n6860), .B2(keyinput44), .C1(n6859), .C2(BS16_N), .A(
        n6858), .ZN(n6869) );
  INV_X1 U7784 ( .A(DATAI_21_), .ZN(n6863) );
  INV_X1 U7785 ( .A(keyinput100), .ZN(n6862) );
  AOI22_X1 U7786 ( .A1(n6863), .A2(keyinput96), .B1(LWORD_REG_4__SCAN_IN), 
        .B2(n6862), .ZN(n6861) );
  OAI221_X1 U7787 ( .B1(n6863), .B2(keyinput96), .C1(n6862), .C2(
        LWORD_REG_4__SCAN_IN), .A(n6861), .ZN(n6868) );
  INV_X1 U7788 ( .A(keyinput68), .ZN(n6865) );
  AOI22_X1 U7789 ( .A1(n6866), .A2(keyinput57), .B1(ADDRESS_REG_5__SCAN_IN), 
        .B2(n6865), .ZN(n6864) );
  OAI221_X1 U7790 ( .B1(n6866), .B2(keyinput57), .C1(n6865), .C2(
        ADDRESS_REG_5__SCAN_IN), .A(n6864), .ZN(n6867) );
  NOR4_X1 U7791 ( .A1(n6870), .A2(n6869), .A3(n6868), .A4(n6867), .ZN(n6871)
         );
  OAI211_X1 U7792 ( .C1(keyinput123), .C2(n6873), .A(n6872), .B(n6871), .ZN(
        n6874) );
  NOR3_X1 U7793 ( .A1(n6876), .A2(n6875), .A3(n6874), .ZN(n6975) );
  INV_X1 U7794 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n6879) );
  INV_X1 U7795 ( .A(keyinput17), .ZN(n6878) );
  AOI22_X1 U7796 ( .A1(n6879), .A2(keyinput120), .B1(BE_N_REG_3__SCAN_IN), 
        .B2(n6878), .ZN(n6877) );
  OAI221_X1 U7797 ( .B1(n6879), .B2(keyinput120), .C1(n6878), .C2(
        BE_N_REG_3__SCAN_IN), .A(n6877), .ZN(n6892) );
  INV_X1 U7798 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n6882) );
  INV_X1 U7799 ( .A(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n6881) );
  AOI22_X1 U7800 ( .A1(n6882), .A2(keyinput13), .B1(n6881), .B2(keyinput125), 
        .ZN(n6880) );
  OAI221_X1 U7801 ( .B1(n6882), .B2(keyinput13), .C1(n6881), .C2(keyinput125), 
        .A(n6880), .ZN(n6891) );
  INV_X1 U7802 ( .A(keyinput39), .ZN(n6884) );
  AOI22_X1 U7803 ( .A1(n6885), .A2(keyinput9), .B1(ADDRESS_REG_23__SCAN_IN), 
        .B2(n6884), .ZN(n6883) );
  OAI221_X1 U7804 ( .B1(n6885), .B2(keyinput9), .C1(n6884), .C2(
        ADDRESS_REG_23__SCAN_IN), .A(n6883), .ZN(n6890) );
  INV_X1 U7805 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n6887) );
  AOI22_X1 U7806 ( .A1(n6888), .A2(keyinput73), .B1(n6887), .B2(keyinput111), 
        .ZN(n6886) );
  OAI221_X1 U7807 ( .B1(n6888), .B2(keyinput73), .C1(n6887), .C2(keyinput111), 
        .A(n6886), .ZN(n6889) );
  NOR4_X1 U7808 ( .A1(n6892), .A2(n6891), .A3(n6890), .A4(n6889), .ZN(n6974)
         );
  INV_X1 U7809 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n6894) );
  AOI22_X1 U7810 ( .A1(n3723), .A2(keyinput23), .B1(n6894), .B2(keyinput47), 
        .ZN(n6893) );
  OAI221_X1 U7811 ( .B1(n3723), .B2(keyinput23), .C1(n6894), .C2(keyinput47), 
        .A(n6893), .ZN(n6907) );
  AOI22_X1 U7812 ( .A1(n6897), .A2(keyinput16), .B1(keyinput32), .B2(n6896), 
        .ZN(n6895) );
  OAI221_X1 U7813 ( .B1(n6897), .B2(keyinput16), .C1(n6896), .C2(keyinput32), 
        .A(n6895), .ZN(n6906) );
  INV_X1 U7814 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n6899) );
  AOI22_X1 U7815 ( .A1(n6900), .A2(keyinput15), .B1(n6899), .B2(keyinput121), 
        .ZN(n6898) );
  OAI221_X1 U7816 ( .B1(n6900), .B2(keyinput15), .C1(n6899), .C2(keyinput121), 
        .A(n6898), .ZN(n6905) );
  INV_X1 U7817 ( .A(keyinput86), .ZN(n6901) );
  XOR2_X1 U7818 ( .A(DATAWIDTH_REG_13__SCAN_IN), .B(n6901), .Z(n6903) );
  XNOR2_X1 U7819 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(keyinput75), .ZN(
        n6902) );
  NAND2_X1 U7820 ( .A1(n6903), .A2(n6902), .ZN(n6904) );
  NOR4_X1 U7821 ( .A1(n6907), .A2(n6906), .A3(n6905), .A4(n6904), .ZN(n6973)
         );
  INV_X1 U7822 ( .A(keyinput80), .ZN(n6909) );
  OAI22_X1 U7823 ( .A1(n6910), .A2(keyinput25), .B1(n6909), .B2(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n6908) );
  AOI221_X1 U7824 ( .B1(n6910), .B2(keyinput25), .C1(DATAWIDTH_REG_25__SCAN_IN), .C2(n6909), .A(n6908), .ZN(n6921) );
  INV_X1 U7825 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n6913) );
  INV_X1 U7826 ( .A(keyinput14), .ZN(n6912) );
  OAI22_X1 U7827 ( .A1(n6913), .A2(keyinput37), .B1(n6912), .B2(
        UWORD_REG_5__SCAN_IN), .ZN(n6911) );
  AOI221_X1 U7828 ( .B1(n6913), .B2(keyinput37), .C1(UWORD_REG_5__SCAN_IN), 
        .C2(n6912), .A(n6911), .ZN(n6920) );
  INV_X1 U7829 ( .A(keyinput26), .ZN(n6915) );
  OAI22_X1 U7830 ( .A1(n5858), .A2(keyinput24), .B1(n6915), .B2(
        LWORD_REG_3__SCAN_IN), .ZN(n6914) );
  AOI221_X1 U7831 ( .B1(n5858), .B2(keyinput24), .C1(LWORD_REG_3__SCAN_IN), 
        .C2(n6915), .A(n6914), .ZN(n6919) );
  OAI22_X1 U7832 ( .A1(n6917), .A2(keyinput127), .B1(n5641), .B2(keyinput88), 
        .ZN(n6916) );
  AOI221_X1 U7833 ( .B1(n6917), .B2(keyinput127), .C1(keyinput88), .C2(n5641), 
        .A(n6916), .ZN(n6918) );
  NAND4_X1 U7834 ( .A1(n6921), .A2(n6920), .A3(n6919), .A4(n6918), .ZN(n6971)
         );
  INV_X1 U7835 ( .A(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n6924) );
  INV_X1 U7836 ( .A(keyinput34), .ZN(n6923) );
  OAI22_X1 U7837 ( .A1(n6924), .A2(keyinput22), .B1(n6923), .B2(DATAI_30_), 
        .ZN(n6922) );
  AOI221_X1 U7838 ( .B1(n6924), .B2(keyinput22), .C1(DATAI_30_), .C2(n6923), 
        .A(n6922), .ZN(n6937) );
  INV_X1 U7839 ( .A(keyinput97), .ZN(n6926) );
  OAI22_X1 U7840 ( .A1(keyinput11), .A2(n6927), .B1(n6926), .B2(
        LWORD_REG_7__SCAN_IN), .ZN(n6925) );
  AOI221_X1 U7841 ( .B1(n6927), .B2(keyinput11), .C1(n6926), .C2(
        LWORD_REG_7__SCAN_IN), .A(n6925), .ZN(n6936) );
  OAI22_X1 U7842 ( .A1(n6930), .A2(keyinput28), .B1(n6929), .B2(keyinput115), 
        .ZN(n6928) );
  AOI221_X1 U7843 ( .B1(n6930), .B2(keyinput28), .C1(keyinput115), .C2(n6929), 
        .A(n6928), .ZN(n6935) );
  INV_X1 U7844 ( .A(keyinput82), .ZN(n6932) );
  OAI22_X1 U7845 ( .A1(keyinput53), .A2(n6933), .B1(n6932), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n6931) );
  AOI221_X1 U7846 ( .B1(n6933), .B2(keyinput53), .C1(n6932), .C2(
        DATAO_REG_25__SCAN_IN), .A(n6931), .ZN(n6934) );
  NAND4_X1 U7847 ( .A1(n6937), .A2(n6936), .A3(n6935), .A4(n6934), .ZN(n6970)
         );
  INV_X1 U7848 ( .A(keyinput92), .ZN(n6939) );
  OAI22_X1 U7849 ( .A1(n6940), .A2(keyinput48), .B1(n6939), .B2(
        MEMORYFETCH_REG_SCAN_IN), .ZN(n6938) );
  AOI221_X1 U7850 ( .B1(n6940), .B2(keyinput48), .C1(MEMORYFETCH_REG_SCAN_IN), 
        .C2(n6939), .A(n6938), .ZN(n6953) );
  INV_X1 U7851 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n6943) );
  INV_X1 U7852 ( .A(keyinput41), .ZN(n6942) );
  OAI22_X1 U7853 ( .A1(n6943), .A2(keyinput19), .B1(n6942), .B2(
        ADDRESS_REG_1__SCAN_IN), .ZN(n6941) );
  AOI221_X1 U7854 ( .B1(n6943), .B2(keyinput19), .C1(ADDRESS_REG_1__SCAN_IN), 
        .C2(n6942), .A(n6941), .ZN(n6952) );
  INV_X1 U7855 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6946) );
  INV_X1 U7856 ( .A(keyinput126), .ZN(n6945) );
  OAI22_X1 U7857 ( .A1(n6946), .A2(keyinput20), .B1(n6945), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n6944) );
  AOI221_X1 U7858 ( .B1(n6946), .B2(keyinput20), .C1(DATAO_REG_29__SCAN_IN), 
        .C2(n6945), .A(n6944), .ZN(n6951) );
  INV_X1 U7859 ( .A(keyinput119), .ZN(n6949) );
  INV_X1 U7860 ( .A(keyinput95), .ZN(n6948) );
  OAI22_X1 U7861 ( .A1(n6949), .A2(ADDRESS_REG_21__SCAN_IN), .B1(n6948), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6947) );
  AOI221_X1 U7862 ( .B1(n6949), .B2(ADDRESS_REG_21__SCAN_IN), .C1(
        DATAO_REG_8__SCAN_IN), .C2(n6948), .A(n6947), .ZN(n6950) );
  NAND4_X1 U7863 ( .A1(n6953), .A2(n6952), .A3(n6951), .A4(n6950), .ZN(n6969)
         );
  INV_X1 U7864 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n6956) );
  OAI22_X1 U7865 ( .A1(n6956), .A2(keyinput59), .B1(n6955), .B2(keyinput74), 
        .ZN(n6954) );
  AOI221_X1 U7866 ( .B1(n6956), .B2(keyinput59), .C1(keyinput74), .C2(n6955), 
        .A(n6954), .ZN(n6967) );
  INV_X1 U7867 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n6959) );
  INV_X1 U7868 ( .A(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n6958) );
  OAI22_X1 U7869 ( .A1(n6959), .A2(keyinput2), .B1(n6958), .B2(keyinput18), 
        .ZN(n6957) );
  AOI221_X1 U7870 ( .B1(n6959), .B2(keyinput2), .C1(keyinput18), .C2(n6958), 
        .A(n6957), .ZN(n6966) );
  INV_X1 U7871 ( .A(keyinput62), .ZN(n6961) );
  OAI22_X1 U7872 ( .A1(n5583), .A2(keyinput49), .B1(n6961), .B2(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n6960) );
  AOI221_X1 U7873 ( .B1(n5583), .B2(keyinput49), .C1(DATAWIDTH_REG_23__SCAN_IN), .C2(n6961), .A(n6960), .ZN(n6965) );
  OAI22_X1 U7874 ( .A1(n4822), .A2(keyinput109), .B1(n6963), .B2(keyinput56), 
        .ZN(n6962) );
  AOI221_X1 U7875 ( .B1(n4822), .B2(keyinput109), .C1(keyinput56), .C2(n6963), 
        .A(n6962), .ZN(n6964) );
  NAND4_X1 U7876 ( .A1(n6967), .A2(n6966), .A3(n6965), .A4(n6964), .ZN(n6968)
         );
  NOR4_X1 U7877 ( .A1(n6971), .A2(n6970), .A3(n6969), .A4(n6968), .ZN(n6972)
         );
  NAND4_X1 U7878 ( .A1(n6975), .A2(n6974), .A3(n6973), .A4(n6972), .ZN(n6976)
         );
  NOR4_X1 U7879 ( .A1(n6979), .A2(n6978), .A3(n6977), .A4(n6976), .ZN(n6983)
         );
  AOI222_X1 U7880 ( .A1(EAX_REG_2__SCAN_IN), .A2(n6981), .B1(n6194), .B2(
        LWORD_REG_2__SCAN_IN), .C1(n6980), .C2(DATAO_REG_2__SCAN_IN), .ZN(
        n6982) );
  XNOR2_X1 U7881 ( .A(n6983), .B(n6982), .ZN(U2921) );
  INV_X1 U4114 ( .A(n3658), .ZN(n3251) );
  CLKBUF_X1 U3558 ( .A(n4314), .Z(n4117) );
  NAND2_X1 U4471 ( .A1(n5653), .A2(n5652), .ZN(n5643) );
  NAND2_X1 U3550 ( .A1(n4473), .A2(n4474), .ZN(n4619) );
  CLKBUF_X2 U3577 ( .A(n3352), .Z(n3299) );
  CLKBUF_X1 U3580 ( .A(n5436), .Z(n4217) );
  AND2_X2 U3586 ( .A1(n3560), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3123)
         );
  OR2_X1 U3596 ( .A1(n3624), .A2(n3251), .ZN(n3247) );
  CLKBUF_X2 U3602 ( .A(n3274), .Z(n3278) );
  NAND2_X1 U3644 ( .A1(n3668), .A2(n3667), .ZN(n3672) );
  NAND2_X1 U3679 ( .A1(n3247), .A2(n3246), .ZN(n3769) );
  CLKBUF_X1 U3688 ( .A(n5626), .Z(n5627) );
  NOR2_X2 U3711 ( .A1(n5598), .A2(n5597), .ZN(n5381) );
  CLKBUF_X1 U3741 ( .A(n5373), .Z(n5596) );
  NAND2_X1 U3760 ( .A1(n5395), .A2(n5633), .ZN(n5935) );
  AOI211_X2 U3859 ( .C1(n5015), .C2(n6392), .A(n5013), .B(n5012), .ZN(n5055)
         );
  NOR2_X4 U3914 ( .A1(n4620), .A2(n4619), .ZN(n4618) );
  OR2_X2 U4140 ( .A1(n5606), .A2(n3727), .ZN(n5598) );
  NAND2_X2 U4142 ( .A1(n4961), .A2(n4962), .ZN(n5061) );
  NOR2_X4 U4197 ( .A1(n4714), .A2(n4715), .ZN(n4961) );
  AOI21_X2 U4200 ( .B1(n5484), .B2(n5483), .A(n5482), .ZN(n5488) );
  CLKBUF_X1 U4580 ( .A(n3391), .Z(n4122) );
  CLKBUF_X1 U4605 ( .A(n3299), .Z(n4295) );
endmodule

