

module b14_C_gen_AntiSAT_k_256_2 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, 
        keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, 
        keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, 
        keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, 
        keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, 
        keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, 
        keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, 
        keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, U3352, U3351, U3350, U3349, U3348, U3347, 
        U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, 
        U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, 
        U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, 
        U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, 
        U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, 
        U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, 
        U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, 
        U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, 
        U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, 
        U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, 
        U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, 
        U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, 
        U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, 
        U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, 
        U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, 
        U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, 
        U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, 
        U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, 
        U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, 
        U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, 
        U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, 
        U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, 
        U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, 
        U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5015, n5016;

  OAI21_X1 U2463 ( .B1(n4563), .B2(n4632), .A(n4434), .ZN(n2822) );
  NOR2_X1 U2464 ( .A1(n4381), .A2(n2812), .ZN(n4395) );
  NOR2_X1 U2465 ( .A1(n4382), .A2(n4383), .ZN(n4381) );
  NOR2_X1 U2466 ( .A1(n4372), .A2(n4371), .ZN(n4370) );
  NAND2_X1 U2467 ( .A1(n2385), .A2(n2384), .ZN(n3005) );
  INV_X1 U2468 ( .A(n3591), .ZN(n2899) );
  INV_X1 U2469 ( .A(n2892), .ZN(n2883) );
  NAND2_X1 U2470 ( .A1(n2251), .A2(n3748), .ZN(n3481) );
  OAI21_X1 U2471 ( .B1(n3135), .B2(n3134), .A(n3847), .ZN(n3212) );
  INV_X1 U2472 ( .A(IR_REG_31__SCAN_IN), .ZN(n2732) );
  OR2_X1 U2473 ( .A1(n2407), .A2(n2732), .ZN(n2408) );
  AOI211_X2 U2475 ( .C1(n4201), .C2(n4590), .A(n4200), .B(n4199), .ZN(n4281)
         );
  AOI21_X2 U2476 ( .B1(n3481), .B2(n3490), .A(n3752), .ZN(n4138) );
  XNOR2_X1 U2477 ( .A(n2408), .B(IR_REG_2__SCAN_IN), .ZN(n4341) );
  NAND2_X2 U2478 ( .A1(n3591), .A2(n4606), .ZN(n3606) );
  AND2_X1 U2479 ( .A1(n2381), .A2(n2382), .ZN(n2418) );
  INV_X1 U2480 ( .A(n2382), .ZN(n3012) );
  AND2_X1 U2481 ( .A1(n3628), .A2(n2244), .ZN(n3679) );
  OAI21_X1 U2482 ( .B1(n2296), .B2(n2237), .A(n2293), .ZN(n4116) );
  OR2_X1 U2483 ( .A1(n3363), .A2(n3864), .ZN(n3409) );
  INV_X4 U2484 ( .A(n3606), .ZN(n2947) );
  INV_X1 U2485 ( .A(n2721), .ZN(n2711) );
  OAI21_X1 U2486 ( .B1(n2866), .B2(n4631), .A(n2865), .ZN(n2258) );
  MUX2_X1 U2487 ( .A(REG1_REG_28__SCAN_IN), .B(n2860), .S(n4634), .Z(n2856) );
  MUX2_X1 U2488 ( .A(REG0_REG_28__SCAN_IN), .B(n2860), .S(n4613), .Z(n2861) );
  NAND2_X1 U2489 ( .A1(n3985), .A2(n3762), .ZN(n2850) );
  AOI21_X1 U2490 ( .B1(n2654), .B2(n2286), .A(n2663), .ZN(n2849) );
  NAND2_X1 U2491 ( .A1(n3986), .A2(n3990), .ZN(n3985) );
  OAI21_X1 U2492 ( .B1(n4023), .B2(n2362), .A(n2363), .ZN(n2645) );
  OAI22_X1 U2493 ( .A1(n4040), .A2(n2638), .B1(n4051), .B2(n4029), .ZN(n4023)
         );
  NAND2_X1 U2494 ( .A1(n2290), .A2(n2287), .ZN(n4040) );
  NAND2_X1 U2495 ( .A1(n3750), .A2(n3454), .ZN(n3470) );
  NAND2_X1 U2496 ( .A1(n4481), .A2(n2830), .ZN(n2832) );
  NAND2_X1 U2497 ( .A1(n3529), .A2(n3528), .ZN(n4351) );
  NAND2_X1 U2498 ( .A1(n2259), .A2(n3862), .ZN(n3363) );
  OAI21_X1 U2499 ( .B1(n3320), .B2(n2499), .A(n2500), .ZN(n4515) );
  NAND2_X1 U2500 ( .A1(n2695), .A2(n3840), .ZN(n3236) );
  OAI21_X1 U2501 ( .B1(n3198), .B2(n2694), .A(n3838), .ZN(n3135) );
  INV_X2 U2502 ( .A(n4182), .ZN(n2222) );
  NAND2_X1 U2503 ( .A1(n3850), .A2(n3841), .ZN(n3785) );
  NAND2_X1 U2504 ( .A1(n3126), .A2(n3192), .ZN(n3850) );
  INV_X2 U2505 ( .A(n3600), .ZN(n3607) );
  AND2_X2 U2506 ( .A1(n3152), .A2(n2869), .ZN(n3591) );
  NAND2_X1 U2507 ( .A1(n2740), .A2(n2739), .ZN(n2869) );
  NAND2_X1 U2508 ( .A1(n2711), .A2(n3903), .ZN(n3152) );
  AND2_X1 U2509 ( .A1(n3037), .A2(n2807), .ZN(n4372) );
  NAND2_X2 U2511 ( .A1(n3012), .A2(n4335), .ZN(n2431) );
  XNOR2_X1 U2512 ( .A(n2684), .B(n2683), .ZN(n3903) );
  XNOR2_X1 U2513 ( .A(n2379), .B(n3620), .ZN(n2381) );
  NOR2_X1 U2514 ( .A1(n2679), .A2(n2678), .ZN(n2730) );
  NAND2_X1 U2515 ( .A1(n3619), .A2(IR_REG_31__SCAN_IN), .ZN(n2379) );
  XNOR2_X1 U2516 ( .A(n2380), .B(n4720), .ZN(n2382) );
  NAND2_X1 U2517 ( .A1(n2596), .A2(n2595), .ZN(n2679) );
  OAI21_X1 U2518 ( .B1(n2299), .B2(IR_REG_28__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2380) );
  NOR2_X1 U2519 ( .A1(n2371), .A2(IR_REG_13__SCAN_IN), .ZN(n2357) );
  INV_X1 U2520 ( .A(IR_REG_16__SCAN_IN), .ZN(n4887) );
  INV_X1 U2521 ( .A(IR_REG_3__SCAN_IN), .ZN(n2424) );
  NOR2_X1 U2522 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2257)
         );
  NOR2_X1 U2523 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2256)
         );
  NOR2_X1 U2524 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2255)
         );
  NOR2_X1 U2525 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2254)
         );
  INV_X1 U2526 ( .A(IR_REG_25__SCAN_IN), .ZN(n4753) );
  NOR2_X2 U2527 ( .A1(n4156), .A2(n3787), .ZN(n4126) );
  NAND2_X4 U2528 ( .A1(n2869), .A2(n2868), .ZN(n2892) );
  NOR2_X2 U2529 ( .A1(n4504), .A2(n4503), .ZN(n4505) );
  NOR2_X2 U2530 ( .A1(n2833), .A2(n4492), .ZN(n4504) );
  INV_X1 U2531 ( .A(n3591), .ZN(n2223) );
  NOR2_X2 U2532 ( .A1(n3138), .A2(n3269), .ZN(n3217) );
  NAND2_X1 U2533 ( .A1(n3012), .A2(n4335), .ZN(n2224) );
  NAND2_X1 U2534 ( .A1(n3012), .A2(n4335), .ZN(n2225) );
  NOR2_X2 U2535 ( .A1(n3487), .A2(n2277), .ZN(n4171) );
  OR2_X2 U2536 ( .A1(n3460), .A2(n3520), .ZN(n3487) );
  NOR2_X2 U2537 ( .A1(n3414), .A2(n3418), .ZN(n3461) );
  NOR2_X4 U2538 ( .A1(n3234), .A2(n3296), .ZN(n4592) );
  OR2_X2 U2539 ( .A1(n3216), .A2(n3238), .ZN(n3234) );
  AND2_X1 U2540 ( .A1(n2872), .A2(n3152), .ZN(n3600) );
  AND2_X1 U2541 ( .A1(n2671), .A2(n2670), .ZN(n3966) );
  AND2_X1 U2542 ( .A1(n4531), .A2(n2398), .ZN(n2392) );
  INV_X1 U2543 ( .A(n2416), .ZN(n2268) );
  INV_X1 U2544 ( .A(IR_REG_18__SCAN_IN), .ZN(n2595) );
  INV_X1 U2545 ( .A(n2594), .ZN(n2596) );
  OAI22_X1 U2546 ( .A1(n4268), .A2(n3606), .B1(n3602), .B2(n3496), .ZN(n3436)
         );
  OAI22_X1 U2547 ( .A1(n2899), .A2(n3171), .B1(n4536), .B2(n2892), .ZN(n2900)
         );
  AND2_X1 U2548 ( .A1(n2632), .A2(REG3_REG_24__SCAN_IN), .ZN(n2647) );
  AOI21_X1 U2549 ( .B1(n3934), .B2(n3051), .A(n2264), .ZN(n3050) );
  XNOR2_X1 U2550 ( .A(n2784), .B(n2783), .ZN(n4446) );
  NOR2_X1 U2551 ( .A1(n3808), .A2(n2285), .ZN(n2284) );
  INV_X1 U2552 ( .A(n2286), .ZN(n2285) );
  OR2_X1 U2553 ( .A1(n4117), .A2(n4224), .ZN(n2615) );
  AND2_X1 U2554 ( .A1(n2871), .A2(n2721), .ZN(n3153) );
  XNOR2_X1 U2555 ( .A(n2247), .B(n3809), .ZN(n2366) );
  NAND2_X1 U2556 ( .A1(n2248), .A2(n3763), .ZN(n2247) );
  NAND2_X1 U2557 ( .A1(n2850), .A2(n3764), .ZN(n2248) );
  NAND2_X1 U2558 ( .A1(n4496), .A2(n4498), .ZN(n4497) );
  INV_X1 U2559 ( .A(n3436), .ZN(n2343) );
  INV_X1 U2560 ( .A(n3225), .ZN(n2975) );
  NOR2_X1 U2561 ( .A1(n4081), .A2(n2616), .ZN(n2292) );
  INV_X1 U2562 ( .A(n4128), .ZN(n3787) );
  NAND2_X1 U2563 ( .A1(n2311), .A2(n2310), .ZN(n2309) );
  INV_X1 U2564 ( .A(n3123), .ZN(n2310) );
  INV_X1 U2565 ( .A(n3122), .ZN(n2311) );
  NAND2_X1 U2566 ( .A1(n3122), .A2(n3123), .ZN(n2308) );
  NAND2_X1 U2567 ( .A1(n2241), .A2(n2326), .ZN(n2325) );
  NAND2_X1 U2568 ( .A1(n3723), .A2(n2327), .ZN(n2326) );
  INV_X1 U2569 ( .A(n3660), .ZN(n2327) );
  OR3_X1 U2570 ( .A1(n2525), .A2(n2524), .A3(n2523), .ZN(n2535) );
  OR2_X1 U2571 ( .A1(n3438), .A2(n2343), .ZN(n2342) );
  NAND2_X1 U2572 ( .A1(n3438), .A2(n2343), .ZN(n2341) );
  AOI21_X1 U2573 ( .B1(n2323), .B2(n2325), .A(n2322), .ZN(n2321) );
  INV_X1 U2574 ( .A(n3623), .ZN(n2322) );
  INV_X1 U2575 ( .A(n2328), .ZN(n2323) );
  INV_X1 U2576 ( .A(n2308), .ZN(n2307) );
  INV_X1 U2577 ( .A(n2306), .ZN(n2305) );
  OAI21_X1 U2578 ( .B1(n2309), .B2(n2307), .A(n3189), .ZN(n2306) );
  INV_X1 U2579 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2524) );
  NAND2_X1 U2580 ( .A1(n3583), .A2(n3581), .ZN(n3680) );
  AOI21_X1 U2581 ( .B1(n2347), .B2(n2350), .A(n2346), .ZN(n2345) );
  NAND2_X1 U2582 ( .A1(n2388), .A2(n2714), .ZN(n2389) );
  NAND2_X1 U2583 ( .A1(n2226), .A2(n3012), .ZN(n2398) );
  NAND2_X1 U2584 ( .A1(n3768), .A2(REG2_REG_1__SCAN_IN), .ZN(n2400) );
  NAND2_X1 U2585 ( .A1(n2419), .A2(REG1_REG_1__SCAN_IN), .ZN(n2399) );
  INV_X1 U2586 ( .A(n4174), .ZN(n4170) );
  XNOR2_X1 U2587 ( .A(n2954), .B(n3607), .ZN(n2958) );
  NOR2_X1 U2588 ( .A1(n2535), .A2(n4884), .ZN(n2542) );
  INV_X1 U2589 ( .A(n4344), .ZN(n3738) );
  INV_X1 U2590 ( .A(n3152), .ZN(n2868) );
  OR2_X1 U2591 ( .A1(n2730), .A2(n2732), .ZN(n2681) );
  OAI21_X1 U2592 ( .B1(n2221), .B2(REG2_REG_2__SCAN_IN), .A(n2265), .ZN(n2264)
         );
  NAND2_X1 U2593 ( .A1(n4375), .A2(n2771), .ZN(n2773) );
  NAND2_X1 U2594 ( .A1(n4398), .A2(n2775), .ZN(n2776) );
  NAND2_X1 U2595 ( .A1(n4437), .A2(n2782), .ZN(n2784) );
  NAND2_X1 U2596 ( .A1(n4446), .A2(REG2_REG_12__SCAN_IN), .ZN(n4445) );
  OAI22_X1 U2597 ( .A1(n3808), .A2(n2662), .B1(n3613), .B2(n3966), .ZN(n2282)
         );
  AND2_X1 U2598 ( .A1(n2653), .A2(n2245), .ZN(n2286) );
  AND2_X1 U2599 ( .A1(n3764), .A2(n3763), .ZN(n3808) );
  NAND2_X1 U2600 ( .A1(n4198), .A2(n4014), .ZN(n2653) );
  AND2_X1 U2601 ( .A1(n3892), .A2(n3762), .ZN(n3990) );
  OR2_X1 U2602 ( .A1(n3793), .A2(n2288), .ZN(n2287) );
  NAND2_X1 U2603 ( .A1(n2618), .A2(n2230), .ZN(n2290) );
  AND2_X1 U2604 ( .A1(n3791), .A2(n2289), .ZN(n2288) );
  AND2_X1 U2605 ( .A1(n2618), .A2(n2292), .ZN(n4080) );
  AND2_X1 U2606 ( .A1(n2294), .A2(n3813), .ZN(n2293) );
  OR2_X1 U2607 ( .A1(n2586), .A2(n2237), .ZN(n2294) );
  OR2_X1 U2608 ( .A1(n2564), .A2(n2563), .ZN(n2577) );
  AND4_X1 U2609 ( .A1(n2582), .A2(n2581), .A3(n2580), .A4(n2579), .ZN(n4149)
         );
  NAND2_X1 U2610 ( .A1(n3470), .A2(n2700), .ZN(n2251) );
  NAND2_X1 U2611 ( .A1(n3451), .A2(n2368), .ZN(n2298) );
  NAND2_X1 U2612 ( .A1(n2551), .A2(REG3_REG_16__SCAN_IN), .ZN(n2564) );
  NAND2_X1 U2613 ( .A1(n2501), .A2(REG3_REG_11__SCAN_IN), .ZN(n2525) );
  OR2_X1 U2614 ( .A1(n2477), .A2(n2476), .ZN(n2490) );
  OAI21_X1 U2615 ( .B1(n3278), .B2(n3277), .A(n3845), .ZN(n3321) );
  INV_X1 U2616 ( .A(n4511), .ZN(n3279) );
  NAND2_X1 U2617 ( .A1(n2252), .A2(n3849), .ZN(n3278) );
  NAND2_X1 U2618 ( .A1(n3295), .A2(n3844), .ZN(n2252) );
  AND2_X1 U2619 ( .A1(n2232), .A2(n3292), .ZN(n2472) );
  NAND2_X1 U2620 ( .A1(n2459), .A2(REG3_REG_8__SCAN_IN), .ZN(n2477) );
  AND4_X1 U2621 ( .A1(n2449), .A2(n2448), .A3(n2447), .A4(n2446), .ZN(n2965)
         );
  AND3_X1 U2622 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2453) );
  OR2_X1 U2623 ( .A1(n2857), .A2(n3968), .ZN(n4190) );
  NAND2_X1 U2624 ( .A1(n3996), .A2(n3613), .ZN(n2857) );
  INV_X1 U2625 ( .A(n3924), .ZN(n3339) );
  NAND2_X1 U2626 ( .A1(n3153), .A2(n3903), .ZN(n4606) );
  INV_X1 U2627 ( .A(n2299), .ZN(n2716) );
  INV_X1 U2628 ( .A(n2377), .ZN(n2269) );
  INV_X1 U2629 ( .A(IR_REG_19__SCAN_IN), .ZN(n2677) );
  AND2_X1 U2630 ( .A1(n2664), .A2(n2656), .ZN(n3991) );
  INV_X1 U2631 ( .A(n3923), .ZN(n3324) );
  OR2_X1 U2632 ( .A1(n2655), .A2(n2648), .ZN(n4017) );
  OR2_X1 U2633 ( .A1(n2606), .A2(n2605), .ZN(n4146) );
  INV_X1 U2634 ( .A(n4513), .ZN(n3921) );
  NAND2_X1 U2635 ( .A1(n2766), .A2(n2765), .ZN(n3935) );
  OR2_X1 U2636 ( .A1(n3005), .A2(REG2_REG_1__SCAN_IN), .ZN(n2766) );
  XNOR2_X1 U2637 ( .A(n2773), .B(n2772), .ZN(n4387) );
  NAND2_X1 U2638 ( .A1(n4387), .A2(REG2_REG_6__SCAN_IN), .ZN(n4386) );
  XNOR2_X1 U2639 ( .A(n2776), .B(n2814), .ZN(n4407) );
  NAND2_X1 U2640 ( .A1(n4407), .A2(REG2_REG_8__SCAN_IN), .ZN(n4406) );
  NAND2_X1 U2641 ( .A1(n4417), .A2(n4418), .ZN(n4416) );
  NAND2_X1 U2642 ( .A1(n4487), .A2(n2791), .ZN(n4496) );
  INV_X1 U2643 ( .A(n3954), .ZN(n4181) );
  NAND2_X1 U2644 ( .A1(n3969), .A2(n2231), .ZN(n2866) );
  INV_X1 U2645 ( .A(IR_REG_6__SCAN_IN), .ZN(n2485) );
  NAND2_X1 U2646 ( .A1(n2352), .A2(n3562), .ZN(n2349) );
  INV_X1 U2647 ( .A(n2364), .ZN(n2346) );
  INV_X1 U2648 ( .A(n3545), .ZN(n2336) );
  AOI21_X1 U2649 ( .B1(n3437), .B2(n2238), .A(n2338), .ZN(n3529) );
  OAI21_X1 U2650 ( .B1(n2341), .B2(n2340), .A(n2339), .ZN(n2338) );
  INV_X1 U2651 ( .A(n3517), .ZN(n2339) );
  AOI21_X1 U2652 ( .B1(n4395), .B2(n4391), .A(n4390), .ZN(n2815) );
  NAND2_X1 U2653 ( .A1(n4413), .A2(n2818), .ZN(n2819) );
  INV_X1 U2654 ( .A(n2625), .ZN(n2289) );
  INV_X1 U2655 ( .A(n2292), .ZN(n2291) );
  AOI21_X1 U2656 ( .B1(n4120), .B2(n2707), .A(n2706), .ZN(n4061) );
  INV_X1 U2657 ( .A(n2587), .ZN(n2295) );
  OR2_X1 U2658 ( .A1(n2471), .A2(n2470), .ZN(n3292) );
  INV_X1 U2659 ( .A(n3828), .ZN(n2250) );
  NOR2_X1 U2660 ( .A1(n3331), .A2(n4510), .ZN(n2280) );
  NAND2_X1 U2661 ( .A1(n3330), .A2(n3329), .ZN(n3331) );
  NOR2_X1 U2662 ( .A1(n4544), .A2(n3165), .ZN(n3111) );
  NAND2_X1 U2663 ( .A1(n2279), .A2(IR_REG_31__SCAN_IN), .ZN(n2387) );
  NAND2_X1 U2664 ( .A1(n2253), .A2(n2378), .ZN(n2279) );
  AND2_X1 U2665 ( .A1(n2375), .A2(n2373), .ZN(n2270) );
  AND2_X1 U2666 ( .A1(n2372), .A2(n2374), .ZN(n2271) );
  INV_X1 U2667 ( .A(n2570), .ZN(n2272) );
  NAND2_X1 U2668 ( .A1(n2358), .A2(n2357), .ZN(n2571) );
  INV_X1 U2669 ( .A(IR_REG_11__SCAN_IN), .ZN(n2515) );
  OR2_X1 U2670 ( .A1(n2508), .A2(IR_REG_10__SCAN_IN), .ZN(n2509) );
  NOR2_X1 U2671 ( .A1(n2440), .A2(IR_REG_5__SCAN_IN), .ZN(n2487) );
  INV_X1 U2672 ( .A(IR_REG_7__SCAN_IN), .ZN(n2484) );
  NOR2_X1 U2673 ( .A1(n2330), .A2(n2329), .ZN(n2328) );
  INV_X1 U2674 ( .A(n2241), .ZN(n2330) );
  INV_X1 U2675 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4884) );
  OR2_X1 U2676 ( .A1(n2989), .A2(n3312), .ZN(n2993) );
  NAND2_X1 U2677 ( .A1(n2876), .A2(n2875), .ZN(n2877) );
  AOI21_X1 U2678 ( .B1(n2947), .B2(n2874), .A(n2878), .ZN(n2880) );
  AOI21_X1 U2679 ( .B1(n2321), .B2(n2324), .A(n2243), .ZN(n2319) );
  INV_X1 U2680 ( .A(n2325), .ZN(n2324) );
  NOR2_X1 U2681 ( .A1(n2626), .A2(n3634), .ZN(n2632) );
  OR2_X1 U2682 ( .A1(n3606), .A2(n3064), .ZN(n2889) );
  OAI21_X1 U2683 ( .B1(n3710), .B2(n2333), .A(n2332), .ZN(n3692) );
  INV_X1 U2684 ( .A(n2334), .ZN(n2333) );
  AOI21_X1 U2685 ( .B1(n2334), .B2(n3713), .A(n2242), .ZN(n2332) );
  NOR2_X1 U2686 ( .A1(n3640), .A2(n2239), .ZN(n2334) );
  NOR2_X1 U2687 ( .A1(n3561), .A2(n3648), .ZN(n2353) );
  NAND2_X1 U2688 ( .A1(n2356), .A2(n2355), .ZN(n2354) );
  INV_X1 U2689 ( .A(n3651), .ZN(n2356) );
  OAI22_X1 U2690 ( .A1(n2894), .A2(n2892), .B1(n2223), .B2(n4545), .ZN(n2893)
         );
  NAND2_X1 U2691 ( .A1(n2902), .A2(n2901), .ZN(n2922) );
  AOI21_X1 U2692 ( .B1(n3668), .B2(n3670), .A(n3669), .ZN(n3710) );
  NOR2_X1 U2693 ( .A1(n3710), .A2(n3711), .ZN(n3709) );
  AOI22_X1 U2694 ( .A1(n3019), .A2(REG2_REG_3__SCAN_IN), .B1(n4340), .B2(n2768), .ZN(n2770) );
  XNOR2_X1 U2695 ( .A(n2815), .B(n2814), .ZN(n4405) );
  NAND2_X1 U2696 ( .A1(n4405), .A2(REG1_REG_8__SCAN_IN), .ZN(n4404) );
  XNOR2_X1 U2697 ( .A(n2819), .B(n2779), .ZN(n4426) );
  NAND2_X1 U2698 ( .A1(n4416), .A2(n2778), .ZN(n2780) );
  NAND2_X1 U2699 ( .A1(n4462), .A2(n2825), .ZN(n2827) );
  OAI21_X1 U2700 ( .B1(n4468), .B2(n2261), .A(n2260), .ZN(n2790) );
  NAND2_X1 U2701 ( .A1(n4477), .A2(n2262), .ZN(n2260) );
  OR2_X1 U2702 ( .A1(n2787), .A2(n2789), .ZN(n2261) );
  NAND2_X1 U2703 ( .A1(n2837), .A2(n2838), .ZN(n3947) );
  OR2_X1 U2704 ( .A1(n2619), .A2(n3703), .ZN(n2626) );
  AOI22_X1 U2705 ( .A1(n4116), .A2(n2607), .B1(n3787), .B2(n4146), .ZN(n4098)
         );
  AND2_X1 U2706 ( .A1(n2588), .A2(REG3_REG_19__SCAN_IN), .ZN(n2600) );
  NOR2_X1 U2707 ( .A1(n2577), .A2(n3716), .ZN(n2588) );
  AND4_X1 U2708 ( .A1(n2569), .A2(n2568), .A3(n2567), .A4(n2566), .ZN(n4178)
         );
  AND2_X1 U2709 ( .A1(n2561), .A2(n2550), .ZN(n2297) );
  INV_X1 U2710 ( .A(n3786), .ZN(n3454) );
  INV_X1 U2711 ( .A(n3496), .ZN(n3418) );
  INV_X1 U2712 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4973) );
  INV_X1 U2713 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2444) );
  NOR2_X1 U2714 ( .A1(n2452), .A2(n2444), .ZN(n2459) );
  NAND2_X1 U2715 ( .A1(n3107), .A2(n3834), .ZN(n3198) );
  NAND2_X1 U2716 ( .A1(n3835), .A2(n3838), .ZN(n3784) );
  NAND2_X1 U2717 ( .A1(n2713), .A2(n2712), .ZN(n4519) );
  INV_X1 U2718 ( .A(n2688), .ZN(n2249) );
  NAND2_X1 U2719 ( .A1(n2250), .A2(n2688), .ZN(n4538) );
  INV_X1 U2720 ( .A(n3154), .ZN(n4546) );
  INV_X1 U2721 ( .A(n4531), .ZN(n4545) );
  INV_X1 U2722 ( .A(n4535), .ZN(n4175) );
  NAND2_X1 U2723 ( .A1(n2250), .A2(n3827), .ZN(n3781) );
  AND2_X1 U2724 ( .A1(n4033), .A2(n4014), .ZN(n4016) );
  NOR2_X1 U2725 ( .A1(n4053), .A2(n4032), .ZN(n4033) );
  INV_X1 U2726 ( .A(n3579), .ZN(n4051) );
  OR2_X1 U2727 ( .A1(n4073), .A2(n4051), .ZN(n4053) );
  INV_X1 U2728 ( .A(n3632), .ZN(n4071) );
  NAND2_X1 U2729 ( .A1(n4103), .A2(n2276), .ZN(n4073) );
  NOR2_X1 U2730 ( .A1(n4071), .A2(n4085), .ZN(n2276) );
  NAND2_X1 U2731 ( .A1(n4103), .A2(n4091), .ZN(n4090) );
  AND2_X1 U2732 ( .A1(n4126), .A2(n4224), .ZN(n4103) );
  NAND2_X1 U2733 ( .A1(n3772), .A2(DATAI_21_), .ZN(n4224) );
  NAND2_X1 U2734 ( .A1(n3772), .A2(DATAI_20_), .ZN(n4128) );
  NAND2_X1 U2735 ( .A1(n4171), .A2(n4170), .ZN(n4168) );
  NAND2_X1 U2736 ( .A1(n4243), .A2(n4346), .ZN(n2277) );
  AND4_X1 U2737 ( .A1(n2556), .A2(n2555), .A3(n2554), .A4(n2553), .ZN(n4244)
         );
  NOR2_X1 U2738 ( .A1(n3487), .A2(n3486), .ZN(n3509) );
  AND4_X1 U2739 ( .A1(n2540), .A2(n2539), .A3(n2538), .A4(n2537), .ZN(n4258)
         );
  INV_X1 U2740 ( .A(n3464), .ZN(n4266) );
  NAND2_X1 U2741 ( .A1(n2280), .A2(n3425), .ZN(n3414) );
  INV_X1 U2742 ( .A(n2280), .ZN(n4522) );
  AND2_X1 U2743 ( .A1(n4592), .A2(n3338), .ZN(n3330) );
  INV_X1 U2744 ( .A(n3282), .ZN(n3338) );
  INV_X1 U2745 ( .A(n4530), .ZN(n4265) );
  INV_X1 U2746 ( .A(n4532), .ZN(n4267) );
  AND2_X1 U2747 ( .A1(n3111), .A2(n3091), .ZN(n3205) );
  AND2_X1 U2748 ( .A1(n3153), .A2(n4338), .ZN(n4530) );
  INV_X1 U2749 ( .A(n4606), .ZN(n4169) );
  NAND2_X1 U2750 ( .A1(n4545), .A2(n4546), .ZN(n4544) );
  INV_X1 U2751 ( .A(n2912), .ZN(n3150) );
  AND3_X1 U2752 ( .A1(n2755), .A2(n2754), .A3(n2910), .ZN(n2855) );
  INV_X1 U2753 ( .A(n2387), .ZN(n2715) );
  XNOR2_X1 U2754 ( .A(n2686), .B(n4785), .ZN(n2871) );
  NAND2_X1 U2755 ( .A1(n2682), .A2(IR_REG_31__SCAN_IN), .ZN(n2684) );
  NAND2_X1 U2756 ( .A1(n3121), .A2(n2309), .ZN(n2304) );
  NAND2_X1 U2757 ( .A1(n3437), .A2(n2342), .ZN(n2337) );
  INV_X1 U2758 ( .A(n3322), .ZN(n3329) );
  AND2_X1 U2759 ( .A1(n2661), .A2(n2660), .ZN(n3729) );
  AND2_X1 U2760 ( .A1(n2321), .A2(n2331), .ZN(n2317) );
  OAI21_X1 U2761 ( .B1(n2331), .B2(n2319), .A(n2314), .ZN(n2313) );
  NAND2_X1 U2762 ( .A1(n2319), .A2(n2315), .ZN(n2314) );
  NAND2_X1 U2763 ( .A1(n2316), .A2(n3611), .ZN(n2315) );
  INV_X1 U2764 ( .A(n2321), .ZN(n2316) );
  NAND2_X1 U2765 ( .A1(n2319), .A2(n3611), .ZN(n2318) );
  AND2_X1 U2766 ( .A1(n3970), .A2(n2665), .ZN(n3978) );
  AOI21_X1 U2767 ( .B1(n2305), .B2(n2307), .A(n2240), .ZN(n2302) );
  INV_X1 U2768 ( .A(n4146), .ZN(n4225) );
  AND4_X1 U2769 ( .A1(n2507), .A2(n2506), .A3(n2505), .A4(n2504), .ZN(n3426)
         );
  AND4_X1 U2770 ( .A1(n2423), .A2(n2422), .A3(n2421), .A4(n2420), .ZN(n2870)
         );
  NAND2_X1 U2771 ( .A1(n3097), .A2(n3096), .ZN(n3095) );
  XNOR2_X1 U2772 ( .A(n2958), .B(n2956), .ZN(n3096) );
  OR2_X1 U2773 ( .A1(n2939), .A2(n2938), .ZN(n4344) );
  NAND2_X1 U2774 ( .A1(n2354), .A2(n2351), .ZN(n3701) );
  INV_X1 U2775 ( .A(n2353), .ZN(n2351) );
  OR2_X1 U2776 ( .A1(n2939), .A2(n2933), .ZN(n3728) );
  INV_X1 U2777 ( .A(n3745), .ZN(n4355) );
  OR2_X1 U2778 ( .A1(n2939), .A2(n2918), .ZN(n3745) );
  INV_X1 U2779 ( .A(n4360), .ZN(n3743) );
  INV_X1 U2780 ( .A(n3729), .ZN(n4011) );
  AND3_X1 U2781 ( .A1(n2651), .A2(n2650), .A3(n2649), .ZN(n2652) );
  NAND2_X1 U2782 ( .A1(n2644), .A2(n2643), .ZN(n3915) );
  AND3_X1 U2783 ( .A1(n2642), .A2(n2641), .A3(n2640), .ZN(n2643) );
  AND3_X1 U2784 ( .A1(n2636), .A2(n2635), .A3(n2634), .ZN(n2637) );
  INV_X1 U2785 ( .A(n4089), .ZN(n4047) );
  OAI211_X1 U2786 ( .C1(n2614), .C2(n4106), .A(n2613), .B(n2612), .ZN(n4086)
         );
  OR2_X1 U2787 ( .A1(n4105), .A2(n2431), .ZN(n2613) );
  INV_X1 U2788 ( .A(n4244), .ZN(n3917) );
  INV_X1 U2789 ( .A(n3426), .ZN(n3922) );
  NAND4_X1 U2790 ( .A1(n2495), .A2(n2494), .A3(n2493), .A4(n2492), .ZN(n4511)
         );
  OR2_X1 U2791 ( .A1(n2431), .A2(n3332), .ZN(n2494) );
  NAND4_X1 U2792 ( .A1(n2482), .A2(n2481), .A3(n2480), .A4(n2479), .ZN(n3923)
         );
  NAND4_X1 U2793 ( .A1(n2464), .A2(n2463), .A3(n2462), .A4(n2461), .ZN(n3924)
         );
  NAND4_X1 U2794 ( .A1(n2457), .A2(n2456), .A3(n2455), .A4(n2454), .ZN(n3925)
         );
  NAND4_X1 U2795 ( .A1(n2439), .A2(n2438), .A3(n2437), .A4(n2436), .ZN(n3926)
         );
  CLKBUF_X2 U2796 ( .A(U4043), .Z(n3928) );
  NAND2_X1 U2797 ( .A1(n3934), .A2(n2263), .ZN(n3052) );
  AND2_X1 U2798 ( .A1(n3051), .A2(n2264), .ZN(n2263) );
  NAND2_X1 U2799 ( .A1(n4386), .A2(n2774), .ZN(n4399) );
  NAND2_X1 U2800 ( .A1(n4406), .A2(n2777), .ZN(n4417) );
  XNOR2_X1 U2801 ( .A(n2780), .B(n2779), .ZN(n4428) );
  AND2_X1 U2802 ( .A1(n4366), .A2(n3907), .ZN(n4456) );
  XNOR2_X1 U2803 ( .A(n2822), .B(n2783), .ZN(n4451) );
  NAND2_X1 U2804 ( .A1(n4445), .A2(n2785), .ZN(n4458) );
  XNOR2_X1 U2805 ( .A(n2827), .B(n4560), .ZN(n4474) );
  NAND2_X1 U2806 ( .A1(n4482), .A2(n4483), .ZN(n4481) );
  NOR2_X1 U2807 ( .A1(n4468), .A2(n2787), .ZN(n4478) );
  XNOR2_X1 U2808 ( .A(n2790), .B(n2831), .ZN(n4488) );
  AND2_X1 U2809 ( .A1(n2841), .A2(n2840), .ZN(n4501) );
  NAND2_X1 U2810 ( .A1(n4497), .A2(n2793), .ZN(n2796) );
  NOR2_X1 U2811 ( .A1(n2796), .A2(n2797), .ZN(n3944) );
  NAND2_X1 U2812 ( .A1(n2283), .A2(n2281), .ZN(n2676) );
  INV_X1 U2813 ( .A(n2282), .ZN(n2281) );
  NAND2_X1 U2814 ( .A1(n2654), .A2(n2284), .ZN(n2283) );
  NAND2_X1 U2815 ( .A1(n2654), .A2(n2653), .ZN(n3989) );
  NOR2_X1 U2816 ( .A1(n4080), .A2(n2625), .ZN(n4060) );
  NAND2_X1 U2817 ( .A1(n4164), .A2(n2587), .ZN(n4153) );
  AND4_X1 U2818 ( .A1(n2530), .A2(n2529), .A3(n2528), .A4(n2527), .ZN(n4268)
         );
  AND4_X1 U2819 ( .A1(n2514), .A2(n2513), .A3(n2512), .A4(n2511), .ZN(n4513)
         );
  NOR2_X1 U2820 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .ZN(n2301)
         );
  XNOR2_X1 U2821 ( .A(n2737), .B(IR_REG_26__SCAN_IN), .ZN(n4336) );
  AND2_X1 U2822 ( .A1(n2928), .A2(STATE_REG_SCAN_IN), .ZN(n4554) );
  NAND2_X1 U2823 ( .A1(n2682), .A2(n2598), .ZN(n3954) );
  MUX2_X1 U2824 ( .A(IR_REG_31__SCAN_IN), .B(n2383), .S(IR_REG_1__SCAN_IN), 
        .Z(n2385) );
  AOI21_X1 U2825 ( .B1(n4361), .B2(n4548), .A(n2274), .ZN(n2273) );
  OAI22_X1 U2826 ( .A1(n4182), .A2(n2275), .B1(n2222), .B2(n4362), .ZN(n2274)
         );
  INV_X1 U2827 ( .A(REG2_REG_30__SCAN_IN), .ZN(n2275) );
  NAND2_X1 U2828 ( .A1(n2258), .A2(n2359), .ZN(U3547) );
  OR2_X1 U2829 ( .A1(n3980), .A2(n4619), .ZN(n2858) );
  OR2_X1 U2830 ( .A1(n3980), .A2(n4580), .ZN(n2862) );
  NAND2_X1 U2831 ( .A1(n4011), .A2(n4000), .ZN(n2662) );
  INV_X1 U2832 ( .A(n2419), .ZN(n2522) );
  INV_X2 U2833 ( .A(n2522), .ZN(n3767) );
  NAND4_X1 U2834 ( .A1(n2415), .A2(n2414), .A3(n2413), .A4(n2412), .ZN(n2874)
         );
  INV_X1 U2835 ( .A(n2892), .ZN(n3564) );
  AND4_X1 U2836 ( .A1(n2400), .A2(n2399), .A3(n2398), .A4(n2397), .ZN(n2894)
         );
  INV_X2 U2837 ( .A(n3564), .ZN(n3602) );
  AND2_X1 U2838 ( .A1(n4335), .A2(REG3_REG_1__SCAN_IN), .ZN(n2226) );
  AND2_X1 U2839 ( .A1(n2424), .A2(n2370), .ZN(n2227) );
  INV_X1 U2840 ( .A(IR_REG_28__SCAN_IN), .ZN(n4906) );
  INV_X1 U2841 ( .A(n3713), .ZN(n2335) );
  AND2_X1 U2842 ( .A1(n3540), .A2(n3539), .ZN(n3713) );
  INV_X1 U2843 ( .A(n4067), .ZN(n2624) );
  INV_X1 U2844 ( .A(n2431), .ZN(n2666) );
  INV_X1 U2845 ( .A(n2358), .ZN(n2440) );
  AND2_X1 U2846 ( .A1(n2354), .A2(n2352), .ZN(n2228) );
  AND2_X1 U2847 ( .A1(n2381), .A2(n3012), .ZN(n2419) );
  NAND2_X1 U2848 ( .A1(n2320), .A2(n2325), .ZN(n3622) );
  XNOR2_X1 U2849 ( .A(n2681), .B(n2680), .ZN(n2721) );
  OR2_X1 U2850 ( .A1(n2920), .A2(n2924), .ZN(n2229) );
  NOR2_X1 U2851 ( .A1(n2291), .A2(n3793), .ZN(n2230) );
  AND2_X1 U2852 ( .A1(n2723), .A2(n2722), .ZN(n2231) );
  NAND2_X1 U2853 ( .A1(n3924), .A2(n3296), .ZN(n2232) );
  NOR2_X1 U2854 ( .A1(n4478), .A2(n4477), .ZN(n2233) );
  AND2_X1 U2855 ( .A1(n4533), .A2(n3154), .ZN(n2234) );
  NAND2_X1 U2856 ( .A1(n2618), .A2(n2617), .ZN(n4079) );
  INV_X1 U2857 ( .A(n2348), .ZN(n2347) );
  NAND2_X1 U2858 ( .A1(n3572), .A2(n2349), .ZN(n2348) );
  AND2_X1 U2859 ( .A1(n2378), .A2(n2714), .ZN(n2235) );
  INV_X1 U2860 ( .A(n3768), .ZN(n2614) );
  NOR2_X1 U2861 ( .A1(n3529), .A2(n3528), .ZN(n3734) );
  INV_X1 U2862 ( .A(n3611), .ZN(n2331) );
  XNOR2_X1 U2863 ( .A(n2735), .B(n2734), .ZN(n2740) );
  NOR2_X1 U2864 ( .A1(n3709), .A2(n3713), .ZN(n2236) );
  AOI21_X1 U2865 ( .B1(n4515), .B2(n4514), .A(n2510), .ZN(n3365) );
  OR2_X1 U2866 ( .A1(n3814), .A2(n2295), .ZN(n2237) );
  NAND2_X1 U2867 ( .A1(n2731), .A2(IR_REG_31__SCAN_IN), .ZN(n2741) );
  NAND2_X1 U2868 ( .A1(n2337), .A2(n2341), .ZN(n3519) );
  INV_X1 U2869 ( .A(n3659), .ZN(n2329) );
  NAND2_X1 U2870 ( .A1(n3692), .A2(n3693), .ZN(n3690) );
  INV_X1 U2871 ( .A(n3425), .ZN(n3371) );
  NAND2_X1 U2872 ( .A1(n2296), .A2(n2586), .ZN(n4164) );
  NAND2_X1 U2873 ( .A1(n2298), .A2(n2550), .ZN(n3489) );
  NOR2_X1 U2874 ( .A1(n4168), .A2(n4154), .ZN(n2278) );
  AND2_X1 U2875 ( .A1(n2342), .A2(n3518), .ZN(n2238) );
  NAND2_X1 U2876 ( .A1(n2344), .A2(n2347), .ZN(n3628) );
  INV_X1 U2877 ( .A(n3562), .ZN(n2355) );
  AND2_X1 U2878 ( .A1(n3711), .A2(n2335), .ZN(n2239) );
  AND2_X1 U2879 ( .A1(n2969), .A2(n2968), .ZN(n2240) );
  NAND2_X1 U2880 ( .A1(n3599), .A2(n3598), .ZN(n2241) );
  NOR2_X1 U2881 ( .A1(n4086), .A2(n4110), .ZN(n2616) );
  AND2_X1 U2882 ( .A1(n2336), .A2(n3544), .ZN(n2242) );
  NAND2_X1 U2883 ( .A1(n3461), .A2(n4266), .ZN(n3460) );
  AND2_X1 U2884 ( .A1(n3605), .A2(n3604), .ZN(n2243) );
  INV_X1 U2885 ( .A(n2352), .ZN(n2350) );
  NOR2_X1 U2886 ( .A1(n3702), .A2(n2353), .ZN(n2352) );
  AND2_X1 U2887 ( .A1(n2364), .A2(n3582), .ZN(n2244) );
  NAND2_X1 U2888 ( .A1(n3729), .A2(n4197), .ZN(n2245) );
  AND2_X1 U2889 ( .A1(n3877), .A2(n3874), .ZN(n3490) );
  INV_X1 U2890 ( .A(n3490), .ZN(n2561) );
  OAI22_X1 U2891 ( .A1(n3287), .A2(n2489), .B1(n3324), .B2(n3338), .ZN(n3320)
         );
  OAI21_X1 U2892 ( .B1(n3384), .B2(n3383), .A(n3382), .ZN(n3437) );
  NAND2_X1 U2893 ( .A1(n3095), .A2(n2959), .ZN(n3121) );
  NAND2_X1 U2894 ( .A1(n2303), .A2(n2302), .ZN(n3224) );
  NAND2_X1 U2895 ( .A1(n2304), .A2(n2308), .ZN(n3188) );
  INV_X1 U2896 ( .A(n3518), .ZN(n2340) );
  AOI21_X1 U2897 ( .B1(n2995), .B2(n2994), .A(n2365), .ZN(n3352) );
  NAND2_X1 U2898 ( .A1(n2300), .A2(n2229), .ZN(n2246) );
  NOR2_X1 U2899 ( .A1(n2571), .A2(n2570), .ZN(n2584) );
  AND4_X1 U2900 ( .A1(n2406), .A2(n2405), .A3(n2404), .A4(n2403), .ZN(n4536)
         );
  XNOR2_X1 U2901 ( .A(n2879), .B(n2880), .ZN(n3085) );
  INV_X1 U2902 ( .A(n2789), .ZN(n2262) );
  AND2_X1 U2903 ( .A1(n2829), .A2(REG2_REG_15__SCAN_IN), .ZN(n2789) );
  INV_X1 U2904 ( .A(IR_REG_14__SCAN_IN), .ZN(n2376) );
  INV_X1 U2905 ( .A(IR_REG_1__SCAN_IN), .ZN(n2267) );
  INV_X1 U2906 ( .A(IR_REG_0__SCAN_IN), .ZN(n2266) );
  NAND2_X1 U2907 ( .A1(n2249), .A2(n3828), .ZN(n4539) );
  AND2_X1 U2908 ( .A1(n3064), .A2(n3154), .ZN(n3828) );
  OAI21_X2 U2909 ( .B1(n3236), .B2(n2696), .A(n3850), .ZN(n3295) );
  NAND2_X1 U2910 ( .A1(n2253), .A2(n2235), .ZN(n2299) );
  INV_X1 U2911 ( .A(n2727), .ZN(n2253) );
  NAND2_X1 U2912 ( .A1(n2716), .A2(n2301), .ZN(n3619) );
  NAND4_X1 U2913 ( .A1(n2257), .A2(n2256), .A3(n2255), .A4(n2254), .ZN(n2371)
         );
  NAND2_X1 U2914 ( .A1(n3409), .A2(n3863), .ZN(n2698) );
  NAND2_X1 U2915 ( .A1(n4509), .A2(n3861), .ZN(n2259) );
  NAND2_X1 U2916 ( .A1(n2883), .A2(n4533), .ZN(n2885) );
  NAND4_X1 U2917 ( .A1(n2396), .A2(n2394), .A3(n2393), .A4(n2395), .ZN(n4533)
         );
  NAND2_X1 U2918 ( .A1(n2221), .A2(REG2_REG_2__SCAN_IN), .ZN(n2265) );
  AND2_X2 U2919 ( .A1(n2267), .A2(n2266), .ZN(n2407) );
  NAND4_X1 U2920 ( .A1(n2269), .A2(n2358), .A3(n4753), .A4(n2357), .ZN(n2727)
         );
  AND2_X2 U2921 ( .A1(n2268), .A2(n2227), .ZN(n2358) );
  NAND3_X1 U2922 ( .A1(n2272), .A2(n2271), .A3(n2270), .ZN(n2377) );
  NAND3_X1 U2923 ( .A1(n2376), .A2(n4887), .A3(n2557), .ZN(n2570) );
  INV_X1 U2924 ( .A(n2273), .ZN(U3261) );
  AOI21_X1 U2925 ( .B1(n4193), .B2(n4190), .A(n4189), .ZN(n4361) );
  NOR2_X2 U2926 ( .A1(n4190), .A2(n4193), .ZN(n4189) );
  INV_X1 U2927 ( .A(n2278), .ZN(n4156) );
  INV_X1 U2928 ( .A(n4163), .ZN(n2296) );
  NAND2_X1 U2929 ( .A1(n2298), .A2(n2297), .ZN(n3492) );
  NAND2_X1 U2930 ( .A1(n2922), .A2(n2921), .ZN(n2300) );
  NAND3_X1 U2931 ( .A1(n2300), .A2(n2229), .A3(n2951), .ZN(n3097) );
  NAND2_X1 U2932 ( .A1(n3121), .A2(n2305), .ZN(n2303) );
  NAND2_X1 U2933 ( .A1(n3658), .A2(n2317), .ZN(n2312) );
  OAI211_X1 U2934 ( .C1(n3658), .C2(n2318), .A(n2312), .B(n2313), .ZN(n3618)
         );
  NAND2_X1 U2935 ( .A1(n3658), .A2(n2328), .ZN(n2320) );
  AOI21_X1 U2936 ( .B1(n3658), .B2(n3659), .A(n3660), .ZN(n3722) );
  NAND2_X1 U2937 ( .A1(n3651), .A2(n2352), .ZN(n2344) );
  OAI21_X1 U2938 ( .B1(n3651), .B2(n2348), .A(n2345), .ZN(n3583) );
  NOR2_X1 U2939 ( .A1(n2571), .A2(n2377), .ZN(n2724) );
  NOR2_X1 U2940 ( .A1(n2440), .A2(n2371), .ZN(n2531) );
  NOR2_X1 U2941 ( .A1(n3211), .A2(n2468), .ZN(n2475) );
  OAI21_X1 U2942 ( .B1(n3133), .B2(n2443), .A(n2442), .ZN(n3211) );
  OR2_X1 U2943 ( .A1(n2225), .A2(n3075), .ZN(n2395) );
  NAND2_X1 U2944 ( .A1(n3768), .A2(REG2_REG_0__SCAN_IN), .ZN(n2396) );
  INV_X1 U2945 ( .A(n2740), .ZN(n2757) );
  OR2_X1 U2946 ( .A1(n2571), .A2(IR_REG_14__SCAN_IN), .ZN(n2548) );
  INV_X1 U2947 ( .A(n2870), .ZN(n3927) );
  NAND2_X2 U2948 ( .A1(n2390), .A2(n2389), .ZN(n2428) );
  NAND2_X1 U2949 ( .A1(n2882), .A2(n2907), .ZN(n2920) );
  INV_X1 U2950 ( .A(n3199), .ZN(n3204) );
  INV_X1 U2951 ( .A(n2810), .ZN(n2772) );
  INV_X1 U2952 ( .A(n4403), .ZN(n2814) );
  INV_X1 U2953 ( .A(n4424), .ZN(n2779) );
  OR2_X1 U2954 ( .A1(n3971), .A2(n4619), .ZN(n2359) );
  OR2_X1 U2955 ( .A1(n3971), .A2(n4580), .ZN(n2360) );
  OR2_X1 U2956 ( .A1(n4613), .A2(n2760), .ZN(n2361) );
  AND2_X1 U2957 ( .A1(n4050), .A2(n3587), .ZN(n2362) );
  NAND2_X1 U2958 ( .A1(n3915), .A2(n4032), .ZN(n2363) );
  XNOR2_X1 U2959 ( .A(n2895), .B(n2896), .ZN(n3066) );
  OR2_X1 U2960 ( .A1(n3576), .A2(n3575), .ZN(n2364) );
  OAI22_X1 U2961 ( .A1(n3104), .A2(n2417), .B1(n3833), .B2(n3091), .ZN(n3197)
         );
  INV_X1 U2962 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2476) );
  NOR2_X1 U2963 ( .A1(n2998), .A2(n2993), .ZN(n2365) );
  INV_X1 U2964 ( .A(IR_REG_17__SCAN_IN), .ZN(n2583) );
  OR2_X1 U2965 ( .A1(n4198), .A2(n4014), .ZN(n2367) );
  NAND2_X1 U2966 ( .A1(n3067), .A2(n2898), .ZN(n3077) );
  AND3_X1 U2967 ( .A1(n3786), .A2(n2549), .A3(n3452), .ZN(n2368) );
  INV_X1 U2968 ( .A(IR_REG_4__SCAN_IN), .ZN(n2370) );
  AND2_X1 U2969 ( .A1(n3408), .A2(n3410), .ZN(n3863) );
  NAND2_X1 U2970 ( .A1(n2409), .A2(n3171), .ZN(n3830) );
  NAND2_X1 U2971 ( .A1(n2874), .A2(n3564), .ZN(n2876) );
  INV_X1 U2972 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2760) );
  OR2_X1 U2973 ( .A1(n2471), .A2(n3242), .ZN(n3291) );
  INV_X1 U2974 ( .A(IR_REG_2__SCAN_IN), .ZN(n2369) );
  NOR2_X1 U2975 ( .A1(n3629), .A2(n3630), .ZN(n3572) );
  OAI22_X1 U2976 ( .A1(n2894), .A2(n3606), .B1(n2892), .B2(n4545), .ZN(n2896)
         );
  INV_X1 U2977 ( .A(n3581), .ZN(n3582) );
  AND2_X1 U2978 ( .A1(n3381), .A2(n3398), .ZN(n3382) );
  INV_X1 U2979 ( .A(n2821), .ZN(n2783) );
  INV_X1 U2980 ( .A(n4172), .ZN(n2586) );
  INV_X1 U2981 ( .A(IR_REG_26__SCAN_IN), .ZN(n2378) );
  INV_X1 U2982 ( .A(IR_REG_15__SCAN_IN), .ZN(n2557) );
  INV_X1 U2983 ( .A(IR_REG_24__SCAN_IN), .ZN(n2734) );
  OAI22_X1 U2984 ( .A1(n2870), .A2(n2892), .B1(n2899), .B2(n3204), .ZN(n2873)
         );
  NAND2_X1 U2985 ( .A1(n2806), .A2(n4339), .ZN(n2807) );
  NOR2_X1 U2986 ( .A1(n2624), .A2(n4091), .ZN(n2625) );
  NAND2_X1 U2987 ( .A1(n2453), .A2(REG3_REG_6__SCAN_IN), .ZN(n2452) );
  INV_X1 U2988 ( .A(n2428), .ZN(n2794) );
  INV_X1 U2989 ( .A(n2690), .ZN(n3162) );
  AND2_X1 U2990 ( .A1(n2487), .A2(n2486), .ZN(n2497) );
  NOR2_X1 U2991 ( .A1(n2756), .A2(n3008), .ZN(n2739) );
  INV_X1 U2992 ( .A(n3832), .ZN(n3091) );
  AND2_X1 U2993 ( .A1(n2977), .A2(n2978), .ZN(n3225) );
  NOR2_X1 U2994 ( .A1(n2490), .A2(n4973), .ZN(n2501) );
  AND2_X1 U2995 ( .A1(n2542), .A2(REG3_REG_15__SCAN_IN), .ZN(n2551) );
  XNOR2_X1 U2996 ( .A(n2900), .B(n3607), .ZN(n2903) );
  AND2_X1 U2997 ( .A1(n2647), .A2(n2646), .ZN(n2655) );
  INV_X1 U2998 ( .A(n3639), .ZN(n4074) );
  NAND2_X1 U2999 ( .A1(n3768), .A2(REG2_REG_3__SCAN_IN), .ZN(n2415) );
  OAI21_X1 U3000 ( .B1(n4508), .B2(n4556), .A(n2843), .ZN(n2844) );
  AND2_X1 U3001 ( .A1(n3942), .A2(REG2_REG_18__SCAN_IN), .ZN(n3943) );
  INV_X1 U3002 ( .A(n2662), .ZN(n2663) );
  INV_X1 U3003 ( .A(n3214), .ZN(n3257) );
  OR2_X1 U3004 ( .A1(n3146), .A2(n2936), .ZN(n4129) );
  INV_X1 U3005 ( .A(n3587), .ZN(n4032) );
  INV_X1 U3006 ( .A(n3644), .ZN(n4154) );
  INV_X1 U3007 ( .A(n4336), .ZN(n2756) );
  XNOR2_X1 U3008 ( .A(n2967), .B(n2968), .ZN(n3189) );
  OR2_X1 U3009 ( .A1(n2608), .A2(n3653), .ZN(n2619) );
  INV_X1 U3010 ( .A(n3728), .ZN(n4350) );
  NAND2_X1 U3011 ( .A1(n2600), .A2(REG3_REG_20__SCAN_IN), .ZN(n2608) );
  OR2_X1 U3012 ( .A1(n2664), .A2(n3612), .ZN(n3970) );
  AOI21_X1 U3013 ( .B1(n4074), .B2(n2666), .A(n2631), .ZN(n4089) );
  INV_X1 U3014 ( .A(n2965), .ZN(n3126) );
  NAND2_X1 U3015 ( .A1(n4451), .A2(REG1_REG_12__SCAN_IN), .ZN(n4450) );
  AND2_X1 U3016 ( .A1(n2841), .A2(n2839), .ZN(n4366) );
  AND2_X1 U3017 ( .A1(n4366), .A2(n3030), .ZN(n4502) );
  AND2_X1 U3018 ( .A1(n4141), .A2(n4142), .ZN(n4172) );
  AND2_X1 U3019 ( .A1(n4182), .A2(n4530), .ZN(n4111) );
  INV_X1 U3020 ( .A(n4186), .ZN(n4161) );
  INV_X1 U3021 ( .A(n4159), .ZN(n4548) );
  NAND2_X1 U3022 ( .A1(n4631), .A2(n2864), .ZN(n2865) );
  AND2_X1 U3023 ( .A1(n2758), .A2(n3015), .ZN(n2912) );
  INV_X1 U3024 ( .A(n3513), .ZN(n4243) );
  NAND2_X1 U3025 ( .A1(n4516), .A2(n4607), .ZN(n4590) );
  AND2_X1 U3026 ( .A1(n3156), .A2(n2871), .ZN(n4601) );
  AND2_X1 U3027 ( .A1(n2932), .A2(n3061), .ZN(n4360) );
  INV_X1 U3028 ( .A(n3966), .ZN(n3987) );
  OAI211_X1 U3029 ( .C1(n4092), .C2(n2431), .A(n2622), .B(n2621), .ZN(n4067)
         );
  INV_X1 U3030 ( .A(n4258), .ZN(n3919) );
  NAND2_X1 U3031 ( .A1(n2846), .A2(n2845), .ZN(n2847) );
  NAND2_X1 U3032 ( .A1(n4182), .A2(n3164), .ZN(n4159) );
  NAND2_X1 U3033 ( .A1(n4634), .A2(n4169), .ZN(n4619) );
  INV_X1 U3034 ( .A(n4634), .ZN(n4631) );
  AND2_X1 U3035 ( .A1(n2360), .A2(n2361), .ZN(n2761) );
  NAND2_X1 U3036 ( .A1(n4613), .A2(n4169), .ZN(n4580) );
  INV_X1 U3037 ( .A(n4613), .ZN(n4611) );
  INV_X1 U3038 ( .A(n4552), .ZN(n4553) );
  INV_X1 U3039 ( .A(n2824), .ZN(n4561) );
  OR2_X1 U3040 ( .A1(n2848), .A2(n2847), .ZN(U3258) );
  NAND2_X1 U3041 ( .A1(n2407), .A2(n2369), .ZN(n2416) );
  NOR2_X1 U3042 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2375)
         );
  NOR2_X1 U3043 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2374)
         );
  NOR2_X1 U3044 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2373)
         );
  NOR2_X1 U3045 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2372)
         );
  INV_X1 U3046 ( .A(IR_REG_30__SCAN_IN), .ZN(n3620) );
  INV_X2 U3047 ( .A(n2381), .ZN(n4335) );
  INV_X1 U3048 ( .A(IR_REG_29__SCAN_IN), .ZN(n4720) );
  AND2_X4 U3049 ( .A1(n4335), .A2(n2382), .ZN(n3768) );
  NAND2_X1 U3050 ( .A1(n2418), .A2(REG0_REG_1__SCAN_IN), .ZN(n2397) );
  INV_X1 U3051 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3071) );
  NAND4_X1 U3052 ( .A1(n2400), .A2(n2399), .A3(n2397), .A4(n2398), .ZN(n2391)
         );
  NAND2_X1 U3053 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2383)
         );
  INV_X1 U3054 ( .A(n2407), .ZN(n2384) );
  INV_X1 U3055 ( .A(n3005), .ZN(n3929) );
  NAND2_X1 U3056 ( .A1(n2715), .A2(IR_REG_28__SCAN_IN), .ZN(n2386) );
  INV_X1 U3057 ( .A(IR_REG_27__SCAN_IN), .ZN(n2714) );
  NAND2_X1 U3058 ( .A1(n2386), .A2(IR_REG_27__SCAN_IN), .ZN(n2390) );
  NAND2_X1 U3059 ( .A1(n2387), .A2(n4906), .ZN(n2388) );
  MUX2_X1 U3060 ( .A(n3929), .B(DATAI_1_), .S(n2428), .Z(n4531) );
  NAND2_X1 U3061 ( .A1(n2391), .A2(n4545), .ZN(n3826) );
  NAND4_X1 U3062 ( .A1(n2392), .A2(n2397), .A3(n2399), .A4(n2400), .ZN(n2689)
         );
  NAND2_X1 U3063 ( .A1(n3826), .A2(n2689), .ZN(n2688) );
  INV_X1 U3064 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3075) );
  NAND2_X1 U3065 ( .A1(n2419), .A2(REG1_REG_0__SCAN_IN), .ZN(n2394) );
  NAND2_X1 U3066 ( .A1(n2418), .A2(REG0_REG_0__SCAN_IN), .ZN(n2393) );
  MUX2_X1 U3067 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2428), .Z(n3154) );
  NAND2_X1 U3068 ( .A1(n2688), .A2(n2234), .ZN(n4529) );
  INV_X1 U3069 ( .A(n2894), .ZN(n2401) );
  NAND2_X1 U3070 ( .A1(n2401), .A2(n4531), .ZN(n2402) );
  NAND2_X1 U3071 ( .A1(n4529), .A2(n2402), .ZN(n3161) );
  INV_X1 U3072 ( .A(n3161), .ZN(n2410) );
  NAND2_X1 U3073 ( .A1(n3768), .A2(REG2_REG_2__SCAN_IN), .ZN(n2406) );
  NAND2_X1 U3074 ( .A1(n2419), .A2(REG1_REG_2__SCAN_IN), .ZN(n2405) );
  NAND2_X1 U3075 ( .A1(n2418), .A2(REG0_REG_2__SCAN_IN), .ZN(n2404) );
  INV_X1 U3076 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3168) );
  OR2_X1 U3077 ( .A1(n2224), .A2(n3168), .ZN(n2403) );
  INV_X1 U3078 ( .A(n4536), .ZN(n2409) );
  MUX2_X1 U3079 ( .A(n2221), .B(DATAI_2_), .S(n2428), .Z(n3165) );
  INV_X1 U3080 ( .A(n3165), .ZN(n3171) );
  NAND2_X1 U3081 ( .A1(n4536), .A2(n3165), .ZN(n2692) );
  NAND2_X1 U3082 ( .A1(n3830), .A2(n2692), .ZN(n2690) );
  NAND2_X1 U3083 ( .A1(n2410), .A2(n2690), .ZN(n3160) );
  NAND2_X1 U3084 ( .A1(n4536), .A2(n3171), .ZN(n2411) );
  NAND2_X1 U3085 ( .A1(n3160), .A2(n2411), .ZN(n3104) );
  NAND2_X1 U3086 ( .A1(n3767), .A2(REG1_REG_3__SCAN_IN), .ZN(n2414) );
  NAND2_X1 U3087 ( .A1(n2418), .A2(REG0_REG_3__SCAN_IN), .ZN(n2413) );
  OR2_X1 U3088 ( .A1(n2431), .A2(REG3_REG_3__SCAN_IN), .ZN(n2412) );
  NAND2_X1 U3089 ( .A1(n2416), .A2(IR_REG_31__SCAN_IN), .ZN(n2425) );
  XNOR2_X1 U3090 ( .A(n2425), .B(IR_REG_3__SCAN_IN), .ZN(n4340) );
  MUX2_X1 U3091 ( .A(n4340), .B(DATAI_3_), .S(n2428), .Z(n3832) );
  NOR2_X1 U3092 ( .A1(n2874), .A2(n3832), .ZN(n2417) );
  INV_X1 U3093 ( .A(n2874), .ZN(n3833) );
  NAND2_X1 U3094 ( .A1(n2418), .A2(REG0_REG_4__SCAN_IN), .ZN(n2423) );
  NAND2_X1 U3095 ( .A1(n2673), .A2(REG1_REG_4__SCAN_IN), .ZN(n2422) );
  NAND2_X1 U3096 ( .A1(n3768), .A2(REG2_REG_4__SCAN_IN), .ZN(n2421) );
  XNOR2_X1 U3097 ( .A(REG3_REG_4__SCAN_IN), .B(REG3_REG_3__SCAN_IN), .ZN(n3206) );
  OR2_X1 U3098 ( .A1(n2431), .A2(n3206), .ZN(n2420) );
  NAND2_X1 U3099 ( .A1(n2425), .A2(n2424), .ZN(n2426) );
  NAND2_X1 U3100 ( .A1(n2426), .A2(IR_REG_31__SCAN_IN), .ZN(n2427) );
  XNOR2_X1 U3101 ( .A(n2427), .B(IR_REG_4__SCAN_IN), .ZN(n4339) );
  INV_X4 U3102 ( .A(n2794), .ZN(n3772) );
  MUX2_X1 U3103 ( .A(n4339), .B(DATAI_4_), .S(n3772), .Z(n3199) );
  NAND2_X1 U3104 ( .A1(n2870), .A2(n3199), .ZN(n3835) );
  NAND2_X1 U3105 ( .A1(n3927), .A2(n3204), .ZN(n3838) );
  NAND2_X1 U3106 ( .A1(n3197), .A2(n3784), .ZN(n2430) );
  NAND2_X1 U3107 ( .A1(n3927), .A2(n3199), .ZN(n2429) );
  NAND2_X1 U3108 ( .A1(n2430), .A2(n2429), .ZN(n3133) );
  INV_X1 U3109 ( .A(n2453), .ZN(n2435) );
  INV_X1 U3110 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2433) );
  NAND2_X1 U3111 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2432) );
  NAND2_X1 U3112 ( .A1(n2433), .A2(n2432), .ZN(n2434) );
  NAND2_X1 U3113 ( .A1(n2435), .A2(n2434), .ZN(n3268) );
  OR2_X1 U3114 ( .A1(n2431), .A2(n3268), .ZN(n2439) );
  NAND2_X1 U3115 ( .A1(n2673), .A2(REG1_REG_5__SCAN_IN), .ZN(n2438) );
  NAND2_X1 U3116 ( .A1(n3768), .A2(REG2_REG_5__SCAN_IN), .ZN(n2437) );
  NAND2_X1 U3117 ( .A1(n2418), .A2(REG0_REG_5__SCAN_IN), .ZN(n2436) );
  NAND2_X1 U3118 ( .A1(n2440), .A2(IR_REG_31__SCAN_IN), .ZN(n2441) );
  XNOR2_X1 U3119 ( .A(n2441), .B(IR_REG_5__SCAN_IN), .ZN(n2809) );
  MUX2_X1 U3120 ( .A(n2809), .B(DATAI_5_), .S(n3772), .Z(n3269) );
  AND2_X1 U3121 ( .A1(n3926), .A2(n3269), .ZN(n2443) );
  INV_X1 U3122 ( .A(n3926), .ZN(n3256) );
  INV_X1 U3123 ( .A(n3269), .ZN(n3098) );
  NAND2_X1 U3124 ( .A1(n3256), .A2(n3098), .ZN(n2442) );
  NAND2_X1 U3125 ( .A1(n2418), .A2(REG0_REG_7__SCAN_IN), .ZN(n2449) );
  NAND2_X1 U3126 ( .A1(n2673), .A2(REG1_REG_7__SCAN_IN), .ZN(n2448) );
  NAND2_X1 U3127 ( .A1(n3768), .A2(REG2_REG_7__SCAN_IN), .ZN(n2447) );
  AND2_X1 U3128 ( .A1(n2452), .A2(n2444), .ZN(n2445) );
  OR2_X1 U3129 ( .A1(n2445), .A2(n2459), .ZN(n3248) );
  OR2_X1 U3130 ( .A1(n2431), .A2(n3248), .ZN(n2446) );
  NAND2_X1 U3131 ( .A1(n2487), .A2(n2485), .ZN(n2450) );
  NAND2_X1 U3132 ( .A1(n2450), .A2(IR_REG_31__SCAN_IN), .ZN(n2465) );
  XNOR2_X1 U3133 ( .A(n2465), .B(IR_REG_7__SCAN_IN), .ZN(n2813) );
  MUX2_X1 U3134 ( .A(n2813), .B(DATAI_7_), .S(n3772), .Z(n3238) );
  INV_X1 U3135 ( .A(n3238), .ZN(n3192) );
  NAND2_X1 U3136 ( .A1(n2965), .A2(n3238), .ZN(n3841) );
  NAND2_X1 U3137 ( .A1(n3126), .A2(n3238), .ZN(n2469) );
  INV_X1 U3138 ( .A(n2469), .ZN(n2451) );
  NOR2_X1 U3139 ( .A1(n3785), .A2(n2451), .ZN(n2471) );
  NAND2_X1 U3140 ( .A1(n2418), .A2(REG0_REG_6__SCAN_IN), .ZN(n2457) );
  OAI21_X1 U3141 ( .B1(n2453), .B2(REG3_REG_6__SCAN_IN), .A(n2452), .ZN(n3254)
         );
  OR2_X1 U3142 ( .A1(n2431), .A2(n3254), .ZN(n2456) );
  NAND2_X1 U3143 ( .A1(n3767), .A2(REG1_REG_6__SCAN_IN), .ZN(n2455) );
  NAND2_X1 U3144 ( .A1(n3768), .A2(REG2_REG_6__SCAN_IN), .ZN(n2454) );
  OR2_X1 U3145 ( .A1(n2487), .A2(n2732), .ZN(n2458) );
  XNOR2_X1 U3146 ( .A(n2458), .B(IR_REG_6__SCAN_IN), .ZN(n2810) );
  MUX2_X1 U3147 ( .A(n2810), .B(DATAI_6_), .S(n3772), .Z(n3214) );
  NOR2_X1 U31480 ( .A1(n3925), .A2(n3214), .ZN(n3242) );
  NAND2_X1 U31490 ( .A1(n2418), .A2(REG0_REG_8__SCAN_IN), .ZN(n2464) );
  OR2_X1 U3150 ( .A1(n2459), .A2(REG3_REG_8__SCAN_IN), .ZN(n2460) );
  NAND2_X1 U3151 ( .A1(n2477), .A2(n2460), .ZN(n3304) );
  OR2_X1 U3152 ( .A1(n2431), .A2(n3304), .ZN(n2463) );
  NAND2_X1 U3153 ( .A1(n3767), .A2(REG1_REG_8__SCAN_IN), .ZN(n2462) );
  NAND2_X1 U3154 ( .A1(n3768), .A2(REG2_REG_8__SCAN_IN), .ZN(n2461) );
  NAND2_X1 U3155 ( .A1(n2465), .A2(n2484), .ZN(n2466) );
  NAND2_X1 U3156 ( .A1(n2466), .A2(IR_REG_31__SCAN_IN), .ZN(n2467) );
  XNOR2_X1 U3157 ( .A(n2467), .B(IR_REG_8__SCAN_IN), .ZN(n4403) );
  MUX2_X1 U3158 ( .A(n4403), .B(DATAI_8_), .S(n3772), .Z(n3296) );
  INV_X1 U3159 ( .A(n3296), .ZN(n3302) );
  AND2_X1 U3160 ( .A1(n3339), .A2(n3302), .ZN(n2473) );
  OR2_X1 U3161 ( .A1(n3291), .A2(n2473), .ZN(n2468) );
  NAND2_X1 U3162 ( .A1(n3925), .A2(n3214), .ZN(n3243) );
  AND2_X1 U3163 ( .A1(n3243), .A2(n2469), .ZN(n2470) );
  NOR2_X1 U3164 ( .A1(n2473), .A2(n2472), .ZN(n2474) );
  NOR2_X1 U3165 ( .A1(n2475), .A2(n2474), .ZN(n3287) );
  NAND2_X1 U3166 ( .A1(n2673), .A2(REG1_REG_9__SCAN_IN), .ZN(n2482) );
  NAND2_X1 U3167 ( .A1(n2477), .A2(n2476), .ZN(n2478) );
  NAND2_X1 U3168 ( .A1(n2490), .A2(n2478), .ZN(n3313) );
  OR2_X1 U3169 ( .A1(n2431), .A2(n3313), .ZN(n2481) );
  NAND2_X1 U3170 ( .A1(n2672), .A2(REG0_REG_9__SCAN_IN), .ZN(n2480) );
  NAND2_X1 U3171 ( .A1(n3768), .A2(REG2_REG_9__SCAN_IN), .ZN(n2479) );
  INV_X1 U3172 ( .A(IR_REG_8__SCAN_IN), .ZN(n2483) );
  AND3_X1 U3173 ( .A1(n2485), .A2(n2484), .A3(n2483), .ZN(n2486) );
  OR2_X1 U3174 ( .A1(n2497), .A2(n2732), .ZN(n2488) );
  XNOR2_X1 U3175 ( .A(n2488), .B(IR_REG_9__SCAN_IN), .ZN(n2817) );
  MUX2_X1 U3176 ( .A(n2817), .B(DATAI_9_), .S(n3772), .Z(n3282) );
  NOR2_X1 U3177 ( .A1(n3923), .A2(n3282), .ZN(n2489) );
  NAND2_X1 U3178 ( .A1(n2672), .A2(REG0_REG_10__SCAN_IN), .ZN(n2495) );
  AND2_X1 U3179 ( .A1(n2490), .A2(n4973), .ZN(n2491) );
  OR2_X1 U3180 ( .A1(n2501), .A2(n2491), .ZN(n3332) );
  NAND2_X1 U3181 ( .A1(n3767), .A2(REG1_REG_10__SCAN_IN), .ZN(n2493) );
  NAND2_X1 U3182 ( .A1(n3768), .A2(REG2_REG_10__SCAN_IN), .ZN(n2492) );
  INV_X1 U3183 ( .A(IR_REG_9__SCAN_IN), .ZN(n2496) );
  NAND2_X1 U3184 ( .A1(n2497), .A2(n2496), .ZN(n2508) );
  NAND2_X1 U3185 ( .A1(n2508), .A2(IR_REG_31__SCAN_IN), .ZN(n2498) );
  XNOR2_X1 U3186 ( .A(n2498), .B(IR_REG_10__SCAN_IN), .ZN(n4424) );
  MUX2_X1 U3187 ( .A(n4424), .B(DATAI_10_), .S(n3772), .Z(n3322) );
  AND2_X1 U3188 ( .A1(n4511), .A2(n3322), .ZN(n2499) );
  NAND2_X1 U3189 ( .A1(n3279), .A2(n3329), .ZN(n2500) );
  NAND2_X1 U3190 ( .A1(n3767), .A2(REG1_REG_11__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U3191 ( .A1(n3768), .A2(REG2_REG_11__SCAN_IN), .ZN(n2506) );
  NAND2_X1 U3192 ( .A1(n2672), .A2(REG0_REG_11__SCAN_IN), .ZN(n2505) );
  OR2_X1 U3193 ( .A1(n2501), .A2(REG3_REG_11__SCAN_IN), .ZN(n2502) );
  AND2_X1 U3194 ( .A1(n2525), .A2(n2502), .ZN(n4521) );
  INV_X1 U3195 ( .A(n4521), .ZN(n2503) );
  OR2_X1 U3196 ( .A1(n2431), .A2(n2503), .ZN(n2504) );
  NAND2_X1 U3197 ( .A1(n2509), .A2(IR_REG_31__SCAN_IN), .ZN(n2516) );
  XNOR2_X1 U3198 ( .A(n2516), .B(IR_REG_11__SCAN_IN), .ZN(n2799) );
  MUX2_X1 U3199 ( .A(n2799), .B(DATAI_11_), .S(n3772), .Z(n4510) );
  NAND2_X1 U3200 ( .A1(n3426), .A2(n4510), .ZN(n3862) );
  INV_X1 U3201 ( .A(n4510), .ZN(n4523) );
  NAND2_X1 U3202 ( .A1(n3922), .A2(n4523), .ZN(n3861) );
  NAND2_X1 U3203 ( .A1(n3862), .A2(n3861), .ZN(n4514) );
  NOR2_X1 U3204 ( .A1(n3922), .A2(n4510), .ZN(n2510) );
  NAND2_X1 U3205 ( .A1(n2672), .A2(REG0_REG_12__SCAN_IN), .ZN(n2514) );
  NAND2_X1 U3206 ( .A1(n3767), .A2(REG1_REG_12__SCAN_IN), .ZN(n2513) );
  NAND2_X1 U3207 ( .A1(n3768), .A2(REG2_REG_12__SCAN_IN), .ZN(n2512) );
  XNOR2_X1 U3208 ( .A(n2525), .B(n2524), .ZN(n3407) );
  OR2_X1 U3209 ( .A1(n2431), .A2(n3407), .ZN(n2511) );
  NAND2_X1 U32100 ( .A1(n2516), .A2(n2515), .ZN(n2517) );
  NAND2_X1 U32110 ( .A1(n2517), .A2(IR_REG_31__SCAN_IN), .ZN(n2518) );
  XNOR2_X1 U32120 ( .A(n2518), .B(IR_REG_12__SCAN_IN), .ZN(n2821) );
  INV_X1 U32130 ( .A(DATAI_12_), .ZN(n4716) );
  MUX2_X1 U32140 ( .A(n2783), .B(n4716), .S(n3772), .Z(n3425) );
  NAND2_X1 U32150 ( .A1(n4513), .A2(n3425), .ZN(n2519) );
  NAND2_X1 U32160 ( .A1(n3365), .A2(n2519), .ZN(n2521) );
  NAND2_X1 U32170 ( .A1(n3921), .A2(n3371), .ZN(n2520) );
  NAND2_X1 U32180 ( .A1(n2521), .A2(n2520), .ZN(n3413) );
  NAND2_X1 U32190 ( .A1(n2672), .A2(REG0_REG_13__SCAN_IN), .ZN(n2530) );
  INV_X1 U32200 ( .A(n2522), .ZN(n2673) );
  NAND2_X1 U32210 ( .A1(n2673), .A2(REG1_REG_13__SCAN_IN), .ZN(n2529) );
  NAND2_X1 U32220 ( .A1(n3768), .A2(REG2_REG_13__SCAN_IN), .ZN(n2528) );
  INV_X1 U32230 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2523) );
  OAI21_X1 U32240 ( .B1(n2525), .B2(n2524), .A(n2523), .ZN(n2526) );
  NAND2_X1 U32250 ( .A1(n2526), .A2(n2535), .ZN(n3387) );
  OR2_X1 U32260 ( .A1(n2431), .A2(n3387), .ZN(n2527) );
  OR2_X1 U32270 ( .A1(n2531), .A2(n2732), .ZN(n2532) );
  XNOR2_X1 U32280 ( .A(n2532), .B(IR_REG_13__SCAN_IN), .ZN(n2824) );
  INV_X1 U32290 ( .A(DATAI_13_), .ZN(n2533) );
  MUX2_X1 U32300 ( .A(n4561), .B(n2533), .S(n3772), .Z(n3496) );
  NAND2_X1 U32310 ( .A1(n4268), .A2(n3496), .ZN(n2534) );
  NAND2_X1 U32320 ( .A1(n3413), .A2(n2534), .ZN(n3451) );
  NAND2_X1 U32330 ( .A1(n2672), .A2(REG0_REG_14__SCAN_IN), .ZN(n2540) );
  NAND2_X1 U32340 ( .A1(n2673), .A2(REG1_REG_14__SCAN_IN), .ZN(n2539) );
  NAND2_X1 U32350 ( .A1(n3768), .A2(REG2_REG_14__SCAN_IN), .ZN(n2538) );
  AND2_X1 U32360 ( .A1(n2535), .A2(n4884), .ZN(n2536) );
  OR2_X1 U32370 ( .A1(n2536), .A2(n2542), .ZN(n3457) );
  OR2_X1 U32380 ( .A1(n2431), .A2(n3457), .ZN(n2537) );
  NAND2_X1 U32390 ( .A1(n2571), .A2(IR_REG_31__SCAN_IN), .ZN(n2541) );
  XNOR2_X1 U32400 ( .A(n2541), .B(IR_REG_14__SCAN_IN), .ZN(n2826) );
  MUX2_X1 U32410 ( .A(n2826), .B(DATAI_14_), .S(n3772), .Z(n3464) );
  NAND2_X1 U32420 ( .A1(n4258), .A2(n3464), .ZN(n3868) );
  NAND2_X1 U32430 ( .A1(n3919), .A2(n4266), .ZN(n3747) );
  NAND2_X1 U32440 ( .A1(n3868), .A2(n3747), .ZN(n3786) );
  NAND2_X1 U32450 ( .A1(n2672), .A2(REG0_REG_15__SCAN_IN), .ZN(n2547) );
  NOR2_X1 U32460 ( .A1(n2542), .A2(REG3_REG_15__SCAN_IN), .ZN(n2543) );
  OR2_X1 U32470 ( .A1(n2551), .A2(n2543), .ZN(n3737) );
  OR2_X1 U32480 ( .A1(n2431), .A2(n3737), .ZN(n2546) );
  NAND2_X1 U32490 ( .A1(n3767), .A2(REG1_REG_15__SCAN_IN), .ZN(n2545) );
  NAND2_X1 U32500 ( .A1(n3768), .A2(REG2_REG_15__SCAN_IN), .ZN(n2544) );
  NAND4_X1 U32510 ( .A1(n2547), .A2(n2546), .A3(n2545), .A4(n2544), .ZN(n3918)
         );
  NAND2_X1 U32520 ( .A1(n2548), .A2(IR_REG_31__SCAN_IN), .ZN(n2558) );
  XNOR2_X1 U32530 ( .A(n2558), .B(IR_REG_15__SCAN_IN), .ZN(n2829) );
  MUX2_X1 U32540 ( .A(n2829), .B(DATAI_15_), .S(n3772), .Z(n3520) );
  NAND2_X1 U32550 ( .A1(n3918), .A2(n3520), .ZN(n2549) );
  INV_X1 U32560 ( .A(n4268), .ZN(n3920) );
  NAND2_X1 U32570 ( .A1(n3920), .A2(n3418), .ZN(n3452) );
  NOR2_X1 U32580 ( .A1(n3919), .A2(n3464), .ZN(n3467) );
  INV_X1 U32590 ( .A(n3918), .ZN(n4345) );
  INV_X1 U32600 ( .A(n3520), .ZN(n4257) );
  AOI22_X1 U32610 ( .A1(n3467), .A2(n2549), .B1(n4345), .B2(n4257), .ZN(n2550)
         );
  NAND2_X1 U32620 ( .A1(n3767), .A2(REG1_REG_16__SCAN_IN), .ZN(n2556) );
  NAND2_X1 U32630 ( .A1(n3768), .A2(REG2_REG_16__SCAN_IN), .ZN(n2555) );
  NAND2_X1 U32640 ( .A1(n2672), .A2(REG0_REG_16__SCAN_IN), .ZN(n2554) );
  OR2_X1 U32650 ( .A1(n2551), .A2(REG3_REG_16__SCAN_IN), .ZN(n2552) );
  NAND2_X1 U32660 ( .A1(n2564), .A2(n2552), .ZN(n4359) );
  OR2_X1 U32670 ( .A1(n2431), .A2(n4359), .ZN(n2553) );
  NAND2_X1 U32680 ( .A1(n2558), .A2(n2557), .ZN(n2559) );
  NAND2_X1 U32690 ( .A1(n2559), .A2(IR_REG_31__SCAN_IN), .ZN(n2560) );
  XNOR2_X1 U32700 ( .A(n2560), .B(IR_REG_16__SCAN_IN), .ZN(n2831) );
  MUX2_X1 U32710 ( .A(n2831), .B(DATAI_16_), .S(n3772), .Z(n3486) );
  NAND2_X1 U32720 ( .A1(n4244), .A2(n3486), .ZN(n3877) );
  INV_X1 U32730 ( .A(n3486), .ZN(n4346) );
  NAND2_X1 U32740 ( .A1(n3917), .A2(n4346), .ZN(n3874) );
  NAND2_X1 U32750 ( .A1(n3917), .A2(n3486), .ZN(n2562) );
  NAND2_X1 U32760 ( .A1(n3492), .A2(n2562), .ZN(n3507) );
  NAND2_X1 U32770 ( .A1(n3767), .A2(REG1_REG_17__SCAN_IN), .ZN(n2569) );
  NAND2_X1 U32780 ( .A1(n3768), .A2(REG2_REG_17__SCAN_IN), .ZN(n2568) );
  NAND2_X1 U32790 ( .A1(n2672), .A2(REG0_REG_17__SCAN_IN), .ZN(n2567) );
  INV_X1 U32800 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2563) );
  NAND2_X1 U32810 ( .A1(n2564), .A2(n2563), .ZN(n2565) );
  NAND2_X1 U32820 ( .A1(n2577), .A2(n2565), .ZN(n3510) );
  OR2_X1 U32830 ( .A1(n2431), .A2(n3510), .ZN(n2566) );
  INV_X1 U32840 ( .A(n2584), .ZN(n2572) );
  NAND2_X1 U32850 ( .A1(n2572), .A2(IR_REG_31__SCAN_IN), .ZN(n2573) );
  XNOR2_X1 U32860 ( .A(n2573), .B(IR_REG_17__SCAN_IN), .ZN(n2835) );
  MUX2_X1 U32870 ( .A(n2835), .B(DATAI_17_), .S(n3772), .Z(n3513) );
  NAND2_X1 U32880 ( .A1(n4178), .A2(n4243), .ZN(n2574) );
  NAND2_X1 U32890 ( .A1(n3507), .A2(n2574), .ZN(n2576) );
  INV_X1 U32900 ( .A(n4178), .ZN(n4349) );
  NAND2_X1 U32910 ( .A1(n4349), .A2(n3513), .ZN(n2575) );
  NAND2_X1 U32920 ( .A1(n2576), .A2(n2575), .ZN(n4163) );
  NAND2_X1 U32930 ( .A1(n2672), .A2(REG0_REG_18__SCAN_IN), .ZN(n2582) );
  NAND2_X1 U32940 ( .A1(n3767), .A2(REG1_REG_18__SCAN_IN), .ZN(n2581) );
  NAND2_X1 U32950 ( .A1(n3768), .A2(REG2_REG_18__SCAN_IN), .ZN(n2580) );
  INV_X1 U32960 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3716) );
  AND2_X1 U32970 ( .A1(n2577), .A2(n3716), .ZN(n2578) );
  OR2_X1 U32980 ( .A1(n2578), .A2(n2588), .ZN(n4166) );
  OR2_X1 U32990 ( .A1(n2431), .A2(n4166), .ZN(n2579) );
  NAND2_X1 U33000 ( .A1(n2584), .A2(n2583), .ZN(n2594) );
  NAND2_X1 U33010 ( .A1(n2594), .A2(IR_REG_31__SCAN_IN), .ZN(n2585) );
  XNOR2_X1 U33020 ( .A(n2585), .B(IR_REG_18__SCAN_IN), .ZN(n3942) );
  MUX2_X1 U33030 ( .A(n3942), .B(DATAI_18_), .S(n3772), .Z(n4174) );
  NAND2_X1 U33040 ( .A1(n4149), .A2(n4174), .ZN(n4141) );
  INV_X1 U33050 ( .A(n4149), .ZN(n3916) );
  NAND2_X1 U33060 ( .A1(n3916), .A2(n4170), .ZN(n4142) );
  NAND2_X1 U33070 ( .A1(n4149), .A2(n4170), .ZN(n2587) );
  NOR2_X1 U33080 ( .A1(n2588), .A2(REG3_REG_19__SCAN_IN), .ZN(n2589) );
  OR2_X1 U33090 ( .A1(n2600), .A2(n2589), .ZN(n3641) );
  OR2_X1 U33100 ( .A1(n3641), .A2(n2431), .ZN(n2593) );
  NAND2_X1 U33110 ( .A1(n3767), .A2(REG1_REG_19__SCAN_IN), .ZN(n2592) );
  NAND2_X1 U33120 ( .A1(n2672), .A2(REG0_REG_19__SCAN_IN), .ZN(n2591) );
  NAND2_X1 U33130 ( .A1(n3768), .A2(REG2_REG_19__SCAN_IN), .ZN(n2590) );
  NAND4_X1 U33140 ( .A1(n2593), .A2(n2592), .A3(n2591), .A4(n2590), .ZN(n4176)
         );
  NAND2_X1 U33150 ( .A1(n2679), .A2(IR_REG_31__SCAN_IN), .ZN(n2597) );
  NAND2_X1 U33160 ( .A1(n2597), .A2(n2677), .ZN(n2682) );
  OR2_X1 U33170 ( .A1(n2597), .A2(n2677), .ZN(n2598) );
  INV_X1 U33180 ( .A(DATAI_19_), .ZN(n2599) );
  MUX2_X1 U33190 ( .A(n3954), .B(n2599), .S(n3772), .Z(n3644) );
  NOR2_X1 U33200 ( .A1(n4176), .A2(n4154), .ZN(n3814) );
  NAND2_X1 U33210 ( .A1(n4176), .A2(n4154), .ZN(n3813) );
  OR2_X1 U33220 ( .A1(n2600), .A2(REG3_REG_20__SCAN_IN), .ZN(n2601) );
  NAND2_X1 U33230 ( .A1(n2608), .A2(n2601), .ZN(n4130) );
  NAND2_X1 U33240 ( .A1(n3768), .A2(REG2_REG_20__SCAN_IN), .ZN(n2602) );
  OAI21_X1 U33250 ( .B1(n4130), .B2(n2431), .A(n2602), .ZN(n2606) );
  NAND2_X1 U33260 ( .A1(n2672), .A2(REG0_REG_20__SCAN_IN), .ZN(n2604) );
  NAND2_X1 U33270 ( .A1(n3767), .A2(REG1_REG_20__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U33280 ( .A1(n2604), .A2(n2603), .ZN(n2605) );
  NAND2_X1 U33290 ( .A1(n4225), .A2(n4128), .ZN(n2607) );
  INV_X1 U33300 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4106) );
  INV_X1 U33310 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3653) );
  NAND2_X1 U33320 ( .A1(n2608), .A2(n3653), .ZN(n2609) );
  NAND2_X1 U33330 ( .A1(n2619), .A2(n2609), .ZN(n4105) );
  NAND2_X1 U33340 ( .A1(n2672), .A2(REG0_REG_21__SCAN_IN), .ZN(n2611) );
  NAND2_X1 U33350 ( .A1(n3767), .A2(REG1_REG_21__SCAN_IN), .ZN(n2610) );
  AND2_X1 U33360 ( .A1(n2611), .A2(n2610), .ZN(n2612) );
  INV_X1 U33370 ( .A(n4086), .ZN(n4117) );
  NAND2_X1 U33380 ( .A1(n4098), .A2(n2615), .ZN(n2618) );
  INV_X1 U33390 ( .A(n4224), .ZN(n4110) );
  INV_X1 U33400 ( .A(n2616), .ZN(n2617) );
  INV_X1 U33410 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3703) );
  NAND2_X1 U33420 ( .A1(n2619), .A2(n3703), .ZN(n2620) );
  NAND2_X1 U33430 ( .A1(n2626), .A2(n2620), .ZN(n4092) );
  AOI22_X1 U33440 ( .A1(n3767), .A2(REG1_REG_22__SCAN_IN), .B1(n2672), .B2(
        REG0_REG_22__SCAN_IN), .ZN(n2622) );
  NAND2_X1 U33450 ( .A1(n3768), .A2(REG2_REG_22__SCAN_IN), .ZN(n2621) );
  NAND2_X1 U33460 ( .A1(n3772), .A2(DATAI_22_), .ZN(n4091) );
  NAND2_X1 U33470 ( .A1(n4067), .A2(n4091), .ZN(n2709) );
  INV_X1 U33480 ( .A(n2709), .ZN(n2623) );
  NOR2_X1 U33490 ( .A1(n4067), .A2(n4091), .ZN(n2708) );
  NOR2_X1 U33500 ( .A1(n2623), .A2(n2708), .ZN(n4081) );
  INV_X1 U33510 ( .A(n4091), .ZN(n4085) );
  INV_X1 U33520 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3634) );
  AND2_X1 U3353 ( .A1(n2626), .A2(n3634), .ZN(n2627) );
  OR2_X1 U33540 ( .A1(n2627), .A2(n2632), .ZN(n3639) );
  NAND2_X1 U3355 ( .A1(n3768), .A2(REG2_REG_23__SCAN_IN), .ZN(n2630) );
  NAND2_X1 U3356 ( .A1(n2672), .A2(REG0_REG_23__SCAN_IN), .ZN(n2629) );
  NAND2_X1 U3357 ( .A1(n3767), .A2(REG1_REG_23__SCAN_IN), .ZN(n2628) );
  NAND3_X1 U3358 ( .A1(n2630), .A2(n2629), .A3(n2628), .ZN(n2631) );
  NAND2_X1 U3359 ( .A1(n3772), .A2(DATAI_23_), .ZN(n3632) );
  NAND2_X1 U3360 ( .A1(n4047), .A2(n4071), .ZN(n3791) );
  NOR2_X1 U3361 ( .A1(n4047), .A2(n4071), .ZN(n3793) );
  NOR2_X1 U3362 ( .A1(n2632), .A2(REG3_REG_24__SCAN_IN), .ZN(n2633) );
  OR2_X1 U3363 ( .A1(n2647), .A2(n2633), .ZN(n4054) );
  NAND2_X1 U3364 ( .A1(n3768), .A2(REG2_REG_24__SCAN_IN), .ZN(n2636) );
  NAND2_X1 U3365 ( .A1(n2672), .A2(REG0_REG_24__SCAN_IN), .ZN(n2635) );
  NAND2_X1 U3366 ( .A1(n2673), .A2(REG1_REG_24__SCAN_IN), .ZN(n2634) );
  OAI21_X1 U3367 ( .B1(n4054), .B2(n2431), .A(n2637), .ZN(n4029) );
  INV_X1 U3368 ( .A(n4029), .ZN(n4070) );
  NAND2_X1 U3369 ( .A1(n3772), .A2(DATAI_24_), .ZN(n3579) );
  NOR2_X1 U3370 ( .A1(n4070), .A2(n3579), .ZN(n2638) );
  INV_X1 U3371 ( .A(REG3_REG_25__SCAN_IN), .ZN(n2639) );
  XNOR2_X1 U3372 ( .A(n2647), .B(n2639), .ZN(n4035) );
  NAND2_X1 U3373 ( .A1(n4035), .A2(n2666), .ZN(n2644) );
  NAND2_X1 U3374 ( .A1(n3768), .A2(REG2_REG_25__SCAN_IN), .ZN(n2642) );
  NAND2_X1 U3375 ( .A1(n3767), .A2(REG1_REG_25__SCAN_IN), .ZN(n2641) );
  NAND2_X1 U3376 ( .A1(n2672), .A2(REG0_REG_25__SCAN_IN), .ZN(n2640) );
  INV_X1 U3377 ( .A(n3915), .ZN(n4050) );
  NAND2_X1 U3378 ( .A1(n3772), .A2(DATAI_25_), .ZN(n3587) );
  INV_X1 U3379 ( .A(n2645), .ZN(n4003) );
  AND2_X1 U3380 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2646) );
  AOI21_X1 U3381 ( .B1(n2647), .B2(REG3_REG_25__SCAN_IN), .A(
        REG3_REG_26__SCAN_IN), .ZN(n2648) );
  NAND2_X1 U3382 ( .A1(n3768), .A2(REG2_REG_26__SCAN_IN), .ZN(n2651) );
  NAND2_X1 U3383 ( .A1(n2672), .A2(REG0_REG_26__SCAN_IN), .ZN(n2650) );
  NAND2_X1 U3384 ( .A1(n2673), .A2(REG1_REG_26__SCAN_IN), .ZN(n2649) );
  OAI21_X1 U3385 ( .B1(n4017), .B2(n2431), .A(n2652), .ZN(n3993) );
  INV_X1 U3386 ( .A(n3993), .ZN(n4198) );
  NAND2_X1 U3387 ( .A1(n3772), .A2(DATAI_26_), .ZN(n4014) );
  NAND2_X1 U3388 ( .A1(n4003), .A2(n2367), .ZN(n2654) );
  INV_X1 U3389 ( .A(n4014), .ZN(n4010) );
  NAND2_X1 U3390 ( .A1(n2655), .A2(REG3_REG_27__SCAN_IN), .ZN(n2664) );
  OR2_X1 U3391 ( .A1(n2655), .A2(REG3_REG_27__SCAN_IN), .ZN(n2656) );
  NAND2_X1 U3392 ( .A1(n3991), .A2(n2666), .ZN(n2661) );
  NAND2_X1 U3393 ( .A1(n3768), .A2(REG2_REG_27__SCAN_IN), .ZN(n2659) );
  NAND2_X1 U3394 ( .A1(n2673), .A2(REG1_REG_27__SCAN_IN), .ZN(n2658) );
  NAND2_X1 U3395 ( .A1(n2672), .A2(REG0_REG_27__SCAN_IN), .ZN(n2657) );
  AND3_X1 U3396 ( .A1(n2659), .A2(n2658), .A3(n2657), .ZN(n2660) );
  NAND2_X1 U3397 ( .A1(n3772), .A2(DATAI_27_), .ZN(n4197) );
  INV_X1 U3398 ( .A(n4197), .ZN(n4000) );
  INV_X1 U3399 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3612) );
  NAND2_X1 U3400 ( .A1(n2664), .A2(n3612), .ZN(n2665) );
  NAND2_X1 U3401 ( .A1(n3978), .A2(n2666), .ZN(n2671) );
  NAND2_X1 U3402 ( .A1(n3768), .A2(REG2_REG_28__SCAN_IN), .ZN(n2669) );
  NAND2_X1 U3403 ( .A1(n2672), .A2(REG0_REG_28__SCAN_IN), .ZN(n2668) );
  NAND2_X1 U3404 ( .A1(n3767), .A2(REG1_REG_28__SCAN_IN), .ZN(n2667) );
  AND3_X1 U3405 ( .A1(n2669), .A2(n2668), .A3(n2667), .ZN(n2670) );
  NAND2_X1 U3406 ( .A1(n3772), .A2(DATAI_28_), .ZN(n3613) );
  NAND2_X1 U3407 ( .A1(n3987), .A2(n3613), .ZN(n3764) );
  INV_X1 U3408 ( .A(n3613), .ZN(n2851) );
  NAND2_X1 U3409 ( .A1(n3966), .A2(n2851), .ZN(n3763) );
  NAND2_X1 U3410 ( .A1(n3772), .A2(DATAI_29_), .ZN(n3774) );
  AOI22_X1 U3411 ( .A1(n2673), .A2(REG1_REG_29__SCAN_IN), .B1(n2672), .B2(
        REG0_REG_29__SCAN_IN), .ZN(n2675) );
  NAND2_X1 U3412 ( .A1(n3768), .A2(REG2_REG_29__SCAN_IN), .ZN(n2674) );
  OAI211_X1 U3413 ( .C1(n3970), .C2(n2431), .A(n2675), .B(n2674), .ZN(n3914)
         );
  XOR2_X1 U3414 ( .A(n3774), .B(n3914), .Z(n3809) );
  XNOR2_X1 U3415 ( .A(n2676), .B(n3809), .ZN(n3964) );
  INV_X1 U3416 ( .A(IR_REG_20__SCAN_IN), .ZN(n2683) );
  NAND2_X1 U3417 ( .A1(n2683), .A2(n2677), .ZN(n2678) );
  INV_X1 U3418 ( .A(IR_REG_21__SCAN_IN), .ZN(n2680) );
  NAND2_X1 U3419 ( .A1(n2730), .A2(n2680), .ZN(n2685) );
  NAND2_X1 U3420 ( .A1(n2685), .A2(IR_REG_31__SCAN_IN), .ZN(n2686) );
  INV_X1 U3421 ( .A(IR_REG_22__SCAN_IN), .ZN(n4785) );
  INV_X1 U3422 ( .A(n2871), .ZN(n4337) );
  XNOR2_X1 U3423 ( .A(n3152), .B(n4337), .ZN(n2687) );
  NAND2_X1 U3424 ( .A1(n2687), .A2(n3954), .ZN(n4516) );
  AND2_X1 U3425 ( .A1(n3903), .A2(n4181), .ZN(n3156) );
  INV_X1 U3426 ( .A(n4601), .ZN(n4607) );
  NAND2_X1 U3427 ( .A1(n3964), .A2(n4590), .ZN(n2723) );
  INV_X1 U3428 ( .A(n4533), .ZN(n3064) );
  NAND2_X1 U3429 ( .A1(n4539), .A2(n2689), .ZN(n2691) );
  NAND2_X1 U3430 ( .A1(n2691), .A2(n3162), .ZN(n3170) );
  NAND2_X1 U3431 ( .A1(n3170), .A2(n2692), .ZN(n2693) );
  XNOR2_X1 U3432 ( .A(n2874), .B(n3832), .ZN(n3105) );
  NAND2_X1 U3433 ( .A1(n2693), .A2(n3105), .ZN(n3107) );
  NAND2_X1 U3434 ( .A1(n3833), .A2(n3832), .ZN(n3834) );
  INV_X1 U3435 ( .A(n3835), .ZN(n2694) );
  AND2_X1 U3436 ( .A1(n3926), .A2(n3098), .ZN(n3134) );
  NAND2_X1 U3437 ( .A1(n3256), .A2(n3269), .ZN(n3847) );
  NAND2_X1 U3438 ( .A1(n3925), .A2(n3257), .ZN(n3848) );
  NAND2_X1 U3439 ( .A1(n3212), .A2(n3848), .ZN(n2695) );
  INV_X1 U3440 ( .A(n3925), .ZN(n3241) );
  NAND2_X1 U3441 ( .A1(n3241), .A2(n3214), .ZN(n3840) );
  INV_X1 U3442 ( .A(n3841), .ZN(n2696) );
  NAND2_X1 U3443 ( .A1(n3339), .A2(n3296), .ZN(n3844) );
  NAND2_X1 U3444 ( .A1(n3924), .A2(n3302), .ZN(n3849) );
  AND2_X1 U3445 ( .A1(n3923), .A2(n3338), .ZN(n3277) );
  NAND2_X1 U3446 ( .A1(n3324), .A2(n3282), .ZN(n3845) );
  NAND2_X1 U3447 ( .A1(n4511), .A2(n3329), .ZN(n3860) );
  NAND2_X1 U3448 ( .A1(n3321), .A2(n3860), .ZN(n2697) );
  NAND2_X1 U3449 ( .A1(n3279), .A2(n3322), .ZN(n3855) );
  NAND2_X1 U3450 ( .A1(n2697), .A2(n3855), .ZN(n4509) );
  NOR2_X1 U3451 ( .A1(n3921), .A2(n3425), .ZN(n3864) );
  NAND2_X1 U3452 ( .A1(n3921), .A2(n3425), .ZN(n3408) );
  NAND2_X1 U3453 ( .A1(n3920), .A2(n3496), .ZN(n3410) );
  NAND2_X1 U3454 ( .A1(n4268), .A2(n3418), .ZN(n3867) );
  NAND2_X2 U3455 ( .A1(n2698), .A2(n3867), .ZN(n3750) );
  NAND2_X1 U3456 ( .A1(n4345), .A2(n3520), .ZN(n3866) );
  NAND2_X1 U3457 ( .A1(n3918), .A2(n4257), .ZN(n3748) );
  NAND2_X1 U34580 ( .A1(n3866), .A2(n3748), .ZN(n3782) );
  INV_X1 U34590 ( .A(n3868), .ZN(n2699) );
  NOR2_X1 U3460 ( .A1(n3782), .A2(n2699), .ZN(n2700) );
  INV_X1 U3461 ( .A(n3874), .ZN(n3752) );
  OR2_X1 U3462 ( .A1(n4178), .A2(n3513), .ZN(n4137) );
  NAND2_X1 U3463 ( .A1(n4176), .A2(n3644), .ZN(n2701) );
  AND2_X1 U3464 ( .A1(n4142), .A2(n2701), .ZN(n2703) );
  AND2_X1 U3465 ( .A1(n4137), .A2(n2703), .ZN(n3751) );
  NAND2_X1 U3466 ( .A1(n4138), .A2(n3751), .ZN(n4120) );
  NAND2_X1 U34670 ( .A1(n4178), .A2(n3513), .ZN(n4139) );
  NAND2_X1 U3468 ( .A1(n4141), .A2(n4139), .ZN(n2704) );
  NOR2_X1 U34690 ( .A1(n4176), .A2(n3644), .ZN(n2702) );
  AOI21_X1 U3470 ( .B1(n2704), .B2(n2703), .A(n2702), .ZN(n4119) );
  NAND2_X1 U34710 ( .A1(n4225), .A2(n3787), .ZN(n2705) );
  NAND2_X1 U3472 ( .A1(n4119), .A2(n2705), .ZN(n3881) );
  INV_X1 U34730 ( .A(n3881), .ZN(n2707) );
  NAND2_X1 U3474 ( .A1(n4146), .A2(n4128), .ZN(n3880) );
  INV_X1 U34750 ( .A(n3880), .ZN(n2706) );
  NOR2_X1 U3476 ( .A1(n4086), .A2(n4224), .ZN(n4062) );
  NOR2_X1 U34770 ( .A1(n2708), .A2(n4062), .ZN(n3885) );
  INV_X1 U3478 ( .A(n3885), .ZN(n2710) );
  NAND2_X1 U34790 ( .A1(n4086), .A2(n4224), .ZN(n3879) );
  INV_X1 U3480 ( .A(n3879), .ZN(n3780) );
  INV_X1 U34810 ( .A(n2708), .ZN(n4063) );
  OAI21_X1 U3482 ( .B1(n4089), .B2(n4071), .A(n2709), .ZN(n3883) );
  AOI21_X1 U34830 ( .B1(n3780), .B2(n4063), .A(n3883), .ZN(n3758) );
  OAI21_X1 U3484 ( .B1(n4061), .B2(n2710), .A(n3758), .ZN(n4043) );
  NOR2_X1 U34850 ( .A1(n4047), .A2(n3632), .ZN(n4041) );
  NOR2_X1 U3486 ( .A1(n4029), .A2(n3579), .ZN(n3802) );
  NOR2_X1 U34870 ( .A1(n4041), .A2(n3802), .ZN(n3756) );
  NAND2_X1 U3488 ( .A1(n4043), .A2(n3756), .ZN(n4025) );
  NAND2_X1 U34890 ( .A1(n3915), .A2(n3587), .ZN(n3800) );
  NAND2_X1 U3490 ( .A1(n4029), .A2(n3579), .ZN(n4024) );
  AND2_X1 U34910 ( .A1(n3800), .A2(n4024), .ZN(n3886) );
  NAND2_X1 U3492 ( .A1(n4025), .A2(n3886), .ZN(n4006) );
  NOR2_X1 U34930 ( .A1(n3993), .A2(n4014), .ZN(n3798) );
  NOR2_X1 U3494 ( .A1(n3915), .A2(n3587), .ZN(n4004) );
  NOR2_X1 U34950 ( .A1(n3798), .A2(n4004), .ZN(n3889) );
  NAND2_X1 U3496 ( .A1(n3993), .A2(n4014), .ZN(n3893) );
  INV_X1 U34970 ( .A(n3893), .ZN(n3799) );
  AOI21_X2 U3498 ( .B1(n4006), .B2(n3889), .A(n3799), .ZN(n3986) );
  NAND2_X1 U34990 ( .A1(n4011), .A2(n4197), .ZN(n3892) );
  NAND2_X1 U3500 ( .A1(n3729), .A2(n4000), .ZN(n3762) );
  NAND2_X1 U35010 ( .A1(n4337), .A2(n4181), .ZN(n2713) );
  INV_X1 U3502 ( .A(n3903), .ZN(n4338) );
  NAND2_X1 U35030 ( .A1(n4338), .A2(n2711), .ZN(n2712) );
  XNOR2_X1 U3504 ( .A(n2715), .B(n2714), .ZN(n4364) );
  NAND2_X1 U35050 ( .A1(n4337), .A2(n2711), .ZN(n2915) );
  INV_X1 U35060 ( .A(n2915), .ZN(n2795) );
  OR2_X1 U35070 ( .A1(n2716), .A2(n2732), .ZN(n2717) );
  XNOR2_X1 U35080 ( .A(n2717), .B(n4906), .ZN(n4343) );
  NAND2_X1 U35090 ( .A1(n2795), .A2(n4343), .ZN(n4535) );
  AOI21_X1 U35100 ( .B1(B_REG_SCAN_IN), .B2(n4364), .A(n4535), .ZN(n3959) );
  NAND2_X1 U35110 ( .A1(n3767), .A2(REG1_REG_30__SCAN_IN), .ZN(n2720) );
  NAND2_X1 U35120 ( .A1(n3768), .A2(REG2_REG_30__SCAN_IN), .ZN(n2719) );
  NAND2_X1 U35130 ( .A1(n2672), .A2(REG0_REG_30__SCAN_IN), .ZN(n2718) );
  NAND3_X1 U35140 ( .A1(n2720), .A2(n2719), .A3(n2718), .ZN(n3913) );
  AOI22_X1 U35150 ( .A1(n2366), .A2(n4519), .B1(n3959), .B2(n3913), .ZN(n3969)
         );
  NOR2_X2 U35160 ( .A1(n2915), .A2(n4343), .ZN(n4532) );
  INV_X1 U35170 ( .A(n3774), .ZN(n3968) );
  AOI22_X1 U35180 ( .A1(n3987), .A2(n4532), .B1(n3968), .B2(n4530), .ZN(n2722)
         );
  NOR2_X1 U35190 ( .A1(n2724), .A2(n2732), .ZN(n2725) );
  MUX2_X1 U35200 ( .A(n2732), .B(n2725), .S(IR_REG_25__SCAN_IN), .Z(n2726) );
  INV_X1 U35210 ( .A(n2726), .ZN(n2728) );
  NAND2_X1 U35220 ( .A1(n2728), .A2(n2727), .ZN(n3008) );
  NAND2_X1 U35230 ( .A1(n3008), .A2(B_REG_SCAN_IN), .ZN(n2736) );
  AND2_X1 U35240 ( .A1(n4785), .A2(n2680), .ZN(n2729) );
  NAND2_X1 U35250 ( .A1(n2730), .A2(n2729), .ZN(n2731) );
  OR2_X1 U35260 ( .A1(n2732), .A2(n4971), .ZN(n2733) );
  NAND2_X1 U35270 ( .A1(n2741), .A2(n2733), .ZN(n2735) );
  MUX2_X1 U35280 ( .A(n2736), .B(B_REG_SCAN_IN), .S(n2740), .Z(n2738) );
  NAND2_X1 U35290 ( .A1(n2727), .A2(IR_REG_31__SCAN_IN), .ZN(n2737) );
  NAND2_X1 U35300 ( .A1(n2738), .A2(n4336), .ZN(n3014) );
  OR2_X1 U35310 ( .A1(n3014), .A2(D_REG_1__SCAN_IN), .ZN(n2911) );
  NAND2_X1 U35320 ( .A1(n3008), .A2(n2756), .ZN(n3017) );
  NAND2_X1 U35330 ( .A1(n2911), .A2(n3017), .ZN(n2755) );
  XNOR2_X1 U35340 ( .A(n2741), .B(n4971), .ZN(n2928) );
  NAND2_X1 U35350 ( .A1(n2869), .A2(n4554), .ZN(n3146) );
  NAND2_X1 U35360 ( .A1(n4601), .A2(n2721), .ZN(n2936) );
  AND2_X1 U35370 ( .A1(n3903), .A2(n3954), .ZN(n2913) );
  OR2_X1 U35380 ( .A1(n2915), .A2(n2913), .ZN(n3148) );
  NAND2_X1 U35390 ( .A1(n2936), .A2(n3148), .ZN(n2742) );
  NOR2_X1 U35400 ( .A1(n3146), .A2(n2742), .ZN(n2754) );
  NOR2_X1 U35410 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_26__SCAN_IN), .ZN(n2746)
         );
  NOR4_X1 U35420 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2745) );
  NOR4_X1 U35430 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2744) );
  NOR4_X1 U35440 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2743) );
  NAND4_X1 U35450 ( .A1(n2746), .A2(n2745), .A3(n2744), .A4(n2743), .ZN(n2752)
         );
  NOR4_X1 U35460 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2750) );
  NOR4_X1 U35470 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_29__SCAN_IN), .ZN(n2749) );
  NOR4_X1 U35480 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2748) );
  NOR4_X1 U35490 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2747) );
  NAND4_X1 U35500 ( .A1(n2750), .A2(n2749), .A3(n2748), .A4(n2747), .ZN(n2751)
         );
  NOR2_X1 U35510 ( .A1(n2752), .A2(n2751), .ZN(n2753) );
  OR2_X1 U35520 ( .A1(n3014), .A2(n2753), .ZN(n2910) );
  OR2_X1 U35530 ( .A1(n3014), .A2(D_REG_0__SCAN_IN), .ZN(n2758) );
  NAND2_X1 U35540 ( .A1(n2757), .A2(n2756), .ZN(n3015) );
  AND2_X2 U35550 ( .A1(n2855), .A2(n3150), .ZN(n4613) );
  NAND2_X1 U35560 ( .A1(n2866), .A2(n4613), .ZN(n2762) );
  NAND2_X1 U35570 ( .A1(n3205), .A2(n3204), .ZN(n3138) );
  NAND2_X1 U35580 ( .A1(n3217), .A2(n3257), .ZN(n3216) );
  AND2_X2 U35590 ( .A1(n4016), .A2(n4197), .ZN(n3996) );
  NAND2_X1 U35600 ( .A1(n2857), .A2(n3968), .ZN(n2759) );
  NAND2_X2 U35610 ( .A1(n4190), .A2(n2759), .ZN(n3971) );
  NAND2_X1 U35620 ( .A1(n2762), .A2(n2761), .ZN(U3515) );
  INV_X2 U35630 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U35640 ( .A(n3942), .ZN(n4556) );
  INV_X1 U35650 ( .A(REG2_REG_18__SCAN_IN), .ZN(n2763) );
  AOI22_X1 U35660 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4556), .B1(n3942), .B2(
        n2763), .ZN(n2797) );
  INV_X1 U35670 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4455) );
  NOR2_X1 U35680 ( .A1(n4455), .A2(n4561), .ZN(n4454) );
  INV_X1 U35690 ( .A(n2799), .ZN(n4563) );
  INV_X1 U35700 ( .A(REG2_REG_11__SCAN_IN), .ZN(n2764) );
  AOI22_X1 U35710 ( .A1(REG2_REG_11__SCAN_IN), .A2(n2799), .B1(n4563), .B2(
        n2764), .ZN(n4439) );
  INV_X1 U35720 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3284) );
  INV_X1 U35730 ( .A(n2817), .ZN(n4564) );
  AOI22_X1 U35740 ( .A1(n2817), .A2(REG2_REG_9__SCAN_IN), .B1(n3284), .B2(
        n4564), .ZN(n4418) );
  INV_X1 U35750 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3249) );
  INV_X1 U35760 ( .A(n2813), .ZN(n4565) );
  AOI22_X1 U35770 ( .A1(n2813), .A2(REG2_REG_7__SCAN_IN), .B1(n3249), .B2(
        n4565), .ZN(n4400) );
  NAND2_X1 U35780 ( .A1(n2809), .A2(REG2_REG_5__SCAN_IN), .ZN(n2771) );
  INV_X1 U35790 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3267) );
  INV_X1 U35800 ( .A(n2809), .ZN(n4567) );
  AOI22_X1 U35810 ( .A1(n2809), .A2(REG2_REG_5__SCAN_IN), .B1(n3267), .B2(
        n4567), .ZN(n4377) );
  NAND2_X1 U3582 ( .A1(n3005), .A2(REG2_REG_1__SCAN_IN), .ZN(n2765) );
  NAND3_X1 U3583 ( .A1(n3935), .A2(REG2_REG_0__SCAN_IN), .A3(IR_REG_0__SCAN_IN), .ZN(n3934) );
  NAND2_X1 U3584 ( .A1(n3929), .A2(REG2_REG_1__SCAN_IN), .ZN(n3051) );
  AOI21_X1 U3585 ( .B1(n2221), .B2(REG2_REG_2__SCAN_IN), .A(n3050), .ZN(n2767)
         );
  XNOR2_X1 U3586 ( .A(n2767), .B(n4340), .ZN(n3019) );
  INV_X1 U3587 ( .A(n2767), .ZN(n2768) );
  INV_X1 U3588 ( .A(n4339), .ZN(n3042) );
  XNOR2_X1 U3589 ( .A(n2770), .B(n4339), .ZN(n3036) );
  NAND2_X1 U3590 ( .A1(n3036), .A2(REG2_REG_4__SCAN_IN), .ZN(n2769) );
  OAI21_X1 U3591 ( .B1(n2770), .B2(n3042), .A(n2769), .ZN(n4376) );
  NAND2_X1 U3592 ( .A1(n4377), .A2(n4376), .ZN(n4375) );
  NAND2_X1 U3593 ( .A1(n2810), .A2(n2773), .ZN(n2774) );
  NAND2_X1 U3594 ( .A1(n4400), .A2(n4399), .ZN(n4398) );
  NAND2_X1 U3595 ( .A1(n2813), .A2(REG2_REG_7__SCAN_IN), .ZN(n2775) );
  NAND2_X1 U3596 ( .A1(n4403), .A2(n2776), .ZN(n2777) );
  NAND2_X1 U3597 ( .A1(n2817), .A2(REG2_REG_9__SCAN_IN), .ZN(n2778) );
  NAND2_X1 U3598 ( .A1(n4424), .A2(n2780), .ZN(n2781) );
  NAND2_X1 U3599 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4428), .ZN(n4427) );
  NAND2_X1 U3600 ( .A1(n2781), .A2(n4427), .ZN(n4438) );
  NAND2_X1 U3601 ( .A1(n4439), .A2(n4438), .ZN(n4437) );
  NAND2_X1 U3602 ( .A1(REG2_REG_11__SCAN_IN), .A2(n2799), .ZN(n2782) );
  NAND2_X1 U3603 ( .A1(n2821), .A2(n2784), .ZN(n2785) );
  OAI22_X1 U3604 ( .A1(n4454), .A2(n4458), .B1(REG2_REG_13__SCAN_IN), .B2(
        n2824), .ZN(n2786) );
  INV_X1 U3605 ( .A(n2826), .ZN(n4560) );
  XNOR2_X1 U3606 ( .A(n2786), .B(n4560), .ZN(n4469) );
  INV_X1 U3607 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4470) );
  NOR2_X1 U3608 ( .A1(n4469), .A2(n4470), .ZN(n4468) );
  NOR2_X1 U3609 ( .A1(n4560), .A2(n2786), .ZN(n2787) );
  NAND2_X1 U3610 ( .A1(REG2_REG_15__SCAN_IN), .A2(n2829), .ZN(n2788) );
  OAI21_X1 U3611 ( .B1(REG2_REG_15__SCAN_IN), .B2(n2829), .A(n2788), .ZN(n4477) );
  INV_X1 U3612 ( .A(n2831), .ZN(n4558) );
  NAND2_X1 U3613 ( .A1(n2790), .A2(n4558), .ZN(n2791) );
  INV_X1 U3614 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4486) );
  NAND2_X1 U3615 ( .A1(n4488), .A2(n4486), .ZN(n4487) );
  NOR2_X1 U3616 ( .A1(n2835), .A2(REG2_REG_17__SCAN_IN), .ZN(n2792) );
  AOI21_X1 U3617 ( .B1(REG2_REG_17__SCAN_IN), .B2(n2835), .A(n2792), .ZN(n4498) );
  INV_X1 U3618 ( .A(n2792), .ZN(n2793) );
  OR2_X1 U3619 ( .A1(n2928), .A2(U3149), .ZN(n3911) );
  NAND2_X1 U3620 ( .A1(n3146), .A2(n3911), .ZN(n2841) );
  AOI21_X1 U3621 ( .B1(n2795), .B2(n2928), .A(n2794), .ZN(n2839) );
  INV_X1 U3622 ( .A(n4364), .ZN(n3030) );
  NOR2_X1 U3623 ( .A1(n4343), .A2(n3030), .ZN(n3907) );
  INV_X1 U3624 ( .A(n4456), .ZN(n4495) );
  AOI211_X1 U3625 ( .C1(n2797), .C2(n2796), .A(n3944), .B(n4495), .ZN(n2848)
         );
  INV_X1 U3626 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U3627 ( .A1(REG1_REG_18__SCAN_IN), .A2(n3942), .B1(n4556), .B2(
        n3948), .ZN(n2838) );
  INV_X1 U3628 ( .A(REG1_REG_13__SCAN_IN), .ZN(n2798) );
  AOI22_X1 U3629 ( .A1(REG1_REG_13__SCAN_IN), .A2(n2824), .B1(n4561), .B2(
        n2798), .ZN(n4464) );
  INV_X1 U3630 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4632) );
  AOI22_X1 U3631 ( .A1(REG1_REG_11__SCAN_IN), .A2(n2799), .B1(n4563), .B2(
        n4632), .ZN(n4436) );
  INV_X1 U3632 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2800) );
  AOI22_X1 U3633 ( .A1(n2817), .A2(REG1_REG_9__SCAN_IN), .B1(n2800), .B2(n4564), .ZN(n4415) );
  XNOR2_X1 U3634 ( .A(n3005), .B(REG1_REG_1__SCAN_IN), .ZN(n3933) );
  AND2_X1 U3635 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3932)
         );
  NAND2_X1 U3636 ( .A1(n3933), .A2(n3932), .ZN(n3931) );
  NAND2_X1 U3637 ( .A1(n3929), .A2(REG1_REG_1__SCAN_IN), .ZN(n2801) );
  NAND2_X1 U3638 ( .A1(n3931), .A2(n2801), .ZN(n3048) );
  INV_X1 U3639 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2802) );
  MUX2_X1 U3640 ( .A(REG1_REG_2__SCAN_IN), .B(n2802), .S(n4341), .Z(n3049) );
  NAND2_X1 U3641 ( .A1(n3048), .A2(n3049), .ZN(n3047) );
  NAND2_X1 U3642 ( .A1(n2221), .A2(REG1_REG_2__SCAN_IN), .ZN(n2803) );
  NAND2_X1 U3643 ( .A1(n3047), .A2(n2803), .ZN(n2804) );
  INV_X1 U3644 ( .A(n4340), .ZN(n3020) );
  XNOR2_X1 U3645 ( .A(n2804), .B(n3020), .ZN(n3023) );
  NAND2_X1 U3646 ( .A1(n3023), .A2(REG1_REG_3__SCAN_IN), .ZN(n3022) );
  NAND2_X1 U3647 ( .A1(n2804), .A2(n4340), .ZN(n2805) );
  NAND2_X1 U3648 ( .A1(n3022), .A2(n2805), .ZN(n2806) );
  XNOR2_X1 U3649 ( .A(n2806), .B(n3042), .ZN(n3038) );
  NAND2_X1 U3650 ( .A1(n3038), .A2(REG1_REG_4__SCAN_IN), .ZN(n3037) );
  NAND2_X1 U3651 ( .A1(n2809), .A2(REG1_REG_5__SCAN_IN), .ZN(n2808) );
  OAI21_X1 U3652 ( .B1(n2809), .B2(REG1_REG_5__SCAN_IN), .A(n2808), .ZN(n4371)
         );
  AOI21_X1 U3653 ( .B1(REG1_REG_5__SCAN_IN), .B2(n2809), .A(n4370), .ZN(n2811)
         );
  XNOR2_X1 U3654 ( .A(n2811), .B(n2772), .ZN(n4382) );
  INV_X1 U3655 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4383) );
  NOR2_X1 U3656 ( .A1(n2811), .A2(n2772), .ZN(n2812) );
  NAND2_X1 U3657 ( .A1(n2813), .A2(REG1_REG_7__SCAN_IN), .ZN(n4391) );
  NOR2_X1 U3658 ( .A1(n2813), .A2(REG1_REG_7__SCAN_IN), .ZN(n4390) );
  NAND2_X1 U3659 ( .A1(n4403), .A2(n2815), .ZN(n2816) );
  NAND2_X1 U3660 ( .A1(n2816), .A2(n4404), .ZN(n4414) );
  NAND2_X1 U3661 ( .A1(n4415), .A2(n4414), .ZN(n4413) );
  NAND2_X1 U3662 ( .A1(n2817), .A2(REG1_REG_9__SCAN_IN), .ZN(n2818) );
  NAND2_X1 U3663 ( .A1(n4424), .A2(n2819), .ZN(n2820) );
  NAND2_X1 U3664 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4426), .ZN(n4425) );
  NAND2_X1 U3665 ( .A1(n2820), .A2(n4425), .ZN(n4435) );
  NAND2_X1 U3666 ( .A1(n4436), .A2(n4435), .ZN(n4434) );
  NAND2_X1 U3667 ( .A1(n2821), .A2(n2822), .ZN(n2823) );
  NAND2_X1 U3668 ( .A1(n2823), .A2(n4450), .ZN(n4463) );
  NAND2_X1 U3669 ( .A1(n4464), .A2(n4463), .ZN(n4462) );
  NAND2_X1 U3670 ( .A1(REG1_REG_13__SCAN_IN), .A2(n2824), .ZN(n2825) );
  NAND2_X1 U3671 ( .A1(n2826), .A2(n2827), .ZN(n2828) );
  NAND2_X1 U3672 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4474), .ZN(n4473) );
  NAND2_X1 U3673 ( .A1(n2828), .A2(n4473), .ZN(n4482) );
  INV_X1 U3674 ( .A(n2829), .ZN(n4559) );
  AOI22_X1 U3675 ( .A1(REG1_REG_15__SCAN_IN), .A2(n2829), .B1(n4559), .B2(
        n4262), .ZN(n4483) );
  NAND2_X1 U3676 ( .A1(REG1_REG_15__SCAN_IN), .A2(n2829), .ZN(n2830) );
  NOR2_X1 U3677 ( .A1(n2831), .A2(n2832), .ZN(n2833) );
  XNOR2_X1 U3678 ( .A(n2832), .B(n2831), .ZN(n4491) );
  NOR2_X1 U3679 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4491), .ZN(n4492) );
  INV_X1 U3680 ( .A(REG1_REG_17__SCAN_IN), .ZN(n2834) );
  INV_X1 U3681 ( .A(n2835), .ZN(n4557) );
  AOI22_X1 U3682 ( .A1(n2835), .A2(n2834), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4557), .ZN(n4503) );
  NOR2_X1 U3683 ( .A1(n2835), .A2(REG1_REG_17__SCAN_IN), .ZN(n2836) );
  NOR2_X1 U3684 ( .A1(n4505), .A2(n2836), .ZN(n2837) );
  OAI211_X1 U3685 ( .C1(n2838), .C2(n2837), .A(n4502), .B(n3947), .ZN(n2846)
         );
  NAND2_X1 U3686 ( .A1(n4366), .A2(n4343), .ZN(n4508) );
  INV_X1 U3687 ( .A(n2839), .ZN(n2840) );
  NOR2_X1 U3688 ( .A1(STATE_REG_SCAN_IN), .A2(n3716), .ZN(n2842) );
  AOI21_X1 U3689 ( .B1(n4501), .B2(ADDR_REG_18__SCAN_IN), .A(n2842), .ZN(n2843) );
  INV_X1 U3690 ( .A(n2844), .ZN(n2845) );
  XNOR2_X1 U3691 ( .A(n2849), .B(n3808), .ZN(n3984) );
  INV_X1 U3692 ( .A(n4590), .ZN(n4250) );
  XNOR2_X1 U3693 ( .A(n2850), .B(n3808), .ZN(n2854) );
  AOI22_X1 U3694 ( .A1(n3914), .A2(n4175), .B1(n2851), .B2(n4530), .ZN(n2852)
         );
  OAI21_X1 U3695 ( .B1(n3729), .B2(n4267), .A(n2852), .ZN(n2853) );
  AOI21_X1 U3696 ( .B1(n2854), .B2(n4519), .A(n2853), .ZN(n3977) );
  OAI21_X1 U3697 ( .B1(n3984), .B2(n4250), .A(n3977), .ZN(n2860) );
  AND2_X2 U3698 ( .A1(n2855), .A2(n2912), .ZN(n4634) );
  INV_X1 U3699 ( .A(n2856), .ZN(n2859) );
  OAI21_X1 U3700 ( .B1(n3996), .B2(n3613), .A(n2857), .ZN(n3980) );
  NAND2_X1 U3701 ( .A1(n2859), .A2(n2858), .ZN(U3546) );
  INV_X1 U3702 ( .A(n2861), .ZN(n2863) );
  NAND2_X1 U3703 ( .A1(n2863), .A2(n2862), .ZN(U3514) );
  INV_X1 U3704 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2864) );
  INV_X1 U3705 ( .A(n4554), .ZN(n2867) );
  NOR2_X1 U3706 ( .A1(n2867), .A2(n2869), .ZN(U4043) );
  NOR2_X1 U3707 ( .A1(n2871), .A2(n4181), .ZN(n2930) );
  INV_X1 U3708 ( .A(n2930), .ZN(n2872) );
  XNOR2_X1 U3709 ( .A(n2873), .B(n3607), .ZN(n2950) );
  OAI22_X1 U3710 ( .A1(n2870), .A2(n3606), .B1(n3602), .B2(n3204), .ZN(n2949)
         );
  XNOR2_X1 U3711 ( .A(n2950), .B(n2949), .ZN(n2924) );
  NAND2_X1 U3712 ( .A1(n3591), .A2(n3832), .ZN(n2875) );
  XNOR2_X1 U3713 ( .A(n2877), .B(n3607), .ZN(n2879) );
  NOR2_X1 U3714 ( .A1(n2892), .A2(n3091), .ZN(n2878) );
  INV_X1 U3715 ( .A(n3085), .ZN(n2882) );
  INV_X1 U3716 ( .A(n2879), .ZN(n2881) );
  NAND2_X1 U3717 ( .A1(n2881), .A2(n2880), .ZN(n2907) );
  NAND2_X1 U3718 ( .A1(n3591), .A2(n3154), .ZN(n2884) );
  AND2_X1 U3719 ( .A1(n2885), .A2(n2884), .ZN(n2890) );
  INV_X1 U3720 ( .A(n2869), .ZN(n2887) );
  NAND2_X1 U3721 ( .A1(n2887), .A2(REG1_REG_0__SCAN_IN), .ZN(n2886) );
  NAND2_X1 U3722 ( .A1(n2890), .A2(n2886), .ZN(n3029) );
  AOI22_X1 U3723 ( .A1(n3564), .A2(n3154), .B1(n2887), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2888) );
  NAND2_X1 U3724 ( .A1(n2889), .A2(n2888), .ZN(n3028) );
  NAND2_X1 U3725 ( .A1(n3029), .A2(n3028), .ZN(n3027) );
  NAND2_X1 U3726 ( .A1(n2890), .A2(n3600), .ZN(n2891) );
  NAND2_X1 U3727 ( .A1(n3027), .A2(n2891), .ZN(n3068) );
  XNOR2_X1 U3728 ( .A(n2893), .B(n3600), .ZN(n2895) );
  NAND2_X1 U3729 ( .A1(n3068), .A2(n3066), .ZN(n3067) );
  INV_X1 U3730 ( .A(n2895), .ZN(n2897) );
  NAND2_X1 U3731 ( .A1(n2897), .A2(n2896), .ZN(n2898) );
  INV_X1 U3732 ( .A(n3077), .ZN(n2902) );
  OAI22_X1 U3733 ( .A1(n4536), .A2(n3606), .B1(n3602), .B2(n3171), .ZN(n2904)
         );
  XNOR2_X1 U3734 ( .A(n2903), .B(n2904), .ZN(n3079) );
  INV_X1 U3735 ( .A(n3079), .ZN(n2901) );
  INV_X1 U3736 ( .A(n2903), .ZN(n2906) );
  INV_X1 U3737 ( .A(n2904), .ZN(n2905) );
  NAND2_X1 U3738 ( .A1(n2906), .A2(n2905), .ZN(n3086) );
  NAND2_X1 U3739 ( .A1(n3086), .A2(n2907), .ZN(n2919) );
  INV_X1 U3740 ( .A(n2919), .ZN(n2908) );
  NAND2_X1 U3741 ( .A1(n2922), .A2(n2908), .ZN(n2909) );
  AND2_X1 U3742 ( .A1(n2920), .A2(n2909), .ZN(n2923) );
  AND2_X1 U3743 ( .A1(n2910), .A2(n3017), .ZN(n3149) );
  NAND3_X1 U3744 ( .A1(n3149), .A2(n2912), .A3(n2911), .ZN(n2939) );
  INV_X1 U3745 ( .A(n3146), .ZN(n3062) );
  INV_X1 U3746 ( .A(n2913), .ZN(n2914) );
  NAND2_X1 U3747 ( .A1(n3153), .A2(n2914), .ZN(n2916) );
  NAND2_X1 U3748 ( .A1(n2916), .A2(n2915), .ZN(n2925) );
  INV_X1 U3749 ( .A(n2925), .ZN(n2917) );
  NAND2_X1 U3750 ( .A1(n3062), .A2(n2917), .ZN(n2918) );
  NOR2_X1 U3751 ( .A1(n2919), .A2(n2924), .ZN(n2921) );
  AOI211_X1 U3752 ( .C1(n2924), .C2(n2923), .A(n3745), .B(n2246), .ZN(n2943)
         );
  NAND2_X1 U3753 ( .A1(n4265), .A2(n2925), .ZN(n2926) );
  NAND2_X1 U3754 ( .A1(n2939), .A2(n2926), .ZN(n2927) );
  NAND2_X1 U3755 ( .A1(n2927), .A2(n3148), .ZN(n3060) );
  NAND2_X1 U3756 ( .A1(n2869), .A2(n2928), .ZN(n2929) );
  OAI21_X1 U3757 ( .B1(n3060), .B2(n2929), .A(STATE_REG_SCAN_IN), .ZN(n2932)
         );
  NAND2_X1 U3758 ( .A1(n4554), .A2(n2930), .ZN(n2931) );
  NOR2_X1 U3759 ( .A1(n2892), .A2(n2931), .ZN(n3908) );
  NAND2_X1 U3760 ( .A1(n2939), .A2(n3908), .ZN(n3061) );
  NOR2_X1 U3761 ( .A1(n4360), .A2(n3206), .ZN(n2942) );
  NAND2_X1 U3762 ( .A1(n3908), .A2(n4343), .ZN(n2933) );
  AND2_X1 U3763 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3039) );
  INV_X1 U3764 ( .A(n3039), .ZN(n2934) );
  OAI21_X1 U3765 ( .B1(n3728), .B2(n3256), .A(n2934), .ZN(n2941) );
  NAND2_X1 U3766 ( .A1(n3062), .A2(n4530), .ZN(n2935) );
  OR2_X1 U3767 ( .A1(n2939), .A2(n2935), .ZN(n2937) );
  AND2_X2 U3768 ( .A1(n2937), .A2(n4129), .ZN(n4347) );
  INV_X1 U3769 ( .A(n4343), .ZN(n3033) );
  NAND2_X1 U3770 ( .A1(n3908), .A2(n3033), .ZN(n2938) );
  OAI22_X1 U3771 ( .A1(n4347), .A2(n3204), .B1(n3833), .B2(n4344), .ZN(n2940)
         );
  OR4_X1 U3772 ( .A1(n2943), .A2(n2942), .A3(n2941), .A4(n2940), .ZN(U3227) );
  NAND2_X1 U3773 ( .A1(n4511), .A2(n2883), .ZN(n2945) );
  NAND2_X1 U3774 ( .A1(n3591), .A2(n3322), .ZN(n2944) );
  NAND2_X1 U3775 ( .A1(n2945), .A2(n2944), .ZN(n2946) );
  XNOR2_X1 U3776 ( .A(n2946), .B(n3600), .ZN(n3347) );
  NOR2_X1 U3777 ( .A1(n3602), .A2(n3329), .ZN(n2948) );
  AOI21_X1 U3778 ( .B1(n2947), .B2(n4511), .A(n2948), .ZN(n3348) );
  XNOR2_X1 U3779 ( .A(n3347), .B(n3348), .ZN(n2998) );
  NAND2_X1 U3780 ( .A1(n2950), .A2(n2949), .ZN(n2951) );
  NAND2_X1 U3781 ( .A1(n3926), .A2(n3564), .ZN(n2953) );
  NAND2_X1 U3782 ( .A1(n3591), .A2(n3269), .ZN(n2952) );
  NAND2_X1 U3783 ( .A1(n2953), .A2(n2952), .ZN(n2954) );
  NOR2_X1 U3784 ( .A1(n3602), .A2(n3098), .ZN(n2955) );
  AOI21_X1 U3785 ( .B1(n2947), .B2(n3926), .A(n2955), .ZN(n2956) );
  INV_X1 U3786 ( .A(n2956), .ZN(n2957) );
  NAND2_X1 U3787 ( .A1(n2958), .A2(n2957), .ZN(n2959) );
  NAND2_X1 U3788 ( .A1(n2947), .A2(n3925), .ZN(n2961) );
  NAND2_X1 U3789 ( .A1(n2883), .A2(n3214), .ZN(n2960) );
  NAND2_X1 U3790 ( .A1(n2961), .A2(n2960), .ZN(n3123) );
  NAND2_X1 U3791 ( .A1(n3925), .A2(n3564), .ZN(n2963) );
  NAND2_X1 U3792 ( .A1(n3591), .A2(n3214), .ZN(n2962) );
  NAND2_X1 U3793 ( .A1(n2963), .A2(n2962), .ZN(n2964) );
  XNOR2_X1 U3794 ( .A(n2964), .B(n3607), .ZN(n3122) );
  OAI22_X1 U3795 ( .A1(n2965), .A2(n3602), .B1(n2899), .B2(n3192), .ZN(n2966)
         );
  XNOR2_X1 U3796 ( .A(n2966), .B(n3600), .ZN(n2967) );
  OAI22_X1 U3797 ( .A1(n2965), .A2(n3606), .B1(n3602), .B2(n3192), .ZN(n2968)
         );
  INV_X1 U3798 ( .A(n2967), .ZN(n2969) );
  INV_X1 U3799 ( .A(n3224), .ZN(n2976) );
  NAND2_X1 U3800 ( .A1(n3924), .A2(n2883), .ZN(n2971) );
  NAND2_X1 U3801 ( .A1(n3591), .A2(n3296), .ZN(n2970) );
  NAND2_X1 U3802 ( .A1(n2971), .A2(n2970), .ZN(n2972) );
  XNOR2_X1 U3803 ( .A(n2972), .B(n3607), .ZN(n2977) );
  NAND2_X1 U3804 ( .A1(n2947), .A2(n3924), .ZN(n2974) );
  NAND2_X1 U3805 ( .A1(n3564), .A2(n3296), .ZN(n2973) );
  NAND2_X1 U3806 ( .A1(n2974), .A2(n2973), .ZN(n2978) );
  NAND2_X1 U3807 ( .A1(n2976), .A2(n2975), .ZN(n2995) );
  INV_X1 U3808 ( .A(n2977), .ZN(n2980) );
  INV_X1 U3809 ( .A(n2978), .ZN(n2979) );
  NAND2_X1 U3810 ( .A1(n2980), .A2(n2979), .ZN(n3310) );
  NAND2_X1 U3811 ( .A1(n3923), .A2(n3564), .ZN(n2982) );
  NAND2_X1 U3812 ( .A1(n3591), .A2(n3282), .ZN(n2981) );
  NAND2_X1 U3813 ( .A1(n2982), .A2(n2981), .ZN(n2983) );
  XNOR2_X1 U3814 ( .A(n2983), .B(n3607), .ZN(n2988) );
  INV_X1 U3815 ( .A(n2988), .ZN(n2985) );
  NOR2_X1 U3816 ( .A1(n3602), .A2(n3338), .ZN(n2984) );
  AOI21_X1 U3817 ( .B1(n2947), .B2(n3923), .A(n2984), .ZN(n2987) );
  NAND2_X1 U3818 ( .A1(n2985), .A2(n2987), .ZN(n2986) );
  AND2_X1 U3819 ( .A1(n3310), .A2(n2986), .ZN(n2992) );
  NAND2_X1 U3820 ( .A1(n2995), .A2(n2992), .ZN(n2990) );
  INV_X1 U3821 ( .A(n2986), .ZN(n2989) );
  XNOR2_X1 U3822 ( .A(n2988), .B(n2987), .ZN(n3312) );
  AND2_X1 U3823 ( .A1(n2990), .A2(n2993), .ZN(n2997) );
  INV_X1 U3824 ( .A(n2998), .ZN(n2991) );
  AND2_X1 U3825 ( .A1(n2992), .A2(n2991), .ZN(n2994) );
  INV_X1 U3826 ( .A(n3352), .ZN(n2996) );
  AOI211_X1 U3827 ( .C1(n2998), .C2(n2997), .A(n3745), .B(n2996), .ZN(n3003)
         );
  NOR2_X1 U3828 ( .A1(n4360), .A2(n3332), .ZN(n3002) );
  NOR2_X1 U3829 ( .A1(STATE_REG_SCAN_IN), .A2(n4973), .ZN(n4432) );
  INV_X1 U3830 ( .A(n4432), .ZN(n2999) );
  OAI21_X1 U3831 ( .B1(n4344), .B2(n3324), .A(n2999), .ZN(n3001) );
  OAI22_X1 U3832 ( .A1(n4347), .A2(n3329), .B1(n3426), .B2(n3728), .ZN(n3000)
         );
  OR4_X1 U3833 ( .A1(n3003), .A2(n3002), .A3(n3001), .A4(n3000), .ZN(U3214) );
  INV_X1 U3834 ( .A(DATAI_1_), .ZN(n3004) );
  MUX2_X1 U3835 ( .A(n3005), .B(n3004), .S(U3149), .Z(n3006) );
  INV_X1 U3836 ( .A(n3006), .ZN(U3351) );
  NAND2_X1 U3837 ( .A1(U3149), .A2(DATAI_25_), .ZN(n3007) );
  OAI21_X1 U3838 ( .B1(n3008), .B2(U3149), .A(n3007), .ZN(U3327) );
  MUX2_X1 U3839 ( .A(n3954), .B(n2599), .S(U3149), .Z(n3009) );
  INV_X1 U3840 ( .A(n3009), .ZN(U3333) );
  INV_X1 U3841 ( .A(DATAI_27_), .ZN(n4793) );
  NAND2_X1 U3842 ( .A1(n4364), .A2(STATE_REG_SCAN_IN), .ZN(n3010) );
  OAI21_X1 U3843 ( .B1(STATE_REG_SCAN_IN), .B2(n4793), .A(n3010), .ZN(U3325)
         );
  INV_X1 U3844 ( .A(DATAI_21_), .ZN(n4732) );
  NAND2_X1 U3845 ( .A1(n2711), .A2(STATE_REG_SCAN_IN), .ZN(n3011) );
  OAI21_X1 U3846 ( .B1(STATE_REG_SCAN_IN), .B2(n4732), .A(n3011), .ZN(U3331)
         );
  INV_X1 U3847 ( .A(DATAI_29_), .ZN(n4878) );
  NAND2_X1 U3848 ( .A1(n3012), .A2(STATE_REG_SCAN_IN), .ZN(n3013) );
  OAI21_X1 U3849 ( .B1(STATE_REG_SCAN_IN), .B2(n4878), .A(n3013), .ZN(U3323)
         );
  NAND2_X1 U3850 ( .A1(n3014), .A2(n3062), .ZN(n4552) );
  INV_X1 U3851 ( .A(D_REG_0__SCAN_IN), .ZN(n4769) );
  INV_X1 U3852 ( .A(n3015), .ZN(n3016) );
  AOI22_X1 U3853 ( .A1(n4552), .A2(n4769), .B1(n3016), .B2(n4554), .ZN(U3458)
         );
  INV_X1 U3854 ( .A(D_REG_1__SCAN_IN), .ZN(n4962) );
  INV_X1 U3855 ( .A(n3017), .ZN(n3018) );
  AOI22_X1 U3856 ( .A1(n4552), .A2(n4962), .B1(n3018), .B2(n4554), .ZN(U3459)
         );
  NOR2_X1 U3857 ( .A1(n4501), .A2(n3928), .ZN(U3148) );
  XNOR2_X1 U3858 ( .A(n3019), .B(REG2_REG_3__SCAN_IN), .ZN(n3026) );
  INV_X1 U3859 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4885) );
  NOR2_X1 U3860 ( .A1(STATE_REG_SCAN_IN), .A2(n4885), .ZN(n3088) );
  NOR2_X1 U3861 ( .A1(n4508), .A2(n3020), .ZN(n3021) );
  AOI211_X1 U3862 ( .C1(n4501), .C2(ADDR_REG_3__SCAN_IN), .A(n3088), .B(n3021), 
        .ZN(n3025) );
  OAI211_X1 U3863 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3023), .A(n4502), .B(n3022), 
        .ZN(n3024) );
  OAI211_X1 U3864 ( .C1(n3026), .C2(n4495), .A(n3025), .B(n3024), .ZN(U3243)
         );
  OAI21_X1 U3865 ( .B1(n3029), .B2(n3028), .A(n3027), .ZN(n3072) );
  NAND3_X1 U3866 ( .A1(n3072), .A2(n3033), .A3(n3030), .ZN(n3035) );
  INV_X1 U3867 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3031) );
  NAND2_X1 U3868 ( .A1(n4364), .A2(n3031), .ZN(n3032) );
  NAND2_X1 U3869 ( .A1(n3033), .A2(n3032), .ZN(n4365) );
  AND2_X1 U3870 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3936)
         );
  AOI22_X1 U3871 ( .A1(n2266), .A2(n4365), .B1(n3907), .B2(n3936), .ZN(n3034)
         );
  NAND3_X1 U3872 ( .A1(n3035), .A2(n3928), .A3(n3034), .ZN(n3058) );
  XOR2_X1 U3873 ( .A(n3036), .B(REG2_REG_4__SCAN_IN), .Z(n3044) );
  OAI211_X1 U3874 ( .C1(REG1_REG_4__SCAN_IN), .C2(n3038), .A(n4502), .B(n3037), 
        .ZN(n3041) );
  AOI21_X1 U3875 ( .B1(n4501), .B2(ADDR_REG_4__SCAN_IN), .A(n3039), .ZN(n3040)
         );
  OAI211_X1 U3876 ( .C1(n4508), .C2(n3042), .A(n3041), .B(n3040), .ZN(n3043)
         );
  AOI21_X1 U3877 ( .B1(n4456), .B2(n3044), .A(n3043), .ZN(n3045) );
  NAND2_X1 U3878 ( .A1(n3058), .A2(n3045), .ZN(U3244) );
  INV_X1 U3879 ( .A(n4508), .ZN(n3930) );
  NAND2_X1 U3880 ( .A1(n4501), .A2(ADDR_REG_2__SCAN_IN), .ZN(n3046) );
  OAI21_X1 U3881 ( .B1(STATE_REG_SCAN_IN), .B2(n3168), .A(n3046), .ZN(n3057)
         );
  OAI211_X1 U3882 ( .C1(n3049), .C2(n3048), .A(n4502), .B(n3047), .ZN(n3055)
         );
  INV_X1 U3883 ( .A(n3050), .ZN(n3053) );
  NAND3_X1 U3884 ( .A1(n4456), .A2(n3053), .A3(n3052), .ZN(n3054) );
  NAND2_X1 U3885 ( .A1(n3055), .A2(n3054), .ZN(n3056) );
  AOI211_X1 U3886 ( .C1(n2221), .C2(n3930), .A(n3057), .B(n3056), .ZN(n3059)
         );
  NAND2_X1 U3887 ( .A1(n3059), .A2(n3058), .ZN(U3242) );
  INV_X1 U3888 ( .A(n3060), .ZN(n3063) );
  NAND3_X1 U3889 ( .A1(n3063), .A2(n3062), .A3(n3061), .ZN(n3082) );
  INV_X1 U3890 ( .A(n3082), .ZN(n3076) );
  INV_X1 U3891 ( .A(n4347), .ZN(n3725) );
  OAI22_X1 U3892 ( .A1(n3064), .A2(n4344), .B1(n3728), .B2(n4536), .ZN(n3065)
         );
  AOI21_X1 U3893 ( .B1(n4531), .B2(n3725), .A(n3065), .ZN(n3070) );
  OAI211_X1 U3894 ( .C1(n3066), .C2(n3068), .A(n3067), .B(n4355), .ZN(n3069)
         );
  OAI211_X1 U3895 ( .C1(n3076), .C2(n3071), .A(n3070), .B(n3069), .ZN(U3219)
         );
  OAI22_X1 U3896 ( .A1(n3072), .A2(n3745), .B1(n3728), .B2(n2894), .ZN(n3073)
         );
  AOI21_X1 U3897 ( .B1(n3154), .B2(n3725), .A(n3073), .ZN(n3074) );
  OAI21_X1 U3898 ( .B1(n3076), .B2(n3075), .A(n3074), .ZN(U3229) );
  INV_X1 U3899 ( .A(n2922), .ZN(n3078) );
  AOI21_X1 U3900 ( .B1(n3079), .B2(n3077), .A(n3078), .ZN(n3084) );
  AOI22_X1 U3901 ( .A1(n4350), .A2(n2874), .B1(n3738), .B2(n2401), .ZN(n3080)
         );
  OAI21_X1 U3902 ( .B1(n4347), .B2(n3171), .A(n3080), .ZN(n3081) );
  AOI21_X1 U3903 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3082), .A(n3081), .ZN(n3083)
         );
  OAI21_X1 U3904 ( .B1(n3084), .B2(n3745), .A(n3083), .ZN(U3234) );
  NAND2_X1 U3905 ( .A1(n2922), .A2(n3086), .ZN(n3087) );
  XOR2_X1 U3906 ( .A(n3085), .B(n3087), .Z(n3094) );
  AOI21_X1 U3907 ( .B1(n4350), .B2(n3927), .A(n3088), .ZN(n3090) );
  NAND2_X1 U3908 ( .A1(n3738), .A2(n2409), .ZN(n3089) );
  OAI211_X1 U3909 ( .C1(n4347), .C2(n3091), .A(n3090), .B(n3089), .ZN(n3092)
         );
  AOI21_X1 U3910 ( .B1(n3743), .B2(n4885), .A(n3092), .ZN(n3093) );
  OAI21_X1 U3911 ( .B1(n3094), .B2(n3745), .A(n3093), .ZN(U3215) );
  OAI211_X1 U3912 ( .C1(n3097), .C2(n3096), .A(n3095), .B(n4355), .ZN(n3103)
         );
  OAI22_X1 U3913 ( .A1(n4347), .A2(n3098), .B1(n3241), .B2(n3728), .ZN(n3101)
         );
  NOR2_X1 U3914 ( .A1(STATE_REG_SCAN_IN), .A2(n2433), .ZN(n4373) );
  INV_X1 U3915 ( .A(n4373), .ZN(n3099) );
  OAI21_X1 U3916 ( .B1(n4344), .B2(n2870), .A(n3099), .ZN(n3100) );
  NOR2_X1 U3917 ( .A1(n3101), .A2(n3100), .ZN(n3102) );
  OAI211_X1 U3918 ( .C1(n4360), .C2(n3268), .A(n3103), .B(n3102), .ZN(U3224)
         );
  INV_X1 U3919 ( .A(n3105), .ZN(n3822) );
  XNOR2_X1 U3920 ( .A(n3104), .B(n3822), .ZN(n3185) );
  INV_X1 U3921 ( .A(n3185), .ZN(n3110) );
  NAND3_X1 U3922 ( .A1(n3170), .A2(n2692), .A3(n3822), .ZN(n3106) );
  NAND2_X1 U3923 ( .A1(n3107), .A2(n3106), .ZN(n3108) );
  INV_X1 U3924 ( .A(n4516), .ZN(n4542) );
  AOI222_X1 U3925 ( .A1(n3108), .A2(n4519), .B1(n3927), .B2(n4175), .C1(n3185), 
        .C2(n4542), .ZN(n3187) );
  AOI22_X1 U3926 ( .A1(n2409), .A2(n4532), .B1(n4530), .B2(n3832), .ZN(n3109)
         );
  OAI211_X1 U3927 ( .C1(n3110), .C2(n4607), .A(n3187), .B(n3109), .ZN(n3119)
         );
  INV_X1 U3928 ( .A(n3205), .ZN(n3113) );
  INV_X1 U3929 ( .A(n3111), .ZN(n3167) );
  NAND2_X1 U3930 ( .A1(n3167), .A2(n3832), .ZN(n3112) );
  NAND2_X1 U3931 ( .A1(n3113), .A2(n3112), .ZN(n3183) );
  INV_X1 U3932 ( .A(REG1_REG_3__SCAN_IN), .ZN(n3114) );
  OAI22_X1 U3933 ( .A1(n4619), .A2(n3183), .B1(n4634), .B2(n3114), .ZN(n3115)
         );
  AOI21_X1 U3934 ( .B1(n3119), .B2(n4634), .A(n3115), .ZN(n3116) );
  INV_X1 U3935 ( .A(n3116), .ZN(U3521) );
  INV_X1 U3936 ( .A(REG0_REG_3__SCAN_IN), .ZN(n3117) );
  OAI22_X1 U3937 ( .A1(n4580), .A2(n3183), .B1(n4613), .B2(n3117), .ZN(n3118)
         );
  AOI21_X1 U3938 ( .B1(n3119), .B2(n4613), .A(n3118), .ZN(n3120) );
  INV_X1 U3939 ( .A(n3120), .ZN(U3473) );
  XOR2_X1 U3940 ( .A(n3123), .B(n3122), .Z(n3124) );
  XNOR2_X1 U3941 ( .A(n3121), .B(n3124), .ZN(n3132) );
  INV_X1 U3942 ( .A(n3254), .ZN(n3130) );
  INV_X1 U3943 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3125) );
  NOR2_X1 U3944 ( .A1(STATE_REG_SCAN_IN), .A2(n3125), .ZN(n4384) );
  AOI21_X1 U3945 ( .B1(n3738), .B2(n3926), .A(n4384), .ZN(n3128) );
  NAND2_X1 U3946 ( .A1(n4350), .A2(n3126), .ZN(n3127) );
  OAI211_X1 U3947 ( .C1(n4347), .C2(n3257), .A(n3128), .B(n3127), .ZN(n3129)
         );
  AOI21_X1 U3948 ( .B1(n3743), .B2(n3130), .A(n3129), .ZN(n3131) );
  OAI21_X1 U3949 ( .B1(n3132), .B2(n3745), .A(n3131), .ZN(U3236) );
  INV_X1 U3950 ( .A(n3134), .ZN(n3837) );
  AND2_X1 U3951 ( .A1(n3837), .A2(n3847), .ZN(n3818) );
  XOR2_X1 U3952 ( .A(n3133), .B(n3818), .Z(n3266) );
  XOR2_X1 U3953 ( .A(n3818), .B(n3135), .Z(n3136) );
  AOI22_X1 U3954 ( .A1(n3136), .A2(n4519), .B1(n4175), .B2(n3925), .ZN(n3276)
         );
  AOI22_X1 U3955 ( .A1(n3927), .A2(n4532), .B1(n4530), .B2(n3269), .ZN(n3137)
         );
  OAI211_X1 U3956 ( .C1(n3266), .C2(n4250), .A(n3276), .B(n3137), .ZN(n3142)
         );
  INV_X1 U3957 ( .A(n3142), .ZN(n3141) );
  INV_X1 U3958 ( .A(n4580), .ZN(n4324) );
  AND2_X1 U3959 ( .A1(n3138), .A2(n3269), .ZN(n3139) );
  NOR2_X1 U3960 ( .A1(n3217), .A2(n3139), .ZN(n3270) );
  AOI22_X1 U3961 ( .A1(n4324), .A2(n3270), .B1(REG0_REG_5__SCAN_IN), .B2(n4611), .ZN(n3140) );
  OAI21_X1 U3962 ( .B1(n3141), .B2(n4611), .A(n3140), .ZN(U3477) );
  INV_X1 U3963 ( .A(REG1_REG_5__SCAN_IN), .ZN(n3145) );
  NAND2_X1 U3964 ( .A1(n3142), .A2(n4634), .ZN(n3144) );
  INV_X1 U3965 ( .A(n4619), .ZN(n4255) );
  NAND2_X1 U3966 ( .A1(n4255), .A2(n3270), .ZN(n3143) );
  OAI211_X1 U3967 ( .C1(n4634), .C2(n3145), .A(n3144), .B(n3143), .ZN(U3523)
         );
  OAI21_X1 U3968 ( .B1(n4962), .B2(n3146), .A(n4552), .ZN(n3147) );
  NAND4_X1 U3969 ( .A1(n3150), .A2(n3149), .A3(n3148), .A4(n3147), .ZN(n3151)
         );
  NAND2_X2 U3970 ( .A1(n3151), .A2(n4129), .ZN(n4182) );
  OR2_X1 U3971 ( .A1(n3152), .A2(n3954), .ZN(n3246) );
  OR2_X1 U3972 ( .A1(n2222), .A2(n3246), .ZN(n4136) );
  NAND2_X1 U3973 ( .A1(n4533), .A2(n4546), .ZN(n3827) );
  INV_X1 U3974 ( .A(n3781), .ZN(n4570) );
  NAND2_X1 U3975 ( .A1(n3154), .A2(n3153), .ZN(n4568) );
  INV_X1 U3976 ( .A(n4519), .ZN(n4537) );
  NAND2_X1 U3977 ( .A1(n4516), .A2(n4537), .ZN(n3155) );
  AOI22_X1 U3978 ( .A1(n3781), .A2(n3155), .B1(n4175), .B2(n2401), .ZN(n4569)
         );
  OAI21_X1 U3979 ( .B1(n3156), .B2(n4568), .A(n4569), .ZN(n3157) );
  INV_X1 U3980 ( .A(n4129), .ZN(n4543) );
  AOI22_X1 U3981 ( .A1(n3157), .A2(n4182), .B1(REG3_REG_0__SCAN_IN), .B2(n4543), .ZN(n3159) );
  NAND2_X1 U3982 ( .A1(n2222), .A2(REG2_REG_0__SCAN_IN), .ZN(n3158) );
  OAI211_X1 U3983 ( .C1(n4136), .C2(n4570), .A(n3159), .B(n3158), .ZN(U3290)
         );
  INV_X1 U3984 ( .A(n4136), .ZN(n4549) );
  NAND2_X1 U3985 ( .A1(n3161), .A2(n3162), .ZN(n3163) );
  NAND2_X1 U3986 ( .A1(n3160), .A2(n3163), .ZN(n4578) );
  AND2_X1 U3987 ( .A1(n4169), .A2(n3954), .ZN(n3164) );
  NAND2_X1 U3988 ( .A1(n4544), .A2(n3165), .ZN(n3166) );
  NAND2_X1 U3989 ( .A1(n3167), .A2(n3166), .ZN(n4618) );
  OAI22_X1 U3990 ( .A1(n4159), .A2(n4618), .B1(n3168), .B2(n4129), .ZN(n3179)
         );
  NAND3_X1 U3991 ( .A1(n2690), .A2(n2689), .A3(n4539), .ZN(n3169) );
  NAND2_X1 U3992 ( .A1(n3170), .A2(n3169), .ZN(n3175) );
  NOR2_X1 U3993 ( .A1(n3171), .A2(n4265), .ZN(n3172) );
  AOI21_X1 U3994 ( .B1(n2874), .B2(n4175), .A(n3172), .ZN(n3173) );
  OAI21_X1 U3995 ( .B1(n2894), .B2(n4267), .A(n3173), .ZN(n3174) );
  AOI21_X1 U3996 ( .B1(n3175), .B2(n4519), .A(n3174), .ZN(n3177) );
  NAND2_X1 U3997 ( .A1(n4578), .A2(n4542), .ZN(n3176) );
  NAND2_X1 U3998 ( .A1(n3177), .A2(n3176), .ZN(n4577) );
  MUX2_X1 U3999 ( .A(REG2_REG_2__SCAN_IN), .B(n4577), .S(n4182), .Z(n3178) );
  AOI211_X1 U4000 ( .C1(n4549), .C2(n4578), .A(n3179), .B(n3178), .ZN(n3180)
         );
  INV_X1 U4001 ( .A(n3180), .ZN(U3288) );
  NAND2_X1 U4002 ( .A1(n4182), .A2(n4532), .ZN(n4107) );
  INV_X1 U4003 ( .A(n4107), .ZN(n3992) );
  AOI22_X1 U4004 ( .A1(n3992), .A2(n2409), .B1(n4111), .B2(n3832), .ZN(n3182)
         );
  AOI22_X1 U4005 ( .A1(n2222), .A2(REG2_REG_3__SCAN_IN), .B1(n4543), .B2(n4885), .ZN(n3181) );
  OAI211_X1 U4006 ( .C1(n4159), .C2(n3183), .A(n3182), .B(n3181), .ZN(n3184)
         );
  AOI21_X1 U4007 ( .B1(n4549), .B2(n3185), .A(n3184), .ZN(n3186) );
  OAI21_X1 U4008 ( .B1(n3187), .B2(n2222), .A(n3186), .ZN(U3287) );
  XNOR2_X1 U4009 ( .A(n3188), .B(n3189), .ZN(n3196) );
  INV_X1 U4010 ( .A(n3248), .ZN(n3194) );
  AND2_X1 U4011 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n4396) );
  AOI21_X1 U4012 ( .B1(n4350), .B2(n3924), .A(n4396), .ZN(n3191) );
  NAND2_X1 U4013 ( .A1(n3738), .A2(n3925), .ZN(n3190) );
  OAI211_X1 U4014 ( .C1(n4347), .C2(n3192), .A(n3191), .B(n3190), .ZN(n3193)
         );
  AOI21_X1 U4015 ( .B1(n3743), .B2(n3194), .A(n3193), .ZN(n3195) );
  OAI21_X1 U4016 ( .B1(n3196), .B2(n3745), .A(n3195), .ZN(U3210) );
  XNOR2_X1 U4017 ( .A(n3784), .B(n3197), .ZN(n3208) );
  XOR2_X1 U4018 ( .A(n3784), .B(n3198), .Z(n3202) );
  AOI22_X1 U4019 ( .A1(n3926), .A2(n4175), .B1(n3199), .B2(n4530), .ZN(n3200)
         );
  OAI21_X1 U4020 ( .B1(n3833), .B2(n4267), .A(n3200), .ZN(n3201) );
  AOI21_X1 U4021 ( .B1(n3202), .B2(n4519), .A(n3201), .ZN(n3203) );
  OAI21_X1 U4022 ( .B1(n3208), .B2(n4516), .A(n3203), .ZN(n4584) );
  OAI211_X1 U4023 ( .C1(n3205), .C2(n3204), .A(n4169), .B(n3138), .ZN(n4583)
         );
  OAI22_X1 U4024 ( .A1(n4583), .A2(n4181), .B1(n4129), .B2(n3206), .ZN(n3207)
         );
  OAI21_X1 U4025 ( .B1(n4584), .B2(n3207), .A(n4182), .ZN(n3210) );
  INV_X1 U4026 ( .A(n3208), .ZN(n4586) );
  AOI22_X1 U4027 ( .A1(n4586), .A2(n4549), .B1(REG2_REG_4__SCAN_IN), .B2(n2222), .ZN(n3209) );
  NAND2_X1 U4028 ( .A1(n3210), .A2(n3209), .ZN(U3286) );
  NAND2_X1 U4029 ( .A1(n3840), .A2(n3848), .ZN(n3783) );
  XOR2_X1 U4030 ( .A(n3783), .B(n3211), .Z(n3261) );
  XOR2_X1 U4031 ( .A(n3212), .B(n3783), .Z(n3213) );
  AOI22_X1 U4032 ( .A1(n3213), .A2(n4519), .B1(n4175), .B2(n3126), .ZN(n3265)
         );
  AOI22_X1 U4033 ( .A1(n3926), .A2(n4532), .B1(n3214), .B2(n4530), .ZN(n3215)
         );
  OAI211_X1 U4034 ( .C1(n3261), .C2(n4250), .A(n3265), .B(n3215), .ZN(n3222)
         );
  OR2_X1 U4035 ( .A1(n3217), .A2(n3257), .ZN(n3218) );
  NAND2_X1 U4036 ( .A1(n3216), .A2(n3218), .ZN(n3253) );
  INV_X1 U4037 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4896) );
  OAI22_X1 U4038 ( .A1(n3253), .A2(n4580), .B1(n4613), .B2(n4896), .ZN(n3219)
         );
  AOI21_X1 U4039 ( .B1(n3222), .B2(n4613), .A(n3219), .ZN(n3220) );
  INV_X1 U4040 ( .A(n3220), .ZN(U3479) );
  OAI22_X1 U4041 ( .A1(n3253), .A2(n4619), .B1(n4634), .B2(n4383), .ZN(n3221)
         );
  AOI21_X1 U4042 ( .B1(n3222), .B2(n4634), .A(n3221), .ZN(n3223) );
  INV_X1 U40430 ( .A(n3223), .ZN(U3524) );
  INV_X1 U4044 ( .A(n3310), .ZN(n3226) );
  NOR2_X1 U4045 ( .A1(n3226), .A2(n3225), .ZN(n3227) );
  XNOR2_X1 U4046 ( .A(n3224), .B(n3227), .ZN(n3233) );
  INV_X1 U4047 ( .A(n3304), .ZN(n3231) );
  INV_X1 U4048 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4968) );
  NOR2_X1 U4049 ( .A1(STATE_REG_SCAN_IN), .A2(n4968), .ZN(n4411) );
  AOI21_X1 U4050 ( .B1(n4350), .B2(n3923), .A(n4411), .ZN(n3229) );
  NAND2_X1 U4051 ( .A1(n3738), .A2(n3126), .ZN(n3228) );
  OAI211_X1 U4052 ( .C1(n4347), .C2(n3302), .A(n3229), .B(n3228), .ZN(n3230)
         );
  AOI21_X1 U4053 ( .B1(n3743), .B2(n3231), .A(n3230), .ZN(n3232) );
  OAI21_X1 U4054 ( .B1(n3233), .B2(n3745), .A(n3232), .ZN(U3218) );
  INV_X1 U4055 ( .A(n3234), .ZN(n3303) );
  AOI211_X1 U4056 ( .C1(n3238), .C2(n3216), .A(n4606), .B(n3303), .ZN(n4589)
         );
  INV_X1 U4057 ( .A(n3785), .ZN(n3235) );
  XNOR2_X1 U4058 ( .A(n3236), .B(n3235), .ZN(n3237) );
  NAND2_X1 U4059 ( .A1(n3237), .A2(n4519), .ZN(n3240) );
  AOI22_X1 U4060 ( .A1(n3924), .A2(n4175), .B1(n4530), .B2(n3238), .ZN(n3239)
         );
  OAI211_X1 U4061 ( .C1(n3241), .C2(n4267), .A(n3240), .B(n3239), .ZN(n4588)
         );
  AOI21_X1 U4062 ( .B1(n4589), .B2(n3954), .A(n4588), .ZN(n3252) );
  OR2_X1 U4063 ( .A1(n3211), .A2(n3242), .ZN(n3244) );
  NAND2_X1 U4064 ( .A1(n3244), .A2(n3243), .ZN(n3245) );
  XOR2_X1 U4065 ( .A(n3785), .B(n3245), .Z(n4591) );
  NAND2_X1 U4066 ( .A1(n4516), .A2(n3246), .ZN(n3247) );
  NAND2_X1 U4067 ( .A1(n4182), .A2(n3247), .ZN(n4186) );
  OAI22_X1 U4068 ( .A1(n4182), .A2(n3249), .B1(n3248), .B2(n4129), .ZN(n3250)
         );
  AOI21_X1 U4069 ( .B1(n4591), .B2(n4161), .A(n3250), .ZN(n3251) );
  OAI21_X1 U4070 ( .B1(n3252), .B2(n2222), .A(n3251), .ZN(U3283) );
  INV_X1 U4071 ( .A(n3253), .ZN(n3260) );
  INV_X1 U4072 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3255) );
  OAI22_X1 U4073 ( .A1(n4182), .A2(n3255), .B1(n3254), .B2(n4129), .ZN(n3259)
         );
  INV_X1 U4074 ( .A(n4111), .ZN(n3283) );
  OAI22_X1 U4075 ( .A1(n3283), .A2(n3257), .B1(n3256), .B2(n4107), .ZN(n3258)
         );
  AOI211_X1 U4076 ( .C1(n4548), .C2(n3260), .A(n3259), .B(n3258), .ZN(n3264)
         );
  INV_X1 U4077 ( .A(n3261), .ZN(n3262) );
  NAND2_X1 U4078 ( .A1(n3262), .A2(n4161), .ZN(n3263) );
  OAI211_X1 U4079 ( .C1(n3265), .C2(n2222), .A(n3264), .B(n3263), .ZN(U3284)
         );
  INV_X1 U4080 ( .A(n3266), .ZN(n3274) );
  OAI22_X1 U4081 ( .A1(n3268), .A2(n4129), .B1(n3267), .B2(n4182), .ZN(n3273)
         );
  AOI22_X1 U4082 ( .A1(n4548), .A2(n3270), .B1(n4111), .B2(n3269), .ZN(n3271)
         );
  OAI21_X1 U4083 ( .B1(n2870), .B2(n4107), .A(n3271), .ZN(n3272) );
  AOI211_X1 U4084 ( .C1(n3274), .C2(n4161), .A(n3273), .B(n3272), .ZN(n3275)
         );
  OAI21_X1 U4085 ( .B1(n2222), .B2(n3276), .A(n3275), .ZN(U3285) );
  INV_X1 U4086 ( .A(n3277), .ZN(n3858) );
  AND2_X1 U4087 ( .A1(n3858), .A2(n3845), .ZN(n3795) );
  XNOR2_X1 U4088 ( .A(n3278), .B(n3795), .ZN(n3280) );
  OAI22_X1 U4089 ( .A1(n3280), .A2(n4537), .B1(n3279), .B2(n4535), .ZN(n3340)
         );
  INV_X1 U4090 ( .A(n3340), .ZN(n3290) );
  INV_X1 U4091 ( .A(n4592), .ZN(n3281) );
  AOI21_X1 U4092 ( .B1(n3282), .B2(n3281), .A(n3330), .ZN(n3344) );
  OAI22_X1 U4093 ( .A1(n3283), .A2(n3338), .B1(n3339), .B2(n4107), .ZN(n3286)
         );
  OAI22_X1 U4094 ( .A1(n3313), .A2(n4129), .B1(n3284), .B2(n4182), .ZN(n3285)
         );
  AOI211_X1 U4095 ( .C1(n3344), .C2(n4548), .A(n3286), .B(n3285), .ZN(n3289)
         );
  XOR2_X1 U4096 ( .A(n3795), .B(n3287), .Z(n3342) );
  NAND2_X1 U4097 ( .A1(n3342), .A2(n4161), .ZN(n3288) );
  OAI211_X1 U4098 ( .C1(n3290), .C2(n2222), .A(n3289), .B(n3288), .ZN(U3281)
         );
  AND2_X1 U4099 ( .A1(n3844), .A2(n3849), .ZN(n3794) );
  OR2_X1 U4100 ( .A1(n3211), .A2(n3291), .ZN(n3293) );
  NAND2_X1 U4101 ( .A1(n3293), .A2(n3292), .ZN(n3294) );
  XOR2_X1 U4102 ( .A(n3794), .B(n3294), .Z(n3301) );
  XOR2_X1 U4103 ( .A(n3794), .B(n3295), .Z(n3299) );
  AOI22_X1 U4104 ( .A1(n3923), .A2(n4175), .B1(n3296), .B2(n4530), .ZN(n3297)
         );
  OAI21_X1 U4105 ( .B1(n2965), .B2(n4267), .A(n3297), .ZN(n3298) );
  AOI21_X1 U4106 ( .B1(n3299), .B2(n4519), .A(n3298), .ZN(n3300) );
  OAI21_X1 U4107 ( .B1(n3301), .B2(n4516), .A(n3300), .ZN(n4594) );
  INV_X1 U4108 ( .A(n4594), .ZN(n3309) );
  INV_X1 U4109 ( .A(n3301), .ZN(n4596) );
  NOR2_X1 U4110 ( .A1(n3303), .A2(n3302), .ZN(n4593) );
  NOR3_X1 U4111 ( .A1(n4593), .A2(n4592), .A3(n4159), .ZN(n3307) );
  INV_X1 U4112 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3305) );
  OAI22_X1 U4113 ( .A1(n4182), .A2(n3305), .B1(n3304), .B2(n4129), .ZN(n3306)
         );
  AOI211_X1 U4114 ( .C1(n4596), .C2(n4549), .A(n3307), .B(n3306), .ZN(n3308)
         );
  OAI21_X1 U4115 ( .B1(n3309), .B2(n2222), .A(n3308), .ZN(U3282) );
  NAND2_X1 U4116 ( .A1(n2995), .A2(n3310), .ZN(n3311) );
  XOR2_X1 U4117 ( .A(n3312), .B(n3311), .Z(n3319) );
  INV_X1 U4118 ( .A(n3313), .ZN(n3317) );
  NOR2_X1 U4119 ( .A1(STATE_REG_SCAN_IN), .A2(n2476), .ZN(n4422) );
  AOI21_X1 U4120 ( .B1(n4350), .B2(n4511), .A(n4422), .ZN(n3315) );
  NAND2_X1 U4121 ( .A1(n3738), .A2(n3924), .ZN(n3314) );
  OAI211_X1 U4122 ( .C1(n4347), .C2(n3338), .A(n3315), .B(n3314), .ZN(n3316)
         );
  AOI21_X1 U4123 ( .B1(n3743), .B2(n3317), .A(n3316), .ZN(n3318) );
  OAI21_X1 U4124 ( .B1(n3319), .B2(n3745), .A(n3318), .ZN(U3228) );
  AND2_X1 U4125 ( .A1(n3855), .A2(n3860), .ZN(n3796) );
  XOR2_X1 U4126 ( .A(n3796), .B(n3320), .Z(n3328) );
  XNOR2_X1 U4127 ( .A(n3321), .B(n3796), .ZN(n3326) );
  AOI22_X1 U4128 ( .A1(n3922), .A2(n4175), .B1(n3322), .B2(n4530), .ZN(n3323)
         );
  OAI21_X1 U4129 ( .B1(n3324), .B2(n4267), .A(n3323), .ZN(n3325) );
  AOI21_X1 U4130 ( .B1(n3326), .B2(n4519), .A(n3325), .ZN(n3327) );
  OAI21_X1 U4131 ( .B1(n3328), .B2(n4516), .A(n3327), .ZN(n4599) );
  INV_X1 U4132 ( .A(n4599), .ZN(n3337) );
  INV_X1 U4133 ( .A(n3328), .ZN(n4602) );
  NOR2_X1 U4134 ( .A1(n3330), .A2(n3329), .ZN(n4598) );
  INV_X1 U4135 ( .A(n3331), .ZN(n4597) );
  NOR3_X1 U4136 ( .A1(n4598), .A2(n4597), .A3(n4159), .ZN(n3335) );
  INV_X1 U4137 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3333) );
  OAI22_X1 U4138 ( .A1(n4182), .A2(n3333), .B1(n3332), .B2(n4129), .ZN(n3334)
         );
  AOI211_X1 U4139 ( .C1(n4602), .C2(n4549), .A(n3335), .B(n3334), .ZN(n3336)
         );
  OAI21_X1 U4140 ( .B1(n3337), .B2(n2222), .A(n3336), .ZN(U3280) );
  OAI22_X1 U4141 ( .A1(n3339), .A2(n4267), .B1(n4265), .B2(n3338), .ZN(n3341)
         );
  AOI211_X1 U4142 ( .C1(n4590), .C2(n3342), .A(n3341), .B(n3340), .ZN(n3346)
         );
  AOI22_X1 U4143 ( .A1(n3344), .A2(n4255), .B1(REG1_REG_9__SCAN_IN), .B2(n4631), .ZN(n3343) );
  OAI21_X1 U4144 ( .B1(n3346), .B2(n4631), .A(n3343), .ZN(U3527) );
  AOI22_X1 U4145 ( .A1(n3344), .A2(n4324), .B1(REG0_REG_9__SCAN_IN), .B2(n4611), .ZN(n3345) );
  OAI21_X1 U4146 ( .B1(n3346), .B2(n4611), .A(n3345), .ZN(U3485) );
  INV_X1 U4147 ( .A(n3347), .ZN(n3350) );
  INV_X1 U4148 ( .A(n3348), .ZN(n3349) );
  NAND2_X1 U4149 ( .A1(n3350), .A2(n3349), .ZN(n3351) );
  NAND2_X1 U4150 ( .A1(n3352), .A2(n3351), .ZN(n3384) );
  OAI22_X1 U4151 ( .A1(n3426), .A2(n3602), .B1(n2899), .B2(n4523), .ZN(n3353)
         );
  XNOR2_X1 U4152 ( .A(n3353), .B(n3600), .ZN(n3396) );
  NOR2_X1 U4153 ( .A1(n3602), .A2(n4523), .ZN(n3354) );
  AOI21_X1 U4154 ( .B1(n3922), .B2(n2947), .A(n3354), .ZN(n3394) );
  INV_X1 U4155 ( .A(n3394), .ZN(n3393) );
  XNOR2_X1 U4156 ( .A(n3396), .B(n3393), .ZN(n3355) );
  XNOR2_X1 U4157 ( .A(n3384), .B(n3355), .ZN(n3361) );
  INV_X1 U4158 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3356) );
  NOR2_X1 U4159 ( .A1(STATE_REG_SCAN_IN), .A2(n3356), .ZN(n4443) );
  AOI21_X1 U4160 ( .B1(n4350), .B2(n3921), .A(n4443), .ZN(n3358) );
  NAND2_X1 U4161 ( .A1(n3738), .A2(n4511), .ZN(n3357) );
  OAI211_X1 U4162 ( .C1(n4347), .C2(n4523), .A(n3358), .B(n3357), .ZN(n3359)
         );
  AOI21_X1 U4163 ( .B1(n3743), .B2(n4521), .A(n3359), .ZN(n3360) );
  OAI21_X1 U4164 ( .B1(n3361), .B2(n3745), .A(n3360), .ZN(U3233) );
  INV_X1 U4165 ( .A(n3408), .ZN(n3362) );
  OR2_X1 U4166 ( .A1(n3362), .A2(n3864), .ZN(n3366) );
  XNOR2_X1 U4167 ( .A(n3363), .B(n3366), .ZN(n3364) );
  OAI22_X1 U4168 ( .A1(n3364), .A2(n4537), .B1(n4268), .B2(n4535), .ZN(n3427)
         );
  INV_X1 U4169 ( .A(n3427), .ZN(n3375) );
  INV_X1 U4170 ( .A(n3366), .ZN(n3797) );
  XNOR2_X1 U4171 ( .A(n3365), .B(n3797), .ZN(n3429) );
  NAND2_X1 U4172 ( .A1(n4522), .A2(n3371), .ZN(n3367) );
  NAND2_X1 U4173 ( .A1(n3414), .A2(n3367), .ZN(n3435) );
  INV_X1 U4174 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3368) );
  OAI22_X1 U4175 ( .A1(n4182), .A2(n3368), .B1(n3407), .B2(n4129), .ZN(n3370)
         );
  NOR2_X1 U4176 ( .A1(n4107), .A2(n3426), .ZN(n3369) );
  AOI211_X1 U4177 ( .C1(n4111), .C2(n3371), .A(n3370), .B(n3369), .ZN(n3372)
         );
  OAI21_X1 U4178 ( .B1(n3435), .B2(n4159), .A(n3372), .ZN(n3373) );
  AOI21_X1 U4179 ( .B1(n3429), .B2(n4161), .A(n3373), .ZN(n3374) );
  OAI21_X1 U4180 ( .B1(n3375), .B2(n2222), .A(n3374), .ZN(U3278) );
  OAI22_X1 U4181 ( .A1(n4513), .A2(n3602), .B1(n2899), .B2(n3425), .ZN(n3376)
         );
  XNOR2_X1 U4182 ( .A(n3376), .B(n3607), .ZN(n3377) );
  OAI22_X1 U4183 ( .A1(n4513), .A2(n3606), .B1(n3602), .B2(n3425), .ZN(n3378)
         );
  NAND2_X1 U4184 ( .A1(n3377), .A2(n3378), .ZN(n3399) );
  OAI21_X1 U4185 ( .B1(n3396), .B2(n3394), .A(n3399), .ZN(n3383) );
  NAND3_X1 U4186 ( .A1(n3399), .A2(n3394), .A3(n3396), .ZN(n3381) );
  INV_X1 U4187 ( .A(n3377), .ZN(n3380) );
  INV_X1 U4188 ( .A(n3378), .ZN(n3379) );
  NAND2_X1 U4189 ( .A1(n3380), .A2(n3379), .ZN(n3398) );
  OAI22_X1 U4190 ( .A1(n4268), .A2(n3602), .B1(n2899), .B2(n3496), .ZN(n3385)
         );
  XNOR2_X1 U4191 ( .A(n3385), .B(n3600), .ZN(n3438) );
  XOR2_X1 U4192 ( .A(n3436), .B(n3438), .Z(n3386) );
  XNOR2_X1 U4193 ( .A(n3437), .B(n3386), .ZN(n3392) );
  INV_X1 U4194 ( .A(n3387), .ZN(n3417) );
  NOR2_X1 U4195 ( .A1(STATE_REG_SCAN_IN), .A2(n2523), .ZN(n4461) );
  AOI21_X1 U4196 ( .B1(n3738), .B2(n3921), .A(n4461), .ZN(n3389) );
  NAND2_X1 U4197 ( .A1(n4350), .A2(n3919), .ZN(n3388) );
  OAI211_X1 U4198 ( .C1(n4347), .C2(n3496), .A(n3389), .B(n3388), .ZN(n3390)
         );
  AOI21_X1 U4199 ( .B1(n3743), .B2(n3417), .A(n3390), .ZN(n3391) );
  OAI21_X1 U4200 ( .B1(n3392), .B2(n3745), .A(n3391), .ZN(U3231) );
  NOR2_X1 U4201 ( .A1(n3384), .A2(n3393), .ZN(n3397) );
  INV_X1 U4202 ( .A(n3384), .ZN(n3395) );
  OAI22_X1 U4203 ( .A1(n3397), .A2(n3396), .B1(n3395), .B2(n3394), .ZN(n3401)
         );
  NAND2_X1 U4204 ( .A1(n3399), .A2(n3398), .ZN(n3400) );
  XNOR2_X1 U4205 ( .A(n3401), .B(n3400), .ZN(n3402) );
  NAND2_X1 U4206 ( .A1(n3402), .A2(n4355), .ZN(n3406) );
  OAI22_X1 U4207 ( .A1(n4347), .A2(n3425), .B1(n4268), .B2(n3728), .ZN(n3404)
         );
  NAND2_X1 U4208 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4447) );
  OAI21_X1 U4209 ( .B1(n4344), .B2(n3426), .A(n4447), .ZN(n3403) );
  NOR2_X1 U4210 ( .A1(n3404), .A2(n3403), .ZN(n3405) );
  OAI211_X1 U4211 ( .C1(n4360), .C2(n3407), .A(n3406), .B(n3405), .ZN(U3221)
         );
  NAND2_X1 U4212 ( .A1(n3409), .A2(n3408), .ZN(n3411) );
  AND2_X1 U4213 ( .A1(n3867), .A2(n3410), .ZN(n3817) );
  XNOR2_X1 U4214 ( .A(n3411), .B(n3817), .ZN(n3412) );
  OAI22_X1 U4215 ( .A1(n3412), .A2(n4537), .B1(n4258), .B2(n4535), .ZN(n3497)
         );
  INV_X1 U4216 ( .A(n3497), .ZN(n3424) );
  XNOR2_X1 U4217 ( .A(n3413), .B(n3817), .ZN(n3499) );
  INV_X1 U4218 ( .A(n3414), .ZN(n3416) );
  INV_X1 U4219 ( .A(n3461), .ZN(n3415) );
  OAI21_X1 U4220 ( .B1(n3416), .B2(n3496), .A(n3415), .ZN(n3504) );
  NOR2_X1 U4221 ( .A1(n3504), .A2(n4159), .ZN(n3422) );
  AOI22_X1 U4222 ( .A1(n2222), .A2(REG2_REG_13__SCAN_IN), .B1(n3417), .B2(
        n4543), .ZN(n3420) );
  NAND2_X1 U4223 ( .A1(n4111), .A2(n3418), .ZN(n3419) );
  OAI211_X1 U4224 ( .C1(n4513), .C2(n4107), .A(n3420), .B(n3419), .ZN(n3421)
         );
  AOI211_X1 U4225 ( .C1(n3499), .C2(n4161), .A(n3422), .B(n3421), .ZN(n3423)
         );
  OAI21_X1 U4226 ( .B1(n2222), .B2(n3424), .A(n3423), .ZN(U3277) );
  INV_X1 U4227 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3430) );
  OAI22_X1 U4228 ( .A1(n3426), .A2(n4267), .B1(n3425), .B2(n4265), .ZN(n3428)
         );
  AOI211_X1 U4229 ( .C1(n4590), .C2(n3429), .A(n3428), .B(n3427), .ZN(n3432)
         );
  MUX2_X1 U4230 ( .A(n3430), .B(n3432), .S(n4634), .Z(n3431) );
  OAI21_X1 U4231 ( .B1(n3435), .B2(n4619), .A(n3431), .ZN(U3530) );
  INV_X1 U4232 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3433) );
  MUX2_X1 U4233 ( .A(n3433), .B(n3432), .S(n4613), .Z(n3434) );
  OAI21_X1 U4234 ( .B1(n3435), .B2(n4580), .A(n3434), .ZN(U3491) );
  OAI22_X1 U4235 ( .A1(n4258), .A2(n3602), .B1(n2899), .B2(n4266), .ZN(n3439)
         );
  XNOR2_X1 U4236 ( .A(n3439), .B(n3600), .ZN(n3444) );
  INV_X1 U4237 ( .A(n3444), .ZN(n3442) );
  NOR2_X1 U4238 ( .A1(n3602), .A2(n4266), .ZN(n3440) );
  AOI21_X1 U4239 ( .B1(n3919), .B2(n2947), .A(n3440), .ZN(n3443) );
  INV_X1 U4240 ( .A(n3443), .ZN(n3441) );
  NAND2_X1 U4241 ( .A1(n3442), .A2(n3441), .ZN(n3518) );
  AND2_X1 U4242 ( .A1(n3444), .A2(n3443), .ZN(n3517) );
  NOR2_X1 U4243 ( .A1(n2340), .A2(n3517), .ZN(n3445) );
  XNOR2_X1 U4244 ( .A(n3519), .B(n3445), .ZN(n3446) );
  NAND2_X1 U4245 ( .A1(n3446), .A2(n4355), .ZN(n3450) );
  OAI22_X1 U4246 ( .A1(n4347), .A2(n4266), .B1(n4268), .B2(n4344), .ZN(n3448)
         );
  NAND2_X1 U4247 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4467) );
  OAI21_X1 U4248 ( .B1(n3728), .B2(n4345), .A(n4467), .ZN(n3447) );
  NOR2_X1 U4249 ( .A1(n3448), .A2(n3447), .ZN(n3449) );
  OAI211_X1 U4250 ( .C1(n4360), .C2(n3457), .A(n3450), .B(n3449), .ZN(U3212)
         );
  NAND2_X1 U4251 ( .A1(n3451), .A2(n3452), .ZN(n3453) );
  NOR2_X1 U4252 ( .A1(n3453), .A2(n3454), .ZN(n3468) );
  AOI21_X1 U4253 ( .B1(n3454), .B2(n3453), .A(n3468), .ZN(n4264) );
  OAI21_X1 U4254 ( .B1(n3454), .B2(n3750), .A(n3470), .ZN(n3455) );
  AOI22_X1 U4255 ( .A1(n3455), .A2(n4519), .B1(n4175), .B2(n3918), .ZN(n3456)
         );
  OAI21_X1 U4256 ( .B1(n4264), .B2(n4516), .A(n3456), .ZN(n4269) );
  NAND2_X1 U4257 ( .A1(n4269), .A2(n4182), .ZN(n3466) );
  INV_X1 U4258 ( .A(n3457), .ZN(n3458) );
  AOI22_X1 U4259 ( .A1(n2222), .A2(REG2_REG_14__SCAN_IN), .B1(n3458), .B2(
        n4543), .ZN(n3459) );
  OAI21_X1 U4260 ( .B1(n4268), .B2(n4107), .A(n3459), .ZN(n3463) );
  OAI21_X1 U4261 ( .B1(n3461), .B2(n4266), .A(n3460), .ZN(n4334) );
  NOR2_X1 U4262 ( .A1(n4334), .A2(n4159), .ZN(n3462) );
  AOI211_X1 U4263 ( .C1(n4111), .C2(n3464), .A(n3463), .B(n3462), .ZN(n3465)
         );
  OAI211_X1 U4264 ( .C1(n4264), .C2(n4136), .A(n3466), .B(n3465), .ZN(U3276)
         );
  NOR2_X1 U4265 ( .A1(n3468), .A2(n3467), .ZN(n3469) );
  XOR2_X1 U4266 ( .A(n3782), .B(n3469), .Z(n4261) );
  INV_X1 U4267 ( .A(n4261), .ZN(n3480) );
  NAND2_X1 U4268 ( .A1(n3470), .A2(n3868), .ZN(n3471) );
  XNOR2_X1 U4269 ( .A(n3471), .B(n3782), .ZN(n3472) );
  OAI22_X1 U4270 ( .A1(n3472), .A2(n4537), .B1(n4244), .B2(n4535), .ZN(n4260)
         );
  NAND2_X1 U4271 ( .A1(n3460), .A2(n3520), .ZN(n3473) );
  NAND2_X1 U4272 ( .A1(n3487), .A2(n3473), .ZN(n4330) );
  INV_X1 U4273 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3474) );
  OAI22_X1 U4274 ( .A1(n4182), .A2(n3474), .B1(n3737), .B2(n4129), .ZN(n3476)
         );
  NOR2_X1 U4275 ( .A1(n4107), .A2(n4258), .ZN(n3475) );
  AOI211_X1 U4276 ( .C1(n4111), .C2(n3520), .A(n3476), .B(n3475), .ZN(n3477)
         );
  OAI21_X1 U4277 ( .B1(n4330), .B2(n4159), .A(n3477), .ZN(n3478) );
  AOI21_X1 U4278 ( .B1(n4260), .B2(n4182), .A(n3478), .ZN(n3479) );
  OAI21_X1 U4279 ( .B1(n3480), .B2(n4186), .A(n3479), .ZN(U3275) );
  XNOR2_X1 U4280 ( .A(n3481), .B(n2561), .ZN(n3485) );
  NAND2_X1 U4281 ( .A1(n3486), .A2(n4530), .ZN(n3483) );
  NAND2_X1 U4282 ( .A1(n3918), .A2(n4532), .ZN(n3482) );
  OAI211_X1 U4283 ( .C1(n4178), .C2(n4535), .A(n3483), .B(n3482), .ZN(n3484)
         );
  AOI21_X1 U4284 ( .B1(n3485), .B2(n4519), .A(n3484), .ZN(n4253) );
  AND2_X1 U4285 ( .A1(n3487), .A2(n3486), .ZN(n3488) );
  NOR2_X1 U4286 ( .A1(n3509), .A2(n3488), .ZN(n4325) );
  OAI22_X1 U4287 ( .A1(n4182), .A2(n4486), .B1(n4359), .B2(n4129), .ZN(n3494)
         );
  NAND2_X1 U4288 ( .A1(n3489), .A2(n3490), .ZN(n3491) );
  NAND2_X1 U4289 ( .A1(n3492), .A2(n3491), .ZN(n4251) );
  NOR2_X1 U4290 ( .A1(n4251), .A2(n4186), .ZN(n3493) );
  AOI211_X1 U4291 ( .C1(n4325), .C2(n4548), .A(n3494), .B(n3493), .ZN(n3495)
         );
  OAI21_X1 U4292 ( .B1(n2222), .B2(n4253), .A(n3495), .ZN(U3274) );
  OAI22_X1 U4293 ( .A1(n4513), .A2(n4267), .B1(n3496), .B2(n4265), .ZN(n3498)
         );
  AOI211_X1 U4294 ( .C1(n3499), .C2(n4590), .A(n3498), .B(n3497), .ZN(n3501)
         );
  MUX2_X1 U4295 ( .A(n2798), .B(n3501), .S(n4634), .Z(n3500) );
  OAI21_X1 U4296 ( .B1(n4619), .B2(n3504), .A(n3500), .ZN(U3531) );
  INV_X1 U4297 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3502) );
  MUX2_X1 U4298 ( .A(n3502), .B(n3501), .S(n4613), .Z(n3503) );
  OAI21_X1 U4299 ( .B1(n3504), .B2(n4580), .A(n3503), .ZN(U3493) );
  AND2_X1 U4300 ( .A1(n4137), .A2(n4139), .ZN(n3819) );
  XNOR2_X1 U4301 ( .A(n4138), .B(n3819), .ZN(n3506) );
  NOR2_X1 U4302 ( .A1(n4149), .A2(n4535), .ZN(n3505) );
  AOI21_X1 U4303 ( .B1(n3506), .B2(n4519), .A(n3505), .ZN(n4247) );
  XNOR2_X1 U4304 ( .A(n3507), .B(n3819), .ZN(n4246) );
  INV_X1 U4305 ( .A(n4171), .ZN(n3508) );
  OAI21_X1 U4306 ( .B1(n3509), .B2(n4243), .A(n3508), .ZN(n4321) );
  INV_X1 U4307 ( .A(n3510), .ZN(n3676) );
  AOI22_X1 U4308 ( .A1(n2222), .A2(REG2_REG_17__SCAN_IN), .B1(n3676), .B2(
        n4543), .ZN(n3511) );
  OAI21_X1 U4309 ( .B1(n4244), .B2(n4107), .A(n3511), .ZN(n3512) );
  AOI21_X1 U4310 ( .B1(n3513), .B2(n4111), .A(n3512), .ZN(n3514) );
  OAI21_X1 U4311 ( .B1(n4321), .B2(n4159), .A(n3514), .ZN(n3515) );
  AOI21_X1 U4312 ( .B1(n4246), .B2(n4161), .A(n3515), .ZN(n3516) );
  OAI21_X1 U4313 ( .B1(n4247), .B2(n2222), .A(n3516), .ZN(U3273) );
  NAND2_X1 U4314 ( .A1(n3918), .A2(n2883), .ZN(n3522) );
  NAND2_X1 U4315 ( .A1(n3591), .A2(n3520), .ZN(n3521) );
  NAND2_X1 U4316 ( .A1(n3522), .A2(n3521), .ZN(n3523) );
  XNOR2_X1 U4317 ( .A(n3523), .B(n3607), .ZN(n3528) );
  NOR2_X1 U4318 ( .A1(n2892), .A2(n4257), .ZN(n3524) );
  AOI21_X1 U4319 ( .B1(n2947), .B2(n3918), .A(n3524), .ZN(n4352) );
  OAI22_X1 U4320 ( .A1(n4244), .A2(n2892), .B1(n2899), .B2(n4346), .ZN(n3525)
         );
  XNOR2_X1 U4321 ( .A(n3525), .B(n3607), .ZN(n3527) );
  OAI22_X1 U4322 ( .A1(n4244), .A2(n3606), .B1(n2892), .B2(n4346), .ZN(n3526)
         );
  NOR2_X1 U4323 ( .A1(n3527), .A2(n3526), .ZN(n3530) );
  AOI21_X1 U4324 ( .B1(n3527), .B2(n3526), .A(n3530), .ZN(n4354) );
  OAI211_X1 U4325 ( .C1(n3734), .C2(n4352), .A(n4354), .B(n4351), .ZN(n3532)
         );
  INV_X1 U4326 ( .A(n3530), .ZN(n3531) );
  NAND2_X1 U4327 ( .A1(n3532), .A2(n3531), .ZN(n3668) );
  OAI22_X1 U4328 ( .A1(n4178), .A2(n2892), .B1(n2899), .B2(n4243), .ZN(n3533)
         );
  XNOR2_X1 U4329 ( .A(n3533), .B(n3607), .ZN(n3535) );
  OAI22_X1 U4330 ( .A1(n4178), .A2(n3606), .B1(n2892), .B2(n4243), .ZN(n3534)
         );
  NAND2_X1 U4331 ( .A1(n3535), .A2(n3534), .ZN(n3670) );
  NOR2_X1 U4332 ( .A1(n3535), .A2(n3534), .ZN(n3669) );
  OAI22_X1 U4333 ( .A1(n4149), .A2(n2892), .B1(n2899), .B2(n4170), .ZN(n3536)
         );
  XNOR2_X1 U4334 ( .A(n3536), .B(n3607), .ZN(n3537) );
  OAI22_X1 U4335 ( .A1(n4149), .A2(n3606), .B1(n2892), .B2(n4170), .ZN(n3538)
         );
  AND2_X1 U4336 ( .A1(n3537), .A2(n3538), .ZN(n3711) );
  INV_X1 U4337 ( .A(n3537), .ZN(n3540) );
  INV_X1 U4338 ( .A(n3538), .ZN(n3539) );
  AOI22_X1 U4339 ( .A1(n2947), .A2(n4176), .B1(n2883), .B2(n4154), .ZN(n3544)
         );
  NAND2_X1 U4340 ( .A1(n4176), .A2(n3564), .ZN(n3542) );
  NAND2_X1 U4341 ( .A1(n3591), .A2(n4154), .ZN(n3541) );
  NAND2_X1 U4342 ( .A1(n3542), .A2(n3541), .ZN(n3543) );
  XNOR2_X1 U4343 ( .A(n3543), .B(n3607), .ZN(n3545) );
  XOR2_X1 U4344 ( .A(n3544), .B(n3545), .Z(n3640) );
  NAND2_X1 U4345 ( .A1(n4146), .A2(n2883), .ZN(n3547) );
  NAND2_X1 U4346 ( .A1(n3591), .A2(n3787), .ZN(n3546) );
  NAND2_X1 U4347 ( .A1(n3547), .A2(n3546), .ZN(n3548) );
  XNOR2_X1 U4348 ( .A(n3548), .B(n3607), .ZN(n3551) );
  NAND2_X1 U4349 ( .A1(n2947), .A2(n4146), .ZN(n3550) );
  NAND2_X1 U4350 ( .A1(n2883), .A2(n3787), .ZN(n3549) );
  NAND2_X1 U4351 ( .A1(n3550), .A2(n3549), .ZN(n3552) );
  NAND2_X1 U4352 ( .A1(n3551), .A2(n3552), .ZN(n3693) );
  INV_X1 U4353 ( .A(n3551), .ZN(n3554) );
  INV_X1 U4354 ( .A(n3552), .ZN(n3553) );
  NAND2_X1 U4355 ( .A1(n3554), .A2(n3553), .ZN(n3694) );
  NAND2_X2 U4356 ( .A1(n3690), .A2(n3694), .ZN(n3651) );
  NAND2_X1 U4357 ( .A1(n4086), .A2(n2883), .ZN(n3556) );
  NAND2_X1 U4358 ( .A1(n3591), .A2(n4110), .ZN(n3555) );
  NAND2_X1 U4359 ( .A1(n3556), .A2(n3555), .ZN(n3557) );
  XNOR2_X1 U4360 ( .A(n3557), .B(n3607), .ZN(n3649) );
  NAND2_X1 U4361 ( .A1(n4086), .A2(n2947), .ZN(n3559) );
  NAND2_X1 U4362 ( .A1(n2883), .A2(n4110), .ZN(n3558) );
  NAND2_X1 U4363 ( .A1(n3559), .A2(n3558), .ZN(n3560) );
  NOR2_X1 U4364 ( .A1(n3649), .A2(n3560), .ZN(n3562) );
  INV_X1 U4365 ( .A(n3649), .ZN(n3561) );
  INV_X1 U4366 ( .A(n3560), .ZN(n3648) );
  AOI22_X1 U4367 ( .A1(n4067), .A2(n3564), .B1(n3591), .B2(n4085), .ZN(n3563)
         );
  XNOR2_X1 U4368 ( .A(n3563), .B(n3607), .ZN(n3568) );
  AOI22_X1 U4369 ( .A1(n4067), .A2(n2947), .B1(n2883), .B2(n4085), .ZN(n3569)
         );
  XNOR2_X1 U4370 ( .A(n3568), .B(n3569), .ZN(n3702) );
  OAI22_X1 U4371 ( .A1(n4089), .A2(n2892), .B1(n2899), .B2(n3632), .ZN(n3565)
         );
  XNOR2_X1 U4372 ( .A(n3565), .B(n3607), .ZN(n3573) );
  OR2_X1 U4373 ( .A1(n4089), .A2(n3606), .ZN(n3567) );
  NAND2_X1 U4374 ( .A1(n2883), .A2(n4071), .ZN(n3566) );
  NAND2_X1 U4375 ( .A1(n3567), .A2(n3566), .ZN(n3574) );
  XNOR2_X1 U4376 ( .A(n3573), .B(n3574), .ZN(n3629) );
  INV_X1 U4377 ( .A(n3568), .ZN(n3571) );
  INV_X1 U4378 ( .A(n3569), .ZN(n3570) );
  NOR2_X1 U4379 ( .A1(n3571), .A2(n3570), .ZN(n3630) );
  INV_X1 U4380 ( .A(n3573), .ZN(n3576) );
  INV_X1 U4381 ( .A(n3574), .ZN(n3575) );
  NAND2_X1 U4382 ( .A1(n4029), .A2(n2947), .ZN(n3578) );
  NAND2_X1 U4383 ( .A1(n2883), .A2(n4051), .ZN(n3577) );
  NAND2_X1 U4384 ( .A1(n3578), .A2(n3577), .ZN(n3581) );
  OAI22_X1 U4385 ( .A1(n4070), .A2(n2892), .B1(n2223), .B2(n3579), .ZN(n3580)
         );
  XOR2_X1 U4386 ( .A(n3607), .B(n3580), .Z(n3682) );
  OAI21_X2 U4387 ( .B1(n3679), .B2(n3682), .A(n3680), .ZN(n3658) );
  NAND2_X1 U4388 ( .A1(n3915), .A2(n3564), .ZN(n3585) );
  NAND2_X1 U4389 ( .A1(n3591), .A2(n4032), .ZN(n3584) );
  NAND2_X1 U4390 ( .A1(n3585), .A2(n3584), .ZN(n3586) );
  XNOR2_X1 U4391 ( .A(n3586), .B(n3600), .ZN(n3590) );
  NOR2_X1 U4392 ( .A1(n2892), .A2(n3587), .ZN(n3588) );
  AOI21_X1 U4393 ( .B1(n3915), .B2(n2947), .A(n3588), .ZN(n3589) );
  NAND2_X1 U4394 ( .A1(n3590), .A2(n3589), .ZN(n3659) );
  NOR2_X1 U4395 ( .A1(n3590), .A2(n3589), .ZN(n3660) );
  NAND2_X1 U4396 ( .A1(n3993), .A2(n2883), .ZN(n3593) );
  NAND2_X1 U4397 ( .A1(n3591), .A2(n4010), .ZN(n3592) );
  NAND2_X1 U4398 ( .A1(n3593), .A2(n3592), .ZN(n3594) );
  XNOR2_X1 U4399 ( .A(n3594), .B(n3600), .ZN(n3599) );
  INV_X1 U4400 ( .A(n3599), .ZN(n3597) );
  NOR2_X1 U4401 ( .A1(n2892), .A2(n4014), .ZN(n3595) );
  AOI21_X1 U4402 ( .B1(n3993), .B2(n2947), .A(n3595), .ZN(n3598) );
  INV_X1 U4403 ( .A(n3598), .ZN(n3596) );
  NAND2_X1 U4404 ( .A1(n3597), .A2(n3596), .ZN(n3723) );
  OAI22_X1 U4405 ( .A1(n3729), .A2(n2892), .B1(n4197), .B2(n2899), .ZN(n3601)
         );
  XNOR2_X1 U4406 ( .A(n3601), .B(n3600), .ZN(n3603) );
  OAI22_X1 U4407 ( .A1(n3729), .A2(n3606), .B1(n4197), .B2(n2892), .ZN(n3604)
         );
  XNOR2_X1 U4408 ( .A(n3603), .B(n3604), .ZN(n3623) );
  INV_X1 U4409 ( .A(n3603), .ZN(n3605) );
  OAI22_X1 U4410 ( .A1(n3966), .A2(n3606), .B1(n2892), .B2(n3613), .ZN(n3608)
         );
  XNOR2_X1 U4411 ( .A(n3608), .B(n3607), .ZN(n3610) );
  OAI22_X1 U4412 ( .A1(n3966), .A2(n2892), .B1(n2899), .B2(n3613), .ZN(n3609)
         );
  XNOR2_X1 U4413 ( .A(n3610), .B(n3609), .ZN(n3611) );
  OAI22_X1 U4414 ( .A1(n3729), .A2(n4344), .B1(STATE_REG_SCAN_IN), .B2(n3612), 
        .ZN(n3616) );
  INV_X1 U4415 ( .A(n3914), .ZN(n3614) );
  OAI22_X1 U4416 ( .A1(n3614), .A2(n3728), .B1(n4347), .B2(n3613), .ZN(n3615)
         );
  AOI211_X1 U4417 ( .C1(n3978), .C2(n3743), .A(n3616), .B(n3615), .ZN(n3617)
         );
  OAI21_X1 U4418 ( .B1(n3618), .B2(n3745), .A(n3617), .ZN(U3217) );
  NAND3_X1 U4419 ( .A1(n3620), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3621) );
  INV_X1 U4420 ( .A(DATAI_31_), .ZN(n4879) );
  OAI22_X1 U4421 ( .A1(n3619), .A2(n3621), .B1(STATE_REG_SCAN_IN), .B2(n4879), 
        .ZN(U3321) );
  XNOR2_X1 U4422 ( .A(n3622), .B(n3623), .ZN(n3627) );
  OAI22_X1 U4423 ( .A1(n4198), .A2(n4344), .B1(n4347), .B2(n4197), .ZN(n3625)
         );
  INV_X1 U4424 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4709) );
  OAI22_X1 U4425 ( .A1(n3966), .A2(n3728), .B1(STATE_REG_SCAN_IN), .B2(n4709), 
        .ZN(n3624) );
  AOI211_X1 U4426 ( .C1(n3991), .C2(n3743), .A(n3625), .B(n3624), .ZN(n3626)
         );
  OAI21_X1 U4427 ( .B1(n3627), .B2(n3745), .A(n3626), .ZN(U3211) );
  OAI21_X1 U4428 ( .B1(n2228), .B2(n3630), .A(n3629), .ZN(n3631) );
  NAND3_X1 U4429 ( .A1(n3628), .A2(n4355), .A3(n3631), .ZN(n3638) );
  OAI22_X1 U4430 ( .A1(n4347), .A2(n3632), .B1(n2624), .B2(n4344), .ZN(n3636)
         );
  NAND2_X1 U4431 ( .A1(n4029), .A2(n4350), .ZN(n3633) );
  OAI21_X1 U4432 ( .B1(STATE_REG_SCAN_IN), .B2(n3634), .A(n3633), .ZN(n3635)
         );
  NOR2_X1 U4433 ( .A1(n3636), .A2(n3635), .ZN(n3637) );
  OAI211_X1 U4434 ( .C1(n4360), .C2(n3639), .A(n3638), .B(n3637), .ZN(U3213)
         );
  XOR2_X1 U4435 ( .A(n3640), .B(n2236), .Z(n3647) );
  INV_X1 U4436 ( .A(n3641), .ZN(n4157) );
  AND2_X1 U4437 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3952) );
  AOI21_X1 U4438 ( .B1(n3738), .B2(n3916), .A(n3952), .ZN(n3643) );
  NAND2_X1 U4439 ( .A1(n4350), .A2(n4146), .ZN(n3642) );
  OAI211_X1 U4440 ( .C1(n4347), .C2(n3644), .A(n3643), .B(n3642), .ZN(n3645)
         );
  AOI21_X1 U4441 ( .B1(n3743), .B2(n4157), .A(n3645), .ZN(n3646) );
  OAI21_X1 U4442 ( .B1(n3647), .B2(n3745), .A(n3646), .ZN(U3216) );
  XNOR2_X1 U4443 ( .A(n3649), .B(n3648), .ZN(n3650) );
  XNOR2_X1 U4444 ( .A(n3651), .B(n3650), .ZN(n3652) );
  NAND2_X1 U4445 ( .A1(n3652), .A2(n4355), .ZN(n3657) );
  OAI22_X1 U4446 ( .A1(n4347), .A2(n4224), .B1(n2624), .B2(n3728), .ZN(n3655)
         );
  OAI22_X1 U4447 ( .A1(n4344), .A2(n4225), .B1(STATE_REG_SCAN_IN), .B2(n3653), 
        .ZN(n3654) );
  NOR2_X1 U4448 ( .A1(n3655), .A2(n3654), .ZN(n3656) );
  OAI211_X1 U4449 ( .C1(n4360), .C2(n4105), .A(n3657), .B(n3656), .ZN(U3220)
         );
  NOR2_X1 U4450 ( .A1(n3660), .A2(n2329), .ZN(n3661) );
  XNOR2_X1 U4451 ( .A(n3658), .B(n3661), .ZN(n3667) );
  INV_X1 U4452 ( .A(n4035), .ZN(n3664) );
  AOI22_X1 U4453 ( .A1(n3993), .A2(n4350), .B1(n3725), .B2(n4032), .ZN(n3663)
         );
  AOI22_X1 U4454 ( .A1(n4029), .A2(n3738), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3662) );
  OAI211_X1 U4455 ( .C1(n4360), .C2(n3664), .A(n3663), .B(n3662), .ZN(n3665)
         );
  INV_X1 U4456 ( .A(n3665), .ZN(n3666) );
  OAI21_X1 U4457 ( .B1(n3667), .B2(n3745), .A(n3666), .ZN(U3222) );
  INV_X1 U4458 ( .A(n3669), .ZN(n3671) );
  NAND2_X1 U4459 ( .A1(n3671), .A2(n3670), .ZN(n3672) );
  XNOR2_X1 U4460 ( .A(n3668), .B(n3672), .ZN(n3678) );
  AND2_X1 U4461 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4500) );
  AOI21_X1 U4462 ( .B1(n3738), .B2(n3917), .A(n4500), .ZN(n3674) );
  NAND2_X1 U4463 ( .A1(n4350), .A2(n3916), .ZN(n3673) );
  OAI211_X1 U4464 ( .C1(n4347), .C2(n4243), .A(n3674), .B(n3673), .ZN(n3675)
         );
  AOI21_X1 U4465 ( .B1(n3743), .B2(n3676), .A(n3675), .ZN(n3677) );
  OAI21_X1 U4466 ( .B1(n3678), .B2(n3745), .A(n3677), .ZN(U3225) );
  INV_X1 U4467 ( .A(n3679), .ZN(n3681) );
  NAND2_X1 U4468 ( .A1(n3681), .A2(n3680), .ZN(n3683) );
  XNOR2_X1 U4469 ( .A(n3683), .B(n3682), .ZN(n3689) );
  INV_X1 U4470 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4868) );
  OAI22_X1 U4471 ( .A1(n4089), .A2(n4344), .B1(STATE_REG_SCAN_IN), .B2(n4868), 
        .ZN(n3684) );
  INV_X1 U4472 ( .A(n3684), .ZN(n3686) );
  AOI22_X1 U4473 ( .A1(n3725), .A2(n4051), .B1(n3915), .B2(n4350), .ZN(n3685)
         );
  OAI211_X1 U4474 ( .C1(n4360), .C2(n4054), .A(n3686), .B(n3685), .ZN(n3687)
         );
  INV_X1 U4475 ( .A(n3687), .ZN(n3688) );
  OAI21_X1 U4476 ( .B1(n3689), .B2(n3745), .A(n3688), .ZN(U3226) );
  INV_X1 U4477 ( .A(n3694), .ZN(n3691) );
  NOR2_X1 U4478 ( .A1(n3690), .A2(n3691), .ZN(n3696) );
  AOI21_X1 U4479 ( .B1(n3694), .B2(n3693), .A(n3692), .ZN(n3695) );
  OAI21_X1 U4480 ( .B1(n3696), .B2(n3695), .A(n4355), .ZN(n3700) );
  OAI22_X1 U4481 ( .A1(n4347), .A2(n4128), .B1(n4117), .B2(n3728), .ZN(n3698)
         );
  INV_X1 U4482 ( .A(n4176), .ZN(n3717) );
  INV_X1 U4483 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4867) );
  OAI22_X1 U4484 ( .A1(n4344), .A2(n3717), .B1(STATE_REG_SCAN_IN), .B2(n4867), 
        .ZN(n3697) );
  NOR2_X1 U4485 ( .A1(n3698), .A2(n3697), .ZN(n3699) );
  OAI211_X1 U4486 ( .C1(n4360), .C2(n4130), .A(n3700), .B(n3699), .ZN(U3230)
         );
  AOI21_X1 U4487 ( .B1(n3702), .B2(n3701), .A(n2228), .ZN(n3708) );
  INV_X1 U4488 ( .A(n4092), .ZN(n3706) );
  OAI22_X1 U4489 ( .A1(n4344), .A2(n4117), .B1(STATE_REG_SCAN_IN), .B2(n3703), 
        .ZN(n3705) );
  OAI22_X1 U4490 ( .A1(n4347), .A2(n4091), .B1(n4089), .B2(n3728), .ZN(n3704)
         );
  AOI211_X1 U4491 ( .C1(n3743), .C2(n3706), .A(n3705), .B(n3704), .ZN(n3707)
         );
  OAI21_X1 U4492 ( .B1(n3708), .B2(n3745), .A(n3707), .ZN(U3232) );
  INV_X1 U4493 ( .A(n3709), .ZN(n3714) );
  OAI21_X1 U4494 ( .B1(n3711), .B2(n3713), .A(n3710), .ZN(n3712) );
  OAI21_X1 U4495 ( .B1(n3714), .B2(n3713), .A(n3712), .ZN(n3715) );
  NAND2_X1 U4496 ( .A1(n3715), .A2(n4355), .ZN(n3721) );
  OAI22_X1 U4497 ( .A1(n4347), .A2(n4170), .B1(n4178), .B2(n4344), .ZN(n3719)
         );
  OAI22_X1 U4498 ( .A1(n3728), .A2(n3717), .B1(STATE_REG_SCAN_IN), .B2(n3716), 
        .ZN(n3718) );
  NOR2_X1 U4499 ( .A1(n3719), .A2(n3718), .ZN(n3720) );
  OAI211_X1 U4500 ( .C1(n4360), .C2(n4166), .A(n3721), .B(n3720), .ZN(U3235)
         );
  NAND2_X1 U4501 ( .A1(n2241), .A2(n3723), .ZN(n3724) );
  XNOR2_X1 U4502 ( .A(n3722), .B(n3724), .ZN(n3733) );
  AOI22_X1 U4503 ( .A1(n3915), .A2(n3738), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3727) );
  NAND2_X1 U4504 ( .A1(n3725), .A2(n4010), .ZN(n3726) );
  OAI211_X1 U4505 ( .C1(n3729), .C2(n3728), .A(n3727), .B(n3726), .ZN(n3731)
         );
  NOR2_X1 U4506 ( .A1(n4360), .A2(n4017), .ZN(n3730) );
  NOR2_X1 U4507 ( .A1(n3731), .A2(n3730), .ZN(n3732) );
  OAI21_X1 U4508 ( .B1(n3733), .B2(n3745), .A(n3732), .ZN(U3237) );
  INV_X1 U4509 ( .A(n3734), .ZN(n3735) );
  NAND2_X1 U4510 ( .A1(n3735), .A2(n4351), .ZN(n3736) );
  XNOR2_X1 U4511 ( .A(n3736), .B(n4352), .ZN(n3746) );
  INV_X1 U4512 ( .A(n3737), .ZN(n3742) );
  AND2_X1 U4513 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4480) );
  AOI21_X1 U4514 ( .B1(n4350), .B2(n3917), .A(n4480), .ZN(n3740) );
  NAND2_X1 U4515 ( .A1(n3738), .A2(n3919), .ZN(n3739) );
  OAI211_X1 U4516 ( .C1(n4347), .C2(n4257), .A(n3740), .B(n3739), .ZN(n3741)
         );
  AOI21_X1 U4517 ( .B1(n3743), .B2(n3742), .A(n3741), .ZN(n3744) );
  OAI21_X1 U4518 ( .B1(n3746), .B2(n3745), .A(n3744), .ZN(U3238) );
  NAND2_X1 U4519 ( .A1(n3868), .A2(n3866), .ZN(n3749) );
  NAND2_X1 U4520 ( .A1(n3748), .A2(n3747), .ZN(n3853) );
  NAND2_X1 U4521 ( .A1(n3853), .A2(n3866), .ZN(n3856) );
  OAI21_X1 U4522 ( .B1(n3750), .B2(n3749), .A(n3856), .ZN(n3753) );
  INV_X1 U4523 ( .A(n3751), .ZN(n3876) );
  AOI211_X1 U4524 ( .C1(n3753), .C2(n3877), .A(n3752), .B(n3876), .ZN(n3754)
         );
  OAI21_X1 U4525 ( .B1(n3754), .B2(n3881), .A(n3880), .ZN(n3755) );
  NAND2_X1 U4526 ( .A1(n3755), .A2(n3885), .ZN(n3757) );
  INV_X1 U4527 ( .A(n3756), .ZN(n3888) );
  AOI21_X1 U4528 ( .B1(n3758), .B2(n3757), .A(n3888), .ZN(n3760) );
  INV_X1 U4529 ( .A(n3886), .ZN(n3759) );
  OAI21_X1 U4530 ( .B1(n3760), .B2(n3759), .A(n3889), .ZN(n3761) );
  AND3_X1 U4531 ( .A1(n3761), .A2(n3990), .A3(n3893), .ZN(n3766) );
  NAND2_X1 U4532 ( .A1(n3763), .A2(n3762), .ZN(n3895) );
  INV_X1 U4533 ( .A(n3764), .ZN(n3765) );
  AOI21_X1 U4534 ( .B1(n3914), .B2(n3774), .A(n3765), .ZN(n3896) );
  OAI21_X1 U4535 ( .B1(n3766), .B2(n3895), .A(n3896), .ZN(n3779) );
  NAND2_X1 U4536 ( .A1(n3772), .A2(DATAI_30_), .ZN(n3776) );
  INV_X1 U4537 ( .A(n3776), .ZN(n4193) );
  NAND2_X1 U4538 ( .A1(n3767), .A2(REG1_REG_31__SCAN_IN), .ZN(n3771) );
  NAND2_X1 U4539 ( .A1(n3768), .A2(REG2_REG_31__SCAN_IN), .ZN(n3770) );
  NAND2_X1 U4540 ( .A1(n2672), .A2(REG0_REG_31__SCAN_IN), .ZN(n3769) );
  NAND3_X1 U4541 ( .A1(n3771), .A2(n3770), .A3(n3769), .ZN(n3960) );
  INV_X1 U4542 ( .A(n3960), .ZN(n3775) );
  INV_X1 U4543 ( .A(n3913), .ZN(n3773) );
  NAND2_X1 U4544 ( .A1(n3772), .A2(DATAI_31_), .ZN(n3961) );
  AND2_X1 U4545 ( .A1(n3960), .A2(n3961), .ZN(n3898) );
  AOI21_X1 U4546 ( .B1(n4193), .B2(n3773), .A(n3898), .ZN(n3807) );
  OAI21_X1 U4547 ( .B1(n3914), .B2(n3774), .A(n3807), .ZN(n3894) );
  AOI21_X1 U4548 ( .B1(n4193), .B2(n3775), .A(n3894), .ZN(n3778) );
  NAND2_X1 U4549 ( .A1(n3913), .A2(n3776), .ZN(n3806) );
  AOI21_X1 U4550 ( .B1(n3806), .B2(n3960), .A(n3961), .ZN(n3777) );
  AOI21_X1 U4551 ( .B1(n3779), .B2(n3778), .A(n3777), .ZN(n3825) );
  INV_X1 U4552 ( .A(n4081), .ZN(n4082) );
  OR2_X1 U4553 ( .A1(n3780), .A2(n4062), .ZN(n4100) );
  NOR4_X1 U4554 ( .A1(n4082), .A2(n3782), .A3(n3781), .A4(n4100), .ZN(n3790)
         );
  NOR4_X1 U4555 ( .A1(n2561), .A2(n4514), .A3(n3784), .A4(n3783), .ZN(n3789)
         );
  NOR4_X1 U4556 ( .A1(n2690), .A2(n2688), .A3(n3786), .A4(n3785), .ZN(n3788)
         );
  XNOR2_X1 U4557 ( .A(n4146), .B(n3787), .ZN(n4121) );
  NAND4_X1 U4558 ( .A1(n3790), .A2(n3789), .A3(n3788), .A4(n4121), .ZN(n3823)
         );
  INV_X1 U4559 ( .A(n3791), .ZN(n3792) );
  OR2_X1 U4560 ( .A1(n3793), .A2(n3792), .ZN(n4064) );
  NAND4_X1 U4561 ( .A1(n3797), .A2(n3796), .A3(n3795), .A4(n3794), .ZN(n3812)
         );
  NOR2_X1 U4562 ( .A1(n3799), .A2(n3798), .ZN(n4007) );
  INV_X1 U4563 ( .A(n3800), .ZN(n3801) );
  OR2_X1 U4564 ( .A1(n4004), .A2(n3801), .ZN(n4026) );
  INV_X1 U4565 ( .A(n4026), .ZN(n3804) );
  INV_X1 U4566 ( .A(n4024), .ZN(n3803) );
  NOR2_X1 U4567 ( .A1(n3803), .A2(n3802), .ZN(n4044) );
  NAND4_X1 U4568 ( .A1(n3990), .A2(n4007), .A3(n3804), .A4(n4044), .ZN(n3811)
         );
  OR2_X1 U4569 ( .A1(n3960), .A2(n3961), .ZN(n3805) );
  AND2_X1 U4570 ( .A1(n3806), .A2(n3805), .ZN(n3897) );
  NAND4_X1 U4571 ( .A1(n3809), .A2(n3808), .A3(n3897), .A4(n3807), .ZN(n3810)
         );
  NOR3_X1 U4572 ( .A1(n3812), .A2(n3811), .A3(n3810), .ZN(n3816) );
  INV_X1 U4573 ( .A(n3813), .ZN(n3815) );
  OR2_X1 U4574 ( .A1(n3815), .A2(n3814), .ZN(n4144) );
  NAND3_X1 U4575 ( .A1(n4064), .A2(n3816), .A3(n4144), .ZN(n3821) );
  NAND4_X1 U4576 ( .A1(n3819), .A2(n3818), .A3(n4172), .A4(n3817), .ZN(n3820)
         );
  NOR4_X1 U4577 ( .A1(n3823), .A2(n3822), .A3(n3821), .A4(n3820), .ZN(n3824)
         );
  MUX2_X1 U4578 ( .A(n3825), .B(n3824), .S(n2721), .Z(n3905) );
  OAI211_X1 U4579 ( .C1(n3828), .C2(n2711), .A(n3827), .B(n3826), .ZN(n3829)
         );
  NAND3_X1 U4580 ( .A1(n3829), .A2(n2692), .A3(n2689), .ZN(n3831) );
  OAI211_X1 U4581 ( .C1(n3833), .C2(n3832), .A(n3831), .B(n3830), .ZN(n3836)
         );
  NAND3_X1 U4582 ( .A1(n3836), .A2(n3835), .A3(n3834), .ZN(n3839) );
  NAND4_X1 U4583 ( .A1(n3839), .A2(n3838), .A3(n3837), .A4(n3848), .ZN(n3842)
         );
  NAND3_X1 U4584 ( .A1(n3842), .A2(n3841), .A3(n3840), .ZN(n3843) );
  NAND3_X1 U4585 ( .A1(n3843), .A2(n3850), .A3(n3849), .ZN(n3846) );
  AND3_X1 U4586 ( .A1(n3846), .A2(n3845), .A3(n3844), .ZN(n3854) );
  INV_X1 U4587 ( .A(n3856), .ZN(n3871) );
  INV_X1 U4588 ( .A(n3847), .ZN(n3851) );
  NAND4_X1 U4589 ( .A1(n3851), .A2(n3850), .A3(n3849), .A4(n3848), .ZN(n3852)
         );
  OAI22_X1 U4590 ( .A1(n3854), .A2(n3853), .B1(n3871), .B2(n3852), .ZN(n3859)
         );
  INV_X1 U4591 ( .A(n3855), .ZN(n3857) );
  AOI22_X1 U4592 ( .A1(n3859), .A2(n3858), .B1(n3857), .B2(n3856), .ZN(n3873)
         );
  NAND3_X1 U4593 ( .A1(n3863), .A2(n3861), .A3(n3860), .ZN(n3872) );
  INV_X1 U4594 ( .A(n3862), .ZN(n3865) );
  OAI21_X1 U4595 ( .B1(n3865), .B2(n3864), .A(n3863), .ZN(n3869) );
  AND4_X1 U4596 ( .A1(n3869), .A2(n3868), .A3(n3867), .A4(n3866), .ZN(n3870)
         );
  OAI22_X1 U4597 ( .A1(n3873), .A2(n3872), .B1(n3871), .B2(n3870), .ZN(n3875)
         );
  NAND2_X1 U4598 ( .A1(n3875), .A2(n3874), .ZN(n3878) );
  AOI21_X1 U4599 ( .B1(n3878), .B2(n3877), .A(n3876), .ZN(n3882) );
  OAI211_X1 U4600 ( .C1(n3882), .C2(n3881), .A(n3880), .B(n3879), .ZN(n3884)
         );
  AOI21_X1 U4601 ( .B1(n3885), .B2(n3884), .A(n3883), .ZN(n3887) );
  OAI21_X1 U4602 ( .B1(n3888), .B2(n3887), .A(n3886), .ZN(n3890) );
  NAND2_X1 U4603 ( .A1(n3890), .A2(n3889), .ZN(n3891) );
  NAND4_X1 U4604 ( .A1(n3896), .A2(n3893), .A3(n3892), .A4(n3891), .ZN(n3902)
         );
  AOI21_X1 U4605 ( .B1(n3896), .B2(n3895), .A(n3894), .ZN(n3901) );
  INV_X1 U4606 ( .A(n3897), .ZN(n3900) );
  INV_X1 U4607 ( .A(n3898), .ZN(n3899) );
  AOI22_X1 U4608 ( .A1(n3902), .A2(n3901), .B1(n3900), .B2(n3899), .ZN(n3904)
         );
  MUX2_X1 U4609 ( .A(n3905), .B(n3904), .S(n3903), .Z(n3906) );
  XNOR2_X1 U4610 ( .A(n3906), .B(n4181), .ZN(n3912) );
  NAND2_X1 U4611 ( .A1(n3908), .A2(n3907), .ZN(n3909) );
  OAI211_X1 U4612 ( .C1(n4337), .C2(n3911), .A(n3909), .B(B_REG_SCAN_IN), .ZN(
        n3910) );
  OAI21_X1 U4613 ( .B1(n3912), .B2(n3911), .A(n3910), .ZN(U3239) );
  MUX2_X1 U4614 ( .A(DATAO_REG_31__SCAN_IN), .B(n3960), .S(n3928), .Z(U3581)
         );
  MUX2_X1 U4615 ( .A(DATAO_REG_30__SCAN_IN), .B(n3913), .S(n3928), .Z(U3580)
         );
  MUX2_X1 U4616 ( .A(DATAO_REG_29__SCAN_IN), .B(n3914), .S(n3928), .Z(U3579)
         );
  MUX2_X1 U4617 ( .A(DATAO_REG_28__SCAN_IN), .B(n3987), .S(n3928), .Z(U3578)
         );
  MUX2_X1 U4618 ( .A(DATAO_REG_27__SCAN_IN), .B(n4011), .S(n3928), .Z(U3577)
         );
  MUX2_X1 U4619 ( .A(DATAO_REG_26__SCAN_IN), .B(n3993), .S(n3928), .Z(U3576)
         );
  MUX2_X1 U4620 ( .A(DATAO_REG_25__SCAN_IN), .B(n3915), .S(n3928), .Z(U3575)
         );
  MUX2_X1 U4621 ( .A(DATAO_REG_24__SCAN_IN), .B(n4029), .S(n3928), .Z(U3574)
         );
  MUX2_X1 U4622 ( .A(DATAO_REG_23__SCAN_IN), .B(n4047), .S(n3928), .Z(U3573)
         );
  MUX2_X1 U4623 ( .A(DATAO_REG_22__SCAN_IN), .B(n4067), .S(n3928), .Z(U3572)
         );
  MUX2_X1 U4624 ( .A(DATAO_REG_21__SCAN_IN), .B(n4086), .S(n3928), .Z(U3571)
         );
  MUX2_X1 U4625 ( .A(DATAO_REG_20__SCAN_IN), .B(n4146), .S(n3928), .Z(U3570)
         );
  MUX2_X1 U4626 ( .A(DATAO_REG_19__SCAN_IN), .B(n4176), .S(n3928), .Z(U3569)
         );
  MUX2_X1 U4627 ( .A(DATAO_REG_18__SCAN_IN), .B(n3916), .S(n3928), .Z(U3568)
         );
  MUX2_X1 U4628 ( .A(DATAO_REG_17__SCAN_IN), .B(n4349), .S(n3928), .Z(U3567)
         );
  MUX2_X1 U4629 ( .A(DATAO_REG_16__SCAN_IN), .B(n3917), .S(n3928), .Z(U3566)
         );
  MUX2_X1 U4630 ( .A(DATAO_REG_15__SCAN_IN), .B(n3918), .S(n3928), .Z(U3565)
         );
  MUX2_X1 U4631 ( .A(DATAO_REG_14__SCAN_IN), .B(n3919), .S(n3928), .Z(U3564)
         );
  MUX2_X1 U4632 ( .A(DATAO_REG_13__SCAN_IN), .B(n3920), .S(n3928), .Z(U3563)
         );
  MUX2_X1 U4633 ( .A(DATAO_REG_12__SCAN_IN), .B(n3921), .S(n3928), .Z(U3562)
         );
  MUX2_X1 U4634 ( .A(DATAO_REG_11__SCAN_IN), .B(n3922), .S(n3928), .Z(U3561)
         );
  MUX2_X1 U4635 ( .A(DATAO_REG_10__SCAN_IN), .B(n4511), .S(n3928), .Z(U3560)
         );
  MUX2_X1 U4636 ( .A(DATAO_REG_9__SCAN_IN), .B(n3923), .S(n3928), .Z(U3559) );
  MUX2_X1 U4637 ( .A(DATAO_REG_8__SCAN_IN), .B(n3924), .S(n3928), .Z(U3558) );
  MUX2_X1 U4638 ( .A(DATAO_REG_7__SCAN_IN), .B(n3126), .S(n3928), .Z(U3557) );
  MUX2_X1 U4639 ( .A(DATAO_REG_6__SCAN_IN), .B(n3925), .S(n3928), .Z(U3556) );
  MUX2_X1 U4640 ( .A(DATAO_REG_5__SCAN_IN), .B(n3926), .S(U4043), .Z(U3555) );
  MUX2_X1 U4641 ( .A(DATAO_REG_4__SCAN_IN), .B(n3927), .S(U4043), .Z(U3554) );
  MUX2_X1 U4642 ( .A(DATAO_REG_3__SCAN_IN), .B(n2874), .S(U4043), .Z(U3553) );
  MUX2_X1 U4643 ( .A(DATAO_REG_2__SCAN_IN), .B(n2409), .S(U4043), .Z(U3552) );
  MUX2_X1 U4644 ( .A(DATAO_REG_1__SCAN_IN), .B(n2401), .S(U4043), .Z(U3551) );
  MUX2_X1 U4645 ( .A(DATAO_REG_0__SCAN_IN), .B(n4533), .S(n3928), .Z(U3550) );
  NAND2_X1 U4646 ( .A1(n3930), .A2(n3929), .ZN(n3940) );
  OAI211_X1 U4647 ( .C1(n3933), .C2(n3932), .A(n4502), .B(n3931), .ZN(n3939)
         );
  OAI211_X1 U4648 ( .C1(n3936), .C2(n3935), .A(n4456), .B(n3934), .ZN(n3938)
         );
  AOI22_X1 U4649 ( .A1(n4501), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3937) );
  NAND4_X1 U4650 ( .A1(n3940), .A2(n3939), .A3(n3938), .A4(n3937), .ZN(U3241)
         );
  INV_X1 U4651 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3941) );
  MUX2_X1 U4652 ( .A(n3941), .B(REG2_REG_19__SCAN_IN), .S(n3954), .Z(n3946) );
  NOR2_X1 U4653 ( .A1(n3944), .A2(n3943), .ZN(n3945) );
  XOR2_X1 U4654 ( .A(n3946), .B(n3945), .Z(n3958) );
  OAI21_X1 U4655 ( .B1(n4556), .B2(n3948), .A(n3947), .ZN(n3951) );
  INV_X1 U4656 ( .A(REG1_REG_19__SCAN_IN), .ZN(n3949) );
  MUX2_X1 U4657 ( .A(REG1_REG_19__SCAN_IN), .B(n3949), .S(n3954), .Z(n3950) );
  XNOR2_X1 U4658 ( .A(n3951), .B(n3950), .ZN(n3956) );
  AOI21_X1 U4659 ( .B1(n4501), .B2(ADDR_REG_19__SCAN_IN), .A(n3952), .ZN(n3953) );
  OAI21_X1 U4660 ( .B1(n4508), .B2(n3954), .A(n3953), .ZN(n3955) );
  AOI21_X1 U4661 ( .B1(n3956), .B2(n4502), .A(n3955), .ZN(n3957) );
  OAI21_X1 U4662 ( .B1(n3958), .B2(n4495), .A(n3957), .ZN(U3259) );
  XNOR2_X1 U4663 ( .A(n4189), .B(n3961), .ZN(n4277) );
  NAND2_X1 U4664 ( .A1(n3960), .A2(n3959), .ZN(n4191) );
  OAI21_X1 U4665 ( .B1(n3961), .B2(n4265), .A(n4191), .ZN(n4274) );
  NAND2_X1 U4666 ( .A1(n4182), .A2(n4274), .ZN(n3963) );
  NAND2_X1 U4667 ( .A1(n2222), .A2(REG2_REG_31__SCAN_IN), .ZN(n3962) );
  OAI211_X1 U4668 ( .C1(n4277), .C2(n4159), .A(n3963), .B(n3962), .ZN(U3260)
         );
  INV_X1 U4669 ( .A(n3964), .ZN(n3976) );
  INV_X1 U4670 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3965) );
  OAI22_X1 U4671 ( .A1(n3966), .A2(n4107), .B1(n4182), .B2(n3965), .ZN(n3967)
         );
  AOI21_X1 U4672 ( .B1(n3968), .B2(n4111), .A(n3967), .ZN(n3975) );
  INV_X1 U4673 ( .A(n3969), .ZN(n3973) );
  OAI22_X1 U4674 ( .A1(n3971), .A2(n4159), .B1(n3970), .B2(n4129), .ZN(n3972)
         );
  OAI21_X1 U4675 ( .B1(n3973), .B2(n3972), .A(n4182), .ZN(n3974) );
  OAI211_X1 U4676 ( .C1(n3976), .C2(n4186), .A(n3975), .B(n3974), .ZN(U3354)
         );
  INV_X1 U4677 ( .A(n3977), .ZN(n3982) );
  AOI22_X1 U4678 ( .A1(n3978), .A2(n4543), .B1(REG2_REG_28__SCAN_IN), .B2(
        n2222), .ZN(n3979) );
  OAI21_X1 U4679 ( .B1(n3980), .B2(n4159), .A(n3979), .ZN(n3981) );
  AOI21_X1 U4680 ( .B1(n3982), .B2(n4182), .A(n3981), .ZN(n3983) );
  OAI21_X1 U4681 ( .B1(n3984), .B2(n4186), .A(n3983), .ZN(U3262) );
  OAI21_X1 U4682 ( .B1(n3986), .B2(n3990), .A(n3985), .ZN(n3988) );
  AOI22_X1 U4683 ( .A1(n3988), .A2(n4519), .B1(n4175), .B2(n3987), .ZN(n4196)
         );
  XOR2_X1 U4684 ( .A(n3990), .B(n3989), .Z(n4201) );
  NAND2_X1 U4685 ( .A1(n4201), .A2(n4161), .ZN(n4002) );
  AOI22_X1 U4686 ( .A1(n3991), .A2(n4543), .B1(n2222), .B2(
        REG2_REG_27__SCAN_IN), .ZN(n3995) );
  NAND2_X1 U4687 ( .A1(n3993), .A2(n3992), .ZN(n3994) );
  NAND2_X1 U4688 ( .A1(n3995), .A2(n3994), .ZN(n3999) );
  INV_X1 U4689 ( .A(n3996), .ZN(n3997) );
  OAI21_X1 U4690 ( .B1(n4016), .B2(n4197), .A(n3997), .ZN(n4284) );
  NOR2_X1 U4691 ( .A1(n4284), .A2(n4159), .ZN(n3998) );
  AOI211_X1 U4692 ( .C1(n4111), .C2(n4000), .A(n3999), .B(n3998), .ZN(n4001)
         );
  OAI211_X1 U4693 ( .C1(n4196), .C2(n2222), .A(n4002), .B(n4001), .ZN(U3263)
         );
  XOR2_X1 U4694 ( .A(n4007), .B(n4003), .Z(n4205) );
  INV_X1 U4695 ( .A(n4205), .ZN(n4022) );
  INV_X1 U4696 ( .A(n4004), .ZN(n4005) );
  NAND2_X1 U4697 ( .A1(n4006), .A2(n4005), .ZN(n4008) );
  XNOR2_X1 U4698 ( .A(n4008), .B(n4007), .ZN(n4009) );
  NAND2_X1 U4699 ( .A1(n4009), .A2(n4519), .ZN(n4013) );
  AOI22_X1 U4700 ( .A1(n4011), .A2(n4175), .B1(n4530), .B2(n4010), .ZN(n4012)
         );
  OAI211_X1 U4701 ( .C1(n4050), .C2(n4267), .A(n4013), .B(n4012), .ZN(n4204)
         );
  NOR2_X1 U4702 ( .A1(n4033), .A2(n4014), .ZN(n4015) );
  OR2_X1 U4703 ( .A1(n4016), .A2(n4015), .ZN(n4288) );
  INV_X1 U4704 ( .A(n4017), .ZN(n4018) );
  AOI22_X1 U4705 ( .A1(REG2_REG_26__SCAN_IN), .A2(n2222), .B1(n4018), .B2(
        n4543), .ZN(n4019) );
  OAI21_X1 U4706 ( .B1(n4288), .B2(n4159), .A(n4019), .ZN(n4020) );
  AOI21_X1 U4707 ( .B1(n4204), .B2(n4182), .A(n4020), .ZN(n4021) );
  OAI21_X1 U4708 ( .B1(n4022), .B2(n4186), .A(n4021), .ZN(U3264) );
  XNOR2_X1 U4709 ( .A(n4023), .B(n4026), .ZN(n4209) );
  INV_X1 U4710 ( .A(n4209), .ZN(n4039) );
  NAND2_X1 U4711 ( .A1(n4025), .A2(n4024), .ZN(n4027) );
  XNOR2_X1 U4712 ( .A(n4027), .B(n4026), .ZN(n4028) );
  NAND2_X1 U4713 ( .A1(n4028), .A2(n4519), .ZN(n4031) );
  AOI22_X1 U4714 ( .A1(n4029), .A2(n4532), .B1(n4032), .B2(n4530), .ZN(n4030)
         );
  OAI211_X1 U4715 ( .C1(n4198), .C2(n4535), .A(n4031), .B(n4030), .ZN(n4208)
         );
  AND2_X1 U4716 ( .A1(n4053), .A2(n4032), .ZN(n4034) );
  OR2_X1 U4717 ( .A1(n4034), .A2(n4033), .ZN(n4292) );
  AOI22_X1 U4718 ( .A1(n2222), .A2(REG2_REG_25__SCAN_IN), .B1(n4035), .B2(
        n4543), .ZN(n4036) );
  OAI21_X1 U4719 ( .B1(n4292), .B2(n4159), .A(n4036), .ZN(n4037) );
  AOI21_X1 U4720 ( .B1(n4208), .B2(n4182), .A(n4037), .ZN(n4038) );
  OAI21_X1 U4721 ( .B1(n4039), .B2(n4186), .A(n4038), .ZN(U3265) );
  XNOR2_X1 U4722 ( .A(n4040), .B(n4044), .ZN(n4213) );
  INV_X1 U4723 ( .A(n4213), .ZN(n4059) );
  INV_X1 U4724 ( .A(n4041), .ZN(n4042) );
  NAND2_X1 U4725 ( .A1(n4043), .A2(n4042), .ZN(n4045) );
  XNOR2_X1 U4726 ( .A(n4045), .B(n4044), .ZN(n4046) );
  NAND2_X1 U4727 ( .A1(n4046), .A2(n4519), .ZN(n4049) );
  AOI22_X1 U4728 ( .A1(n4047), .A2(n4532), .B1(n4530), .B2(n4051), .ZN(n4048)
         );
  OAI211_X1 U4729 ( .C1(n4050), .C2(n4535), .A(n4049), .B(n4048), .ZN(n4212)
         );
  NAND2_X1 U4730 ( .A1(n4073), .A2(n4051), .ZN(n4052) );
  NAND2_X1 U4731 ( .A1(n4053), .A2(n4052), .ZN(n4296) );
  INV_X1 U4732 ( .A(n4054), .ZN(n4055) );
  AOI22_X1 U4733 ( .A1(n2222), .A2(REG2_REG_24__SCAN_IN), .B1(n4055), .B2(
        n4543), .ZN(n4056) );
  OAI21_X1 U4734 ( .B1(n4296), .B2(n4159), .A(n4056), .ZN(n4057) );
  AOI21_X1 U4735 ( .B1(n4212), .B2(n4182), .A(n4057), .ZN(n4058) );
  OAI21_X1 U4736 ( .B1(n4059), .B2(n4186), .A(n4058), .ZN(U3266) );
  XOR2_X1 U4737 ( .A(n4064), .B(n4060), .Z(n4217) );
  INV_X1 U4738 ( .A(n4217), .ZN(n4078) );
  INV_X1 U4739 ( .A(n4061), .ZN(n4101) );
  NOR2_X1 U4740 ( .A1(n4101), .A2(n4100), .ZN(n4099) );
  NOR2_X1 U4741 ( .A1(n4099), .A2(n4062), .ZN(n4083) );
  OAI21_X1 U4742 ( .B1(n4083), .B2(n4082), .A(n4063), .ZN(n4065) );
  XNOR2_X1 U4743 ( .A(n4065), .B(n4064), .ZN(n4066) );
  NAND2_X1 U4744 ( .A1(n4066), .A2(n4519), .ZN(n4069) );
  AOI22_X1 U4745 ( .A1(n4067), .A2(n4532), .B1(n4530), .B2(n4071), .ZN(n4068)
         );
  OAI211_X1 U4746 ( .C1(n4070), .C2(n4535), .A(n4069), .B(n4068), .ZN(n4216)
         );
  NAND2_X1 U4747 ( .A1(n4090), .A2(n4071), .ZN(n4072) );
  NAND2_X1 U4748 ( .A1(n4073), .A2(n4072), .ZN(n4300) );
  AOI22_X1 U4749 ( .A1(n2222), .A2(REG2_REG_23__SCAN_IN), .B1(n4074), .B2(
        n4543), .ZN(n4075) );
  OAI21_X1 U4750 ( .B1(n4300), .B2(n4159), .A(n4075), .ZN(n4076) );
  AOI21_X1 U4751 ( .B1(n4216), .B2(n4182), .A(n4076), .ZN(n4077) );
  OAI21_X1 U4752 ( .B1(n4078), .B2(n4186), .A(n4077), .ZN(U3267) );
  AOI21_X1 U4753 ( .B1(n4081), .B2(n4079), .A(n4080), .ZN(n4221) );
  INV_X1 U4754 ( .A(n4221), .ZN(n4097) );
  XNOR2_X1 U4755 ( .A(n4083), .B(n4082), .ZN(n4084) );
  NAND2_X1 U4756 ( .A1(n4084), .A2(n4519), .ZN(n4088) );
  AOI22_X1 U4757 ( .A1(n4086), .A2(n4532), .B1(n4085), .B2(n4530), .ZN(n4087)
         );
  OAI211_X1 U4758 ( .C1(n4089), .C2(n4535), .A(n4088), .B(n4087), .ZN(n4220)
         );
  OAI21_X1 U4759 ( .B1(n4103), .B2(n4091), .A(n4090), .ZN(n4304) );
  NOR2_X1 U4760 ( .A1(n4304), .A2(n4159), .ZN(n4095) );
  INV_X1 U4761 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4093) );
  OAI22_X1 U4762 ( .A1(n4182), .A2(n4093), .B1(n4092), .B2(n4129), .ZN(n4094)
         );
  AOI211_X1 U4763 ( .C1(n4220), .C2(n4182), .A(n4095), .B(n4094), .ZN(n4096)
         );
  OAI21_X1 U4764 ( .B1(n4097), .B2(n4186), .A(n4096), .ZN(U3268) );
  XNOR2_X1 U4765 ( .A(n4098), .B(n4100), .ZN(n4228) );
  INV_X1 U4766 ( .A(n4228), .ZN(n4115) );
  AOI21_X1 U4767 ( .B1(n4101), .B2(n4100), .A(n4099), .ZN(n4102) );
  OAI22_X1 U4768 ( .A1(n4102), .A2(n4537), .B1(n2624), .B2(n4535), .ZN(n4226)
         );
  INV_X1 U4769 ( .A(n4103), .ZN(n4104) );
  OAI21_X1 U4770 ( .B1(n4126), .B2(n4224), .A(n4104), .ZN(n4308) );
  OAI22_X1 U4771 ( .A1(n4182), .A2(n4106), .B1(n4105), .B2(n4129), .ZN(n4109)
         );
  NOR2_X1 U4772 ( .A1(n4107), .A2(n4225), .ZN(n4108) );
  AOI211_X1 U4773 ( .C1(n4111), .C2(n4110), .A(n4109), .B(n4108), .ZN(n4112)
         );
  OAI21_X1 U4774 ( .B1(n4308), .B2(n4159), .A(n4112), .ZN(n4113) );
  AOI21_X1 U4775 ( .B1(n4226), .B2(n4182), .A(n4113), .ZN(n4114) );
  OAI21_X1 U4776 ( .B1(n4115), .B2(n4186), .A(n4114), .ZN(U3269) );
  XOR2_X1 U4777 ( .A(n4121), .B(n4116), .Z(n4231) );
  OAI22_X1 U4778 ( .A1(n4117), .A2(n4535), .B1(n4265), .B2(n4128), .ZN(n4118)
         );
  AOI21_X1 U4779 ( .B1(n4532), .B2(n4176), .A(n4118), .ZN(n4125) );
  NAND2_X1 U4780 ( .A1(n4120), .A2(n4119), .ZN(n4122) );
  XNOR2_X1 U4781 ( .A(n4122), .B(n4121), .ZN(n4123) );
  NAND2_X1 U4782 ( .A1(n4123), .A2(n4519), .ZN(n4124) );
  OAI211_X1 U4783 ( .C1(n4231), .C2(n4516), .A(n4125), .B(n4124), .ZN(n4232)
         );
  NAND2_X1 U4784 ( .A1(n4232), .A2(n4182), .ZN(n4135) );
  INV_X1 U4785 ( .A(n4126), .ZN(n4127) );
  OAI21_X1 U4786 ( .B1(n2278), .B2(n4128), .A(n4127), .ZN(n4312) );
  INV_X1 U4787 ( .A(n4312), .ZN(n4133) );
  INV_X1 U4788 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4131) );
  OAI22_X1 U4789 ( .A1(n4182), .A2(n4131), .B1(n4130), .B2(n4129), .ZN(n4132)
         );
  AOI21_X1 U4790 ( .B1(n4133), .B2(n4548), .A(n4132), .ZN(n4134) );
  OAI211_X1 U4791 ( .C1(n4231), .C2(n4136), .A(n4135), .B(n4134), .ZN(U3270)
         );
  NAND2_X1 U4792 ( .A1(n4138), .A2(n4137), .ZN(n4140) );
  NAND2_X1 U4793 ( .A1(n4140), .A2(n4139), .ZN(n4173) );
  INV_X1 U4794 ( .A(n4141), .ZN(n4143) );
  OAI21_X1 U4795 ( .B1(n4173), .B2(n4143), .A(n4142), .ZN(n4145) );
  INV_X1 U4796 ( .A(n4144), .ZN(n4152) );
  XNOR2_X1 U4797 ( .A(n4145), .B(n4152), .ZN(n4151) );
  NAND2_X1 U4798 ( .A1(n4154), .A2(n4530), .ZN(n4148) );
  NAND2_X1 U4799 ( .A1(n4146), .A2(n4175), .ZN(n4147) );
  OAI211_X1 U4800 ( .C1(n4149), .C2(n4267), .A(n4148), .B(n4147), .ZN(n4150)
         );
  AOI21_X1 U4801 ( .B1(n4151), .B2(n4519), .A(n4150), .ZN(n4238) );
  XNOR2_X1 U4802 ( .A(n4153), .B(n4152), .ZN(n4236) );
  NAND2_X1 U4803 ( .A1(n4168), .A2(n4154), .ZN(n4155) );
  NAND2_X1 U4804 ( .A1(n4156), .A2(n4155), .ZN(n4316) );
  AOI22_X1 U4805 ( .A1(n2222), .A2(REG2_REG_19__SCAN_IN), .B1(n4157), .B2(
        n4543), .ZN(n4158) );
  OAI21_X1 U4806 ( .B1(n4316), .B2(n4159), .A(n4158), .ZN(n4160) );
  AOI21_X1 U4807 ( .B1(n4236), .B2(n4161), .A(n4160), .ZN(n4162) );
  OAI21_X1 U4808 ( .B1(n4238), .B2(n2222), .A(n4162), .ZN(U3271) );
  INV_X1 U4809 ( .A(n4164), .ZN(n4165) );
  AOI21_X1 U4810 ( .B1(n4172), .B2(n4163), .A(n4165), .ZN(n4242) );
  INV_X1 U4811 ( .A(n4166), .ZN(n4167) );
  AOI22_X1 U4812 ( .A1(n2222), .A2(REG2_REG_18__SCAN_IN), .B1(n4167), .B2(
        n4543), .ZN(n4185) );
  OAI211_X1 U4813 ( .C1(n4171), .C2(n4170), .A(n4169), .B(n4168), .ZN(n4240)
         );
  XNOR2_X1 U4814 ( .A(n4173), .B(n4172), .ZN(n4180) );
  AOI22_X1 U4815 ( .A1(n4176), .A2(n4175), .B1(n4174), .B2(n4530), .ZN(n4177)
         );
  OAI21_X1 U4816 ( .B1(n4178), .B2(n4267), .A(n4177), .ZN(n4179) );
  AOI21_X1 U4817 ( .B1(n4180), .B2(n4519), .A(n4179), .ZN(n4241) );
  OAI21_X1 U4818 ( .B1(n4181), .B2(n4240), .A(n4241), .ZN(n4183) );
  NAND2_X1 U4819 ( .A1(n4183), .A2(n4182), .ZN(n4184) );
  OAI211_X1 U4820 ( .C1(n4242), .C2(n4186), .A(n4185), .B(n4184), .ZN(U3272)
         );
  NAND2_X1 U4821 ( .A1(n4634), .A2(n4274), .ZN(n4188) );
  NAND2_X1 U4822 ( .A1(n4631), .A2(REG1_REG_31__SCAN_IN), .ZN(n4187) );
  OAI211_X1 U4823 ( .C1(n4277), .C2(n4619), .A(n4188), .B(n4187), .ZN(U3549)
         );
  INV_X1 U4824 ( .A(n4361), .ZN(n4280) );
  INV_X1 U4825 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4194) );
  INV_X1 U4826 ( .A(n4191), .ZN(n4192) );
  AOI21_X1 U4827 ( .B1(n4193), .B2(n4530), .A(n4192), .ZN(n4362) );
  MUX2_X1 U4828 ( .A(n4194), .B(n4362), .S(n4634), .Z(n4195) );
  OAI21_X1 U4829 ( .B1(n4280), .B2(n4619), .A(n4195), .ZN(U3548) );
  INV_X1 U4830 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4202) );
  INV_X1 U4831 ( .A(n4196), .ZN(n4200) );
  OAI22_X1 U4832 ( .A1(n4198), .A2(n4267), .B1(n4197), .B2(n4265), .ZN(n4199)
         );
  MUX2_X1 U4833 ( .A(n4202), .B(n4281), .S(n4634), .Z(n4203) );
  OAI21_X1 U4834 ( .B1(n4619), .B2(n4284), .A(n4203), .ZN(U3545) );
  INV_X1 U4835 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4206) );
  AOI21_X1 U4836 ( .B1(n4205), .B2(n4590), .A(n4204), .ZN(n4285) );
  MUX2_X1 U4837 ( .A(n4206), .B(n4285), .S(n4634), .Z(n4207) );
  OAI21_X1 U4838 ( .B1(n4619), .B2(n4288), .A(n4207), .ZN(U3544) );
  INV_X1 U4839 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4210) );
  AOI21_X1 U4840 ( .B1(n4209), .B2(n4590), .A(n4208), .ZN(n4289) );
  MUX2_X1 U4841 ( .A(n4210), .B(n4289), .S(n4634), .Z(n4211) );
  OAI21_X1 U4842 ( .B1(n4619), .B2(n4292), .A(n4211), .ZN(U3543) );
  INV_X1 U4843 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4214) );
  AOI21_X1 U4844 ( .B1(n4213), .B2(n4590), .A(n4212), .ZN(n4293) );
  MUX2_X1 U4845 ( .A(n4214), .B(n4293), .S(n4634), .Z(n4215) );
  OAI21_X1 U4846 ( .B1(n4619), .B2(n4296), .A(n4215), .ZN(U3542) );
  INV_X1 U4847 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4218) );
  AOI21_X1 U4848 ( .B1(n4217), .B2(n4590), .A(n4216), .ZN(n4297) );
  MUX2_X1 U4849 ( .A(n4218), .B(n4297), .S(n4634), .Z(n4219) );
  OAI21_X1 U4850 ( .B1(n4619), .B2(n4300), .A(n4219), .ZN(U3541) );
  INV_X1 U4851 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4222) );
  AOI21_X1 U4852 ( .B1(n4221), .B2(n4590), .A(n4220), .ZN(n4301) );
  MUX2_X1 U4853 ( .A(n4222), .B(n4301), .S(n4634), .Z(n4223) );
  OAI21_X1 U4854 ( .B1(n4619), .B2(n4304), .A(n4223), .ZN(U3540) );
  INV_X1 U4855 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4229) );
  OAI22_X1 U4856 ( .A1(n4225), .A2(n4267), .B1(n4224), .B2(n4265), .ZN(n4227)
         );
  AOI211_X1 U4857 ( .C1(n4228), .C2(n4590), .A(n4227), .B(n4226), .ZN(n4305)
         );
  MUX2_X1 U4858 ( .A(n4229), .B(n4305), .S(n4634), .Z(n4230) );
  OAI21_X1 U4859 ( .B1(n4619), .B2(n4308), .A(n4230), .ZN(U3539) );
  INV_X1 U4860 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4234) );
  INV_X1 U4861 ( .A(n4231), .ZN(n4233) );
  AOI21_X1 U4862 ( .B1(n4601), .B2(n4233), .A(n4232), .ZN(n4309) );
  MUX2_X1 U4863 ( .A(n4234), .B(n4309), .S(n4634), .Z(n4235) );
  OAI21_X1 U4864 ( .B1(n4619), .B2(n4312), .A(n4235), .ZN(U3538) );
  NAND2_X1 U4865 ( .A1(n4236), .A2(n4590), .ZN(n4237) );
  AND2_X1 U4866 ( .A1(n4238), .A2(n4237), .ZN(n4313) );
  MUX2_X1 U4867 ( .A(n3949), .B(n4313), .S(n4634), .Z(n4239) );
  OAI21_X1 U4868 ( .B1(n4619), .B2(n4316), .A(n4239), .ZN(U3537) );
  OAI211_X1 U4869 ( .C1(n4242), .C2(n4250), .A(n4241), .B(n4240), .ZN(n4317)
         );
  MUX2_X1 U4870 ( .A(REG1_REG_18__SCAN_IN), .B(n4317), .S(n4634), .Z(U3536) );
  OAI22_X1 U4871 ( .A1(n4244), .A2(n4267), .B1(n4243), .B2(n4265), .ZN(n4245)
         );
  AOI21_X1 U4872 ( .B1(n4246), .B2(n4590), .A(n4245), .ZN(n4248) );
  AND2_X1 U4873 ( .A1(n4248), .A2(n4247), .ZN(n4318) );
  MUX2_X1 U4874 ( .A(n2834), .B(n4318), .S(n4634), .Z(n4249) );
  OAI21_X1 U4875 ( .B1(n4619), .B2(n4321), .A(n4249), .ZN(U3535) );
  OR2_X1 U4876 ( .A1(n4251), .A2(n4250), .ZN(n4252) );
  NAND2_X1 U4877 ( .A1(n4253), .A2(n4252), .ZN(n4322) );
  MUX2_X1 U4878 ( .A(n4322), .B(REG1_REG_16__SCAN_IN), .S(n4631), .Z(n4254) );
  AOI21_X1 U4879 ( .B1(n4255), .B2(n4325), .A(n4254), .ZN(n4256) );
  INV_X1 U4880 ( .A(n4256), .ZN(U3534) );
  INV_X1 U4881 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4262) );
  OAI22_X1 U4882 ( .A1(n4258), .A2(n4267), .B1(n4257), .B2(n4265), .ZN(n4259)
         );
  AOI211_X1 U4883 ( .C1(n4261), .C2(n4590), .A(n4260), .B(n4259), .ZN(n4327)
         );
  MUX2_X1 U4884 ( .A(n4262), .B(n4327), .S(n4634), .Z(n4263) );
  OAI21_X1 U4885 ( .B1(n4619), .B2(n4330), .A(n4263), .ZN(U3533) );
  INV_X1 U4886 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4272) );
  INV_X1 U4887 ( .A(n4264), .ZN(n4271) );
  OAI22_X1 U4888 ( .A1(n4268), .A2(n4267), .B1(n4266), .B2(n4265), .ZN(n4270)
         );
  AOI211_X1 U4889 ( .C1(n4601), .C2(n4271), .A(n4270), .B(n4269), .ZN(n4331)
         );
  MUX2_X1 U4890 ( .A(n4272), .B(n4331), .S(n4634), .Z(n4273) );
  OAI21_X1 U4891 ( .B1(n4619), .B2(n4334), .A(n4273), .ZN(U3532) );
  NAND2_X1 U4892 ( .A1(n4613), .A2(n4274), .ZN(n4276) );
  NAND2_X1 U4893 ( .A1(n4611), .A2(REG0_REG_31__SCAN_IN), .ZN(n4275) );
  OAI211_X1 U4894 ( .C1(n4277), .C2(n4580), .A(n4276), .B(n4275), .ZN(U3517)
         );
  INV_X1 U4895 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4278) );
  MUX2_X1 U4896 ( .A(n4278), .B(n4362), .S(n4613), .Z(n4279) );
  OAI21_X1 U4897 ( .B1(n4280), .B2(n4580), .A(n4279), .ZN(U3516) );
  INV_X1 U4898 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4282) );
  MUX2_X1 U4899 ( .A(n4282), .B(n4281), .S(n4613), .Z(n4283) );
  OAI21_X1 U4900 ( .B1(n4284), .B2(n4580), .A(n4283), .ZN(U3513) );
  INV_X1 U4901 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4286) );
  MUX2_X1 U4902 ( .A(n4286), .B(n4285), .S(n4613), .Z(n4287) );
  OAI21_X1 U4903 ( .B1(n4288), .B2(n4580), .A(n4287), .ZN(U3512) );
  INV_X1 U4904 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4290) );
  MUX2_X1 U4905 ( .A(n4290), .B(n4289), .S(n4613), .Z(n4291) );
  OAI21_X1 U4906 ( .B1(n4292), .B2(n4580), .A(n4291), .ZN(U3511) );
  INV_X1 U4907 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4294) );
  MUX2_X1 U4908 ( .A(n4294), .B(n4293), .S(n4613), .Z(n4295) );
  OAI21_X1 U4909 ( .B1(n4296), .B2(n4580), .A(n4295), .ZN(U3510) );
  INV_X1 U4910 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4298) );
  MUX2_X1 U4911 ( .A(n4298), .B(n4297), .S(n4613), .Z(n4299) );
  OAI21_X1 U4912 ( .B1(n4300), .B2(n4580), .A(n4299), .ZN(U3509) );
  INV_X1 U4913 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4302) );
  MUX2_X1 U4914 ( .A(n4302), .B(n4301), .S(n4613), .Z(n4303) );
  OAI21_X1 U4915 ( .B1(n4304), .B2(n4580), .A(n4303), .ZN(U3508) );
  INV_X1 U4916 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4306) );
  MUX2_X1 U4917 ( .A(n4306), .B(n4305), .S(n4613), .Z(n4307) );
  OAI21_X1 U4918 ( .B1(n4308), .B2(n4580), .A(n4307), .ZN(U3507) );
  INV_X1 U4919 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4310) );
  MUX2_X1 U4920 ( .A(n4310), .B(n4309), .S(n4613), .Z(n4311) );
  OAI21_X1 U4921 ( .B1(n4312), .B2(n4580), .A(n4311), .ZN(U3506) );
  INV_X1 U4922 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4314) );
  MUX2_X1 U4923 ( .A(n4314), .B(n4313), .S(n4613), .Z(n4315) );
  OAI21_X1 U4924 ( .B1(n4316), .B2(n4580), .A(n4315), .ZN(U3505) );
  MUX2_X1 U4925 ( .A(REG0_REG_18__SCAN_IN), .B(n4317), .S(n4613), .Z(U3503) );
  INV_X1 U4926 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4319) );
  MUX2_X1 U4927 ( .A(n4319), .B(n4318), .S(n4613), .Z(n4320) );
  OAI21_X1 U4928 ( .B1(n4321), .B2(n4580), .A(n4320), .ZN(U3501) );
  MUX2_X1 U4929 ( .A(n4322), .B(REG0_REG_16__SCAN_IN), .S(n4611), .Z(n4323) );
  AOI21_X1 U4930 ( .B1(n4325), .B2(n4324), .A(n4323), .ZN(n4326) );
  INV_X1 U4931 ( .A(n4326), .ZN(U3499) );
  INV_X1 U4932 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4328) );
  MUX2_X1 U4933 ( .A(n4328), .B(n4327), .S(n4613), .Z(n4329) );
  OAI21_X1 U4934 ( .B1(n4330), .B2(n4580), .A(n4329), .ZN(U3497) );
  INV_X1 U4935 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4332) );
  MUX2_X1 U4936 ( .A(n4332), .B(n4331), .S(n4613), .Z(n4333) );
  OAI21_X1 U4937 ( .B1(n4334), .B2(n4580), .A(n4333), .ZN(U3495) );
  MUX2_X1 U4938 ( .A(DATAI_30_), .B(n4335), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4939 ( .A(n4336), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4940 ( .A(n2740), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U4941 ( .A(DATAI_22_), .B(n4337), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U4942 ( .A(DATAI_20_), .B(n4338), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4943 ( .A(DATAI_4_), .B(n4339), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4944 ( .A(DATAI_3_), .B(n4340), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U4945 ( .A(n2221), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  INV_X1 U4946 ( .A(DATAI_28_), .ZN(n4342) );
  AOI22_X1 U4947 ( .A1(STATE_REG_SCAN_IN), .A2(n4343), .B1(n4342), .B2(U3149), 
        .ZN(U3324) );
  INV_X1 U4948 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4988) );
  NOR2_X1 U4949 ( .A1(STATE_REG_SCAN_IN), .A2(n4988), .ZN(n4490) );
  OAI22_X1 U4950 ( .A1(n4347), .A2(n4346), .B1(n4345), .B2(n4344), .ZN(n4348)
         );
  AOI211_X1 U4951 ( .C1(n4350), .C2(n4349), .A(n4490), .B(n4348), .ZN(n4358)
         );
  AOI21_X1 U4952 ( .B1(n4352), .B2(n4351), .A(n3734), .ZN(n4353) );
  XOR2_X1 U4953 ( .A(n4354), .B(n4353), .Z(n4356) );
  NAND2_X1 U4954 ( .A1(n4356), .A2(n4355), .ZN(n4357) );
  OAI211_X1 U4955 ( .C1(n4360), .C2(n4359), .A(n4358), .B(n4357), .ZN(U3223)
         );
  INV_X1 U4956 ( .A(n4365), .ZN(n4363) );
  OAI211_X1 U4957 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4364), .A(n4366), .B(n4363), 
        .ZN(n4369) );
  INV_X1 U4958 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4614) );
  AOI22_X1 U4959 ( .A1(n4366), .A2(n4365), .B1(n4502), .B2(n4614), .ZN(n4368)
         );
  AOI22_X1 U4960 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4501), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4367) );
  OAI221_X1 U4961 ( .B1(IR_REG_0__SCAN_IN), .B2(n4369), .C1(n2266), .C2(n4368), 
        .A(n4367), .ZN(U3240) );
  INV_X1 U4962 ( .A(n4502), .ZN(n4380) );
  AOI211_X1 U4963 ( .C1(n4372), .C2(n4371), .A(n4370), .B(n4380), .ZN(n4374)
         );
  AOI211_X1 U4964 ( .C1(n4501), .C2(ADDR_REG_5__SCAN_IN), .A(n4374), .B(n4373), 
        .ZN(n4379) );
  OAI211_X1 U4965 ( .C1(n4377), .C2(n4376), .A(n4456), .B(n4375), .ZN(n4378)
         );
  OAI211_X1 U4966 ( .C1(n4508), .C2(n4567), .A(n4379), .B(n4378), .ZN(U3245)
         );
  AOI211_X1 U4967 ( .C1(n4383), .C2(n4382), .A(n4381), .B(n4380), .ZN(n4385)
         );
  AOI211_X1 U4968 ( .C1(n4501), .C2(ADDR_REG_6__SCAN_IN), .A(n4385), .B(n4384), 
        .ZN(n4389) );
  OAI211_X1 U4969 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4387), .A(n4456), .B(n4386), 
        .ZN(n4388) );
  OAI211_X1 U4970 ( .C1(n4508), .C2(n2772), .A(n4389), .B(n4388), .ZN(U3246)
         );
  INV_X1 U4971 ( .A(n4390), .ZN(n4392) );
  NAND2_X1 U4972 ( .A1(n4392), .A2(n4391), .ZN(n4394) );
  OAI21_X1 U4973 ( .B1(n4395), .B2(n4394), .A(n4502), .ZN(n4393) );
  AOI21_X1 U4974 ( .B1(n4395), .B2(n4394), .A(n4393), .ZN(n4397) );
  AOI211_X1 U4975 ( .C1(n4501), .C2(ADDR_REG_7__SCAN_IN), .A(n4397), .B(n4396), 
        .ZN(n4402) );
  OAI211_X1 U4976 ( .C1(n4400), .C2(n4399), .A(n4456), .B(n4398), .ZN(n4401)
         );
  OAI211_X1 U4977 ( .C1(n4508), .C2(n4565), .A(n4402), .B(n4401), .ZN(U3247)
         );
  OAI211_X1 U4978 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4405), .A(n4502), .B(n4404), 
        .ZN(n4409) );
  OAI211_X1 U4979 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4407), .A(n4456), .B(n4406), 
        .ZN(n4408) );
  OAI211_X1 U4980 ( .C1(n4508), .C2(n2814), .A(n4409), .B(n4408), .ZN(n4410)
         );
  AOI211_X1 U4981 ( .C1(n4501), .C2(ADDR_REG_8__SCAN_IN), .A(n4411), .B(n4410), 
        .ZN(n4412) );
  INV_X1 U4982 ( .A(n4412), .ZN(U3248) );
  OAI211_X1 U4983 ( .C1(n4415), .C2(n4414), .A(n4502), .B(n4413), .ZN(n4420)
         );
  OAI211_X1 U4984 ( .C1(n4418), .C2(n4417), .A(n4456), .B(n4416), .ZN(n4419)
         );
  OAI211_X1 U4985 ( .C1(n4508), .C2(n4564), .A(n4420), .B(n4419), .ZN(n4421)
         );
  AOI211_X1 U4986 ( .C1(n4501), .C2(ADDR_REG_9__SCAN_IN), .A(n4422), .B(n4421), 
        .ZN(n4423) );
  INV_X1 U4987 ( .A(n4423), .ZN(U3249) );
  OAI211_X1 U4988 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4426), .A(n4502), .B(n4425), .ZN(n4430) );
  OAI211_X1 U4989 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4428), .A(n4456), .B(n4427), .ZN(n4429) );
  OAI211_X1 U4990 ( .C1(n4508), .C2(n2779), .A(n4430), .B(n4429), .ZN(n4431)
         );
  AOI211_X1 U4991 ( .C1(n4501), .C2(ADDR_REG_10__SCAN_IN), .A(n4432), .B(n4431), .ZN(n4433) );
  INV_X1 U4992 ( .A(n4433), .ZN(U3250) );
  OAI211_X1 U4993 ( .C1(n4436), .C2(n4435), .A(n4502), .B(n4434), .ZN(n4441)
         );
  OAI211_X1 U4994 ( .C1(n4439), .C2(n4438), .A(n4456), .B(n4437), .ZN(n4440)
         );
  OAI211_X1 U4995 ( .C1(n4508), .C2(n4563), .A(n4441), .B(n4440), .ZN(n4442)
         );
  AOI211_X1 U4996 ( .C1(n4501), .C2(ADDR_REG_11__SCAN_IN), .A(n4443), .B(n4442), .ZN(n4444) );
  INV_X1 U4997 ( .A(n4444), .ZN(U3251) );
  OAI211_X1 U4998 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4446), .A(n4456), .B(n4445), .ZN(n4448) );
  NAND2_X1 U4999 ( .A1(n4448), .A2(n4447), .ZN(n4449) );
  AOI21_X1 U5000 ( .B1(n4501), .B2(ADDR_REG_12__SCAN_IN), .A(n4449), .ZN(n4453) );
  OAI211_X1 U5001 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4451), .A(n4502), .B(n4450), .ZN(n4452) );
  OAI211_X1 U5002 ( .C1(n4508), .C2(n2783), .A(n4453), .B(n4452), .ZN(U3252)
         );
  AOI21_X1 U5003 ( .B1(n4455), .B2(n4561), .A(n4454), .ZN(n4459) );
  OAI21_X1 U5004 ( .B1(n4459), .B2(n4458), .A(n4456), .ZN(n4457) );
  AOI21_X1 U5005 ( .B1(n4459), .B2(n4458), .A(n4457), .ZN(n4460) );
  AOI211_X1 U5006 ( .C1(n4501), .C2(ADDR_REG_13__SCAN_IN), .A(n4461), .B(n4460), .ZN(n4466) );
  OAI211_X1 U5007 ( .C1(n4464), .C2(n4463), .A(n4502), .B(n4462), .ZN(n4465)
         );
  OAI211_X1 U5008 ( .C1(n4508), .C2(n4561), .A(n4466), .B(n4465), .ZN(U3253)
         );
  INV_X1 U5009 ( .A(n4467), .ZN(n4472) );
  AOI211_X1 U5010 ( .C1(n4470), .C2(n4469), .A(n4468), .B(n4495), .ZN(n4471)
         );
  AOI211_X1 U5011 ( .C1(n4501), .C2(ADDR_REG_14__SCAN_IN), .A(n4472), .B(n4471), .ZN(n4476) );
  OAI211_X1 U5012 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4474), .A(n4502), .B(n4473), .ZN(n4475) );
  OAI211_X1 U5013 ( .C1(n4508), .C2(n4560), .A(n4476), .B(n4475), .ZN(U3254)
         );
  AOI211_X1 U5014 ( .C1(n4478), .C2(n4477), .A(n2233), .B(n4495), .ZN(n4479)
         );
  AOI211_X1 U5015 ( .C1(n4501), .C2(ADDR_REG_15__SCAN_IN), .A(n4480), .B(n4479), .ZN(n4485) );
  OAI211_X1 U5016 ( .C1(n4483), .C2(n4482), .A(n4502), .B(n4481), .ZN(n4484)
         );
  OAI211_X1 U5017 ( .C1(n4508), .C2(n4559), .A(n4485), .B(n4484), .ZN(U3255)
         );
  AOI221_X1 U5018 ( .B1(n4488), .B2(n4487), .C1(n4486), .C2(n4487), .A(n4495), 
        .ZN(n4489) );
  AOI211_X1 U5019 ( .C1(n4501), .C2(ADDR_REG_16__SCAN_IN), .A(n4490), .B(n4489), .ZN(n4494) );
  OAI221_X1 U5020 ( .B1(n4492), .B2(REG1_REG_16__SCAN_IN), .C1(n4492), .C2(
        n4491), .A(n4502), .ZN(n4493) );
  OAI211_X1 U5021 ( .C1(n4508), .C2(n4558), .A(n4494), .B(n4493), .ZN(U3256)
         );
  AOI221_X1 U5022 ( .B1(n4498), .B2(n4497), .C1(n4496), .C2(n4497), .A(n4495), 
        .ZN(n4499) );
  AOI211_X1 U5023 ( .C1(n4501), .C2(ADDR_REG_17__SCAN_IN), .A(n4500), .B(n4499), .ZN(n4507) );
  OAI221_X1 U5024 ( .B1(n4505), .B2(n4504), .C1(n4505), .C2(n4503), .A(n4502), 
        .ZN(n4506) );
  OAI211_X1 U5025 ( .C1(n4508), .C2(n4557), .A(n4507), .B(n4506), .ZN(U3257)
         );
  XOR2_X1 U5026 ( .A(n4514), .B(n4509), .Z(n4520) );
  AOI22_X1 U5027 ( .A1(n4511), .A2(n4532), .B1(n4530), .B2(n4510), .ZN(n4512)
         );
  OAI21_X1 U5028 ( .B1(n4513), .B2(n4535), .A(n4512), .ZN(n4518) );
  XOR2_X1 U5029 ( .A(n4515), .B(n4514), .Z(n4608) );
  NOR2_X1 U5030 ( .A1(n4608), .A2(n4516), .ZN(n4517) );
  AOI211_X1 U5031 ( .C1(n4520), .C2(n4519), .A(n4518), .B(n4517), .ZN(n4604)
         );
  AOI22_X1 U5032 ( .A1(n4521), .A2(n4543), .B1(REG2_REG_11__SCAN_IN), .B2(
        n2222), .ZN(n4527) );
  INV_X1 U5033 ( .A(n4608), .ZN(n4525) );
  OAI21_X1 U5034 ( .B1(n4597), .B2(n4523), .A(n4522), .ZN(n4605) );
  INV_X1 U5035 ( .A(n4605), .ZN(n4524) );
  AOI22_X1 U5036 ( .A1(n4525), .A2(n4549), .B1(n4548), .B2(n4524), .ZN(n4526)
         );
  OAI211_X1 U5037 ( .C1(n2222), .C2(n4604), .A(n4527), .B(n4526), .ZN(U3279)
         );
  OR2_X1 U5038 ( .A1(n2688), .A2(n2234), .ZN(n4528) );
  AND2_X1 U5039 ( .A1(n4529), .A2(n4528), .ZN(n4576) );
  AOI22_X1 U5040 ( .A1(n4533), .A2(n4532), .B1(n4531), .B2(n4530), .ZN(n4534)
         );
  OAI21_X1 U5041 ( .B1(n4536), .B2(n4535), .A(n4534), .ZN(n4541) );
  AOI21_X1 U5042 ( .B1(n4539), .B2(n4538), .A(n4537), .ZN(n4540) );
  AOI211_X1 U5043 ( .C1(n4576), .C2(n4542), .A(n4541), .B(n4540), .ZN(n4573)
         );
  AOI22_X1 U5044 ( .A1(REG3_REG_1__SCAN_IN), .A2(n4543), .B1(
        REG2_REG_1__SCAN_IN), .B2(n2222), .ZN(n4551) );
  OAI21_X1 U5045 ( .B1(n4546), .B2(n4545), .A(n4544), .ZN(n4572) );
  INV_X1 U5046 ( .A(n4572), .ZN(n4547) );
  AOI22_X1 U5047 ( .A1(n4549), .A2(n4576), .B1(n4548), .B2(n4547), .ZN(n4550)
         );
  OAI211_X1 U5048 ( .C1(n2222), .C2(n4573), .A(n4551), .B(n4550), .ZN(U3289)
         );
  INV_X1 U5049 ( .A(D_REG_31__SCAN_IN), .ZN(n4926) );
  NOR2_X1 U5050 ( .A1(n4553), .A2(n4926), .ZN(U3291) );
  AND2_X1 U5051 ( .A1(n4552), .A2(D_REG_30__SCAN_IN), .ZN(U3292) );
  INV_X1 U5052 ( .A(D_REG_29__SCAN_IN), .ZN(n4907) );
  NOR2_X1 U5053 ( .A1(n4553), .A2(n4907), .ZN(U3293) );
  INV_X1 U5054 ( .A(D_REG_28__SCAN_IN), .ZN(n4764) );
  NOR2_X1 U5055 ( .A1(n4553), .A2(n4764), .ZN(U3294) );
  INV_X1 U5056 ( .A(D_REG_27__SCAN_IN), .ZN(n4929) );
  NOR2_X1 U5057 ( .A1(n4553), .A2(n4929), .ZN(U3295) );
  AND2_X1 U5058 ( .A1(n4552), .A2(D_REG_26__SCAN_IN), .ZN(U3296) );
  INV_X1 U5059 ( .A(D_REG_25__SCAN_IN), .ZN(n4754) );
  NOR2_X1 U5060 ( .A1(n4553), .A2(n4754), .ZN(U3297) );
  INV_X1 U5061 ( .A(D_REG_24__SCAN_IN), .ZN(n4920) );
  NOR2_X1 U5062 ( .A1(n4553), .A2(n4920), .ZN(U3298) );
  INV_X1 U5063 ( .A(D_REG_23__SCAN_IN), .ZN(n4728) );
  NOR2_X1 U5064 ( .A1(n4553), .A2(n4728), .ZN(U3299) );
  INV_X1 U5065 ( .A(D_REG_22__SCAN_IN), .ZN(n4740) );
  NOR2_X1 U5066 ( .A1(n4553), .A2(n4740), .ZN(U3300) );
  INV_X1 U5067 ( .A(D_REG_21__SCAN_IN), .ZN(n4738) );
  NOR2_X1 U5068 ( .A1(n4553), .A2(n4738), .ZN(U3301) );
  INV_X1 U5069 ( .A(D_REG_20__SCAN_IN), .ZN(n4944) );
  NOR2_X1 U5070 ( .A1(n4553), .A2(n4944), .ZN(U3302) );
  AND2_X1 U5071 ( .A1(n4552), .A2(D_REG_19__SCAN_IN), .ZN(U3303) );
  INV_X1 U5072 ( .A(D_REG_18__SCAN_IN), .ZN(n4718) );
  NOR2_X1 U5073 ( .A1(n4553), .A2(n4718), .ZN(U3304) );
  AND2_X1 U5074 ( .A1(n4552), .A2(D_REG_17__SCAN_IN), .ZN(U3305) );
  INV_X1 U5075 ( .A(D_REG_16__SCAN_IN), .ZN(n4943) );
  NOR2_X1 U5076 ( .A1(n4553), .A2(n4943), .ZN(U3306) );
  INV_X1 U5077 ( .A(D_REG_15__SCAN_IN), .ZN(n4923) );
  NOR2_X1 U5078 ( .A1(n4553), .A2(n4923), .ZN(U3307) );
  INV_X1 U5079 ( .A(D_REG_14__SCAN_IN), .ZN(n4913) );
  NOR2_X1 U5080 ( .A1(n4553), .A2(n4913), .ZN(U3308) );
  INV_X1 U5081 ( .A(D_REG_13__SCAN_IN), .ZN(n4921) );
  NOR2_X1 U5082 ( .A1(n4553), .A2(n4921), .ZN(U3309) );
  INV_X1 U5083 ( .A(D_REG_12__SCAN_IN), .ZN(n4927) );
  NOR2_X1 U5084 ( .A1(n4553), .A2(n4927), .ZN(U3310) );
  INV_X1 U5085 ( .A(D_REG_11__SCAN_IN), .ZN(n4924) );
  NOR2_X1 U5086 ( .A1(n4553), .A2(n4924), .ZN(U3311) );
  INV_X1 U5087 ( .A(D_REG_10__SCAN_IN), .ZN(n4940) );
  NOR2_X1 U5088 ( .A1(n4553), .A2(n4940), .ZN(U3312) );
  AND2_X1 U5089 ( .A1(n4552), .A2(D_REG_9__SCAN_IN), .ZN(U3313) );
  INV_X1 U5090 ( .A(D_REG_8__SCAN_IN), .ZN(n4912) );
  NOR2_X1 U5091 ( .A1(n4553), .A2(n4912), .ZN(U3314) );
  AND2_X1 U5092 ( .A1(n4552), .A2(D_REG_7__SCAN_IN), .ZN(U3315) );
  AND2_X1 U5093 ( .A1(n4552), .A2(D_REG_6__SCAN_IN), .ZN(U3316) );
  INV_X1 U5094 ( .A(D_REG_5__SCAN_IN), .ZN(n4930) );
  NOR2_X1 U5095 ( .A1(n4553), .A2(n4930), .ZN(U3317) );
  AND2_X1 U5096 ( .A1(n4552), .A2(D_REG_4__SCAN_IN), .ZN(U3318) );
  INV_X1 U5097 ( .A(D_REG_3__SCAN_IN), .ZN(n4941) );
  NOR2_X1 U5098 ( .A1(n4553), .A2(n4941), .ZN(U3319) );
  INV_X1 U5099 ( .A(D_REG_2__SCAN_IN), .ZN(n4775) );
  NOR2_X1 U5100 ( .A1(n4553), .A2(n4775), .ZN(U3320) );
  INV_X1 U5101 ( .A(DATAI_23_), .ZN(n4976) );
  AOI21_X1 U5102 ( .B1(U3149), .B2(n4976), .A(n4554), .ZN(U3329) );
  INV_X1 U5103 ( .A(DATAI_18_), .ZN(n4555) );
  AOI22_X1 U5104 ( .A1(STATE_REG_SCAN_IN), .A2(n4556), .B1(n4555), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U5105 ( .A(DATAI_17_), .ZN(n4954) );
  AOI22_X1 U5106 ( .A1(STATE_REG_SCAN_IN), .A2(n4557), .B1(n4954), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5107 ( .A(DATAI_16_), .ZN(n4958) );
  AOI22_X1 U5108 ( .A1(STATE_REG_SCAN_IN), .A2(n4558), .B1(n4958), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5109 ( .A(DATAI_15_), .ZN(n4983) );
  AOI22_X1 U5110 ( .A1(STATE_REG_SCAN_IN), .A2(n4559), .B1(n4983), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5111 ( .A(DATAI_14_), .ZN(n4974) );
  AOI22_X1 U5112 ( .A1(STATE_REG_SCAN_IN), .A2(n4560), .B1(n4974), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U5113 ( .A1(STATE_REG_SCAN_IN), .A2(n4561), .B1(n2533), .B2(U3149), 
        .ZN(U3339) );
  AOI22_X1 U5114 ( .A1(STATE_REG_SCAN_IN), .A2(n2783), .B1(n4716), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5115 ( .A(DATAI_11_), .ZN(n4562) );
  AOI22_X1 U5116 ( .A1(STATE_REG_SCAN_IN), .A2(n4563), .B1(n4562), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5117 ( .A(DATAI_10_), .ZN(n4948) );
  AOI22_X1 U5118 ( .A1(STATE_REG_SCAN_IN), .A2(n2779), .B1(n4948), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5119 ( .A(DATAI_9_), .ZN(n4915) );
  AOI22_X1 U5120 ( .A1(STATE_REG_SCAN_IN), .A2(n4564), .B1(n4915), .B2(U3149), 
        .ZN(U3343) );
  INV_X1 U5121 ( .A(DATAI_8_), .ZN(n4946) );
  AOI22_X1 U5122 ( .A1(STATE_REG_SCAN_IN), .A2(n2814), .B1(n4946), .B2(U3149), 
        .ZN(U3344) );
  INV_X1 U5123 ( .A(DATAI_7_), .ZN(n4957) );
  AOI22_X1 U5124 ( .A1(STATE_REG_SCAN_IN), .A2(n4565), .B1(n4957), .B2(U3149), 
        .ZN(U3345) );
  INV_X1 U5125 ( .A(DATAI_6_), .ZN(n4566) );
  AOI22_X1 U5126 ( .A1(STATE_REG_SCAN_IN), .A2(n2772), .B1(n4566), .B2(U3149), 
        .ZN(U3346) );
  INV_X1 U5127 ( .A(DATAI_5_), .ZN(n4985) );
  AOI22_X1 U5128 ( .A1(STATE_REG_SCAN_IN), .A2(n4567), .B1(n4985), .B2(U3149), 
        .ZN(U3347) );
  OAI211_X1 U5129 ( .C1(n4570), .C2(n4607), .A(n4569), .B(n4568), .ZN(n4571)
         );
  INV_X1 U5130 ( .A(n4571), .ZN(n4615) );
  INV_X1 U5131 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4780) );
  AOI22_X1 U5132 ( .A1(n4613), .A2(n4615), .B1(n4780), .B2(n4611), .ZN(U3467)
         );
  NOR2_X1 U5133 ( .A1(n4572), .A2(n4606), .ZN(n4575) );
  INV_X1 U5134 ( .A(n4573), .ZN(n4574) );
  AOI211_X1 U5135 ( .C1(n4576), .C2(n4601), .A(n4575), .B(n4574), .ZN(n4617)
         );
  INV_X1 U5136 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4731) );
  AOI22_X1 U5137 ( .A1(n4613), .A2(n4617), .B1(n4731), .B2(n4611), .ZN(U3469)
         );
  AOI21_X1 U5138 ( .B1(n4601), .B2(n4578), .A(n4577), .ZN(n4622) );
  INV_X1 U5139 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4579) );
  OAI22_X1 U5140 ( .A1(n4580), .A2(n4618), .B1(n4613), .B2(n4579), .ZN(n4581)
         );
  INV_X1 U5141 ( .A(n4581), .ZN(n4582) );
  OAI21_X1 U5142 ( .B1(n4622), .B2(n4611), .A(n4582), .ZN(U3471) );
  INV_X1 U5143 ( .A(n4583), .ZN(n4585) );
  AOI211_X1 U5144 ( .C1(n4586), .C2(n4601), .A(n4585), .B(n4584), .ZN(n4624)
         );
  INV_X1 U5145 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4587) );
  AOI22_X1 U5146 ( .A1(n4613), .A2(n4624), .B1(n4587), .B2(n4611), .ZN(U3475)
         );
  AOI211_X1 U5147 ( .C1(n4591), .C2(n4590), .A(n4589), .B(n4588), .ZN(n4626)
         );
  INV_X1 U5148 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4894) );
  AOI22_X1 U5149 ( .A1(n4613), .A2(n4626), .B1(n4894), .B2(n4611), .ZN(U3481)
         );
  NOR3_X1 U5150 ( .A1(n4593), .A2(n4592), .A3(n4606), .ZN(n4595) );
  AOI211_X1 U5151 ( .C1(n4596), .C2(n4601), .A(n4595), .B(n4594), .ZN(n4628)
         );
  INV_X1 U5152 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4893) );
  AOI22_X1 U5153 ( .A1(n4613), .A2(n4628), .B1(n4893), .B2(n4611), .ZN(U3483)
         );
  NOR3_X1 U5154 ( .A1(n4598), .A2(n4597), .A3(n4606), .ZN(n4600) );
  AOI211_X1 U5155 ( .C1(n4602), .C2(n4601), .A(n4600), .B(n4599), .ZN(n4630)
         );
  INV_X1 U5156 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4603) );
  AOI22_X1 U5157 ( .A1(n4613), .A2(n4630), .B1(n4603), .B2(n4611), .ZN(U3487)
         );
  INV_X1 U5158 ( .A(n4604), .ZN(n4610) );
  OAI22_X1 U5159 ( .A1(n4608), .A2(n4607), .B1(n4606), .B2(n4605), .ZN(n4609)
         );
  NOR2_X1 U5160 ( .A1(n4610), .A2(n4609), .ZN(n4633) );
  INV_X1 U5161 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4612) );
  AOI22_X1 U5162 ( .A1(n4613), .A2(n4633), .B1(n4612), .B2(n4611), .ZN(U3489)
         );
  AOI22_X1 U5163 ( .A1(n4634), .A2(n4615), .B1(n4614), .B2(n4631), .ZN(U3518)
         );
  INV_X1 U5164 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4616) );
  AOI22_X1 U5165 ( .A1(n4634), .A2(n4617), .B1(n4616), .B2(n4631), .ZN(U3519)
         );
  OAI22_X1 U5166 ( .A1(n4619), .A2(n4618), .B1(n4634), .B2(n2802), .ZN(n4620)
         );
  INV_X1 U5167 ( .A(n4620), .ZN(n4621) );
  OAI21_X1 U5168 ( .B1(n4622), .B2(n4631), .A(n4621), .ZN(U3520) );
  INV_X1 U5169 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4623) );
  AOI22_X1 U5170 ( .A1(n4634), .A2(n4624), .B1(n4623), .B2(n4631), .ZN(U3522)
         );
  INV_X1 U5171 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4625) );
  AOI22_X1 U5172 ( .A1(n4634), .A2(n4626), .B1(n4625), .B2(n4631), .ZN(U3525)
         );
  INV_X1 U5173 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4627) );
  AOI22_X1 U5174 ( .A1(n4634), .A2(n4628), .B1(n4627), .B2(n4631), .ZN(U3526)
         );
  INV_X1 U5175 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4629) );
  AOI22_X1 U5176 ( .A1(n4634), .A2(n4630), .B1(n4629), .B2(n4631), .ZN(U3528)
         );
  AOI22_X1 U5177 ( .A1(n4634), .A2(n4633), .B1(n4632), .B2(n4631), .ZN(U3529)
         );
  OAI22_X1 U5178 ( .A1(DATAI_16_), .A2(keyinput_g15), .B1(DATAI_18_), .B2(
        keyinput_g13), .ZN(n4635) );
  AOI221_X1 U5179 ( .B1(DATAI_16_), .B2(keyinput_g15), .C1(keyinput_g13), .C2(
        DATAI_18_), .A(n4635), .ZN(n4642) );
  OAI22_X1 U5180 ( .A1(REG3_REG_24__SCAN_IN), .A2(keyinput_g49), .B1(
        keyinput_g3), .B2(DATAI_28_), .ZN(n4636) );
  AOI221_X1 U5181 ( .B1(REG3_REG_24__SCAN_IN), .B2(keyinput_g49), .C1(
        DATAI_28_), .C2(keyinput_g3), .A(n4636), .ZN(n4641) );
  OAI22_X1 U5182 ( .A1(REG3_REG_4__SCAN_IN), .A2(keyinput_g50), .B1(
        keyinput_g11), .B2(DATAI_20_), .ZN(n4637) );
  AOI221_X1 U5183 ( .B1(REG3_REG_4__SCAN_IN), .B2(keyinput_g50), .C1(DATAI_20_), .C2(keyinput_g11), .A(n4637), .ZN(n4640) );
  OAI22_X1 U5184 ( .A1(IR_REG_16__SCAN_IN), .A2(keyinput_g71), .B1(DATAI_11_), 
        .B2(keyinput_g20), .ZN(n4638) );
  AOI221_X1 U5185 ( .B1(IR_REG_16__SCAN_IN), .B2(keyinput_g71), .C1(
        keyinput_g20), .C2(DATAI_11_), .A(n4638), .ZN(n4639) );
  NAND4_X1 U5186 ( .A1(n4642), .A2(n4641), .A3(n4640), .A4(n4639), .ZN(n4670)
         );
  OAI22_X1 U5187 ( .A1(IR_REG_26__SCAN_IN), .A2(keyinput_g81), .B1(
        keyinput_g103), .B2(D_REG_16__SCAN_IN), .ZN(n4643) );
  AOI221_X1 U5188 ( .B1(IR_REG_26__SCAN_IN), .B2(keyinput_g81), .C1(
        D_REG_16__SCAN_IN), .C2(keyinput_g103), .A(n4643), .ZN(n4650) );
  OAI22_X1 U5189 ( .A1(STATE_REG_SCAN_IN), .A2(keyinput_g32), .B1(DATAI_1_), 
        .B2(keyinput_g30), .ZN(n4644) );
  AOI221_X1 U5190 ( .B1(STATE_REG_SCAN_IN), .B2(keyinput_g32), .C1(
        keyinput_g30), .C2(DATAI_1_), .A(n4644), .ZN(n4649) );
  OAI22_X1 U5191 ( .A1(D_REG_9__SCAN_IN), .A2(keyinput_g96), .B1(keyinput_g48), 
        .B2(REG3_REG_17__SCAN_IN), .ZN(n4645) );
  AOI221_X1 U5192 ( .B1(D_REG_9__SCAN_IN), .B2(keyinput_g96), .C1(
        REG3_REG_17__SCAN_IN), .C2(keyinput_g48), .A(n4645), .ZN(n4648) );
  OAI22_X1 U5193 ( .A1(D_REG_6__SCAN_IN), .A2(keyinput_g93), .B1(DATAI_6_), 
        .B2(keyinput_g25), .ZN(n4646) );
  AOI221_X1 U5194 ( .B1(D_REG_6__SCAN_IN), .B2(keyinput_g93), .C1(keyinput_g25), .C2(DATAI_6_), .A(n4646), .ZN(n4647) );
  NAND4_X1 U5195 ( .A1(n4650), .A2(n4649), .A3(n4648), .A4(n4647), .ZN(n4669)
         );
  OAI22_X1 U5196 ( .A1(REG0_REG_3__SCAN_IN), .A2(keyinput_g122), .B1(
        keyinput_g123), .B2(REG0_REG_4__SCAN_IN), .ZN(n4651) );
  AOI221_X1 U5197 ( .B1(REG0_REG_3__SCAN_IN), .B2(keyinput_g122), .C1(
        REG0_REG_4__SCAN_IN), .C2(keyinput_g123), .A(n4651), .ZN(n4658) );
  OAI22_X1 U5198 ( .A1(IR_REG_19__SCAN_IN), .A2(keyinput_g74), .B1(
        keyinput_g67), .B2(IR_REG_12__SCAN_IN), .ZN(n4652) );
  AOI221_X1 U5199 ( .B1(IR_REG_19__SCAN_IN), .B2(keyinput_g74), .C1(
        IR_REG_12__SCAN_IN), .C2(keyinput_g67), .A(n4652), .ZN(n4657) );
  OAI22_X1 U5200 ( .A1(D_REG_29__SCAN_IN), .A2(keyinput_g116), .B1(
        D_REG_14__SCAN_IN), .B2(keyinput_g101), .ZN(n4653) );
  AOI221_X1 U5201 ( .B1(D_REG_29__SCAN_IN), .B2(keyinput_g116), .C1(
        keyinput_g101), .C2(D_REG_14__SCAN_IN), .A(n4653), .ZN(n4656) );
  OAI22_X1 U5202 ( .A1(D_REG_13__SCAN_IN), .A2(keyinput_g100), .B1(
        D_REG_24__SCAN_IN), .B2(keyinput_g111), .ZN(n4654) );
  AOI221_X1 U5203 ( .B1(D_REG_13__SCAN_IN), .B2(keyinput_g100), .C1(
        keyinput_g111), .C2(D_REG_24__SCAN_IN), .A(n4654), .ZN(n4655) );
  NAND4_X1 U5204 ( .A1(n4658), .A2(n4657), .A3(n4656), .A4(n4655), .ZN(n4668)
         );
  OAI22_X1 U5205 ( .A1(D_REG_12__SCAN_IN), .A2(keyinput_g99), .B1(
        D_REG_27__SCAN_IN), .B2(keyinput_g114), .ZN(n4659) );
  AOI221_X1 U5206 ( .B1(D_REG_12__SCAN_IN), .B2(keyinput_g99), .C1(
        keyinput_g114), .C2(D_REG_27__SCAN_IN), .A(n4659), .ZN(n4666) );
  OAI22_X1 U5207 ( .A1(REG3_REG_23__SCAN_IN), .A2(keyinput_g36), .B1(
        REG3_REG_12__SCAN_IN), .B2(keyinput_g44), .ZN(n4660) );
  AOI221_X1 U5208 ( .B1(REG3_REG_23__SCAN_IN), .B2(keyinput_g36), .C1(
        keyinput_g44), .C2(REG3_REG_12__SCAN_IN), .A(n4660), .ZN(n4665) );
  OAI22_X1 U5209 ( .A1(IR_REG_10__SCAN_IN), .A2(keyinput_g65), .B1(
        REG3_REG_16__SCAN_IN), .B2(keyinput_g46), .ZN(n4661) );
  AOI221_X1 U5210 ( .B1(IR_REG_10__SCAN_IN), .B2(keyinput_g65), .C1(
        keyinput_g46), .C2(REG3_REG_16__SCAN_IN), .A(n4661), .ZN(n4664) );
  OAI22_X1 U5211 ( .A1(IR_REG_24__SCAN_IN), .A2(keyinput_g79), .B1(
        IR_REG_5__SCAN_IN), .B2(keyinput_g60), .ZN(n4662) );
  AOI221_X1 U5212 ( .B1(IR_REG_24__SCAN_IN), .B2(keyinput_g79), .C1(
        keyinput_g60), .C2(IR_REG_5__SCAN_IN), .A(n4662), .ZN(n4663) );
  NAND4_X1 U5213 ( .A1(n4666), .A2(n4665), .A3(n4664), .A4(n4663), .ZN(n4667)
         );
  NOR4_X1 U5214 ( .A1(n4670), .A2(n4669), .A3(n4668), .A4(n4667), .ZN(n5013)
         );
  OAI22_X1 U5215 ( .A1(IR_REG_21__SCAN_IN), .A2(keyinput_g76), .B1(
        keyinput_g121), .B2(REG0_REG_2__SCAN_IN), .ZN(n4671) );
  AOI221_X1 U5216 ( .B1(IR_REG_21__SCAN_IN), .B2(keyinput_g76), .C1(
        REG0_REG_2__SCAN_IN), .C2(keyinput_g121), .A(n4671), .ZN(n4678) );
  OAI22_X1 U5217 ( .A1(DATAI_29_), .A2(keyinput_g2), .B1(keyinput_g12), .B2(
        DATAI_19_), .ZN(n4672) );
  AOI221_X1 U5218 ( .B1(DATAI_29_), .B2(keyinput_g2), .C1(DATAI_19_), .C2(
        keyinput_g12), .A(n4672), .ZN(n4677) );
  OAI22_X1 U5219 ( .A1(IR_REG_0__SCAN_IN), .A2(keyinput_g55), .B1(
        D_REG_26__SCAN_IN), .B2(keyinput_g113), .ZN(n4673) );
  AOI221_X1 U5220 ( .B1(IR_REG_0__SCAN_IN), .B2(keyinput_g55), .C1(
        keyinput_g113), .C2(D_REG_26__SCAN_IN), .A(n4673), .ZN(n4676) );
  OAI22_X1 U5221 ( .A1(IR_REG_3__SCAN_IN), .A2(keyinput_g58), .B1(keyinput_g94), .B2(D_REG_7__SCAN_IN), .ZN(n4674) );
  AOI221_X1 U5222 ( .B1(IR_REG_3__SCAN_IN), .B2(keyinput_g58), .C1(
        D_REG_7__SCAN_IN), .C2(keyinput_g94), .A(n4674), .ZN(n4675) );
  NAND4_X1 U5223 ( .A1(n4678), .A2(n4677), .A3(n4676), .A4(n4675), .ZN(n4804)
         );
  OAI22_X1 U5224 ( .A1(D_REG_4__SCAN_IN), .A2(keyinput_g91), .B1(keyinput_g53), 
        .B2(REG3_REG_20__SCAN_IN), .ZN(n4679) );
  AOI221_X1 U5225 ( .B1(D_REG_4__SCAN_IN), .B2(keyinput_g91), .C1(
        REG3_REG_20__SCAN_IN), .C2(keyinput_g53), .A(n4679), .ZN(n4704) );
  OAI22_X1 U5226 ( .A1(REG3_REG_10__SCAN_IN), .A2(keyinput_g37), .B1(DATAI_15_), .B2(keyinput_g16), .ZN(n4680) );
  AOI221_X1 U5227 ( .B1(REG3_REG_10__SCAN_IN), .B2(keyinput_g37), .C1(
        keyinput_g16), .C2(DATAI_15_), .A(n4680), .ZN(n4683) );
  OAI22_X1 U5228 ( .A1(IR_REG_30__SCAN_IN), .A2(keyinput_g85), .B1(
        REG0_REG_5__SCAN_IN), .B2(keyinput_g124), .ZN(n4681) );
  AOI221_X1 U5229 ( .B1(IR_REG_30__SCAN_IN), .B2(keyinput_g85), .C1(
        keyinput_g124), .C2(REG0_REG_5__SCAN_IN), .A(n4681), .ZN(n4682) );
  OAI211_X1 U5230 ( .C1(n2476), .C2(keyinput_g51), .A(n4683), .B(n4682), .ZN(
        n4684) );
  AOI21_X1 U5231 ( .B1(n2476), .B2(keyinput_g51), .A(n4684), .ZN(n4703) );
  AOI22_X1 U5232 ( .A1(DATAI_9_), .A2(keyinput_g22), .B1(IR_REG_6__SCAN_IN), 
        .B2(keyinput_g61), .ZN(n4685) );
  OAI221_X1 U5233 ( .B1(DATAI_9_), .B2(keyinput_g22), .C1(IR_REG_6__SCAN_IN), 
        .C2(keyinput_g61), .A(n4685), .ZN(n4692) );
  AOI22_X1 U5234 ( .A1(DATAI_31_), .A2(keyinput_g0), .B1(DATAI_2_), .B2(
        keyinput_g29), .ZN(n4686) );
  OAI221_X1 U5235 ( .B1(DATAI_31_), .B2(keyinput_g0), .C1(DATAI_2_), .C2(
        keyinput_g29), .A(n4686), .ZN(n4691) );
  AOI22_X1 U5236 ( .A1(REG3_REG_3__SCAN_IN), .A2(keyinput_g38), .B1(
        D_REG_19__SCAN_IN), .B2(keyinput_g106), .ZN(n4687) );
  OAI221_X1 U5237 ( .B1(REG3_REG_3__SCAN_IN), .B2(keyinput_g38), .C1(
        D_REG_19__SCAN_IN), .C2(keyinput_g106), .A(n4687), .ZN(n4690) );
  AOI22_X1 U5238 ( .A1(D_REG_31__SCAN_IN), .A2(keyinput_g118), .B1(
        IR_REG_20__SCAN_IN), .B2(keyinput_g75), .ZN(n4688) );
  OAI221_X1 U5239 ( .B1(D_REG_31__SCAN_IN), .B2(keyinput_g118), .C1(
        IR_REG_20__SCAN_IN), .C2(keyinput_g75), .A(n4688), .ZN(n4689) );
  NOR4_X1 U5240 ( .A1(n4692), .A2(n4691), .A3(n4690), .A4(n4689), .ZN(n4702)
         );
  AOI22_X1 U5241 ( .A1(DATAI_3_), .A2(keyinput_g28), .B1(DATAI_17_), .B2(
        keyinput_g14), .ZN(n4693) );
  OAI221_X1 U5242 ( .B1(DATAI_3_), .B2(keyinput_g28), .C1(DATAI_17_), .C2(
        keyinput_g14), .A(n4693), .ZN(n4700) );
  AOI22_X1 U5243 ( .A1(DATAI_22_), .A2(keyinput_g9), .B1(D_REG_30__SCAN_IN), 
        .B2(keyinput_g117), .ZN(n4694) );
  OAI221_X1 U5244 ( .B1(DATAI_22_), .B2(keyinput_g9), .C1(D_REG_30__SCAN_IN), 
        .C2(keyinput_g117), .A(n4694), .ZN(n4699) );
  AOI22_X1 U5245 ( .A1(REG0_REG_7__SCAN_IN), .A2(keyinput_g126), .B1(
        IR_REG_1__SCAN_IN), .B2(keyinput_g56), .ZN(n4695) );
  OAI221_X1 U5246 ( .B1(REG0_REG_7__SCAN_IN), .B2(keyinput_g126), .C1(
        IR_REG_1__SCAN_IN), .C2(keyinput_g56), .A(n4695), .ZN(n4698) );
  AOI22_X1 U5247 ( .A1(D_REG_5__SCAN_IN), .A2(keyinput_g92), .B1(
        IR_REG_8__SCAN_IN), .B2(keyinput_g63), .ZN(n4696) );
  OAI221_X1 U5248 ( .B1(D_REG_5__SCAN_IN), .B2(keyinput_g92), .C1(
        IR_REG_8__SCAN_IN), .C2(keyinput_g63), .A(n4696), .ZN(n4697) );
  NOR4_X1 U5249 ( .A1(n4700), .A2(n4699), .A3(n4698), .A4(n4697), .ZN(n4701)
         );
  NAND4_X1 U5250 ( .A1(n4704), .A2(n4703), .A3(n4702), .A4(n4701), .ZN(n4803)
         );
  AOI22_X1 U5251 ( .A1(REG3_REG_7__SCAN_IN), .A2(keyinput_g33), .B1(
        D_REG_17__SCAN_IN), .B2(keyinput_g104), .ZN(n4705) );
  OAI221_X1 U5252 ( .B1(REG3_REG_7__SCAN_IN), .B2(keyinput_g33), .C1(
        D_REG_17__SCAN_IN), .C2(keyinput_g104), .A(n4705), .ZN(n4713) );
  AOI22_X1 U5253 ( .A1(IR_REG_15__SCAN_IN), .A2(keyinput_g70), .B1(
        IR_REG_2__SCAN_IN), .B2(keyinput_g57), .ZN(n4706) );
  OAI221_X1 U5254 ( .B1(IR_REG_15__SCAN_IN), .B2(keyinput_g70), .C1(
        IR_REG_2__SCAN_IN), .C2(keyinput_g57), .A(n4706), .ZN(n4712) );
  AOI22_X1 U5255 ( .A1(REG3_REG_28__SCAN_IN), .A2(keyinput_g40), .B1(
        IR_REG_31__SCAN_IN), .B2(keyinput_g86), .ZN(n4707) );
  OAI221_X1 U5256 ( .B1(REG3_REG_28__SCAN_IN), .B2(keyinput_g40), .C1(
        IR_REG_31__SCAN_IN), .C2(keyinput_g86), .A(n4707), .ZN(n4711) );
  AOI22_X1 U5257 ( .A1(n4893), .A2(keyinput_g127), .B1(n4709), .B2(
        keyinput_g34), .ZN(n4708) );
  OAI221_X1 U5258 ( .B1(n4893), .B2(keyinput_g127), .C1(n4709), .C2(
        keyinput_g34), .A(n4708), .ZN(n4710) );
  NOR4_X1 U5259 ( .A1(n4713), .A2(n4712), .A3(n4711), .A4(n4710), .ZN(n4751)
         );
  INV_X1 U5260 ( .A(DATAI_26_), .ZN(n4986) );
  AOI22_X1 U5261 ( .A1(n4986), .A2(keyinput_g5), .B1(n4884), .B2(keyinput_g35), 
        .ZN(n4714) );
  OAI221_X1 U5262 ( .B1(n4986), .B2(keyinput_g5), .C1(n4884), .C2(keyinput_g35), .A(n4714), .ZN(n4724) );
  AOI22_X1 U5263 ( .A1(n4716), .A2(keyinput_g19), .B1(n2376), .B2(keyinput_g69), .ZN(n4715) );
  OAI221_X1 U5264 ( .B1(n4716), .B2(keyinput_g19), .C1(n2376), .C2(
        keyinput_g69), .A(n4715), .ZN(n4723) );
  AOI22_X1 U5265 ( .A1(n4718), .A2(keyinput_g105), .B1(n4944), .B2(
        keyinput_g107), .ZN(n4717) );
  OAI221_X1 U5266 ( .B1(n4718), .B2(keyinput_g105), .C1(n4944), .C2(
        keyinput_g107), .A(n4717), .ZN(n4722) );
  AOI22_X1 U5267 ( .A1(n4720), .A2(keyinput_g84), .B1(n4940), .B2(keyinput_g97), .ZN(n4719) );
  OAI221_X1 U5268 ( .B1(n4720), .B2(keyinput_g84), .C1(n4940), .C2(
        keyinput_g97), .A(n4719), .ZN(n4721) );
  NOR4_X1 U5269 ( .A1(n4724), .A2(n4723), .A3(n4722), .A4(n4721), .ZN(n4750)
         );
  INV_X1 U5270 ( .A(DATAI_30_), .ZN(n4726) );
  AOI22_X1 U5271 ( .A1(n4726), .A2(keyinput_g1), .B1(n2484), .B2(keyinput_g62), 
        .ZN(n4725) );
  OAI221_X1 U5272 ( .B1(n4726), .B2(keyinput_g1), .C1(n2484), .C2(keyinput_g62), .A(n4725), .ZN(n4736) );
  AOI22_X1 U5273 ( .A1(n4985), .A2(keyinput_g26), .B1(n4728), .B2(
        keyinput_g110), .ZN(n4727) );
  OAI221_X1 U5274 ( .B1(n4985), .B2(keyinput_g26), .C1(n4728), .C2(
        keyinput_g110), .A(n4727), .ZN(n4735) );
  AOI22_X1 U5275 ( .A1(n4941), .A2(keyinput_g90), .B1(keyinput_g52), .B2(n3075), .ZN(n4729) );
  OAI221_X1 U5276 ( .B1(n4941), .B2(keyinput_g90), .C1(n3075), .C2(
        keyinput_g52), .A(n4729), .ZN(n4734) );
  AOI22_X1 U5277 ( .A1(n4732), .A2(keyinput_g10), .B1(keyinput_g120), .B2(
        n4731), .ZN(n4730) );
  OAI221_X1 U5278 ( .B1(n4732), .B2(keyinput_g10), .C1(n4731), .C2(
        keyinput_g120), .A(n4730), .ZN(n4733) );
  NOR4_X1 U5279 ( .A1(n4736), .A2(n4735), .A3(n4734), .A4(n4733), .ZN(n4749)
         );
  AOI22_X1 U5280 ( .A1(n4738), .A2(keyinput_g108), .B1(keyinput_g95), .B2(
        n4912), .ZN(n4737) );
  OAI221_X1 U5281 ( .B1(n4738), .B2(keyinput_g108), .C1(n4912), .C2(
        keyinput_g95), .A(n4737), .ZN(n4747) );
  AOI22_X1 U5282 ( .A1(n4924), .A2(keyinput_g98), .B1(n4740), .B2(
        keyinput_g109), .ZN(n4739) );
  OAI221_X1 U5283 ( .B1(n4924), .B2(keyinput_g98), .C1(n4740), .C2(
        keyinput_g109), .A(n4739), .ZN(n4746) );
  AOI22_X1 U5284 ( .A1(n2639), .A2(keyinput_g45), .B1(n2583), .B2(keyinput_g72), .ZN(n4741) );
  OAI221_X1 U5285 ( .B1(n2639), .B2(keyinput_g45), .C1(n2583), .C2(
        keyinput_g72), .A(n4741), .ZN(n4745) );
  XNOR2_X1 U5286 ( .A(IR_REG_18__SCAN_IN), .B(keyinput_g73), .ZN(n4743) );
  XNOR2_X1 U5287 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput_g39), .ZN(n4742) );
  NAND2_X1 U5288 ( .A1(n4743), .A2(n4742), .ZN(n4744) );
  NOR4_X1 U5289 ( .A1(n4747), .A2(n4746), .A3(n4745), .A4(n4744), .ZN(n4748)
         );
  NAND4_X1 U5290 ( .A1(n4751), .A2(n4750), .A3(n4749), .A4(n4748), .ZN(n4802)
         );
  AOI22_X1 U5291 ( .A1(n4974), .A2(keyinput_g17), .B1(n2515), .B2(keyinput_g66), .ZN(n4752) );
  OAI221_X1 U5292 ( .B1(n4974), .B2(keyinput_g17), .C1(n2515), .C2(
        keyinput_g66), .A(n4752), .ZN(n4757) );
  XNOR2_X1 U5293 ( .A(n4753), .B(keyinput_g80), .ZN(n4756) );
  XNOR2_X1 U5294 ( .A(n4754), .B(keyinput_g112), .ZN(n4755) );
  OR3_X1 U5295 ( .A1(n4757), .A2(n4756), .A3(n4755), .ZN(n4762) );
  INV_X1 U5296 ( .A(DATAI_25_), .ZN(n4982) );
  AOI22_X1 U5297 ( .A1(n4982), .A2(keyinput_g6), .B1(keyinput_g8), .B2(n4976), 
        .ZN(n4758) );
  OAI221_X1 U5298 ( .B1(n4982), .B2(keyinput_g6), .C1(n4976), .C2(keyinput_g8), 
        .A(n4758), .ZN(n4761) );
  INV_X1 U5299 ( .A(IR_REG_23__SCAN_IN), .ZN(n4971) );
  AOI22_X1 U5300 ( .A1(n4971), .A2(keyinput_g78), .B1(keyinput_g47), .B2(n2433), .ZN(n4759) );
  OAI221_X1 U5301 ( .B1(n4971), .B2(keyinput_g78), .C1(n2433), .C2(
        keyinput_g47), .A(n4759), .ZN(n4760) );
  NOR3_X1 U5302 ( .A1(n4762), .A2(n4761), .A3(n4760), .ZN(n4800) );
  AOI22_X1 U5303 ( .A1(n4764), .A2(keyinput_g115), .B1(keyinput_g41), .B2(
        n4968), .ZN(n4763) );
  OAI221_X1 U5304 ( .B1(n4764), .B2(keyinput_g115), .C1(n4968), .C2(
        keyinput_g41), .A(n4763), .ZN(n4773) );
  INV_X1 U5305 ( .A(DATAI_0_), .ZN(n4969) );
  INV_X1 U5306 ( .A(DATAI_24_), .ZN(n4766) );
  AOI22_X1 U5307 ( .A1(n4969), .A2(keyinput_g31), .B1(keyinput_g7), .B2(n4766), 
        .ZN(n4765) );
  OAI221_X1 U5308 ( .B1(n4969), .B2(keyinput_g31), .C1(n4766), .C2(keyinput_g7), .A(n4765), .ZN(n4772) );
  AOI22_X1 U5309 ( .A1(n4923), .A2(keyinput_g102), .B1(keyinput_g125), .B2(
        n4896), .ZN(n4767) );
  OAI221_X1 U5310 ( .B1(n4923), .B2(keyinput_g102), .C1(n4896), .C2(
        keyinput_g125), .A(n4767), .ZN(n4771) );
  AOI22_X1 U5311 ( .A1(n4769), .A2(keyinput_g87), .B1(keyinput_g43), .B2(n3653), .ZN(n4768) );
  OAI221_X1 U5312 ( .B1(n4769), .B2(keyinput_g87), .C1(n3653), .C2(
        keyinput_g43), .A(n4768), .ZN(n4770) );
  NOR4_X1 U5313 ( .A1(n4773), .A2(n4772), .A3(n4771), .A4(n4770), .ZN(n4799)
         );
  INV_X1 U5314 ( .A(DATAI_4_), .ZN(n4898) );
  AOI22_X1 U5315 ( .A1(n4775), .A2(keyinput_g89), .B1(keyinput_g27), .B2(n4898), .ZN(n4774) );
  OAI221_X1 U5316 ( .B1(n4775), .B2(keyinput_g89), .C1(n4898), .C2(
        keyinput_g27), .A(n4774), .ZN(n4784) );
  XOR2_X1 U5317 ( .A(n2533), .B(keyinput_g18), .Z(n4779) );
  XNOR2_X1 U5318 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_g59), .ZN(n4778) );
  XNOR2_X1 U5319 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_g64), .ZN(n4777) );
  XNOR2_X1 U5320 ( .A(IR_REG_13__SCAN_IN), .B(keyinput_g68), .ZN(n4776) );
  NAND4_X1 U5321 ( .A1(n4779), .A2(n4778), .A3(n4777), .A4(n4776), .ZN(n4783)
         );
  XNOR2_X1 U5322 ( .A(keyinput_g54), .B(n2523), .ZN(n4782) );
  XNOR2_X1 U5323 ( .A(keyinput_g119), .B(n4780), .ZN(n4781) );
  NOR4_X1 U5324 ( .A1(n4784), .A2(n4783), .A3(n4782), .A4(n4781), .ZN(n4798)
         );
  XOR2_X1 U5325 ( .A(DATAI_7_), .B(keyinput_g24), .Z(n4788) );
  XNOR2_X1 U5326 ( .A(n4906), .B(keyinput_g83), .ZN(n4787) );
  XNOR2_X1 U5327 ( .A(n4785), .B(keyinput_g77), .ZN(n4786) );
  NOR3_X1 U5328 ( .A1(n4788), .A2(n4787), .A3(n4786), .ZN(n4791) );
  XNOR2_X1 U5329 ( .A(DATAI_10_), .B(keyinput_g21), .ZN(n4790) );
  XNOR2_X1 U5330 ( .A(IR_REG_27__SCAN_IN), .B(keyinput_g82), .ZN(n4789) );
  NAND3_X1 U5331 ( .A1(n4791), .A2(n4790), .A3(n4789), .ZN(n4796) );
  AOI22_X1 U5332 ( .A1(n4946), .A2(keyinput_g23), .B1(n4793), .B2(keyinput_g4), 
        .ZN(n4792) );
  OAI221_X1 U5333 ( .B1(n4946), .B2(keyinput_g23), .C1(n4793), .C2(keyinput_g4), .A(n4792), .ZN(n4795) );
  XNOR2_X1 U5334 ( .A(n4962), .B(keyinput_g88), .ZN(n4794) );
  NOR3_X1 U5335 ( .A1(n4796), .A2(n4795), .A3(n4794), .ZN(n4797) );
  NAND4_X1 U5336 ( .A1(n4800), .A2(n4799), .A3(n4798), .A4(n4797), .ZN(n4801)
         );
  NOR4_X1 U5337 ( .A1(n4804), .A2(n4803), .A3(n4802), .A4(n4801), .ZN(n5012)
         );
  AOI22_X1 U5338 ( .A1(REG3_REG_21__SCAN_IN), .A2(keyinput_f43), .B1(
        IR_REG_0__SCAN_IN), .B2(keyinput_f55), .ZN(n4805) );
  OAI221_X1 U5339 ( .B1(REG3_REG_21__SCAN_IN), .B2(keyinput_f43), .C1(
        IR_REG_0__SCAN_IN), .C2(keyinput_f55), .A(n4805), .ZN(n4812) );
  AOI22_X1 U5340 ( .A1(REG3_REG_4__SCAN_IN), .A2(keyinput_f50), .B1(
        REG3_REG_7__SCAN_IN), .B2(keyinput_f33), .ZN(n4806) );
  OAI221_X1 U5341 ( .B1(REG3_REG_4__SCAN_IN), .B2(keyinput_f50), .C1(
        REG3_REG_7__SCAN_IN), .C2(keyinput_f33), .A(n4806), .ZN(n4811) );
  AOI22_X1 U5342 ( .A1(REG3_REG_17__SCAN_IN), .A2(keyinput_f48), .B1(
        D_REG_30__SCAN_IN), .B2(keyinput_f117), .ZN(n4807) );
  OAI221_X1 U5343 ( .B1(REG3_REG_17__SCAN_IN), .B2(keyinput_f48), .C1(
        D_REG_30__SCAN_IN), .C2(keyinput_f117), .A(n4807), .ZN(n4810) );
  AOI22_X1 U5344 ( .A1(D_REG_19__SCAN_IN), .A2(keyinput_f106), .B1(
        D_REG_26__SCAN_IN), .B2(keyinput_f113), .ZN(n4808) );
  OAI221_X1 U5345 ( .B1(D_REG_19__SCAN_IN), .B2(keyinput_f106), .C1(
        D_REG_26__SCAN_IN), .C2(keyinput_f113), .A(n4808), .ZN(n4809) );
  NOR4_X1 U5346 ( .A1(n4812), .A2(n4811), .A3(n4810), .A4(n4809), .ZN(n5006)
         );
  OAI22_X1 U5347 ( .A1(D_REG_17__SCAN_IN), .A2(keyinput_f104), .B1(
        D_REG_9__SCAN_IN), .B2(keyinput_f96), .ZN(n4813) );
  AOI221_X1 U5348 ( .B1(D_REG_17__SCAN_IN), .B2(keyinput_f104), .C1(
        keyinput_f96), .C2(D_REG_9__SCAN_IN), .A(n4813), .ZN(n4820) );
  OAI22_X1 U5349 ( .A1(D_REG_7__SCAN_IN), .A2(keyinput_f94), .B1(
        D_REG_6__SCAN_IN), .B2(keyinput_f93), .ZN(n4814) );
  AOI221_X1 U5350 ( .B1(D_REG_7__SCAN_IN), .B2(keyinput_f94), .C1(keyinput_f93), .C2(D_REG_6__SCAN_IN), .A(n4814), .ZN(n4819) );
  OAI22_X1 U5351 ( .A1(D_REG_4__SCAN_IN), .A2(keyinput_f91), .B1(
        IR_REG_30__SCAN_IN), .B2(keyinput_f85), .ZN(n4815) );
  AOI221_X1 U5352 ( .B1(D_REG_4__SCAN_IN), .B2(keyinput_f91), .C1(keyinput_f85), .C2(IR_REG_30__SCAN_IN), .A(n4815), .ZN(n4818) );
  OAI22_X1 U5353 ( .A1(IR_REG_31__SCAN_IN), .A2(keyinput_f86), .B1(
        IR_REG_14__SCAN_IN), .B2(keyinput_f69), .ZN(n4816) );
  AOI221_X1 U5354 ( .B1(IR_REG_31__SCAN_IN), .B2(keyinput_f86), .C1(
        keyinput_f69), .C2(IR_REG_14__SCAN_IN), .A(n4816), .ZN(n4817) );
  NAND4_X1 U5355 ( .A1(n4820), .A2(n4819), .A3(n4818), .A4(n4817), .ZN(n4826)
         );
  AOI22_X1 U5356 ( .A1(DATAI_1_), .A2(keyinput_f30), .B1(DATAI_2_), .B2(
        keyinput_f29), .ZN(n4821) );
  OAI221_X1 U5357 ( .B1(DATAI_1_), .B2(keyinput_f30), .C1(DATAI_2_), .C2(
        keyinput_f29), .A(n4821), .ZN(n4825) );
  AOI22_X1 U5358 ( .A1(DATAI_24_), .A2(keyinput_f7), .B1(DATAI_28_), .B2(
        keyinput_f3), .ZN(n4822) );
  OAI221_X1 U5359 ( .B1(DATAI_24_), .B2(keyinput_f7), .C1(DATAI_28_), .C2(
        keyinput_f3), .A(n4822), .ZN(n4824) );
  XOR2_X1 U5360 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_f60), .Z(n4823) );
  NOR4_X1 U5361 ( .A1(n4826), .A2(n4825), .A3(n4824), .A4(n4823), .ZN(n4838)
         );
  OAI22_X1 U5362 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput_f34), .B1(
        keyinput_f12), .B2(DATAI_19_), .ZN(n4827) );
  AOI221_X1 U5363 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput_f34), .C1(
        DATAI_19_), .C2(keyinput_f12), .A(n4827), .ZN(n4837) );
  OAI22_X1 U5364 ( .A1(IR_REG_15__SCAN_IN), .A2(keyinput_f70), .B1(DATAI_11_), 
        .B2(keyinput_f20), .ZN(n4828) );
  AOI221_X1 U5365 ( .B1(IR_REG_15__SCAN_IN), .B2(keyinput_f70), .C1(
        keyinput_f20), .C2(DATAI_11_), .A(n4828), .ZN(n4835) );
  OAI22_X1 U5366 ( .A1(DATAI_6_), .A2(keyinput_f25), .B1(REG0_REG_4__SCAN_IN), 
        .B2(keyinput_f123), .ZN(n4829) );
  AOI221_X1 U5367 ( .B1(DATAI_6_), .B2(keyinput_f25), .C1(keyinput_f123), .C2(
        REG0_REG_4__SCAN_IN), .A(n4829), .ZN(n4834) );
  OAI22_X1 U5368 ( .A1(REG0_REG_5__SCAN_IN), .A2(keyinput_f124), .B1(
        REG0_REG_0__SCAN_IN), .B2(keyinput_f119), .ZN(n4830) );
  AOI221_X1 U5369 ( .B1(REG0_REG_5__SCAN_IN), .B2(keyinput_f124), .C1(
        keyinput_f119), .C2(REG0_REG_0__SCAN_IN), .A(n4830), .ZN(n4833) );
  OAI22_X1 U5370 ( .A1(IR_REG_8__SCAN_IN), .A2(keyinput_f63), .B1(
        keyinput_f120), .B2(REG0_REG_1__SCAN_IN), .ZN(n4831) );
  AOI221_X1 U5371 ( .B1(IR_REG_8__SCAN_IN), .B2(keyinput_f63), .C1(
        REG0_REG_1__SCAN_IN), .C2(keyinput_f120), .A(n4831), .ZN(n4832) );
  AND4_X1 U5372 ( .A1(n4835), .A2(n4834), .A3(n4833), .A4(n4832), .ZN(n4836)
         );
  AND3_X1 U5373 ( .A1(n4838), .A2(n4837), .A3(n4836), .ZN(n5005) );
  AOI22_X1 U5374 ( .A1(DATAI_13_), .A2(keyinput_f18), .B1(IR_REG_12__SCAN_IN), 
        .B2(keyinput_f67), .ZN(n4839) );
  OAI221_X1 U5375 ( .B1(DATAI_13_), .B2(keyinput_f18), .C1(IR_REG_12__SCAN_IN), 
        .C2(keyinput_f67), .A(n4839), .ZN(n4846) );
  AOI22_X1 U5376 ( .A1(REG3_REG_13__SCAN_IN), .A2(keyinput_f54), .B1(
        IR_REG_19__SCAN_IN), .B2(keyinput_f74), .ZN(n4840) );
  OAI221_X1 U5377 ( .B1(REG3_REG_13__SCAN_IN), .B2(keyinput_f54), .C1(
        IR_REG_19__SCAN_IN), .C2(keyinput_f74), .A(n4840), .ZN(n4845) );
  AOI22_X1 U5378 ( .A1(D_REG_28__SCAN_IN), .A2(keyinput_f115), .B1(
        IR_REG_18__SCAN_IN), .B2(keyinput_f73), .ZN(n4841) );
  OAI221_X1 U5379 ( .B1(D_REG_28__SCAN_IN), .B2(keyinput_f115), .C1(
        IR_REG_18__SCAN_IN), .C2(keyinput_f73), .A(n4841), .ZN(n4844) );
  AOI22_X1 U5380 ( .A1(D_REG_23__SCAN_IN), .A2(keyinput_f110), .B1(
        D_REG_22__SCAN_IN), .B2(keyinput_f109), .ZN(n4842) );
  OAI221_X1 U5381 ( .B1(D_REG_23__SCAN_IN), .B2(keyinput_f110), .C1(
        D_REG_22__SCAN_IN), .C2(keyinput_f109), .A(n4842), .ZN(n4843) );
  NOR4_X1 U5382 ( .A1(n4846), .A2(n4845), .A3(n4844), .A4(n4843), .ZN(n4876)
         );
  AOI22_X1 U5383 ( .A1(D_REG_21__SCAN_IN), .A2(keyinput_f108), .B1(
        D_REG_25__SCAN_IN), .B2(keyinput_f112), .ZN(n4847) );
  OAI221_X1 U5384 ( .B1(D_REG_21__SCAN_IN), .B2(keyinput_f108), .C1(
        D_REG_25__SCAN_IN), .C2(keyinput_f112), .A(n4847), .ZN(n4854) );
  AOI22_X1 U5385 ( .A1(D_REG_2__SCAN_IN), .A2(keyinput_f89), .B1(
        D_REG_18__SCAN_IN), .B2(keyinput_f105), .ZN(n4848) );
  OAI221_X1 U5386 ( .B1(D_REG_2__SCAN_IN), .B2(keyinput_f89), .C1(
        D_REG_18__SCAN_IN), .C2(keyinput_f105), .A(n4848), .ZN(n4853) );
  AOI22_X1 U5387 ( .A1(REG3_REG_12__SCAN_IN), .A2(keyinput_f44), .B1(
        REG3_REG_23__SCAN_IN), .B2(keyinput_f36), .ZN(n4849) );
  OAI221_X1 U5388 ( .B1(REG3_REG_12__SCAN_IN), .B2(keyinput_f44), .C1(
        REG3_REG_23__SCAN_IN), .C2(keyinput_f36), .A(n4849), .ZN(n4852) );
  AOI22_X1 U5389 ( .A1(IR_REG_27__SCAN_IN), .A2(keyinput_f82), .B1(
        IR_REG_29__SCAN_IN), .B2(keyinput_f84), .ZN(n4850) );
  OAI221_X1 U5390 ( .B1(IR_REG_27__SCAN_IN), .B2(keyinput_f82), .C1(
        IR_REG_29__SCAN_IN), .C2(keyinput_f84), .A(n4850), .ZN(n4851) );
  NOR4_X1 U5391 ( .A1(n4854), .A2(n4853), .A3(n4852), .A4(n4851), .ZN(n4875)
         );
  AOI22_X1 U5392 ( .A1(IR_REG_17__SCAN_IN), .A2(keyinput_f72), .B1(
        IR_REG_21__SCAN_IN), .B2(keyinput_f76), .ZN(n4855) );
  OAI221_X1 U5393 ( .B1(IR_REG_17__SCAN_IN), .B2(keyinput_f72), .C1(
        IR_REG_21__SCAN_IN), .C2(keyinput_f76), .A(n4855), .ZN(n4862) );
  AOI22_X1 U5394 ( .A1(DATAI_21_), .A2(keyinput_f10), .B1(IR_REG_24__SCAN_IN), 
        .B2(keyinput_f79), .ZN(n4856) );
  OAI221_X1 U5395 ( .B1(DATAI_21_), .B2(keyinput_f10), .C1(IR_REG_24__SCAN_IN), 
        .C2(keyinput_f79), .A(n4856), .ZN(n4861) );
  AOI22_X1 U5396 ( .A1(DATAI_30_), .A2(keyinput_f1), .B1(DATAI_12_), .B2(
        keyinput_f19), .ZN(n4857) );
  OAI221_X1 U5397 ( .B1(DATAI_30_), .B2(keyinput_f1), .C1(DATAI_12_), .C2(
        keyinput_f19), .A(n4857), .ZN(n4860) );
  AOI22_X1 U5398 ( .A1(D_REG_0__SCAN_IN), .A2(keyinput_f87), .B1(
        IR_REG_26__SCAN_IN), .B2(keyinput_f81), .ZN(n4858) );
  OAI221_X1 U5399 ( .B1(D_REG_0__SCAN_IN), .B2(keyinput_f87), .C1(
        IR_REG_26__SCAN_IN), .C2(keyinput_f81), .A(n4858), .ZN(n4859) );
  NOR4_X1 U5400 ( .A1(n4862), .A2(n4861), .A3(n4860), .A4(n4859), .ZN(n4874)
         );
  AOI22_X1 U5401 ( .A1(IR_REG_9__SCAN_IN), .A2(keyinput_f64), .B1(
        IR_REG_13__SCAN_IN), .B2(keyinput_f68), .ZN(n4863) );
  OAI221_X1 U5402 ( .B1(IR_REG_9__SCAN_IN), .B2(keyinput_f64), .C1(
        IR_REG_13__SCAN_IN), .C2(keyinput_f68), .A(n4863), .ZN(n4872) );
  AOI22_X1 U5403 ( .A1(DATAI_27_), .A2(keyinput_f4), .B1(U3149), .B2(
        keyinput_f32), .ZN(n4864) );
  OAI221_X1 U5404 ( .B1(DATAI_27_), .B2(keyinput_f4), .C1(U3149), .C2(
        keyinput_f32), .A(n4864), .ZN(n4871) );
  AOI22_X1 U5405 ( .A1(n3075), .A2(keyinput_f52), .B1(n3612), .B2(keyinput_f40), .ZN(n4865) );
  OAI221_X1 U5406 ( .B1(n3075), .B2(keyinput_f52), .C1(n3612), .C2(
        keyinput_f40), .A(n4865), .ZN(n4870) );
  AOI22_X1 U5407 ( .A1(n4868), .A2(keyinput_f49), .B1(keyinput_f53), .B2(n4867), .ZN(n4866) );
  OAI221_X1 U5408 ( .B1(n4868), .B2(keyinput_f49), .C1(n4867), .C2(
        keyinput_f53), .A(n4866), .ZN(n4869) );
  NOR4_X1 U5409 ( .A1(n4872), .A2(n4871), .A3(n4870), .A4(n4869), .ZN(n4873)
         );
  NAND4_X1 U5410 ( .A1(n4876), .A2(n4875), .A3(n4874), .A4(n4873), .ZN(n5003)
         );
  AOI22_X1 U5411 ( .A1(n4879), .A2(keyinput_f0), .B1(n4878), .B2(keyinput_f2), 
        .ZN(n4877) );
  OAI221_X1 U5412 ( .B1(n4879), .B2(keyinput_f0), .C1(n4878), .C2(keyinput_f2), 
        .A(n4877), .ZN(n4891) );
  INV_X1 U5413 ( .A(DATAI_22_), .ZN(n4882) );
  INV_X1 U5414 ( .A(DATAI_20_), .ZN(n4881) );
  AOI22_X1 U5415 ( .A1(n4882), .A2(keyinput_f9), .B1(keyinput_f11), .B2(n4881), 
        .ZN(n4880) );
  OAI221_X1 U5416 ( .B1(n4882), .B2(keyinput_f9), .C1(n4881), .C2(keyinput_f11), .A(n4880), .ZN(n4890) );
  AOI22_X1 U5417 ( .A1(n4885), .A2(keyinput_f38), .B1(n4884), .B2(keyinput_f35), .ZN(n4883) );
  OAI221_X1 U5418 ( .B1(n4885), .B2(keyinput_f38), .C1(n4884), .C2(
        keyinput_f35), .A(n4883), .ZN(n4889) );
  AOI22_X1 U5419 ( .A1(n4887), .A2(keyinput_f71), .B1(n2267), .B2(keyinput_f56), .ZN(n4886) );
  OAI221_X1 U5420 ( .B1(n4887), .B2(keyinput_f71), .C1(n2267), .C2(
        keyinput_f56), .A(n4886), .ZN(n4888) );
  NOR4_X1 U5421 ( .A1(n4891), .A2(n4890), .A3(n4889), .A4(n4888), .ZN(n4938)
         );
  AOI22_X1 U5422 ( .A1(n4894), .A2(keyinput_f126), .B1(n4893), .B2(
        keyinput_f127), .ZN(n4892) );
  OAI221_X1 U5423 ( .B1(n4894), .B2(keyinput_f126), .C1(n4893), .C2(
        keyinput_f127), .A(n4892), .ZN(n4904) );
  AOI22_X1 U5424 ( .A1(n4896), .A2(keyinput_f125), .B1(n2485), .B2(
        keyinput_f61), .ZN(n4895) );
  OAI221_X1 U5425 ( .B1(n4896), .B2(keyinput_f125), .C1(n2485), .C2(
        keyinput_f61), .A(n4895), .ZN(n4903) );
  AOI22_X1 U5426 ( .A1(n3117), .A2(keyinput_f122), .B1(keyinput_f27), .B2(
        n4898), .ZN(n4897) );
  OAI221_X1 U5427 ( .B1(n3117), .B2(keyinput_f122), .C1(n4898), .C2(
        keyinput_f27), .A(n4897), .ZN(n4902) );
  XOR2_X1 U5428 ( .A(n2433), .B(keyinput_f47), .Z(n4900) );
  XNOR2_X1 U5429 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_f58), .ZN(n4899) );
  NAND2_X1 U5430 ( .A1(n4900), .A2(n4899), .ZN(n4901) );
  NOR4_X1 U5431 ( .A1(n4904), .A2(n4903), .A3(n4902), .A4(n4901), .ZN(n4937)
         );
  AOI22_X1 U5432 ( .A1(n2476), .A2(keyinput_f51), .B1(n2515), .B2(keyinput_f66), .ZN(n4905) );
  OAI221_X1 U5433 ( .B1(n2476), .B2(keyinput_f51), .C1(n2515), .C2(
        keyinput_f66), .A(n4905), .ZN(n4910) );
  XNOR2_X1 U5434 ( .A(n4906), .B(keyinput_f83), .ZN(n4909) );
  XNOR2_X1 U5435 ( .A(n4907), .B(keyinput_f116), .ZN(n4908) );
  OR3_X1 U5436 ( .A1(n4910), .A2(n4909), .A3(n4908), .ZN(n4918) );
  AOI22_X1 U5437 ( .A1(n4913), .A2(keyinput_f101), .B1(keyinput_f95), .B2(
        n4912), .ZN(n4911) );
  OAI221_X1 U5438 ( .B1(n4913), .B2(keyinput_f101), .C1(n4912), .C2(
        keyinput_f95), .A(n4911), .ZN(n4917) );
  AOI22_X1 U5439 ( .A1(n2484), .A2(keyinput_f62), .B1(keyinput_f22), .B2(n4915), .ZN(n4914) );
  OAI221_X1 U5440 ( .B1(n2484), .B2(keyinput_f62), .C1(n4915), .C2(
        keyinput_f22), .A(n4914), .ZN(n4916) );
  NOR3_X1 U5441 ( .A1(n4918), .A2(n4917), .A3(n4916), .ZN(n4936) );
  AOI22_X1 U5442 ( .A1(n4921), .A2(keyinput_f100), .B1(keyinput_f111), .B2(
        n4920), .ZN(n4919) );
  OAI221_X1 U5443 ( .B1(n4921), .B2(keyinput_f100), .C1(n4920), .C2(
        keyinput_f111), .A(n4919), .ZN(n4934) );
  AOI22_X1 U5444 ( .A1(n4924), .A2(keyinput_f98), .B1(keyinput_f102), .B2(
        n4923), .ZN(n4922) );
  OAI221_X1 U5445 ( .B1(n4924), .B2(keyinput_f98), .C1(n4923), .C2(
        keyinput_f102), .A(n4922), .ZN(n4933) );
  AOI22_X1 U5446 ( .A1(n4927), .A2(keyinput_f99), .B1(keyinput_f118), .B2(
        n4926), .ZN(n4925) );
  OAI221_X1 U5447 ( .B1(n4927), .B2(keyinput_f99), .C1(n4926), .C2(
        keyinput_f118), .A(n4925), .ZN(n4932) );
  AOI22_X1 U5448 ( .A1(n4930), .A2(keyinput_f92), .B1(keyinput_f114), .B2(
        n4929), .ZN(n4928) );
  OAI221_X1 U5449 ( .B1(n4930), .B2(keyinput_f92), .C1(n4929), .C2(
        keyinput_f114), .A(n4928), .ZN(n4931) );
  NOR4_X1 U5450 ( .A1(n4934), .A2(n4933), .A3(n4932), .A4(n4931), .ZN(n4935)
         );
  NAND4_X1 U5451 ( .A1(n4938), .A2(n4937), .A3(n4936), .A4(n4935), .ZN(n5002)
         );
  AOI22_X1 U5452 ( .A1(n4941), .A2(keyinput_f90), .B1(keyinput_f97), .B2(n4940), .ZN(n4939) );
  OAI221_X1 U5453 ( .B1(n4941), .B2(keyinput_f90), .C1(n4940), .C2(
        keyinput_f97), .A(n4939), .ZN(n4952) );
  AOI22_X1 U5454 ( .A1(n4944), .A2(keyinput_f107), .B1(keyinput_f103), .B2(
        n4943), .ZN(n4942) );
  OAI221_X1 U5455 ( .B1(n4944), .B2(keyinput_f107), .C1(n4943), .C2(
        keyinput_f103), .A(n4942), .ZN(n4951) );
  AOI22_X1 U5456 ( .A1(n2639), .A2(keyinput_f45), .B1(keyinput_f23), .B2(n4946), .ZN(n4945) );
  OAI221_X1 U5457 ( .B1(n2639), .B2(keyinput_f45), .C1(n4946), .C2(
        keyinput_f23), .A(n4945), .ZN(n4950) );
  AOI22_X1 U5458 ( .A1(n2683), .A2(keyinput_f75), .B1(keyinput_f21), .B2(n4948), .ZN(n4947) );
  OAI221_X1 U5459 ( .B1(n2683), .B2(keyinput_f75), .C1(n4948), .C2(
        keyinput_f21), .A(n4947), .ZN(n4949) );
  NOR4_X1 U5460 ( .A1(n4952), .A2(n4951), .A3(n4950), .A4(n4949), .ZN(n5000)
         );
  INV_X1 U5461 ( .A(DATAI_3_), .ZN(n4955) );
  AOI22_X1 U5462 ( .A1(n4955), .A2(keyinput_f28), .B1(n4954), .B2(keyinput_f14), .ZN(n4953) );
  OAI221_X1 U5463 ( .B1(n4955), .B2(keyinput_f28), .C1(n4954), .C2(
        keyinput_f14), .A(n4953), .ZN(n4966) );
  AOI22_X1 U5464 ( .A1(n4958), .A2(keyinput_f15), .B1(keyinput_f24), .B2(n4957), .ZN(n4956) );
  OAI221_X1 U5465 ( .B1(n4958), .B2(keyinput_f15), .C1(n4957), .C2(
        keyinput_f24), .A(n4956), .ZN(n4965) );
  XNOR2_X1 U5466 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_f59), .ZN(n4961) );
  XNOR2_X1 U5467 ( .A(IR_REG_22__SCAN_IN), .B(keyinput_f77), .ZN(n4960) );
  XNOR2_X1 U5468 ( .A(DATAI_18_), .B(keyinput_f13), .ZN(n4959) );
  NAND3_X1 U5469 ( .A1(n4961), .A2(n4960), .A3(n4959), .ZN(n4964) );
  XNOR2_X1 U5470 ( .A(n4962), .B(keyinput_f88), .ZN(n4963) );
  NOR4_X1 U5471 ( .A1(n4966), .A2(n4965), .A3(n4964), .A4(n4963), .ZN(n4999)
         );
  AOI22_X1 U5472 ( .A1(n4969), .A2(keyinput_f31), .B1(n4968), .B2(keyinput_f41), .ZN(n4967) );
  OAI221_X1 U5473 ( .B1(n4969), .B2(keyinput_f31), .C1(n4968), .C2(
        keyinput_f41), .A(n4967), .ZN(n4980) );
  AOI22_X1 U5474 ( .A1(n2369), .A2(keyinput_f57), .B1(n4971), .B2(keyinput_f78), .ZN(n4970) );
  OAI221_X1 U5475 ( .B1(n2369), .B2(keyinput_f57), .C1(n4971), .C2(
        keyinput_f78), .A(n4970), .ZN(n4979) );
  AOI22_X1 U5476 ( .A1(n4974), .A2(keyinput_f17), .B1(n4973), .B2(keyinput_f37), .ZN(n4972) );
  OAI221_X1 U5477 ( .B1(n4974), .B2(keyinput_f17), .C1(n4973), .C2(
        keyinput_f37), .A(n4972), .ZN(n4978) );
  AOI22_X1 U5478 ( .A1(n4976), .A2(keyinput_f8), .B1(keyinput_f121), .B2(n4579), .ZN(n4975) );
  OAI221_X1 U5479 ( .B1(n4976), .B2(keyinput_f8), .C1(n4579), .C2(
        keyinput_f121), .A(n4975), .ZN(n4977) );
  NOR4_X1 U5480 ( .A1(n4980), .A2(n4979), .A3(n4978), .A4(n4977), .ZN(n4998)
         );
  AOI22_X1 U5481 ( .A1(n4983), .A2(keyinput_f16), .B1(n4982), .B2(keyinput_f6), 
        .ZN(n4981) );
  OAI221_X1 U5482 ( .B1(n4983), .B2(keyinput_f16), .C1(n4982), .C2(keyinput_f6), .A(n4981), .ZN(n4996) );
  AOI22_X1 U5483 ( .A1(n4986), .A2(keyinput_f5), .B1(n4985), .B2(keyinput_f26), 
        .ZN(n4984) );
  OAI221_X1 U5484 ( .B1(n4986), .B2(keyinput_f5), .C1(n4985), .C2(keyinput_f26), .A(n4984), .ZN(n4995) );
  INV_X1 U5485 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4989) );
  AOI22_X1 U5486 ( .A1(n4989), .A2(keyinput_f39), .B1(keyinput_f46), .B2(n4988), .ZN(n4987) );
  OAI221_X1 U5487 ( .B1(n4989), .B2(keyinput_f39), .C1(n4988), .C2(
        keyinput_f46), .A(n4987), .ZN(n4994) );
  INV_X1 U5488 ( .A(IR_REG_10__SCAN_IN), .ZN(n4990) );
  XOR2_X1 U5489 ( .A(n4990), .B(keyinput_f65), .Z(n4992) );
  XNOR2_X1 U5490 ( .A(IR_REG_25__SCAN_IN), .B(keyinput_f80), .ZN(n4991) );
  NAND2_X1 U5491 ( .A1(n4992), .A2(n4991), .ZN(n4993) );
  NOR4_X1 U5492 ( .A1(n4996), .A2(n4995), .A3(n4994), .A4(n4993), .ZN(n4997)
         );
  NAND4_X1 U5493 ( .A1(n5000), .A2(n4999), .A3(n4998), .A4(n4997), .ZN(n5001)
         );
  NOR3_X1 U5494 ( .A1(n5003), .A2(n5002), .A3(n5001), .ZN(n5004) );
  NAND3_X1 U5495 ( .A1(n5006), .A2(n5005), .A3(n5004), .ZN(n5008) );
  AOI21_X1 U5496 ( .B1(keyinput_f42), .B2(n5008), .A(REG3_REG_1__SCAN_IN), 
        .ZN(n5010) );
  INV_X1 U5497 ( .A(keyinput_f42), .ZN(n5007) );
  AOI21_X1 U5498 ( .B1(n5008), .B2(n5007), .A(keyinput_g42), .ZN(n5009) );
  AOI22_X1 U5499 ( .A1(keyinput_g42), .A2(n5010), .B1(REG3_REG_1__SCAN_IN), 
        .B2(n5009), .ZN(n5011) );
  AOI21_X1 U5500 ( .B1(n5013), .B2(n5012), .A(n5011), .ZN(n5016) );
  AOI22_X1 U5501 ( .A1(STATE_REG_SCAN_IN), .A2(IR_REG_0__SCAN_IN), .B1(
        DATAI_0_), .B2(U3149), .ZN(n5015) );
  XNOR2_X1 U5502 ( .A(n5016), .B(n5015), .ZN(U3352) );
  CLKBUF_X1 U2474 ( .A(n2418), .Z(n2672) );
  CLKBUF_X1 U2510 ( .A(n4341), .Z(n2221) );
endmodule

