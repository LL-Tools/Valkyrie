

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325;

  INV_X1 U4893 ( .A(n9560), .ZN(n9533) );
  INV_X1 U4894 ( .A(n5984), .ZN(n6301) );
  INV_X1 U4895 ( .A(n5968), .ZN(n6395) );
  NAND2_X1 U4896 ( .A1(n5882), .A2(n5881), .ZN(n8865) );
  INV_X1 U4897 ( .A(n5596), .ZN(n6457) );
  INV_X1 U4898 ( .A(n7330), .ZN(n6460) );
  AND2_X1 U4899 ( .A1(n5899), .A2(n9013), .ZN(n5902) );
  CLKBUF_X2 U4900 ( .A(n9701), .Z(n4390) );
  INV_X1 U4901 ( .A(n5901), .ZN(n6569) );
  INV_X1 U4902 ( .A(n4395), .ZN(n6227) );
  AOI21_X1 U4903 ( .B1(n8299), .B2(n8298), .A(n6277), .ZN(n6292) );
  INV_X1 U4904 ( .A(n8142), .ZN(n6812) );
  INV_X1 U4905 ( .A(n8233), .ZN(n5900) );
  INV_X1 U4906 ( .A(n8087), .ZN(n6322) );
  INV_X1 U4907 ( .A(n5944), .ZN(n6556) );
  INV_X1 U4908 ( .A(n8865), .ZN(n8734) );
  INV_X1 U4909 ( .A(n4990), .ZN(n6445) );
  AND2_X2 U4910 ( .A1(n8203), .A2(n4944), .ZN(n5009) );
  NAND2_X2 U4911 ( .A1(n5478), .A2(n7861), .ZN(n4958) );
  AOI21_X1 U4912 ( .B1(n5484), .B2(n9637), .A(n5483), .ZN(n9515) );
  INV_X1 U4913 ( .A(n5598), .ZN(n10053) );
  OR2_X1 U4914 ( .A1(n4949), .A2(n5187), .ZN(n4951) );
  BUF_X1 U4915 ( .A(n4980), .Z(n4391) );
  AOI21_X1 U4916 ( .B1(n6298), .B2(n6297), .A(n8256), .ZN(n8321) );
  AND3_X2 U4917 ( .A1(n5937), .A2(n5936), .A3(n5935), .ZN(n6894) );
  INV_X1 U4918 ( .A(n5010), .ZN(n4964) );
  XNOR2_X1 U4920 ( .A(n6357), .B(n6356), .ZN(n7956) );
  INV_X1 U4921 ( .A(n4945), .ZN(n8203) );
  NAND3_X1 U4922 ( .A1(n4963), .A2(n4962), .A3(n4961), .ZN(n5598) );
  NAND2_X2 U4923 ( .A1(n7170), .A2(n7169), .ZN(n7412) );
  AOI211_X2 U4924 ( .C1(n10006), .C2(n9736), .A(n9538), .B(n9537), .ZN(n9539)
         );
  NOR2_X4 U4925 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5933) );
  INV_X1 U4926 ( .A(n4980), .ZN(n4389) );
  XNOR2_X2 U4927 ( .A(n4940), .B(P1_IR_REG_30__SCAN_IN), .ZN(n4944) );
  NAND2_X4 U4928 ( .A1(n4777), .A2(n6508), .ZN(n5984) );
  XNOR2_X2 U4929 ( .A(n5867), .B(n5866), .ZN(n8223) );
  NAND2_X1 U4930 ( .A1(n4803), .A2(n4802), .ZN(n8248) );
  NAND2_X1 U4931 ( .A1(n7618), .A2(n7619), .ZN(n7617) );
  NAND2_X1 U4932 ( .A1(n5350), .A2(n5349), .ZN(n9618) );
  NAND2_X1 U4933 ( .A1(n7972), .A2(n8014), .ZN(n8154) );
  NAND2_X1 U4934 ( .A1(n7341), .A2(n10129), .ZN(n8014) );
  NAND2_X1 U4935 ( .A1(n7310), .A2(n9373), .ZN(n9172) );
  INV_X2 U4936 ( .A(n5592), .ZN(n6462) );
  NAND2_X1 U4937 ( .A1(n5096), .A2(n5095), .ZN(n5106) );
  AND2_X1 U4938 ( .A1(n6497), .A2(n10191), .ZN(n6896) );
  NAND4_X1 U4939 ( .A1(n4996), .A2(n4995), .A3(n4994), .A4(n4993), .ZN(n9469)
         );
  INV_X1 U4940 ( .A(n6998), .ZN(n5607) );
  NAND4_X2 U4941 ( .A1(n5932), .A2(n5931), .A3(n5930), .A4(n5929), .ZN(n6491)
         );
  NAND4_X2 U4942 ( .A1(n5958), .A2(n5957), .A3(n5956), .A4(n5955), .ZN(n10111)
         );
  OR2_X1 U4943 ( .A1(n4398), .A2(n5918), .ZN(n5922) );
  OR2_X1 U4944 ( .A1(n5954), .A2(n6681), .ZN(n5929) );
  CLKBUF_X3 U4945 ( .A(n5954), .Z(n4398) );
  CLKBUF_X3 U4946 ( .A(n5954), .Z(n4397) );
  NAND2_X1 U4947 ( .A1(n9022), .A2(n8233), .ZN(n5953) );
  BUF_X1 U4948 ( .A(n5943), .Z(n4395) );
  NAND2_X2 U4949 ( .A1(n5900), .A2(n9022), .ZN(n5968) );
  NAND2_X1 U4950 ( .A1(n5944), .A2(n5868), .ZN(n5943) );
  INV_X2 U4951 ( .A(n5902), .ZN(n9022) );
  INV_X8 U4952 ( .A(n4825), .ZN(n5868) );
  INV_X1 U4953 ( .A(n4980), .ZN(n4825) );
  OAI21_X1 U4954 ( .B1(n9447), .B2(n9446), .A(n9445), .ZN(n9455) );
  AND2_X1 U4955 ( .A1(n4702), .A2(n4703), .ZN(n6482) );
  OR2_X1 U4956 ( .A1(n9407), .A2(n9443), .ZN(n9446) );
  OAI21_X1 U4957 ( .B1(n9406), .B2(n9332), .A(n9331), .ZN(n4568) );
  AOI21_X1 U4958 ( .B1(n8140), .B2(n8139), .A(n8138), .ZN(n4744) );
  NAND2_X2 U4959 ( .A1(n5748), .A2(n9133), .ZN(n9034) );
  OAI21_X1 U4960 ( .B1(n4581), .B2(n4580), .A(n9396), .ZN(n9282) );
  AOI21_X1 U4961 ( .B1(n8229), .B2(n10156), .A(n8228), .ZN(n8908) );
  AOI21_X1 U4962 ( .B1(n9277), .B2(n6439), .A(n4416), .ZN(n4580) );
  NAND2_X1 U4963 ( .A1(n4834), .A2(n4833), .ZN(n8740) );
  AND2_X1 U4964 ( .A1(n8759), .A2(n8758), .ZN(n8761) );
  AOI21_X1 U4965 ( .B1(n4750), .B2(n8725), .A(n4749), .ZN(n4748) );
  XNOR2_X1 U4966 ( .A(n6276), .B(n6274), .ZN(n8299) );
  NAND2_X1 U4967 ( .A1(n8248), .A2(n6265), .ZN(n6276) );
  NAND2_X1 U4968 ( .A1(n8113), .A2(n8112), .ZN(n8823) );
  NAND2_X1 U4969 ( .A1(n8209), .A2(n8208), .ZN(n8806) );
  OR2_X1 U4970 ( .A1(n9563), .A2(n9545), .ZN(n9541) );
  NAND2_X1 U4971 ( .A1(n4767), .A2(n4765), .ZN(n8840) );
  NAND2_X1 U4972 ( .A1(n5870), .A2(n5869), .ZN(n8724) );
  NAND2_X1 U4973 ( .A1(n5400), .A2(n5399), .ZN(n9563) );
  NAND2_X1 U4974 ( .A1(n5911), .A2(n5910), .ZN(n8935) );
  NAND2_X1 U4975 ( .A1(n5381), .A2(n5380), .ZN(n9756) );
  XNOR2_X1 U4976 ( .A(n5412), .B(n5411), .ZN(n7730) );
  NOR2_X1 U4977 ( .A1(n9653), .A2(n9772), .ZN(n9639) );
  NAND2_X1 U4978 ( .A1(n4680), .A2(n5392), .ZN(n5412) );
  AND2_X1 U4979 ( .A1(n9296), .A2(n9608), .ZN(n9243) );
  OR2_X1 U4980 ( .A1(n5394), .A2(n5393), .ZN(n4680) );
  NAND2_X1 U4981 ( .A1(n7362), .A2(n7363), .ZN(n4781) );
  NAND2_X1 U4982 ( .A1(n4764), .A2(n4762), .ZN(n7878) );
  NAND2_X1 U4983 ( .A1(n4879), .A2(n4885), .ZN(n7453) );
  NAND2_X1 U4984 ( .A1(n5333), .A2(n5332), .ZN(n9772) );
  XNOR2_X1 U4985 ( .A(n5377), .B(n5376), .ZN(n7502) );
  OAI21_X1 U4986 ( .B1(n5362), .B2(n5361), .A(n5360), .ZN(n5377) );
  OR2_X1 U4987 ( .A1(n5513), .A2(n5512), .ZN(n7758) );
  NAND2_X1 U4988 ( .A1(n5322), .A2(n5321), .ZN(n9657) );
  OAI21_X1 U4989 ( .B1(n5340), .B2(n4642), .A(n5344), .ZN(n5362) );
  NAND2_X1 U4990 ( .A1(n7190), .A2(n7189), .ZN(n7188) );
  XNOR2_X1 U4991 ( .A(n5630), .B(n5631), .ZN(n7190) );
  NAND2_X1 U4992 ( .A1(n4685), .A2(n5298), .ZN(n5316) );
  AND2_X1 U4993 ( .A1(n8024), .A2(n8026), .ZN(n10154) );
  OAI21_X1 U4994 ( .B1(n5279), .B2(n5278), .A(n5277), .ZN(n5296) );
  NAND2_X1 U4995 ( .A1(n5083), .A2(n9310), .ZN(n7325) );
  NAND2_X1 U4996 ( .A1(n8022), .A2(n8020), .ZN(n8156) );
  NAND2_X1 U4997 ( .A1(n6151), .A2(n6150), .ZN(n8989) );
  NAND2_X1 U4998 ( .A1(n6118), .A2(n6117), .ZN(n10162) );
  OR2_X1 U4999 ( .A1(n7562), .A2(n7561), .ZN(n8022) );
  NAND2_X1 U5000 ( .A1(n5168), .A2(n5167), .ZN(n9058) );
  NAND2_X1 U5001 ( .A1(n4645), .A2(n4643), .ZN(n5279) );
  NAND2_X1 U5002 ( .A1(n6136), .A2(n6135), .ZN(n8033) );
  NAND2_X1 U5003 ( .A1(n6103), .A2(n6102), .ZN(n7562) );
  OAI21_X1 U5004 ( .B1(n7234), .B2(n9377), .A(n9419), .ZN(n7327) );
  AND2_X1 U5005 ( .A1(n8006), .A2(n8007), .ZN(n8150) );
  NAND2_X1 U5006 ( .A1(n5202), .A2(n5201), .ZN(n5220) );
  NOR2_X2 U5007 ( .A1(n7144), .A2(n10248), .ZN(n6504) );
  INV_X2 U5008 ( .A(n8881), .ZN(n4392) );
  AND2_X1 U5009 ( .A1(n7996), .A2(n7999), .ZN(n8893) );
  INV_X2 U5010 ( .A(n10260), .ZN(n4393) );
  AND2_X2 U5011 ( .A1(n7133), .A2(n10008), .ZN(n10024) );
  CLKBUF_X3 U5012 ( .A(n5596), .Z(n6463) );
  AND2_X1 U5013 ( .A1(n9415), .A2(n9414), .ZN(n9302) );
  NAND2_X1 U5014 ( .A1(n4590), .A2(n7199), .ZN(n7198) );
  INV_X1 U5015 ( .A(n6912), .ZN(n6902) );
  AND4_X1 U5016 ( .A1(n6108), .A2(n6107), .A3(n6106), .A4(n6105), .ZN(n7561)
         );
  AND4_X1 U5017 ( .A1(n6073), .A2(n6072), .A3(n6071), .A4(n6070), .ZN(n10129)
         );
  AND4_X1 U5018 ( .A1(n6059), .A2(n6058), .A3(n6057), .A4(n6056), .ZN(n7268)
         );
  AND4_X1 U5019 ( .A1(n6024), .A2(n6023), .A3(n6022), .A4(n6021), .ZN(n7102)
         );
  NAND4_X1 U5020 ( .A1(n5972), .A2(n5971), .A3(n5970), .A4(n5969), .ZN(n8337)
         );
  AND3_X1 U5021 ( .A1(n5008), .A2(n5007), .A3(n5006), .ZN(n10057) );
  AND4_X1 U5022 ( .A1(n6043), .A2(n6042), .A3(n6041), .A4(n6040), .ZN(n7168)
         );
  NAND4_X1 U5023 ( .A1(n5992), .A2(n5991), .A3(n5990), .A4(n5989), .ZN(n10139)
         );
  NAND4_X2 U5024 ( .A1(n5923), .A2(n5922), .A3(n5921), .A4(n5920), .ZN(n6497)
         );
  NOR2_X1 U5025 ( .A1(n4398), .A2(n10151), .ZN(n6002) );
  INV_X1 U5026 ( .A(n8098), .ZN(n8097) );
  OR2_X1 U5027 ( .A1(n6428), .A2(n6531), .ZN(n4962) );
  NAND2_X1 U5028 ( .A1(n4958), .A2(n5868), .ZN(n4986) );
  NAND2_X1 U5029 ( .A1(n8145), .A2(n8171), .ZN(n6508) );
  CLKBUF_X2 U5030 ( .A(n5943), .Z(n4394) );
  XNOR2_X1 U5031 ( .A(n5875), .B(n5877), .ZN(n8104) );
  XNOR2_X1 U5032 ( .A(n4510), .B(n5305), .ZN(n9701) );
  NAND2_X1 U5033 ( .A1(n4632), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4631) );
  OR2_X1 U5034 ( .A1(n6051), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6081) );
  OAI21_X1 U5035 ( .B1(n5876), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6357) );
  XNOR2_X1 U5036 ( .A(n5865), .B(n5864), .ZN(n6394) );
  AND4_X1 U5037 ( .A1(n4919), .A2(n4436), .A3(n4950), .A4(n5101), .ZN(n4941)
         );
  NAND2_X1 U5038 ( .A1(n5898), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4507) );
  INV_X1 U5039 ( .A(n5112), .ZN(n5101) );
  NAND2_X2 U5040 ( .A1(n5868), .A2(P2_U3152), .ZN(n9018) );
  INV_X2 U5041 ( .A(n9016), .ZN(n9021) );
  NAND2_X1 U5042 ( .A1(n4775), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5867) );
  AND3_X1 U5043 ( .A1(n4856), .A2(n4858), .A3(n5864), .ZN(n5894) );
  NOR2_X1 U5044 ( .A1(n4934), .A2(n4933), .ZN(n5303) );
  NAND2_X1 U5045 ( .A1(n4430), .A2(n4876), .ZN(n5112) );
  NOR2_X1 U5046 ( .A1(n6352), .A2(n4857), .ZN(n4856) );
  NAND2_X2 U5047 ( .A1(n4827), .A2(n4826), .ZN(n4980) );
  NAND4_X1 U5048 ( .A1(n4410), .A2(n5861), .A3(n4470), .A4(n4469), .ZN(n6352)
         );
  AND4_X1 U5049 ( .A1(n5857), .A2(n5976), .A3(n5856), .A4(n6032), .ZN(n5858)
         );
  AND2_X1 U5050 ( .A1(n5862), .A2(n6361), .ZN(n5863) );
  NOR2_X1 U5051 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5854) );
  NOR2_X1 U5052 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5853) );
  NOR2_X1 U5053 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n4470) );
  NOR2_X1 U5054 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5852) );
  INV_X4 U5055 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NOR2_X1 U5056 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5857) );
  INV_X1 U5057 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5280) );
  INV_X1 U5058 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5872) );
  INV_X1 U5059 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5976) );
  NOR2_X1 U5060 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5861) );
  NOR2_X1 U5061 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n4469) );
  INV_X1 U5062 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4931) );
  INV_X1 U5063 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6361) );
  NOR2_X1 U5064 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4932) );
  INV_X1 U5065 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6032) );
  INV_X2 U5066 ( .A(n5871), .ZN(n4858) );
  OAI21_X2 U5067 ( .B1(n5106), .B2(n5105), .A(n5107), .ZN(n5124) );
  OAI222_X1 U5068 ( .A1(P2_U3152), .A2(n8223), .B1(n9021), .B2(n7884), .C1(
        n7883), .C2(n9018), .ZN(P2_U3331) );
  OAI21_X2 U5069 ( .B1(n5106), .B2(n4870), .A(n4867), .ZN(n5143) );
  NAND2_X4 U5070 ( .A1(n4945), .A2(n9876), .ZN(n5210) );
  XNOR2_X2 U5071 ( .A(n4951), .B(n4950), .ZN(n5478) );
  NAND2_X1 U5072 ( .A1(n5900), .A2(n9022), .ZN(n4396) );
  XNOR2_X2 U5073 ( .A(n4507), .B(n4506), .ZN(n8233) );
  NAND2_X1 U5074 ( .A1(n5183), .A2(n5182), .ZN(n5201) );
  NAND2_X1 U5075 ( .A1(n4478), .A2(n4477), .ZN(n4476) );
  NAND2_X1 U5076 ( .A1(n7982), .A2(n8098), .ZN(n4478) );
  NAND2_X1 U5077 ( .A1(n7983), .A2(n8097), .ZN(n4477) );
  AOI21_X1 U5078 ( .B1(n4487), .B2(n8119), .A(n8098), .ZN(n4486) );
  OAI21_X1 U5079 ( .B1(n8057), .B2(n4488), .A(n8056), .ZN(n4487) );
  OR2_X1 U5080 ( .A1(n8121), .A2(n8055), .ZN(n4488) );
  NOR2_X1 U5081 ( .A1(n4484), .A2(n4483), .ZN(n4482) );
  NOR2_X1 U5082 ( .A1(n8163), .A2(n4400), .ZN(n4484) );
  INV_X1 U5083 ( .A(n8067), .ZN(n4483) );
  AOI21_X1 U5084 ( .B1(n4871), .B2(n4869), .A(n4868), .ZN(n4867) );
  INV_X1 U5085 ( .A(n4871), .ZN(n4870) );
  INV_X1 U5086 ( .A(n5107), .ZN(n4869) );
  NAND2_X1 U5087 ( .A1(n5863), .A2(n5866), .ZN(n4857) );
  INV_X1 U5088 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5864) );
  NAND2_X2 U5089 ( .A1(n5839), .A2(n5582), .ZN(n5649) );
  AOI21_X1 U5090 ( .B1(n4647), .B2(n4650), .A(n4644), .ZN(n4643) );
  INV_X1 U5091 ( .A(n5262), .ZN(n4644) );
  AND2_X1 U5092 ( .A1(n9224), .A2(n9223), .ZN(n4579) );
  OR2_X1 U5093 ( .A1(n8061), .A2(n8097), .ZN(n4489) );
  AOI21_X1 U5094 ( .B1(n4565), .B2(n9240), .A(n9323), .ZN(n4561) );
  NAND2_X1 U5095 ( .A1(n4480), .A2(n4479), .ZN(n8070) );
  NAND2_X1 U5096 ( .A1(n7956), .A2(n7955), .ZN(n8098) );
  OR2_X1 U5097 ( .A1(n8134), .A2(n8090), .ZN(n8137) );
  OR2_X1 U5098 ( .A1(n8390), .A2(n8095), .ZN(n8099) );
  NOR2_X1 U5099 ( .A1(n8958), .A2(n8966), .ZN(n4544) );
  OR2_X1 U5100 ( .A1(n8975), .A2(n7963), .ZN(n8107) );
  OR2_X1 U5101 ( .A1(n8984), .A2(n7800), .ZN(n7968) );
  OR2_X1 U5102 ( .A1(n8989), .A2(n7711), .ZN(n8030) );
  INV_X1 U5103 ( .A(n8002), .ZN(n4758) );
  OR2_X1 U5104 ( .A1(n8905), .A2(n8682), .ZN(n8084) );
  NAND2_X1 U5105 ( .A1(n5646), .A2(n7455), .ZN(n4898) );
  INV_X1 U5106 ( .A(n9050), .ZN(n5684) );
  OR2_X1 U5107 ( .A1(n6464), .A2(n9534), .ZN(n9391) );
  AND2_X1 U5108 ( .A1(n9431), .A2(n9385), .ZN(n4699) );
  AND2_X1 U5109 ( .A1(n4442), .A2(n4604), .ZN(n4602) );
  INV_X1 U5110 ( .A(n5151), .ZN(n5149) );
  NAND2_X1 U5111 ( .A1(n7325), .A2(n4690), .ZN(n10012) );
  NOR2_X1 U5112 ( .A1(n4692), .A2(n4691), .ZN(n4690) );
  INV_X1 U5113 ( .A(n9192), .ZN(n4691) );
  INV_X1 U5114 ( .A(n9187), .ZN(n4692) );
  OR2_X1 U5115 ( .A1(n9398), .A2(n5539), .ZN(n5839) );
  NAND2_X1 U5116 ( .A1(n4667), .A2(n4665), .ZN(n6414) );
  AOI21_X1 U5117 ( .B1(n4669), .B2(n4671), .A(n4666), .ZN(n4665) );
  INV_X1 U5118 ( .A(n6411), .ZN(n4666) );
  XNOR2_X1 U5119 ( .A(n6414), .B(n6412), .ZN(n6422) );
  NAND2_X1 U5120 ( .A1(n5431), .A2(n5430), .ZN(n5444) );
  AOI21_X1 U5121 ( .B1(n4681), .B2(n4678), .A(n4677), .ZN(n4676) );
  AND2_X1 U5122 ( .A1(n5430), .A2(n5416), .ZN(n5428) );
  NAND2_X1 U5123 ( .A1(n5379), .A2(n5378), .ZN(n5394) );
  NAND2_X1 U5124 ( .A1(n5331), .A2(n5330), .ZN(n5340) );
  AND2_X1 U5125 ( .A1(n5262), .A2(n5246), .ZN(n5260) );
  NAND2_X1 U5126 ( .A1(n5240), .A2(n5224), .ZN(n5241) );
  NAND2_X1 U5127 ( .A1(n4658), .A2(n4656), .ZN(n5202) );
  AOI21_X1 U5128 ( .B1(n4659), .B2(n4407), .A(n4657), .ZN(n4656) );
  AND2_X1 U5129 ( .A1(n5201), .A2(n5185), .ZN(n5199) );
  NOR2_X1 U5130 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4977) );
  AOI21_X1 U5131 ( .B1(n4434), .B2(n4823), .A(n4821), .ZN(n4820) );
  INV_X1 U5132 ( .A(n6351), .ZN(n4821) );
  NAND2_X1 U5133 ( .A1(n6332), .A2(n8191), .ZN(n4823) );
  NOR2_X1 U5134 ( .A1(n8685), .A2(n8920), .ZN(n4546) );
  AND2_X1 U5135 ( .A1(n4549), .A2(n4548), .ZN(n4547) );
  NOR2_X1 U5136 ( .A1(n8685), .A2(n8920), .ZN(n4549) );
  NOR2_X1 U5137 ( .A1(n4865), .A2(n4863), .ZN(n4862) );
  INV_X1 U5138 ( .A(n8207), .ZN(n4863) );
  NOR2_X1 U5139 ( .A1(n8969), .A2(n4866), .ZN(n4865) );
  OR2_X1 U5140 ( .A1(n8975), .A2(n8841), .ZN(n8207) );
  AND2_X1 U5141 ( .A1(n6624), .A2(n6401), .ZN(n8877) );
  NAND2_X1 U5142 ( .A1(n6494), .A2(n8141), .ZN(n10156) );
  NAND2_X1 U5143 ( .A1(n8222), .A2(n4399), .ZN(n4852) );
  NAND2_X1 U5144 ( .A1(n4779), .A2(n8145), .ZN(n10248) );
  NAND2_X1 U5145 ( .A1(n5895), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5896) );
  NAND3_X1 U5146 ( .A1(n5859), .A2(n5977), .A3(n5858), .ZN(n5871) );
  AND4_X1 U5147 ( .A1(n6114), .A2(n5854), .A3(n5853), .A4(n5852), .ZN(n5859)
         );
  INV_X1 U5148 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5856) );
  AND2_X1 U5149 ( .A1(n5823), .A2(n5822), .ZN(n6470) );
  NAND2_X1 U5150 ( .A1(n4435), .A2(n4518), .ZN(n4515) );
  INV_X1 U5151 ( .A(n5009), .ZN(n5460) );
  INV_X1 U5152 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4950) );
  AND2_X1 U5153 ( .A1(n5455), .A2(n5479), .ZN(n9517) );
  NAND2_X1 U5154 ( .A1(n5427), .A2(n4699), .ZN(n9532) );
  NOR2_X1 U5155 ( .A1(n4427), .A2(n4608), .ZN(n4607) );
  NOR2_X1 U5156 ( .A1(n9709), .A2(n4708), .ZN(n4707) );
  INV_X1 U5157 ( .A(n9218), .ZN(n4708) );
  NAND2_X1 U5158 ( .A1(n5477), .A2(n5476), .ZN(n9637) );
  INV_X1 U5159 ( .A(n6428), .ZN(n5306) );
  INV_X1 U5160 ( .A(n4986), .ZN(n5164) );
  NAND2_X1 U5161 ( .A1(n5552), .A2(n5551), .ZN(n5582) );
  AND2_X1 U5162 ( .A1(n7568), .A2(n10228), .ZN(n8993) );
  OAI22_X1 U5163 ( .A1(n7986), .A2(n4476), .B1(n8097), .B2(n7985), .ZN(n4475)
         );
  OAI21_X1 U5164 ( .B1(n4476), .B2(n7998), .A(n4473), .ZN(n4472) );
  AND2_X1 U5165 ( .A1(n7996), .A2(n7997), .ZN(n4473) );
  NAND2_X1 U5166 ( .A1(n4589), .A2(n4587), .ZN(n9180) );
  OAI21_X1 U5167 ( .B1(n9172), .B2(n9303), .A(n4588), .ZN(n4587) );
  NAND2_X1 U5168 ( .A1(n9173), .A2(n9284), .ZN(n4589) );
  AOI21_X1 U5169 ( .B1(n9191), .B2(n9190), .A(n9189), .ZN(n4597) );
  OAI21_X1 U5170 ( .B1(n4505), .B2(n4504), .A(n4503), .ZN(n4502) );
  AND2_X1 U5171 ( .A1(n8042), .A2(n4441), .ZN(n4503) );
  OAI21_X1 U5172 ( .B1(n8029), .B2(n8097), .A(n8158), .ZN(n4504) );
  NOR2_X1 U5173 ( .A1(n8028), .A2(n8098), .ZN(n4505) );
  AND2_X1 U5174 ( .A1(n8045), .A2(n8851), .ZN(n4501) );
  OAI21_X1 U5175 ( .B1(n4573), .B2(n4577), .A(n4579), .ZN(n4572) );
  NOR2_X1 U5176 ( .A1(n9209), .A2(n4573), .ZN(n4570) );
  AND2_X1 U5177 ( .A1(n4578), .A2(n9208), .ZN(n4577) );
  NAND2_X1 U5178 ( .A1(n9220), .A2(n4411), .ZN(n4575) );
  NAND2_X1 U5179 ( .A1(n4489), .A2(n4485), .ZN(n8065) );
  NOR2_X1 U5180 ( .A1(n4486), .A2(n8757), .ZN(n4485) );
  AOI21_X1 U5181 ( .B1(n4482), .B2(n4400), .A(n4432), .ZN(n4479) );
  NAND2_X1 U5182 ( .A1(n4562), .A2(n4561), .ZN(n9260) );
  NAND2_X1 U5183 ( .A1(n4498), .A2(n4500), .ZN(n4497) );
  INV_X1 U5184 ( .A(n8101), .ZN(n4499) );
  AND2_X1 U5185 ( .A1(n4872), .A2(n4918), .ZN(n4871) );
  NAND2_X1 U5186 ( .A1(n5105), .A2(n5107), .ZN(n4872) );
  INV_X1 U5187 ( .A(n4670), .ZN(n4669) );
  OAI21_X1 U5188 ( .B1(n6404), .B2(n4671), .A(n6426), .ZN(n4670) );
  NAND2_X1 U5189 ( .A1(n5222), .A2(n5221), .ZN(n5240) );
  NAND2_X1 U5190 ( .A1(n5161), .A2(n8653), .ZN(n5178) );
  XNOR2_X1 U5191 ( .A(n5984), .B(n6894), .ZN(n5940) );
  NAND2_X1 U5192 ( .A1(n6491), .A2(n8142), .ZN(n5941) );
  INV_X1 U5193 ( .A(n6190), .ZN(n4794) );
  NAND2_X1 U5194 ( .A1(n8137), .A2(n8100), .ZN(n8167) );
  OR2_X1 U5195 ( .A1(n8935), .A2(n8271), .ZN(n8124) );
  OR2_X1 U5196 ( .A1(n8926), .A2(n8260), .ZN(n8126) );
  OR2_X1 U5197 ( .A1(n8969), .A2(n8859), .ZN(n8109) );
  INV_X1 U5198 ( .A(n8007), .ZN(n4754) );
  INV_X1 U5199 ( .A(n4760), .ZN(n4755) );
  OR2_X1 U5200 ( .A1(n8685), .A2(n8204), .ZN(n8130) );
  OR2_X1 U5201 ( .A1(n8724), .A2(n8730), .ZN(n8731) );
  NOR2_X1 U5202 ( .A1(n8952), .A2(n4543), .ZN(n4542) );
  INV_X1 U5203 ( .A(n4544), .ZN(n4543) );
  INV_X1 U5204 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U5205 ( .A1(n7284), .A2(n4884), .ZN(n4883) );
  INV_X1 U5206 ( .A(n7285), .ZN(n4884) );
  NAND2_X1 U5207 ( .A1(n5638), .A2(n7285), .ZN(n4882) );
  OAI21_X1 U5208 ( .B1(n5684), .B2(n4905), .A(n4903), .ZN(n5702) );
  AOI21_X1 U5209 ( .B1(n9053), .B2(n4906), .A(n4904), .ZN(n4903) );
  INV_X1 U5210 ( .A(n4906), .ZN(n4905) );
  INV_X1 U5211 ( .A(n9109), .ZN(n4904) );
  AOI21_X1 U5212 ( .B1(n9270), .B2(n6439), .A(n4582), .ZN(n4581) );
  OR2_X1 U5213 ( .A1(n9761), .A2(n9581), .ZN(n9336) );
  OR2_X1 U5214 ( .A1(n5334), .A2(n9044), .ZN(n5352) );
  AND2_X1 U5215 ( .A1(n9851), .A2(n9787), .ZN(n9299) );
  NOR2_X1 U5216 ( .A1(n9685), .A2(n4636), .ZN(n4635) );
  OR2_X1 U5217 ( .A1(n9727), .A2(n9802), .ZN(n4636) );
  OR2_X1 U5218 ( .A1(n5170), .A2(n9054), .ZN(n5193) );
  OR2_X1 U5219 ( .A1(n7603), .A2(n10017), .ZN(n9346) );
  NOR2_X1 U5220 ( .A1(n5539), .A2(n4509), .ZN(n5584) );
  AND2_X1 U5221 ( .A1(n5445), .A2(n5434), .ZN(n5443) );
  NAND2_X1 U5222 ( .A1(n5544), .A2(n4902), .ZN(n4901) );
  INV_X1 U5223 ( .A(n5341), .ZN(n4642) );
  INV_X1 U5224 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n4930) );
  NAND2_X1 U5225 ( .A1(n5296), .A2(n5295), .ZN(n4685) );
  INV_X1 U5226 ( .A(n5294), .ZN(n5295) );
  NOR2_X1 U5227 ( .A1(n5160), .A2(n4664), .ZN(n4663) );
  INV_X1 U5228 ( .A(n5144), .ZN(n4664) );
  XNOR2_X1 U5229 ( .A(n5158), .B(n8590), .ZN(n5157) );
  AOI21_X1 U5230 ( .B1(n4791), .B2(n4795), .A(n4789), .ZN(n4788) );
  INV_X1 U5231 ( .A(n7770), .ZN(n4789) );
  NAND2_X1 U5232 ( .A1(n8311), .A2(n4408), .ZN(n10119) );
  XNOR2_X1 U5233 ( .A(n5940), .B(n5941), .ZN(n6825) );
  AOI21_X1 U5234 ( .B1(n4807), .B2(n7853), .A(n4805), .ZN(n4804) );
  INV_X1 U5235 ( .A(n6255), .ZN(n4805) );
  OR2_X1 U5236 ( .A1(n6282), .A2(n6281), .ZN(n6284) );
  INV_X1 U5237 ( .A(n4917), .ZN(n4808) );
  AND2_X1 U5238 ( .A1(n8291), .A2(n4808), .ZN(n4807) );
  INV_X1 U5239 ( .A(n8104), .ZN(n8171) );
  INV_X1 U5240 ( .A(n8100), .ZN(n8138) );
  INV_X1 U5241 ( .A(n8168), .ZN(n8139) );
  OAI21_X1 U5242 ( .B1(n4492), .B2(n4490), .A(n4493), .ZN(n8173) );
  INV_X1 U5243 ( .A(n4494), .ZN(n4493) );
  INV_X1 U5244 ( .A(n8082), .ZN(n4492) );
  NAND2_X1 U5245 ( .A1(n8083), .A2(n4491), .ZN(n4490) );
  AND4_X1 U5246 ( .A1(n6206), .A2(n6205), .A3(n6204), .A4(n6203), .ZN(n7963)
         );
  NOR2_X1 U5247 ( .A1(n6709), .A2(n6708), .ZN(n6707) );
  NOR2_X1 U5248 ( .A1(n6707), .A2(n4718), .ZN(n6657) );
  AND2_X1 U5249 ( .A1(n6644), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4718) );
  OR2_X1 U5250 ( .A1(n6657), .A2(n6656), .ZN(n4717) );
  OR2_X1 U5251 ( .A1(n6672), .A2(n6671), .ZN(n4722) );
  AND2_X1 U5252 ( .A1(n4722), .A2(n4721), .ZN(n6751) );
  NAND2_X1 U5253 ( .A1(n6748), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4721) );
  OR2_X1 U5254 ( .A1(n6751), .A2(n6750), .ZN(n4720) );
  NOR2_X1 U5255 ( .A1(n8926), .A2(n8731), .ZN(n8716) );
  INV_X1 U5256 ( .A(n4831), .ZN(n4830) );
  OAI21_X1 U5257 ( .B1(n8708), .B2(n4832), .A(n8701), .ZN(n4831) );
  INV_X1 U5258 ( .A(n8215), .ZN(n4832) );
  NAND2_X1 U5259 ( .A1(n8214), .A2(n8260), .ZN(n8215) );
  OR2_X1 U5260 ( .A1(n8724), .A2(n8751), .ZN(n8213) );
  NAND2_X1 U5261 ( .A1(n8709), .A2(n8708), .ZN(n8707) );
  NOR2_X1 U5262 ( .A1(n8940), .A2(n8947), .ZN(n8768) );
  AOI21_X1 U5263 ( .B1(n4835), .B2(n8776), .A(n4433), .ZN(n4833) );
  AND2_X1 U5264 ( .A1(n8123), .A2(n8117), .ZN(n4771) );
  NAND2_X1 U5265 ( .A1(n4769), .A2(n8120), .ZN(n4768) );
  NAND2_X1 U5266 ( .A1(n8123), .A2(n4770), .ZN(n4769) );
  NAND2_X1 U5267 ( .A1(n4541), .A2(n8251), .ZN(n4837) );
  AND2_X1 U5268 ( .A1(n8120), .A2(n8119), .ZN(n8776) );
  AND2_X1 U5269 ( .A1(n8757), .A2(n4837), .ZN(n4835) );
  NAND2_X1 U5270 ( .A1(n8823), .A2(n8117), .ZN(n4774) );
  OR2_X1 U5271 ( .A1(n6230), .A2(n8547), .ZN(n6246) );
  OR2_X1 U5272 ( .A1(n8966), .A2(n8842), .ZN(n8208) );
  NAND2_X1 U5273 ( .A1(n4860), .A2(n4859), .ZN(n8209) );
  NOR2_X1 U5274 ( .A1(n4861), .A2(n4418), .ZN(n4859) );
  AND2_X1 U5275 ( .A1(n8862), .A2(n8870), .ZN(n8863) );
  AND2_X1 U5276 ( .A1(n8838), .A2(n8863), .ZN(n8834) );
  AND2_X1 U5277 ( .A1(n8980), .A2(n8330), .ZN(n8205) );
  OR3_X1 U5278 ( .A1(n6181), .A2(n6180), .A3(n6179), .ZN(n6182) );
  AOI21_X1 U5279 ( .B1(n7722), .B2(n7969), .A(n4763), .ZN(n4762) );
  INV_X1 U5280 ( .A(n8030), .ZN(n4763) );
  NAND2_X1 U5281 ( .A1(n7799), .A2(n7798), .ZN(n7871) );
  OR2_X1 U5282 ( .A1(n6121), .A2(n5885), .ZN(n6137) );
  NAND2_X1 U5283 ( .A1(n7087), .A2(n7086), .ZN(n8890) );
  INV_X1 U5284 ( .A(n8893), .ZN(n7086) );
  OAI21_X1 U5285 ( .B1(n7099), .B2(n7092), .A(n7984), .ZN(n8876) );
  AND3_X1 U5286 ( .A1(n5965), .A2(n5964), .A3(n5963), .ZN(n6912) );
  OR2_X1 U5287 ( .A1(n4394), .A2(n9019), .ZN(n8076) );
  AND2_X1 U5288 ( .A1(n8086), .A2(n8085), .ZN(n8904) );
  OR2_X1 U5289 ( .A1(n4395), .A2(n8235), .ZN(n8085) );
  NAND2_X1 U5290 ( .A1(n6244), .A2(n6243), .ZN(n8958) );
  OR2_X1 U5291 ( .A1(n4395), .A2(n7245), .ZN(n6243) );
  NAND2_X1 U5292 ( .A1(n6178), .A2(n6177), .ZN(n8984) );
  AND3_X1 U5293 ( .A1(n5983), .A2(n5982), .A3(n5981), .ZN(n10202) );
  OR2_X1 U5294 ( .A1(n4394), .A2(n6538), .ZN(n5981) );
  NAND2_X1 U5295 ( .A1(n6505), .A2(n6347), .ZN(n10213) );
  INV_X1 U5296 ( .A(n5863), .ZN(n4855) );
  INV_X1 U5297 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5855) );
  NAND2_X1 U5298 ( .A1(n5026), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5066) );
  NAND2_X1 U5299 ( .A1(n5134), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5151) );
  NAND2_X1 U5300 ( .A1(n4898), .A2(n5651), .ZN(n7635) );
  INV_X1 U5301 ( .A(n4898), .ZN(n4895) );
  NAND2_X1 U5302 ( .A1(n4511), .A2(n4886), .ZN(n9050) );
  AOI21_X1 U5303 ( .B1(n4888), .B2(n4890), .A(n4426), .ZN(n4886) );
  NAND2_X1 U5304 ( .A1(n7617), .A2(n4888), .ZN(n4511) );
  NAND2_X1 U5305 ( .A1(n5047), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5051) );
  AND2_X1 U5306 ( .A1(n5806), .A2(n5805), .ZN(n9089) );
  OAI22_X1 U5307 ( .A1(n7389), .A2(n6457), .B1(n7056), .B2(n5649), .ZN(n5583)
         );
  OR2_X1 U5308 ( .A1(n5086), .A2(n7638), .ZN(n5117) );
  NAND2_X1 U5309 ( .A1(n4892), .A2(n4896), .ZN(n7618) );
  NAND2_X1 U5310 ( .A1(n7634), .A2(n5652), .ZN(n4896) );
  NOR2_X1 U5311 ( .A1(n4894), .A2(n4897), .ZN(n4893) );
  INV_X1 U5312 ( .A(n9034), .ZN(n4537) );
  AND2_X1 U5313 ( .A1(n4443), .A2(n5660), .ZN(n4891) );
  OAI22_X1 U5314 ( .A1(n7312), .A2(n6457), .B1(n5607), .B2(n5649), .ZN(n5608)
         );
  OR2_X1 U5315 ( .A1(n9332), .A2(n5584), .ZN(n7131) );
  NAND2_X1 U5316 ( .A1(n5419), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5454) );
  INV_X1 U5317 ( .A(n5420), .ZN(n5419) );
  OR2_X1 U5318 ( .A1(n5234), .A2(n5233), .ZN(n5253) );
  NAND2_X1 U5319 ( .A1(n5207), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5234) );
  INV_X1 U5320 ( .A(n5208), .ZN(n5207) );
  AND2_X1 U5321 ( .A1(n5409), .A2(n5408), .ZN(n9545) );
  OR2_X1 U5322 ( .A1(n5210), .A2(n6612), .ZN(n4968) );
  AND2_X1 U5323 ( .A1(n6959), .A2(n4741), .ZN(n6792) );
  NAND2_X1 U5324 ( .A1(n6594), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4741) );
  OR2_X1 U5325 ( .A1(n6792), .A2(n6791), .ZN(n4740) );
  INV_X1 U5326 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4520) );
  NOR2_X1 U5327 ( .A1(n6871), .A2(n4735), .ZN(n6874) );
  NOR2_X1 U5328 ( .A1(n6863), .A2(n4736), .ZN(n4735) );
  NOR2_X1 U5329 ( .A1(n6874), .A2(n6873), .ZN(n7219) );
  OR2_X1 U5330 ( .A1(n7650), .A2(n7649), .ZN(n4733) );
  AOI21_X1 U5331 ( .B1(n9517), .B2(n4964), .A(n5461), .ZN(n9534) );
  OAI22_X1 U5332 ( .A1(n9540), .A2(n5535), .B1(n9836), .B2(n9533), .ZN(n9524)
         );
  NAND2_X1 U5333 ( .A1(n5359), .A2(n9297), .ZN(n9599) );
  NAND2_X1 U5334 ( .A1(n9606), .A2(n5528), .ZN(n4609) );
  AOI21_X1 U5335 ( .B1(n5526), .B2(n4605), .A(n4421), .ZN(n4604) );
  INV_X1 U5336 ( .A(n5524), .ZN(n4605) );
  NOR2_X1 U5337 ( .A1(n9225), .A2(n4706), .ZN(n4705) );
  INV_X1 U5338 ( .A(n9369), .ZN(n4706) );
  NAND2_X1 U5339 ( .A1(n7698), .A2(n5215), .ZN(n7753) );
  OR2_X1 U5340 ( .A1(n7747), .A2(n9816), .ZN(n7762) );
  NOR2_X1 U5341 ( .A1(n9311), .A2(n4599), .ZN(n4598) );
  INV_X1 U5342 ( .A(n5496), .ZN(n4599) );
  OAI21_X1 U5343 ( .B1(n7383), .B2(n4612), .A(n4610), .ZN(n7329) );
  NAND2_X1 U5344 ( .A1(n7383), .A2(n5494), .ZN(n7384) );
  OR2_X1 U5345 ( .A1(n10032), .A2(n5539), .ZN(n9695) );
  NAND2_X1 U5346 ( .A1(n9532), .A2(n9390), .ZN(n6442) );
  NAND2_X1 U5347 ( .A1(n5232), .A2(n5231), .ZN(n7846) );
  AND4_X1 U5348 ( .A1(n5072), .A2(n5071), .A3(n5070), .A4(n5069), .ZN(n7483)
         );
  OR2_X1 U5349 ( .A1(n9332), .A2(n9449), .ZN(n10062) );
  NAND2_X1 U5350 ( .A1(n9869), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4940) );
  OR2_X1 U5351 ( .A1(n4941), .A2(n5187), .ZN(n4942) );
  XNOR2_X1 U5352 ( .A(n6427), .B(n6426), .ZN(n8202) );
  NAND2_X1 U5353 ( .A1(n4668), .A2(n6406), .ZN(n6427) );
  NAND2_X1 U5354 ( .A1(n6405), .A2(n6404), .ZN(n4668) );
  NAND2_X1 U5355 ( .A1(n4675), .A2(n4681), .ZN(n5429) );
  NAND2_X1 U5356 ( .A1(n5394), .A2(n4683), .ZN(n4675) );
  INV_X1 U5357 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5541) );
  AND2_X1 U5358 ( .A1(n5378), .A2(n5366), .ZN(n5376) );
  XNOR2_X1 U5359 ( .A(n5362), .B(n5361), .ZN(n7426) );
  NAND2_X1 U5360 ( .A1(n5468), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U5361 ( .A1(n4646), .A2(n4649), .ZN(n5261) );
  NAND2_X1 U5362 ( .A1(n5220), .A2(n4652), .ZN(n4646) );
  OAI21_X1 U5363 ( .B1(n5145), .B2(n4407), .A(n4659), .ZN(n5200) );
  NOR2_X1 U5364 ( .A1(n5112), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5465) );
  INV_X1 U5365 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8525) );
  NOR2_X1 U5366 ( .A1(n5015), .A2(n4877), .ZN(n5033) );
  NOR2_X1 U5367 ( .A1(n9901), .A2(n10304), .ZN(n9902) );
  INV_X1 U5368 ( .A(n4512), .ZN(n6839) );
  OAI21_X1 U5369 ( .B1(n5592), .B2(n4514), .A(n4513), .ZN(n4512) );
  AOI21_X1 U5370 ( .B1(n5596), .B2(n10034), .A(n5594), .ZN(n4513) );
  INV_X1 U5371 ( .A(n5593), .ZN(n4514) );
  OR2_X1 U5372 ( .A1(n4394), .A2(n7883), .ZN(n6314) );
  XNOR2_X1 U5373 ( .A(n6292), .B(n6280), .ZN(n8238) );
  INV_X1 U5374 ( .A(n4820), .ZN(n4811) );
  AND2_X1 U5375 ( .A1(n4815), .A2(n4814), .ZN(n4813) );
  INV_X1 U5376 ( .A(n4816), .ZN(n4815) );
  NAND2_X1 U5377 ( .A1(n4820), .A2(n4822), .ZN(n4814) );
  OAI21_X1 U5378 ( .B1(n6386), .B2(n4817), .A(n6385), .ZN(n4816) );
  NAND2_X1 U5379 ( .A1(n4819), .A2(n4823), .ZN(n4818) );
  INV_X1 U5380 ( .A(n6386), .ZN(n4819) );
  NAND2_X1 U5381 ( .A1(n6201), .A2(n6200), .ZN(n8975) );
  OR2_X1 U5382 ( .A1(n5953), .A2(n5967), .ZN(n5970) );
  NAND2_X1 U5383 ( .A1(n8087), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5958) );
  AND2_X1 U5384 ( .A1(n6641), .A2(n6640), .ZN(n8382) );
  AND2_X1 U5385 ( .A1(n4551), .A2(n4550), .ZN(n8906) );
  NAND2_X1 U5386 ( .A1(n8683), .A2(n8905), .ZN(n4551) );
  AND2_X1 U5387 ( .A1(n4752), .A2(n4412), .ZN(n8712) );
  NAND2_X1 U5388 ( .A1(n4752), .A2(n4750), .ZN(n8711) );
  NAND2_X1 U5389 ( .A1(n8227), .A2(n8226), .ZN(n8228) );
  AOI22_X1 U5390 ( .A1(n8906), .A2(n10215), .B1(n8905), .B2(n10213), .ZN(n8907) );
  NAND2_X1 U5391 ( .A1(n8674), .A2(n4851), .ZN(n4850) );
  NOR2_X1 U5392 ( .A1(n8222), .A2(n4399), .ZN(n4851) );
  NOR2_X1 U5393 ( .A1(n10260), .A2(n8993), .ZN(n4853) );
  OR2_X1 U5394 ( .A1(n8907), .A2(n10260), .ZN(n4845) );
  NAND2_X1 U5395 ( .A1(n5206), .A2(n5205), .ZN(n9030) );
  AND2_X1 U5396 ( .A1(n9148), .A2(n4922), .ZN(n6479) );
  NAND2_X1 U5397 ( .A1(n4567), .A2(n4566), .ZN(n9447) );
  NAND2_X1 U5398 ( .A1(n9403), .A2(n4390), .ZN(n4566) );
  NAND2_X1 U5399 ( .A1(n4568), .A2(n4509), .ZN(n4567) );
  NAND2_X1 U5400 ( .A1(n9444), .A2(n9443), .ZN(n9445) );
  INV_X1 U5401 ( .A(n7373), .ZN(n9467) );
  NAND2_X1 U5402 ( .A1(n4618), .A2(n9287), .ZN(n4617) );
  NAND2_X1 U5403 ( .A1(n9753), .A2(n4616), .ZN(n9556) );
  OR2_X1 U5404 ( .A1(n5848), .A2(n5847), .ZN(n10008) );
  AND2_X1 U5405 ( .A1(n8189), .A2(n9731), .ZN(n8184) );
  NAND2_X1 U5406 ( .A1(n10076), .A2(n9803), .ZN(n9864) );
  XNOR2_X1 U5407 ( .A(n6419), .B(n6418), .ZN(n9868) );
  NAND2_X1 U5408 ( .A1(n6416), .A2(n6415), .ZN(n6419) );
  NOR2_X1 U5409 ( .A1(n8415), .A2(n10305), .ZN(n10304) );
  NOR2_X1 U5410 ( .A1(n10319), .A2(n10318), .ZN(n10317) );
  AOI21_X1 U5411 ( .B1(n4474), .B2(n4471), .A(n8000), .ZN(n8005) );
  NAND2_X1 U5412 ( .A1(n4472), .A2(n8097), .ZN(n4471) );
  AOI21_X1 U5413 ( .B1(n9191), .B2(n9375), .A(n9365), .ZN(n4594) );
  NOR2_X1 U5414 ( .A1(n9284), .A2(n4593), .ZN(n4592) );
  INV_X1 U5415 ( .A(n9344), .ZN(n4593) );
  AND2_X1 U5416 ( .A1(n9193), .A2(n9284), .ZN(n4596) );
  NAND2_X1 U5417 ( .A1(n4403), .A2(n4574), .ZN(n4573) );
  NAND2_X1 U5418 ( .A1(n4578), .A2(n4576), .ZN(n4574) );
  OR2_X1 U5419 ( .A1(n9207), .A2(n9284), .ZN(n4576) );
  NAND2_X1 U5420 ( .A1(n4502), .A2(n4501), .ZN(n8046) );
  NAND2_X1 U5421 ( .A1(n4575), .A2(n4571), .ZN(n9228) );
  NOR2_X1 U5422 ( .A1(n4417), .A2(n4586), .ZN(n4585) );
  NOR2_X1 U5423 ( .A1(n9541), .A2(n9284), .ZN(n4586) );
  INV_X1 U5424 ( .A(n5125), .ZN(n4868) );
  INV_X1 U5425 ( .A(n7999), .ZN(n4761) );
  NOR2_X1 U5426 ( .A1(n4908), .A2(n4907), .ZN(n4906) );
  INV_X1 U5427 ( .A(n9110), .ZN(n4908) );
  INV_X1 U5428 ( .A(n5685), .ZN(n4907) );
  OR2_X1 U5429 ( .A1(n9269), .A2(n9284), .ZN(n4582) );
  INV_X1 U5430 ( .A(n6406), .ZN(n4671) );
  NOR2_X1 U5431 ( .A1(n4679), .A2(n4674), .ZN(n4673) );
  INV_X1 U5432 ( .A(n5378), .ZN(n4674) );
  INV_X1 U5433 ( .A(n4681), .ZN(n4679) );
  INV_X1 U5434 ( .A(n4683), .ZN(n4678) );
  INV_X1 U5435 ( .A(n5428), .ZN(n4677) );
  INV_X1 U5436 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4927) );
  INV_X1 U5437 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n4928) );
  NAND2_X1 U5438 ( .A1(n5300), .A2(n5299), .ZN(n5317) );
  AOI21_X1 U5439 ( .B1(n4649), .B2(n4651), .A(n4648), .ZN(n4647) );
  INV_X1 U5440 ( .A(n5260), .ZN(n4648) );
  INV_X1 U5441 ( .A(n5199), .ZN(n4657) );
  NOR2_X1 U5442 ( .A1(n4499), .A2(n8091), .ZN(n4491) );
  OAI211_X1 U5443 ( .C1(n4499), .C2(n4496), .A(n4495), .B(n8145), .ZN(n4494)
         );
  INV_X1 U5444 ( .A(n8102), .ZN(n4496) );
  OR2_X1 U5445 ( .A1(n4499), .A2(n4497), .ZN(n4495) );
  NOR2_X1 U5446 ( .A1(n6081), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n6115) );
  INV_X1 U5447 ( .A(SI_11_), .ZN(n8590) );
  OR2_X1 U5448 ( .A1(n6316), .A2(n8195), .ZN(n6336) );
  AND2_X1 U5449 ( .A1(n8124), .A2(n8062), .ZN(n8212) );
  INV_X1 U5450 ( .A(n4772), .ZN(n4770) );
  NOR2_X1 U5451 ( .A1(n8160), .A2(n4773), .ZN(n4772) );
  NOR2_X1 U5452 ( .A1(n4559), .A2(n8984), .ZN(n4557) );
  NAND2_X1 U5453 ( .A1(n7717), .A2(n4560), .ZN(n4559) );
  INV_X1 U5454 ( .A(n8033), .ZN(n4560) );
  OR2_X1 U5455 ( .A1(n7574), .A2(n7969), .ZN(n7723) );
  NAND2_X1 U5456 ( .A1(n7345), .A2(n7405), .ZN(n8015) );
  OR2_X1 U5457 ( .A1(n7345), .A2(n7405), .ZN(n7973) );
  NOR2_X1 U5458 ( .A1(n10125), .A2(n10085), .ZN(n4554) );
  NAND2_X1 U5459 ( .A1(n8875), .A2(n4760), .ZN(n4759) );
  NAND2_X1 U5460 ( .A1(n6903), .A2(n6902), .ZN(n7978) );
  INV_X1 U5461 ( .A(n8337), .ZN(n6903) );
  NAND2_X1 U5462 ( .A1(n6490), .A2(n6830), .ZN(n7990) );
  OR2_X1 U5463 ( .A1(n7161), .A2(n10135), .ZN(n8883) );
  NAND2_X1 U5464 ( .A1(n6358), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6379) );
  AND2_X1 U5465 ( .A1(n4402), .A2(n5873), .ZN(n4797) );
  CLKBUF_X1 U5466 ( .A(n5871), .Z(n6353) );
  NOR2_X1 U5467 ( .A1(n6013), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n6033) );
  INV_X1 U5468 ( .A(n4889), .ZN(n4888) );
  OAI21_X1 U5469 ( .B1(n4891), .B2(n4890), .A(n7791), .ZN(n4889) );
  INV_X1 U5470 ( .A(n5668), .ZN(n4890) );
  NOR2_X1 U5471 ( .A1(n7634), .A2(n5652), .ZN(n4897) );
  INV_X1 U5472 ( .A(n7455), .ZN(n4894) );
  NAND2_X1 U5473 ( .A1(n9101), .A2(n4536), .ZN(n4527) );
  OR2_X1 U5474 ( .A1(n5776), .A2(n9043), .ZN(n5782) );
  NAND2_X1 U5475 ( .A1(n9063), .A2(n4519), .ZN(n4518) );
  INV_X1 U5476 ( .A(n5806), .ZN(n4519) );
  CLKBUF_X1 U5477 ( .A(n5653), .Z(n6456) );
  NOR2_X1 U5478 ( .A1(n7543), .A2(n4737), .ZN(n7646) );
  AND2_X1 U5479 ( .A1(n7544), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4737) );
  NOR2_X1 U5480 ( .A1(n9501), .A2(n4624), .ZN(n4622) );
  INV_X1 U5481 ( .A(n4699), .ZN(n4696) );
  INV_X1 U5482 ( .A(n9272), .ZN(n4695) );
  NOR2_X1 U5483 ( .A1(n4640), .A2(n9563), .ZN(n4639) );
  INV_X1 U5484 ( .A(n4641), .ZN(n4640) );
  NOR2_X1 U5485 ( .A1(n9756), .A2(n9761), .ZN(n4641) );
  INV_X1 U5486 ( .A(n5529), .ZN(n4608) );
  OR2_X1 U5487 ( .A1(n9618), .A2(n9603), .ZN(n9297) );
  NOR2_X1 U5488 ( .A1(n5514), .A2(n7758), .ZN(n4924) );
  INV_X1 U5489 ( .A(n5193), .ZN(n5191) );
  AND2_X1 U5490 ( .A1(n7644), .A2(n7462), .ZN(n4630) );
  INV_X1 U5491 ( .A(n5494), .ZN(n4611) );
  NAND2_X1 U5492 ( .A1(n7476), .A2(n5497), .ZN(n10010) );
  NOR2_X1 U5493 ( .A1(n5411), .A2(n4684), .ZN(n4683) );
  INV_X1 U5494 ( .A(n5392), .ZN(n4684) );
  AOI21_X1 U5495 ( .B1(n4683), .B2(n5393), .A(n4682), .ZN(n4681) );
  INV_X1 U5496 ( .A(n5410), .ZN(n4682) );
  NAND2_X1 U5497 ( .A1(n5466), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5475) );
  OR2_X1 U5498 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(n5462), .ZN(n5463) );
  OAI21_X1 U5499 ( .B1(n5316), .B2(n5315), .A(n5317), .ZN(n5329) );
  AND2_X1 U5500 ( .A1(n5330), .A2(n5320), .ZN(n5328) );
  INV_X1 U5501 ( .A(n5219), .ZN(n4653) );
  INV_X1 U5502 ( .A(n5159), .ZN(n4661) );
  INV_X1 U5503 ( .A(n4660), .ZN(n4659) );
  OAI21_X1 U5504 ( .B1(n4663), .B2(n4407), .A(n5178), .ZN(n4660) );
  NAND2_X1 U5505 ( .A1(n5098), .A2(n5097), .ZN(n5107) );
  INV_X1 U5506 ( .A(SI_7_), .ZN(n8589) );
  NOR2_X1 U5507 ( .A1(n4843), .A2(n4844), .ZN(n4842) );
  NAND2_X1 U5508 ( .A1(n5039), .A2(n4839), .ZN(n4838) );
  NAND2_X1 U5509 ( .A1(n4926), .A2(n4878), .ZN(n4877) );
  INV_X1 U5510 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4878) );
  INV_X1 U5511 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4926) );
  NAND2_X1 U5512 ( .A1(n4389), .A2(n4424), .ZN(n4956) );
  NAND2_X1 U5513 ( .A1(n4781), .A2(n4780), .ZN(n7551) );
  AND2_X1 U5514 ( .A1(n6162), .A2(n6146), .ZN(n4780) );
  NAND2_X1 U5515 ( .A1(n5891), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6282) );
  INV_X1 U5516 ( .A(n6269), .ZN(n5891) );
  NAND2_X1 U5517 ( .A1(n4434), .A2(n4823), .ZN(n4817) );
  INV_X1 U5518 ( .A(n4823), .ZN(n4822) );
  INV_X1 U5519 ( .A(n4800), .ZN(n4799) );
  OAI21_X1 U5520 ( .B1(n4408), .B2(n4801), .A(n10120), .ZN(n4800) );
  INV_X1 U5521 ( .A(n6048), .ZN(n4801) );
  NAND2_X1 U5522 ( .A1(n4779), .A2(n4778), .ZN(n8142) );
  NOR2_X1 U5523 ( .A1(n8170), .A2(n8734), .ZN(n4778) );
  NAND2_X1 U5524 ( .A1(n6242), .A2(n6241), .ZN(n4809) );
  NAND2_X1 U5525 ( .A1(n4786), .A2(n6096), .ZN(n10096) );
  INV_X1 U5526 ( .A(n10099), .ZN(n4786) );
  INV_X1 U5527 ( .A(n4792), .ZN(n4791) );
  OAI21_X1 U5528 ( .B1(n7625), .B2(n4793), .A(n6209), .ZN(n4792) );
  NAND2_X1 U5529 ( .A1(n6198), .A2(n4794), .ZN(n4793) );
  OR2_X1 U5530 ( .A1(n7625), .A2(n4796), .ZN(n4795) );
  INV_X1 U5531 ( .A(n6198), .ZN(n4796) );
  NOR2_X1 U5532 ( .A1(n4686), .A2(n8167), .ZN(n8169) );
  NOR2_X1 U5533 ( .A1(n8165), .A2(n8166), .ZN(n4687) );
  AND2_X1 U5534 ( .A1(n6289), .A2(n6288), .ZN(n8236) );
  AND3_X1 U5535 ( .A1(n6250), .A2(n6249), .A3(n6248), .ZN(n8827) );
  AND2_X1 U5536 ( .A1(n4717), .A2(n4716), .ZN(n6695) );
  NAND2_X1 U5537 ( .A1(n6632), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4716) );
  AND2_X1 U5538 ( .A1(n4720), .A2(n4719), .ZN(n6931) );
  NAND2_X1 U5539 ( .A1(n6928), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4719) );
  NOR2_X1 U5540 ( .A1(n6983), .A2(n4724), .ZN(n6987) );
  AND2_X1 U5541 ( .A1(n6984), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4724) );
  NOR2_X1 U5542 ( .A1(n6987), .A2(n6986), .ZN(n7070) );
  NOR2_X1 U5543 ( .A1(n7070), .A2(n4723), .ZN(n7072) );
  AND2_X1 U5544 ( .A1(n7071), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4723) );
  NOR2_X1 U5545 ( .A1(n7072), .A2(n7073), .ZN(n7252) );
  NAND2_X1 U5546 ( .A1(n7511), .A2(n4710), .ZN(n7513) );
  OR2_X1 U5547 ( .A1(n7512), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4710) );
  NAND2_X1 U5548 ( .A1(n7513), .A2(n7514), .ZN(n7826) );
  NAND2_X1 U5549 ( .A1(n7826), .A2(n4709), .ZN(n7886) );
  OR2_X1 U5550 ( .A1(n7829), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4709) );
  NOR2_X1 U5551 ( .A1(n8357), .A2(n4468), .ZN(n8361) );
  NAND2_X1 U5552 ( .A1(n8361), .A2(n8360), .ZN(n8374) );
  AND2_X1 U5553 ( .A1(n6400), .A2(n6399), .ZN(n8682) );
  OR2_X1 U5554 ( .A1(n4395), .A2(n7914), .ZN(n6345) );
  NAND2_X1 U5555 ( .A1(n4829), .A2(n4828), .ZN(n8676) );
  AOI21_X1 U5556 ( .B1(n4830), .B2(n4832), .A(n4456), .ZN(n4828) );
  NAND2_X1 U5557 ( .A1(n8726), .A2(n8163), .ZN(n4752) );
  INV_X1 U5558 ( .A(n8212), .ZN(n8748) );
  NAND2_X1 U5559 ( .A1(n4774), .A2(n4772), .ZN(n8793) );
  NAND2_X1 U5560 ( .A1(n5890), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6258) );
  AND2_X1 U5561 ( .A1(n8118), .A2(n8114), .ZN(n8805) );
  INV_X1 U5562 ( .A(n8825), .ZN(n8112) );
  AOI21_X1 U5563 ( .B1(n8106), .B2(n7966), .A(n4766), .ZN(n4765) );
  INV_X1 U5564 ( .A(n8107), .ZN(n4766) );
  AND4_X1 U5565 ( .A1(n6172), .A2(n6171), .A3(n6170), .A4(n6169), .ZN(n8857)
         );
  NAND2_X1 U5566 ( .A1(n5887), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6215) );
  INV_X1 U5567 ( .A(n6182), .ZN(n5887) );
  NOR2_X1 U5568 ( .A1(n10168), .A2(n4556), .ZN(n8862) );
  NAND2_X1 U5569 ( .A1(n4557), .A2(n7813), .ZN(n4556) );
  OR2_X1 U5570 ( .A1(n7807), .A2(n7966), .ZN(n8853) );
  NOR2_X1 U5571 ( .A1(n10168), .A2(n4555), .ZN(n7872) );
  INV_X1 U5572 ( .A(n4557), .ZN(n4555) );
  AND4_X1 U5573 ( .A1(n6142), .A2(n6141), .A3(n6140), .A4(n6139), .ZN(n8032)
         );
  NAND2_X1 U5574 ( .A1(n7723), .A2(n7722), .ZN(n7804) );
  NOR2_X1 U5575 ( .A1(n7416), .A2(n7345), .ZN(n7417) );
  INV_X1 U5576 ( .A(n8156), .ZN(n7569) );
  AND4_X1 U5577 ( .A1(n6127), .A2(n6126), .A3(n6125), .A4(n6124), .ZN(n7576)
         );
  NAND2_X1 U5578 ( .A1(n7407), .A2(n7406), .ZN(n7411) );
  NAND2_X2 U5579 ( .A1(n7973), .A2(n8015), .ZN(n8155) );
  OAI21_X1 U5580 ( .B1(n8875), .B2(n4756), .A(n4753), .ZN(n7271) );
  INV_X1 U5581 ( .A(n4757), .ZN(n4756) );
  NAND2_X1 U5582 ( .A1(n4552), .A2(n8885), .ZN(n7416) );
  NOR2_X1 U5583 ( .A1(n4553), .A2(n7341), .ZN(n4552) );
  INV_X1 U5584 ( .A(n4554), .ZN(n4553) );
  NAND2_X1 U5585 ( .A1(n8885), .A2(n4554), .ZN(n7275) );
  NAND2_X1 U5586 ( .A1(n4759), .A2(n8002), .ZN(n7175) );
  NOR2_X1 U5587 ( .A1(n8883), .A2(n10214), .ZN(n8885) );
  AND2_X1 U5588 ( .A1(n8885), .A2(n10222), .ZN(n7181) );
  INV_X1 U5589 ( .A(n10156), .ZN(n8854) );
  AND2_X1 U5590 ( .A1(n4539), .A2(n4538), .ZN(n7160) );
  NOR2_X1 U5591 ( .A1(n6902), .A2(n6913), .ZN(n4538) );
  NAND2_X1 U5592 ( .A1(n7160), .A2(n10202), .ZN(n7161) );
  NAND2_X1 U5593 ( .A1(n4539), .A2(n10195), .ZN(n7037) );
  OR2_X1 U5594 ( .A1(n6497), .A2(n7109), .ZN(n7110) );
  OR2_X1 U5595 ( .A1(n10186), .A2(n6374), .ZN(n6919) );
  NAND2_X1 U5596 ( .A1(n8094), .A2(n8093), .ZN(n8390) );
  OR2_X1 U5597 ( .A1(n4394), .A2(n6574), .ZN(n8093) );
  XNOR2_X1 U5598 ( .A(n8899), .B(n8390), .ZN(n8898) );
  NAND2_X1 U5599 ( .A1(n8834), .A2(n4415), .ZN(n8947) );
  INV_X1 U5600 ( .A(n10213), .ZN(n10255) );
  OR2_X1 U5601 ( .A1(n6853), .A2(n6852), .ZN(n6921) );
  NAND2_X1 U5602 ( .A1(n4540), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5865) );
  NAND2_X1 U5603 ( .A1(n4856), .A2(n4858), .ZN(n4540) );
  NAND2_X1 U5604 ( .A1(n6379), .A2(n6378), .ZN(n6381) );
  INV_X1 U5605 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6356) );
  INV_X1 U5606 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5879) );
  NAND2_X1 U5607 ( .A1(n4858), .A2(n4402), .ZN(n6210) );
  OR2_X1 U5608 ( .A1(n6049), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n6051) );
  OR2_X1 U5609 ( .A1(n5979), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n6013) );
  NAND2_X1 U5610 ( .A1(n5638), .A2(n7285), .ZN(n4885) );
  INV_X1 U5611 ( .A(n5066), .ZN(n5064) );
  NAND2_X1 U5612 ( .A1(n4529), .A2(n4530), .ZN(n9041) );
  INV_X1 U5613 ( .A(n4531), .ZN(n4530) );
  OAI21_X1 U5614 ( .B1(n4536), .B2(n4532), .A(n9101), .ZN(n4531) );
  AND2_X1 U5615 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5047) );
  NAND2_X1 U5616 ( .A1(n7029), .A2(n5626), .ZN(n5630) );
  OR2_X1 U5617 ( .A1(n9071), .A2(n9072), .ZN(n9080) );
  XNOR2_X1 U5618 ( .A(n5618), .B(n6460), .ZN(n5619) );
  NAND2_X1 U5619 ( .A1(n5617), .A2(n5616), .ZN(n5618) );
  INV_X1 U5620 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6767) );
  OR2_X1 U5621 ( .A1(n5117), .A2(n6767), .ZN(n5135) );
  NAND2_X1 U5622 ( .A1(n5323), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5334) );
  INV_X1 U5623 ( .A(n5324), .ZN(n5323) );
  OR2_X1 U5624 ( .A1(n5309), .A2(n9036), .ZN(n5324) );
  NAND2_X1 U5625 ( .A1(n5684), .A2(n5683), .ZN(n9051) );
  AND2_X1 U5626 ( .A1(n5772), .A2(n4534), .ZN(n4533) );
  NAND2_X1 U5627 ( .A1(n9101), .A2(n4532), .ZN(n4534) );
  NOR2_X1 U5628 ( .A1(n4528), .A2(n4527), .ZN(n4526) );
  INV_X1 U5629 ( .A(n5792), .ZN(n4528) );
  AND2_X1 U5630 ( .A1(n9121), .A2(n9123), .ZN(n5792) );
  NAND2_X1 U5631 ( .A1(n4521), .A2(n4533), .ZN(n9122) );
  NAND2_X1 U5632 ( .A1(n4537), .A2(n4522), .ZN(n4521) );
  INV_X1 U5633 ( .A(n4527), .ZN(n4522) );
  INV_X1 U5634 ( .A(n5403), .ZN(n5401) );
  NAND2_X1 U5635 ( .A1(n5713), .A2(n5712), .ZN(n9157) );
  NAND2_X1 U5636 ( .A1(n4569), .A2(n9293), .ZN(n9406) );
  NAND2_X1 U5637 ( .A1(n9286), .A2(n9285), .ZN(n4569) );
  AND4_X1 U5638 ( .A1(n5239), .A2(n5238), .A3(n5237), .A4(n5236), .ZN(n9074)
         );
  OR2_X1 U5639 ( .A1(n4990), .A2(n4972), .ZN(n4974) );
  NOR2_X1 U5640 ( .A1(n6803), .A2(n4452), .ZN(n9938) );
  NOR2_X1 U5641 ( .A1(n4877), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n4875) );
  NAND2_X1 U5642 ( .A1(n9938), .A2(n9939), .ZN(n9937) );
  NOR2_X1 U5643 ( .A1(n7219), .A2(n4450), .ZN(n9964) );
  NAND2_X1 U5644 ( .A1(n9964), .A2(n9963), .ZN(n9962) );
  OR2_X1 U5645 ( .A1(n5304), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5165) );
  OR2_X1 U5646 ( .A1(n5165), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5186) );
  NOR2_X1 U5647 ( .A1(n9971), .A2(n4738), .ZN(n7223) );
  AND2_X1 U5648 ( .A1(n9976), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4738) );
  NOR2_X1 U5649 ( .A1(n7223), .A2(n7222), .ZN(n7543) );
  XNOR2_X1 U5650 ( .A(n7646), .B(n7645), .ZN(n7545) );
  NOR2_X1 U5651 ( .A1(n9484), .A2(n4728), .ZN(n9989) );
  AND2_X1 U5652 ( .A1(n9487), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4728) );
  NOR2_X1 U5653 ( .A1(n9989), .A2(n9988), .ZN(n9987) );
  OR2_X1 U5654 ( .A1(n5582), .A2(n7499), .ZN(n6968) );
  AND2_X1 U5655 ( .A1(n4622), .A2(n9290), .ZN(n4621) );
  INV_X1 U5656 ( .A(n4622), .ZN(n4618) );
  OR2_X1 U5657 ( .A1(n5487), .A2(n9290), .ZN(n4619) );
  OAI21_X1 U5658 ( .B1(n5427), .B2(n4697), .A(n4694), .ZN(n6443) );
  INV_X1 U5659 ( .A(n4698), .ZN(n4697) );
  AOI21_X1 U5660 ( .B1(n4696), .B2(n4698), .A(n4695), .ZN(n4694) );
  NOR2_X1 U5661 ( .A1(n6441), .A2(n9274), .ZN(n4698) );
  OAI21_X1 U5662 ( .B1(n5533), .B2(n4615), .A(n4614), .ZN(n9540) );
  INV_X1 U5663 ( .A(n4616), .ZN(n4615) );
  AOI21_X1 U5664 ( .B1(n4616), .B2(n9583), .A(n4425), .ZN(n4614) );
  NAND2_X1 U5665 ( .A1(n9589), .A2(n4637), .ZN(n9525) );
  NOR2_X1 U5666 ( .A1(n4638), .A2(n9265), .ZN(n4637) );
  INV_X1 U5667 ( .A(n4639), .ZN(n4638) );
  AND2_X1 U5668 ( .A1(n9558), .A2(n5534), .ZN(n4616) );
  NAND2_X1 U5669 ( .A1(n9589), .A2(n4641), .ZN(n9572) );
  OR2_X1 U5670 ( .A1(n5369), .A2(n6521), .ZN(n5382) );
  NOR2_X1 U5671 ( .A1(n9298), .A2(n9340), .ZN(n4693) );
  AOI21_X1 U5672 ( .B1(n4602), .B2(n4606), .A(n4423), .ZN(n4601) );
  OR2_X1 U5673 ( .A1(n9722), .A2(n4634), .ZN(n9653) );
  NAND2_X1 U5674 ( .A1(n5485), .A2(n4635), .ZN(n4634) );
  AND2_X1 U5675 ( .A1(n9333), .A2(n9234), .ZN(n9661) );
  NOR2_X1 U5676 ( .A1(n9722), .A2(n4633), .ZN(n9674) );
  INV_X1 U5677 ( .A(n4635), .ZN(n4633) );
  NAND2_X1 U5678 ( .A1(n5252), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5267) );
  OR2_X1 U5679 ( .A1(n5267), .A2(n9083), .ZN(n5287) );
  OR2_X1 U5680 ( .A1(n9222), .A2(n9225), .ZN(n9697) );
  NOR2_X1 U5681 ( .A1(n7762), .A2(n9030), .ZN(n7843) );
  AND2_X1 U5682 ( .A1(n9206), .A2(n9343), .ZN(n9318) );
  OR2_X1 U5683 ( .A1(n7662), .A2(n9058), .ZN(n7747) );
  AND4_X1 U5684 ( .A1(n5176), .A2(n5175), .A3(n5174), .A4(n5173), .ZN(n9113)
         );
  AND2_X1 U5685 ( .A1(n7333), .A2(n4626), .ZN(n7663) );
  NOR2_X1 U5686 ( .A1(n4628), .A2(n7603), .ZN(n4626) );
  NAND2_X1 U5687 ( .A1(n7333), .A2(n4630), .ZN(n10002) );
  NOR2_X1 U5688 ( .A1(n7393), .A2(n7394), .ZN(n7392) );
  AND2_X1 U5689 ( .A1(n7392), .A2(n7469), .ZN(n7333) );
  AND4_X1 U5690 ( .A1(n5014), .A2(n5013), .A3(n5012), .A4(n5011), .ZN(n7389)
         );
  OR2_X1 U5691 ( .A1(n7317), .A2(n7371), .ZN(n7393) );
  NOR2_X1 U5692 ( .A1(n7204), .A2(n6998), .ZN(n7318) );
  OR2_X1 U5693 ( .A1(n9284), .A2(n5539), .ZN(n5848) );
  OR2_X1 U5694 ( .A1(n4388), .A2(n10034), .ZN(n7204) );
  INV_X1 U5695 ( .A(n9695), .ZN(n10003) );
  NAND2_X1 U5696 ( .A1(n5451), .A2(n5450), .ZN(n6464) );
  NAND2_X1 U5697 ( .A1(n5436), .A2(n5435), .ZN(n9737) );
  AND4_X1 U5698 ( .A1(n5056), .A2(n5055), .A3(n5054), .A4(n5053), .ZN(n7373)
         );
  AND2_X1 U5699 ( .A1(n5832), .A2(n9449), .ZN(n9819) );
  AND2_X1 U5700 ( .A1(n6881), .A2(n5570), .ZN(n9803) );
  XNOR2_X1 U5701 ( .A(n6423), .B(SI_30_), .ZN(n8234) );
  NAND2_X1 U5702 ( .A1(n5444), .A2(n5443), .ZN(n5446) );
  AND2_X1 U5703 ( .A1(n6406), .A2(n5449), .ZN(n6404) );
  INV_X1 U5704 ( .A(n4901), .ZN(n4900) );
  XNOR2_X1 U5705 ( .A(n5444), .B(n5443), .ZN(n7859) );
  INV_X1 U5706 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5544) );
  INV_X1 U5707 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5228) );
  INV_X1 U5708 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U5709 ( .A1(n4654), .A2(n5219), .ZN(n5242) );
  NAND2_X1 U5710 ( .A1(n4655), .A2(n5216), .ZN(n4654) );
  INV_X1 U5711 ( .A(n5220), .ZN(n4655) );
  NAND2_X1 U5712 ( .A1(n4662), .A2(n5159), .ZN(n5180) );
  NAND2_X1 U5713 ( .A1(n5145), .A2(n4663), .ZN(n4662) );
  CLKBUF_X1 U5714 ( .A(n6080), .Z(n5130) );
  INV_X1 U5715 ( .A(n5022), .ZN(n4844) );
  XNOR2_X1 U5716 ( .A(n5040), .B(SI_5_), .ZN(n5058) );
  NAND2_X1 U5717 ( .A1(n5020), .A2(n5019), .ZN(n5023) );
  NAND2_X1 U5718 ( .A1(n4876), .A2(n4926), .ZN(n5017) );
  NOR2_X1 U5719 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4925) );
  AND2_X1 U5720 ( .A1(n8311), .A2(n6030), .ZN(n10087) );
  AND4_X1 U5721 ( .A1(n6188), .A2(n6187), .A3(n6186), .A4(n6185), .ZN(n7800)
         );
  NAND2_X1 U5722 ( .A1(n4781), .A2(n6146), .ZN(n7553) );
  INV_X1 U5723 ( .A(n6824), .ZN(n5939) );
  AOI21_X1 U5724 ( .B1(n4804), .B2(n4806), .A(n4464), .ZN(n4802) );
  INV_X1 U5725 ( .A(n4807), .ZN(n4806) );
  OR2_X1 U5726 ( .A1(n4394), .A2(n7305), .ZN(n6256) );
  NOR2_X1 U5727 ( .A1(n8257), .A2(n8258), .ZN(n8256) );
  NAND2_X1 U5728 ( .A1(n6167), .A2(n6166), .ZN(n8980) );
  NAND2_X1 U5729 ( .A1(n8283), .A2(n5998), .ZN(n10142) );
  NAND2_X1 U5730 ( .A1(n4790), .A2(n6198), .ZN(n7626) );
  NAND2_X1 U5731 ( .A1(n7687), .A2(n6190), .ZN(n4790) );
  OR2_X1 U5732 ( .A1(n4394), .A2(n7593), .ZN(n5910) );
  OR2_X1 U5733 ( .A1(n4394), .A2(n7933), .ZN(n6266) );
  INV_X1 U5734 ( .A(n4784), .ZN(n4783) );
  OAI21_X1 U5735 ( .B1(n6096), .B2(n4785), .A(n7116), .ZN(n4784) );
  NAND2_X1 U5736 ( .A1(n6393), .A2(n6383), .ZN(n10098) );
  AND4_X1 U5737 ( .A1(n6236), .A2(n6235), .A3(n6234), .A4(n6233), .ZN(n8293)
         );
  INV_X1 U5738 ( .A(n10138), .ZN(n10130) );
  AND2_X1 U5739 ( .A1(n8241), .A2(n8877), .ZN(n10140) );
  AND2_X1 U5740 ( .A1(n5907), .A2(n5906), .ZN(n8322) );
  INV_X1 U5741 ( .A(n10098), .ZN(n10145) );
  AND4_X1 U5742 ( .A1(n6156), .A2(n6155), .A3(n6154), .A4(n6153), .ZN(n7711)
         );
  AND2_X1 U5743 ( .A1(n8241), .A2(n8879), .ZN(n10138) );
  NAND2_X1 U5744 ( .A1(n6626), .A2(n10190), .ZN(n10176) );
  INV_X1 U5745 ( .A(n8877), .ZN(n8856) );
  INV_X1 U5746 ( .A(n8322), .ZN(n8751) );
  INV_X1 U5747 ( .A(n8236), .ZN(n8779) );
  OR2_X1 U5748 ( .A1(n6626), .A2(n6488), .ZN(n8338) );
  INV_X1 U5749 ( .A(n4717), .ZN(n6655) );
  INV_X1 U5750 ( .A(n4722), .ZN(n6747) );
  INV_X1 U5751 ( .A(n4720), .ZN(n6927) );
  XNOR2_X1 U5752 ( .A(n7886), .B(n7887), .ZN(n7828) );
  INV_X1 U5753 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8388) );
  XNOR2_X1 U5754 ( .A(n4711), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8380) );
  NAND2_X1 U5755 ( .A1(n8374), .A2(n4712), .ZN(n4711) );
  OR2_X1 U5756 ( .A1(n8375), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n4712) );
  INV_X1 U5757 ( .A(n8904), .ZN(n8134) );
  NAND2_X1 U5758 ( .A1(n8707), .A2(n8215), .ZN(n8693) );
  OAI21_X1 U5759 ( .B1(n8709), .B2(n4832), .A(n4830), .ZN(n8692) );
  OR2_X1 U5760 ( .A1(n4395), .A2(n7823), .ZN(n6299) );
  OR2_X1 U5761 ( .A1(n4395), .A2(n7731), .ZN(n5869) );
  NAND2_X1 U5762 ( .A1(n6279), .A2(n6278), .ZN(n8940) );
  OR2_X1 U5763 ( .A1(n4395), .A2(n7504), .ZN(n6278) );
  OR2_X1 U5764 ( .A1(n8774), .A2(n8776), .ZN(n4836) );
  NAND2_X1 U5765 ( .A1(n8834), .A2(n8820), .ZN(n8809) );
  AND2_X1 U5766 ( .A1(n4860), .A2(n4864), .ZN(n8816) );
  NAND2_X1 U5767 ( .A1(n8847), .A2(n8207), .ZN(n8833) );
  NAND2_X1 U5768 ( .A1(n7713), .A2(n7712), .ZN(n7716) );
  NAND2_X1 U5769 ( .A1(n8890), .A2(n7088), .ZN(n7090) );
  NAND2_X1 U5770 ( .A1(n8875), .A2(n7999), .ZN(n7173) );
  CLKBUF_X1 U5771 ( .A(n8890), .Z(n8891) );
  OR2_X1 U5772 ( .A1(n10176), .A2(n6850), .ZN(n8888) );
  INV_X1 U5773 ( .A(n6504), .ZN(n8780) );
  INV_X1 U5774 ( .A(n8869), .ZN(n10161) );
  AND2_X1 U5775 ( .A1(n6390), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10190) );
  NAND2_X1 U5776 ( .A1(n4858), .A2(n4776), .ZN(n4775) );
  NOR2_X1 U5777 ( .A1(n6352), .A2(n4855), .ZN(n4776) );
  NOR2_X1 U5778 ( .A1(n5871), .A2(n6352), .ZN(n6362) );
  INV_X1 U5779 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6979) );
  INV_X1 U5780 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6950) );
  INV_X1 U5781 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n8464) );
  INV_X1 U5782 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6745) );
  INV_X1 U5783 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6611) );
  INV_X1 U5784 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6561) );
  INV_X1 U5785 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n8604) );
  INV_X1 U5786 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n8529) );
  NAND2_X1 U5787 ( .A1(n5934), .A2(n4713), .ZN(n6692) );
  AOI22_X1 U5788 ( .A1(n4431), .A2(P2_IR_REG_0__SCAN_IN), .B1(n4715), .B2(
        n4714), .ZN(n4713) );
  AND4_X1 U5789 ( .A1(n5091), .A2(n5090), .A3(n5089), .A4(n5088), .ZN(n10016)
         );
  AND2_X1 U5790 ( .A1(n5388), .A2(n5387), .ZN(n6522) );
  AND4_X1 U5791 ( .A1(n5156), .A2(n5155), .A3(n5154), .A4(n5153), .ZN(n7746)
         );
  NAND2_X1 U5792 ( .A1(n7617), .A2(n5660), .ZN(n7679) );
  NAND2_X1 U5793 ( .A1(n6476), .A2(n6475), .ZN(n6477) );
  NAND2_X1 U5794 ( .A1(n7635), .A2(n7634), .ZN(n7632) );
  NAND2_X1 U5795 ( .A1(n5604), .A2(n5603), .ZN(n5606) );
  NAND2_X1 U5796 ( .A1(n9088), .A2(n5806), .ZN(n9062) );
  CLKBUF_X1 U5797 ( .A(n9069), .Z(n9071) );
  AND4_X1 U5798 ( .A1(n5141), .A2(n5140), .A3(n5139), .A4(n5138), .ZN(n10017)
         );
  INV_X1 U5799 ( .A(n9651), .ZN(n9776) );
  NAND2_X1 U5800 ( .A1(n4537), .A2(n4536), .ZN(n4535) );
  NAND2_X1 U5801 ( .A1(n5190), .A2(n5189), .ZN(n9816) );
  AND3_X1 U5802 ( .A1(n5338), .A2(n5337), .A3(n5336), .ZN(n9777) );
  NAND2_X1 U5803 ( .A1(n4525), .A2(n4523), .ZN(n9127) );
  NAND2_X1 U5804 ( .A1(n5792), .A2(n4524), .ZN(n4523) );
  NAND2_X1 U5805 ( .A1(n4537), .A2(n4526), .ZN(n4525) );
  INV_X1 U5806 ( .A(n4533), .ZN(n4524) );
  CLKBUF_X1 U5807 ( .A(n9120), .Z(n9126) );
  NAND2_X1 U5808 ( .A1(n7617), .A2(n4891), .ZN(n4887) );
  INV_X1 U5809 ( .A(n9806), .ZN(n9721) );
  INV_X1 U5810 ( .A(n9170), .ZN(n9142) );
  OR2_X1 U5811 ( .A1(n5838), .A2(n6834), .ZN(n9092) );
  AND2_X1 U5812 ( .A1(n9149), .A2(n9146), .ZN(n5817) );
  AND4_X1 U5813 ( .A1(n5258), .A2(n5257), .A3(n5256), .A4(n5255), .ZN(n9699)
         );
  AND2_X1 U5814 ( .A1(n5843), .A2(n9449), .ZN(n9167) );
  INV_X1 U5815 ( .A(n9545), .ZN(n9578) );
  INV_X1 U5816 ( .A(n6522), .ZN(n9600) );
  AOI22_X1 U5817 ( .A1(n5009), .A2(P1_REG2_REG_1__SCAN_IN), .B1(n9876), .B2(
        n4874), .ZN(n4947) );
  OR2_X1 U5818 ( .A1(n5210), .A2(n10077), .ZN(n4946) );
  OR2_X1 U5819 ( .A1(n6968), .A2(P1_U3084), .ZN(n9471) );
  OR2_X1 U5820 ( .A1(n4990), .A2(n6884), .ZN(n4966) );
  INV_X1 U5821 ( .A(n4740), .ZN(n6790) );
  AND2_X1 U5822 ( .A1(n4740), .A2(n4739), .ZN(n9923) );
  NAND2_X1 U5823 ( .A1(n6596), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4739) );
  NAND2_X1 U5824 ( .A1(n9948), .A2(n9949), .ZN(n9947) );
  NAND2_X1 U5825 ( .A1(n9937), .A2(n4729), .ZN(n9948) );
  NAND2_X1 U5826 ( .A1(n6772), .A2(n6771), .ZN(n4729) );
  INV_X1 U5827 ( .A(n4733), .ZN(n7936) );
  OAI21_X1 U5828 ( .B1(n7650), .B2(n4731), .A(n4730), .ZN(n9472) );
  NAND2_X1 U5829 ( .A1(n4734), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4731) );
  NAND2_X1 U5830 ( .A1(n7937), .A2(n4734), .ZN(n4730) );
  INV_X1 U5831 ( .A(n9473), .ZN(n4734) );
  INV_X1 U5832 ( .A(n7937), .ZN(n4732) );
  INV_X1 U5833 ( .A(n9966), .ZN(n9986) );
  XNOR2_X1 U5834 ( .A(n4726), .B(n4725), .ZN(n7949) );
  INV_X1 U5835 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n4725) );
  OR2_X1 U5836 ( .A1(n9987), .A2(n4727), .ZN(n4726) );
  AND2_X1 U5837 ( .A1(n9993), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4727) );
  NOR2_X1 U5838 ( .A1(n9502), .A2(n9695), .ZN(n9733) );
  NAND2_X1 U5839 ( .A1(n5427), .A2(n9385), .ZN(n9531) );
  NAND2_X1 U5840 ( .A1(n5533), .A2(n5532), .ZN(n9753) );
  NAND2_X1 U5841 ( .A1(n4609), .A2(n5529), .ZN(n9588) );
  NAND2_X1 U5842 ( .A1(n4603), .A2(n4604), .ZN(n9647) );
  OR2_X1 U5843 ( .A1(n5525), .A2(n4606), .ZN(n4603) );
  NAND2_X1 U5844 ( .A1(n5308), .A2(n5307), .ZN(n9670) );
  NAND2_X1 U5845 ( .A1(n5266), .A2(n5265), .ZN(n9802) );
  NAND2_X1 U5846 ( .A1(n5251), .A2(n5250), .ZN(n9727) );
  NAND2_X1 U5847 ( .A1(n7753), .A2(n9218), .ZN(n7840) );
  NAND2_X1 U5848 ( .A1(n5148), .A2(n5147), .ZN(n7794) );
  NAND2_X1 U5849 ( .A1(n7328), .A2(n5496), .ZN(n7478) );
  AND2_X1 U5850 ( .A1(n7384), .A2(n5495), .ZN(n7231) );
  NAND2_X1 U5851 ( .A1(n9629), .A2(n7134), .ZN(n9623) );
  AND4_X1 U5852 ( .A1(n5032), .A2(n5031), .A3(n5030), .A4(n5029), .ZN(n10063)
         );
  INV_X1 U5853 ( .A(n9706), .ZN(n9714) );
  OR2_X1 U5854 ( .A1(n7133), .A2(n4509), .ZN(n9724) );
  INV_X1 U5855 ( .A(n9623), .ZN(n10028) );
  INV_X1 U5856 ( .A(n10008), .ZN(n10035) );
  INV_X1 U5857 ( .A(n9657), .ZN(n9851) );
  INV_X1 U5858 ( .A(n7448), .ZN(n7462) );
  INV_X1 U5859 ( .A(n5635), .ZN(n7469) );
  INV_X1 U5860 ( .A(n10047), .ZN(n10048) );
  AND2_X1 U5861 ( .A1(n5582), .A2(n5555), .ZN(n10051) );
  NAND2_X1 U5862 ( .A1(n4941), .A2(n4939), .ZN(n9869) );
  XNOR2_X1 U5863 ( .A(n6405), .B(n6404), .ZN(n7911) );
  XNOR2_X1 U5864 ( .A(n5548), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U5865 ( .A1(n5547), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U5866 ( .A1(n5547), .A2(n5543), .ZN(n7733) );
  XNOR2_X1 U5867 ( .A(n5470), .B(n8603), .ZN(n9405) );
  NAND2_X1 U5868 ( .A1(n5474), .A2(n5473), .ZN(n9398) );
  NAND2_X1 U5869 ( .A1(n5472), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n5473) );
  INV_X1 U5870 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5305) );
  OAI21_X1 U5871 ( .B1(n5304), .B2(n5462), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4510) );
  INV_X1 U5872 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n8634) );
  INV_X1 U5873 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8436) );
  INV_X1 U5874 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6609) );
  INV_X1 U5875 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6555) );
  INV_X1 U5876 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6551) );
  XNOR2_X1 U5877 ( .A(n4960), .B(n4959), .ZN(n6592) );
  NOR2_X1 U5878 ( .A1(n9904), .A2(n10317), .ZN(n10303) );
  AOI21_X1 U5879 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10301), .ZN(n10300) );
  NOR2_X1 U5880 ( .A1(n10300), .A2(n10299), .ZN(n10298) );
  NAND2_X1 U5881 ( .A1(n4813), .A2(n4818), .ZN(n4812) );
  NOR2_X1 U5882 ( .A1(n8908), .A2(n4392), .ZN(n8230) );
  AND2_X1 U5883 ( .A1(n8908), .A2(n8907), .ZN(n4854) );
  NAND2_X1 U5884 ( .A1(n4848), .A2(n4393), .ZN(n4847) );
  INV_X1 U5885 ( .A(n6454), .ZN(n6455) );
  MUX2_X1 U5886 ( .A(n8185), .B(n8184), .S(n10076), .Z(n8186) );
  NOR2_X1 U5887 ( .A1(n5572), .A2(n5571), .ZN(n5573) );
  NAND2_X1 U5888 ( .A1(n5576), .A2(n10076), .ZN(n5574) );
  AND2_X1 U5889 ( .A1(n8689), .A2(n8204), .ZN(n4399) );
  NAND2_X1 U5890 ( .A1(n6267), .A2(n6266), .ZN(n8946) );
  INV_X1 U5891 ( .A(n8946), .ZN(n4541) );
  AND2_X1 U5892 ( .A1(n7958), .A2(n8098), .ZN(n4400) );
  NAND2_X1 U5893 ( .A1(n4809), .A2(n4807), .ZN(n8246) );
  AND2_X1 U5894 ( .A1(n4600), .A2(n4601), .ZN(n4401) );
  XNOR2_X1 U5895 ( .A(n8920), .B(n8681), .ZN(n8701) );
  INV_X1 U5896 ( .A(n8701), .ZN(n4747) );
  INV_X1 U5897 ( .A(n9709), .ZN(n4578) );
  AND2_X1 U5898 ( .A1(n5872), .A2(n4798), .ZN(n4402) );
  NAND2_X1 U5899 ( .A1(n5796), .A2(n5795), .ZN(n6516) );
  XNOR2_X1 U5900 ( .A(n5037), .B(SI_4_), .ZN(n5035) );
  AND2_X1 U5901 ( .A1(n9221), .A2(n9712), .ZN(n4403) );
  INV_X1 U5902 ( .A(n5539), .ZN(n9443) );
  XNOR2_X1 U5903 ( .A(n5475), .B(P1_IR_REG_20__SCAN_IN), .ZN(n5539) );
  NAND2_X1 U5904 ( .A1(n4836), .A2(n4835), .ZN(n8756) );
  INV_X1 U5905 ( .A(n9583), .ZN(n5532) );
  AND2_X1 U5906 ( .A1(n9361), .A2(n9253), .ZN(n9583) );
  NAND2_X1 U5907 ( .A1(n6425), .A2(n6424), .ZN(n9501) );
  AND2_X1 U5908 ( .A1(n6213), .A2(n6212), .ZN(n8838) );
  INV_X1 U5909 ( .A(n8838), .ZN(n8969) );
  AND2_X1 U5910 ( .A1(n9657), .A2(n9769), .ZN(n9298) );
  INV_X1 U5911 ( .A(n4628), .ZN(n4627) );
  NAND2_X1 U5912 ( .A1(n4630), .A2(n4629), .ZN(n4628) );
  AND2_X1 U5913 ( .A1(n4845), .A2(n4463), .ZN(n4404) );
  INV_X1 U5914 ( .A(n9284), .ZN(n4588) );
  INV_X1 U5915 ( .A(n8920), .ZN(n8216) );
  INV_X1 U5916 ( .A(n6452), .ZN(n4625) );
  NAND2_X1 U5917 ( .A1(n4759), .A2(n4757), .ZN(n7269) );
  AND2_X1 U5918 ( .A1(n8834), .A2(n4542), .ZN(n4405) );
  INV_X1 U5919 ( .A(n8260), .ZN(n8728) );
  AND2_X1 U5920 ( .A1(n6311), .A2(n6310), .ZN(n8260) );
  OR2_X1 U5921 ( .A1(n10168), .A2(n8033), .ZN(n4406) );
  NAND2_X1 U5922 ( .A1(n6346), .A2(n6345), .ZN(n8685) );
  NOR2_X1 U5923 ( .A1(n9722), .A2(n4636), .ZN(n9673) );
  INV_X1 U5924 ( .A(n5210), .ZN(n5456) );
  INV_X1 U5925 ( .A(n5953), .ZN(n5901) );
  INV_X1 U5926 ( .A(n4398), .ZN(n6318) );
  NAND2_X1 U5927 ( .A1(n7994), .A2(n7978), .ZN(n6905) );
  OR2_X1 U5928 ( .A1(n5179), .A2(n4661), .ZN(n4407) );
  INV_X1 U5929 ( .A(n9543), .ZN(n4584) );
  AOI21_X1 U5930 ( .B1(n9868), .B2(n5164), .A(n6421), .ZN(n9287) );
  AND2_X1 U5931 ( .A1(n10086), .A2(n6030), .ZN(n4408) );
  INV_X1 U5932 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4714) );
  NOR2_X1 U5933 ( .A1(n10162), .A2(n8334), .ZN(n4409) );
  AND2_X1 U5934 ( .A1(n8002), .A2(n8001), .ZN(n8151) );
  AND3_X1 U5935 ( .A1(n5951), .A2(n5950), .A3(n5949), .ZN(n10195) );
  AND3_X1 U5936 ( .A1(n5873), .A2(n5872), .A3(n5860), .ZN(n4410) );
  AND2_X1 U5937 ( .A1(n4403), .A2(n9284), .ZN(n4411) );
  NAND2_X1 U5938 ( .A1(n5259), .A2(n9369), .ZN(n9696) );
  NAND2_X1 U5939 ( .A1(n5314), .A2(n9234), .ZN(n9645) );
  AND2_X1 U5940 ( .A1(n4900), .A2(n4915), .ZN(n4899) );
  NAND2_X1 U5941 ( .A1(n4535), .A2(n5755), .ZN(n9100) );
  XNOR2_X1 U5942 ( .A(n4983), .B(n4957), .ZN(n4982) );
  OR2_X1 U5943 ( .A1(n8724), .A2(n8322), .ZN(n4412) );
  AND2_X1 U5944 ( .A1(n5144), .A2(n5129), .ZN(n4413) );
  NAND4_X1 U5945 ( .A1(n4968), .A2(n4967), .A3(n4966), .A4(n4965), .ZN(n5593)
         );
  INV_X1 U5946 ( .A(n8127), .ZN(n4749) );
  NAND2_X2 U5947 ( .A1(n4944), .A2(n4945), .ZN(n5010) );
  AND2_X1 U5948 ( .A1(n4836), .A2(n4837), .ZN(n8755) );
  AND2_X1 U5949 ( .A1(n4704), .A2(n10076), .ZN(n4414) );
  OR2_X1 U5950 ( .A1(n9737), .A2(n9546), .ZN(n9390) );
  NAND2_X1 U5951 ( .A1(n5368), .A2(n5367), .ZN(n9761) );
  NAND2_X1 U5952 ( .A1(n6257), .A2(n6256), .ZN(n8952) );
  OR2_X1 U5953 ( .A1(n5553), .A2(n4901), .ZN(n5540) );
  INV_X1 U5954 ( .A(n4650), .ZN(n4649) );
  OAI21_X1 U5955 ( .B1(n5216), .B2(n4651), .A(n5240), .ZN(n4650) );
  AND2_X1 U5956 ( .A1(n4542), .A2(n4541), .ZN(n4415) );
  OR2_X1 U5957 ( .A1(n9278), .A2(n4588), .ZN(n4416) );
  OR2_X1 U5958 ( .A1(n8958), .A2(n8827), .ZN(n8118) );
  INV_X1 U5959 ( .A(n8118), .ZN(n4773) );
  NAND2_X1 U5960 ( .A1(n5446), .A2(n5445), .ZN(n6405) );
  AND2_X1 U5961 ( .A1(n9267), .A2(n9263), .ZN(n4417) );
  NOR2_X1 U5962 ( .A1(n8820), .A2(n8293), .ZN(n4418) );
  AND2_X1 U5963 ( .A1(n9244), .A2(n9608), .ZN(n9634) );
  INV_X1 U5964 ( .A(n9265), .ZN(n9836) );
  NAND2_X1 U5965 ( .A1(n5418), .A2(n5417), .ZN(n9265) );
  AND2_X1 U5966 ( .A1(n6229), .A2(n6228), .ZN(n8820) );
  INV_X1 U5967 ( .A(n8820), .ZN(n8966) );
  AND2_X1 U5968 ( .A1(n4774), .A2(n8118), .ZN(n4419) );
  AND2_X1 U5969 ( .A1(n6012), .A2(n5998), .ZN(n4420) );
  INV_X1 U5970 ( .A(n4751), .ZN(n4750) );
  NAND2_X1 U5971 ( .A1(n8713), .A2(n4412), .ZN(n4751) );
  INV_X1 U5972 ( .A(n9507), .ZN(n4704) );
  INV_X1 U5973 ( .A(n4550), .ZN(n8668) );
  NAND2_X1 U5974 ( .A1(n8716), .A2(n4547), .ZN(n4550) );
  OR2_X1 U5975 ( .A1(n8946), .A2(n8251), .ZN(n8120) );
  AND2_X1 U5976 ( .A1(n9670), .A2(n9651), .ZN(n4421) );
  AND2_X1 U5977 ( .A1(n9192), .A2(n10011), .ZN(n9311) );
  AND2_X1 U5978 ( .A1(n9267), .A2(n9266), .ZN(n4422) );
  NOR2_X1 U5979 ( .A1(n9657), .A2(n9787), .ZN(n4423) );
  AND2_X1 U5980 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4424) );
  NOR2_X1 U5981 ( .A1(n9563), .A2(n9578), .ZN(n4425) );
  NOR2_X1 U5982 ( .A1(n5675), .A2(n5674), .ZN(n4426) );
  AND2_X1 U5983 ( .A1(n9761), .A2(n9614), .ZN(n4427) );
  AND2_X1 U5984 ( .A1(n4481), .A2(n4482), .ZN(n4428) );
  INV_X1 U5985 ( .A(n8091), .ZN(n4498) );
  NAND2_X1 U5986 ( .A1(n7981), .A2(n7995), .ZN(n8147) );
  OR2_X1 U5987 ( .A1(n5553), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4429) );
  AND2_X1 U5988 ( .A1(n4875), .A2(n4520), .ZN(n4430) );
  INV_X1 U5989 ( .A(n4624), .ZN(n4623) );
  NAND2_X1 U5990 ( .A1(n5486), .A2(n4625), .ZN(n4624) );
  INV_X1 U5991 ( .A(n9053), .ZN(n5683) );
  NAND2_X1 U5992 ( .A1(n9589), .A2(n9592), .ZN(n9571) );
  AND2_X1 U5993 ( .A1(n8030), .A2(n8031), .ZN(n8037) );
  INV_X1 U5994 ( .A(n8037), .ZN(n7714) );
  AND2_X1 U5995 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4431) );
  NAND2_X1 U5996 ( .A1(n4412), .A2(n8126), .ZN(n4432) );
  NOR2_X1 U5997 ( .A1(n8211), .A2(n8236), .ZN(n4433) );
  OR2_X1 U5998 ( .A1(n6333), .A2(n6313), .ZN(n4434) );
  INV_X1 U5999 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5873) );
  NAND2_X1 U6000 ( .A1(n9063), .A2(n9089), .ZN(n4435) );
  AND2_X1 U6001 ( .A1(n4899), .A2(n4952), .ZN(n4436) );
  AND2_X1 U6002 ( .A1(n8084), .A2(n8132), .ZN(n8222) );
  AND2_X1 U6003 ( .A1(n9230), .A2(n9234), .ZN(n4437) );
  NOR2_X1 U6004 ( .A1(n9737), .A2(n9458), .ZN(n4438) );
  AND2_X1 U6005 ( .A1(n10063), .A2(n7469), .ZN(n4439) );
  AND2_X1 U6006 ( .A1(n9753), .A2(n5534), .ZN(n4440) );
  AND2_X1 U6007 ( .A1(n8043), .A2(n7806), .ZN(n4441) );
  AND2_X1 U6008 ( .A1(n9390), .A2(n9271), .ZN(n9431) );
  NAND2_X1 U6009 ( .A1(n9657), .A2(n9787), .ZN(n4442) );
  NAND2_X1 U6010 ( .A1(n7677), .A2(n5666), .ZN(n4443) );
  AND2_X1 U6011 ( .A1(n4518), .A2(n6518), .ZN(n4444) );
  AND2_X1 U6012 ( .A1(n5623), .A2(n5622), .ZN(n4445) );
  AND2_X1 U6013 ( .A1(n7172), .A2(n7088), .ZN(n4446) );
  INV_X1 U6014 ( .A(n6097), .ZN(n4785) );
  AND2_X1 U6015 ( .A1(n7714), .A2(n7712), .ZN(n4447) );
  AND2_X1 U6016 ( .A1(n4813), .A2(n4811), .ZN(n4448) );
  NAND2_X1 U6017 ( .A1(n4858), .A2(n4797), .ZN(n5878) );
  INV_X1 U6018 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5895) );
  AND2_X1 U6019 ( .A1(n9589), .A2(n4639), .ZN(n4449) );
  INV_X1 U6020 ( .A(n8681), .ZN(n8714) );
  AND2_X1 U6021 ( .A1(n6325), .A2(n6324), .ZN(n8681) );
  AND2_X1 U6022 ( .A1(n7220), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4450) );
  AND2_X1 U6023 ( .A1(n9051), .A2(n5685), .ZN(n4451) );
  AND2_X1 U6024 ( .A1(n6776), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4452) );
  OAI21_X1 U6025 ( .B1(n7687), .B2(n4795), .A(n4791), .ZN(n7769) );
  NAND2_X1 U6026 ( .A1(n4887), .A2(n5668), .ZN(n7790) );
  AND2_X1 U6027 ( .A1(n8853), .A2(n8106), .ZN(n4453) );
  OR2_X1 U6028 ( .A1(n9722), .A2(n9727), .ZN(n4454) );
  NAND2_X1 U6029 ( .A1(n8077), .A2(n8076), .ZN(n8905) );
  INV_X1 U6030 ( .A(n8905), .ZN(n4548) );
  NOR2_X1 U6031 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6114) );
  AND2_X1 U6032 ( .A1(n7526), .A2(n5500), .ZN(n7666) );
  NAND2_X1 U6033 ( .A1(n6315), .A2(n6314), .ZN(n8920) );
  NAND2_X1 U6034 ( .A1(n4876), .A2(n4875), .ZN(n5073) );
  NAND2_X1 U6035 ( .A1(n5285), .A2(n5284), .ZN(n9685) );
  AND4_X1 U6036 ( .A1(n6221), .A2(n6220), .A3(n6219), .A4(n6218), .ZN(n8859)
         );
  INV_X1 U6037 ( .A(n8859), .ZN(n4866) );
  AND3_X1 U6038 ( .A1(n6273), .A2(n6272), .A3(n6271), .ZN(n8251) );
  AND2_X1 U6039 ( .A1(n6343), .A2(n6342), .ZN(n8204) );
  NAND2_X1 U6040 ( .A1(n5133), .A2(n5132), .ZN(n7603) );
  NAND2_X1 U6041 ( .A1(n8834), .A2(n4544), .ZN(n4545) );
  AND2_X1 U6042 ( .A1(n4733), .A2(n4732), .ZN(n4455) );
  INV_X1 U6043 ( .A(n4652), .ZN(n4651) );
  NOR2_X1 U6044 ( .A1(n5241), .A2(n4653), .ZN(n4652) );
  NAND2_X1 U6045 ( .A1(n4895), .A2(n5652), .ZN(n7631) );
  NAND2_X1 U6046 ( .A1(n6430), .A2(n6429), .ZN(n6452) );
  AND2_X1 U6047 ( .A1(n9639), .A2(n9846), .ZN(n9589) );
  NAND2_X1 U6048 ( .A1(n5104), .A2(n5103), .ZN(n7496) );
  AND2_X1 U6049 ( .A1(n8216), .A2(n8681), .ZN(n4456) );
  AND2_X1 U6050 ( .A1(n7802), .A2(n7966), .ZN(n8206) );
  INV_X1 U6051 ( .A(n5755), .ZN(n4532) );
  NOR2_X1 U6052 ( .A1(n4394), .A2(n8464), .ZN(n4457) );
  OR2_X1 U6053 ( .A1(n9299), .A2(n9232), .ZN(n4458) );
  AND2_X1 U6054 ( .A1(n4852), .A2(n4853), .ZN(n4459) );
  AND2_X1 U6055 ( .A1(n4809), .A2(n4808), .ZN(n4460) );
  AND2_X1 U6056 ( .A1(n6403), .A2(n6402), .ZN(n4461) );
  INV_X1 U6057 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5875) );
  OR2_X1 U6058 ( .A1(n6921), .A2(n6854), .ZN(n10260) );
  NAND2_X1 U6059 ( .A1(n7333), .A2(n7462), .ZN(n7332) );
  NOR2_X1 U6060 ( .A1(n7176), .A2(n4758), .ZN(n4757) );
  XNOR2_X1 U6061 ( .A(n5883), .B(P2_IR_REG_20__SCAN_IN), .ZN(n8170) );
  INV_X1 U6062 ( .A(n8170), .ZN(n8145) );
  AND2_X1 U6063 ( .A1(n7333), .A2(n4627), .ZN(n4462) );
  OR2_X1 U6064 ( .A1(n4393), .A2(n8570), .ZN(n4463) );
  NAND2_X1 U6065 ( .A1(n5142), .A2(n9346), .ZN(n7668) );
  NAND2_X1 U6066 ( .A1(n7325), .A2(n9187), .ZN(n7474) );
  XOR2_X1 U6067 ( .A(n6264), .B(n6262), .Z(n4464) );
  INV_X1 U6068 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4902) );
  NAND2_X1 U6069 ( .A1(n6300), .A2(n6299), .ZN(n8926) );
  INV_X1 U6070 ( .A(n8926), .ZN(n8214) );
  NAND2_X1 U6071 ( .A1(n4873), .A2(n5622), .ZN(n7028) );
  AND2_X1 U6072 ( .A1(n9183), .A2(n5495), .ZN(n4613) );
  NAND2_X1 U6073 ( .A1(n4919), .A2(n5101), .ZN(n5553) );
  INV_X1 U6074 ( .A(n4558), .ZN(n7873) );
  NOR2_X1 U6075 ( .A1(n10168), .A2(n4559), .ZN(n4558) );
  NAND2_X1 U6076 ( .A1(n6362), .A2(n6361), .ZN(n4465) );
  OR2_X1 U6077 ( .A1(n6353), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n4466) );
  INV_X1 U6078 ( .A(n4864), .ZN(n4861) );
  NAND2_X1 U6079 ( .A1(n8969), .A2(n4866), .ZN(n4864) );
  NAND2_X1 U6080 ( .A1(n8179), .A2(n8734), .ZN(n6494) );
  NAND2_X1 U6081 ( .A1(n5116), .A2(n5115), .ZN(n10027) );
  INV_X1 U6082 ( .A(n10027), .ZN(n4629) );
  NOR2_X1 U6083 ( .A1(n8392), .A2(n8104), .ZN(n4467) );
  AND2_X1 U6084 ( .A1(n8358), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4468) );
  NAND2_X1 U6085 ( .A1(n6894), .A2(n7109), .ZN(n7036) );
  INV_X1 U6086 ( .A(n7036), .ZN(n4539) );
  INV_X1 U6087 ( .A(n4390), .ZN(n4509) );
  INV_X1 U6088 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4798) );
  INV_X1 U6089 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4715) );
  INV_X1 U6090 ( .A(n5908), .ZN(n4779) );
  BUF_X1 U6091 ( .A(n5898), .Z(n9013) );
  INV_X1 U6092 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4954) );
  INV_X1 U6093 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n4736) );
  INV_X1 U6094 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4506) );
  NAND3_X1 U6095 ( .A1(n4475), .A2(n7993), .A3(n7996), .ZN(n4474) );
  NAND2_X1 U6096 ( .A1(n8066), .A2(n4482), .ZN(n4480) );
  OR2_X1 U6097 ( .A1(n8066), .A2(n4400), .ZN(n4481) );
  INV_X1 U6098 ( .A(n8092), .ZN(n4500) );
  INV_X1 U6099 ( .A(n8878), .ZN(n7155) );
  NAND3_X1 U6100 ( .A1(n6004), .A2(n6003), .A3(n4508), .ZN(n8878) );
  AOI21_X1 U6101 ( .B1(n5901), .B2(P2_REG0_REG_5__SCAN_IN), .A(n6002), .ZN(
        n4508) );
  NAND2_X1 U6102 ( .A1(n5595), .A2(n6838), .ZN(n5605) );
  NAND4_X1 U6103 ( .A1(n6838), .A2(n5604), .A3(n5595), .A4(n5603), .ZN(n6887)
         );
  NAND2_X1 U6104 ( .A1(n6887), .A2(n6886), .ZN(n6885) );
  NAND2_X1 U6105 ( .A1(n4873), .A2(n4445), .ZN(n7029) );
  AND2_X2 U6106 ( .A1(n5581), .A2(n5582), .ZN(n5596) );
  NAND2_X2 U6107 ( .A1(n5585), .A2(n5653), .ZN(n5592) );
  NAND3_X1 U6108 ( .A1(n5796), .A2(n5795), .A3(n4518), .ZN(n4517) );
  NAND2_X1 U6109 ( .A1(n6517), .A2(n6518), .ZN(n6515) );
  NAND2_X1 U6110 ( .A1(n6517), .A2(n4444), .ZN(n4516) );
  NAND3_X1 U6111 ( .A1(n4517), .A2(n4516), .A3(n4515), .ZN(n9147) );
  NAND3_X1 U6112 ( .A1(n6515), .A2(n9089), .A3(n6516), .ZN(n9088) );
  NAND2_X1 U6113 ( .A1(n9034), .A2(n5755), .ZN(n4529) );
  INV_X1 U6114 ( .A(n9035), .ZN(n4536) );
  INV_X1 U6115 ( .A(n10195), .ZN(n6913) );
  INV_X1 U6116 ( .A(n4545), .ZN(n8808) );
  NAND2_X1 U6117 ( .A1(n8716), .A2(n8216), .ZN(n8695) );
  NAND2_X1 U6118 ( .A1(n8716), .A2(n4546), .ZN(n8683) );
  NAND2_X1 U6119 ( .A1(n9231), .A2(n9230), .ZN(n9237) );
  NAND3_X1 U6120 ( .A1(n9241), .A2(n4563), .A3(n4565), .ZN(n4562) );
  NAND2_X1 U6121 ( .A1(n4564), .A2(n4458), .ZN(n4563) );
  NAND2_X1 U6122 ( .A1(n9231), .A2(n4437), .ZN(n4564) );
  INV_X1 U6123 ( .A(n9248), .ZN(n4565) );
  NOR2_X1 U6124 ( .A1(n4570), .A2(n4572), .ZN(n4571) );
  OAI21_X1 U6125 ( .B1(n4583), .B2(n4422), .A(n9271), .ZN(n9275) );
  AOI21_X1 U6126 ( .B1(n9264), .B2(n4585), .A(n4584), .ZN(n4583) );
  NAND2_X1 U6127 ( .A1(n7309), .A2(n7311), .ZN(n7310) );
  NAND2_X1 U6128 ( .A1(n7198), .A2(n4971), .ZN(n7003) );
  INV_X1 U6129 ( .A(n9305), .ZN(n4590) );
  XNOR2_X2 U6130 ( .A(n5597), .B(n10053), .ZN(n9305) );
  NAND3_X1 U6131 ( .A1(n4595), .A2(n4591), .A3(n9201), .ZN(n9216) );
  OAI21_X1 U6132 ( .B1(n4594), .B2(n9186), .A(n4592), .ZN(n4591) );
  OAI21_X1 U6133 ( .B1(n4597), .B2(n9194), .A(n4596), .ZN(n4595) );
  AND3_X1 U6134 ( .A1(n4919), .A2(n5101), .A3(n4436), .ZN(n4949) );
  NAND2_X1 U6135 ( .A1(n7328), .A2(n4598), .ZN(n7476) );
  NAND2_X1 U6136 ( .A1(n5525), .A2(n4602), .ZN(n4600) );
  NAND2_X1 U6137 ( .A1(n5525), .A2(n5524), .ZN(n9662) );
  INV_X1 U6138 ( .A(n5526), .ZN(n4606) );
  NAND2_X1 U6139 ( .A1(n4609), .A2(n4607), .ZN(n5531) );
  AOI21_X1 U6140 ( .B1(n4613), .B2(n4611), .A(n4439), .ZN(n4610) );
  INV_X1 U6141 ( .A(n4613), .ZN(n4612) );
  NAND2_X1 U6142 ( .A1(n7384), .A2(n4613), .ZN(n7230) );
  AND2_X1 U6143 ( .A1(n5487), .A2(n4623), .ZN(n9499) );
  NAND2_X1 U6144 ( .A1(n5487), .A2(n4621), .ZN(n4620) );
  NAND2_X1 U6145 ( .A1(n5487), .A2(n5486), .ZN(n6451) );
  NAND3_X1 U6146 ( .A1(n4620), .A2(n4619), .A3(n4617), .ZN(n6432) );
  XNOR2_X2 U6147 ( .A(n4631), .B(n4952), .ZN(n7861) );
  NAND3_X1 U6148 ( .A1(n4919), .A2(n4899), .A3(n5101), .ZN(n4632) );
  NAND2_X1 U6149 ( .A1(n5220), .A2(n4647), .ZN(n4645) );
  NAND2_X1 U6150 ( .A1(n5145), .A2(n4659), .ZN(n4658) );
  NAND2_X1 U6151 ( .A1(n5145), .A2(n5144), .ZN(n4824) );
  NAND2_X1 U6152 ( .A1(n6405), .A2(n4669), .ZN(n4667) );
  NAND2_X1 U6153 ( .A1(n5379), .A2(n4673), .ZN(n4672) );
  NAND2_X1 U6154 ( .A1(n4672), .A2(n4676), .ZN(n5431) );
  NAND2_X1 U6155 ( .A1(n8099), .A2(n8096), .ZN(n8168) );
  NAND3_X1 U6156 ( .A1(n8099), .A2(n8096), .A3(n4687), .ZN(n4686) );
  NAND2_X1 U6157 ( .A1(n8390), .A2(n8095), .ZN(n8100) );
  OAI21_X1 U6158 ( .B1(n8909), .B2(n8993), .A(n4854), .ZN(n8997) );
  NAND2_X1 U6159 ( .A1(n7198), .A2(n4688), .ZN(n7200) );
  NAND2_X1 U6160 ( .A1(n4689), .A2(n9305), .ZN(n4688) );
  INV_X1 U6161 ( .A(n7199), .ZN(n4689) );
  NAND2_X1 U6162 ( .A1(n5314), .A2(n4693), .ZN(n9633) );
  NAND2_X1 U6163 ( .A1(n9633), .A2(n5339), .ZN(n9607) );
  NOR2_X1 U6164 ( .A1(n9512), .A2(n9507), .ZN(n4702) );
  NAND2_X1 U6165 ( .A1(n4700), .A2(n6484), .ZN(n6487) );
  NAND3_X1 U6166 ( .A1(n4703), .A2(n4701), .A3(n4414), .ZN(n4700) );
  INV_X1 U6167 ( .A(n9512), .ZN(n4701) );
  NAND2_X1 U6168 ( .A1(n9506), .A2(n10066), .ZN(n4703) );
  NAND2_X1 U6169 ( .A1(n5259), .A2(n4705), .ZN(n9677) );
  NAND2_X1 U6170 ( .A1(n9677), .A2(n9335), .ZN(n5293) );
  NAND2_X1 U6171 ( .A1(n7753), .A2(n4707), .ZN(n7842) );
  MUX2_X1 U6172 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6629), .S(n6692), .Z(n6683)
         );
  XNOR2_X1 U6173 ( .A(n7935), .B(n7942), .ZN(n7650) );
  NAND2_X1 U6174 ( .A1(n4742), .A2(n8175), .ZN(n8176) );
  NAND2_X1 U6175 ( .A1(n4743), .A2(n8143), .ZN(n4742) );
  XNOR2_X1 U6176 ( .A(n4744), .B(n8865), .ZN(n4743) );
  OAI21_X1 U6177 ( .B1(n8726), .B2(n4751), .A(n4748), .ZN(n8700) );
  NAND3_X1 U6178 ( .A1(n4746), .A2(n8128), .A3(n4745), .ZN(n8679) );
  NAND3_X1 U6179 ( .A1(n4748), .A2(n4751), .A3(n4747), .ZN(n4745) );
  NAND3_X1 U6180 ( .A1(n8726), .A2(n4748), .A3(n4747), .ZN(n4746) );
  AOI21_X1 U6181 ( .B1(n4757), .B2(n4755), .A(n4754), .ZN(n4753) );
  NOR2_X1 U6182 ( .A1(n7172), .A2(n4761), .ZN(n4760) );
  NAND2_X1 U6183 ( .A1(n7574), .A2(n7722), .ZN(n4764) );
  NAND2_X1 U6184 ( .A1(n7807), .A2(n8106), .ZN(n4767) );
  AOI21_X1 U6185 ( .B1(n8823), .B2(n4771), .A(n4768), .ZN(n8759) );
  OR2_X1 U6186 ( .A1(n4394), .A2(n6548), .ZN(n5964) );
  OAI21_X1 U6187 ( .B1(n7152), .B2(n8147), .A(n7995), .ZN(n7099) );
  NAND2_X1 U6188 ( .A1(n7091), .A2(n7978), .ZN(n7152) );
  NAND3_X1 U6189 ( .A1(n5908), .A2(n6494), .A3(n8104), .ZN(n4777) );
  NAND2_X1 U6190 ( .A1(n8283), .A2(n4420), .ZN(n10144) );
  NAND2_X1 U6191 ( .A1(n8282), .A2(n5994), .ZN(n8283) );
  NAND2_X1 U6192 ( .A1(n10099), .A2(n6097), .ZN(n4782) );
  NAND2_X1 U6193 ( .A1(n4782), .A2(n4783), .ZN(n7119) );
  NAND2_X1 U6194 ( .A1(n4787), .A2(n4788), .ZN(n6226) );
  NAND2_X1 U6195 ( .A1(n7687), .A2(n4791), .ZN(n4787) );
  OAI21_X2 U6196 ( .B1(n8311), .B2(n4801), .A(n4799), .ZN(n7012) );
  NAND2_X1 U6197 ( .A1(n6242), .A2(n4804), .ZN(n4803) );
  NAND2_X1 U6198 ( .A1(n8190), .A2(n4448), .ZN(n4810) );
  OAI211_X1 U6199 ( .C1(n8190), .C2(n4812), .A(n4810), .B(n4461), .ZN(P2_U3222) );
  AOI21_X1 U6200 ( .B1(n8190), .B2(n6331), .A(n8191), .ZN(n8200) );
  XNOR2_X1 U6201 ( .A(n4824), .B(n5157), .ZN(n6562) );
  NAND3_X1 U6202 ( .A1(n8479), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4826) );
  NAND3_X1 U6203 ( .A1(n8388), .A2(n4954), .A3(n4953), .ZN(n4827) );
  NAND2_X1 U6204 ( .A1(n8709), .A2(n4830), .ZN(n4829) );
  NAND2_X1 U6205 ( .A1(n8774), .A2(n4835), .ZN(n4834) );
  NAND2_X1 U6206 ( .A1(n5023), .A2(n4842), .ZN(n4840) );
  INV_X1 U6207 ( .A(n5035), .ZN(n4839) );
  NAND3_X1 U6208 ( .A1(n4840), .A2(n5058), .A3(n4838), .ZN(n5043) );
  OAI21_X1 U6209 ( .B1(n5023), .B2(n4839), .A(n4841), .ZN(n5059) );
  AOI21_X1 U6210 ( .B1(n4844), .B2(n5035), .A(n4843), .ZN(n4841) );
  NAND2_X1 U6211 ( .A1(n5023), .A2(n5022), .ZN(n5036) );
  INV_X1 U6212 ( .A(n5039), .ZN(n4843) );
  INV_X1 U6213 ( .A(n8908), .ZN(n4848) );
  NAND3_X1 U6214 ( .A1(n4847), .A2(n4846), .A3(n4404), .ZN(P2_U3517) );
  NAND3_X1 U6215 ( .A1(n4849), .A2(n4459), .A3(n4850), .ZN(n4846) );
  OR2_X2 U6216 ( .A1(n8674), .A2(n8166), .ZN(n4849) );
  NAND3_X1 U6217 ( .A1(n4850), .A2(n4852), .A3(n4849), .ZN(n8909) );
  NAND2_X1 U6218 ( .A1(n8847), .A2(n4862), .ZN(n4860) );
  NAND2_X1 U6219 ( .A1(n10162), .A2(n7576), .ZN(n8026) );
  NAND2_X1 U6220 ( .A1(n8890), .A2(n4446), .ZN(n7170) );
  NAND2_X1 U6221 ( .A1(n4447), .A2(n7713), .ZN(n7799) );
  NAND2_X1 U6222 ( .A1(n6973), .A2(n6974), .ZN(n4873) );
  OR2_X1 U6223 ( .A1(n4944), .A2(n4945), .ZN(n4990) );
  NOR2_X1 U6224 ( .A1(n4945), .A2(n4943), .ZN(n4874) );
  INV_X1 U6225 ( .A(n5015), .ZN(n4876) );
  NAND2_X1 U6226 ( .A1(n4880), .A2(n7188), .ZN(n4879) );
  NAND2_X1 U6227 ( .A1(n4881), .A2(n4882), .ZN(n4880) );
  NAND2_X1 U6228 ( .A1(n5633), .A2(n4883), .ZN(n4881) );
  NAND2_X1 U6229 ( .A1(n7188), .A2(n5633), .ZN(n7283) );
  NAND2_X1 U6230 ( .A1(n5646), .A2(n4893), .ZN(n4892) );
  OAI21_X1 U6231 ( .B1(n8155), .B2(n7403), .A(n7973), .ZN(n7570) );
  NAND2_X1 U6232 ( .A1(n7353), .A2(n8014), .ZN(n7403) );
  AND2_X1 U6233 ( .A1(n8238), .A2(n8237), .ZN(n8268) );
  INV_X1 U6234 ( .A(n7411), .ZN(n7408) );
  CLKBUF_X1 U6235 ( .A(n6510), .Z(n6511) );
  AND2_X1 U6236 ( .A1(n8154), .A2(n7264), .ZN(n7348) );
  NAND2_X1 U6237 ( .A1(n7110), .A2(n7990), .ZN(n6906) );
  OR2_X1 U6238 ( .A1(n10248), .A2(n8912), .ZN(n8915) );
  INV_X1 U6239 ( .A(n10248), .ZN(n10215) );
  NAND2_X1 U6240 ( .A1(n6491), .A2(n6894), .ZN(n6492) );
  NAND2_X1 U6241 ( .A1(n8849), .A2(n8848), .ZN(n8847) );
  NAND2_X1 U6242 ( .A1(n5143), .A2(n4413), .ZN(n5145) );
  XNOR2_X1 U6243 ( .A(n5143), .B(n4413), .ZN(n6080) );
  AND2_X1 U6244 ( .A1(n7564), .A2(n10166), .ZN(n7565) );
  AOI21_X1 U6245 ( .B1(n6479), .B2(n6478), .A(n6477), .ZN(n6480) );
  NAND2_X2 U6246 ( .A1(n6083), .A2(n6082), .ZN(n7345) );
  INV_X1 U6247 ( .A(n7956), .ZN(n8179) );
  NAND2_X1 U6248 ( .A1(n7956), .A2(n8104), .ZN(n5908) );
  AND2_X1 U6249 ( .A1(n9120), .A2(n5794), .ZN(n5795) );
  INV_X1 U6250 ( .A(n9398), .ZN(n9411) );
  INV_X1 U6251 ( .A(n4944), .ZN(n9876) );
  OAI22_X1 U6252 ( .A1(n8788), .A2(n8210), .B1(n8292), .B2(n8792), .ZN(n8774)
         );
  NAND2_X2 U6253 ( .A1(n6503), .A2(n8888), .ZN(n8881) );
  OR2_X1 U6254 ( .A1(n6921), .A2(n6920), .ZN(n10273) );
  NOR2_X1 U6255 ( .A1(n7413), .A2(n7569), .ZN(n4909) );
  NAND2_X1 U6256 ( .A1(n9405), .A2(n4509), .ZN(n9284) );
  OR2_X1 U6257 ( .A1(n5575), .A2(n7129), .ZN(n10081) );
  INV_X2 U6258 ( .A(n10075), .ZN(n10076) );
  INV_X1 U6259 ( .A(n9405), .ZN(n9452) );
  OR2_X1 U6260 ( .A1(n9529), .A2(n9170), .ZN(n4910) );
  AND3_X1 U6261 ( .A1(n6468), .A2(n9160), .A3(n6467), .ZN(n4911) );
  OR2_X1 U6262 ( .A1(n5486), .A2(n9534), .ZN(n4912) );
  NOR2_X1 U6263 ( .A1(n5520), .A2(n9690), .ZN(n4913) );
  NOR2_X1 U6264 ( .A1(n5739), .A2(n5735), .ZN(n4914) );
  AND2_X1 U6265 ( .A1(n5541), .A2(n4938), .ZN(n4915) );
  AND2_X1 U6266 ( .A1(n6290), .A2(n8237), .ZN(n4916) );
  AND2_X1 U6267 ( .A1(n6240), .A2(n6239), .ZN(n4917) );
  AND2_X1 U6268 ( .A1(n5125), .A2(n5111), .ZN(n4918) );
  NOR2_X1 U6269 ( .A1(n5486), .A2(n9864), .ZN(n5571) );
  AND4_X1 U6270 ( .A1(n5303), .A2(n4937), .A3(n4936), .A4(n4935), .ZN(n4919)
         );
  OR2_X1 U6271 ( .A1(n9287), .A2(n9815), .ZN(n4920) );
  NAND2_X1 U6272 ( .A1(n9710), .A2(n5518), .ZN(n4921) );
  AND2_X1 U6273 ( .A1(n5829), .A2(n5830), .ZN(n4922) );
  INV_X1 U6274 ( .A(n8989), .ZN(n7717) );
  AND2_X1 U6275 ( .A1(n9030), .A2(n9817), .ZN(n4923) );
  INV_X1 U6276 ( .A(n7969), .ZN(n7573) );
  NAND2_X1 U6277 ( .A1(n5002), .A2(n5001), .ZN(n5020) );
  MUX2_X1 U6278 ( .A(n9247), .B(n9246), .S(n9284), .Z(n9248) );
  INV_X1 U6279 ( .A(n8132), .ZN(n8133) );
  AOI21_X1 U6280 ( .B1(n8134), .B2(n4467), .A(n8133), .ZN(n8135) );
  NAND2_X1 U6281 ( .A1(n4388), .A2(n5653), .ZN(n5599) );
  INV_X1 U6282 ( .A(n6215), .ZN(n5889) );
  INV_X1 U6283 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5860) );
  INV_X1 U6284 ( .A(n9225), .ZN(n5273) );
  INV_X1 U6285 ( .A(n9302), .ZN(n5490) );
  INV_X1 U6286 ( .A(n6137), .ZN(n5886) );
  NAND2_X1 U6287 ( .A1(n5889), .A2(n5888), .ZN(n6230) );
  INV_X1 U6288 ( .A(n6246), .ZN(n5890) );
  CLKBUF_X1 U6289 ( .A(n6492), .Z(n7988) );
  INV_X1 U6290 ( .A(n5135), .ZN(n5134) );
  NAND2_X1 U6291 ( .A1(n5601), .A2(n6460), .ZN(n5604) );
  INV_X1 U6292 ( .A(n5253), .ZN(n5252) );
  INV_X1 U6293 ( .A(n5352), .ZN(n5351) );
  OR2_X1 U6294 ( .A1(n5382), .A2(n9095), .ZN(n5403) );
  INV_X1 U6295 ( .A(n5287), .ZN(n5286) );
  NAND2_X1 U6296 ( .A1(n7699), .A2(n9318), .ZN(n7698) );
  INV_X1 U6297 ( .A(n6464), .ZN(n5486) );
  INV_X1 U6298 ( .A(SI_12_), .ZN(n8653) );
  INV_X1 U6299 ( .A(n5157), .ZN(n5160) );
  INV_X1 U6300 ( .A(n7554), .ZN(n6162) );
  AND2_X1 U6301 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n5884) );
  INV_X1 U6302 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U6303 ( .A1(n5886), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U6304 ( .A1(n8142), .A2(n8141), .ZN(n8143) );
  AND2_X1 U6305 ( .A1(n6336), .A2(n6317), .ZN(n8698) );
  NOR2_X1 U6306 ( .A1(n7348), .A2(n7347), .ZN(n7350) );
  NAND2_X1 U6307 ( .A1(n7990), .A2(n6492), .ZN(n6510) );
  NAND2_X1 U6308 ( .A1(n8702), .A2(n8877), .ZN(n8227) );
  OR2_X1 U6309 ( .A1(n6133), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U6310 ( .A1(n5064), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5086) );
  NAND2_X1 U6311 ( .A1(n5401), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U6312 ( .A1(n5351), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5369) );
  NAND2_X1 U6313 ( .A1(n5191), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5208) );
  INV_X1 U6314 ( .A(n5487), .ZN(n9526) );
  NAND2_X1 U6315 ( .A1(n5286), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5309) );
  NAND2_X1 U6316 ( .A1(n5149), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U6317 ( .A1(n9174), .A2(n9177), .ZN(n7235) );
  OR2_X1 U6318 ( .A1(n6414), .A2(n6413), .ZN(n6415) );
  INV_X1 U6319 ( .A(n5274), .ZN(n5278) );
  NOR2_X1 U6320 ( .A1(n5186), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5204) );
  INV_X1 U6321 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5187) );
  INV_X1 U6322 ( .A(n6291), .ZN(n6280) );
  AND2_X1 U6323 ( .A1(n6067), .A2(n5884), .ZN(n6084) );
  NOR2_X1 U6324 ( .A1(n6018), .A2(n6017), .ZN(n6037) );
  NAND2_X1 U6325 ( .A1(n8238), .A2(n4916), .ZN(n6296) );
  OR2_X1 U6326 ( .A1(n6284), .A2(n5912), .ZN(n5914) );
  INV_X1 U6327 ( .A(n7853), .ZN(n6241) );
  OR2_X1 U6328 ( .A1(n10098), .A2(n6812), .ZN(n8315) );
  AND2_X1 U6329 ( .A1(n6393), .A2(n6392), .ZN(n8241) );
  OR2_X1 U6330 ( .A1(n6387), .A2(n4398), .ZN(n6343) );
  OR2_X1 U6331 ( .A1(n6258), .A2(n8606), .ZN(n6269) );
  INV_X1 U6332 ( .A(n6624), .ZN(n6558) );
  AND2_X1 U6333 ( .A1(n8179), .A2(n8171), .ZN(n6624) );
  OR2_X1 U6334 ( .A1(n10248), .A2(n8865), .ZN(n6850) );
  AND2_X1 U6335 ( .A1(n6624), .A2(n8178), .ZN(n6918) );
  OR2_X1 U6336 ( .A1(n7412), .A2(n8150), .ZN(n7265) );
  OR2_X1 U6337 ( .A1(n6558), .A2(n6401), .ZN(n8858) );
  INV_X1 U6338 ( .A(n6918), .ZN(n6811) );
  OR2_X1 U6339 ( .A1(n5454), .A2(n5453), .ZN(n5479) );
  INV_X1 U6340 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7638) );
  INV_X1 U6341 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9054) );
  INV_X1 U6342 ( .A(n9327), .ZN(n6439) );
  INV_X1 U6343 ( .A(n9819), .ZN(n10015) );
  NAND2_X1 U6344 ( .A1(n5519), .A2(n4921), .ZN(n9690) );
  NAND2_X1 U6345 ( .A1(n10081), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5577) );
  INV_X1 U6346 ( .A(n10062), .ZN(n9818) );
  INV_X1 U6347 ( .A(n9637), .ZN(n10020) );
  INV_X1 U6348 ( .A(n6422), .ZN(n6423) );
  XNOR2_X1 U6349 ( .A(n5217), .B(SI_14_), .ZN(n5216) );
  NAND2_X1 U6350 ( .A1(n6084), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6121) );
  AND2_X1 U6351 ( .A1(n6037), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6067) );
  AND2_X1 U6352 ( .A1(n6388), .A2(n6500), .ZN(n8263) );
  AND2_X1 U6353 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6000) );
  AND2_X1 U6354 ( .A1(n8263), .A2(n10213), .ZN(n10136) );
  NAND2_X1 U6355 ( .A1(n6318), .A2(n5966), .ZN(n5971) );
  INV_X1 U6356 ( .A(n8377), .ZN(n8381) );
  INV_X1 U6357 ( .A(n8858), .ZN(n8879) );
  AND2_X1 U6358 ( .A1(n8109), .A2(n8108), .ZN(n8832) );
  NAND2_X1 U6359 ( .A1(n8881), .A2(n6506), .ZN(n8869) );
  OR3_X1 U6360 ( .A1(n6919), .A2(n6918), .A3(n10176), .ZN(n6920) );
  AND2_X1 U6361 ( .A1(n8917), .A2(n8916), .ZN(n8918) );
  NOR2_X1 U6362 ( .A1(n8806), .A2(n8805), .ZN(n8963) );
  AND2_X1 U6363 ( .A1(n7265), .A2(n7171), .ZN(n10233) );
  INV_X1 U6364 ( .A(n8993), .ZN(n10259) );
  AND2_X1 U6365 ( .A1(n6364), .A2(n7822), .ZN(n10175) );
  XNOR2_X1 U6366 ( .A(n6359), .B(P2_IR_REG_24__SCAN_IN), .ZN(n7592) );
  INV_X1 U6367 ( .A(n4958), .ZN(n6576) );
  INV_X1 U6368 ( .A(n9167), .ZN(n9139) );
  INV_X1 U6369 ( .A(n9092), .ZN(n9164) );
  AND2_X1 U6370 ( .A1(n5442), .A2(n5441), .ZN(n9546) );
  AND4_X1 U6371 ( .A1(n5292), .A2(n5291), .A3(n5290), .A4(n5289), .ZN(n9700)
         );
  OR2_X1 U6372 ( .A1(n6587), .A2(n6586), .ZN(n9491) );
  INV_X1 U6373 ( .A(n9492), .ZN(n9998) );
  INV_X1 U6374 ( .A(n9431), .ZN(n9530) );
  AND2_X1 U6375 ( .A1(n9336), .A2(n9249), .ZN(n9598) );
  INV_X1 U6376 ( .A(n9724), .ZN(n10006) );
  OAI22_X1 U6377 ( .A1(n4625), .A2(n9815), .B1(n10083), .B2(n6453), .ZN(n6454)
         );
  INV_X1 U6378 ( .A(n10051), .ZN(n7126) );
  NAND2_X1 U6379 ( .A1(n5080), .A2(n5079), .ZN(n5093) );
  INV_X1 U6380 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n9884) );
  NOR2_X1 U6381 ( .A1(n9898), .A2(n10310), .ZN(n9899) );
  INV_X1 U6382 ( .A(n8389), .ZN(n8350) );
  AND2_X1 U6383 ( .A1(n6391), .A2(n8182), .ZN(n10152) );
  INV_X1 U6384 ( .A(n10140), .ZN(n10095) );
  INV_X1 U6385 ( .A(n10136), .ZN(n8327) );
  INV_X1 U6386 ( .A(n8204), .ZN(n8702) );
  NAND2_X1 U6387 ( .A1(n8881), .A2(n6509), .ZN(n8874) );
  NOR2_X1 U6388 ( .A1(n10176), .A2(n10175), .ZN(n10184) );
  INV_X1 U6389 ( .A(n10184), .ZN(n10187) );
  INV_X1 U6390 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6761) );
  INV_X1 U6391 ( .A(n7603), .ZN(n7686) );
  NAND2_X1 U6392 ( .A1(n6469), .A2(n4911), .ZN(n6481) );
  INV_X1 U6393 ( .A(n9160), .ZN(n9144) );
  NAND2_X1 U6394 ( .A1(n5426), .A2(n5425), .ZN(n9560) );
  OR2_X1 U6395 ( .A1(n5313), .A2(n5312), .ZN(n9651) );
  INV_X1 U6396 ( .A(n10016), .ZN(n9464) );
  NAND2_X1 U6397 ( .A1(n9629), .A2(n7331), .ZN(n9706) );
  NAND2_X1 U6398 ( .A1(n10083), .A2(n9803), .ZN(n9815) );
  INV_X2 U6399 ( .A(n10081), .ZN(n10083) );
  INV_X1 U6400 ( .A(n9618), .ZN(n9846) );
  INV_X1 U6401 ( .A(n7846), .ZN(n9171) );
  OR2_X1 U6402 ( .A1(n5575), .A2(n9867), .ZN(n10075) );
  AND2_X1 U6403 ( .A1(n10051), .A2(n10040), .ZN(n10047) );
  INV_X1 U6404 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n8557) );
  INV_X1 U6405 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6565) );
  INV_X1 U6406 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6534) );
  NOR2_X1 U6407 ( .A1(n10312), .A2(n10311), .ZN(n10310) );
  NOR2_X1 U6408 ( .A1(n10303), .A2(n10302), .ZN(n10301) );
  INV_X1 U6409 ( .A(n9471), .ZN(P1_U4006) );
  NAND2_X1 U6410 ( .A1(n5574), .A2(n5573), .ZN(P1_U3519) );
  NAND2_X1 U6411 ( .A1(n4977), .A2(n4925), .ZN(n5015) );
  NAND2_X1 U6412 ( .A1(n5225), .A2(n5228), .ZN(n5247) );
  INV_X1 U6413 ( .A(n5247), .ZN(n4929) );
  NAND3_X1 U6414 ( .A1(n4929), .A2(n4928), .A3(n4927), .ZN(n4934) );
  NAND4_X1 U6415 ( .A1(n4932), .A2(n4931), .A3(n4930), .A4(n5280), .ZN(n4933)
         );
  NOR2_X1 U6416 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n4937) );
  NOR2_X1 U6417 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4936) );
  NOR2_X1 U6418 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n4935) );
  INV_X1 U6419 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4938) );
  INV_X1 U6420 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4939) );
  XNOR2_X2 U6421 ( .A(n4942), .B(P1_IR_REG_29__SCAN_IN), .ZN(n4945) );
  INV_X1 U6422 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7206) );
  OR2_X1 U6423 ( .A1(n5010), .A2(n7206), .ZN(n4948) );
  INV_X1 U6424 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n4943) );
  NAND3_X2 U6425 ( .A1(n4948), .A2(n4947), .A3(n4946), .ZN(n5597) );
  INV_X1 U6426 ( .A(n5597), .ZN(n6842) );
  INV_X1 U6427 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4952) );
  INV_X1 U6428 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4953) );
  AND2_X1 U6429 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n4955) );
  NAND2_X1 U6430 ( .A1(n4980), .A2(n4955), .ZN(n4969) );
  NAND2_X1 U6431 ( .A1(n4956), .A2(n4969), .ZN(n4983) );
  INV_X1 U6432 ( .A(SI_1_), .ZN(n4957) );
  MUX2_X1 U6433 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4391), .Z(n4981) );
  XNOR2_X1 U6434 ( .A(n4982), .B(n4981), .ZN(n6536) );
  OR2_X1 U6435 ( .A1(n4986), .A2(n6536), .ZN(n4963) );
  NAND2_X4 U6436 ( .A1(n4958), .A2(n4825), .ZN(n6428) );
  INV_X1 U6437 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6531) );
  INV_X1 U6438 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4960) );
  NAND2_X1 U6439 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4959) );
  OR2_X1 U6440 ( .A1(n4958), .A2(n6592), .ZN(n4961) );
  NAND2_X1 U6441 ( .A1(n6842), .A2(n4388), .ZN(n4971) );
  INV_X1 U6442 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6612) );
  NAND2_X1 U6443 ( .A1(n5009), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n4967) );
  INV_X1 U6444 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6884) );
  NAND2_X1 U6445 ( .A1(n4964), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n4965) );
  INV_X1 U6446 ( .A(SI_0_), .ZN(n5924) );
  INV_X1 U6447 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8622) );
  OAI21_X1 U6448 ( .B1(n4825), .B2(n5924), .A(n8622), .ZN(n4970) );
  AND2_X1 U6449 ( .A1(n4970), .A2(n4969), .ZN(n6527) );
  MUX2_X1 U6450 ( .A(P1_IR_REG_0__SCAN_IN), .B(n6527), .S(n4958), .Z(n10034)
         );
  INV_X1 U6451 ( .A(n10034), .ZN(n7205) );
  NOR2_X2 U6452 ( .A1(n5593), .A2(n7205), .ZN(n7199) );
  NAND2_X1 U6453 ( .A1(n5009), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4976) );
  INV_X1 U6454 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7135) );
  OR2_X1 U6455 ( .A1(n5010), .A2(n7135), .ZN(n4975) );
  INV_X1 U6456 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n4972) );
  OR2_X1 U6457 ( .A1(n5210), .A2(n6590), .ZN(n4973) );
  AND4_X2 U6458 ( .A1(n4976), .A2(n4975), .A3(n4974), .A4(n4973), .ZN(n7312)
         );
  INV_X1 U6459 ( .A(n7312), .ZN(n9470) );
  OR2_X1 U6460 ( .A1(n4977), .A2(n5187), .ZN(n4979) );
  INV_X1 U6461 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4978) );
  NAND2_X1 U6462 ( .A1(n4979), .A2(n4978), .ZN(n5003) );
  OAI21_X1 U6463 ( .B1(n4979), .B2(n4978), .A(n5003), .ZN(n6957) );
  INV_X1 U6464 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6529) );
  OR2_X1 U6465 ( .A1(n6428), .A2(n6529), .ZN(n4988) );
  INV_X1 U6466 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6540) );
  MUX2_X1 U6467 ( .A(n6540), .B(n6529), .S(n4980), .Z(n4999) );
  XNOR2_X1 U6468 ( .A(n4999), .B(SI_2_), .ZN(n4997) );
  NAND2_X1 U6469 ( .A1(n4982), .A2(n4981), .ZN(n4985) );
  NAND2_X1 U6470 ( .A1(n4983), .A2(SI_1_), .ZN(n4984) );
  NAND2_X1 U6471 ( .A1(n4985), .A2(n4984), .ZN(n4998) );
  XNOR2_X1 U6472 ( .A(n4997), .B(n4998), .ZN(n6541) );
  OR2_X1 U6473 ( .A1(n4986), .A2(n6541), .ZN(n4987) );
  OAI211_X1 U6474 ( .C1(n4958), .C2(n6957), .A(n4988), .B(n4987), .ZN(n6998)
         );
  NAND2_X1 U6475 ( .A1(n9470), .A2(n5607), .ZN(n9415) );
  NAND2_X1 U6476 ( .A1(n7312), .A2(n6998), .ZN(n9414) );
  NAND2_X1 U6477 ( .A1(n7003), .A2(n9302), .ZN(n4989) );
  NAND2_X1 U6478 ( .A1(n4989), .A2(n9414), .ZN(n7309) );
  NAND2_X1 U6479 ( .A1(n5009), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4996) );
  INV_X1 U6480 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n4991) );
  OR2_X1 U6481 ( .A1(n4990), .A2(n4991), .ZN(n4995) );
  INV_X1 U6482 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n4992) );
  OR2_X1 U6483 ( .A1(n5210), .A2(n4992), .ZN(n4994) );
  OR2_X1 U6484 ( .A1(n5010), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n4993) );
  NAND2_X1 U6485 ( .A1(n4998), .A2(n4997), .ZN(n5002) );
  INV_X1 U6486 ( .A(n4999), .ZN(n5000) );
  NAND2_X1 U6487 ( .A1(n5000), .A2(SI_2_), .ZN(n5001) );
  MUX2_X1 U6488 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n4391), .Z(n5021) );
  INV_X1 U6489 ( .A(SI_3_), .ZN(n8636) );
  XNOR2_X1 U6490 ( .A(n5021), .B(n8636), .ZN(n5019) );
  XNOR2_X1 U6491 ( .A(n5020), .B(n5019), .ZN(n6549) );
  OR2_X1 U6492 ( .A1(n4986), .A2(n6549), .ZN(n5008) );
  INV_X1 U6493 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6532) );
  OR2_X1 U6494 ( .A1(n6428), .A2(n6532), .ZN(n5007) );
  NAND2_X1 U6495 ( .A1(n5003), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5005) );
  INV_X1 U6496 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5004) );
  XNOR2_X1 U6497 ( .A(n5005), .B(n5004), .ZN(n6789) );
  OR2_X1 U6498 ( .A1(n4958), .A2(n6789), .ZN(n5006) );
  XNOR2_X1 U6499 ( .A(n9469), .B(n10057), .ZN(n9304) );
  INV_X1 U6500 ( .A(n9304), .ZN(n7311) );
  INV_X1 U6501 ( .A(n9469), .ZN(n7372) );
  INV_X1 U6502 ( .A(n10057), .ZN(n7321) );
  NAND2_X1 U6503 ( .A1(n7372), .A2(n7321), .ZN(n9373) );
  NAND2_X1 U6504 ( .A1(n6445), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5014) );
  INV_X1 U6505 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6598) );
  OR2_X1 U6506 ( .A1(n5210), .A2(n6598), .ZN(n5013) );
  INV_X1 U6507 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6582) );
  OR2_X1 U6508 ( .A1(n5460), .A2(n6582), .ZN(n5012) );
  XNOR2_X1 U6509 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7369) );
  OR2_X1 U6510 ( .A1(n5010), .A2(n7369), .ZN(n5011) );
  INV_X1 U6511 ( .A(n7389), .ZN(n9468) );
  NAND2_X1 U6512 ( .A1(n5015), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5016) );
  MUX2_X1 U6513 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5016), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5018) );
  NAND2_X1 U6514 ( .A1(n5018), .A2(n5017), .ZN(n6597) );
  INV_X1 U6515 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6530) );
  OR2_X1 U6516 ( .A1(n6428), .A2(n6530), .ZN(n5025) );
  NAND2_X1 U6517 ( .A1(n5021), .A2(SI_3_), .ZN(n5022) );
  INV_X1 U6518 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6538) );
  MUX2_X1 U6519 ( .A(n6538), .B(n6530), .S(n4391), .Z(n5037) );
  XNOR2_X1 U6520 ( .A(n5036), .B(n5035), .ZN(n6539) );
  OR2_X1 U6521 ( .A1(n4986), .A2(n6539), .ZN(n5024) );
  OAI211_X1 U6522 ( .C1(n4958), .C2(n6597), .A(n5025), .B(n5024), .ZN(n7371)
         );
  INV_X1 U6523 ( .A(n7371), .ZN(n7056) );
  NAND2_X1 U6524 ( .A1(n9468), .A2(n7056), .ZN(n9379) );
  NAND2_X1 U6525 ( .A1(n9172), .A2(n9379), .ZN(n9173) );
  NAND2_X1 U6526 ( .A1(n7389), .A2(n7371), .ZN(n9176) );
  NAND2_X1 U6527 ( .A1(n9173), .A2(n9176), .ZN(n7234) );
  NAND2_X1 U6528 ( .A1(n6445), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5032) );
  INV_X1 U6529 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6775) );
  OR2_X1 U6530 ( .A1(n5460), .A2(n6775), .ZN(n5031) );
  INV_X1 U6531 ( .A(n5051), .ZN(n5026) );
  INV_X1 U6532 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n8449) );
  NAND2_X1 U6533 ( .A1(n5051), .A2(n8449), .ZN(n5027) );
  NAND2_X1 U6534 ( .A1(n5066), .A2(n5027), .ZN(n7464) );
  OR2_X1 U6535 ( .A1(n5010), .A2(n7464), .ZN(n5030) );
  INV_X1 U6536 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5028) );
  OR2_X1 U6537 ( .A1(n5210), .A2(n5028), .ZN(n5029) );
  OR2_X1 U6538 ( .A1(n5033), .A2(n5187), .ZN(n5034) );
  XNOR2_X1 U6539 ( .A(n5034), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6776) );
  INV_X1 U6540 ( .A(n6776), .ZN(n6802) );
  INV_X1 U6541 ( .A(n5037), .ZN(n5038) );
  NAND2_X1 U6542 ( .A1(n5038), .A2(SI_4_), .ZN(n5039) );
  INV_X1 U6543 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6546) );
  INV_X1 U6544 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6533) );
  MUX2_X1 U6545 ( .A(n6546), .B(n6533), .S(n5868), .Z(n5040) );
  INV_X1 U6546 ( .A(n5040), .ZN(n5041) );
  NAND2_X1 U6547 ( .A1(n5041), .A2(SI_5_), .ZN(n5042) );
  NAND2_X1 U6548 ( .A1(n5043), .A2(n5042), .ZN(n5076) );
  INV_X1 U6549 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6544) );
  MUX2_X1 U6550 ( .A(n6544), .B(n6534), .S(n5868), .Z(n5077) );
  XNOR2_X1 U6551 ( .A(n5077), .B(SI_6_), .ZN(n5075) );
  XNOR2_X1 U6552 ( .A(n5076), .B(n5075), .ZN(n6545) );
  OR2_X1 U6553 ( .A1(n4986), .A2(n6545), .ZN(n5045) );
  OR2_X1 U6554 ( .A1(n6428), .A2(n6534), .ZN(n5044) );
  OAI211_X1 U6555 ( .C1(n4958), .C2(n6802), .A(n5045), .B(n5044), .ZN(n5635)
         );
  NAND2_X1 U6556 ( .A1(n10063), .A2(n5635), .ZN(n9188) );
  NAND2_X1 U6557 ( .A1(n5009), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5056) );
  INV_X1 U6558 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5046) );
  OR2_X1 U6559 ( .A1(n5210), .A2(n5046), .ZN(n5055) );
  INV_X1 U6560 ( .A(n5047), .ZN(n5049) );
  INV_X1 U6561 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5048) );
  NAND2_X1 U6562 ( .A1(n5049), .A2(n5048), .ZN(n5050) );
  NAND2_X1 U6563 ( .A1(n5051), .A2(n5050), .ZN(n7395) );
  OR2_X1 U6564 ( .A1(n5010), .A2(n7395), .ZN(n5054) );
  INV_X1 U6565 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5052) );
  OR2_X1 U6566 ( .A1(n4990), .A2(n5052), .ZN(n5053) );
  NAND2_X1 U6567 ( .A1(n5017), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5057) );
  XNOR2_X1 U6568 ( .A(n5057), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6774) );
  INV_X1 U6569 ( .A(n6774), .ZN(n6589) );
  XNOR2_X1 U6570 ( .A(n5059), .B(n5058), .ZN(n6547) );
  OR2_X1 U6571 ( .A1(n4986), .A2(n6547), .ZN(n5061) );
  OR2_X1 U6572 ( .A1(n6428), .A2(n6533), .ZN(n5060) );
  OAI211_X1 U6573 ( .C1(n4958), .C2(n6589), .A(n5061), .B(n5060), .ZN(n7394)
         );
  NAND2_X1 U6574 ( .A1(n7373), .A2(n7394), .ZN(n9177) );
  NAND2_X1 U6575 ( .A1(n9188), .A2(n9177), .ZN(n9377) );
  INV_X1 U6576 ( .A(n7394), .ZN(n10061) );
  NAND2_X1 U6577 ( .A1(n9467), .A2(n10061), .ZN(n9174) );
  INV_X1 U6578 ( .A(n9174), .ZN(n9178) );
  NAND2_X1 U6579 ( .A1(n9188), .A2(n9178), .ZN(n5062) );
  INV_X1 U6580 ( .A(n10063), .ZN(n9466) );
  NAND2_X1 U6581 ( .A1(n9466), .A2(n7469), .ZN(n9300) );
  AND2_X1 U6582 ( .A1(n5062), .A2(n9300), .ZN(n9419) );
  INV_X1 U6583 ( .A(n7327), .ZN(n5083) );
  NAND2_X1 U6584 ( .A1(n5009), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5072) );
  INV_X1 U6585 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5063) );
  OR2_X1 U6586 ( .A1(n5210), .A2(n5063), .ZN(n5071) );
  INV_X1 U6587 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5065) );
  NAND2_X1 U6588 ( .A1(n5066), .A2(n5065), .ZN(n5067) );
  NAND2_X1 U6589 ( .A1(n5086), .A2(n5067), .ZN(n7458) );
  OR2_X1 U6590 ( .A1(n5010), .A2(n7458), .ZN(n5070) );
  INV_X1 U6591 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5068) );
  OR2_X1 U6592 ( .A1(n4990), .A2(n5068), .ZN(n5069) );
  NAND2_X1 U6593 ( .A1(n5073), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5074) );
  XNOR2_X1 U6594 ( .A(n5074), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9933) );
  INV_X1 U6595 ( .A(n9933), .ZN(n6772) );
  NAND2_X1 U6596 ( .A1(n5076), .A2(n5075), .ZN(n5080) );
  INV_X1 U6597 ( .A(n5077), .ZN(n5078) );
  NAND2_X1 U6598 ( .A1(n5078), .A2(SI_6_), .ZN(n5079) );
  MUX2_X1 U6599 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5868), .Z(n5094) );
  XNOR2_X1 U6600 ( .A(n5094), .B(n8589), .ZN(n5092) );
  XNOR2_X1 U6601 ( .A(n5093), .B(n5092), .ZN(n6543) );
  OR2_X1 U6602 ( .A1(n6543), .A2(n4986), .ZN(n5082) );
  INV_X1 U6603 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6535) );
  OR2_X1 U6604 ( .A1(n6428), .A2(n6535), .ZN(n5081) );
  OAI211_X1 U6605 ( .C1(n4958), .C2(n6772), .A(n5082), .B(n5081), .ZN(n7448)
         );
  NAND2_X1 U6606 ( .A1(n7483), .A2(n7448), .ZN(n9187) );
  INV_X1 U6607 ( .A(n7483), .ZN(n9465) );
  NAND2_X1 U6608 ( .A1(n9465), .A2(n7462), .ZN(n9418) );
  NAND2_X1 U6609 ( .A1(n9187), .A2(n9418), .ZN(n9309) );
  NAND2_X1 U6610 ( .A1(n6445), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5091) );
  INV_X1 U6611 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5084) );
  OR2_X1 U6612 ( .A1(n5210), .A2(n5084), .ZN(n5090) );
  INV_X1 U6613 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5085) );
  OR2_X1 U6614 ( .A1(n5460), .A2(n5085), .ZN(n5089) );
  NAND2_X1 U6615 ( .A1(n5086), .A2(n7638), .ZN(n5087) );
  NAND2_X1 U6616 ( .A1(n5117), .A2(n5087), .ZN(n7640) );
  OR2_X1 U6617 ( .A1(n5010), .A2(n7640), .ZN(n5088) );
  NAND2_X1 U6618 ( .A1(n5093), .A2(n5092), .ZN(n5096) );
  NAND2_X1 U6619 ( .A1(n5094), .A2(SI_7_), .ZN(n5095) );
  MUX2_X1 U6620 ( .A(n8529), .B(n6551), .S(n5868), .Z(n5098) );
  INV_X1 U6621 ( .A(SI_8_), .ZN(n5097) );
  INV_X1 U6622 ( .A(n5098), .ZN(n5099) );
  NAND2_X1 U6623 ( .A1(n5099), .A2(SI_8_), .ZN(n5100) );
  NAND2_X1 U6624 ( .A1(n5107), .A2(n5100), .ZN(n5105) );
  XNOR2_X1 U6625 ( .A(n5106), .B(n5105), .ZN(n6550) );
  NAND2_X1 U6626 ( .A1(n6550), .A2(n5164), .ZN(n5104) );
  NAND2_X1 U6627 ( .A1(n5112), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5102) );
  XNOR2_X1 U6628 ( .A(n5102), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9946) );
  AOI22_X1 U6629 ( .A1(n5306), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6576), .B2(
        n9946), .ZN(n5103) );
  NAND2_X1 U6630 ( .A1(n10016), .A2(n7496), .ZN(n9192) );
  MUX2_X1 U6631 ( .A(n8604), .B(n6555), .S(n5868), .Z(n5109) );
  INV_X1 U6632 ( .A(SI_9_), .ZN(n5108) );
  NAND2_X1 U6633 ( .A1(n5109), .A2(n5108), .ZN(n5125) );
  INV_X1 U6634 ( .A(n5109), .ZN(n5110) );
  NAND2_X1 U6635 ( .A1(n5110), .A2(SI_9_), .ZN(n5111) );
  XNOR2_X2 U6636 ( .A(n5124), .B(n4918), .ZN(n6553) );
  NAND2_X1 U6637 ( .A1(n6553), .A2(n5164), .ZN(n5116) );
  OR2_X1 U6638 ( .A1(n5465), .A2(n5187), .ZN(n5113) );
  MUX2_X1 U6639 ( .A(n5113), .B(P1_IR_REG_31__SCAN_IN), .S(n8525), .Z(n5114)
         );
  NAND2_X1 U6640 ( .A1(n5465), .A2(n8525), .ZN(n5304) );
  NAND2_X1 U6641 ( .A1(n5114), .A2(n5304), .ZN(n6863) );
  INV_X1 U6642 ( .A(n6863), .ZN(n6872) );
  AOI22_X1 U6643 ( .A1(n5306), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6576), .B2(
        n6872), .ZN(n5115) );
  NAND2_X1 U6644 ( .A1(n5009), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5123) );
  INV_X1 U6645 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6862) );
  OR2_X1 U6646 ( .A1(n5210), .A2(n6862), .ZN(n5122) );
  NAND2_X1 U6647 ( .A1(n5117), .A2(n6767), .ZN(n5118) );
  NAND2_X1 U6648 ( .A1(n5135), .A2(n5118), .ZN(n10009) );
  OR2_X1 U6649 ( .A1(n5010), .A2(n10009), .ZN(n5121) );
  INV_X1 U6650 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5119) );
  OR2_X1 U6651 ( .A1(n4990), .A2(n5119), .ZN(n5120) );
  NAND4_X1 U6652 ( .A1(n5123), .A2(n5122), .A3(n5121), .A4(n5120), .ZN(n9463)
         );
  INV_X1 U6653 ( .A(n9463), .ZN(n7639) );
  OR2_X1 U6654 ( .A1(n10027), .A2(n7639), .ZN(n9308) );
  INV_X1 U6655 ( .A(n7496), .ZN(n7644) );
  NAND2_X1 U6656 ( .A1(n9464), .A2(n7644), .ZN(n10011) );
  AND2_X1 U6657 ( .A1(n9308), .A2(n10011), .ZN(n9347) );
  NAND2_X1 U6658 ( .A1(n10012), .A2(n9347), .ZN(n7522) );
  MUX2_X1 U6659 ( .A(n6561), .B(n6565), .S(n5868), .Z(n5127) );
  INV_X1 U6660 ( .A(SI_10_), .ZN(n5126) );
  NAND2_X1 U6661 ( .A1(n5127), .A2(n5126), .ZN(n5144) );
  INV_X1 U6662 ( .A(n5127), .ZN(n5128) );
  NAND2_X1 U6663 ( .A1(n5128), .A2(SI_10_), .ZN(n5129) );
  NAND2_X1 U6664 ( .A1(n5130), .A2(n5164), .ZN(n5133) );
  NAND2_X1 U6665 ( .A1(n5304), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5131) );
  XNOR2_X1 U6666 ( .A(n5131), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7220) );
  AOI22_X1 U6667 ( .A1(n5306), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6576), .B2(
        n7220), .ZN(n5132) );
  NAND2_X1 U6668 ( .A1(n5009), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5141) );
  INV_X1 U6669 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6868) );
  NAND2_X1 U6670 ( .A1(n5135), .A2(n6868), .ZN(n5136) );
  NAND2_X1 U6671 ( .A1(n5151), .A2(n5136), .ZN(n7681) );
  OR2_X1 U6672 ( .A1(n5010), .A2(n7681), .ZN(n5140) );
  INV_X1 U6673 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5137) );
  OR2_X1 U6674 ( .A1(n4990), .A2(n5137), .ZN(n5139) );
  INV_X1 U6675 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6861) );
  OR2_X1 U6676 ( .A1(n5210), .A2(n6861), .ZN(n5138) );
  NAND2_X1 U6677 ( .A1(n7603), .A2(n10017), .ZN(n9195) );
  NAND2_X1 U6678 ( .A1(n10027), .A2(n7639), .ZN(n9307) );
  AND2_X1 U6679 ( .A1(n9195), .A2(n9307), .ZN(n9344) );
  NAND2_X1 U6680 ( .A1(n7522), .A2(n9344), .ZN(n5142) );
  MUX2_X1 U6681 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n5868), .Z(n5158) );
  NAND2_X1 U6682 ( .A1(n6562), .A2(n5164), .ZN(n5148) );
  NAND2_X1 U6683 ( .A1(n5165), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5146) );
  XNOR2_X1 U6684 ( .A(n5146), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9958) );
  AOI22_X1 U6685 ( .A1(n5306), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6576), .B2(
        n9958), .ZN(n5147) );
  NAND2_X1 U6686 ( .A1(n6445), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5156) );
  INV_X1 U6687 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7661) );
  OR2_X1 U6688 ( .A1(n5460), .A2(n7661), .ZN(n5155) );
  OR2_X1 U6689 ( .A1(n5210), .A2(n9915), .ZN(n5154) );
  INV_X1 U6690 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5150) );
  NAND2_X1 U6691 ( .A1(n5151), .A2(n5150), .ZN(n5152) );
  NAND2_X1 U6692 ( .A1(n5170), .A2(n5152), .ZN(n7792) );
  OR2_X1 U6693 ( .A1(n5010), .A2(n7792), .ZN(n5153) );
  NAND2_X1 U6694 ( .A1(n7794), .A2(n7746), .ZN(n9202) );
  NAND2_X1 U6695 ( .A1(n7668), .A2(n9202), .ZN(n7736) );
  NAND2_X1 U6696 ( .A1(n5158), .A2(SI_11_), .ZN(n5159) );
  MUX2_X1 U6697 ( .A(n6611), .B(n6609), .S(n5868), .Z(n5161) );
  INV_X1 U6698 ( .A(n5161), .ZN(n5162) );
  NAND2_X1 U6699 ( .A1(n5162), .A2(SI_12_), .ZN(n5163) );
  NAND2_X1 U6700 ( .A1(n5178), .A2(n5163), .ZN(n5179) );
  XNOR2_X1 U6701 ( .A(n5180), .B(n5179), .ZN(n6113) );
  NAND2_X1 U6702 ( .A1(n6113), .A2(n5164), .ZN(n5168) );
  NAND2_X1 U6703 ( .A1(n5186), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5166) );
  XNOR2_X1 U6704 ( .A(n5166), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9976) );
  AOI22_X1 U6705 ( .A1(n5306), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6576), .B2(
        n9976), .ZN(n5167) );
  NAND2_X1 U6706 ( .A1(n5009), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5176) );
  INV_X1 U6707 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5169) );
  OR2_X1 U6708 ( .A1(n5210), .A2(n5169), .ZN(n5175) );
  NAND2_X1 U6709 ( .A1(n5170), .A2(n9054), .ZN(n5171) );
  NAND2_X1 U6710 ( .A1(n5193), .A2(n5171), .ZN(n9056) );
  OR2_X1 U6711 ( .A1(n5010), .A2(n9056), .ZN(n5174) );
  INV_X1 U6712 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5172) );
  OR2_X1 U6713 ( .A1(n4990), .A2(n5172), .ZN(n5173) );
  OR2_X1 U6714 ( .A1(n9058), .A2(n9113), .ZN(n9203) );
  OR2_X1 U6715 ( .A1(n7794), .A2(n7746), .ZN(n7735) );
  AND2_X1 U6716 ( .A1(n9203), .A2(n7735), .ZN(n9212) );
  NAND2_X1 U6717 ( .A1(n7736), .A2(n9212), .ZN(n5177) );
  NAND2_X1 U6718 ( .A1(n9058), .A2(n9113), .ZN(n9210) );
  NAND2_X1 U6719 ( .A1(n5177), .A2(n9210), .ZN(n7699) );
  INV_X1 U6720 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5181) );
  MUX2_X1 U6721 ( .A(n6745), .B(n5181), .S(n5868), .Z(n5183) );
  INV_X1 U6722 ( .A(SI_13_), .ZN(n5182) );
  INV_X1 U6723 ( .A(n5183), .ZN(n5184) );
  NAND2_X1 U6724 ( .A1(n5184), .A2(SI_13_), .ZN(n5185) );
  XNOR2_X1 U6725 ( .A(n5200), .B(n5199), .ZN(n6743) );
  NAND2_X1 U6726 ( .A1(n6743), .A2(n5164), .ZN(n5190) );
  OR2_X1 U6727 ( .A1(n5204), .A2(n5187), .ZN(n5188) );
  XNOR2_X1 U6728 ( .A(n5188), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7544) );
  AOI22_X1 U6729 ( .A1(n5306), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6576), .B2(
        n7544), .ZN(n5189) );
  NAND2_X1 U6730 ( .A1(n6445), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5198) );
  INV_X1 U6731 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7213) );
  OR2_X1 U6732 ( .A1(n5210), .A2(n7213), .ZN(n5197) );
  INV_X1 U6733 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7702) );
  OR2_X1 U6734 ( .A1(n5460), .A2(n7702), .ZN(n5196) );
  INV_X1 U6735 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6736 ( .A1(n5193), .A2(n5192), .ZN(n5194) );
  NAND2_X1 U6737 ( .A1(n5208), .A2(n5194), .ZN(n9112) );
  OR2_X1 U6738 ( .A1(n5010), .A2(n9112), .ZN(n5195) );
  NAND4_X1 U6739 ( .A1(n5198), .A2(n5197), .A3(n5196), .A4(n5195), .ZN(n9460)
         );
  INV_X1 U6740 ( .A(n9460), .ZN(n9055) );
  OR2_X1 U6741 ( .A1(n9816), .A2(n9055), .ZN(n9206) );
  NAND2_X1 U6742 ( .A1(n9816), .A2(n9055), .ZN(n9343) );
  MUX2_X1 U6743 ( .A(n6761), .B(n8436), .S(n5868), .Z(n5217) );
  XNOR2_X1 U6744 ( .A(n5220), .B(n5216), .ZN(n6760) );
  NAND2_X1 U6745 ( .A1(n6760), .A2(n5164), .ZN(n5206) );
  INV_X1 U6746 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5203) );
  NAND2_X1 U6747 ( .A1(n5204), .A2(n5203), .ZN(n5248) );
  NAND2_X1 U6748 ( .A1(n5248), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5226) );
  XNOR2_X1 U6749 ( .A(n5226), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7653) );
  AOI22_X1 U6750 ( .A1(n5306), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7653), .B2(
        n6576), .ZN(n5205) );
  NAND2_X1 U6751 ( .A1(n6445), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5214) );
  INV_X1 U6752 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7763) );
  OR2_X1 U6753 ( .A1(n5460), .A2(n7763), .ZN(n5213) );
  INV_X1 U6754 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7541) );
  NAND2_X1 U6755 ( .A1(n5208), .A2(n7541), .ZN(n5209) );
  NAND2_X1 U6756 ( .A1(n5234), .A2(n5209), .ZN(n9027) );
  OR2_X1 U6757 ( .A1(n5010), .A2(n9027), .ZN(n5212) );
  INV_X1 U6758 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7537) );
  OR2_X1 U6759 ( .A1(n5210), .A2(n7537), .ZN(n5211) );
  NAND4_X1 U6760 ( .A1(n5214), .A2(n5213), .A3(n5212), .A4(n5211), .ZN(n9817)
         );
  INV_X1 U6761 ( .A(n9817), .ZN(n7703) );
  OR2_X1 U6762 ( .A1(n9030), .A2(n7703), .ZN(n9218) );
  NAND2_X1 U6763 ( .A1(n9030), .A2(n7703), .ZN(n9352) );
  NAND2_X1 U6764 ( .A1(n9218), .A2(n9352), .ZN(n7760) );
  INV_X1 U6765 ( .A(n9343), .ZN(n9217) );
  NOR2_X1 U6766 ( .A1(n7760), .A2(n9217), .ZN(n5215) );
  INV_X1 U6767 ( .A(n5217), .ZN(n5218) );
  NAND2_X1 U6768 ( .A1(n5218), .A2(SI_14_), .ZN(n5219) );
  MUX2_X1 U6769 ( .A(n8464), .B(n8557), .S(n5868), .Z(n5222) );
  INV_X1 U6770 ( .A(SI_15_), .ZN(n5221) );
  INV_X1 U6771 ( .A(n5222), .ZN(n5223) );
  NAND2_X1 U6772 ( .A1(n5223), .A2(SI_15_), .ZN(n5224) );
  XNOR2_X1 U6773 ( .A(n5242), .B(n5241), .ZN(n6940) );
  NAND2_X1 U6774 ( .A1(n6940), .A2(n5164), .ZN(n5232) );
  NAND2_X1 U6775 ( .A1(n5226), .A2(n5225), .ZN(n5227) );
  NAND2_X1 U6776 ( .A1(n5227), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5229) );
  XNOR2_X1 U6777 ( .A(n5229), .B(n5228), .ZN(n7942) );
  OAI22_X1 U6778 ( .A1(n7942), .A2(n4958), .B1(n6428), .B2(n8557), .ZN(n5230)
         );
  INV_X1 U6779 ( .A(n5230), .ZN(n5231) );
  NAND2_X1 U6780 ( .A1(n6445), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5239) );
  OR2_X1 U6781 ( .A1(n5460), .A2(n7649), .ZN(n5238) );
  INV_X1 U6782 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7931) );
  OR2_X1 U6783 ( .A1(n5210), .A2(n7931), .ZN(n5237) );
  INV_X1 U6784 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5233) );
  NAND2_X1 U6785 ( .A1(n5234), .A2(n5233), .ZN(n5235) );
  NAND2_X1 U6786 ( .A1(n5253), .A2(n5235), .ZN(n9163) );
  OR2_X1 U6787 ( .A1(n5010), .A2(n9163), .ZN(n5236) );
  OR2_X1 U6788 ( .A1(n7846), .A2(n9074), .ZN(n9355) );
  NAND2_X1 U6789 ( .A1(n7846), .A2(n9074), .ZN(n9353) );
  NAND2_X1 U6790 ( .A1(n9355), .A2(n9353), .ZN(n9709) );
  NAND2_X1 U6791 ( .A1(n7842), .A2(n9353), .ZN(n9707) );
  MUX2_X1 U6792 ( .A(n6950), .B(n8634), .S(n5868), .Z(n5244) );
  INV_X1 U6793 ( .A(SI_16_), .ZN(n5243) );
  NAND2_X1 U6794 ( .A1(n5244), .A2(n5243), .ZN(n5262) );
  INV_X1 U6795 ( .A(n5244), .ZN(n5245) );
  NAND2_X1 U6796 ( .A1(n5245), .A2(SI_16_), .ZN(n5246) );
  XNOR2_X1 U6797 ( .A(n5261), .B(n5260), .ZN(n6942) );
  NAND2_X1 U6798 ( .A1(n6942), .A2(n5164), .ZN(n5251) );
  OR2_X1 U6799 ( .A1(n5248), .A2(n5247), .ZN(n5264) );
  NAND2_X1 U6800 ( .A1(n5264), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5249) );
  XNOR2_X1 U6801 ( .A(n5249), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9477) );
  AOI22_X1 U6802 ( .A1(n6576), .A2(n9477), .B1(n5306), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n5250) );
  NAND2_X1 U6803 ( .A1(n6445), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5258) );
  INV_X1 U6804 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9716) );
  OR2_X1 U6805 ( .A1(n5460), .A2(n9716), .ZN(n5257) );
  INV_X1 U6806 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9073) );
  NAND2_X1 U6807 ( .A1(n5253), .A2(n9073), .ZN(n5254) );
  NAND2_X1 U6808 ( .A1(n5267), .A2(n5254), .ZN(n9715) );
  OR2_X1 U6809 ( .A1(n5010), .A2(n9715), .ZN(n5256) );
  INV_X1 U6810 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9813) );
  OR2_X1 U6811 ( .A1(n5210), .A2(n9813), .ZN(n5255) );
  OR2_X1 U6812 ( .A1(n9727), .A2(n9699), .ZN(n9354) );
  NAND2_X1 U6813 ( .A1(n9727), .A2(n9699), .ZN(n9369) );
  NAND2_X1 U6814 ( .A1(n9354), .A2(n9369), .ZN(n9708) );
  INV_X1 U6815 ( .A(n9708), .ZN(n9712) );
  NAND2_X1 U6816 ( .A1(n9707), .A2(n9712), .ZN(n5259) );
  INV_X1 U6817 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5263) );
  MUX2_X1 U6818 ( .A(n6979), .B(n5263), .S(n5868), .Z(n5275) );
  XNOR2_X1 U6819 ( .A(n5275), .B(SI_17_), .ZN(n5274) );
  XNOR2_X1 U6820 ( .A(n5279), .B(n5274), .ZN(n6952) );
  NAND2_X1 U6821 ( .A1(n6952), .A2(n5164), .ZN(n5266) );
  OAI21_X1 U6822 ( .B1(n5264), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5281) );
  XNOR2_X1 U6823 ( .A(n5281), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9487) );
  AOI22_X1 U6824 ( .A1(n9487), .A2(n6576), .B1(n5306), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n5265) );
  NAND2_X1 U6825 ( .A1(n5009), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5272) );
  INV_X1 U6826 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n8539) );
  OR2_X1 U6827 ( .A1(n4990), .A2(n8539), .ZN(n5271) );
  INV_X1 U6828 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9083) );
  NAND2_X1 U6829 ( .A1(n5267), .A2(n9083), .ZN(n5268) );
  NAND2_X1 U6830 ( .A1(n5287), .A2(n5268), .ZN(n9693) );
  OR2_X1 U6831 ( .A1(n5010), .A2(n9693), .ZN(n5270) );
  INV_X1 U6832 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n8462) );
  OR2_X1 U6833 ( .A1(n5210), .A2(n8462), .ZN(n5269) );
  NAND4_X1 U6834 ( .A1(n5272), .A2(n5271), .A3(n5270), .A4(n5269), .ZN(n9806)
         );
  AND2_X1 U6835 ( .A1(n9802), .A2(n9721), .ZN(n9225) );
  INV_X1 U6836 ( .A(n5275), .ZN(n5276) );
  NAND2_X1 U6837 ( .A1(n5276), .A2(SI_17_), .ZN(n5277) );
  MUX2_X1 U6838 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5868), .Z(n5297) );
  XNOR2_X1 U6839 ( .A(n5297), .B(SI_18_), .ZN(n5294) );
  XNOR2_X1 U6840 ( .A(n5296), .B(n5294), .ZN(n7024) );
  NAND2_X1 U6841 ( .A1(n7024), .A2(n5164), .ZN(n5285) );
  NAND2_X1 U6842 ( .A1(n5281), .A2(n5280), .ZN(n5282) );
  NAND2_X1 U6843 ( .A1(n5282), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5283) );
  XNOR2_X1 U6844 ( .A(n5283), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9993) );
  AOI22_X1 U6845 ( .A1(n9993), .A2(n6576), .B1(n5306), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n5284) );
  NAND2_X1 U6846 ( .A1(n6445), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5292) );
  INV_X1 U6847 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9683) );
  OR2_X1 U6848 ( .A1(n5460), .A2(n9683), .ZN(n5291) );
  INV_X1 U6849 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8582) );
  NAND2_X1 U6850 ( .A1(n5287), .A2(n8582), .ZN(n5288) );
  NAND2_X1 U6851 ( .A1(n5309), .A2(n5288), .ZN(n9682) );
  OR2_X1 U6852 ( .A1(n5010), .A2(n9682), .ZN(n5290) );
  INV_X1 U6853 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9798) );
  OR2_X1 U6854 ( .A1(n5210), .A2(n9798), .ZN(n5289) );
  OR2_X1 U6855 ( .A1(n9685), .A2(n9700), .ZN(n9229) );
  OR2_X1 U6856 ( .A1(n9802), .A2(n9721), .ZN(n9676) );
  AND2_X1 U6857 ( .A1(n9229), .A2(n9676), .ZN(n9335) );
  NAND2_X1 U6858 ( .A1(n9685), .A2(n9700), .ZN(n9233) );
  NAND2_X1 U6859 ( .A1(n5293), .A2(n9233), .ZN(n9660) );
  NAND2_X1 U6860 ( .A1(n5297), .A2(SI_18_), .ZN(n5298) );
  INV_X1 U6861 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7062) );
  INV_X1 U6862 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7061) );
  MUX2_X1 U6863 ( .A(n7062), .B(n7061), .S(n5868), .Z(n5300) );
  INV_X1 U6864 ( .A(SI_19_), .ZN(n5299) );
  INV_X1 U6865 ( .A(n5300), .ZN(n5301) );
  NAND2_X1 U6866 ( .A1(n5301), .A2(SI_19_), .ZN(n5302) );
  NAND2_X1 U6867 ( .A1(n5317), .A2(n5302), .ZN(n5315) );
  XNOR2_X1 U6868 ( .A(n5316), .B(n5315), .ZN(n7060) );
  NAND2_X1 U6869 ( .A1(n7060), .A2(n5164), .ZN(n5308) );
  INV_X1 U6870 ( .A(n5303), .ZN(n5462) );
  AOI22_X1 U6871 ( .A1(n5306), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n4509), .B2(
        n6576), .ZN(n5307) );
  INV_X1 U6872 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9036) );
  NAND2_X1 U6873 ( .A1(n5309), .A2(n9036), .ZN(n5310) );
  NAND2_X1 U6874 ( .A1(n5324), .A2(n5310), .ZN(n9663) );
  INV_X1 U6875 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9853) );
  OAI22_X1 U6876 ( .A1(n9663), .A2(n5010), .B1(n4990), .B2(n9853), .ZN(n5313)
         );
  INV_X1 U6877 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9793) );
  NAND2_X1 U6878 ( .A1(n5009), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5311) );
  OAI21_X1 U6879 ( .B1(n5210), .B2(n9793), .A(n5311), .ZN(n5312) );
  OR2_X1 U6880 ( .A1(n9670), .A2(n9776), .ZN(n9333) );
  NAND2_X1 U6881 ( .A1(n9670), .A2(n9776), .ZN(n9234) );
  NAND2_X1 U6882 ( .A1(n9660), .A2(n9661), .ZN(n5314) );
  INV_X1 U6883 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7245) );
  INV_X1 U6884 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7229) );
  MUX2_X1 U6885 ( .A(n7245), .B(n7229), .S(n5868), .Z(n5318) );
  INV_X1 U6886 ( .A(SI_20_), .ZN(n8609) );
  NAND2_X1 U6887 ( .A1(n5318), .A2(n8609), .ZN(n5330) );
  INV_X1 U6888 ( .A(n5318), .ZN(n5319) );
  NAND2_X1 U6889 ( .A1(n5319), .A2(SI_20_), .ZN(n5320) );
  XNOR2_X1 U6890 ( .A(n5329), .B(n5328), .ZN(n7228) );
  NAND2_X1 U6891 ( .A1(n7228), .A2(n5164), .ZN(n5322) );
  OR2_X1 U6892 ( .A1(n6428), .A2(n7229), .ZN(n5321) );
  INV_X1 U6893 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9849) );
  INV_X1 U6894 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9104) );
  NAND2_X1 U6895 ( .A1(n5324), .A2(n9104), .ZN(n5325) );
  NAND2_X1 U6896 ( .A1(n5334), .A2(n5325), .ZN(n9648) );
  OR2_X1 U6897 ( .A1(n9648), .A2(n5010), .ZN(n5327) );
  AOI22_X1 U6898 ( .A1(n5456), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n5009), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n5326) );
  OAI211_X1 U6899 ( .C1(n4990), .C2(n9849), .A(n5327), .B(n5326), .ZN(n9787)
         );
  INV_X1 U6900 ( .A(n9787), .ZN(n9769) );
  NAND2_X1 U6901 ( .A1(n5329), .A2(n5328), .ZN(n5331) );
  INV_X1 U6902 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7305) );
  INV_X1 U6903 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7401) );
  MUX2_X1 U6904 ( .A(n7305), .B(n7401), .S(n5868), .Z(n5342) );
  XNOR2_X1 U6905 ( .A(n5342), .B(SI_21_), .ZN(n5341) );
  XNOR2_X1 U6906 ( .A(n5340), .B(n5341), .ZN(n7304) );
  NAND2_X1 U6907 ( .A1(n7304), .A2(n5164), .ZN(n5333) );
  OR2_X1 U6908 ( .A1(n6428), .A2(n7401), .ZN(n5332) );
  INV_X1 U6909 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9044) );
  NAND2_X1 U6910 ( .A1(n5334), .A2(n9044), .ZN(n5335) );
  AND2_X1 U6911 ( .A1(n5352), .A2(n5335), .ZN(n9640) );
  NAND2_X1 U6912 ( .A1(n9640), .A2(n4964), .ZN(n5338) );
  AOI22_X1 U6913 ( .A1(n5009), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n6445), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n5337) );
  INV_X1 U6914 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n8465) );
  OR2_X1 U6915 ( .A1(n5210), .A2(n8465), .ZN(n5336) );
  OR2_X1 U6916 ( .A1(n9772), .A2(n9777), .ZN(n9244) );
  NAND2_X1 U6917 ( .A1(n9772), .A2(n9777), .ZN(n9608) );
  INV_X1 U6918 ( .A(n9634), .ZN(n9628) );
  NOR2_X1 U6919 ( .A1(n9628), .A2(n9299), .ZN(n5339) );
  INV_X1 U6920 ( .A(n5342), .ZN(n5343) );
  NAND2_X1 U6921 ( .A1(n5343), .A2(SI_21_), .ZN(n5344) );
  INV_X1 U6922 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7933) );
  INV_X1 U6923 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7427) );
  MUX2_X1 U6924 ( .A(n7933), .B(n7427), .S(n5868), .Z(n5346) );
  INV_X1 U6925 ( .A(SI_22_), .ZN(n5345) );
  NAND2_X1 U6926 ( .A1(n5346), .A2(n5345), .ZN(n5360) );
  INV_X1 U6927 ( .A(n5346), .ZN(n5347) );
  NAND2_X1 U6928 ( .A1(n5347), .A2(SI_22_), .ZN(n5348) );
  NAND2_X1 U6929 ( .A1(n5360), .A2(n5348), .ZN(n5361) );
  NAND2_X1 U6930 ( .A1(n7426), .A2(n5164), .ZN(n5350) );
  OR2_X1 U6931 ( .A1(n6428), .A2(n7427), .ZN(n5349) );
  INV_X1 U6932 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9128) );
  NAND2_X1 U6933 ( .A1(n5352), .A2(n9128), .ZN(n5353) );
  NAND2_X1 U6934 ( .A1(n5369), .A2(n5353), .ZN(n9619) );
  OR2_X1 U6935 ( .A1(n9619), .A2(n5010), .ZN(n5358) );
  INV_X1 U6936 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9767) );
  NAND2_X1 U6937 ( .A1(n6445), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5355) );
  NAND2_X1 U6938 ( .A1(n5009), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5354) );
  OAI211_X1 U6939 ( .C1(n5210), .C2(n9767), .A(n5355), .B(n5354), .ZN(n5356)
         );
  INV_X1 U6940 ( .A(n5356), .ZN(n5357) );
  NAND2_X1 U6941 ( .A1(n5358), .A2(n5357), .ZN(n9636) );
  INV_X1 U6942 ( .A(n9636), .ZN(n9603) );
  NAND2_X1 U6943 ( .A1(n9618), .A2(n9603), .ZN(n9296) );
  NAND2_X1 U6944 ( .A1(n9607), .A2(n9243), .ZN(n5359) );
  INV_X1 U6945 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7504) );
  INV_X1 U6946 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7501) );
  MUX2_X1 U6947 ( .A(n7504), .B(n7501), .S(n5868), .Z(n5364) );
  INV_X1 U6948 ( .A(SI_23_), .ZN(n5363) );
  NAND2_X1 U6949 ( .A1(n5364), .A2(n5363), .ZN(n5378) );
  INV_X1 U6950 ( .A(n5364), .ZN(n5365) );
  NAND2_X1 U6951 ( .A1(n5365), .A2(SI_23_), .ZN(n5366) );
  NAND2_X1 U6952 ( .A1(n7502), .A2(n5164), .ZN(n5368) );
  OR2_X1 U6953 ( .A1(n6428), .A2(n7501), .ZN(n5367) );
  INV_X1 U6954 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6521) );
  NAND2_X1 U6955 ( .A1(n5369), .A2(n6521), .ZN(n5370) );
  NAND2_X1 U6956 ( .A1(n5382), .A2(n5370), .ZN(n9594) );
  OR2_X1 U6957 ( .A1(n9594), .A2(n5010), .ZN(n5375) );
  INV_X1 U6958 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n8593) );
  NAND2_X1 U6959 ( .A1(n6445), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5372) );
  INV_X1 U6960 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9593) );
  OR2_X1 U6961 ( .A1(n5460), .A2(n9593), .ZN(n5371) );
  OAI211_X1 U6962 ( .C1(n5210), .C2(n8593), .A(n5372), .B(n5371), .ZN(n5373)
         );
  INV_X1 U6963 ( .A(n5373), .ZN(n5374) );
  NAND2_X1 U6964 ( .A1(n5375), .A2(n5374), .ZN(n9614) );
  INV_X1 U6965 ( .A(n9614), .ZN(n9581) );
  NAND2_X1 U6966 ( .A1(n9761), .A2(n9581), .ZN(n9249) );
  NAND2_X1 U6967 ( .A1(n9599), .A2(n9598), .ZN(n9597) );
  NAND2_X1 U6968 ( .A1(n9597), .A2(n9336), .ZN(n9577) );
  NAND2_X1 U6969 ( .A1(n5377), .A2(n5376), .ZN(n5379) );
  INV_X1 U6970 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7593) );
  INV_X1 U6971 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7590) );
  MUX2_X1 U6972 ( .A(n7593), .B(n7590), .S(n5868), .Z(n5390) );
  XNOR2_X1 U6973 ( .A(n5390), .B(SI_24_), .ZN(n5389) );
  XNOR2_X1 U6974 ( .A(n5394), .B(n5389), .ZN(n5909) );
  NAND2_X1 U6975 ( .A1(n5909), .A2(n5164), .ZN(n5381) );
  OR2_X1 U6976 ( .A1(n6428), .A2(n7590), .ZN(n5380) );
  INV_X1 U6977 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9095) );
  NAND2_X1 U6978 ( .A1(n5382), .A2(n9095), .ZN(n5383) );
  AND2_X1 U6979 ( .A1(n5403), .A2(n5383), .ZN(n9574) );
  NAND2_X1 U6980 ( .A1(n9574), .A2(n4964), .ZN(n5388) );
  INV_X1 U6981 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n8454) );
  NAND2_X1 U6982 ( .A1(n6445), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U6983 ( .A1(n5009), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5384) );
  OAI211_X1 U6984 ( .C1(n5210), .C2(n8454), .A(n5385), .B(n5384), .ZN(n5386)
         );
  INV_X1 U6985 ( .A(n5386), .ZN(n5387) );
  OR2_X2 U6986 ( .A1(n9756), .A2(n6522), .ZN(n9361) );
  NAND2_X1 U6987 ( .A1(n9756), .A2(n6522), .ZN(n9253) );
  NAND2_X1 U6988 ( .A1(n9577), .A2(n9583), .ZN(n9576) );
  NAND2_X1 U6989 ( .A1(n9576), .A2(n9361), .ZN(n9557) );
  INV_X1 U6990 ( .A(n5389), .ZN(n5393) );
  INV_X1 U6991 ( .A(n5390), .ZN(n5391) );
  NAND2_X1 U6992 ( .A1(n5391), .A2(SI_24_), .ZN(n5392) );
  INV_X1 U6993 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7731) );
  INV_X1 U6994 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8552) );
  MUX2_X1 U6995 ( .A(n7731), .B(n8552), .S(n5868), .Z(n5396) );
  INV_X1 U6996 ( .A(SI_25_), .ZN(n5395) );
  NAND2_X1 U6997 ( .A1(n5396), .A2(n5395), .ZN(n5410) );
  INV_X1 U6998 ( .A(n5396), .ZN(n5397) );
  NAND2_X1 U6999 ( .A1(n5397), .A2(SI_25_), .ZN(n5398) );
  NAND2_X1 U7000 ( .A1(n5410), .A2(n5398), .ZN(n5411) );
  NAND2_X1 U7001 ( .A1(n7730), .A2(n5164), .ZN(n5400) );
  OR2_X1 U7002 ( .A1(n6428), .A2(n8552), .ZN(n5399) );
  INV_X1 U7003 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U7004 ( .A1(n5403), .A2(n5402), .ZN(n5404) );
  NAND2_X1 U7005 ( .A1(n5420), .A2(n5404), .ZN(n9564) );
  OR2_X1 U7006 ( .A1(n9564), .A2(n5010), .ZN(n5409) );
  INV_X1 U7007 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9750) );
  NAND2_X1 U7008 ( .A1(n6445), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U7009 ( .A1(n5009), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5405) );
  OAI211_X1 U7010 ( .C1(n5210), .C2(n9750), .A(n5406), .B(n5405), .ZN(n5407)
         );
  INV_X1 U7011 ( .A(n5407), .ZN(n5408) );
  NAND2_X1 U7012 ( .A1(n9563), .A2(n9545), .ZN(n9262) );
  NAND2_X1 U7013 ( .A1(n9557), .A2(n9262), .ZN(n9542) );
  INV_X1 U7014 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7823) );
  INV_X1 U7015 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7788) );
  MUX2_X1 U7016 ( .A(n7823), .B(n7788), .S(n5868), .Z(n5414) );
  INV_X1 U7017 ( .A(SI_26_), .ZN(n5413) );
  NAND2_X1 U7018 ( .A1(n5414), .A2(n5413), .ZN(n5430) );
  INV_X1 U7019 ( .A(n5414), .ZN(n5415) );
  NAND2_X1 U7020 ( .A1(n5415), .A2(SI_26_), .ZN(n5416) );
  XNOR2_X1 U7021 ( .A(n5429), .B(n5428), .ZN(n7787) );
  NAND2_X1 U7022 ( .A1(n7787), .A2(n5164), .ZN(n5418) );
  OR2_X1 U7023 ( .A1(n6428), .A2(n7788), .ZN(n5417) );
  INV_X1 U7024 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9151) );
  NAND2_X1 U7025 ( .A1(n5420), .A2(n9151), .ZN(n5421) );
  NAND2_X1 U7026 ( .A1(n5454), .A2(n5421), .ZN(n9549) );
  OR2_X1 U7027 ( .A1(n9549), .A2(n5010), .ZN(n5426) );
  INV_X1 U7028 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9745) );
  NAND2_X1 U7029 ( .A1(n6445), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U7030 ( .A1(n5009), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5422) );
  OAI211_X1 U7031 ( .C1(n5210), .C2(n9745), .A(n5423), .B(n5422), .ZN(n5424)
         );
  INV_X1 U7032 ( .A(n5424), .ZN(n5425) );
  OR2_X1 U7033 ( .A1(n9265), .A2(n9533), .ZN(n9261) );
  AND2_X1 U7034 ( .A1(n9261), .A2(n9541), .ZN(n9393) );
  NAND2_X1 U7035 ( .A1(n9542), .A2(n9393), .ZN(n5427) );
  NAND2_X1 U7036 ( .A1(n9265), .A2(n9533), .ZN(n9385) );
  INV_X1 U7037 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7883) );
  INV_X1 U7038 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7860) );
  MUX2_X1 U7039 ( .A(n7883), .B(n7860), .S(n5868), .Z(n5432) );
  INV_X1 U7040 ( .A(SI_27_), .ZN(n8541) );
  NAND2_X1 U7041 ( .A1(n5432), .A2(n8541), .ZN(n5445) );
  INV_X1 U7042 ( .A(n5432), .ZN(n5433) );
  NAND2_X1 U7043 ( .A1(n5433), .A2(SI_27_), .ZN(n5434) );
  NAND2_X1 U7044 ( .A1(n7859), .A2(n5164), .ZN(n5436) );
  OR2_X1 U7045 ( .A1(n6428), .A2(n7860), .ZN(n5435) );
  XNOR2_X1 U7046 ( .A(n5454), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9527) );
  NAND2_X1 U7047 ( .A1(n9527), .A2(n4964), .ZN(n5442) );
  INV_X1 U7048 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U7049 ( .A1(n6445), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5438) );
  NAND2_X1 U7050 ( .A1(n5456), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5437) );
  OAI211_X1 U7051 ( .C1(n5460), .C2(n5439), .A(n5438), .B(n5437), .ZN(n5440)
         );
  INV_X1 U7052 ( .A(n5440), .ZN(n5441) );
  NAND2_X1 U7053 ( .A1(n9737), .A2(n9546), .ZN(n9271) );
  INV_X1 U7054 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7914) );
  INV_X1 U7055 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7910) );
  MUX2_X1 U7056 ( .A(n7914), .B(n7910), .S(n5868), .Z(n5447) );
  INV_X1 U7057 ( .A(SI_28_), .ZN(n8620) );
  NAND2_X1 U7058 ( .A1(n5447), .A2(n8620), .ZN(n6406) );
  INV_X1 U7059 ( .A(n5447), .ZN(n5448) );
  NAND2_X1 U7060 ( .A1(n5448), .A2(SI_28_), .ZN(n5449) );
  NAND2_X1 U7061 ( .A1(n7911), .A2(n5164), .ZN(n5451) );
  OR2_X1 U7062 ( .A1(n6428), .A2(n7910), .ZN(n5450) );
  INV_X1 U7063 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5842) );
  INV_X1 U7064 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5452) );
  OAI21_X1 U7065 ( .B1(n5454), .B2(n5842), .A(n5452), .ZN(n5455) );
  NAND2_X1 U7066 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5453) );
  INV_X1 U7067 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U7068 ( .A1(n6445), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U7069 ( .A1(n5456), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5457) );
  OAI211_X1 U7070 ( .C1(n5460), .C2(n5459), .A(n5458), .B(n5457), .ZN(n5461)
         );
  NAND2_X1 U7071 ( .A1(n6464), .A2(n9534), .ZN(n9272) );
  NAND2_X1 U7072 ( .A1(n9391), .A2(n9272), .ZN(n9295) );
  XNOR2_X1 U7073 ( .A(n6442), .B(n9295), .ZN(n5484) );
  NOR2_X1 U7074 ( .A1(n5463), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U7075 ( .A1(n5465), .A2(n5464), .ZN(n5466) );
  INV_X1 U7076 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U7077 ( .A1(n5475), .A2(n5467), .ZN(n5468) );
  INV_X1 U7078 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U7079 ( .A1(n5471), .A2(n5469), .ZN(n5474) );
  NAND2_X1 U7080 ( .A1(n5474), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U7081 ( .A1(n9452), .A2(n4509), .ZN(n5477) );
  INV_X1 U7082 ( .A(n5471), .ZN(n5472) );
  OR2_X1 U7083 ( .A1(n9398), .A2(n9443), .ZN(n5476) );
  NAND2_X1 U7084 ( .A1(n9452), .A2(n9411), .ZN(n9332) );
  INV_X1 U7085 ( .A(n9332), .ZN(n5832) );
  INV_X1 U7086 ( .A(n5478), .ZN(n9449) );
  INV_X1 U7087 ( .A(n5479), .ZN(n9508) );
  INV_X1 U7088 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6453) );
  NAND2_X1 U7089 ( .A1(n6445), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5481) );
  NAND2_X1 U7090 ( .A1(n5009), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5480) );
  OAI211_X1 U7091 ( .C1(n5210), .C2(n6453), .A(n5481), .B(n5480), .ZN(n5482)
         );
  AOI21_X1 U7092 ( .B1(n9508), .B2(n4964), .A(n5482), .ZN(n6982) );
  OAI22_X1 U7093 ( .A1(n9546), .A2(n10015), .B1(n6982), .B2(n10062), .ZN(n5483) );
  NAND2_X1 U7094 ( .A1(n7318), .A2(n10057), .ZN(n7317) );
  INV_X1 U7095 ( .A(n7794), .ZN(n9912) );
  NAND2_X1 U7096 ( .A1(n7663), .A2(n9912), .ZN(n7662) );
  NAND2_X1 U7097 ( .A1(n7843), .A2(n9171), .ZN(n9722) );
  INV_X1 U7098 ( .A(n9685), .ZN(n9859) );
  INV_X1 U7099 ( .A(n9670), .ZN(n9855) );
  AND2_X1 U7100 ( .A1(n9851), .A2(n9855), .ZN(n5485) );
  INV_X1 U7101 ( .A(n9761), .ZN(n9592) );
  NOR2_X2 U7102 ( .A1(n9525), .A2(n9737), .ZN(n5487) );
  NAND2_X1 U7103 ( .A1(n9405), .A2(n9398), .ZN(n10032) );
  NAND2_X1 U7104 ( .A1(n6464), .A2(n9526), .ZN(n5488) );
  NAND3_X1 U7105 ( .A1(n6451), .A2(n10003), .A3(n5488), .ZN(n9516) );
  AND2_X1 U7106 ( .A1(n5593), .A2(n10034), .ZN(n7197) );
  NAND2_X1 U7107 ( .A1(n9305), .A2(n7197), .ZN(n7196) );
  NAND2_X1 U7108 ( .A1(n5597), .A2(n4388), .ZN(n5489) );
  NAND2_X1 U7109 ( .A1(n7196), .A2(n5489), .ZN(n6999) );
  INV_X1 U7110 ( .A(n6999), .ZN(n5491) );
  NAND2_X1 U7111 ( .A1(n5491), .A2(n5490), .ZN(n7001) );
  NAND2_X1 U7112 ( .A1(n7312), .A2(n5607), .ZN(n5492) );
  NAND2_X1 U7113 ( .A1(n7001), .A2(n5492), .ZN(n7307) );
  NAND2_X1 U7114 ( .A1(n7307), .A2(n9304), .ZN(n7306) );
  NAND2_X1 U7115 ( .A1(n7372), .A2(n10057), .ZN(n5493) );
  NAND2_X1 U7116 ( .A1(n7306), .A2(n5493), .ZN(n7048) );
  NAND2_X1 U7117 ( .A1(n9176), .A2(n9379), .ZN(n7051) );
  NAND2_X1 U7118 ( .A1(n7048), .A2(n7051), .ZN(n7383) );
  NAND2_X1 U7119 ( .A1(n7389), .A2(n7056), .ZN(n7382) );
  AND2_X1 U7120 ( .A1(n7235), .A2(n7382), .ZN(n5494) );
  NAND2_X1 U7121 ( .A1(n9467), .A2(n7394), .ZN(n5495) );
  NAND2_X1 U7122 ( .A1(n9188), .A2(n9300), .ZN(n9183) );
  NAND2_X1 U7123 ( .A1(n7329), .A2(n9309), .ZN(n7328) );
  NAND2_X1 U7124 ( .A1(n7483), .A2(n7462), .ZN(n5496) );
  NAND2_X1 U7125 ( .A1(n9464), .A2(n7496), .ZN(n5497) );
  OR2_X1 U7126 ( .A1(n10027), .A2(n9463), .ZN(n5499) );
  AND2_X1 U7127 ( .A1(n10027), .A2(n9463), .ZN(n5498) );
  AOI21_X1 U7128 ( .B1(n10010), .B2(n5499), .A(n5498), .ZN(n7527) );
  NAND2_X1 U7129 ( .A1(n9346), .A2(n9195), .ZN(n9313) );
  NAND2_X1 U7130 ( .A1(n7527), .A2(n9313), .ZN(n7526) );
  INV_X1 U7131 ( .A(n10017), .ZN(n9462) );
  OR2_X1 U7132 ( .A1(n7603), .A2(n9462), .ZN(n5500) );
  NAND2_X1 U7133 ( .A1(n7735), .A2(n9202), .ZN(n9314) );
  AND2_X1 U7134 ( .A1(n9816), .A2(n9460), .ZN(n5508) );
  INV_X1 U7135 ( .A(n9113), .ZN(n9820) );
  NAND2_X1 U7136 ( .A1(n9058), .A2(n9820), .ZN(n5507) );
  INV_X1 U7137 ( .A(n5507), .ZN(n5501) );
  NAND2_X1 U7138 ( .A1(n9203), .A2(n9210), .ZN(n9315) );
  OR2_X1 U7139 ( .A1(n5501), .A2(n9315), .ZN(n7695) );
  OR2_X1 U7140 ( .A1(n5508), .A2(n7695), .ZN(n5506) );
  AND2_X1 U7141 ( .A1(n9314), .A2(n5506), .ZN(n5502) );
  OR2_X1 U7142 ( .A1(n9816), .A2(n9460), .ZN(n5505) );
  AND2_X1 U7143 ( .A1(n5502), .A2(n5505), .ZN(n7757) );
  NOR2_X1 U7144 ( .A1(n9030), .A2(n9817), .ZN(n5514) );
  INV_X1 U7145 ( .A(n5514), .ZN(n5503) );
  AND2_X1 U7146 ( .A1(n7757), .A2(n5503), .ZN(n5504) );
  NAND2_X1 U7147 ( .A1(n7666), .A2(n5504), .ZN(n5516) );
  INV_X1 U7148 ( .A(n5505), .ZN(n5513) );
  INV_X1 U7149 ( .A(n5506), .ZN(n5511) );
  INV_X1 U7150 ( .A(n7746), .ZN(n9461) );
  NAND2_X1 U7151 ( .A1(n7794), .A2(n9461), .ZN(n7739) );
  AND2_X1 U7152 ( .A1(n7739), .A2(n5507), .ZN(n7694) );
  INV_X1 U7153 ( .A(n5508), .ZN(n5509) );
  AND2_X1 U7154 ( .A1(n7694), .A2(n5509), .ZN(n5510) );
  OR2_X1 U7155 ( .A1(n5511), .A2(n5510), .ZN(n5512) );
  NOR2_X1 U7156 ( .A1(n4924), .A2(n4923), .ZN(n5515) );
  NAND2_X1 U7157 ( .A1(n5516), .A2(n5515), .ZN(n7839) );
  INV_X1 U7158 ( .A(n9699), .ZN(n9459) );
  NAND2_X1 U7159 ( .A1(n9727), .A2(n9459), .ZN(n5518) );
  NAND2_X1 U7160 ( .A1(n9712), .A2(n5518), .ZN(n5519) );
  AND2_X1 U7161 ( .A1(n9709), .A2(n5519), .ZN(n9689) );
  OR2_X1 U7162 ( .A1(n9802), .A2(n9806), .ZN(n5517) );
  AND2_X1 U7163 ( .A1(n9689), .A2(n5517), .ZN(n5521) );
  INV_X1 U7164 ( .A(n5517), .ZN(n5520) );
  INV_X1 U7165 ( .A(n9074), .ZN(n9807) );
  NAND2_X1 U7166 ( .A1(n7846), .A2(n9807), .ZN(n9710) );
  AOI21_X1 U7167 ( .B1(n7839), .B2(n5521), .A(n4913), .ZN(n5523) );
  NAND2_X1 U7168 ( .A1(n9802), .A2(n9806), .ZN(n5522) );
  NAND2_X1 U7169 ( .A1(n5523), .A2(n5522), .ZN(n9681) );
  NAND2_X1 U7170 ( .A1(n9229), .A2(n9233), .ZN(n9680) );
  NAND2_X1 U7171 ( .A1(n9681), .A2(n9680), .ZN(n5525) );
  INV_X1 U7172 ( .A(n9700), .ZN(n9786) );
  NAND2_X1 U7173 ( .A1(n9685), .A2(n9786), .ZN(n5524) );
  OR2_X1 U7174 ( .A1(n9670), .A2(n9651), .ZN(n5526) );
  NAND2_X1 U7175 ( .A1(n4401), .A2(n9628), .ZN(n9627) );
  INV_X1 U7176 ( .A(n9777), .ZN(n9613) );
  NAND2_X1 U7177 ( .A1(n9772), .A2(n9613), .ZN(n5527) );
  NAND2_X1 U7178 ( .A1(n9627), .A2(n5527), .ZN(n9606) );
  OR2_X1 U7179 ( .A1(n9636), .A2(n9618), .ZN(n5528) );
  NAND2_X1 U7180 ( .A1(n9618), .A2(n9636), .ZN(n5529) );
  OR2_X1 U7181 ( .A1(n9761), .A2(n9614), .ZN(n5530) );
  NAND2_X1 U7182 ( .A1(n5531), .A2(n5530), .ZN(n9584) );
  INV_X1 U7183 ( .A(n9584), .ZN(n5533) );
  NAND2_X1 U7184 ( .A1(n9756), .A2(n9600), .ZN(n5534) );
  NAND2_X1 U7185 ( .A1(n9541), .A2(n9262), .ZN(n9558) );
  NOR2_X1 U7186 ( .A1(n9265), .A2(n9560), .ZN(n5535) );
  NOR2_X1 U7187 ( .A1(n9524), .A2(n9431), .ZN(n5536) );
  INV_X1 U7188 ( .A(n9546), .ZN(n9458) );
  NOR2_X1 U7189 ( .A1(n5536), .A2(n4438), .ZN(n5537) );
  NAND2_X1 U7190 ( .A1(n5537), .A2(n9295), .ZN(n6438) );
  OAI21_X1 U7191 ( .B1(n5537), .B2(n9295), .A(n6438), .ZN(n9523) );
  NAND2_X1 U7192 ( .A1(n9452), .A2(n4390), .ZN(n5840) );
  MUX2_X1 U7193 ( .A(n9452), .B(n5840), .S(n5839), .Z(n7672) );
  INV_X1 U7194 ( .A(n7672), .ZN(n10066) );
  OR2_X1 U7195 ( .A1(n9523), .A2(n7672), .ZN(n5538) );
  NAND3_X1 U7196 ( .A1(n9515), .A2(n9516), .A3(n5538), .ZN(n5576) );
  NAND2_X1 U7197 ( .A1(n5540), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5542) );
  NAND2_X1 U7198 ( .A1(n5542), .A2(n5541), .ZN(n5547) );
  OR2_X1 U7199 ( .A1(n5542), .A2(n5541), .ZN(n5543) );
  NAND2_X1 U7200 ( .A1(n7733), .A2(P1_B_REG_SCAN_IN), .ZN(n5546) );
  NAND2_X1 U7201 ( .A1(n4429), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5545) );
  XNOR2_X1 U7202 ( .A(n5545), .B(n5544), .ZN(n7591) );
  INV_X1 U7203 ( .A(n7591), .ZN(n5568) );
  MUX2_X1 U7204 ( .A(n5546), .B(P1_B_REG_SCAN_IN), .S(n5568), .Z(n5549) );
  NAND2_X1 U7205 ( .A1(n5549), .A2(n5552), .ZN(n10040) );
  INV_X1 U7206 ( .A(n7733), .ZN(n5550) );
  OAI22_X1 U7207 ( .A1(n10040), .A2(P1_D_REG_1__SCAN_IN), .B1(n5552), .B2(
        n5550), .ZN(n7127) );
  NOR2_X1 U7208 ( .A1(n7733), .A2(n7591), .ZN(n5551) );
  NAND2_X1 U7209 ( .A1(n5553), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5554) );
  XNOR2_X1 U7210 ( .A(n5554), .B(n4902), .ZN(n6489) );
  AND2_X1 U7211 ( .A1(n6489), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5555) );
  INV_X1 U7212 ( .A(n10040), .ZN(n5566) );
  NOR2_X1 U7213 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .ZN(
        n8431) );
  NOR4_X1 U7214 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n5558) );
  NOR4_X1 U7215 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5557) );
  NOR4_X1 U7216 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5556) );
  AND4_X1 U7217 ( .A1(n8431), .A2(n5558), .A3(n5557), .A4(n5556), .ZN(n5564)
         );
  NOR4_X1 U7218 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n5562) );
  NOR4_X1 U7219 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n5561) );
  NOR4_X1 U7220 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n5560) );
  NOR4_X1 U7221 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5559) );
  AND4_X1 U7222 ( .A1(n5562), .A2(n5561), .A3(n5560), .A4(n5559), .ZN(n5563)
         );
  NAND2_X1 U7223 ( .A1(n5564), .A2(n5563), .ZN(n5565) );
  NAND2_X1 U7224 ( .A1(n5566), .A2(n5565), .ZN(n7128) );
  AND3_X1 U7225 ( .A1(n7127), .A2(n10051), .A3(n7128), .ZN(n5567) );
  OAI211_X1 U7226 ( .C1(n5848), .C2(n9411), .A(n5567), .B(n7131), .ZN(n5575)
         );
  OAI22_X1 U7227 ( .A1(n10040), .A2(P1_D_REG_0__SCAN_IN), .B1(n5552), .B2(
        n5568), .ZN(n7129) );
  INV_X1 U7228 ( .A(n7129), .ZN(n9867) );
  INV_X1 U7229 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n5569) );
  NOR2_X1 U7230 ( .A1(n10076), .A2(n5569), .ZN(n5572) );
  INV_X1 U7231 ( .A(n10032), .ZN(n6881) );
  INV_X1 U7232 ( .A(n5584), .ZN(n5570) );
  NAND2_X1 U7233 ( .A1(n5576), .A2(n10083), .ZN(n5580) );
  OAI21_X1 U7234 ( .B1(n5486), .B2(n9815), .A(n5577), .ZN(n5578) );
  INV_X1 U7235 ( .A(n5578), .ZN(n5579) );
  NAND2_X1 U7236 ( .A1(n5580), .A2(n5579), .ZN(P1_U3551) );
  INV_X2 U7237 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U7238 ( .A(n5839), .ZN(n5581) );
  AND2_X4 U7239 ( .A1(n5840), .A2(n5839), .ZN(n7330) );
  XNOR2_X1 U7240 ( .A(n5583), .B(n6460), .ZN(n5625) );
  INV_X1 U7241 ( .A(n5649), .ZN(n5653) );
  NAND2_X1 U7242 ( .A1(n9405), .A2(n5584), .ZN(n5585) );
  OR2_X1 U7243 ( .A1(n7389), .A2(n5592), .ZN(n5587) );
  NAND2_X1 U7244 ( .A1(n7371), .A2(n6463), .ZN(n5586) );
  NAND2_X1 U7245 ( .A1(n5587), .A2(n5586), .ZN(n5624) );
  XNOR2_X1 U7246 ( .A(n5625), .B(n5624), .ZN(n7031) );
  INV_X1 U7247 ( .A(n7031), .ZN(n5623) );
  NAND2_X1 U7248 ( .A1(n5593), .A2(n5596), .ZN(n5590) );
  NOR2_X1 U7249 ( .A1(n5582), .A2(n6612), .ZN(n5588) );
  AOI21_X1 U7250 ( .B1(n10034), .B2(n5653), .A(n5588), .ZN(n5589) );
  NAND2_X1 U7251 ( .A1(n5590), .A2(n5589), .ZN(n6837) );
  INV_X1 U7252 ( .A(n6837), .ZN(n5591) );
  NAND2_X1 U7253 ( .A1(n5591), .A2(n6460), .ZN(n5595) );
  INV_X1 U7254 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n8650) );
  NOR2_X1 U7255 ( .A1(n5582), .A2(n8650), .ZN(n5594) );
  NAND2_X1 U7256 ( .A1(n6839), .A2(n6837), .ZN(n6838) );
  NAND2_X1 U7257 ( .A1(n5597), .A2(n5596), .ZN(n5600) );
  NAND2_X1 U7258 ( .A1(n5600), .A2(n5599), .ZN(n5602) );
  INV_X1 U7259 ( .A(n5602), .ZN(n5601) );
  NAND2_X1 U7260 ( .A1(n5602), .A2(n7330), .ZN(n5603) );
  AOI22_X1 U7261 ( .A1(n5597), .A2(n6462), .B1(n4388), .B2(n5596), .ZN(n6886)
         );
  NAND2_X1 U7262 ( .A1(n5605), .A2(n5606), .ZN(n6889) );
  NAND2_X1 U7263 ( .A1(n6885), .A2(n6889), .ZN(n6945) );
  XNOR2_X1 U7264 ( .A(n5608), .B(n7330), .ZN(n5611) );
  OR2_X1 U7265 ( .A1(n7312), .A2(n5592), .ZN(n5610) );
  NAND2_X1 U7266 ( .A1(n6998), .A2(n5596), .ZN(n5609) );
  NAND2_X1 U7267 ( .A1(n5610), .A2(n5609), .ZN(n5612) );
  XNOR2_X1 U7268 ( .A(n5611), .B(n5612), .ZN(n6944) );
  NAND2_X1 U7269 ( .A1(n6945), .A2(n6944), .ZN(n5615) );
  INV_X1 U7270 ( .A(n5612), .ZN(n5613) );
  NAND2_X1 U7271 ( .A1(n5611), .A2(n5613), .ZN(n5614) );
  NAND2_X1 U7272 ( .A1(n5615), .A2(n5614), .ZN(n6973) );
  NAND2_X1 U7273 ( .A1(n9469), .A2(n5596), .ZN(n5617) );
  OR2_X1 U7274 ( .A1(n10057), .A2(n5649), .ZN(n5616) );
  AOI22_X1 U7275 ( .A1(n9469), .A2(n6462), .B1(n7321), .B2(n5596), .ZN(n5620)
         );
  XNOR2_X1 U7276 ( .A(n5619), .B(n5620), .ZN(n6974) );
  INV_X1 U7277 ( .A(n5619), .ZN(n5621) );
  NAND2_X1 U7278 ( .A1(n5621), .A2(n5620), .ZN(n5622) );
  NAND2_X1 U7279 ( .A1(n5625), .A2(n5624), .ZN(n5626) );
  OAI22_X1 U7280 ( .A1(n7373), .A2(n6457), .B1(n10061), .B2(n5649), .ZN(n5627)
         );
  XNOR2_X1 U7281 ( .A(n5627), .B(n7330), .ZN(n5631) );
  OR2_X1 U7282 ( .A1(n7373), .A2(n5592), .ZN(n5629) );
  NAND2_X1 U7283 ( .A1(n7394), .A2(n6463), .ZN(n5628) );
  AND2_X1 U7284 ( .A1(n5629), .A2(n5628), .ZN(n7189) );
  INV_X1 U7285 ( .A(n5630), .ZN(n5632) );
  NAND2_X1 U7286 ( .A1(n5632), .A2(n5631), .ZN(n5633) );
  OAI22_X1 U7287 ( .A1(n10063), .A2(n6457), .B1(n7469), .B2(n5649), .ZN(n5634)
         );
  XNOR2_X1 U7288 ( .A(n5634), .B(n7330), .ZN(n7284) );
  OR2_X1 U7289 ( .A1(n10063), .A2(n5592), .ZN(n5637) );
  NAND2_X1 U7290 ( .A1(n5635), .A2(n6463), .ZN(n5636) );
  NAND2_X1 U7291 ( .A1(n5637), .A2(n5636), .ZN(n7285) );
  INV_X1 U7292 ( .A(n7284), .ZN(n5638) );
  OAI22_X1 U7293 ( .A1(n7483), .A2(n6457), .B1(n7462), .B2(n5649), .ZN(n5639)
         );
  XNOR2_X1 U7294 ( .A(n5639), .B(n7330), .ZN(n5642) );
  OR2_X1 U7295 ( .A1(n7483), .A2(n5592), .ZN(n5641) );
  NAND2_X1 U7296 ( .A1(n7448), .A2(n6463), .ZN(n5640) );
  AND2_X1 U7297 ( .A1(n5641), .A2(n5640), .ZN(n5643) );
  NAND2_X1 U7298 ( .A1(n5642), .A2(n5643), .ZN(n7454) );
  NAND2_X1 U7299 ( .A1(n7453), .A2(n7454), .ZN(n5646) );
  INV_X1 U7300 ( .A(n5642), .ZN(n5645) );
  INV_X1 U7301 ( .A(n5643), .ZN(n5644) );
  NAND2_X1 U7302 ( .A1(n5645), .A2(n5644), .ZN(n7455) );
  OR2_X1 U7303 ( .A1(n10016), .A2(n5592), .ZN(n5648) );
  NAND2_X1 U7304 ( .A1(n7496), .A2(n6463), .ZN(n5647) );
  NAND2_X1 U7305 ( .A1(n5648), .A2(n5647), .ZN(n5651) );
  OAI22_X1 U7306 ( .A1(n10016), .A2(n6457), .B1(n7644), .B2(n5649), .ZN(n5650)
         );
  XNOR2_X1 U7307 ( .A(n5650), .B(n7330), .ZN(n7634) );
  INV_X1 U7308 ( .A(n5651), .ZN(n5652) );
  NAND2_X1 U7309 ( .A1(n10027), .A2(n6456), .ZN(n5655) );
  NAND2_X1 U7310 ( .A1(n9463), .A2(n6463), .ZN(n5654) );
  NAND2_X1 U7311 ( .A1(n5655), .A2(n5654), .ZN(n5656) );
  XNOR2_X1 U7312 ( .A(n5656), .B(n6460), .ZN(n5657) );
  AOI22_X1 U7313 ( .A1(n10027), .A2(n6463), .B1(n6462), .B2(n9463), .ZN(n5658)
         );
  XNOR2_X1 U7314 ( .A(n5657), .B(n5658), .ZN(n7619) );
  INV_X1 U7315 ( .A(n5657), .ZN(n5659) );
  NAND2_X1 U7316 ( .A1(n5659), .A2(n5658), .ZN(n5660) );
  NAND2_X1 U7317 ( .A1(n7603), .A2(n6456), .ZN(n5662) );
  OR2_X1 U7318 ( .A1(n10017), .A2(n6457), .ZN(n5661) );
  NAND2_X1 U7319 ( .A1(n5662), .A2(n5661), .ZN(n5663) );
  XNOR2_X1 U7320 ( .A(n5663), .B(n7330), .ZN(n7677) );
  NAND2_X1 U7321 ( .A1(n7603), .A2(n6463), .ZN(n5665) );
  OR2_X1 U7322 ( .A1(n10017), .A2(n5592), .ZN(n5664) );
  AND2_X1 U7323 ( .A1(n5665), .A2(n5664), .ZN(n5666) );
  INV_X1 U7324 ( .A(n7677), .ZN(n5667) );
  INV_X1 U7325 ( .A(n5666), .ZN(n7676) );
  NAND2_X1 U7326 ( .A1(n5667), .A2(n7676), .ZN(n5668) );
  NAND2_X1 U7327 ( .A1(n7794), .A2(n6456), .ZN(n5670) );
  OR2_X1 U7328 ( .A1(n7746), .A2(n6457), .ZN(n5669) );
  NAND2_X1 U7329 ( .A1(n5670), .A2(n5669), .ZN(n5671) );
  XNOR2_X1 U7330 ( .A(n5671), .B(n6460), .ZN(n5673) );
  NOR2_X1 U7331 ( .A1(n7746), .A2(n5592), .ZN(n5672) );
  AOI21_X1 U7332 ( .B1(n7794), .B2(n6463), .A(n5672), .ZN(n5674) );
  XNOR2_X1 U7333 ( .A(n5673), .B(n5674), .ZN(n7791) );
  INV_X1 U7334 ( .A(n5673), .ZN(n5675) );
  NAND2_X1 U7335 ( .A1(n9058), .A2(n6456), .ZN(n5677) );
  OR2_X1 U7336 ( .A1(n9113), .A2(n6457), .ZN(n5676) );
  NAND2_X1 U7337 ( .A1(n5677), .A2(n5676), .ZN(n5678) );
  XNOR2_X1 U7338 ( .A(n5678), .B(n7330), .ZN(n5681) );
  NOR2_X1 U7339 ( .A1(n9113), .A2(n5592), .ZN(n5679) );
  AOI21_X1 U7340 ( .B1(n9058), .B2(n6463), .A(n5679), .ZN(n5680) );
  NAND2_X1 U7341 ( .A1(n5681), .A2(n5680), .ZN(n5685) );
  OR2_X1 U7342 ( .A1(n5681), .A2(n5680), .ZN(n5682) );
  NAND2_X1 U7343 ( .A1(n5685), .A2(n5682), .ZN(n9053) );
  NAND2_X1 U7344 ( .A1(n9816), .A2(n6456), .ZN(n5687) );
  NAND2_X1 U7345 ( .A1(n9460), .A2(n6463), .ZN(n5686) );
  NAND2_X1 U7346 ( .A1(n5687), .A2(n5686), .ZN(n5688) );
  XNOR2_X1 U7347 ( .A(n5688), .B(n7330), .ZN(n5690) );
  AND2_X1 U7348 ( .A1(n9460), .A2(n6462), .ZN(n5689) );
  AOI21_X1 U7349 ( .B1(n9816), .B2(n6463), .A(n5689), .ZN(n5691) );
  NAND2_X1 U7350 ( .A1(n5690), .A2(n5691), .ZN(n9110) );
  INV_X1 U7351 ( .A(n5690), .ZN(n5693) );
  INV_X1 U7352 ( .A(n5691), .ZN(n5692) );
  NAND2_X1 U7353 ( .A1(n5693), .A2(n5692), .ZN(n9109) );
  INV_X1 U7354 ( .A(n5702), .ZN(n5698) );
  NAND2_X1 U7355 ( .A1(n9030), .A2(n6456), .ZN(n5695) );
  NAND2_X1 U7356 ( .A1(n9817), .A2(n6463), .ZN(n5694) );
  NAND2_X1 U7357 ( .A1(n5695), .A2(n5694), .ZN(n5696) );
  XNOR2_X1 U7358 ( .A(n5696), .B(n6460), .ZN(n5701) );
  INV_X1 U7359 ( .A(n5701), .ZN(n5697) );
  NAND2_X1 U7360 ( .A1(n5698), .A2(n5697), .ZN(n9024) );
  NAND2_X1 U7361 ( .A1(n9030), .A2(n6463), .ZN(n5700) );
  NAND2_X1 U7362 ( .A1(n9817), .A2(n6462), .ZN(n5699) );
  NAND2_X1 U7363 ( .A1(n5700), .A2(n5699), .ZN(n9026) );
  NAND2_X1 U7364 ( .A1(n9024), .A2(n9026), .ZN(n5710) );
  NAND2_X1 U7365 ( .A1(n5702), .A2(n5701), .ZN(n5709) );
  NAND2_X1 U7366 ( .A1(n7846), .A2(n6456), .ZN(n5704) );
  OR2_X1 U7367 ( .A1(n9074), .A2(n6457), .ZN(n5703) );
  NAND2_X1 U7368 ( .A1(n5704), .A2(n5703), .ZN(n5705) );
  XNOR2_X1 U7369 ( .A(n5705), .B(n7330), .ZN(n5711) );
  AND2_X1 U7370 ( .A1(n5709), .A2(n5711), .ZN(n5706) );
  NAND2_X1 U7371 ( .A1(n5710), .A2(n5706), .ZN(n9156) );
  NAND2_X1 U7372 ( .A1(n7846), .A2(n6463), .ZN(n5708) );
  OR2_X1 U7373 ( .A1(n9074), .A2(n5592), .ZN(n5707) );
  NAND2_X1 U7374 ( .A1(n5708), .A2(n5707), .ZN(n9158) );
  NAND2_X1 U7375 ( .A1(n9156), .A2(n9158), .ZN(n5741) );
  NAND2_X1 U7376 ( .A1(n5710), .A2(n5709), .ZN(n5713) );
  INV_X1 U7377 ( .A(n5711), .ZN(n5712) );
  NAND2_X1 U7378 ( .A1(n5741), .A2(n9157), .ZN(n9069) );
  INV_X1 U7379 ( .A(n9069), .ZN(n5729) );
  NAND2_X1 U7380 ( .A1(n9727), .A2(n6456), .ZN(n5715) );
  OR2_X1 U7381 ( .A1(n9699), .A2(n6457), .ZN(n5714) );
  NAND2_X1 U7382 ( .A1(n5715), .A2(n5714), .ZN(n5716) );
  XNOR2_X1 U7383 ( .A(n5716), .B(n7330), .ZN(n5731) );
  NOR2_X1 U7384 ( .A1(n9699), .A2(n5592), .ZN(n5717) );
  AOI21_X1 U7385 ( .B1(n9727), .B2(n6463), .A(n5717), .ZN(n5730) );
  XNOR2_X1 U7386 ( .A(n5731), .B(n5730), .ZN(n9072) );
  NAND2_X1 U7387 ( .A1(n9802), .A2(n6456), .ZN(n5719) );
  NAND2_X1 U7388 ( .A1(n9806), .A2(n6463), .ZN(n5718) );
  NAND2_X1 U7389 ( .A1(n5719), .A2(n5718), .ZN(n5720) );
  XNOR2_X1 U7390 ( .A(n5720), .B(n6460), .ZN(n5724) );
  INV_X1 U7391 ( .A(n5724), .ZN(n5722) );
  AND2_X1 U7392 ( .A1(n9806), .A2(n6462), .ZN(n5721) );
  AOI21_X1 U7393 ( .B1(n9802), .B2(n6463), .A(n5721), .ZN(n5723) );
  NAND2_X1 U7394 ( .A1(n5722), .A2(n5723), .ZN(n5732) );
  INV_X1 U7395 ( .A(n5732), .ZN(n5725) );
  XNOR2_X1 U7396 ( .A(n5724), .B(n5723), .ZN(n9082) );
  NOR2_X1 U7397 ( .A1(n5725), .A2(n9082), .ZN(n5734) );
  OR2_X1 U7398 ( .A1(n9072), .A2(n5734), .ZN(n5739) );
  NAND2_X1 U7399 ( .A1(n9685), .A2(n6456), .ZN(n5727) );
  OR2_X1 U7400 ( .A1(n9700), .A2(n6457), .ZN(n5726) );
  NAND2_X1 U7401 ( .A1(n5727), .A2(n5726), .ZN(n5728) );
  XNOR2_X1 U7402 ( .A(n5728), .B(n7330), .ZN(n5744) );
  INV_X1 U7403 ( .A(n5744), .ZN(n5735) );
  NAND2_X1 U7404 ( .A1(n5729), .A2(n4914), .ZN(n9135) );
  NAND2_X1 U7405 ( .A1(n5731), .A2(n5730), .ZN(n9079) );
  AND2_X1 U7406 ( .A1(n9079), .A2(n5732), .ZN(n5733) );
  OR2_X1 U7407 ( .A1(n5734), .A2(n5733), .ZN(n5743) );
  OR2_X1 U7408 ( .A1(n5735), .A2(n5743), .ZN(n9134) );
  NAND2_X1 U7409 ( .A1(n9685), .A2(n6463), .ZN(n5737) );
  OR2_X1 U7410 ( .A1(n9700), .A2(n5592), .ZN(n5736) );
  NAND2_X1 U7411 ( .A1(n5737), .A2(n5736), .ZN(n9138) );
  AND2_X1 U7412 ( .A1(n9134), .A2(n9138), .ZN(n5738) );
  NAND2_X1 U7413 ( .A1(n9135), .A2(n5738), .ZN(n5748) );
  INV_X1 U7414 ( .A(n5739), .ZN(n5740) );
  AND2_X1 U7415 ( .A1(n5740), .A2(n9157), .ZN(n5742) );
  NAND2_X1 U7416 ( .A1(n5742), .A2(n5741), .ZN(n5747) );
  INV_X1 U7417 ( .A(n5743), .ZN(n5745) );
  NOR2_X1 U7418 ( .A1(n5745), .A2(n5744), .ZN(n5746) );
  NAND2_X1 U7419 ( .A1(n5747), .A2(n5746), .ZN(n9133) );
  NAND2_X1 U7420 ( .A1(n9670), .A2(n6456), .ZN(n5750) );
  NAND2_X1 U7421 ( .A1(n9651), .A2(n6463), .ZN(n5749) );
  NAND2_X1 U7422 ( .A1(n5750), .A2(n5749), .ZN(n5751) );
  XNOR2_X1 U7423 ( .A(n5751), .B(n7330), .ZN(n5754) );
  AND2_X1 U7424 ( .A1(n9651), .A2(n6462), .ZN(n5752) );
  AOI21_X1 U7425 ( .B1(n9670), .B2(n6463), .A(n5752), .ZN(n5753) );
  XNOR2_X1 U7426 ( .A(n5754), .B(n5753), .ZN(n9035) );
  NAND2_X1 U7427 ( .A1(n5754), .A2(n5753), .ZN(n5755) );
  NAND2_X1 U7428 ( .A1(n9657), .A2(n6456), .ZN(n5757) );
  NAND2_X1 U7429 ( .A1(n9787), .A2(n6463), .ZN(n5756) );
  NAND2_X1 U7430 ( .A1(n5757), .A2(n5756), .ZN(n5758) );
  XNOR2_X1 U7431 ( .A(n5758), .B(n6460), .ZN(n5761) );
  NAND2_X1 U7432 ( .A1(n9657), .A2(n6463), .ZN(n5760) );
  NAND2_X1 U7433 ( .A1(n9787), .A2(n6462), .ZN(n5759) );
  NAND2_X1 U7434 ( .A1(n5760), .A2(n5759), .ZN(n5762) );
  NAND2_X1 U7435 ( .A1(n5761), .A2(n5762), .ZN(n9101) );
  INV_X1 U7436 ( .A(n5761), .ZN(n5764) );
  INV_X1 U7437 ( .A(n5762), .ZN(n5763) );
  NAND2_X1 U7438 ( .A1(n5764), .A2(n5763), .ZN(n9102) );
  NAND2_X1 U7439 ( .A1(n9772), .A2(n6456), .ZN(n5766) );
  OR2_X1 U7440 ( .A1(n9777), .A2(n6457), .ZN(n5765) );
  NAND2_X1 U7441 ( .A1(n5766), .A2(n5765), .ZN(n5767) );
  XNOR2_X1 U7442 ( .A(n5767), .B(n6460), .ZN(n5775) );
  INV_X1 U7443 ( .A(n5775), .ZN(n5769) );
  NOR2_X1 U7444 ( .A1(n9777), .A2(n5592), .ZN(n5768) );
  AOI21_X1 U7445 ( .B1(n9772), .B2(n6463), .A(n5768), .ZN(n5774) );
  NAND2_X1 U7446 ( .A1(n5769), .A2(n5774), .ZN(n5773) );
  AND2_X1 U7447 ( .A1(n9102), .A2(n5773), .ZN(n5780) );
  AND2_X1 U7448 ( .A1(n9636), .A2(n6462), .ZN(n5770) );
  AOI21_X1 U7449 ( .B1(n9618), .B2(n6463), .A(n5770), .ZN(n5781) );
  INV_X1 U7450 ( .A(n5781), .ZN(n5771) );
  AND2_X1 U7451 ( .A1(n5780), .A2(n5771), .ZN(n5772) );
  INV_X1 U7452 ( .A(n5773), .ZN(n5776) );
  XNOR2_X1 U7453 ( .A(n5775), .B(n5774), .ZN(n9043) );
  OR2_X1 U7454 ( .A1(n5781), .A2(n5782), .ZN(n9121) );
  NAND2_X1 U7455 ( .A1(n9618), .A2(n6456), .ZN(n5778) );
  NAND2_X1 U7456 ( .A1(n9636), .A2(n6463), .ZN(n5777) );
  NAND2_X1 U7457 ( .A1(n5778), .A2(n5777), .ZN(n5779) );
  XNOR2_X1 U7458 ( .A(n5779), .B(n7330), .ZN(n9123) );
  NAND2_X1 U7459 ( .A1(n9122), .A2(n5792), .ZN(n5785) );
  NAND2_X1 U7460 ( .A1(n9041), .A2(n5780), .ZN(n5784) );
  AND2_X1 U7461 ( .A1(n5782), .A2(n5781), .ZN(n5783) );
  NAND2_X1 U7462 ( .A1(n5784), .A2(n5783), .ZN(n9120) );
  NAND2_X1 U7463 ( .A1(n5785), .A2(n9120), .ZN(n5789) );
  NAND2_X1 U7464 ( .A1(n9761), .A2(n6456), .ZN(n5787) );
  NAND2_X1 U7465 ( .A1(n9614), .A2(n6463), .ZN(n5786) );
  NAND2_X1 U7466 ( .A1(n5787), .A2(n5786), .ZN(n5788) );
  XNOR2_X1 U7467 ( .A(n5788), .B(n7330), .ZN(n5793) );
  NAND2_X1 U7468 ( .A1(n5789), .A2(n5793), .ZN(n6517) );
  NAND2_X1 U7469 ( .A1(n9761), .A2(n6463), .ZN(n5791) );
  NAND2_X1 U7470 ( .A1(n9614), .A2(n6462), .ZN(n5790) );
  NAND2_X1 U7471 ( .A1(n5791), .A2(n5790), .ZN(n6518) );
  INV_X1 U7472 ( .A(n9127), .ZN(n5796) );
  INV_X1 U7473 ( .A(n5793), .ZN(n5794) );
  NAND2_X1 U7474 ( .A1(n9756), .A2(n6456), .ZN(n5798) );
  NAND2_X1 U7475 ( .A1(n9600), .A2(n6463), .ZN(n5797) );
  NAND2_X1 U7476 ( .A1(n5798), .A2(n5797), .ZN(n5799) );
  XNOR2_X1 U7477 ( .A(n5799), .B(n7330), .ZN(n5801) );
  NOR2_X1 U7478 ( .A1(n6522), .A2(n5592), .ZN(n5800) );
  AOI21_X1 U7479 ( .B1(n9756), .B2(n6463), .A(n5800), .ZN(n5802) );
  NAND2_X1 U7480 ( .A1(n5801), .A2(n5802), .ZN(n5806) );
  INV_X1 U7481 ( .A(n5801), .ZN(n5804) );
  INV_X1 U7482 ( .A(n5802), .ZN(n5803) );
  NAND2_X1 U7483 ( .A1(n5804), .A2(n5803), .ZN(n5805) );
  NAND2_X1 U7484 ( .A1(n9563), .A2(n6456), .ZN(n5808) );
  NAND2_X1 U7485 ( .A1(n9578), .A2(n6463), .ZN(n5807) );
  NAND2_X1 U7486 ( .A1(n5808), .A2(n5807), .ZN(n5809) );
  XNOR2_X1 U7487 ( .A(n5809), .B(n6460), .ZN(n5814) );
  AOI22_X1 U7488 ( .A1(n9563), .A2(n6463), .B1(n6462), .B2(n9578), .ZN(n5815)
         );
  XNOR2_X1 U7489 ( .A(n5814), .B(n5815), .ZN(n9063) );
  NAND2_X1 U7490 ( .A1(n9265), .A2(n6456), .ZN(n5811) );
  NAND2_X1 U7491 ( .A1(n9560), .A2(n6463), .ZN(n5810) );
  NAND2_X1 U7492 ( .A1(n5811), .A2(n5810), .ZN(n5812) );
  XNOR2_X1 U7493 ( .A(n5812), .B(n6460), .ZN(n5828) );
  AND2_X1 U7494 ( .A1(n9560), .A2(n6462), .ZN(n5813) );
  AOI21_X1 U7495 ( .B1(n9265), .B2(n6463), .A(n5813), .ZN(n5826) );
  XNOR2_X1 U7496 ( .A(n5828), .B(n5826), .ZN(n9149) );
  INV_X1 U7497 ( .A(n5814), .ZN(n5816) );
  NAND2_X1 U7498 ( .A1(n5816), .A2(n5815), .ZN(n9146) );
  NAND2_X1 U7499 ( .A1(n9147), .A2(n5817), .ZN(n9148) );
  NAND2_X1 U7500 ( .A1(n9737), .A2(n6456), .ZN(n5819) );
  OR2_X1 U7501 ( .A1(n9546), .A2(n6457), .ZN(n5818) );
  NAND2_X1 U7502 ( .A1(n5819), .A2(n5818), .ZN(n5820) );
  XNOR2_X1 U7503 ( .A(n5820), .B(n7330), .ZN(n5823) );
  INV_X1 U7504 ( .A(n5823), .ZN(n5825) );
  NOR2_X1 U7505 ( .A1(n9546), .A2(n5592), .ZN(n5821) );
  AOI21_X1 U7506 ( .B1(n9737), .B2(n6463), .A(n5821), .ZN(n5822) );
  INV_X1 U7507 ( .A(n5822), .ZN(n5824) );
  AOI21_X1 U7508 ( .B1(n5825), .B2(n5824), .A(n6470), .ZN(n5829) );
  INV_X1 U7509 ( .A(n5826), .ZN(n5827) );
  NAND2_X1 U7510 ( .A1(n5828), .A2(n5827), .ZN(n5830) );
  AOI21_X1 U7511 ( .B1(n9148), .B2(n5830), .A(n5829), .ZN(n5834) );
  INV_X1 U7512 ( .A(n7127), .ZN(n5831) );
  NAND3_X1 U7513 ( .A1(n9867), .A2(n5831), .A3(n7128), .ZN(n5837) );
  OR2_X1 U7514 ( .A1(n5837), .A2(n7126), .ZN(n5846) );
  OR2_X1 U7515 ( .A1(n9803), .A2(n5832), .ZN(n5833) );
  NOR2_X2 U7516 ( .A1(n5846), .A2(n5833), .ZN(n9160) );
  OAI21_X1 U7517 ( .B1(n6479), .B2(n5834), .A(n9160), .ZN(n5851) );
  INV_X1 U7518 ( .A(n9803), .ZN(n10071) );
  NAND2_X1 U7519 ( .A1(n10071), .A2(n5837), .ZN(n6835) );
  AND3_X1 U7520 ( .A1(n7131), .A2(n5582), .A3(n6489), .ZN(n5835) );
  AOI21_X1 U7521 ( .B1(n6835), .B2(n5835), .A(P1_U3084), .ZN(n5838) );
  OR2_X1 U7522 ( .A1(n10032), .A2(n9443), .ZN(n10031) );
  NOR2_X1 U7523 ( .A1(n10031), .A2(n7126), .ZN(n5836) );
  AND2_X1 U7524 ( .A1(n5837), .A2(n5836), .ZN(n6834) );
  OR2_X1 U7525 ( .A1(n5840), .A2(n5839), .ZN(n6880) );
  NOR2_X1 U7526 ( .A1(n5846), .A2(n6880), .ZN(n5843) );
  NAND2_X1 U7527 ( .A1(n9560), .A2(n9167), .ZN(n5841) );
  OAI21_X1 U7528 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n5842), .A(n5841), .ZN(n5845) );
  NAND2_X1 U7529 ( .A1(n5843), .A2(n5478), .ZN(n9162) );
  NOR2_X1 U7530 ( .A1(n9534), .A2(n9162), .ZN(n5844) );
  AOI211_X1 U7531 ( .C1(n9527), .C2(n9092), .A(n5845), .B(n5844), .ZN(n5850)
         );
  INV_X1 U7532 ( .A(n9737), .ZN(n9529) );
  INV_X1 U7533 ( .A(n5846), .ZN(n5849) );
  INV_X1 U7534 ( .A(n10031), .ZN(n7134) );
  NAND2_X1 U7535 ( .A1(n10051), .A2(n9398), .ZN(n5847) );
  AOI21_X2 U7536 ( .B1(n5849), .B2(n7134), .A(n10035), .ZN(n9170) );
  NAND3_X1 U7537 ( .A1(n5851), .A2(n5850), .A3(n4910), .ZN(P1_U3212) );
  AND2_X2 U7538 ( .A1(n5933), .A2(n5855), .ZN(n5977) );
  INV_X1 U7539 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5866) );
  NAND2_X2 U7540 ( .A1(n6394), .A2(n8223), .ZN(n5944) );
  NAND2_X2 U7541 ( .A1(n5944), .A2(n4389), .ZN(n6031) );
  INV_X2 U7542 ( .A(n6031), .ZN(n6164) );
  NAND2_X1 U7543 ( .A1(n7730), .A2(n6164), .ZN(n5870) );
  INV_X1 U7544 ( .A(n8724), .ZN(n8732) );
  INV_X1 U7545 ( .A(n5878), .ZN(n5874) );
  NAND2_X1 U7546 ( .A1(n5874), .A2(n5861), .ZN(n5876) );
  NAND2_X1 U7547 ( .A1(n5876), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U7548 ( .A1(n5878), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5880) );
  NAND2_X1 U7549 ( .A1(n5880), .A2(n5879), .ZN(n5882) );
  OR2_X1 U7550 ( .A1(n5880), .A2(n5879), .ZN(n5881) );
  NAND2_X1 U7551 ( .A1(n5882), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5883) );
  XNOR2_X1 U7552 ( .A(n8732), .B(n5984), .ZN(n6298) );
  NAND2_X1 U7553 ( .A1(n6000), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7554 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n5885) );
  INV_X1 U7555 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6180) );
  INV_X1 U7556 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6179) );
  AND2_X1 U7557 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n5888) );
  INV_X1 U7558 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8547) );
  INV_X1 U7559 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8606) );
  INV_X1 U7560 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n6281) );
  INV_X1 U7561 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5912) );
  INV_X1 U7562 ( .A(n5914), .ZN(n5892) );
  NAND2_X1 U7563 ( .A1(n5892), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6304) );
  INV_X1 U7564 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8259) );
  NAND2_X1 U7565 ( .A1(n5914), .A2(n8259), .ZN(n5893) );
  NAND2_X1 U7566 ( .A1(n6304), .A2(n5893), .ZN(n8733) );
  NAND2_X1 U7567 ( .A1(n5894), .A2(n5895), .ZN(n5898) );
  OAI21_X1 U7568 ( .B1(n5894), .B2(n4714), .A(P2_IR_REG_29__SCAN_IN), .ZN(
        n5897) );
  NAND2_X1 U7569 ( .A1(n5897), .A2(n5896), .ZN(n5899) );
  NAND2_X2 U7570 ( .A1(n5900), .A2(n5902), .ZN(n5954) );
  OR2_X1 U7571 ( .A1(n8733), .A2(n4398), .ZN(n5907) );
  INV_X1 U7572 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8492) );
  NAND2_X1 U7573 ( .A1(n5901), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5904) );
  AND2_X4 U7574 ( .A1(n8233), .A2(n5902), .ZN(n8087) );
  NAND2_X1 U7575 ( .A1(n8087), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5903) );
  OAI211_X1 U7576 ( .C1(n5968), .C2(n8492), .A(n5904), .B(n5903), .ZN(n5905)
         );
  INV_X1 U7577 ( .A(n5905), .ZN(n5906) );
  NAND2_X1 U7578 ( .A1(n8751), .A2(n8142), .ZN(n6297) );
  NAND2_X1 U7579 ( .A1(n5909), .A2(n6164), .ZN(n5911) );
  XNOR2_X1 U7580 ( .A(n8935), .B(n5984), .ZN(n6293) );
  INV_X1 U7581 ( .A(n6293), .ZN(n8269) );
  NAND2_X1 U7582 ( .A1(n6284), .A2(n5912), .ZN(n5913) );
  AND2_X1 U7583 ( .A1(n5914), .A2(n5913), .ZN(n8743) );
  INV_X1 U7584 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8542) );
  NAND2_X1 U7585 ( .A1(n6395), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5916) );
  NAND2_X1 U7586 ( .A1(n8087), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5915) );
  OAI211_X1 U7587 ( .C1(n8542), .C2(n6569), .A(n5916), .B(n5915), .ZN(n5917)
         );
  AOI21_X1 U7588 ( .B1(n8743), .B2(n6318), .A(n5917), .ZN(n8271) );
  NOR2_X1 U7589 ( .A1(n8271), .A2(n6812), .ZN(n6294) );
  INV_X1 U7590 ( .A(n6294), .ZN(n8273) );
  NAND2_X1 U7591 ( .A1(n8087), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5923) );
  INV_X1 U7592 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n5918) );
  INV_X1 U7593 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6843) );
  OR2_X1 U7594 ( .A1(n5968), .A2(n6843), .ZN(n5921) );
  INV_X1 U7595 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5919) );
  OR2_X1 U7596 ( .A1(n5953), .A2(n5919), .ZN(n5920) );
  NOR2_X1 U7597 ( .A1(n5868), .A2(n5924), .ZN(n5926) );
  INV_X1 U7598 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5925) );
  XNOR2_X1 U7599 ( .A(n5926), .B(n5925), .ZN(n9023) );
  MUX2_X1 U7600 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9023), .S(n5944), .Z(n10191)
         );
  NAND2_X1 U7601 ( .A1(n6896), .A2(n8142), .ZN(n6813) );
  OR2_X1 U7602 ( .A1(n10191), .A2(n5984), .ZN(n5927) );
  NAND2_X1 U7603 ( .A1(n6813), .A2(n5927), .ZN(n6824) );
  NAND2_X1 U7604 ( .A1(n8087), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5932) );
  INV_X1 U7605 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5928) );
  OR2_X1 U7606 ( .A1(n5953), .A2(n5928), .ZN(n5931) );
  INV_X1 U7607 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6642) );
  OR2_X1 U7608 ( .A1(n4396), .A2(n6642), .ZN(n5930) );
  INV_X1 U7609 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6681) );
  INV_X1 U7610 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6537) );
  OR2_X1 U7611 ( .A1(n5943), .A2(n6537), .ZN(n5937) );
  OR2_X1 U7612 ( .A1(n6031), .A2(n6536), .ZN(n5936) );
  INV_X1 U7613 ( .A(n5933), .ZN(n5934) );
  OR2_X1 U7614 ( .A1(n5944), .A2(n6692), .ZN(n5935) );
  INV_X1 U7615 ( .A(n6825), .ZN(n5938) );
  NAND2_X1 U7616 ( .A1(n5939), .A2(n5938), .ZN(n6827) );
  NAND2_X1 U7617 ( .A1(n5941), .A2(n5940), .ZN(n5942) );
  AND2_X1 U7618 ( .A1(n6827), .A2(n5942), .ZN(n6819) );
  OR2_X1 U7619 ( .A1(n6031), .A2(n6541), .ZN(n5951) );
  OR2_X1 U7620 ( .A1(n4394), .A2(n6540), .ZN(n5950) );
  NOR2_X1 U7621 ( .A1(n5933), .A2(n4714), .ZN(n5945) );
  MUX2_X1 U7622 ( .A(n4714), .B(n5945), .S(P2_IR_REG_2__SCAN_IN), .Z(n5946) );
  INV_X1 U7623 ( .A(n5946), .ZN(n5948) );
  INV_X1 U7624 ( .A(n5977), .ZN(n5947) );
  NAND2_X1 U7625 ( .A1(n5948), .A2(n5947), .ZN(n6717) );
  OR2_X1 U7626 ( .A1(n5944), .A2(n6717), .ZN(n5949) );
  XNOR2_X1 U7627 ( .A(n10195), .B(n5984), .ZN(n10105) );
  INV_X1 U7628 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5952) );
  OR2_X1 U7629 ( .A1(n5953), .A2(n5952), .ZN(n5957) );
  INV_X1 U7630 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6643) );
  OR2_X1 U7631 ( .A1(n5968), .A2(n6643), .ZN(n5956) );
  INV_X1 U7632 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6706) );
  OR2_X1 U7633 ( .A1(n4397), .A2(n6706), .ZN(n5955) );
  NAND2_X1 U7634 ( .A1(n10111), .A2(n8142), .ZN(n5959) );
  OR2_X1 U7635 ( .A1(n10105), .A2(n5959), .ZN(n5961) );
  NAND2_X1 U7636 ( .A1(n5959), .A2(n10105), .ZN(n5960) );
  AND2_X1 U7637 ( .A1(n5961), .A2(n5960), .ZN(n6818) );
  NAND2_X1 U7638 ( .A1(n6819), .A2(n6818), .ZN(n6817) );
  NAND2_X1 U7639 ( .A1(n6817), .A2(n5961), .ZN(n5975) );
  OR2_X1 U7640 ( .A1(n6031), .A2(n6549), .ZN(n5965) );
  INV_X1 U7641 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6548) );
  OR2_X1 U7642 ( .A1(n5977), .A2(n4714), .ZN(n5962) );
  XNOR2_X1 U7643 ( .A(n5962), .B(n5976), .ZN(n6666) );
  OR2_X1 U7644 ( .A1(n5944), .A2(n6666), .ZN(n5963) );
  XNOR2_X1 U7645 ( .A(n6912), .B(n5984), .ZN(n8286) );
  NAND2_X1 U7646 ( .A1(n8087), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5972) );
  INV_X1 U7647 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5966) );
  INV_X1 U7648 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5967) );
  INV_X1 U7649 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6645) );
  OR2_X1 U7650 ( .A1(n5968), .A2(n6645), .ZN(n5969) );
  NAND2_X1 U7651 ( .A1(n8337), .A2(n8142), .ZN(n5973) );
  OR2_X1 U7652 ( .A1(n8286), .A2(n5973), .ZN(n5993) );
  NAND2_X1 U7653 ( .A1(n5973), .A2(n8286), .ZN(n5974) );
  AND2_X1 U7654 ( .A1(n5993), .A2(n5974), .ZN(n10107) );
  NAND2_X1 U7655 ( .A1(n5975), .A2(n10107), .ZN(n8282) );
  OR2_X1 U7656 ( .A1(n6539), .A2(n6031), .ZN(n5983) );
  NAND2_X1 U7657 ( .A1(n5977), .A2(n5976), .ZN(n5979) );
  NAND2_X1 U7658 ( .A1(n5979), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5978) );
  MUX2_X1 U7659 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5978), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5980) );
  NAND2_X1 U7660 ( .A1(n5980), .A2(n6013), .ZN(n6705) );
  OR2_X1 U7661 ( .A1(n5944), .A2(n6705), .ZN(n5982) );
  XNOR2_X1 U7662 ( .A(n10202), .B(n6301), .ZN(n5995) );
  NAND2_X1 U7663 ( .A1(n6395), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5992) );
  INV_X1 U7664 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6633) );
  OR2_X1 U7665 ( .A1(n6322), .A2(n6633), .ZN(n5991) );
  INV_X1 U7666 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5985) );
  OR2_X1 U7667 ( .A1(n5953), .A2(n5985), .ZN(n5990) );
  INV_X1 U7668 ( .A(n6000), .ZN(n5988) );
  INV_X1 U7669 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7670 ( .A1(n5966), .A2(n5986), .ZN(n5987) );
  NAND2_X1 U7671 ( .A1(n5988), .A2(n5987), .ZN(n8279) );
  OR2_X1 U7672 ( .A1(n4397), .A2(n8279), .ZN(n5989) );
  NAND2_X1 U7673 ( .A1(n10139), .A2(n8142), .ZN(n5997) );
  XNOR2_X1 U7674 ( .A(n5995), .B(n5997), .ZN(n8285) );
  AND2_X1 U7675 ( .A1(n8285), .A2(n5993), .ZN(n5994) );
  INV_X1 U7676 ( .A(n5995), .ZN(n5996) );
  NAND2_X1 U7677 ( .A1(n5997), .A2(n5996), .ZN(n5998) );
  NAND2_X1 U7678 ( .A1(n6395), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6004) );
  INV_X1 U7679 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5999) );
  OR2_X1 U7680 ( .A1(n6322), .A2(n5999), .ZN(n6003) );
  OAI21_X1 U7681 ( .B1(n6000), .B2(P2_REG3_REG_5__SCAN_IN), .A(n6018), .ZN(
        n10151) );
  INV_X1 U7682 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6001) );
  NOR2_X1 U7683 ( .A1(n7155), .A2(n6812), .ZN(n6008) );
  OR2_X1 U7684 ( .A1(n6547), .A2(n6031), .ZN(n6007) );
  NAND2_X1 U7685 ( .A1(n6013), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6005) );
  XNOR2_X1 U7686 ( .A(n6005), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6669) );
  AOI22_X1 U7687 ( .A1(n6227), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6556), .B2(
        n6669), .ZN(n6006) );
  NAND2_X1 U7688 ( .A1(n6007), .A2(n6006), .ZN(n10135) );
  XNOR2_X1 U7689 ( .A(n10135), .B(n5984), .ZN(n6009) );
  NAND2_X1 U7690 ( .A1(n6008), .A2(n6009), .ZN(n6025) );
  INV_X1 U7691 ( .A(n6008), .ZN(n6010) );
  INV_X1 U7692 ( .A(n6009), .ZN(n8314) );
  NAND2_X1 U7693 ( .A1(n6010), .A2(n8314), .ZN(n6011) );
  NAND2_X1 U7694 ( .A1(n6025), .A2(n6011), .ZN(n10141) );
  INV_X1 U7695 ( .A(n10141), .ZN(n6012) );
  OR2_X1 U7696 ( .A1(n6545), .A2(n6031), .ZN(n6016) );
  OR2_X1 U7697 ( .A1(n6033), .A2(n4714), .ZN(n6014) );
  XNOR2_X1 U7698 ( .A(n6014), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6676) );
  AOI22_X1 U7699 ( .A1(n6227), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6556), .B2(
        n6676), .ZN(n6015) );
  NAND2_X1 U7700 ( .A1(n6016), .A2(n6015), .ZN(n10214) );
  XNOR2_X1 U7701 ( .A(n10214), .B(n5984), .ZN(n6027) );
  NAND2_X1 U7702 ( .A1(n8087), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6024) );
  INV_X1 U7703 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n8882) );
  OR2_X1 U7704 ( .A1(n5968), .A2(n8882), .ZN(n6023) );
  AND2_X1 U7705 ( .A1(n6018), .A2(n6017), .ZN(n6019) );
  OR2_X1 U7706 ( .A1(n6019), .A2(n6037), .ZN(n8887) );
  OR2_X1 U7707 ( .A1(n4397), .A2(n8887), .ZN(n6022) );
  INV_X1 U7708 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6020) );
  OR2_X1 U7709 ( .A1(n6569), .A2(n6020), .ZN(n6021) );
  OR2_X1 U7710 ( .A1(n7102), .A2(n6812), .ZN(n6028) );
  XNOR2_X1 U7711 ( .A(n6027), .B(n6028), .ZN(n8313) );
  AND2_X1 U7712 ( .A1(n8313), .A2(n6025), .ZN(n6026) );
  NAND2_X1 U7713 ( .A1(n10144), .A2(n6026), .ZN(n8311) );
  INV_X1 U7714 ( .A(n6027), .ZN(n6029) );
  NAND2_X1 U7715 ( .A1(n6029), .A2(n6028), .ZN(n6030) );
  OR2_X1 U7716 ( .A1(n6543), .A2(n6031), .ZN(n6036) );
  NAND2_X1 U7717 ( .A1(n6033), .A2(n6032), .ZN(n6049) );
  NAND2_X1 U7718 ( .A1(n6049), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6034) );
  XNOR2_X1 U7719 ( .A(n6034), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6748) );
  AOI22_X1 U7720 ( .A1(n6227), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6556), .B2(
        n6748), .ZN(n6035) );
  NAND2_X1 U7721 ( .A1(n6036), .A2(n6035), .ZN(n10085) );
  XNOR2_X1 U7722 ( .A(n10085), .B(n5984), .ZN(n10117) );
  NAND2_X1 U7723 ( .A1(n8087), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6043) );
  NOR2_X1 U7724 ( .A1(n6037), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6038) );
  OR2_X1 U7725 ( .A1(n6067), .A2(n6038), .ZN(n10092) );
  OR2_X1 U7726 ( .A1(n4397), .A2(n10092), .ZN(n6042) );
  INV_X1 U7727 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6039) );
  OR2_X1 U7728 ( .A1(n5953), .A2(n6039), .ZN(n6041) );
  INV_X1 U7729 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7094) );
  OR2_X1 U7730 ( .A1(n5968), .A2(n7094), .ZN(n6040) );
  NOR2_X1 U7731 ( .A1(n7168), .A2(n6812), .ZN(n6044) );
  NAND2_X1 U7732 ( .A1(n10117), .A2(n6044), .ZN(n6048) );
  INV_X1 U7733 ( .A(n10117), .ZN(n6046) );
  INV_X1 U7734 ( .A(n6044), .ZN(n6045) );
  NAND2_X1 U7735 ( .A1(n6046), .A2(n6045), .ZN(n6047) );
  AND2_X1 U7736 ( .A1(n6048), .A2(n6047), .ZN(n10086) );
  NAND2_X1 U7737 ( .A1(n6550), .A2(n6164), .ZN(n6054) );
  NAND2_X1 U7738 ( .A1(n6051), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6050) );
  MUX2_X1 U7739 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6050), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n6052) );
  NAND2_X1 U7740 ( .A1(n6052), .A2(n6081), .ZN(n6935) );
  INV_X1 U7741 ( .A(n6935), .ZN(n6928) );
  AOI22_X1 U7742 ( .A1(n6227), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6556), .B2(
        n6928), .ZN(n6053) );
  NAND2_X1 U7743 ( .A1(n6054), .A2(n6053), .ZN(n10125) );
  XNOR2_X1 U7744 ( .A(n10125), .B(n5984), .ZN(n6060) );
  NAND2_X1 U7745 ( .A1(n8087), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6059) );
  XNOR2_X1 U7746 ( .A(n6067), .B(P2_REG3_REG_8__SCAN_IN), .ZN(n10134) );
  OR2_X1 U7747 ( .A1(n4398), .A2(n10134), .ZN(n6058) );
  INV_X1 U7748 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6055) );
  OR2_X1 U7749 ( .A1(n6569), .A2(n6055), .ZN(n6057) );
  INV_X1 U7750 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7180) );
  OR2_X1 U7751 ( .A1(n5968), .A2(n7180), .ZN(n6056) );
  NOR2_X1 U7752 ( .A1(n7268), .A2(n6812), .ZN(n6061) );
  NAND2_X1 U7753 ( .A1(n6060), .A2(n6061), .ZN(n6074) );
  INV_X1 U7754 ( .A(n6060), .ZN(n7013) );
  INV_X1 U7755 ( .A(n6061), .ZN(n6062) );
  NAND2_X1 U7756 ( .A1(n7013), .A2(n6062), .ZN(n6063) );
  AND2_X1 U7757 ( .A1(n6074), .A2(n6063), .ZN(n10120) );
  NAND2_X1 U7758 ( .A1(n6553), .A2(n6164), .ZN(n6066) );
  NAND2_X1 U7759 ( .A1(n6081), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6064) );
  XNOR2_X1 U7760 ( .A(n6064), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6984) );
  AOI22_X1 U7761 ( .A1(n6227), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6556), .B2(
        n6984), .ZN(n6065) );
  NAND2_X2 U7762 ( .A1(n6066), .A2(n6065), .ZN(n7341) );
  XNOR2_X1 U7763 ( .A(n7341), .B(n6301), .ZN(n6078) );
  NAND2_X1 U7764 ( .A1(n8087), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6073) );
  INV_X1 U7765 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7278) );
  OR2_X1 U7766 ( .A1(n5968), .A2(n7278), .ZN(n6072) );
  AOI21_X1 U7767 ( .B1(n6067), .B2(P2_REG3_REG_8__SCAN_IN), .A(
        P2_REG3_REG_9__SCAN_IN), .ZN(n6068) );
  OR2_X1 U7768 ( .A1(n6084), .A2(n6068), .ZN(n7277) );
  OR2_X1 U7769 ( .A1(n4397), .A2(n7277), .ZN(n6071) );
  INV_X1 U7770 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n6069) );
  OR2_X1 U7771 ( .A1(n6569), .A2(n6069), .ZN(n6070) );
  NOR2_X1 U7772 ( .A1(n10129), .A2(n6812), .ZN(n6076) );
  XNOR2_X1 U7773 ( .A(n6078), .B(n6076), .ZN(n7022) );
  AND2_X1 U7774 ( .A1(n7022), .A2(n6074), .ZN(n6075) );
  NAND2_X1 U7775 ( .A1(n7012), .A2(n6075), .ZN(n7015) );
  INV_X1 U7776 ( .A(n6076), .ZN(n6077) );
  NAND2_X1 U7777 ( .A1(n6078), .A2(n6077), .ZN(n6079) );
  NAND2_X1 U7778 ( .A1(n7015), .A2(n6079), .ZN(n10099) );
  NAND2_X1 U7779 ( .A1(n6080), .A2(n6164), .ZN(n6083) );
  OR2_X1 U7780 ( .A1(n6115), .A2(n4714), .ZN(n6099) );
  XNOR2_X1 U7781 ( .A(n6099), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7071) );
  AOI22_X1 U7782 ( .A1(n7071), .A2(n6556), .B1(n6227), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n6082) );
  XNOR2_X1 U7783 ( .A(n7345), .B(n5984), .ZN(n6092) );
  NAND2_X1 U7784 ( .A1(n8087), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6091) );
  INV_X1 U7785 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7357) );
  OR2_X1 U7786 ( .A1(n5968), .A2(n7357), .ZN(n6090) );
  INV_X1 U7787 ( .A(n6084), .ZN(n6085) );
  INV_X1 U7788 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8483) );
  NAND2_X1 U7789 ( .A1(n6085), .A2(n8483), .ZN(n6086) );
  NAND2_X1 U7790 ( .A1(n6121), .A2(n6086), .ZN(n10104) );
  OR2_X1 U7791 ( .A1(n4398), .A2(n10104), .ZN(n6089) );
  INV_X1 U7792 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n6087) );
  OR2_X1 U7793 ( .A1(n6569), .A2(n6087), .ZN(n6088) );
  AND4_X2 U7794 ( .A1(n6091), .A2(n6090), .A3(n6089), .A4(n6088), .ZN(n7405)
         );
  NOR2_X1 U7795 ( .A1(n7405), .A2(n6812), .ZN(n6093) );
  NAND2_X1 U7796 ( .A1(n6092), .A2(n6093), .ZN(n6097) );
  INV_X1 U7797 ( .A(n6092), .ZN(n7118) );
  INV_X1 U7798 ( .A(n6093), .ZN(n6094) );
  NAND2_X1 U7799 ( .A1(n7118), .A2(n6094), .ZN(n6095) );
  NAND2_X1 U7800 ( .A1(n6097), .A2(n6095), .ZN(n10100) );
  INV_X1 U7801 ( .A(n10100), .ZN(n6096) );
  NAND2_X1 U7802 ( .A1(n6562), .A2(n6164), .ZN(n6103) );
  INV_X1 U7803 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7804 ( .A1(n6099), .A2(n6098), .ZN(n6100) );
  NAND2_X1 U7805 ( .A1(n6100), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6101) );
  XNOR2_X1 U7806 ( .A(n6101), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7253) );
  AOI22_X1 U7807 ( .A1(n7253), .A2(n6556), .B1(n6227), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n6102) );
  XNOR2_X1 U7808 ( .A(n7562), .B(n6301), .ZN(n6109) );
  NAND2_X1 U7809 ( .A1(n8087), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6108) );
  INV_X1 U7810 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7420) );
  OR2_X1 U7811 ( .A1(n5968), .A2(n7420), .ZN(n6107) );
  INV_X1 U7812 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6120) );
  XNOR2_X1 U7813 ( .A(n6121), .B(n6120), .ZN(n7419) );
  OR2_X1 U7814 ( .A1(n4398), .A2(n7419), .ZN(n6106) );
  INV_X1 U7815 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n6104) );
  OR2_X1 U7816 ( .A1(n6569), .A2(n6104), .ZN(n6105) );
  NOR2_X1 U7817 ( .A1(n7561), .A2(n6812), .ZN(n6110) );
  XNOR2_X1 U7818 ( .A(n6109), .B(n6110), .ZN(n7116) );
  INV_X1 U7819 ( .A(n6109), .ZN(n6111) );
  NAND2_X1 U7820 ( .A1(n6111), .A2(n6110), .ZN(n6112) );
  NAND2_X1 U7821 ( .A1(n7119), .A2(n6112), .ZN(n7295) );
  NAND2_X1 U7822 ( .A1(n6113), .A2(n6164), .ZN(n6118) );
  NAND2_X1 U7823 ( .A1(n6115), .A2(n6114), .ZN(n6133) );
  NAND2_X1 U7824 ( .A1(n6133), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6116) );
  XNOR2_X1 U7825 ( .A(n6116), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7433) );
  AOI22_X1 U7826 ( .A1(n7433), .A2(n6556), .B1(n6227), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n6117) );
  XNOR2_X1 U7827 ( .A(n10162), .B(n6301), .ZN(n6128) );
  NAND2_X1 U7828 ( .A1(n6395), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6127) );
  INV_X1 U7829 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7254) );
  OR2_X1 U7830 ( .A1(n6322), .A2(n7254), .ZN(n6126) );
  INV_X1 U7831 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6119) );
  OAI21_X1 U7832 ( .B1(n6121), .B2(n6120), .A(n6119), .ZN(n6122) );
  NAND2_X1 U7833 ( .A1(n6122), .A2(n6137), .ZN(n10158) );
  OR2_X1 U7834 ( .A1(n4397), .A2(n10158), .ZN(n6125) );
  INV_X1 U7835 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n6123) );
  OR2_X1 U7836 ( .A1(n5953), .A2(n6123), .ZN(n6124) );
  OR2_X1 U7837 ( .A1(n7576), .A2(n6812), .ZN(n6129) );
  NAND2_X1 U7838 ( .A1(n6128), .A2(n6129), .ZN(n7294) );
  NAND2_X1 U7839 ( .A1(n7295), .A2(n7294), .ZN(n6132) );
  INV_X1 U7840 ( .A(n6128), .ZN(n6131) );
  INV_X1 U7841 ( .A(n6129), .ZN(n6130) );
  NAND2_X1 U7842 ( .A1(n6131), .A2(n6130), .ZN(n7293) );
  NAND2_X1 U7843 ( .A1(n6132), .A2(n7293), .ZN(n7362) );
  NAND2_X1 U7844 ( .A1(n6743), .A2(n6164), .ZN(n6136) );
  NAND2_X1 U7845 ( .A1(n6134), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6148) );
  XNOR2_X1 U7846 ( .A(n6148), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7512) );
  AOI22_X1 U7847 ( .A1(n7512), .A2(n6556), .B1(n6227), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n6135) );
  XNOR2_X1 U7848 ( .A(n8033), .B(n6301), .ZN(n6143) );
  NAND2_X1 U7849 ( .A1(n5901), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6142) );
  INV_X1 U7850 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7582) );
  OR2_X1 U7851 ( .A1(n5968), .A2(n7582), .ZN(n6141) );
  INV_X1 U7852 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7614) );
  OR2_X1 U7853 ( .A1(n6322), .A2(n7614), .ZN(n6140) );
  INV_X1 U7854 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U7855 ( .A1(n6137), .A2(n8638), .ZN(n6138) );
  NAND2_X1 U7856 ( .A1(n6181), .A2(n6138), .ZN(n7581) );
  OR2_X1 U7857 ( .A1(n4397), .A2(n7581), .ZN(n6139) );
  NOR2_X1 U7858 ( .A1(n8032), .A2(n6812), .ZN(n6144) );
  XNOR2_X1 U7859 ( .A(n6143), .B(n6144), .ZN(n7363) );
  INV_X1 U7860 ( .A(n6143), .ZN(n6145) );
  NAND2_X1 U7861 ( .A1(n6145), .A2(n6144), .ZN(n6146) );
  NAND2_X1 U7862 ( .A1(n6760), .A2(n6164), .ZN(n6151) );
  INV_X1 U7863 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7864 ( .A1(n6148), .A2(n6147), .ZN(n6149) );
  NAND2_X1 U7865 ( .A1(n6149), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6174) );
  XNOR2_X1 U7866 ( .A(n6174), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7829) );
  AOI22_X1 U7867 ( .A1(n7829), .A2(n6556), .B1(n6227), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n6150) );
  XNOR2_X1 U7868 ( .A(n8989), .B(n6301), .ZN(n6157) );
  NAND2_X1 U7869 ( .A1(n5901), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6156) );
  INV_X1 U7870 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7510) );
  OR2_X1 U7871 ( .A1(n6322), .A2(n7510), .ZN(n6155) );
  INV_X1 U7872 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6152) );
  OR2_X1 U7873 ( .A1(n5968), .A2(n6152), .ZN(n6154) );
  XNOR2_X1 U7874 ( .A(n6181), .B(n6180), .ZN(n7555) );
  OR2_X1 U7875 ( .A1(n4398), .A2(n7555), .ZN(n6153) );
  OR2_X1 U7876 ( .A1(n7711), .A2(n6812), .ZN(n6158) );
  NAND2_X1 U7877 ( .A1(n6157), .A2(n6158), .ZN(n6163) );
  INV_X1 U7878 ( .A(n6157), .ZN(n6160) );
  INV_X1 U7879 ( .A(n6158), .ZN(n6159) );
  NAND2_X1 U7880 ( .A1(n6160), .A2(n6159), .ZN(n6161) );
  NAND2_X1 U7881 ( .A1(n6163), .A2(n6161), .ZN(n7554) );
  NAND2_X1 U7882 ( .A1(n7551), .A2(n6163), .ZN(n7687) );
  NAND2_X1 U7883 ( .A1(n6942), .A2(n6164), .ZN(n6167) );
  NAND2_X1 U7884 ( .A1(n6353), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6165) );
  XNOR2_X1 U7885 ( .A(n6165), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8345) );
  AOI22_X1 U7886 ( .A1(n6227), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6556), .B2(
        n8345), .ZN(n6166) );
  XNOR2_X1 U7887 ( .A(n8980), .B(n5984), .ZN(n6193) );
  INV_X1 U7888 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7815) );
  OR2_X1 U7889 ( .A1(n5968), .A2(n7815), .ZN(n6172) );
  INV_X1 U7890 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8649) );
  OR2_X1 U7891 ( .A1(n6322), .A2(n8649), .ZN(n6171) );
  INV_X1 U7892 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7899) );
  NAND2_X1 U7893 ( .A1(n6182), .A2(n7899), .ZN(n6168) );
  NAND2_X1 U7894 ( .A1(n6215), .A2(n6168), .ZN(n7814) );
  OR2_X1 U7895 ( .A1(n4397), .A2(n7814), .ZN(n6170) );
  INV_X1 U7896 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8632) );
  OR2_X1 U7897 ( .A1(n6569), .A2(n8632), .ZN(n6169) );
  NOR2_X1 U7898 ( .A1(n8857), .A2(n6812), .ZN(n6194) );
  NAND2_X1 U7899 ( .A1(n6193), .A2(n6194), .ZN(n7777) );
  NAND2_X1 U7900 ( .A1(n6940), .A2(n6164), .ZN(n6178) );
  INV_X1 U7901 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7902 ( .A1(n6174), .A2(n6173), .ZN(n6175) );
  NAND2_X1 U7903 ( .A1(n6175), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6176) );
  XNOR2_X1 U7904 ( .A(n6176), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7893) );
  AOI21_X1 U7905 ( .B1(n7893), .B2(n6556), .A(n4457), .ZN(n6177) );
  XNOR2_X1 U7906 ( .A(n8984), .B(n5984), .ZN(n6191) );
  NAND2_X1 U7907 ( .A1(n6395), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6188) );
  INV_X1 U7908 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7827) );
  OR2_X1 U7909 ( .A1(n6322), .A2(n7827), .ZN(n6187) );
  OAI21_X1 U7910 ( .B1(n6181), .B2(n6180), .A(n6179), .ZN(n6183) );
  NAND2_X1 U7911 ( .A1(n6183), .A2(n6182), .ZN(n7874) );
  OR2_X1 U7912 ( .A1(n4398), .A2(n7874), .ZN(n6186) );
  INV_X1 U7913 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n6184) );
  OR2_X1 U7914 ( .A1(n6569), .A2(n6184), .ZN(n6185) );
  NOR2_X1 U7915 ( .A1(n7800), .A2(n6812), .ZN(n6192) );
  NAND2_X1 U7916 ( .A1(n6191), .A2(n6192), .ZN(n6189) );
  AND2_X1 U7917 ( .A1(n7777), .A2(n6189), .ZN(n6190) );
  INV_X1 U7918 ( .A(n6191), .ZN(n7778) );
  INV_X1 U7919 ( .A(n6192), .ZN(n7779) );
  NAND3_X1 U7920 ( .A1(n7777), .A2(n7778), .A3(n7779), .ZN(n6197) );
  INV_X1 U7921 ( .A(n6193), .ZN(n6196) );
  INV_X1 U7922 ( .A(n6194), .ZN(n6195) );
  NAND2_X1 U7923 ( .A1(n6196), .A2(n6195), .ZN(n7776) );
  AND2_X1 U7924 ( .A1(n6197), .A2(n7776), .ZN(n6198) );
  NAND2_X1 U7925 ( .A1(n6952), .A2(n6164), .ZN(n6201) );
  NAND2_X1 U7926 ( .A1(n4466), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6199) );
  XNOR2_X1 U7927 ( .A(n6199), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8358) );
  AOI22_X1 U7928 ( .A1(n6227), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6556), .B2(
        n8358), .ZN(n6200) );
  XNOR2_X1 U7929 ( .A(n8975), .B(n5984), .ZN(n6208) );
  INV_X1 U7930 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n6202) );
  OR2_X1 U7931 ( .A1(n6322), .A2(n6202), .ZN(n6206) );
  INV_X1 U7932 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8868) );
  OR2_X1 U7933 ( .A1(n5968), .A2(n8868), .ZN(n6205) );
  INV_X1 U7934 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8652) );
  XNOR2_X1 U7935 ( .A(n6215), .B(n8652), .ZN(n8867) );
  OR2_X1 U7936 ( .A1(n4398), .A2(n8867), .ZN(n6204) );
  INV_X1 U7937 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8596) );
  OR2_X1 U7938 ( .A1(n6569), .A2(n8596), .ZN(n6203) );
  NOR2_X1 U7939 ( .A1(n7963), .A2(n6812), .ZN(n6207) );
  XNOR2_X1 U7940 ( .A(n6208), .B(n6207), .ZN(n7625) );
  NAND2_X1 U7941 ( .A1(n6208), .A2(n6207), .ZN(n6209) );
  NAND2_X1 U7942 ( .A1(n7024), .A2(n6164), .ZN(n6213) );
  NAND2_X1 U7943 ( .A1(n6210), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6211) );
  XNOR2_X1 U7944 ( .A(n6211), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8375) );
  AOI22_X1 U7945 ( .A1(n6227), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6556), .B2(
        n8375), .ZN(n6212) );
  XNOR2_X1 U7946 ( .A(n8838), .B(n5984), .ZN(n6222) );
  INV_X1 U7947 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8359) );
  OR2_X1 U7948 ( .A1(n6322), .A2(n8359), .ZN(n6221) );
  INV_X1 U7949 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8531) );
  OR2_X1 U7950 ( .A1(n6569), .A2(n8531), .ZN(n6220) );
  INV_X1 U7951 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6214) );
  OAI21_X1 U7952 ( .B1(n6215), .B2(n8652), .A(n6214), .ZN(n6216) );
  NAND2_X1 U7953 ( .A1(n6216), .A2(n6230), .ZN(n7771) );
  OR2_X1 U7954 ( .A1(n4397), .A2(n7771), .ZN(n6219) );
  INV_X1 U7955 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n6217) );
  OR2_X1 U7956 ( .A1(n4396), .A2(n6217), .ZN(n6218) );
  NOR2_X1 U7957 ( .A1(n8859), .A2(n6812), .ZN(n6223) );
  XNOR2_X1 U7958 ( .A(n6222), .B(n6223), .ZN(n7770) );
  INV_X1 U7959 ( .A(n6222), .ZN(n6224) );
  NAND2_X1 U7960 ( .A1(n6224), .A2(n6223), .ZN(n6225) );
  NAND2_X1 U7961 ( .A1(n6226), .A2(n6225), .ZN(n7852) );
  INV_X1 U7962 ( .A(n7852), .ZN(n6242) );
  NAND2_X1 U7963 ( .A1(n7060), .A2(n6164), .ZN(n6229) );
  AOI22_X1 U7964 ( .A1(n6227), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8734), .B2(
        n6556), .ZN(n6228) );
  XNOR2_X1 U7965 ( .A(n8820), .B(n6301), .ZN(n6237) );
  NAND2_X1 U7966 ( .A1(n6230), .A2(n8547), .ZN(n6231) );
  AND2_X1 U7967 ( .A1(n6246), .A2(n6231), .ZN(n8817) );
  NAND2_X1 U7968 ( .A1(n8817), .A2(n6318), .ZN(n6236) );
  NAND2_X1 U7969 ( .A1(n6395), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6235) );
  NAND2_X1 U7970 ( .A1(n5901), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6234) );
  INV_X1 U7971 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n6232) );
  OR2_X1 U7972 ( .A1(n6322), .A2(n6232), .ZN(n6233) );
  NOR2_X1 U7973 ( .A1(n8293), .A2(n6812), .ZN(n6238) );
  AND2_X1 U7974 ( .A1(n6237), .A2(n6238), .ZN(n7853) );
  INV_X1 U7975 ( .A(n6237), .ZN(n6240) );
  INV_X1 U7976 ( .A(n6238), .ZN(n6239) );
  NAND2_X1 U7977 ( .A1(n7228), .A2(n6164), .ZN(n6244) );
  XNOR2_X1 U7978 ( .A(n8958), .B(n5984), .ZN(n6251) );
  INV_X1 U7979 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U7980 ( .A1(n6246), .A2(n6245), .ZN(n6247) );
  NAND2_X1 U7981 ( .A1(n6258), .A2(n6247), .ZN(n8811) );
  OR2_X1 U7982 ( .A1(n8811), .A2(n4397), .ZN(n6250) );
  AOI22_X1 U7983 ( .A1(n8087), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n6395), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n6249) );
  NAND2_X1 U7984 ( .A1(n5901), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6248) );
  NOR2_X1 U7985 ( .A1(n8827), .A2(n6812), .ZN(n6252) );
  NAND2_X1 U7986 ( .A1(n6251), .A2(n6252), .ZN(n6255) );
  INV_X1 U7987 ( .A(n6251), .ZN(n8247) );
  INV_X1 U7988 ( .A(n6252), .ZN(n6253) );
  NAND2_X1 U7989 ( .A1(n8247), .A2(n6253), .ZN(n6254) );
  AND2_X1 U7990 ( .A1(n6255), .A2(n6254), .ZN(n8291) );
  NAND2_X1 U7991 ( .A1(n7304), .A2(n6164), .ZN(n6257) );
  XNOR2_X1 U7992 ( .A(n8952), .B(n5984), .ZN(n6264) );
  NAND2_X1 U7993 ( .A1(n6258), .A2(n8606), .ZN(n6259) );
  NAND2_X1 U7994 ( .A1(n6269), .A2(n6259), .ZN(n8789) );
  AOI22_X1 U7995 ( .A1(n8087), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n6395), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n6261) );
  NAND2_X1 U7996 ( .A1(n5901), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6260) );
  OAI211_X1 U7997 ( .C1(n8789), .C2(n4398), .A(n6261), .B(n6260), .ZN(n8804)
         );
  NAND2_X1 U7998 ( .A1(n8804), .A2(n8142), .ZN(n6262) );
  INV_X1 U7999 ( .A(n6262), .ZN(n6263) );
  NAND2_X1 U8000 ( .A1(n6264), .A2(n6263), .ZN(n6265) );
  NAND2_X1 U8001 ( .A1(n7426), .A2(n6164), .ZN(n6267) );
  XNOR2_X1 U8002 ( .A(n8946), .B(n6301), .ZN(n6274) );
  INV_X1 U8003 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n6268) );
  NAND2_X1 U8004 ( .A1(n6269), .A2(n6268), .ZN(n6270) );
  NAND2_X1 U8005 ( .A1(n6282), .A2(n6270), .ZN(n8302) );
  OR2_X1 U8006 ( .A1(n8302), .A2(n4397), .ZN(n6273) );
  AOI22_X1 U8007 ( .A1(n8087), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n6395), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n6272) );
  INV_X1 U8008 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8484) );
  OR2_X1 U8009 ( .A1(n6569), .A2(n8484), .ZN(n6271) );
  OR2_X1 U8010 ( .A1(n8251), .A2(n6812), .ZN(n8298) );
  INV_X1 U8011 ( .A(n6274), .ZN(n6275) );
  NOR2_X1 U8012 ( .A1(n6276), .A2(n6275), .ZN(n6277) );
  NAND2_X1 U8013 ( .A1(n7502), .A2(n6164), .ZN(n6279) );
  XNOR2_X1 U8014 ( .A(n8940), .B(n5984), .ZN(n6291) );
  INV_X1 U8015 ( .A(n8271), .ZN(n8729) );
  OR2_X1 U8016 ( .A1(n6293), .A2(n8729), .ZN(n6290) );
  NAND2_X1 U8017 ( .A1(n6282), .A2(n6281), .ZN(n6283) );
  NAND2_X1 U8018 ( .A1(n6284), .A2(n6283), .ZN(n8764) );
  OR2_X1 U8019 ( .A1(n8764), .A2(n4397), .ZN(n6289) );
  INV_X1 U8020 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8623) );
  NAND2_X1 U8021 ( .A1(n6395), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6286) );
  NAND2_X1 U8022 ( .A1(n5901), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6285) );
  OAI211_X1 U8023 ( .C1(n6322), .C2(n8623), .A(n6286), .B(n6285), .ZN(n6287)
         );
  INV_X1 U8024 ( .A(n6287), .ZN(n6288) );
  NOR2_X1 U8025 ( .A1(n8236), .A2(n6812), .ZN(n8237) );
  AND2_X1 U8026 ( .A1(n6292), .A2(n6291), .ZN(n8267) );
  OAI21_X1 U8027 ( .B1(n6294), .B2(n6293), .A(n8267), .ZN(n6295) );
  OAI211_X1 U8028 ( .C1(n8269), .C2(n8273), .A(n6296), .B(n6295), .ZN(n8257)
         );
  XNOR2_X1 U8029 ( .A(n6298), .B(n6297), .ZN(n8258) );
  NAND2_X1 U8030 ( .A1(n7787), .A2(n6164), .ZN(n6300) );
  XNOR2_X1 U8031 ( .A(n8926), .B(n6301), .ZN(n8192) );
  INV_X1 U8032 ( .A(n6304), .ZN(n6302) );
  NAND2_X1 U8033 ( .A1(n6302), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6316) );
  INV_X1 U8034 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U8035 ( .A1(n6304), .A2(n6303), .ZN(n6305) );
  NAND2_X1 U8036 ( .A1(n6316), .A2(n6305), .ZN(n8718) );
  OR2_X1 U8037 ( .A1(n8718), .A2(n4398), .ZN(n6311) );
  INV_X1 U8038 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n6308) );
  NAND2_X1 U8039 ( .A1(n8087), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6307) );
  INV_X1 U8040 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8583) );
  OR2_X1 U8041 ( .A1(n6569), .A2(n8583), .ZN(n6306) );
  OAI211_X1 U8042 ( .C1(n4396), .C2(n6308), .A(n6307), .B(n6306), .ZN(n6309)
         );
  INV_X1 U8043 ( .A(n6309), .ZN(n6310) );
  NAND2_X1 U8044 ( .A1(n8728), .A2(n8142), .ZN(n6312) );
  NOR2_X1 U8045 ( .A1(n8192), .A2(n6312), .ZN(n6313) );
  AOI21_X1 U8046 ( .B1(n8192), .B2(n6312), .A(n6313), .ZN(n8320) );
  NAND2_X1 U8047 ( .A1(n8321), .A2(n8320), .ZN(n8190) );
  INV_X1 U8048 ( .A(n6313), .ZN(n6331) );
  NAND2_X1 U8049 ( .A1(n7859), .A2(n6164), .ZN(n6315) );
  XNOR2_X1 U8050 ( .A(n8920), .B(n5984), .ZN(n6326) );
  INV_X1 U8051 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8195) );
  NAND2_X1 U8052 ( .A1(n6316), .A2(n8195), .ZN(n6317) );
  NAND2_X1 U8053 ( .A1(n8698), .A2(n6318), .ZN(n6325) );
  INV_X1 U8054 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6321) );
  NAND2_X1 U8055 ( .A1(n6395), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6320) );
  NAND2_X1 U8056 ( .A1(n5901), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6319) );
  OAI211_X1 U8057 ( .C1(n6322), .C2(n6321), .A(n6320), .B(n6319), .ZN(n6323)
         );
  INV_X1 U8058 ( .A(n6323), .ZN(n6324) );
  NOR2_X1 U8059 ( .A1(n8681), .A2(n6812), .ZN(n6327) );
  NAND2_X1 U8060 ( .A1(n6326), .A2(n6327), .ZN(n6332) );
  INV_X1 U8061 ( .A(n6326), .ZN(n6329) );
  INV_X1 U8062 ( .A(n6327), .ZN(n6328) );
  NAND2_X1 U8063 ( .A1(n6329), .A2(n6328), .ZN(n6330) );
  NAND2_X1 U8064 ( .A1(n6332), .A2(n6330), .ZN(n8191) );
  INV_X1 U8065 ( .A(n6332), .ZN(n6333) );
  INV_X1 U8066 ( .A(n6336), .ZN(n6334) );
  NAND2_X1 U8067 ( .A1(n6334), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8217) );
  INV_X1 U8068 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U8069 ( .A1(n6336), .A2(n6335), .ZN(n6337) );
  NAND2_X1 U8070 ( .A1(n8217), .A2(n6337), .ZN(n6387) );
  INV_X1 U8071 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6340) );
  NAND2_X1 U8072 ( .A1(n6395), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6339) );
  NAND2_X1 U8073 ( .A1(n8087), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6338) );
  OAI211_X1 U8074 ( .C1(n6340), .C2(n6569), .A(n6339), .B(n6338), .ZN(n6341)
         );
  INV_X1 U8075 ( .A(n6341), .ZN(n6342) );
  NOR2_X1 U8076 ( .A1(n8204), .A2(n6812), .ZN(n6344) );
  XNOR2_X1 U8077 ( .A(n6344), .B(n5984), .ZN(n6350) );
  NAND2_X1 U8078 ( .A1(n7911), .A2(n6164), .ZN(n6346) );
  INV_X1 U8079 ( .A(n8685), .ZN(n8689) );
  OR2_X1 U8080 ( .A1(n5908), .A2(n8145), .ZN(n6505) );
  OR2_X1 U8081 ( .A1(n5908), .A2(n8865), .ZN(n6347) );
  NOR3_X1 U8082 ( .A1(n8689), .A2(n6350), .A3(n10213), .ZN(n6348) );
  AOI21_X1 U8083 ( .B1(n6350), .B2(n8689), .A(n6348), .ZN(n6386) );
  NAND3_X1 U8084 ( .A1(n8685), .A2(n10255), .A3(n6350), .ZN(n6349) );
  OAI21_X1 U8085 ( .B1(n8685), .B2(n6350), .A(n6349), .ZN(n6351) );
  NOR2_X1 U8086 ( .A1(n8689), .A2(n10255), .ZN(n8913) );
  OR2_X1 U8087 ( .A1(n6353), .A2(n6352), .ZN(n6354) );
  NAND2_X1 U8088 ( .A1(n6354), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6355) );
  XNOR2_X1 U8089 ( .A(n6355), .B(P2_IR_REG_25__SCAN_IN), .ZN(n6376) );
  INV_X1 U8090 ( .A(n6376), .ZN(n7732) );
  INV_X1 U8091 ( .A(P2_B_REG_SCAN_IN), .ZN(n8639) );
  NAND2_X1 U8092 ( .A1(n6357), .A2(n6356), .ZN(n6358) );
  INV_X1 U8093 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6378) );
  NAND2_X1 U8094 ( .A1(n6381), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6359) );
  XNOR2_X1 U8095 ( .A(n8639), .B(n7592), .ZN(n6360) );
  NAND2_X1 U8096 ( .A1(n7732), .A2(n6360), .ZN(n6364) );
  NAND2_X1 U8097 ( .A1(n4465), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6363) );
  XNOR2_X1 U8098 ( .A(n6363), .B(P2_IR_REG_26__SCAN_IN), .ZN(n7822) );
  INV_X1 U8099 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10188) );
  NOR2_X1 U8100 ( .A1(n7822), .A2(n6376), .ZN(n10189) );
  AOI21_X1 U8101 ( .B1(n10175), .B2(n10188), .A(n10189), .ZN(n6853) );
  NOR4_X1 U8102 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6368) );
  NOR4_X1 U8103 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6367) );
  NOR4_X1 U8104 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n6366) );
  NOR4_X1 U8105 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6365) );
  NAND4_X1 U8106 ( .A1(n6368), .A2(n6367), .A3(n6366), .A4(n6365), .ZN(n6373)
         );
  NOR2_X1 U8107 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .ZN(
        n8430) );
  NOR4_X1 U8108 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n6371) );
  NOR4_X1 U8109 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6370) );
  NOR4_X1 U8110 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6369) );
  NAND4_X1 U8111 ( .A1(n8430), .A2(n6371), .A3(n6370), .A4(n6369), .ZN(n6372)
         );
  OAI21_X1 U8112 ( .B1(n6373), .B2(n6372), .A(n10175), .ZN(n6851) );
  AND2_X1 U8113 ( .A1(n6853), .A2(n6851), .ZN(n6502) );
  NOR2_X1 U8114 ( .A1(n7592), .A2(n7822), .ZN(n10186) );
  INV_X1 U8115 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10185) );
  AND2_X1 U8116 ( .A1(n10175), .A2(n10185), .ZN(n6374) );
  INV_X1 U8117 ( .A(n6919), .ZN(n6375) );
  NAND2_X1 U8118 ( .A1(n6502), .A2(n6375), .ZN(n6382) );
  NAND2_X1 U8119 ( .A1(n6382), .A2(n6850), .ZN(n6388) );
  AND2_X1 U8120 ( .A1(n7822), .A2(n6376), .ZN(n6377) );
  NAND2_X1 U8121 ( .A1(n7592), .A2(n6377), .ZN(n6626) );
  OR2_X1 U8122 ( .A1(n6379), .A2(n6378), .ZN(n6380) );
  NAND2_X1 U8123 ( .A1(n6381), .A2(n6380), .ZN(n6390) );
  INV_X1 U8124 ( .A(n10176), .ZN(n6500) );
  NAND2_X1 U8125 ( .A1(n8913), .A2(n8263), .ZN(n6384) );
  NOR2_X1 U8126 ( .A1(n6382), .A2(n10176), .ZN(n6393) );
  NOR2_X1 U8127 ( .A1(n10213), .A2(n6624), .ZN(n6383) );
  NAND2_X1 U8128 ( .A1(n6384), .A2(n10098), .ZN(n6385) );
  INV_X1 U8129 ( .A(n6387), .ZN(n8686) );
  NAND2_X1 U8130 ( .A1(n8145), .A2(n8865), .ZN(n8178) );
  NAND3_X1 U8131 ( .A1(n6388), .A2(n6626), .A3(n6811), .ZN(n6389) );
  NAND2_X1 U8132 ( .A1(n6389), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6391) );
  OR2_X1 U8133 ( .A1(n6390), .A2(P2_U3152), .ZN(n8182) );
  INV_X1 U8134 ( .A(n10152), .ZN(n8303) );
  INV_X1 U8135 ( .A(n8178), .ZN(n6392) );
  INV_X1 U8136 ( .A(n6394), .ZN(n6401) );
  OR2_X1 U8137 ( .A1(n8217), .A2(n4397), .ZN(n6400) );
  INV_X1 U8138 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8570) );
  NAND2_X1 U8139 ( .A1(n8087), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6397) );
  NAND2_X1 U8140 ( .A1(n6395), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6396) );
  OAI211_X1 U8141 ( .C1(n8570), .C2(n6569), .A(n6397), .B(n6396), .ZN(n6398)
         );
  INV_X1 U8142 ( .A(n6398), .ZN(n6399) );
  INV_X1 U8143 ( .A(n8682), .ZN(n8329) );
  AOI22_X1 U8144 ( .A1(n8686), .A2(n8303), .B1(n10138), .B2(n8329), .ZN(n6403)
         );
  AOI22_X1 U8145 ( .A1(n10140), .A2(n8714), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6402) );
  INV_X1 U8146 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6436) );
  INV_X1 U8147 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9019) );
  INV_X1 U8148 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8607) );
  MUX2_X1 U8149 ( .A(n9019), .B(n8607), .S(n5868), .Z(n6408) );
  INV_X1 U8150 ( .A(SI_29_), .ZN(n6407) );
  NAND2_X1 U8151 ( .A1(n6408), .A2(n6407), .ZN(n6411) );
  INV_X1 U8152 ( .A(n6408), .ZN(n6409) );
  NAND2_X1 U8153 ( .A1(n6409), .A2(SI_29_), .ZN(n6410) );
  AND2_X1 U8154 ( .A1(n6411), .A2(n6410), .ZN(n6426) );
  MUX2_X1 U8155 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n5868), .Z(n6412) );
  NAND2_X1 U8156 ( .A1(n6422), .A2(SI_30_), .ZN(n6416) );
  INV_X1 U8157 ( .A(n6412), .ZN(n6413) );
  MUX2_X1 U8158 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n4391), .Z(n6417) );
  XNOR2_X1 U8159 ( .A(n6417), .B(SI_31_), .ZN(n6418) );
  INV_X1 U8160 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6420) );
  NOR2_X1 U8161 ( .A1(n6428), .A2(n6420), .ZN(n6421) );
  NAND2_X1 U8162 ( .A1(n8234), .A2(n5164), .ZN(n6425) );
  INV_X1 U8163 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9875) );
  OR2_X1 U8164 ( .A1(n6428), .A2(n9875), .ZN(n6424) );
  INV_X1 U8165 ( .A(n9501), .ZN(n6431) );
  NAND2_X1 U8166 ( .A1(n8202), .A2(n5164), .ZN(n6430) );
  OR2_X1 U8167 ( .A1(n6428), .A2(n8607), .ZN(n6429) );
  NAND2_X1 U8168 ( .A1(n6432), .A2(n10003), .ZN(n8189) );
  NAND2_X1 U8169 ( .A1(n5009), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6434) );
  INV_X1 U8170 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8185) );
  OR2_X1 U8171 ( .A1(n4990), .A2(n8185), .ZN(n6433) );
  OAI211_X1 U8172 ( .C1(n5210), .C2(n6436), .A(n6434), .B(n6433), .ZN(n9288)
         );
  INV_X1 U8173 ( .A(n7861), .ZN(n9448) );
  AND2_X1 U8174 ( .A1(n9448), .A2(P1_B_REG_SCAN_IN), .ZN(n6435) );
  NOR2_X1 U8175 ( .A1(n10062), .A2(n6435), .ZN(n6448) );
  NAND2_X1 U8176 ( .A1(n9288), .A2(n6448), .ZN(n9731) );
  MUX2_X1 U8177 ( .A(n6436), .B(n8184), .S(n10083), .Z(n6437) );
  NAND2_X1 U8178 ( .A1(n6437), .A2(n4920), .ZN(P1_U3554) );
  NAND2_X1 U8179 ( .A1(n6438), .A2(n4912), .ZN(n6440) );
  OR2_X1 U8180 ( .A1(n6452), .A2(n6982), .ZN(n9392) );
  NAND2_X1 U8181 ( .A1(n6452), .A2(n6982), .ZN(n9437) );
  NAND2_X1 U8182 ( .A1(n9392), .A2(n9437), .ZN(n9327) );
  XNOR2_X1 U8183 ( .A(n6440), .B(n6439), .ZN(n9506) );
  INV_X1 U8184 ( .A(n9391), .ZN(n6441) );
  XNOR2_X1 U8185 ( .A(n6443), .B(n6439), .ZN(n6444) );
  NAND2_X1 U8186 ( .A1(n6444), .A2(n9637), .ZN(n6450) );
  INV_X1 U8187 ( .A(n9534), .ZN(n9457) );
  INV_X1 U8188 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9734) );
  NAND2_X1 U8189 ( .A1(n5009), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6447) );
  NAND2_X1 U8190 ( .A1(n6445), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6446) );
  OAI211_X1 U8191 ( .C1(n5210), .C2(n9734), .A(n6447), .B(n6446), .ZN(n9456)
         );
  AOI22_X1 U8192 ( .A1(n9457), .A2(n9819), .B1(n6448), .B2(n9456), .ZN(n6449)
         );
  NAND2_X1 U8193 ( .A1(n6450), .A2(n6449), .ZN(n9512) );
  AOI211_X1 U8194 ( .C1(n6452), .C2(n6451), .A(n9695), .B(n9499), .ZN(n9507)
         );
  OAI21_X1 U8195 ( .B1(n6482), .B2(n10081), .A(n6455), .ZN(P1_U3552) );
  INV_X1 U8196 ( .A(n6479), .ZN(n6469) );
  NAND2_X1 U8197 ( .A1(n6464), .A2(n6456), .ZN(n6459) );
  OR2_X1 U8198 ( .A1(n9534), .A2(n6457), .ZN(n6458) );
  NAND2_X1 U8199 ( .A1(n6459), .A2(n6458), .ZN(n6461) );
  XNOR2_X1 U8200 ( .A(n6461), .B(n6460), .ZN(n6466) );
  AOI22_X1 U8201 ( .A1(n6464), .A2(n6463), .B1(n6462), .B2(n9457), .ZN(n6465)
         );
  XNOR2_X1 U8202 ( .A(n6466), .B(n6465), .ZN(n6471) );
  INV_X1 U8203 ( .A(n6471), .ZN(n6468) );
  INV_X1 U8204 ( .A(n6470), .ZN(n6467) );
  AND2_X1 U8205 ( .A1(n6471), .A2(n9160), .ZN(n6478) );
  NAND3_X1 U8206 ( .A1(n6471), .A2(n9160), .A3(n6470), .ZN(n6476) );
  AOI22_X1 U8207 ( .A1(n9517), .A2(n9092), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6472) );
  OAI21_X1 U8208 ( .B1(n6982), .B2(n9162), .A(n6472), .ZN(n6474) );
  NOR2_X1 U8209 ( .A1(n5486), .A2(n9170), .ZN(n6473) );
  AOI211_X1 U8210 ( .C1(n9167), .C2(n9458), .A(n6474), .B(n6473), .ZN(n6475)
         );
  NAND2_X1 U8211 ( .A1(n6481), .A2(n6480), .ZN(P1_U3218) );
  INV_X1 U8212 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U8213 ( .A1(n10075), .A2(n6483), .ZN(n6484) );
  INV_X1 U8214 ( .A(n9864), .ZN(n6485) );
  NAND2_X1 U8215 ( .A1(n6452), .A2(n6485), .ZN(n6486) );
  NAND2_X1 U8216 ( .A1(n6487), .A2(n6486), .ZN(P1_U3520) );
  INV_X1 U8217 ( .A(n10190), .ZN(n6488) );
  INV_X2 U8218 ( .A(n8338), .ZN(P2_U3966) );
  INV_X1 U8219 ( .A(n6489), .ZN(n7499) );
  INV_X1 U8220 ( .A(n10191), .ZN(n7109) );
  INV_X1 U8221 ( .A(n6491), .ZN(n6490) );
  INV_X1 U8222 ( .A(n7988), .ZN(n6496) );
  INV_X1 U8223 ( .A(n7110), .ZN(n6493) );
  NAND2_X1 U8224 ( .A1(n6511), .A2(n6493), .ZN(n6495) );
  NAND2_X1 U8225 ( .A1(n8170), .A2(n8171), .ZN(n8141) );
  OAI211_X1 U8226 ( .C1(n6906), .C2(n6496), .A(n6495), .B(n10156), .ZN(n6499)
         );
  AOI22_X1 U8227 ( .A1(n8877), .A2(n6497), .B1(n10111), .B2(n8879), .ZN(n6498)
         );
  NAND2_X1 U8228 ( .A1(n6499), .A2(n6498), .ZN(n6857) );
  NAND3_X1 U8229 ( .A1(n6500), .A2(n6919), .A3(n6811), .ZN(n6854) );
  INV_X1 U8230 ( .A(n6854), .ZN(n6501) );
  NAND2_X1 U8231 ( .A1(n6502), .A2(n6501), .ZN(n6503) );
  MUX2_X1 U8232 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6857), .S(n8881), .Z(n6514)
         );
  OR2_X1 U8233 ( .A1(n6503), .A2(n8734), .ZN(n7144) );
  OAI21_X1 U8234 ( .B1(n7109), .B2(n6894), .A(n7036), .ZN(n6856) );
  OAI22_X1 U8235 ( .A1(n8780), .A2(n6856), .B1(n6681), .B2(n8888), .ZN(n6513)
         );
  INV_X1 U8236 ( .A(n6505), .ZN(n6506) );
  NAND2_X1 U8237 ( .A1(n6508), .A2(n7956), .ZN(n6507) );
  NAND3_X1 U8238 ( .A1(n6558), .A2(n6507), .A3(n8865), .ZN(n7568) );
  OR2_X1 U8239 ( .A1(n6508), .A2(n8865), .ZN(n7142) );
  NAND2_X1 U8240 ( .A1(n7568), .A2(n7142), .ZN(n6509) );
  NAND2_X1 U8241 ( .A1(n6510), .A2(n6896), .ZN(n6895) );
  OAI21_X1 U8242 ( .B1(n6511), .B2(n6896), .A(n6895), .ZN(n6855) );
  OAI22_X1 U8243 ( .A1(n6894), .A2(n8869), .B1(n8874), .B2(n6855), .ZN(n6512)
         );
  OR3_X1 U8244 ( .A1(n6514), .A2(n6513), .A3(n6512), .ZN(P2_U3295) );
  INV_X1 U8245 ( .A(n6515), .ZN(n6520) );
  AOI21_X1 U8246 ( .B1(n6516), .B2(n6517), .A(n6518), .ZN(n6519) );
  AOI211_X1 U8247 ( .C1(n6520), .C2(n6516), .A(n9144), .B(n6519), .ZN(n6526)
         );
  NOR2_X1 U8248 ( .A1(n9592), .A2(n9170), .ZN(n6525) );
  OAI22_X1 U8249 ( .A1(n9603), .A2(n9139), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6521), .ZN(n6524) );
  OAI22_X1 U8250 ( .A1(n6522), .A2(n9162), .B1(n9164), .B2(n9594), .ZN(n6523)
         );
  OR4_X1 U8251 ( .A1(n6526), .A2(n6525), .A3(n6524), .A4(n6523), .ZN(P1_U3214)
         );
  AND2_X1 U8252 ( .A1(P1_STATE_REG_SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6614) );
  AOI21_X1 U8253 ( .B1(n6527), .B2(P1_U3084), .A(n6614), .ZN(n6528) );
  INV_X1 U8254 ( .A(n6528), .ZN(P1_U3353) );
  NOR2_X1 U8255 ( .A1(n5868), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9871) );
  INV_X2 U8256 ( .A(n9871), .ZN(n9874) );
  AND2_X1 U8257 ( .A1(n5868), .A2(P1_U3084), .ZN(n7907) );
  INV_X2 U8258 ( .A(n7907), .ZN(n9878) );
  OAI222_X1 U8259 ( .A1(n9874), .A2(n6529), .B1(n9878), .B2(n6541), .C1(
        P1_U3084), .C2(n6957), .ZN(P1_U3351) );
  OAI222_X1 U8260 ( .A1(n9874), .A2(n6530), .B1(n9878), .B2(n6539), .C1(
        P1_U3084), .C2(n6597), .ZN(P1_U3349) );
  OAI222_X1 U8261 ( .A1(n9874), .A2(n6531), .B1(n9878), .B2(n6536), .C1(
        P1_U3084), .C2(n6592), .ZN(P1_U3352) );
  OAI222_X1 U8262 ( .A1(n9874), .A2(n6532), .B1(n9878), .B2(n6549), .C1(
        P1_U3084), .C2(n6789), .ZN(P1_U3350) );
  OAI222_X1 U8263 ( .A1(n9874), .A2(n6533), .B1(n9878), .B2(n6547), .C1(
        P1_U3084), .C2(n6589), .ZN(P1_U3348) );
  OAI222_X1 U8264 ( .A1(n9874), .A2(n6534), .B1(n9878), .B2(n6545), .C1(
        P1_U3084), .C2(n6802), .ZN(P1_U3347) );
  OAI222_X1 U8265 ( .A1(n9874), .A2(n6535), .B1(n9878), .B2(n6543), .C1(
        P1_U3084), .C2(n6772), .ZN(P1_U3346) );
  NOR2_X1 U8266 ( .A1(n5868), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9016) );
  OAI222_X1 U8267 ( .A1(n9018), .A2(n6537), .B1(n9021), .B2(n6536), .C1(n6692), 
        .C2(P2_U3152), .ZN(P2_U3357) );
  OAI222_X1 U8268 ( .A1(n6705), .A2(P2_U3152), .B1(n9021), .B2(n6539), .C1(
        n6538), .C2(n9018), .ZN(P2_U3354) );
  OAI222_X1 U8269 ( .A1(n6717), .A2(P2_U3152), .B1(n9021), .B2(n6541), .C1(
        n6540), .C2(n9018), .ZN(P2_U3356) );
  INV_X1 U8270 ( .A(n6748), .ZN(n6755) );
  INV_X1 U8271 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6542) );
  OAI222_X1 U8272 ( .A1(n6755), .A2(P2_U3152), .B1(n9021), .B2(n6543), .C1(
        n6542), .C2(n9018), .ZN(P2_U3351) );
  INV_X1 U8273 ( .A(n6676), .ZN(n6729) );
  OAI222_X1 U8274 ( .A1(n6729), .A2(P2_U3152), .B1(n9021), .B2(n6545), .C1(
        n6544), .C2(n9018), .ZN(P2_U3352) );
  INV_X1 U8275 ( .A(n6669), .ZN(n6675) );
  OAI222_X1 U8276 ( .A1(n6675), .A2(P2_U3152), .B1(n9021), .B2(n6547), .C1(
        n6546), .C2(n9018), .ZN(P2_U3353) );
  OAI222_X1 U8277 ( .A1(n6666), .A2(P2_U3152), .B1(n9021), .B2(n6549), .C1(
        n6548), .C2(n9018), .ZN(P2_U3355) );
  INV_X1 U8278 ( .A(n6550), .ZN(n6552) );
  INV_X1 U8279 ( .A(n9946), .ZN(n6770) );
  OAI222_X1 U8280 ( .A1(n9874), .A2(n6551), .B1(n9878), .B2(n6552), .C1(
        P1_U3084), .C2(n6770), .ZN(P1_U3345) );
  OAI222_X1 U8281 ( .A1(n6935), .A2(P2_U3152), .B1(n9021), .B2(n6552), .C1(
        n8529), .C2(n9018), .ZN(P2_U3350) );
  INV_X1 U8282 ( .A(n6984), .ZN(n6991) );
  INV_X1 U8283 ( .A(n6553), .ZN(n6554) );
  OAI222_X1 U8284 ( .A1(P2_U3152), .A2(n6991), .B1(n9021), .B2(n6554), .C1(
        n8604), .C2(n9018), .ZN(P2_U3349) );
  OAI222_X1 U8285 ( .A1(n9874), .A2(n6555), .B1(n6863), .B2(P1_U3084), .C1(
        n9878), .C2(n6554), .ZN(P1_U3344) );
  NAND2_X1 U8286 ( .A1(n10176), .A2(n8182), .ZN(n6557) );
  NAND2_X1 U8287 ( .A1(n6557), .A2(n6556), .ZN(n6560) );
  OR2_X1 U8288 ( .A1(n10176), .A2(n6558), .ZN(n6559) );
  AND2_X1 U8289 ( .A1(n6560), .A2(n6559), .ZN(n8389) );
  NOR2_X1 U8290 ( .A1(n8350), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8291 ( .A(n7071), .ZN(n6997) );
  INV_X1 U8292 ( .A(n5130), .ZN(n6564) );
  OAI222_X1 U8293 ( .A1(P2_U3152), .A2(n6997), .B1(n9021), .B2(n6564), .C1(
        n6561), .C2(n9018), .ZN(P2_U3348) );
  INV_X1 U8294 ( .A(n6562), .ZN(n6567) );
  INV_X1 U8295 ( .A(n9958), .ZN(n7211) );
  INV_X1 U8296 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6563) );
  OAI222_X1 U8297 ( .A1(n9878), .A2(n6567), .B1(n7211), .B2(P1_U3084), .C1(
        n6563), .C2(n9874), .ZN(P1_U3342) );
  INV_X1 U8298 ( .A(n7220), .ZN(n6870) );
  OAI222_X1 U8299 ( .A1(n9874), .A2(n6565), .B1(n6870), .B2(P1_U3084), .C1(
        n9878), .C2(n6564), .ZN(P1_U3343) );
  INV_X1 U8300 ( .A(n7253), .ZN(n7077) );
  INV_X1 U8301 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6566) );
  OAI222_X1 U8302 ( .A1(P2_U3152), .A2(n7077), .B1(n9021), .B2(n6567), .C1(
        n6566), .C2(n9018), .ZN(P2_U3347) );
  INV_X1 U8303 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U8304 ( .A1(n8087), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6571) );
  INV_X1 U8305 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6568) );
  OR2_X1 U8306 ( .A1(n6569), .A2(n6568), .ZN(n6570) );
  OAI211_X1 U8307 ( .C1(n4396), .C2(n8394), .A(n6571), .B(n6570), .ZN(n8392)
         );
  NAND2_X1 U8308 ( .A1(n8392), .A2(P2_U3966), .ZN(n6572) );
  OAI21_X1 U8309 ( .B1(P2_U3966), .B2(n6420), .A(n6572), .ZN(P2_U3583) );
  INV_X1 U8310 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6574) );
  NAND2_X1 U8311 ( .A1(n9288), .A2(P1_U4006), .ZN(n6573) );
  OAI21_X1 U8312 ( .B1(P1_U4006), .B2(n6574), .A(n6573), .ZN(P1_U3586) );
  OR2_X1 U8313 ( .A1(n9332), .A2(n7499), .ZN(n6575) );
  NAND2_X1 U8314 ( .A1(n6575), .A2(n6968), .ZN(n6587) );
  OR2_X1 U8315 ( .A1(n6587), .A2(n6576), .ZN(n6613) );
  NAND2_X1 U8316 ( .A1(n6613), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8317 ( .A(P1_U3083), .ZN(n6577) );
  NAND2_X1 U8318 ( .A1(n6577), .A2(n6968), .ZN(n9984) );
  INV_X1 U8319 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6607) );
  OR2_X1 U8320 ( .A1(n5478), .A2(P1_U3084), .ZN(n7908) );
  NOR2_X1 U8321 ( .A1(n6587), .A2(n7908), .ZN(n6600) );
  INV_X1 U8322 ( .A(n6600), .ZN(n6578) );
  NOR2_X1 U8323 ( .A1(n6578), .A2(n7861), .ZN(n9966) );
  NOR2_X1 U8324 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6774), .ZN(n6579) );
  AOI21_X1 U8325 ( .B1(n6774), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6579), .ZN(
        n6584) );
  INV_X1 U8326 ( .A(n6597), .ZN(n9928) );
  INV_X1 U8327 ( .A(n6789), .ZN(n6596) );
  INV_X1 U8328 ( .A(n6957), .ZN(n6594) );
  INV_X1 U8329 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6580) );
  MUX2_X1 U8330 ( .A(n6580), .B(P1_REG2_REG_1__SCAN_IN), .S(n6592), .Z(n6731)
         );
  AND2_X1 U8331 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6967) );
  NAND2_X1 U8332 ( .A1(n6731), .A2(n6967), .ZN(n6730) );
  OAI21_X1 U8333 ( .B1(n6592), .B2(n6580), .A(n6730), .ZN(n6960) );
  INV_X1 U8334 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6581) );
  MUX2_X1 U8335 ( .A(n6581), .B(P1_REG2_REG_2__SCAN_IN), .S(n6957), .Z(n6961)
         );
  NAND2_X1 U8336 ( .A1(n6960), .A2(n6961), .ZN(n6959) );
  INV_X1 U8337 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7319) );
  XNOR2_X1 U8338 ( .A(n6789), .B(n7319), .ZN(n6791) );
  MUX2_X1 U8339 ( .A(n6582), .B(P1_REG2_REG_4__SCAN_IN), .S(n6597), .Z(n9922)
         );
  NAND2_X1 U8340 ( .A1(n9923), .A2(n9922), .ZN(n9921) );
  OAI21_X1 U8341 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n9928), .A(n9921), .ZN(
        n6583) );
  NAND2_X1 U8342 ( .A1(n6583), .A2(n6584), .ZN(n6773) );
  OAI21_X1 U8343 ( .B1(n6584), .B2(n6583), .A(n6773), .ZN(n6605) );
  NOR2_X1 U8344 ( .A1(n7861), .A2(P1_U3084), .ZN(n6585) );
  NAND2_X1 U8345 ( .A1(n6585), .A2(n5478), .ZN(n6586) );
  NAND2_X1 U8346 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3084), .ZN(n6588) );
  OAI21_X1 U8347 ( .B1(n9491), .B2(n6589), .A(n6588), .ZN(n6604) );
  INV_X1 U8348 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6590) );
  MUX2_X1 U8349 ( .A(n6590), .B(P1_REG1_REG_2__SCAN_IN), .S(n6957), .Z(n6956)
         );
  INV_X1 U8350 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10077) );
  MUX2_X1 U8351 ( .A(n10077), .B(P1_REG1_REG_1__SCAN_IN), .S(n6592), .Z(n6735)
         );
  AND2_X1 U8352 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6591) );
  NAND2_X1 U8353 ( .A1(n6735), .A2(n6591), .ZN(n6736) );
  INV_X1 U8354 ( .A(n6592), .ZN(n6732) );
  NAND2_X1 U8355 ( .A1(n6732), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6593) );
  NAND2_X1 U8356 ( .A1(n6736), .A2(n6593), .ZN(n6955) );
  NAND2_X1 U8357 ( .A1(n6956), .A2(n6955), .ZN(n6954) );
  NAND2_X1 U8358 ( .A1(n6594), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U8359 ( .A1(n6954), .A2(n6595), .ZN(n6785) );
  XNOR2_X1 U8360 ( .A(n6789), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n6784) );
  AND2_X1 U8361 ( .A1(n6785), .A2(n6784), .ZN(n6787) );
  AOI21_X1 U8362 ( .B1(n6596), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6787), .ZN(
        n9920) );
  MUX2_X1 U8363 ( .A(n6598), .B(P1_REG1_REG_4__SCAN_IN), .S(n6597), .Z(n9919)
         );
  NAND2_X1 U8364 ( .A1(n9920), .A2(n9919), .ZN(n9918) );
  OAI21_X1 U8365 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9928), .A(n9918), .ZN(
        n6602) );
  NAND2_X1 U8366 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6774), .ZN(n6599) );
  OAI21_X1 U8367 ( .B1(n6774), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6599), .ZN(
        n6601) );
  NOR2_X1 U8368 ( .A1(n6602), .A2(n6601), .ZN(n6763) );
  NAND2_X1 U8369 ( .A1(n6600), .A2(n7861), .ZN(n9492) );
  AOI211_X1 U8370 ( .C1(n6602), .C2(n6601), .A(n6763), .B(n9492), .ZN(n6603)
         );
  AOI211_X1 U8371 ( .C1(n9966), .C2(n6605), .A(n6604), .B(n6603), .ZN(n6606)
         );
  OAI21_X1 U8372 ( .B1(n9984), .B2(n6607), .A(n6606), .ZN(P1_U3246) );
  NAND2_X1 U8373 ( .A1(n5593), .A2(P1_U4006), .ZN(n6608) );
  OAI21_X1 U8374 ( .B1(P1_U4006), .B2(n5925), .A(n6608), .ZN(P1_U3555) );
  INV_X1 U8375 ( .A(n6113), .ZN(n6610) );
  INV_X1 U8376 ( .A(n9976), .ZN(n7210) );
  OAI222_X1 U8377 ( .A1(n9874), .A2(n6609), .B1(n9878), .B2(n6610), .C1(
        P1_U3084), .C2(n7210), .ZN(P1_U3341) );
  INV_X1 U8378 ( .A(n7433), .ZN(n7263) );
  OAI222_X1 U8379 ( .A1(n9018), .A2(n6611), .B1(n9021), .B2(n6610), .C1(n7263), 
        .C2(P2_U3152), .ZN(P2_U3346) );
  INV_X1 U8380 ( .A(n9984), .ZN(n9997) );
  INV_X1 U8381 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n8619) );
  NAND3_X1 U8382 ( .A1(n9998), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6612), .ZN(
        n6621) );
  OAI22_X1 U8383 ( .A1(n7861), .A2(n6967), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n6612), .ZN(n6619) );
  INV_X1 U8384 ( .A(n6613), .ZN(n6618) );
  INV_X1 U8385 ( .A(n7908), .ZN(n6616) );
  INV_X1 U8386 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10039) );
  NAND2_X1 U8387 ( .A1(n9448), .A2(n10039), .ZN(n6615) );
  AOI21_X1 U8388 ( .B1(n6616), .B2(n6615), .A(n6614), .ZN(n6969) );
  INV_X1 U8389 ( .A(n6969), .ZN(n6617) );
  OAI211_X1 U8390 ( .C1(n5478), .C2(n6619), .A(n6618), .B(n6617), .ZN(n6620)
         );
  OAI211_X1 U8391 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n8619), .A(n6621), .B(n6620), .ZN(n6622) );
  AOI21_X1 U8392 ( .B1(n9997), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n6622), .ZN(
        n6623) );
  INV_X1 U8393 ( .A(n6623), .ZN(P1_U3241) );
  OR2_X1 U8394 ( .A1(n6394), .A2(P2_U3152), .ZN(n7912) );
  OR2_X1 U8395 ( .A1(n10176), .A2(n6624), .ZN(n6625) );
  OAI211_X1 U8396 ( .C1(n6626), .C2(n7912), .A(n6625), .B(n8182), .ZN(n6635)
         );
  NAND2_X1 U8397 ( .A1(n6635), .A2(n5944), .ZN(n6627) );
  NAND2_X1 U8398 ( .A1(n6627), .A2(n8338), .ZN(n6641) );
  NAND2_X1 U8399 ( .A1(n6641), .A2(n6394), .ZN(n8376) );
  INV_X1 U8400 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6628) );
  NOR2_X1 U8401 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6628), .ZN(n6639) );
  INV_X1 U8402 ( .A(n6705), .ZN(n6648) );
  INV_X1 U8403 ( .A(n6666), .ZN(n6632) );
  INV_X1 U8404 ( .A(n6717), .ZN(n6644) );
  INV_X1 U8405 ( .A(n6692), .ZN(n6630) );
  INV_X1 U8406 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6629) );
  NAND2_X1 U8407 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n6684) );
  NOR2_X1 U8408 ( .A1(n6683), .A2(n6684), .ZN(n6682) );
  AOI21_X1 U8409 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(n6630), .A(n6682), .ZN(
        n6709) );
  INV_X1 U8410 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6631) );
  MUX2_X1 U8411 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6631), .S(n6717), .Z(n6708)
         );
  XOR2_X1 U8412 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6666), .Z(n6656) );
  MUX2_X1 U8413 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6633), .S(n6705), .Z(n6694)
         );
  NOR2_X1 U8414 ( .A1(n6695), .A2(n6694), .ZN(n6693) );
  AOI21_X1 U8415 ( .B1(n6648), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6693), .ZN(
        n6637) );
  XNOR2_X1 U8416 ( .A(n6669), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n6636) );
  AND2_X1 U8417 ( .A1(n5944), .A2(n8223), .ZN(n6634) );
  NAND2_X1 U8418 ( .A1(n6635), .A2(n6634), .ZN(n8377) );
  NOR2_X1 U8419 ( .A1(n6637), .A2(n6636), .ZN(n6668) );
  AOI211_X1 U8420 ( .C1(n6637), .C2(n6636), .A(n8377), .B(n6668), .ZN(n6638)
         );
  AOI211_X1 U8421 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n8350), .A(n6639), .B(
        n6638), .ZN(n6654) );
  NOR2_X1 U8422 ( .A1(n6394), .A2(n8223), .ZN(n6640) );
  MUX2_X1 U8423 ( .A(n6642), .B(P2_REG2_REG_1__SCAN_IN), .S(n6692), .Z(n6688)
         );
  NAND3_X1 U8424 ( .A1(n6688), .A2(P2_REG2_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n6687) );
  OAI21_X1 U8425 ( .B1(n6642), .B2(n6692), .A(n6687), .ZN(n6713) );
  MUX2_X1 U8426 ( .A(n6643), .B(P2_REG2_REG_2__SCAN_IN), .S(n6717), .Z(n6714)
         );
  NAND2_X1 U8427 ( .A1(n6713), .A2(n6714), .ZN(n6712) );
  NAND2_X1 U8428 ( .A1(n6644), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6662) );
  MUX2_X1 U8429 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6645), .S(n6666), .Z(n6661)
         );
  AOI21_X1 U8430 ( .B1(n6712), .B2(n6662), .A(n6661), .ZN(n6660) );
  NOR2_X1 U8431 ( .A1(n6666), .A2(n6645), .ZN(n6697) );
  INV_X1 U8432 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6646) );
  MUX2_X1 U8433 ( .A(n6646), .B(P2_REG2_REG_4__SCAN_IN), .S(n6705), .Z(n6647)
         );
  OAI21_X1 U8434 ( .B1(n6660), .B2(n6697), .A(n6647), .ZN(n6702) );
  NAND2_X1 U8435 ( .A1(n6648), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6650) );
  INV_X1 U8436 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n8470) );
  MUX2_X1 U8437 ( .A(n8470), .B(P2_REG2_REG_5__SCAN_IN), .S(n6669), .Z(n6649)
         );
  AOI21_X1 U8438 ( .B1(n6702), .B2(n6650), .A(n6649), .ZN(n6724) );
  INV_X1 U8439 ( .A(n6724), .ZN(n6652) );
  NAND3_X1 U8440 ( .A1(n6702), .A2(n6650), .A3(n6649), .ZN(n6651) );
  NAND3_X1 U8441 ( .A1(n8382), .A2(n6652), .A3(n6651), .ZN(n6653) );
  OAI211_X1 U8442 ( .C1(n8376), .C2(n6675), .A(n6654), .B(n6653), .ZN(P2_U3250) );
  NOR2_X1 U8443 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5966), .ZN(n6659) );
  AOI211_X1 U8444 ( .C1(n6657), .C2(n6656), .A(n6655), .B(n8377), .ZN(n6658)
         );
  AOI211_X1 U8445 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n8350), .A(n6659), .B(
        n6658), .ZN(n6665) );
  INV_X1 U8446 ( .A(n6660), .ZN(n6700) );
  NAND3_X1 U8447 ( .A1(n6712), .A2(n6662), .A3(n6661), .ZN(n6663) );
  NAND3_X1 U8448 ( .A1(n8382), .A2(n6700), .A3(n6663), .ZN(n6664) );
  OAI211_X1 U8449 ( .C1(n8376), .C2(n6666), .A(n6665), .B(n6664), .ZN(P2_U3248) );
  INV_X1 U8450 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6667) );
  NOR2_X1 U8451 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6667), .ZN(n6674) );
  AOI21_X1 U8452 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n6669), .A(n6668), .ZN(
        n6720) );
  XNOR2_X1 U8453 ( .A(n6676), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n6719) );
  NOR2_X1 U8454 ( .A1(n6720), .A2(n6719), .ZN(n6718) );
  AOI21_X1 U8455 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n6676), .A(n6718), .ZN(
        n6672) );
  INV_X1 U8456 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6670) );
  MUX2_X1 U8457 ( .A(n6670), .B(P2_REG1_REG_7__SCAN_IN), .S(n6748), .Z(n6671)
         );
  AOI211_X1 U8458 ( .C1(n6672), .C2(n6671), .A(n8377), .B(n6747), .ZN(n6673)
         );
  AOI211_X1 U8459 ( .C1(P2_ADDR_REG_7__SCAN_IN), .C2(n8350), .A(n6674), .B(
        n6673), .ZN(n6680) );
  NOR2_X1 U8460 ( .A1(n6675), .A2(n8470), .ZN(n6723) );
  MUX2_X1 U8461 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n8882), .S(n6676), .Z(n6722)
         );
  OAI21_X1 U8462 ( .B1(n6724), .B2(n6723), .A(n6722), .ZN(n6726) );
  OAI21_X1 U8463 ( .B1(n8882), .B2(n6729), .A(n6726), .ZN(n6678) );
  MUX2_X1 U8464 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7094), .S(n6748), .Z(n6677)
         );
  NAND2_X1 U8465 ( .A1(n6677), .A2(n6678), .ZN(n6754) );
  OAI211_X1 U8466 ( .C1(n6678), .C2(n6677), .A(n8382), .B(n6754), .ZN(n6679)
         );
  OAI211_X1 U8467 ( .C1(n8376), .C2(n6755), .A(n6680), .B(n6679), .ZN(P2_U3252) );
  NOR2_X1 U8468 ( .A1(n6681), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6686) );
  AOI211_X1 U8469 ( .C1(n6684), .C2(n6683), .A(n6682), .B(n8377), .ZN(n6685)
         );
  AOI211_X1 U8470 ( .C1(P2_ADDR_REG_1__SCAN_IN), .C2(n8350), .A(n6686), .B(
        n6685), .ZN(n6691) );
  AND2_X1 U8471 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n6689) );
  OAI211_X1 U8472 ( .C1(n6689), .C2(n6688), .A(n8382), .B(n6687), .ZN(n6690)
         );
  OAI211_X1 U8473 ( .C1(n8376), .C2(n6692), .A(n6691), .B(n6690), .ZN(P2_U3246) );
  AND2_X1 U8474 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n8281) );
  AOI211_X1 U8475 ( .C1(n6695), .C2(n6694), .A(n8377), .B(n6693), .ZN(n6696)
         );
  AOI211_X1 U8476 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n8350), .A(n8281), .B(
        n6696), .ZN(n6704) );
  INV_X1 U8477 ( .A(n6697), .ZN(n6699) );
  MUX2_X1 U8478 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6646), .S(n6705), .Z(n6698)
         );
  NAND3_X1 U8479 ( .A1(n6700), .A2(n6699), .A3(n6698), .ZN(n6701) );
  NAND3_X1 U8480 ( .A1(n8382), .A2(n6702), .A3(n6701), .ZN(n6703) );
  OAI211_X1 U8481 ( .C1(n8376), .C2(n6705), .A(n6704), .B(n6703), .ZN(P2_U3249) );
  NOR2_X1 U8482 ( .A1(n6706), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6711) );
  AOI211_X1 U8483 ( .C1(n6709), .C2(n6708), .A(n6707), .B(n8377), .ZN(n6710)
         );
  AOI211_X1 U8484 ( .C1(P2_ADDR_REG_2__SCAN_IN), .C2(n8350), .A(n6711), .B(
        n6710), .ZN(n6716) );
  OAI211_X1 U8485 ( .C1(n6714), .C2(n6713), .A(n8382), .B(n6712), .ZN(n6715)
         );
  OAI211_X1 U8486 ( .C1(n8376), .C2(n6717), .A(n6716), .B(n6715), .ZN(P2_U3247) );
  AND2_X1 U8487 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8310) );
  AOI211_X1 U8488 ( .C1(n6720), .C2(n6719), .A(n8377), .B(n6718), .ZN(n6721)
         );
  AOI211_X1 U8489 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n8350), .A(n8310), .B(
        n6721), .ZN(n6728) );
  OR3_X1 U8490 ( .A1(n6724), .A2(n6723), .A3(n6722), .ZN(n6725) );
  NAND3_X1 U8491 ( .A1(n8382), .A2(n6726), .A3(n6725), .ZN(n6727) );
  OAI211_X1 U8492 ( .C1(n8376), .C2(n6729), .A(n6728), .B(n6727), .ZN(P2_U3251) );
  OAI211_X1 U8493 ( .C1(n6731), .C2(n6967), .A(n9966), .B(n6730), .ZN(n6734)
         );
  INV_X1 U8494 ( .A(n9491), .ZN(n9992) );
  NAND2_X1 U8495 ( .A1(n9992), .A2(n6732), .ZN(n6733) );
  OAI211_X1 U8496 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n7206), .A(n6734), .B(n6733), .ZN(n6741) );
  NAND2_X1 U8497 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n6739) );
  INV_X1 U8498 ( .A(n6735), .ZN(n6738) );
  INV_X1 U8499 ( .A(n6736), .ZN(n6737) );
  AOI211_X1 U8500 ( .C1(n6739), .C2(n6738), .A(n6737), .B(n9492), .ZN(n6740)
         );
  AOI211_X1 U8501 ( .C1(P1_ADDR_REG_1__SCAN_IN), .C2(n9997), .A(n6741), .B(
        n6740), .ZN(n6742) );
  INV_X1 U8502 ( .A(n6742), .ZN(P1_U3242) );
  INV_X1 U8503 ( .A(n6743), .ZN(n6746) );
  AOI22_X1 U8504 ( .A1(n7544), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9871), .ZN(n6744) );
  OAI21_X1 U8505 ( .B1(n6746), .B2(n9878), .A(n6744), .ZN(P1_U3340) );
  INV_X1 U8506 ( .A(n7512), .ZN(n7506) );
  OAI222_X1 U8507 ( .A1(P2_U3152), .A2(n7506), .B1(n9021), .B2(n6746), .C1(
        n6745), .C2(n9018), .ZN(P2_U3345) );
  NAND2_X1 U8508 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n10127) );
  INV_X1 U8509 ( .A(n10127), .ZN(n6753) );
  INV_X1 U8510 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6749) );
  MUX2_X1 U8511 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6749), .S(n6935), .Z(n6750)
         );
  AOI211_X1 U8512 ( .C1(n6751), .C2(n6750), .A(n6927), .B(n8377), .ZN(n6752)
         );
  AOI211_X1 U8513 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n8350), .A(n6753), .B(
        n6752), .ZN(n6759) );
  OAI21_X1 U8514 ( .B1(n6755), .B2(n7094), .A(n6754), .ZN(n6757) );
  MUX2_X1 U8515 ( .A(n7180), .B(P2_REG2_REG_8__SCAN_IN), .S(n6935), .Z(n6756)
         );
  NAND2_X1 U8516 ( .A1(n6756), .A2(n6757), .ZN(n6934) );
  OAI211_X1 U8517 ( .C1(n6757), .C2(n6756), .A(n8382), .B(n6934), .ZN(n6758)
         );
  OAI211_X1 U8518 ( .C1(n8376), .C2(n6935), .A(n6759), .B(n6758), .ZN(P2_U3253) );
  INV_X1 U8519 ( .A(n6760), .ZN(n6762) );
  INV_X1 U8520 ( .A(n7653), .ZN(n7645) );
  OAI222_X1 U8521 ( .A1(n9878), .A2(n6762), .B1(n7645), .B2(P1_U3084), .C1(
        n8436), .C2(n9874), .ZN(P1_U3339) );
  INV_X1 U8522 ( .A(n7829), .ZN(n7509) );
  OAI222_X1 U8523 ( .A1(P2_U3152), .A2(n7509), .B1(n9021), .B2(n6762), .C1(
        n6761), .C2(n9018), .ZN(P2_U3344) );
  AOI22_X1 U8524 ( .A1(n9946), .A2(P1_REG1_REG_8__SCAN_IN), .B1(n5084), .B2(
        n6770), .ZN(n9952) );
  AOI22_X1 U8525 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n9933), .B1(n6772), .B2(
        n5063), .ZN(n9936) );
  AOI21_X1 U8526 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n6774), .A(n6763), .ZN(
        n6800) );
  NOR2_X1 U8527 ( .A1(n6776), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6764) );
  AOI21_X1 U8528 ( .B1(n6776), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6764), .ZN(
        n6799) );
  NAND2_X1 U8529 ( .A1(n6800), .A2(n6799), .ZN(n6798) );
  OAI21_X1 U8530 ( .B1(n6776), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6798), .ZN(
        n9935) );
  NAND2_X1 U8531 ( .A1(n9936), .A2(n9935), .ZN(n9934) );
  OAI21_X1 U8532 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n9933), .A(n9934), .ZN(
        n9951) );
  NAND2_X1 U8533 ( .A1(n9952), .A2(n9951), .ZN(n9950) );
  OAI21_X1 U8534 ( .B1(n9946), .B2(P1_REG1_REG_8__SCAN_IN), .A(n9950), .ZN(
        n6766) );
  MUX2_X1 U8535 ( .A(n6862), .B(P1_REG1_REG_9__SCAN_IN), .S(n6863), .Z(n6765)
         );
  NAND2_X1 U8536 ( .A1(n6765), .A2(n6766), .ZN(n6864) );
  OAI21_X1 U8537 ( .B1(n6766), .B2(n6765), .A(n6864), .ZN(n6782) );
  NAND2_X1 U8538 ( .A1(n9997), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n6769) );
  NOR2_X1 U8539 ( .A1(n6767), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7622) );
  INV_X1 U8540 ( .A(n7622), .ZN(n6768) );
  OAI211_X1 U8541 ( .C1(n9491), .C2(n6863), .A(n6769), .B(n6768), .ZN(n6781)
         );
  AOI22_X1 U8542 ( .A1(n9946), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n5085), .B2(
        n6770), .ZN(n9949) );
  INV_X1 U8543 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6771) );
  AOI22_X1 U8544 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n9933), .B1(n6772), .B2(
        n6771), .ZN(n9939) );
  OAI21_X1 U8545 ( .B1(n6774), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6773), .ZN(
        n6805) );
  MUX2_X1 U8546 ( .A(n6775), .B(P1_REG2_REG_6__SCAN_IN), .S(n6776), .Z(n6804)
         );
  NOR2_X1 U8547 ( .A1(n6805), .A2(n6804), .ZN(n6803) );
  OAI21_X1 U8548 ( .B1(n9946), .B2(P1_REG2_REG_8__SCAN_IN), .A(n9947), .ZN(
        n6779) );
  NAND2_X1 U8549 ( .A1(n6872), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6777) );
  OAI21_X1 U8550 ( .B1(n6872), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6777), .ZN(
        n6778) );
  NOR2_X1 U8551 ( .A1(n6778), .A2(n6779), .ZN(n6871) );
  AOI211_X1 U8552 ( .C1(n6779), .C2(n6778), .A(n6871), .B(n9986), .ZN(n6780)
         );
  AOI211_X1 U8553 ( .C1(n9998), .C2(n6782), .A(n6781), .B(n6780), .ZN(n6783)
         );
  INV_X1 U8554 ( .A(n6783), .ZN(P1_U3250) );
  INV_X1 U8555 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6797) );
  NOR2_X1 U8556 ( .A1(n6785), .A2(n6784), .ZN(n6786) );
  NOR2_X1 U8557 ( .A1(n6787), .A2(n6786), .ZN(n6795) );
  NAND2_X1 U8558 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3084), .ZN(n6788) );
  OAI21_X1 U8559 ( .B1(n9491), .B2(n6789), .A(n6788), .ZN(n6794) );
  AOI211_X1 U8560 ( .C1(n6792), .C2(n6791), .A(n6790), .B(n9986), .ZN(n6793)
         );
  AOI211_X1 U8561 ( .C1(n9998), .C2(n6795), .A(n6794), .B(n6793), .ZN(n6796)
         );
  OAI21_X1 U8562 ( .B1(n9984), .B2(n6797), .A(n6796), .ZN(P1_U3244) );
  INV_X1 U8563 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6810) );
  OAI21_X1 U8564 ( .B1(n6800), .B2(n6799), .A(n6798), .ZN(n6808) );
  NOR2_X1 U8565 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8449), .ZN(n7289) );
  INV_X1 U8566 ( .A(n7289), .ZN(n6801) );
  OAI21_X1 U8567 ( .B1(n9491), .B2(n6802), .A(n6801), .ZN(n6807) );
  AOI211_X1 U8568 ( .C1(n6805), .C2(n6804), .A(n6803), .B(n9986), .ZN(n6806)
         );
  AOI211_X1 U8569 ( .C1(n9998), .C2(n6808), .A(n6807), .B(n6806), .ZN(n6809)
         );
  OAI21_X1 U8570 ( .B1(n9984), .B2(n6810), .A(n6809), .ZN(P1_U3247) );
  NAND2_X1 U8571 ( .A1(n8263), .A2(n6811), .ZN(n6829) );
  AOI22_X1 U8572 ( .A1(n10138), .A2(n6491), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n6829), .ZN(n6816) );
  INV_X1 U8573 ( .A(n6497), .ZN(n6833) );
  OAI22_X1 U8574 ( .A1(n8315), .A2(n6833), .B1(n7109), .B2(n10098), .ZN(n6814)
         );
  NAND2_X1 U8575 ( .A1(n6814), .A2(n6813), .ZN(n6815) );
  OAI211_X1 U8576 ( .C1(n8327), .C2(n7109), .A(n6816), .B(n6815), .ZN(P2_U3234) );
  INV_X1 U8577 ( .A(n6491), .ZN(n6897) );
  AOI22_X1 U8578 ( .A1(n10138), .A2(n8337), .B1(n10136), .B2(n6913), .ZN(n6823) );
  OAI21_X1 U8579 ( .B1(n6819), .B2(n6818), .A(n6817), .ZN(n6820) );
  INV_X1 U8580 ( .A(n6820), .ZN(n6821) );
  AOI22_X1 U8581 ( .A1(n10145), .A2(n6821), .B1(n6829), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n6822) );
  OAI211_X1 U8582 ( .C1(n10095), .C2(n6897), .A(n6823), .B(n6822), .ZN(
        P2_U3239) );
  NAND2_X1 U8583 ( .A1(n6825), .A2(n6824), .ZN(n6826) );
  AOI21_X1 U8584 ( .B1(n6827), .B2(n6826), .A(n10098), .ZN(n6828) );
  AOI21_X1 U8585 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n6829), .A(n6828), .ZN(
        n6832) );
  INV_X1 U8586 ( .A(n6894), .ZN(n6830) );
  AOI22_X1 U8587 ( .A1(n10138), .A2(n10111), .B1(n10136), .B2(n6830), .ZN(
        n6831) );
  OAI211_X1 U8588 ( .C1(n6833), .C2(n10095), .A(n6832), .B(n6831), .ZN(
        P2_U3224) );
  INV_X1 U8589 ( .A(n6834), .ZN(n6836) );
  NAND4_X1 U8590 ( .A1(n6836), .A2(n10051), .A3(n6835), .A4(n7131), .ZN(n6946)
         );
  AOI22_X1 U8591 ( .A1(n9142), .A2(n10034), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n6946), .ZN(n6841) );
  OAI21_X1 U8592 ( .B1(n6839), .B2(n6837), .A(n6838), .ZN(n6965) );
  NAND2_X1 U8593 ( .A1(n6965), .A2(n9160), .ZN(n6840) );
  OAI211_X1 U8594 ( .C1(n6842), .C2(n9162), .A(n6841), .B(n6840), .ZN(P1_U3230) );
  AOI22_X1 U8595 ( .A1(n8382), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n8381), .ZN(n6847) );
  NAND2_X1 U8596 ( .A1(n8382), .A2(n6843), .ZN(n6844) );
  OAI211_X1 U8597 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n8377), .A(n6844), .B(
        n8376), .ZN(n6845) );
  INV_X1 U8598 ( .A(n6845), .ZN(n6846) );
  MUX2_X1 U8599 ( .A(n6847), .B(n6846), .S(P2_IR_REG_0__SCAN_IN), .Z(n6849) );
  AOI22_X1 U8600 ( .A1(n8350), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n6848) );
  NAND2_X1 U8601 ( .A1(n6849), .A2(n6848), .ZN(P2_U3245) );
  NAND2_X1 U8602 ( .A1(n6851), .A2(n6850), .ZN(n6852) );
  INV_X1 U8603 ( .A(n6855), .ZN(n6859) );
  OR3_X1 U8604 ( .A1(n8179), .A2(n8170), .A3(n8865), .ZN(n10228) );
  OAI22_X1 U8605 ( .A1(n6856), .A2(n10248), .B1(n6894), .B2(n10255), .ZN(n6858) );
  AOI211_X1 U8606 ( .C1(n6859), .C2(n10259), .A(n6858), .B(n6857), .ZN(n6926)
         );
  OR2_X1 U8607 ( .A1(n4393), .A2(n5928), .ZN(n6860) );
  OAI21_X1 U8608 ( .B1(n10260), .B2(n6926), .A(n6860), .ZN(P2_U3454) );
  INV_X1 U8609 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6879) );
  MUX2_X1 U8610 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6861), .S(n7220), .Z(n6867)
         );
  NAND2_X1 U8611 ( .A1(n6863), .A2(n6862), .ZN(n6865) );
  NAND2_X1 U8612 ( .A1(n6865), .A2(n6864), .ZN(n6866) );
  NAND2_X1 U8613 ( .A1(n6867), .A2(n6866), .ZN(n7212) );
  OAI21_X1 U8614 ( .B1(n6867), .B2(n6866), .A(n7212), .ZN(n6877) );
  NOR2_X1 U8615 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6868), .ZN(n7683) );
  INV_X1 U8616 ( .A(n7683), .ZN(n6869) );
  OAI21_X1 U8617 ( .B1(n9491), .B2(n6870), .A(n6869), .ZN(n6876) );
  XNOR2_X1 U8618 ( .A(n7220), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n6873) );
  AOI211_X1 U8619 ( .C1(n6874), .C2(n6873), .A(n7219), .B(n9986), .ZN(n6875)
         );
  AOI211_X1 U8620 ( .C1(n9998), .C2(n6877), .A(n6876), .B(n6875), .ZN(n6878)
         );
  OAI21_X1 U8621 ( .B1(n9984), .B2(n6879), .A(n6878), .ZN(P1_U3251) );
  AND2_X1 U8622 ( .A1(n5593), .A2(n7205), .ZN(n9409) );
  NOR2_X1 U8623 ( .A1(n9409), .A2(n7199), .ZN(n9301) );
  INV_X1 U8624 ( .A(n6880), .ZN(n9450) );
  NOR3_X1 U8625 ( .A1(n9301), .A2(n9450), .A3(n6881), .ZN(n6882) );
  AOI21_X1 U8626 ( .B1(n9818), .B2(n5597), .A(n6882), .ZN(n10037) );
  OAI21_X1 U8627 ( .B1(n7205), .B2(n10032), .A(n10037), .ZN(n9828) );
  NAND2_X1 U8628 ( .A1(n9828), .A2(n10076), .ZN(n6883) );
  OAI21_X1 U8629 ( .B1(n10076), .B2(n6884), .A(n6883), .ZN(P1_U3454) );
  INV_X1 U8630 ( .A(n6885), .ZN(n6890) );
  AOI21_X1 U8631 ( .B1(n6887), .B2(n6889), .A(n6886), .ZN(n6888) );
  AOI21_X1 U8632 ( .B1(n6890), .B2(n6889), .A(n6888), .ZN(n6893) );
  AOI22_X1 U8633 ( .A1(n9142), .A2(n4388), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n6946), .ZN(n6892) );
  INV_X1 U8634 ( .A(n9162), .ZN(n9116) );
  AOI22_X1 U8635 ( .A1(n9116), .A2(n9470), .B1(n9167), .B2(n5593), .ZN(n6891)
         );
  OAI211_X1 U8636 ( .C1(n6893), .C2(n9144), .A(n6892), .B(n6891), .ZN(P1_U3220) );
  NAND2_X1 U8637 ( .A1(n6895), .A2(n6894), .ZN(n6900) );
  INV_X1 U8638 ( .A(n6896), .ZN(n6898) );
  NAND2_X1 U8639 ( .A1(n6898), .A2(n6897), .ZN(n6899) );
  NAND2_X1 U8640 ( .A1(n6900), .A2(n6899), .ZN(n7043) );
  OR2_X2 U8641 ( .A1(n10111), .A2(n10195), .ZN(n7989) );
  NAND2_X1 U8642 ( .A1(n10111), .A2(n10195), .ZN(n7991) );
  NAND2_X2 U8643 ( .A1(n7989), .A2(n7991), .ZN(n8146) );
  NAND2_X1 U8644 ( .A1(n7043), .A2(n8146), .ZN(n7042) );
  OR2_X1 U8645 ( .A1(n10111), .A2(n6913), .ZN(n6901) );
  NAND2_X1 U8646 ( .A1(n7042), .A2(n6901), .ZN(n6904) );
  NAND2_X1 U8647 ( .A1(n8337), .A2(n6912), .ZN(n7994) );
  NAND2_X1 U8648 ( .A1(n6904), .A2(n6905), .ZN(n7082) );
  OAI21_X1 U8649 ( .B1(n6904), .B2(n6905), .A(n7082), .ZN(n7148) );
  INV_X1 U8650 ( .A(n7148), .ZN(n6916) );
  AOI22_X1 U8651 ( .A1(n8877), .A2(n10111), .B1(n10139), .B2(n8879), .ZN(n6911) );
  INV_X1 U8652 ( .A(n6905), .ZN(n6907) );
  INV_X1 U8653 ( .A(n8146), .ZN(n7040) );
  AND2_X1 U8654 ( .A1(n6906), .A2(n7988), .ZN(n7039) );
  NAND2_X1 U8655 ( .A1(n7040), .A2(n7039), .ZN(n7038) );
  NAND2_X1 U8656 ( .A1(n7038), .A2(n7989), .ZN(n6908) );
  NAND2_X1 U8657 ( .A1(n6908), .A2(n6907), .ZN(n7091) );
  OAI21_X1 U8658 ( .B1(n6907), .B2(n6908), .A(n7091), .ZN(n6909) );
  NAND2_X1 U8659 ( .A1(n6909), .A2(n10156), .ZN(n6910) );
  OAI211_X1 U8660 ( .C1(n6916), .C2(n7568), .A(n6911), .B(n6910), .ZN(n7149)
         );
  INV_X1 U8661 ( .A(n7149), .ZN(n6915) );
  AOI211_X1 U8662 ( .C1(n6902), .C2(n7037), .A(n10248), .B(n7160), .ZN(n7145)
         );
  AOI21_X1 U8663 ( .B1(n6902), .B2(n10213), .A(n7145), .ZN(n6914) );
  OAI211_X1 U8664 ( .C1(n6916), .C2(n10228), .A(n6915), .B(n6914), .ZN(n6922)
         );
  NAND2_X1 U8665 ( .A1(n6922), .A2(n4393), .ZN(n6917) );
  OAI21_X1 U8666 ( .B1(n4393), .B2(n5967), .A(n6917), .ZN(P2_U3460) );
  INV_X1 U8667 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6924) );
  NAND2_X1 U8668 ( .A1(n6922), .A2(n10275), .ZN(n6923) );
  OAI21_X1 U8669 ( .B1(n10275), .B2(n6924), .A(n6923), .ZN(P2_U3523) );
  OR2_X1 U8670 ( .A1(n10275), .A2(n6629), .ZN(n6925) );
  OAI21_X1 U8671 ( .B1(n10273), .B2(n6926), .A(n6925), .ZN(P2_U3521) );
  NAND2_X1 U8672 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7016) );
  INV_X1 U8673 ( .A(n7016), .ZN(n6933) );
  INV_X1 U8674 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6929) );
  MUX2_X1 U8675 ( .A(n6929), .B(P2_REG1_REG_9__SCAN_IN), .S(n6984), .Z(n6930)
         );
  NOR2_X1 U8676 ( .A1(n6931), .A2(n6930), .ZN(n6983) );
  AOI211_X1 U8677 ( .C1(n6931), .C2(n6930), .A(n6983), .B(n8377), .ZN(n6932)
         );
  AOI211_X1 U8678 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n8350), .A(n6933), .B(
        n6932), .ZN(n6939) );
  OAI21_X1 U8679 ( .B1(n6935), .B2(n7180), .A(n6934), .ZN(n6937) );
  MUX2_X1 U8680 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7278), .S(n6984), .Z(n6936)
         );
  NAND2_X1 U8681 ( .A1(n6936), .A2(n6937), .ZN(n6990) );
  OAI211_X1 U8682 ( .C1(n6937), .C2(n6936), .A(n8382), .B(n6990), .ZN(n6938)
         );
  OAI211_X1 U8683 ( .C1(n8376), .C2(n6991), .A(n6939), .B(n6938), .ZN(P2_U3254) );
  INV_X1 U8684 ( .A(n7893), .ZN(n7887) );
  INV_X1 U8685 ( .A(n6940), .ZN(n6941) );
  OAI222_X1 U8686 ( .A1(n7887), .A2(P2_U3152), .B1(n9021), .B2(n6941), .C1(
        n8464), .C2(n9018), .ZN(P2_U3343) );
  OAI222_X1 U8687 ( .A1(n9874), .A2(n8557), .B1(n9878), .B2(n6941), .C1(
        P1_U3084), .C2(n7942), .ZN(P1_U3338) );
  INV_X1 U8688 ( .A(n6942), .ZN(n6951) );
  INV_X1 U8689 ( .A(n9477), .ZN(n6943) );
  OAI222_X1 U8690 ( .A1(n9878), .A2(n6951), .B1(n6943), .B2(P1_U3084), .C1(
        n8634), .C2(n9874), .ZN(P1_U3337) );
  XOR2_X1 U8691 ( .A(n6945), .B(n6944), .Z(n6949) );
  AOI22_X1 U8692 ( .A1(n9142), .A2(n6998), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n6946), .ZN(n6948) );
  AOI22_X1 U8693 ( .A1(n9116), .A2(n9469), .B1(n9167), .B2(n5597), .ZN(n6947)
         );
  OAI211_X1 U8694 ( .C1(n6949), .C2(n9144), .A(n6948), .B(n6947), .ZN(P1_U3235) );
  INV_X1 U8695 ( .A(n8345), .ZN(n7903) );
  OAI222_X1 U8696 ( .A1(P2_U3152), .A2(n7903), .B1(n9021), .B2(n6951), .C1(
        n6950), .C2(n9018), .ZN(P2_U3342) );
  INV_X1 U8697 ( .A(n6952), .ZN(n6980) );
  AOI22_X1 U8698 ( .A1(n9487), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9871), .ZN(n6953) );
  OAI21_X1 U8699 ( .B1(n6980), .B2(n9878), .A(n6953), .ZN(P1_U3336) );
  OAI211_X1 U8700 ( .C1(n6956), .C2(n6955), .A(n9998), .B(n6954), .ZN(n6964)
         );
  OAI22_X1 U8701 ( .A1(n9491), .A2(n6957), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7135), .ZN(n6958) );
  INV_X1 U8702 ( .A(n6958), .ZN(n6963) );
  OAI211_X1 U8703 ( .C1(n6961), .C2(n6960), .A(n9966), .B(n6959), .ZN(n6962)
         );
  NAND3_X1 U8704 ( .A1(n6964), .A2(n6963), .A3(n6962), .ZN(n6971) );
  INV_X1 U8705 ( .A(n6965), .ZN(n6966) );
  MUX2_X1 U8706 ( .A(n6967), .B(n6966), .S(n7861), .Z(n6970) );
  AOI211_X1 U8707 ( .C1(n6970), .C2(n9449), .A(n6969), .B(n6968), .ZN(n9926)
         );
  AOI211_X1 U8708 ( .C1(n9997), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n6971), .B(
        n9926), .ZN(n6972) );
  INV_X1 U8709 ( .A(n6972), .ZN(P1_U3243) );
  XOR2_X1 U8710 ( .A(n6973), .B(n6974), .Z(n6978) );
  MUX2_X1 U8711 ( .A(n9092), .B(P1_U3084), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n6976) );
  OAI22_X1 U8712 ( .A1(n9139), .A2(n7312), .B1(n10057), .B2(n9170), .ZN(n6975)
         );
  AOI211_X1 U8713 ( .C1(n9116), .C2(n9468), .A(n6976), .B(n6975), .ZN(n6977)
         );
  OAI21_X1 U8714 ( .B1(n6978), .B2(n9144), .A(n6977), .ZN(P1_U3216) );
  INV_X1 U8715 ( .A(n8358), .ZN(n8353) );
  OAI222_X1 U8716 ( .A1(P2_U3152), .A2(n8353), .B1(n9021), .B2(n6980), .C1(
        n6979), .C2(n9018), .ZN(P2_U3341) );
  NAND2_X1 U8717 ( .A1(n9471), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6981) );
  OAI21_X1 U8718 ( .B1(n6982), .B2(n9471), .A(n6981), .ZN(P1_U3584) );
  NOR2_X1 U8719 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8483), .ZN(n6989) );
  INV_X1 U8720 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6985) );
  MUX2_X1 U8721 ( .A(n6985), .B(P2_REG1_REG_10__SCAN_IN), .S(n7071), .Z(n6986)
         );
  AOI211_X1 U8722 ( .C1(n6987), .C2(n6986), .A(n7070), .B(n8377), .ZN(n6988)
         );
  AOI211_X1 U8723 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n8350), .A(n6989), .B(
        n6988), .ZN(n6996) );
  OAI21_X1 U8724 ( .B1(n6991), .B2(n7278), .A(n6990), .ZN(n6994) );
  MUX2_X1 U8725 ( .A(n7357), .B(P2_REG2_REG_10__SCAN_IN), .S(n7071), .Z(n6992)
         );
  INV_X1 U8726 ( .A(n6992), .ZN(n6993) );
  NAND2_X1 U8727 ( .A1(n6993), .A2(n6994), .ZN(n7064) );
  OAI211_X1 U8728 ( .C1(n6994), .C2(n6993), .A(n8382), .B(n7064), .ZN(n6995)
         );
  OAI211_X1 U8729 ( .C1(n8376), .C2(n6997), .A(n6996), .B(n6995), .ZN(P2_U3255) );
  AOI211_X1 U8730 ( .C1(n6998), .C2(n7204), .A(n9695), .B(n7318), .ZN(n7137)
         );
  NAND2_X1 U8731 ( .A1(n6999), .A2(n9302), .ZN(n7000) );
  NAND2_X1 U8732 ( .A1(n7001), .A2(n7000), .ZN(n7002) );
  NAND2_X1 U8733 ( .A1(n7002), .A2(n10066), .ZN(n7007) );
  AOI22_X1 U8734 ( .A1(n9818), .A2(n9469), .B1(n5597), .B2(n9819), .ZN(n7006)
         );
  XNOR2_X1 U8735 ( .A(n9302), .B(n7003), .ZN(n7004) );
  NAND2_X1 U8736 ( .A1(n7004), .A2(n9637), .ZN(n7005) );
  NAND3_X1 U8737 ( .A1(n7007), .A2(n7006), .A3(n7005), .ZN(n7138) );
  NOR2_X1 U8738 ( .A1(n7137), .A2(n7138), .ZN(n7011) );
  OAI22_X1 U8739 ( .A1(n9864), .A2(n5607), .B1(n10076), .B2(n4972), .ZN(n7008)
         );
  INV_X1 U8740 ( .A(n7008), .ZN(n7009) );
  OAI21_X1 U8741 ( .B1(n7011), .B2(n10075), .A(n7009), .ZN(P1_U3460) );
  INV_X1 U8742 ( .A(n9815), .ZN(n7604) );
  AOI22_X1 U8743 ( .A1(n7604), .A2(n6998), .B1(n10081), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n7010) );
  OAI21_X1 U8744 ( .B1(n7011), .B2(n10081), .A(n7010), .ZN(P1_U3525) );
  INV_X1 U8745 ( .A(n7012), .ZN(n10122) );
  NOR3_X1 U8746 ( .A1(n8315), .A2(n7268), .A3(n7013), .ZN(n7014) );
  AOI21_X1 U8747 ( .B1(n10122), .B2(n10145), .A(n7014), .ZN(n7023) );
  INV_X1 U8748 ( .A(n7015), .ZN(n7020) );
  INV_X1 U8749 ( .A(n7268), .ZN(n10084) );
  NAND2_X1 U8750 ( .A1(n10140), .A2(n10084), .ZN(n7017) );
  OAI211_X1 U8751 ( .C1(n10152), .C2(n7277), .A(n7017), .B(n7016), .ZN(n7019)
         );
  INV_X1 U8752 ( .A(n7341), .ZN(n10234) );
  OAI22_X1 U8753 ( .A1(n10130), .A2(n7405), .B1(n8327), .B2(n10234), .ZN(n7018) );
  AOI211_X1 U8754 ( .C1(n7020), .C2(n10145), .A(n7019), .B(n7018), .ZN(n7021)
         );
  OAI21_X1 U8755 ( .B1(n7023), .B2(n7022), .A(n7021), .ZN(P2_U3233) );
  INV_X1 U8756 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7025) );
  INV_X1 U8757 ( .A(n7024), .ZN(n7027) );
  INV_X1 U8758 ( .A(n9993), .ZN(n7940) );
  OAI222_X1 U8759 ( .A1(n9874), .A2(n7025), .B1(n9878), .B2(n7027), .C1(
        P1_U3084), .C2(n7940), .ZN(P1_U3335) );
  INV_X1 U8760 ( .A(n8375), .ZN(n8362) );
  INV_X1 U8761 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7026) );
  OAI222_X1 U8762 ( .A1(n8362), .A2(P2_U3152), .B1(n9021), .B2(n7027), .C1(
        n7026), .C2(n9018), .ZN(P2_U3340) );
  INV_X1 U8763 ( .A(n7029), .ZN(n7030) );
  AOI211_X1 U8764 ( .C1(n7031), .C2(n7028), .A(n9144), .B(n7030), .ZN(n7035)
         );
  AOI22_X1 U8765 ( .A1(n9116), .A2(n9467), .B1(n9167), .B2(n9469), .ZN(n7033)
         );
  INV_X1 U8766 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n8461) );
  NOR2_X1 U8767 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8461), .ZN(n9927) );
  AOI21_X1 U8768 ( .B1(n9142), .B2(n7371), .A(n9927), .ZN(n7032) );
  OAI211_X1 U8769 ( .C1(n9164), .C2(n7369), .A(n7033), .B(n7032), .ZN(n7034)
         );
  OR2_X1 U8770 ( .A1(n7035), .A2(n7034), .ZN(P1_U3228) );
  OAI22_X1 U8771 ( .A1(n6643), .A2(n8881), .B1(n6706), .B2(n8888), .ZN(n7047)
         );
  OAI21_X1 U8772 ( .B1(n4539), .B2(n10195), .A(n7037), .ZN(n10196) );
  OAI21_X1 U8773 ( .B1(n7040), .B2(n7039), .A(n7038), .ZN(n7041) );
  AOI222_X1 U8774 ( .A1(n10156), .A2(n7041), .B1(n8337), .B2(n8879), .C1(n6491), .C2(n8877), .ZN(n10197) );
  OAI22_X1 U8775 ( .A1(n8780), .A2(n10196), .B1(n4392), .B2(n10197), .ZN(n7046) );
  OAI21_X1 U8776 ( .B1(n7043), .B2(n8146), .A(n7042), .ZN(n10200) );
  INV_X1 U8777 ( .A(n10200), .ZN(n7044) );
  OAI22_X1 U8778 ( .A1(n10195), .A2(n8869), .B1(n8874), .B2(n7044), .ZN(n7045)
         );
  OR3_X1 U8779 ( .A1(n7047), .A2(n7046), .A3(n7045), .ZN(P2_U3294) );
  OAI21_X1 U8780 ( .B1(n7048), .B2(n7051), .A(n7383), .ZN(n7379) );
  AOI21_X1 U8781 ( .B1(n7317), .B2(n7371), .A(n9695), .ZN(n7049) );
  NAND2_X1 U8782 ( .A1(n7049), .A2(n7393), .ZN(n7377) );
  AOI22_X1 U8783 ( .A1(n9467), .A2(n9818), .B1(n9819), .B2(n9469), .ZN(n7050)
         );
  NAND2_X1 U8784 ( .A1(n7377), .A2(n7050), .ZN(n7053) );
  XNOR2_X1 U8785 ( .A(n9172), .B(n7051), .ZN(n7052) );
  NOR2_X1 U8786 ( .A1(n7052), .A2(n10020), .ZN(n7368) );
  AOI211_X1 U8787 ( .C1(n10066), .C2(n7379), .A(n7053), .B(n7368), .ZN(n7059)
         );
  AOI22_X1 U8788 ( .A1(n7604), .A2(n7371), .B1(n10081), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n7054) );
  OAI21_X1 U8789 ( .B1(n7059), .B2(n10081), .A(n7054), .ZN(P1_U3527) );
  INV_X1 U8790 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7055) );
  OAI22_X1 U8791 ( .A1(n9864), .A2(n7056), .B1(n10076), .B2(n7055), .ZN(n7057)
         );
  INV_X1 U8792 ( .A(n7057), .ZN(n7058) );
  OAI21_X1 U8793 ( .B1(n7059), .B2(n10075), .A(n7058), .ZN(P1_U3466) );
  INV_X1 U8794 ( .A(n7060), .ZN(n7063) );
  OAI222_X1 U8795 ( .A1(n9874), .A2(n7061), .B1(n9878), .B2(n7063), .C1(n4390), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  OAI222_X1 U8796 ( .A1(n8865), .A2(P2_U3152), .B1(n9021), .B2(n7063), .C1(
        n7062), .C2(n9018), .ZN(P2_U3339) );
  NAND2_X1 U8797 ( .A1(n7071), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7065) );
  NAND2_X1 U8798 ( .A1(n7065), .A2(n7064), .ZN(n7068) );
  MUX2_X1 U8799 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n7420), .S(n7253), .Z(n7066)
         );
  INV_X1 U8800 ( .A(n7066), .ZN(n7067) );
  NOR2_X1 U8801 ( .A1(n7068), .A2(n7067), .ZN(n7247) );
  AOI21_X1 U8802 ( .B1(n7068), .B2(n7067), .A(n7247), .ZN(n7080) );
  INV_X1 U8803 ( .A(n8382), .ZN(n8368) );
  NOR2_X1 U8804 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6120), .ZN(n7123) );
  AOI21_X1 U8805 ( .B1(n8350), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7123), .ZN(
        n7076) );
  INV_X1 U8806 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7069) );
  MUX2_X1 U8807 ( .A(n7069), .B(P2_REG1_REG_11__SCAN_IN), .S(n7253), .Z(n7073)
         );
  AOI21_X1 U8808 ( .B1(n7073), .B2(n7072), .A(n7252), .ZN(n7074) );
  NAND2_X1 U8809 ( .A1(n8381), .A2(n7074), .ZN(n7075) );
  OAI211_X1 U8810 ( .C1(n8376), .C2(n7077), .A(n7076), .B(n7075), .ZN(n7078)
         );
  INV_X1 U8811 ( .A(n7078), .ZN(n7079) );
  OAI21_X1 U8812 ( .B1(n7080), .B2(n8368), .A(n7079), .ZN(P2_U3256) );
  OR2_X1 U8813 ( .A1(n10085), .A2(n7168), .ZN(n8002) );
  NAND2_X1 U8814 ( .A1(n10085), .A2(n7168), .ZN(n8001) );
  OR2_X1 U8815 ( .A1(n8337), .A2(n6902), .ZN(n7081) );
  NAND2_X1 U8816 ( .A1(n7082), .A2(n7081), .ZN(n7159) );
  OR2_X1 U8817 ( .A1(n10139), .A2(n10202), .ZN(n7981) );
  NAND2_X1 U8818 ( .A1(n10139), .A2(n10202), .ZN(n7995) );
  NAND2_X1 U8819 ( .A1(n7159), .A2(n8147), .ZN(n7158) );
  INV_X1 U8820 ( .A(n10202), .ZN(n7164) );
  OR2_X1 U8821 ( .A1(n10139), .A2(n7164), .ZN(n7083) );
  NAND2_X1 U8822 ( .A1(n7158), .A2(n7083), .ZN(n7106) );
  NAND2_X1 U8823 ( .A1(n7155), .A2(n10135), .ZN(n7984) );
  INV_X1 U8824 ( .A(n10135), .ZN(n10209) );
  NAND2_X1 U8825 ( .A1(n8878), .A2(n10209), .ZN(n7997) );
  NAND2_X1 U8826 ( .A1(n7984), .A2(n7997), .ZN(n8149) );
  NAND2_X1 U8827 ( .A1(n7106), .A2(n8149), .ZN(n7085) );
  OR2_X1 U8828 ( .A1(n8878), .A2(n10135), .ZN(n7084) );
  NAND2_X1 U8829 ( .A1(n7085), .A2(n7084), .ZN(n8892) );
  INV_X1 U8830 ( .A(n8892), .ZN(n7087) );
  OR2_X1 U8831 ( .A1(n10214), .A2(n7102), .ZN(n7996) );
  NAND2_X1 U8832 ( .A1(n7102), .A2(n10214), .ZN(n7999) );
  INV_X1 U8833 ( .A(n7102), .ZN(n10137) );
  NAND2_X1 U8834 ( .A1(n10214), .A2(n10137), .ZN(n7088) );
  INV_X1 U8835 ( .A(n7170), .ZN(n7089) );
  AOI21_X1 U8836 ( .B1(n8151), .B2(n7090), .A(n7089), .ZN(n10221) );
  INV_X1 U8837 ( .A(n7997), .ZN(n7092) );
  NAND2_X1 U8838 ( .A1(n8876), .A2(n8893), .ZN(n8875) );
  XNOR2_X1 U8839 ( .A(n7173), .B(n8151), .ZN(n7093) );
  AOI222_X1 U8840 ( .A1(n10137), .A2(n8877), .B1(n10084), .B2(n8879), .C1(
        n10156), .C2(n7093), .ZN(n10224) );
  MUX2_X1 U8841 ( .A(n7094), .B(n10224), .S(n8881), .Z(n7098) );
  INV_X1 U8842 ( .A(n10085), .ZN(n10222) );
  INV_X1 U8843 ( .A(n7181), .ZN(n7095) );
  OAI21_X1 U8844 ( .B1(n10222), .B2(n8885), .A(n7095), .ZN(n10223) );
  OAI22_X1 U8845 ( .A1(n8780), .A2(n10223), .B1(n10092), .B2(n8888), .ZN(n7096) );
  AOI21_X1 U8846 ( .B1(n10161), .B2(n10085), .A(n7096), .ZN(n7097) );
  OAI211_X1 U8847 ( .C1(n10221), .C2(n8874), .A(n7098), .B(n7097), .ZN(
        P2_U3289) );
  INV_X1 U8848 ( .A(n10139), .ZN(n7101) );
  XOR2_X1 U8849 ( .A(n8149), .B(n7099), .Z(n7100) );
  OAI222_X1 U8850 ( .A1(n8858), .A2(n7102), .B1(n8856), .B2(n7101), .C1(n8854), 
        .C2(n7100), .ZN(n10210) );
  XNOR2_X1 U8851 ( .A(n7161), .B(n10209), .ZN(n7103) );
  NAND2_X1 U8852 ( .A1(n7103), .A2(n10215), .ZN(n10208) );
  OAI22_X1 U8853 ( .A1(n10208), .A2(n8734), .B1(n8888), .B2(n10151), .ZN(n7104) );
  NOR2_X1 U8854 ( .A1(n10210), .A2(n7104), .ZN(n7105) );
  MUX2_X1 U8855 ( .A(n8470), .B(n7105), .S(n8881), .Z(n7108) );
  XNOR2_X1 U8856 ( .A(n7106), .B(n8149), .ZN(n10212) );
  INV_X1 U8857 ( .A(n8874), .ZN(n10172) );
  AOI22_X1 U8858 ( .A1(n10212), .A2(n10172), .B1(n10161), .B2(n10135), .ZN(
        n7107) );
  NAND2_X1 U8859 ( .A1(n7108), .A2(n7107), .ZN(P2_U3291) );
  NAND2_X1 U8860 ( .A1(n6497), .A2(n7109), .ZN(n7987) );
  NAND2_X1 U8861 ( .A1(n7110), .A2(n7987), .ZN(n10192) );
  INV_X1 U8862 ( .A(n10192), .ZN(n7115) );
  AOI22_X1 U8863 ( .A1(n10192), .A2(n10156), .B1(n8879), .B2(n6491), .ZN(
        n10194) );
  INV_X1 U8864 ( .A(n8888), .ZN(n10159) );
  NAND2_X1 U8865 ( .A1(n10159), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7111) );
  AOI21_X1 U8866 ( .B1(n10194), .B2(n7111), .A(n4392), .ZN(n7112) );
  AOI21_X1 U8867 ( .B1(n4392), .B2(P2_REG2_REG_0__SCAN_IN), .A(n7112), .ZN(
        n7114) );
  OAI21_X1 U8868 ( .B1(n6504), .B2(n10161), .A(n10191), .ZN(n7113) );
  OAI211_X1 U8869 ( .C1(n7115), .C2(n8874), .A(n7114), .B(n7113), .ZN(P2_U3296) );
  INV_X1 U8870 ( .A(n7562), .ZN(n10247) );
  INV_X1 U8871 ( .A(n7116), .ZN(n7117) );
  AOI21_X1 U8872 ( .B1(n10096), .B2(n7117), .A(n10098), .ZN(n7121) );
  NOR3_X1 U8873 ( .A1(n8315), .A2(n7405), .A3(n7118), .ZN(n7120) );
  OAI21_X1 U8874 ( .B1(n7121), .B2(n7120), .A(n7119), .ZN(n7125) );
  INV_X1 U8875 ( .A(n7576), .ZN(n8334) );
  OAI22_X1 U8876 ( .A1(n10095), .A2(n7405), .B1(n10152), .B2(n7419), .ZN(n7122) );
  AOI211_X1 U8877 ( .C1(n10138), .C2(n8334), .A(n7123), .B(n7122), .ZN(n7124)
         );
  OAI211_X1 U8878 ( .C1(n10247), .C2(n8327), .A(n7125), .B(n7124), .ZN(
        P2_U3238) );
  OR2_X1 U8879 ( .A1(n7127), .A2(n7126), .ZN(n10049) );
  NAND2_X1 U8880 ( .A1(n7129), .A2(n7128), .ZN(n7130) );
  NOR2_X1 U8881 ( .A1(n10049), .A2(n7130), .ZN(n7132) );
  NAND2_X1 U8882 ( .A1(n7132), .A2(n7131), .ZN(n7133) );
  INV_X2 U8883 ( .A(n10024), .ZN(n9629) );
  OAI22_X1 U8884 ( .A1(n9623), .A2(n5607), .B1(n7135), .B2(n10008), .ZN(n7136)
         );
  AOI21_X1 U8885 ( .B1(n7137), .B2(n10006), .A(n7136), .ZN(n7141) );
  MUX2_X1 U8886 ( .A(n7138), .B(P1_REG2_REG_2__SCAN_IN), .S(n10024), .Z(n7139)
         );
  INV_X1 U8887 ( .A(n7139), .ZN(n7140) );
  NAND2_X1 U8888 ( .A1(n7141), .A2(n7140), .ZN(P1_U3289) );
  INV_X1 U8889 ( .A(n7142), .ZN(n7143) );
  AND2_X1 U8890 ( .A1(n8881), .A2(n7143), .ZN(n7818) );
  INV_X1 U8891 ( .A(n7144), .ZN(n10171) );
  AOI22_X1 U8892 ( .A1(n10171), .A2(n7145), .B1(n10159), .B2(n5966), .ZN(n7146) );
  OAI21_X1 U8893 ( .B1(n6645), .B2(n8881), .A(n7146), .ZN(n7147) );
  AOI21_X1 U8894 ( .B1(n7818), .B2(n7148), .A(n7147), .ZN(n7151) );
  AOI22_X1 U8895 ( .A1(n8881), .A2(n7149), .B1(n10161), .B2(n6902), .ZN(n7150)
         );
  NAND2_X1 U8896 ( .A1(n7151), .A2(n7150), .ZN(P2_U3293) );
  INV_X1 U8897 ( .A(n8147), .ZN(n7153) );
  XNOR2_X1 U8898 ( .A(n7152), .B(n7153), .ZN(n7157) );
  NAND2_X1 U8899 ( .A1(n8337), .A2(n8877), .ZN(n7154) );
  OAI21_X1 U8900 ( .B1(n7155), .B2(n8858), .A(n7154), .ZN(n7156) );
  AOI21_X1 U8901 ( .B1(n7157), .B2(n10156), .A(n7156), .ZN(n10204) );
  OAI21_X1 U8902 ( .B1(n7159), .B2(n8147), .A(n7158), .ZN(n10207) );
  AOI22_X1 U8903 ( .A1(n10172), .A2(n10207), .B1(n10161), .B2(n7164), .ZN(
        n7167) );
  INV_X1 U8904 ( .A(n7160), .ZN(n7163) );
  INV_X1 U8905 ( .A(n7161), .ZN(n7162) );
  AOI21_X1 U8906 ( .B1(n7164), .B2(n7163), .A(n7162), .ZN(n10201) );
  OAI22_X1 U8907 ( .A1(n8881), .A2(n6646), .B1(n8279), .B2(n8888), .ZN(n7165)
         );
  AOI21_X1 U8908 ( .B1(n6504), .B2(n10201), .A(n7165), .ZN(n7166) );
  OAI211_X1 U8909 ( .C1(n4392), .C2(n10204), .A(n7167), .B(n7166), .ZN(
        P2_U3292) );
  INV_X1 U8910 ( .A(n7168), .ZN(n10126) );
  OR2_X1 U8911 ( .A1(n10085), .A2(n10126), .ZN(n7169) );
  OR2_X1 U8912 ( .A1(n10125), .A2(n7268), .ZN(n8006) );
  NAND2_X1 U8913 ( .A1(n10125), .A2(n7268), .ZN(n8007) );
  NAND2_X1 U8914 ( .A1(n7412), .A2(n8150), .ZN(n7171) );
  INV_X1 U8915 ( .A(n10233), .ZN(n7187) );
  INV_X1 U8916 ( .A(n7818), .ZN(n7587) );
  INV_X1 U8917 ( .A(n8150), .ZN(n7176) );
  INV_X1 U8918 ( .A(n8151), .ZN(n7172) );
  INV_X1 U8919 ( .A(n7269), .ZN(n7174) );
  AOI21_X1 U8920 ( .B1(n7176), .B2(n7175), .A(n7174), .ZN(n7179) );
  INV_X1 U8921 ( .A(n10129), .ZN(n8336) );
  AOI22_X1 U8922 ( .A1(n8877), .A2(n10126), .B1(n8336), .B2(n8879), .ZN(n7178)
         );
  INV_X1 U8923 ( .A(n7568), .ZN(n7811) );
  NAND2_X1 U8924 ( .A1(n10233), .A2(n7811), .ZN(n7177) );
  OAI211_X1 U8925 ( .C1(n7179), .C2(n8854), .A(n7178), .B(n7177), .ZN(n10231)
         );
  NAND2_X1 U8926 ( .A1(n10231), .A2(n8881), .ZN(n7186) );
  OAI22_X1 U8927 ( .A1(n8881), .A2(n7180), .B1(n10134), .B2(n8888), .ZN(n7184)
         );
  INV_X1 U8928 ( .A(n10125), .ZN(n10229) );
  OR2_X1 U8929 ( .A1(n7181), .A2(n10229), .ZN(n7182) );
  NAND2_X1 U8930 ( .A1(n7275), .A2(n7182), .ZN(n10230) );
  NOR2_X1 U8931 ( .A1(n8780), .A2(n10230), .ZN(n7183) );
  AOI211_X1 U8932 ( .C1(n10161), .C2(n10125), .A(n7184), .B(n7183), .ZN(n7185)
         );
  OAI211_X1 U8933 ( .C1(n7187), .C2(n7587), .A(n7186), .B(n7185), .ZN(P2_U3288) );
  OAI21_X1 U8934 ( .B1(n7190), .B2(n7189), .A(n7188), .ZN(n7194) );
  AOI22_X1 U8935 ( .A1(n9142), .A2(n7394), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        P1_U3084), .ZN(n7192) );
  AOI22_X1 U8936 ( .A1(n9116), .A2(n9466), .B1(n9167), .B2(n9468), .ZN(n7191)
         );
  OAI211_X1 U8937 ( .C1(n9164), .C2(n7395), .A(n7192), .B(n7191), .ZN(n7193)
         );
  AOI21_X1 U8938 ( .B1(n7194), .B2(n9160), .A(n7193), .ZN(n7195) );
  INV_X1 U8939 ( .A(n7195), .ZN(P1_U3225) );
  AOI22_X1 U8940 ( .A1(n10028), .A2(n4388), .B1(n10024), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7209) );
  OAI21_X1 U8941 ( .B1(n9305), .B2(n7197), .A(n7196), .ZN(n7203) );
  AOI22_X1 U8942 ( .A1(n9470), .A2(n9818), .B1(n9819), .B2(n5593), .ZN(n7202)
         );
  NAND2_X1 U8943 ( .A1(n7200), .A2(n9637), .ZN(n7201) );
  OAI211_X1 U8944 ( .C1(n7203), .C2(n7672), .A(n7202), .B(n7201), .ZN(n10054)
         );
  OAI211_X1 U8945 ( .C1(n7205), .C2(n10053), .A(n10003), .B(n7204), .ZN(n10052) );
  OAI22_X1 U8946 ( .A1(n10052), .A2(n4509), .B1(n10008), .B2(n7206), .ZN(n7207) );
  OAI21_X1 U8947 ( .B1(n10054), .B2(n7207), .A(n9629), .ZN(n7208) );
  NAND2_X1 U8948 ( .A1(n7209), .A2(n7208), .ZN(P1_U3290) );
  INV_X1 U8949 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7227) );
  AOI22_X1 U8950 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n9976), .B1(n7210), .B2(
        n5169), .ZN(n9978) );
  INV_X1 U8951 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9915) );
  AOI22_X1 U8952 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n9958), .B1(n7211), .B2(
        n9915), .ZN(n9961) );
  OAI21_X1 U8953 ( .B1(n7220), .B2(P1_REG1_REG_10__SCAN_IN), .A(n7212), .ZN(
        n9960) );
  NAND2_X1 U8954 ( .A1(n9961), .A2(n9960), .ZN(n9959) );
  OAI21_X1 U8955 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9958), .A(n9959), .ZN(
        n9979) );
  NAND2_X1 U8956 ( .A1(n9978), .A2(n9979), .ZN(n9977) );
  OAI21_X1 U8957 ( .B1(n9976), .B2(P1_REG1_REG_12__SCAN_IN), .A(n9977), .ZN(
        n7215) );
  XNOR2_X1 U8958 ( .A(n7544), .B(n7213), .ZN(n7214) );
  NAND2_X1 U8959 ( .A1(n7214), .A2(n7215), .ZN(n7538) );
  OAI21_X1 U8960 ( .B1(n7215), .B2(n7214), .A(n7538), .ZN(n7216) );
  NAND2_X1 U8961 ( .A1(n7216), .A2(n9998), .ZN(n7226) );
  AND2_X1 U8962 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9115) );
  NAND2_X1 U8963 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n9976), .ZN(n7217) );
  OAI21_X1 U8964 ( .B1(n9976), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7217), .ZN(
        n9972) );
  NOR2_X1 U8965 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n9958), .ZN(n7218) );
  AOI21_X1 U8966 ( .B1(n9958), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7218), .ZN(
        n9963) );
  OAI21_X1 U8967 ( .B1(n9958), .B2(P1_REG2_REG_11__SCAN_IN), .A(n9962), .ZN(
        n9973) );
  NOR2_X1 U8968 ( .A1(n9972), .A2(n9973), .ZN(n9971) );
  MUX2_X1 U8969 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n7702), .S(n7544), .Z(n7221)
         );
  INV_X1 U8970 ( .A(n7221), .ZN(n7222) );
  AOI211_X1 U8971 ( .C1(n7223), .C2(n7222), .A(n7543), .B(n9986), .ZN(n7224)
         );
  AOI211_X1 U8972 ( .C1(n9992), .C2(n7544), .A(n9115), .B(n7224), .ZN(n7225)
         );
  OAI211_X1 U8973 ( .C1(n9984), .C2(n7227), .A(n7226), .B(n7225), .ZN(P1_U3254) );
  INV_X1 U8974 ( .A(n7228), .ZN(n7246) );
  OAI222_X1 U8975 ( .A1(n9878), .A2(n7246), .B1(P1_U3084), .B2(n9443), .C1(
        n7229), .C2(n9874), .ZN(P1_U3333) );
  OAI21_X1 U8976 ( .B1(n7231), .B2(n9183), .A(n7230), .ZN(n7471) );
  OAI21_X1 U8977 ( .B1(n7392), .B2(n7469), .A(n10003), .ZN(n7232) );
  NOR2_X1 U8978 ( .A1(n7232), .A2(n7333), .ZN(n7463) );
  OAI22_X1 U8979 ( .A1(n7483), .A2(n10062), .B1(n7373), .B2(n10015), .ZN(n7233) );
  AOI211_X1 U8980 ( .C1(n7471), .C2(n10066), .A(n7463), .B(n7233), .ZN(n7238)
         );
  INV_X1 U8981 ( .A(n7235), .ZN(n7388) );
  INV_X1 U8982 ( .A(n9177), .ZN(n9175) );
  AOI21_X1 U8983 ( .B1(n7234), .B2(n7388), .A(n9175), .ZN(n7236) );
  XNOR2_X1 U8984 ( .A(n7236), .B(n9183), .ZN(n7237) );
  NAND2_X1 U8985 ( .A1(n7237), .A2(n9637), .ZN(n7473) );
  NAND2_X1 U8986 ( .A1(n7238), .A2(n7473), .ZN(n7243) );
  OAI22_X1 U8987 ( .A1(n9815), .A2(n7469), .B1(n10083), .B2(n5028), .ZN(n7239)
         );
  AOI21_X1 U8988 ( .B1(n7243), .B2(n10083), .A(n7239), .ZN(n7240) );
  INV_X1 U8989 ( .A(n7240), .ZN(P1_U3529) );
  INV_X1 U8990 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7241) );
  OAI22_X1 U8991 ( .A1(n9864), .A2(n7469), .B1(n10076), .B2(n7241), .ZN(n7242)
         );
  AOI21_X1 U8992 ( .B1(n7243), .B2(n10076), .A(n7242), .ZN(n7244) );
  INV_X1 U8993 ( .A(n7244), .ZN(P1_U3472) );
  OAI222_X1 U8994 ( .A1(P2_U3152), .A2(n8145), .B1(n9021), .B2(n7246), .C1(
        n7245), .C2(n9018), .ZN(P2_U3338) );
  NOR2_X1 U8995 ( .A1(n7253), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7248) );
  NOR2_X1 U8996 ( .A1(n7248), .A2(n7247), .ZN(n7251) );
  INV_X1 U8997 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7249) );
  MUX2_X1 U8998 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7249), .S(n7433), .Z(n7250)
         );
  NAND2_X1 U8999 ( .A1(n7433), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7429) );
  OAI211_X1 U9000 ( .C1(n7433), .C2(P2_REG2_REG_12__SCAN_IN), .A(n7251), .B(
        n7429), .ZN(n7428) );
  OAI211_X1 U9001 ( .C1(n7251), .C2(n7250), .A(n7428), .B(n8382), .ZN(n7262)
         );
  AOI21_X1 U9002 ( .B1(n7253), .B2(P2_REG1_REG_11__SCAN_IN), .A(n7252), .ZN(
        n7256) );
  MUX2_X1 U9003 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7254), .S(n7433), .Z(n7255)
         );
  NAND2_X1 U9004 ( .A1(n7256), .A2(n7255), .ZN(n7432) );
  OAI21_X1 U9005 ( .B1(n7256), .B2(n7255), .A(n7432), .ZN(n7260) );
  NAND2_X1 U9006 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7300) );
  INV_X1 U9007 ( .A(n7300), .ZN(n7259) );
  INV_X1 U9008 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7257) );
  NOR2_X1 U9009 ( .A1(n8389), .A2(n7257), .ZN(n7258) );
  AOI211_X1 U9010 ( .C1(n8381), .C2(n7260), .A(n7259), .B(n7258), .ZN(n7261)
         );
  OAI211_X1 U9011 ( .C1(n8376), .C2(n7263), .A(n7262), .B(n7261), .ZN(P2_U3257) );
  NAND2_X1 U9012 ( .A1(n10125), .A2(n10084), .ZN(n7264) );
  AND2_X1 U9013 ( .A1(n7265), .A2(n7264), .ZN(n7267) );
  OR2_X1 U9014 ( .A1(n7341), .A2(n10129), .ZN(n7972) );
  NAND2_X1 U9015 ( .A1(n7265), .A2(n7348), .ZN(n7266) );
  OAI21_X1 U9016 ( .B1(n7267), .B2(n8154), .A(n7266), .ZN(n10239) );
  OAI22_X1 U9017 ( .A1(n7405), .A2(n8858), .B1(n7268), .B2(n8856), .ZN(n7274)
         );
  INV_X1 U9018 ( .A(n8154), .ZN(n7270) );
  NAND2_X1 U9019 ( .A1(n7271), .A2(n7270), .ZN(n7353) );
  NAND3_X1 U9020 ( .A1(n7269), .A2(n8007), .A3(n8154), .ZN(n7272) );
  AOI21_X1 U9021 ( .B1(n7353), .B2(n7272), .A(n8854), .ZN(n7273) );
  AOI211_X1 U9022 ( .C1(n10239), .C2(n7811), .A(n7274), .B(n7273), .ZN(n10236)
         );
  NAND2_X1 U9023 ( .A1(n7275), .A2(n7341), .ZN(n7276) );
  NAND2_X1 U9024 ( .A1(n7416), .A2(n7276), .ZN(n10235) );
  OAI22_X1 U9025 ( .A1(n8881), .A2(n7278), .B1(n7277), .B2(n8888), .ZN(n7279)
         );
  AOI21_X1 U9026 ( .B1(n10161), .B2(n7341), .A(n7279), .ZN(n7280) );
  OAI21_X1 U9027 ( .B1(n8780), .B2(n10235), .A(n7280), .ZN(n7281) );
  AOI21_X1 U9028 ( .B1(n10239), .B2(n7818), .A(n7281), .ZN(n7282) );
  OAI21_X1 U9029 ( .B1(n10236), .B2(n4392), .A(n7282), .ZN(P2_U3287) );
  XOR2_X1 U9030 ( .A(n7285), .B(n7284), .Z(n7286) );
  XNOR2_X1 U9031 ( .A(n7283), .B(n7286), .ZN(n7292) );
  INV_X1 U9032 ( .A(n7464), .ZN(n7287) );
  AOI22_X1 U9033 ( .A1(n9116), .A2(n9465), .B1(n7287), .B2(n9092), .ZN(n7291)
         );
  NOR2_X1 U9034 ( .A1(n9170), .A2(n7469), .ZN(n7288) );
  AOI211_X1 U9035 ( .C1(n9167), .C2(n9467), .A(n7289), .B(n7288), .ZN(n7290)
         );
  OAI211_X1 U9036 ( .C1(n7292), .C2(n9144), .A(n7291), .B(n7290), .ZN(P1_U3237) );
  NAND2_X1 U9037 ( .A1(n7294), .A2(n7293), .ZN(n7296) );
  XOR2_X1 U9038 ( .A(n7296), .B(n7295), .Z(n7303) );
  OR2_X1 U9039 ( .A1(n8032), .A2(n8858), .ZN(n7298) );
  OR2_X1 U9040 ( .A1(n7561), .A2(n8856), .ZN(n7297) );
  NAND2_X1 U9041 ( .A1(n7298), .A2(n7297), .ZN(n10155) );
  NAND2_X1 U9042 ( .A1(n8241), .A2(n10155), .ZN(n7299) );
  OAI211_X1 U9043 ( .C1(n10152), .C2(n10158), .A(n7300), .B(n7299), .ZN(n7301)
         );
  AOI21_X1 U9044 ( .B1(n10136), .B2(n10162), .A(n7301), .ZN(n7302) );
  OAI21_X1 U9045 ( .B1(n7303), .B2(n10098), .A(n7302), .ZN(P2_U3226) );
  INV_X1 U9046 ( .A(n7304), .ZN(n7402) );
  OAI222_X1 U9047 ( .A1(P2_U3152), .A2(n8104), .B1(n9021), .B2(n7402), .C1(
        n7305), .C2(n9018), .ZN(P2_U3337) );
  OAI21_X1 U9048 ( .B1(n7307), .B2(n9304), .A(n7306), .ZN(n7308) );
  NAND2_X1 U9049 ( .A1(n7308), .A2(n10066), .ZN(n7316) );
  OAI21_X1 U9050 ( .B1(n7311), .B2(n7309), .A(n7310), .ZN(n7314) );
  OAI22_X1 U9051 ( .A1(n7389), .A2(n10062), .B1(n7312), .B2(n10015), .ZN(n7313) );
  AOI21_X1 U9052 ( .B1(n7314), .B2(n9637), .A(n7313), .ZN(n7315) );
  AND2_X1 U9053 ( .A1(n7316), .A2(n7315), .ZN(n10060) );
  OAI211_X1 U9054 ( .C1(n7318), .C2(n10057), .A(n10003), .B(n7317), .ZN(n10056) );
  OAI22_X1 U9055 ( .A1(n9629), .A2(n7319), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10008), .ZN(n7320) );
  AOI21_X1 U9056 ( .B1(n10028), .B2(n7321), .A(n7320), .ZN(n7322) );
  OAI21_X1 U9057 ( .B1(n9724), .B2(n10056), .A(n7322), .ZN(n7323) );
  INV_X1 U9058 ( .A(n7323), .ZN(n7324) );
  OAI21_X1 U9059 ( .B1(n10060), .B2(n10024), .A(n7324), .ZN(P1_U3288) );
  INV_X1 U9060 ( .A(n7325), .ZN(n7326) );
  AOI21_X1 U9061 ( .B1(n9309), .B2(n7327), .A(n7326), .ZN(n7445) );
  NAND2_X1 U9062 ( .A1(n9629), .A2(n9637), .ZN(n9730) );
  OAI21_X1 U9063 ( .B1(n7329), .B2(n9309), .A(n7328), .ZN(n7447) );
  NOR2_X1 U9064 ( .A1(n9450), .A2(n7330), .ZN(n7331) );
  NAND2_X1 U9065 ( .A1(n7447), .A2(n9714), .ZN(n7340) );
  OAI211_X1 U9066 ( .C1(n7333), .C2(n7462), .A(n10003), .B(n7332), .ZN(n7443)
         );
  INV_X1 U9067 ( .A(n7443), .ZN(n7338) );
  NAND2_X1 U9068 ( .A1(n9629), .A2(n9818), .ZN(n9720) );
  NAND2_X1 U9069 ( .A1(n9629), .A2(n9819), .ZN(n9631) );
  INV_X1 U9070 ( .A(n9631), .ZN(n9718) );
  OAI22_X1 U9071 ( .A1(n9629), .A2(n6771), .B1(n7458), .B2(n10008), .ZN(n7334)
         );
  AOI21_X1 U9072 ( .B1(n9718), .B2(n9466), .A(n7334), .ZN(n7336) );
  NAND2_X1 U9073 ( .A1(n10028), .A2(n7448), .ZN(n7335) );
  OAI211_X1 U9074 ( .C1(n10016), .C2(n9720), .A(n7336), .B(n7335), .ZN(n7337)
         );
  AOI21_X1 U9075 ( .B1(n7338), .B2(n10006), .A(n7337), .ZN(n7339) );
  OAI211_X1 U9076 ( .C1(n7445), .C2(n9730), .A(n7340), .B(n7339), .ZN(P1_U3284) );
  OR2_X1 U9077 ( .A1(n7341), .A2(n8336), .ZN(n7349) );
  INV_X1 U9078 ( .A(n7349), .ZN(n7342) );
  OR2_X1 U9079 ( .A1(n8150), .A2(n7342), .ZN(n7346) );
  OR2_X1 U9080 ( .A1(n7412), .A2(n7346), .ZN(n7344) );
  OR2_X1 U9081 ( .A1(n7342), .A2(n7348), .ZN(n7343) );
  NAND2_X1 U9082 ( .A1(n7344), .A2(n7343), .ZN(n7352) );
  INV_X1 U9083 ( .A(n8155), .ZN(n7347) );
  OR2_X1 U9084 ( .A1(n7346), .A2(n7347), .ZN(n7413) );
  OR2_X1 U9085 ( .A1(n7412), .A2(n7413), .ZN(n7409) );
  NAND2_X1 U9086 ( .A1(n7350), .A2(n7349), .ZN(n7407) );
  AND2_X1 U9087 ( .A1(n7409), .A2(n7407), .ZN(n7351) );
  OAI21_X1 U9088 ( .B1(n7352), .B2(n8155), .A(n7351), .ZN(n10240) );
  XOR2_X1 U9089 ( .A(n8155), .B(n7403), .Z(n7355) );
  OAI22_X1 U9090 ( .A1(n7561), .A2(n8858), .B1(n10129), .B2(n8856), .ZN(n7354)
         );
  AOI21_X1 U9091 ( .B1(n7355), .B2(n10156), .A(n7354), .ZN(n7356) );
  OAI21_X1 U9092 ( .B1(n10240), .B2(n7568), .A(n7356), .ZN(n10243) );
  NAND2_X1 U9093 ( .A1(n10243), .A2(n8881), .ZN(n7361) );
  OAI22_X1 U9094 ( .A1(n8881), .A2(n7357), .B1(n10104), .B2(n8888), .ZN(n7359)
         );
  XNOR2_X1 U9095 ( .A(n7416), .B(n7345), .ZN(n10242) );
  NOR2_X1 U9096 ( .A1(n8780), .A2(n10242), .ZN(n7358) );
  AOI211_X1 U9097 ( .C1(n10161), .C2(n7345), .A(n7359), .B(n7358), .ZN(n7360)
         );
  OAI211_X1 U9098 ( .C1(n10240), .C2(n7587), .A(n7361), .B(n7360), .ZN(
        P2_U3286) );
  XNOR2_X1 U9099 ( .A(n7362), .B(n7363), .ZN(n7367) );
  INV_X1 U9100 ( .A(n7711), .ZN(n8332) );
  AND2_X1 U9101 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7438) );
  OAI22_X1 U9102 ( .A1(n10095), .A2(n7576), .B1(n10152), .B2(n7581), .ZN(n7364) );
  AOI211_X1 U9103 ( .C1(n10138), .C2(n8332), .A(n7438), .B(n7364), .ZN(n7366)
         );
  NAND2_X1 U9104 ( .A1(n10136), .A2(n8033), .ZN(n7365) );
  OAI211_X1 U9105 ( .C1(n7367), .C2(n10098), .A(n7366), .B(n7365), .ZN(
        P2_U3236) );
  INV_X1 U9106 ( .A(n7368), .ZN(n7381) );
  OAI22_X1 U9107 ( .A1(n9629), .A2(n6582), .B1(n7369), .B2(n10008), .ZN(n7370)
         );
  AOI21_X1 U9108 ( .B1(n10028), .B2(n7371), .A(n7370), .ZN(n7376) );
  OAI22_X1 U9109 ( .A1(n7373), .A2(n9720), .B1(n9631), .B2(n7372), .ZN(n7374)
         );
  INV_X1 U9110 ( .A(n7374), .ZN(n7375) );
  OAI211_X1 U9111 ( .C1(n7377), .C2(n9724), .A(n7376), .B(n7375), .ZN(n7378)
         );
  AOI21_X1 U9112 ( .B1(n7379), .B2(n9714), .A(n7378), .ZN(n7380) );
  OAI21_X1 U9113 ( .B1(n7381), .B2(n10024), .A(n7380), .ZN(P1_U3287) );
  NAND2_X1 U9114 ( .A1(n7383), .A2(n7382), .ZN(n7386) );
  INV_X1 U9115 ( .A(n7384), .ZN(n7385) );
  AOI21_X1 U9116 ( .B1(n7388), .B2(n7386), .A(n7385), .ZN(n10067) );
  AOI22_X1 U9117 ( .A1(n10028), .A2(n7394), .B1(n10024), .B2(
        P1_REG2_REG_5__SCAN_IN), .ZN(n7387) );
  OAI21_X1 U9118 ( .B1(n10063), .B2(n9720), .A(n7387), .ZN(n7399) );
  XNOR2_X1 U9119 ( .A(n7234), .B(n7388), .ZN(n7391) );
  NOR2_X1 U9120 ( .A1(n7389), .A2(n10015), .ZN(n7390) );
  AOI21_X1 U9121 ( .B1(n7391), .B2(n9637), .A(n7390), .ZN(n10068) );
  AOI211_X1 U9122 ( .C1(n7394), .C2(n7393), .A(n9695), .B(n7392), .ZN(n10065)
         );
  INV_X1 U9123 ( .A(n7395), .ZN(n7396) );
  AOI22_X1 U9124 ( .A1(n10065), .A2(n4390), .B1(n10035), .B2(n7396), .ZN(n7397) );
  AOI21_X1 U9125 ( .B1(n10068), .B2(n7397), .A(n10024), .ZN(n7398) );
  AOI211_X1 U9126 ( .C1(n9714), .C2(n10067), .A(n7399), .B(n7398), .ZN(n7400)
         );
  INV_X1 U9127 ( .A(n7400), .ZN(P1_U3286) );
  OAI222_X1 U9128 ( .A1(n9878), .A2(n7402), .B1(P1_U3084), .B2(n9398), .C1(
        n7401), .C2(n9874), .ZN(P1_U3332) );
  NAND2_X1 U9129 ( .A1(n7562), .A2(n7561), .ZN(n8020) );
  XNOR2_X1 U9130 ( .A(n7570), .B(n7569), .ZN(n7404) );
  OAI222_X1 U9131 ( .A1(n8858), .A2(n7576), .B1(n8856), .B2(n7405), .C1(n8854), 
        .C2(n7404), .ZN(n10250) );
  INV_X1 U9132 ( .A(n10250), .ZN(n7425) );
  INV_X1 U9133 ( .A(n7405), .ZN(n8335) );
  NAND2_X1 U9134 ( .A1(n7345), .A2(n8335), .ZN(n7406) );
  NAND2_X1 U9135 ( .A1(n7409), .A2(n7408), .ZN(n7410) );
  OR2_X1 U9136 ( .A1(n7410), .A2(n8156), .ZN(n7415) );
  NAND2_X1 U9137 ( .A1(n8156), .A2(n7411), .ZN(n7563) );
  INV_X1 U9138 ( .A(n7412), .ZN(n7414) );
  NAND2_X1 U9139 ( .A1(n7414), .A2(n4909), .ZN(n7566) );
  AND2_X1 U9140 ( .A1(n7563), .A2(n7566), .ZN(n10164) );
  AND2_X1 U9141 ( .A1(n7415), .A2(n10164), .ZN(n10252) );
  AND2_X1 U9142 ( .A1(n7417), .A2(n10247), .ZN(n10169) );
  NOR2_X1 U9143 ( .A1(n7417), .A2(n10247), .ZN(n7418) );
  OR2_X1 U9144 ( .A1(n10169), .A2(n7418), .ZN(n10249) );
  OAI22_X1 U9145 ( .A1(n8881), .A2(n7420), .B1(n7419), .B2(n8888), .ZN(n7421)
         );
  AOI21_X1 U9146 ( .B1(n10161), .B2(n7562), .A(n7421), .ZN(n7422) );
  OAI21_X1 U9147 ( .B1(n10249), .B2(n8780), .A(n7422), .ZN(n7423) );
  AOI21_X1 U9148 ( .B1(n10252), .B2(n10172), .A(n7423), .ZN(n7424) );
  OAI21_X1 U9149 ( .B1(n7425), .B2(n4392), .A(n7424), .ZN(P2_U3285) );
  INV_X1 U9150 ( .A(n7426), .ZN(n7934) );
  OAI222_X1 U9151 ( .A1(n9874), .A2(n7427), .B1(n9878), .B2(n7934), .C1(n9405), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  NAND2_X1 U9152 ( .A1(n7429), .A2(n7428), .ZN(n7431) );
  AOI22_X1 U9153 ( .A1(n7512), .A2(n7582), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7506), .ZN(n7430) );
  NOR2_X1 U9154 ( .A1(n7431), .A2(n7430), .ZN(n7505) );
  AOI21_X1 U9155 ( .B1(n7431), .B2(n7430), .A(n7505), .ZN(n7442) );
  OAI21_X1 U9156 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n7433), .A(n7432), .ZN(
        n7435) );
  AOI22_X1 U9157 ( .A1(n7512), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n7614), .B2(
        n7506), .ZN(n7434) );
  NAND2_X1 U9158 ( .A1(n7434), .A2(n7435), .ZN(n7511) );
  OAI21_X1 U9159 ( .B1(n7435), .B2(n7434), .A(n7511), .ZN(n7439) );
  INV_X1 U9160 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7436) );
  NOR2_X1 U9161 ( .A1(n8389), .A2(n7436), .ZN(n7437) );
  AOI211_X1 U9162 ( .C1(n8381), .C2(n7439), .A(n7438), .B(n7437), .ZN(n7441)
         );
  INV_X1 U9163 ( .A(n8376), .ZN(n7518) );
  NAND2_X1 U9164 ( .A1(n7518), .A2(n7512), .ZN(n7440) );
  OAI211_X1 U9165 ( .C1(n7442), .C2(n8368), .A(n7441), .B(n7440), .ZN(P2_U3258) );
  AOI22_X1 U9166 ( .A1(n9818), .A2(n9464), .B1(n9466), .B2(n9819), .ZN(n7444)
         );
  OAI211_X1 U9167 ( .C1(n7445), .C2(n10020), .A(n7444), .B(n7443), .ZN(n7446)
         );
  AOI21_X1 U9168 ( .B1(n10066), .B2(n7447), .A(n7446), .ZN(n7452) );
  AOI22_X1 U9169 ( .A1(n7604), .A2(n7448), .B1(n10081), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7449) );
  OAI21_X1 U9170 ( .B1(n7452), .B2(n10081), .A(n7449), .ZN(P1_U3530) );
  OAI22_X1 U9171 ( .A1(n9864), .A2(n7462), .B1(n10076), .B2(n5068), .ZN(n7450)
         );
  INV_X1 U9172 ( .A(n7450), .ZN(n7451) );
  OAI21_X1 U9173 ( .B1(n7452), .B2(n10075), .A(n7451), .ZN(P1_U3475) );
  NAND2_X1 U9174 ( .A1(n7455), .A2(n7454), .ZN(n7456) );
  XNOR2_X1 U9175 ( .A(n7453), .B(n7456), .ZN(n7457) );
  NAND2_X1 U9176 ( .A1(n7457), .A2(n9160), .ZN(n7461) );
  AND2_X1 U9177 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9932) );
  OAI22_X1 U9178 ( .A1(n9164), .A2(n7458), .B1(n9162), .B2(n10016), .ZN(n7459)
         );
  AOI211_X1 U9179 ( .C1(n9167), .C2(n9466), .A(n9932), .B(n7459), .ZN(n7460)
         );
  OAI211_X1 U9180 ( .C1(n7462), .C2(n9170), .A(n7461), .B(n7460), .ZN(P1_U3211) );
  NAND2_X1 U9181 ( .A1(n7463), .A2(n10006), .ZN(n7468) );
  OAI22_X1 U9182 ( .A1(n9629), .A2(n6775), .B1(n7464), .B2(n10008), .ZN(n7466)
         );
  NOR2_X1 U9183 ( .A1(n9720), .A2(n7483), .ZN(n7465) );
  AOI211_X1 U9184 ( .C1(n9718), .C2(n9467), .A(n7466), .B(n7465), .ZN(n7467)
         );
  OAI211_X1 U9185 ( .C1(n7469), .C2(n9623), .A(n7468), .B(n7467), .ZN(n7470)
         );
  AOI21_X1 U9186 ( .B1(n7471), .B2(n9714), .A(n7470), .ZN(n7472) );
  OAI21_X1 U9187 ( .B1(n10024), .B2(n7473), .A(n7472), .ZN(P1_U3285) );
  XNOR2_X1 U9188 ( .A(n7474), .B(n9311), .ZN(n7475) );
  NAND2_X1 U9189 ( .A1(n7475), .A2(n9637), .ZN(n7490) );
  INV_X1 U9190 ( .A(n7476), .ZN(n7477) );
  AOI21_X1 U9191 ( .B1(n9311), .B2(n7478), .A(n7477), .ZN(n7492) );
  NAND2_X1 U9192 ( .A1(n7492), .A2(n9714), .ZN(n7487) );
  AOI21_X1 U9193 ( .B1(n7332), .B2(n7496), .A(n9695), .ZN(n7479) );
  NAND2_X1 U9194 ( .A1(n7479), .A2(n10002), .ZN(n7488) );
  INV_X1 U9195 ( .A(n7488), .ZN(n7485) );
  INV_X1 U9196 ( .A(n9720), .ZN(n7744) );
  OAI22_X1 U9197 ( .A1(n9629), .A2(n5085), .B1(n7640), .B2(n10008), .ZN(n7480)
         );
  AOI21_X1 U9198 ( .B1(n7744), .B2(n9463), .A(n7480), .ZN(n7482) );
  NAND2_X1 U9199 ( .A1(n10028), .A2(n7496), .ZN(n7481) );
  OAI211_X1 U9200 ( .C1(n7483), .C2(n9631), .A(n7482), .B(n7481), .ZN(n7484)
         );
  AOI21_X1 U9201 ( .B1(n7485), .B2(n10006), .A(n7484), .ZN(n7486) );
  OAI211_X1 U9202 ( .C1(n10024), .C2(n7490), .A(n7487), .B(n7486), .ZN(
        P1_U3283) );
  AOI22_X1 U9203 ( .A1(n9465), .A2(n9819), .B1(n9818), .B2(n9463), .ZN(n7489)
         );
  NAND3_X1 U9204 ( .A1(n7490), .A2(n7489), .A3(n7488), .ZN(n7491) );
  AOI21_X1 U9205 ( .B1(n7492), .B2(n10066), .A(n7491), .ZN(n7498) );
  INV_X1 U9206 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7493) );
  OAI22_X1 U9207 ( .A1(n9864), .A2(n7644), .B1(n10076), .B2(n7493), .ZN(n7494)
         );
  INV_X1 U9208 ( .A(n7494), .ZN(n7495) );
  OAI21_X1 U9209 ( .B1(n7498), .B2(n10075), .A(n7495), .ZN(P1_U3478) );
  AOI22_X1 U9210 ( .A1(n7604), .A2(n7496), .B1(n10081), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n7497) );
  OAI21_X1 U9211 ( .B1(n7498), .B2(n10081), .A(n7497), .ZN(P1_U3531) );
  NAND2_X1 U9212 ( .A1(n7502), .A2(n7907), .ZN(n7500) );
  NAND2_X1 U9213 ( .A1(n7499), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9454) );
  OAI211_X1 U9214 ( .C1(n7501), .C2(n9874), .A(n7500), .B(n9454), .ZN(P1_U3330) );
  NAND2_X1 U9215 ( .A1(n7502), .A2(n9016), .ZN(n7503) );
  OAI211_X1 U9216 ( .C1(n7504), .C2(n9018), .A(n7503), .B(n8182), .ZN(P2_U3335) );
  AOI21_X1 U9217 ( .B1(n7506), .B2(n7582), .A(n7505), .ZN(n7508) );
  AOI22_X1 U9218 ( .A1(n7829), .A2(n6152), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7509), .ZN(n7507) );
  NOR2_X1 U9219 ( .A1(n7508), .A2(n7507), .ZN(n7830) );
  AOI21_X1 U9220 ( .B1(n7508), .B2(n7507), .A(n7830), .ZN(n7521) );
  AOI22_X1 U9221 ( .A1(n7829), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n7510), .B2(
        n7509), .ZN(n7514) );
  OAI21_X1 U9222 ( .B1(n7514), .B2(n7513), .A(n7826), .ZN(n7515) );
  NAND2_X1 U9223 ( .A1(n7515), .A2(n8381), .ZN(n7520) );
  INV_X1 U9224 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7516) );
  NAND2_X1 U9225 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7556) );
  OAI21_X1 U9226 ( .B1(n8389), .B2(n7516), .A(n7556), .ZN(n7517) );
  AOI21_X1 U9227 ( .B1(n7518), .B2(n7829), .A(n7517), .ZN(n7519) );
  OAI211_X1 U9228 ( .C1(n7521), .C2(n8368), .A(n7520), .B(n7519), .ZN(P2_U3259) );
  NAND2_X1 U9229 ( .A1(n7522), .A2(n9307), .ZN(n7524) );
  INV_X1 U9230 ( .A(n9313), .ZN(n7523) );
  XNOR2_X1 U9231 ( .A(n7524), .B(n7523), .ZN(n7525) );
  NAND2_X1 U9232 ( .A1(n7525), .A2(n9637), .ZN(n7598) );
  OAI21_X1 U9233 ( .B1(n7527), .B2(n9313), .A(n7526), .ZN(n7600) );
  NAND2_X1 U9234 ( .A1(n7600), .A2(n9714), .ZN(n7536) );
  OAI21_X1 U9235 ( .B1(n4462), .B2(n7686), .A(n10003), .ZN(n7528) );
  OR2_X1 U9236 ( .A1(n7528), .A2(n7663), .ZN(n7596) );
  INV_X1 U9237 ( .A(n7596), .ZN(n7534) );
  INV_X1 U9238 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7529) );
  OAI22_X1 U9239 ( .A1(n9629), .A2(n7529), .B1(n7681), .B2(n10008), .ZN(n7530)
         );
  AOI21_X1 U9240 ( .B1(n7744), .B2(n9461), .A(n7530), .ZN(n7532) );
  NAND2_X1 U9241 ( .A1(n10028), .A2(n7603), .ZN(n7531) );
  OAI211_X1 U9242 ( .C1(n7639), .C2(n9631), .A(n7532), .B(n7531), .ZN(n7533)
         );
  AOI21_X1 U9243 ( .B1(n7534), .B2(n10006), .A(n7533), .ZN(n7535) );
  OAI211_X1 U9244 ( .C1(n10024), .C2(n7598), .A(n7536), .B(n7535), .ZN(
        P1_U3281) );
  INV_X1 U9245 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7550) );
  MUX2_X1 U9246 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n7537), .S(n7653), .Z(n7540)
         );
  OAI21_X1 U9247 ( .B1(n7544), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7538), .ZN(
        n7539) );
  NAND2_X1 U9248 ( .A1(n7540), .A2(n7539), .ZN(n7652) );
  OAI21_X1 U9249 ( .B1(n7540), .B2(n7539), .A(n7652), .ZN(n7548) );
  NOR2_X1 U9250 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7541), .ZN(n9029) );
  INV_X1 U9251 ( .A(n9029), .ZN(n7542) );
  OAI21_X1 U9252 ( .B1(n9491), .B2(n7645), .A(n7542), .ZN(n7547) );
  NOR2_X1 U9253 ( .A1(n7763), .A2(n7545), .ZN(n7647) );
  AOI211_X1 U9254 ( .C1(n7545), .C2(n7763), .A(n7647), .B(n9986), .ZN(n7546)
         );
  AOI211_X1 U9255 ( .C1(n9998), .C2(n7548), .A(n7547), .B(n7546), .ZN(n7549)
         );
  OAI21_X1 U9256 ( .B1(n9984), .B2(n7550), .A(n7549), .ZN(P1_U3255) );
  INV_X1 U9257 ( .A(n7551), .ZN(n7552) );
  AOI21_X1 U9258 ( .B1(n7554), .B2(n7553), .A(n7552), .ZN(n7560) );
  INV_X1 U9259 ( .A(n7555), .ZN(n7718) );
  INV_X1 U9260 ( .A(n8032), .ZN(n8333) );
  AOI22_X1 U9261 ( .A1(n7718), .A2(n8303), .B1(n10140), .B2(n8333), .ZN(n7557)
         );
  OAI211_X1 U9262 ( .C1(n7800), .C2(n10130), .A(n7557), .B(n7556), .ZN(n7558)
         );
  AOI21_X1 U9263 ( .B1(n10136), .B2(n8989), .A(n7558), .ZN(n7559) );
  OAI21_X1 U9264 ( .B1(n7560), .B2(n10098), .A(n7559), .ZN(P2_U3217) );
  INV_X1 U9265 ( .A(n7561), .ZN(n10093) );
  NAND2_X1 U9266 ( .A1(n7562), .A2(n10093), .ZN(n10163) );
  AND2_X1 U9267 ( .A1(n10163), .A2(n7563), .ZN(n7564) );
  OR2_X1 U9268 ( .A1(n10162), .A2(n7576), .ZN(n8024) );
  INV_X1 U9269 ( .A(n10154), .ZN(n10166) );
  AOI21_X2 U9270 ( .B1(n7566), .B2(n7565), .A(n4409), .ZN(n7567) );
  XNOR2_X1 U9271 ( .A(n8033), .B(n8032), .ZN(n7969) );
  NAND2_X1 U9272 ( .A1(n7567), .A2(n7969), .ZN(n7713) );
  OAI21_X1 U9273 ( .B1(n7567), .B2(n7969), .A(n7713), .ZN(n7609) );
  OR2_X1 U9274 ( .A1(n7609), .A2(n7568), .ZN(n7580) );
  NAND2_X1 U9275 ( .A1(n7570), .A2(n7569), .ZN(n7571) );
  NAND2_X1 U9276 ( .A1(n7571), .A2(n8022), .ZN(n10153) );
  NAND2_X1 U9277 ( .A1(n10153), .A2(n10154), .ZN(n7572) );
  NAND2_X1 U9278 ( .A1(n7572), .A2(n8024), .ZN(n7574) );
  NAND2_X1 U9279 ( .A1(n7574), .A2(n7969), .ZN(n7575) );
  NAND2_X1 U9280 ( .A1(n7723), .A2(n7575), .ZN(n7578) );
  OAI22_X1 U9281 ( .A1(n7711), .A2(n8858), .B1(n7576), .B2(n8856), .ZN(n7577)
         );
  AOI21_X1 U9282 ( .B1(n7578), .B2(n10156), .A(n7577), .ZN(n7579) );
  NAND2_X1 U9283 ( .A1(n7580), .A2(n7579), .ZN(n7611) );
  OAI22_X1 U9284 ( .A1(n8881), .A2(n7582), .B1(n7581), .B2(n8888), .ZN(n7583)
         );
  AOI21_X1 U9285 ( .B1(n8033), .B2(n10161), .A(n7583), .ZN(n7586) );
  INV_X1 U9286 ( .A(n10162), .ZN(n10256) );
  NAND2_X1 U9287 ( .A1(n10169), .A2(n10256), .ZN(n10168) );
  NAND2_X1 U9288 ( .A1(n10168), .A2(n8033), .ZN(n7584) );
  AND2_X1 U9289 ( .A1(n4406), .A2(n7584), .ZN(n7607) );
  NAND2_X1 U9290 ( .A1(n7607), .A2(n6504), .ZN(n7585) );
  OAI211_X1 U9291 ( .C1(n7609), .C2(n7587), .A(n7586), .B(n7585), .ZN(n7588)
         );
  AOI21_X1 U9292 ( .B1(n8881), .B2(n7611), .A(n7588), .ZN(n7589) );
  INV_X1 U9293 ( .A(n7589), .ZN(P2_U3283) );
  INV_X1 U9294 ( .A(n5909), .ZN(n7594) );
  OAI222_X1 U9295 ( .A1(n9878), .A2(n7594), .B1(P1_U3084), .B2(n7591), .C1(
        n7590), .C2(n9874), .ZN(P1_U3329) );
  INV_X1 U9296 ( .A(n7592), .ZN(n7595) );
  OAI222_X1 U9297 ( .A1(P2_U3152), .A2(n7595), .B1(n9021), .B2(n7594), .C1(
        n7593), .C2(n9018), .ZN(P2_U3334) );
  AOI22_X1 U9298 ( .A1(n9461), .A2(n9818), .B1(n9819), .B2(n9463), .ZN(n7597)
         );
  NAND3_X1 U9299 ( .A1(n7598), .A2(n7597), .A3(n7596), .ZN(n7599) );
  AOI21_X1 U9300 ( .B1(n7600), .B2(n10066), .A(n7599), .ZN(n7606) );
  OAI22_X1 U9301 ( .A1(n7686), .A2(n9864), .B1(n10076), .B2(n5137), .ZN(n7601)
         );
  INV_X1 U9302 ( .A(n7601), .ZN(n7602) );
  OAI21_X1 U9303 ( .B1(n7606), .B2(n10075), .A(n7602), .ZN(P1_U3484) );
  AOI22_X1 U9304 ( .A1(n7604), .A2(n7603), .B1(n10081), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7605) );
  OAI21_X1 U9305 ( .B1(n7606), .B2(n10081), .A(n7605), .ZN(P1_U3533) );
  AOI22_X1 U9306 ( .A1(n7607), .A2(n10215), .B1(n8033), .B2(n10213), .ZN(n7608) );
  OAI21_X1 U9307 ( .B1(n7609), .B2(n10228), .A(n7608), .ZN(n7610) );
  NOR2_X1 U9308 ( .A1(n7611), .A2(n7610), .ZN(n7615) );
  INV_X1 U9309 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7612) );
  MUX2_X1 U9310 ( .A(n7615), .B(n7612), .S(n10260), .Z(n7613) );
  INV_X1 U9311 ( .A(n7613), .ZN(P2_U3490) );
  MUX2_X1 U9312 ( .A(n7615), .B(n7614), .S(n10273), .Z(n7616) );
  INV_X1 U9313 ( .A(n7616), .ZN(P2_U3533) );
  OAI21_X1 U9314 ( .B1(n7619), .B2(n7618), .A(n7617), .ZN(n7620) );
  NAND2_X1 U9315 ( .A1(n7620), .A2(n9160), .ZN(n7624) );
  OAI22_X1 U9316 ( .A1(n9164), .A2(n10009), .B1(n9162), .B2(n10017), .ZN(n7621) );
  AOI211_X1 U9317 ( .C1(n9167), .C2(n9464), .A(n7622), .B(n7621), .ZN(n7623)
         );
  OAI211_X1 U9318 ( .C1(n4629), .C2(n9170), .A(n7624), .B(n7623), .ZN(P1_U3229) );
  XNOR2_X1 U9319 ( .A(n7626), .B(n7625), .ZN(n7630) );
  OAI22_X1 U9320 ( .A1(n10130), .A2(n8859), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8652), .ZN(n7628) );
  OAI22_X1 U9321 ( .A1(n10095), .A2(n8857), .B1(n10152), .B2(n8867), .ZN(n7627) );
  AOI211_X1 U9322 ( .C1(n8975), .C2(n10136), .A(n7628), .B(n7627), .ZN(n7629)
         );
  OAI21_X1 U9323 ( .B1(n7630), .B2(n10098), .A(n7629), .ZN(P2_U3230) );
  INV_X1 U9324 ( .A(n7631), .ZN(n7633) );
  NOR2_X1 U9325 ( .A1(n7633), .A2(n7632), .ZN(n7637) );
  AOI21_X1 U9326 ( .B1(n7631), .B2(n7635), .A(n7634), .ZN(n7636) );
  OAI21_X1 U9327 ( .B1(n7637), .B2(n7636), .A(n9160), .ZN(n7643) );
  NOR2_X1 U9328 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7638), .ZN(n9945) );
  OAI22_X1 U9329 ( .A1(n9164), .A2(n7640), .B1(n9162), .B2(n7639), .ZN(n7641)
         );
  AOI211_X1 U9330 ( .C1(n9167), .C2(n9465), .A(n9945), .B(n7641), .ZN(n7642)
         );
  OAI211_X1 U9331 ( .C1(n7644), .C2(n9170), .A(n7643), .B(n7642), .ZN(P1_U3219) );
  NOR2_X1 U9332 ( .A1(n7646), .A2(n7645), .ZN(n7648) );
  NOR2_X1 U9333 ( .A1(n7648), .A2(n7647), .ZN(n7935) );
  INV_X1 U9334 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7649) );
  AOI211_X1 U9335 ( .C1(n7650), .C2(n7649), .A(n7936), .B(n9986), .ZN(n7660)
         );
  INV_X1 U9336 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7658) );
  INV_X1 U9337 ( .A(n7942), .ZN(n7651) );
  AND2_X1 U9338 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9166) );
  AOI21_X1 U9339 ( .B1(n9992), .B2(n7651), .A(n9166), .ZN(n7657) );
  OAI21_X1 U9340 ( .B1(n7653), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7652), .ZN(
        n7941) );
  XNOR2_X1 U9341 ( .A(n7942), .B(n7941), .ZN(n7654) );
  AND2_X1 U9342 ( .A1(n7654), .A2(n7931), .ZN(n7655) );
  NOR2_X1 U9343 ( .A1(n7931), .A2(n7654), .ZN(n7943) );
  OR3_X1 U9344 ( .A1(n9492), .A2(n7655), .A3(n7943), .ZN(n7656) );
  OAI211_X1 U9345 ( .C1(n9984), .C2(n7658), .A(n7657), .B(n7656), .ZN(n7659)
         );
  OR2_X1 U9346 ( .A1(n7660), .A2(n7659), .ZN(P1_U3256) );
  OAI22_X1 U9347 ( .A1(n9629), .A2(n7661), .B1(n7792), .B2(n10008), .ZN(n7665)
         );
  OAI211_X1 U9348 ( .C1(n7663), .C2(n9912), .A(n10003), .B(n7662), .ZN(n9911)
         );
  NOR2_X1 U9349 ( .A1(n9911), .A2(n9724), .ZN(n7664) );
  AOI211_X1 U9350 ( .C1(n10028), .C2(n7794), .A(n7665), .B(n7664), .ZN(n7675)
         );
  NAND2_X1 U9351 ( .A1(n7666), .A2(n9314), .ZN(n7740) );
  OR2_X1 U9352 ( .A1(n7666), .A2(n9314), .ZN(n7667) );
  NAND2_X1 U9353 ( .A1(n7740), .A2(n7667), .ZN(n7673) );
  XNOR2_X1 U9354 ( .A(n7668), .B(n9314), .ZN(n7670) );
  OAI22_X1 U9355 ( .A1(n9113), .A2(n10062), .B1(n10017), .B2(n10015), .ZN(
        n7669) );
  AOI21_X1 U9356 ( .B1(n7670), .B2(n9637), .A(n7669), .ZN(n7671) );
  OAI21_X1 U9357 ( .B1(n7673), .B2(n7672), .A(n7671), .ZN(n9913) );
  NAND2_X1 U9358 ( .A1(n9913), .A2(n9629), .ZN(n7674) );
  NAND2_X1 U9359 ( .A1(n7675), .A2(n7674), .ZN(P1_U3280) );
  XNOR2_X1 U9360 ( .A(n7677), .B(n7676), .ZN(n7678) );
  XNOR2_X1 U9361 ( .A(n7679), .B(n7678), .ZN(n7680) );
  NAND2_X1 U9362 ( .A1(n7680), .A2(n9160), .ZN(n7685) );
  OAI22_X1 U9363 ( .A1(n9164), .A2(n7681), .B1(n9162), .B2(n7746), .ZN(n7682)
         );
  AOI211_X1 U9364 ( .C1(n9167), .C2(n9463), .A(n7683), .B(n7682), .ZN(n7684)
         );
  OAI211_X1 U9365 ( .C1(n7686), .C2(n9170), .A(n7685), .B(n7684), .ZN(P1_U3215) );
  INV_X1 U9366 ( .A(n8984), .ZN(n7877) );
  NAND2_X1 U9367 ( .A1(n10145), .A2(n7779), .ZN(n7689) );
  INV_X1 U9368 ( .A(n8315), .ZN(n10118) );
  INV_X1 U9369 ( .A(n7800), .ZN(n8331) );
  NAND2_X1 U9370 ( .A1(n10118), .A2(n8331), .ZN(n7688) );
  XNOR2_X1 U9371 ( .A(n7687), .B(n7778), .ZN(n7780) );
  MUX2_X1 U9372 ( .A(n7689), .B(n7688), .S(n7780), .Z(n7693) );
  INV_X1 U9373 ( .A(n8857), .ZN(n8330) );
  NOR2_X1 U9374 ( .A1(n10152), .A2(n7874), .ZN(n7691) );
  OAI22_X1 U9375 ( .A1(n10095), .A2(n7711), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6179), .ZN(n7690) );
  AOI211_X1 U9376 ( .C1(n10138), .C2(n8330), .A(n7691), .B(n7690), .ZN(n7692)
         );
  OAI211_X1 U9377 ( .C1(n7877), .C2(n8327), .A(n7693), .B(n7692), .ZN(P2_U3243) );
  NAND2_X1 U9378 ( .A1(n7740), .A2(n7694), .ZN(n7696) );
  AND2_X1 U9379 ( .A1(n7696), .A2(n7695), .ZN(n7697) );
  XNOR2_X1 U9380 ( .A(n7697), .B(n9318), .ZN(n9826) );
  INV_X1 U9381 ( .A(n9826), .ZN(n7710) );
  OAI21_X1 U9382 ( .B1(n9318), .B2(n7699), .A(n7698), .ZN(n7700) );
  AND2_X1 U9383 ( .A1(n7700), .A2(n9637), .ZN(n9825) );
  AOI21_X1 U9384 ( .B1(n7747), .B2(n9816), .A(n9695), .ZN(n7701) );
  NAND2_X1 U9385 ( .A1(n7701), .A2(n7762), .ZN(n9822) );
  OAI22_X1 U9386 ( .A1(n9629), .A2(n7702), .B1(n9112), .B2(n10008), .ZN(n7705)
         );
  NOR2_X1 U9387 ( .A1(n9720), .A2(n7703), .ZN(n7704) );
  AOI211_X1 U9388 ( .C1(n9718), .C2(n9820), .A(n7705), .B(n7704), .ZN(n7707)
         );
  NAND2_X1 U9389 ( .A1(n9816), .A2(n10028), .ZN(n7706) );
  OAI211_X1 U9390 ( .C1(n9822), .C2(n9724), .A(n7707), .B(n7706), .ZN(n7708)
         );
  AOI21_X1 U9391 ( .B1(n9825), .B2(n9629), .A(n7708), .ZN(n7709) );
  OAI21_X1 U9392 ( .B1(n7710), .B2(n9706), .A(n7709), .ZN(P1_U3278) );
  NAND2_X1 U9393 ( .A1(n8989), .A2(n7711), .ZN(n8031) );
  NAND2_X1 U9394 ( .A1(n8033), .A2(n8333), .ZN(n7712) );
  INV_X1 U9395 ( .A(n7799), .ZN(n7715) );
  AOI21_X1 U9396 ( .B1(n8037), .B2(n7716), .A(n7715), .ZN(n8994) );
  AOI21_X1 U9397 ( .B1(n8989), .B2(n4406), .A(n4558), .ZN(n8990) );
  AOI22_X1 U9398 ( .A1(n4392), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7718), .B2(
        n10159), .ZN(n7719) );
  OAI21_X1 U9399 ( .B1(n7717), .B2(n8869), .A(n7719), .ZN(n7728) );
  INV_X1 U9400 ( .A(n7723), .ZN(n7720) );
  AND2_X1 U9401 ( .A1(n8033), .A2(n8032), .ZN(n7721) );
  OAI21_X1 U9402 ( .B1(n7720), .B2(n7721), .A(n7714), .ZN(n7724) );
  NOR2_X1 U9403 ( .A1(n7714), .A2(n7721), .ZN(n7722) );
  AND3_X1 U9404 ( .A1(n7724), .A2(n7804), .A3(n10156), .ZN(n7726) );
  OAI22_X1 U9405 ( .A1(n7800), .A2(n8858), .B1(n8032), .B2(n8856), .ZN(n7725)
         );
  NOR2_X1 U9406 ( .A1(n7726), .A2(n7725), .ZN(n8992) );
  NOR2_X1 U9407 ( .A1(n8992), .A2(n4392), .ZN(n7727) );
  AOI211_X1 U9408 ( .C1(n8990), .C2(n6504), .A(n7728), .B(n7727), .ZN(n7729)
         );
  OAI21_X1 U9409 ( .B1(n8994), .B2(n8874), .A(n7729), .ZN(P2_U3282) );
  INV_X1 U9410 ( .A(n7730), .ZN(n7734) );
  OAI222_X1 U9411 ( .A1(n7732), .A2(P2_U3152), .B1(n9021), .B2(n7734), .C1(
        n7731), .C2(n9018), .ZN(P2_U3333) );
  OAI222_X1 U9412 ( .A1(n9874), .A2(n8552), .B1(n9878), .B2(n7734), .C1(n7733), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  NAND2_X1 U9413 ( .A1(n7736), .A2(n7735), .ZN(n7737) );
  XNOR2_X1 U9414 ( .A(n7737), .B(n9315), .ZN(n7738) );
  NAND2_X1 U9415 ( .A1(n7738), .A2(n9637), .ZN(n7864) );
  NAND2_X1 U9416 ( .A1(n7740), .A2(n7739), .ZN(n7741) );
  XOR2_X1 U9417 ( .A(n9315), .B(n7741), .Z(n7866) );
  NAND2_X1 U9418 ( .A1(n7866), .A2(n9714), .ZN(n7752) );
  INV_X1 U9419 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7742) );
  OAI22_X1 U9420 ( .A1(n9629), .A2(n7742), .B1(n9056), .B2(n10008), .ZN(n7743)
         );
  AOI21_X1 U9421 ( .B1(n7744), .B2(n9460), .A(n7743), .ZN(n7745) );
  OAI21_X1 U9422 ( .B1(n7746), .B2(n9631), .A(n7745), .ZN(n7750) );
  AOI21_X1 U9423 ( .B1(n7662), .B2(n9058), .A(n9695), .ZN(n7748) );
  NAND2_X1 U9424 ( .A1(n7748), .A2(n7747), .ZN(n7862) );
  NOR2_X1 U9425 ( .A1(n7862), .A2(n9724), .ZN(n7749) );
  AOI211_X1 U9426 ( .C1(n10028), .C2(n9058), .A(n7750), .B(n7749), .ZN(n7751)
         );
  OAI211_X1 U9427 ( .C1(n10024), .C2(n7864), .A(n7752), .B(n7751), .ZN(
        P1_U3279) );
  NAND2_X1 U9428 ( .A1(n7753), .A2(n9637), .ZN(n7756) );
  INV_X1 U9429 ( .A(n7760), .ZN(n9319) );
  AOI21_X1 U9430 ( .B1(n7698), .B2(n9343), .A(n9319), .ZN(n7755) );
  AOI22_X1 U9431 ( .A1(n9807), .A2(n9818), .B1(n9819), .B2(n9460), .ZN(n7754)
         );
  OAI21_X1 U9432 ( .B1(n7756), .B2(n7755), .A(n7754), .ZN(n7915) );
  INV_X1 U9433 ( .A(n7915), .ZN(n7768) );
  NAND2_X1 U9434 ( .A1(n7666), .A2(n7757), .ZN(n7759) );
  AND2_X1 U9435 ( .A1(n7759), .A2(n7758), .ZN(n7761) );
  XNOR2_X1 U9436 ( .A(n7761), .B(n7760), .ZN(n7917) );
  NAND2_X1 U9437 ( .A1(n7917), .A2(n9714), .ZN(n7767) );
  AOI211_X1 U9438 ( .C1(n9030), .C2(n7762), .A(n9695), .B(n7843), .ZN(n7916)
         );
  INV_X1 U9439 ( .A(n9030), .ZN(n7922) );
  NOR2_X1 U9440 ( .A1(n7922), .A2(n9623), .ZN(n7765) );
  OAI22_X1 U9441 ( .A1(n9629), .A2(n7763), .B1(n9027), .B2(n10008), .ZN(n7764)
         );
  AOI211_X1 U9442 ( .C1(n7916), .C2(n10006), .A(n7765), .B(n7764), .ZN(n7766)
         );
  OAI211_X1 U9443 ( .C1(n10024), .C2(n7768), .A(n7767), .B(n7766), .ZN(
        P1_U3277) );
  XNOR2_X1 U9444 ( .A(n7769), .B(n7770), .ZN(n7775) );
  INV_X1 U9445 ( .A(n7771), .ZN(n8836) );
  INV_X1 U9446 ( .A(n7963), .ZN(n8841) );
  AOI22_X1 U9447 ( .A1(n8836), .A2(n8303), .B1(n10140), .B2(n8841), .ZN(n7772)
         );
  NAND2_X1 U9448 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8363) );
  OAI211_X1 U9449 ( .C1(n8293), .C2(n10130), .A(n7772), .B(n8363), .ZN(n7773)
         );
  AOI21_X1 U9450 ( .B1(n8969), .B2(n10136), .A(n7773), .ZN(n7774) );
  OAI21_X1 U9451 ( .B1(n7775), .B2(n10098), .A(n7774), .ZN(P2_U3240) );
  NAND2_X1 U9452 ( .A1(n7777), .A2(n7776), .ZN(n7782) );
  OAI22_X1 U9453 ( .A1(n7780), .A2(n7779), .B1(n7778), .B2(n7687), .ZN(n7781)
         );
  XOR2_X1 U9454 ( .A(n7782), .B(n7781), .Z(n7786) );
  OAI22_X1 U9455 ( .A1(n7963), .A2(n8858), .B1(n7800), .B2(n8856), .ZN(n7809)
         );
  AOI22_X1 U9456 ( .A1(n8241), .A2(n7809), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3152), .ZN(n7783) );
  OAI21_X1 U9457 ( .B1(n10152), .B2(n7814), .A(n7783), .ZN(n7784) );
  AOI21_X1 U9458 ( .B1(n8980), .B2(n10136), .A(n7784), .ZN(n7785) );
  OAI21_X1 U9459 ( .B1(n7786), .B2(n10098), .A(n7785), .ZN(P2_U3228) );
  INV_X1 U9460 ( .A(n7787), .ZN(n7824) );
  INV_X1 U9461 ( .A(n5552), .ZN(n7789) );
  OAI222_X1 U9462 ( .A1(n9878), .A2(n7824), .B1(P1_U3084), .B2(n7789), .C1(
        n7788), .C2(n9874), .ZN(P1_U3327) );
  XNOR2_X1 U9463 ( .A(n7790), .B(n7791), .ZN(n7797) );
  AND2_X1 U9464 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9957) );
  OAI22_X1 U9465 ( .A1(n9164), .A2(n7792), .B1(n9162), .B2(n9113), .ZN(n7793)
         );
  AOI211_X1 U9466 ( .C1(n9167), .C2(n9462), .A(n9957), .B(n7793), .ZN(n7796)
         );
  NAND2_X1 U9467 ( .A1(n7794), .A2(n9142), .ZN(n7795) );
  OAI211_X1 U9468 ( .C1(n7797), .C2(n9144), .A(n7796), .B(n7795), .ZN(P1_U3234) );
  OR2_X1 U9469 ( .A1(n8989), .A2(n8332), .ZN(n7798) );
  NAND2_X1 U9470 ( .A1(n8984), .A2(n7800), .ZN(n7967) );
  NAND2_X1 U9471 ( .A1(n7968), .A2(n7967), .ZN(n7971) );
  NOR2_X1 U9472 ( .A1(n8984), .A2(n8331), .ZN(n7801) );
  AOI21_X2 U9473 ( .B1(n7871), .B2(n7971), .A(n7801), .ZN(n7802) );
  OR2_X1 U9474 ( .A1(n8980), .A2(n8857), .ZN(n8044) );
  NAND2_X1 U9475 ( .A1(n8980), .A2(n8857), .ZN(n8852) );
  NAND2_X1 U9476 ( .A1(n8044), .A2(n8852), .ZN(n7966) );
  NOR2_X1 U9477 ( .A1(n7802), .A2(n7966), .ZN(n7803) );
  OR2_X1 U9478 ( .A1(n8206), .A2(n7803), .ZN(n8983) );
  INV_X1 U9479 ( .A(n8983), .ZN(n7819) );
  INV_X1 U9480 ( .A(n7971), .ZN(n8041) );
  NAND2_X1 U9481 ( .A1(n7878), .A2(n8041), .ZN(n7805) );
  NAND2_X1 U9482 ( .A1(n7805), .A2(n7968), .ZN(n7807) );
  INV_X1 U9483 ( .A(n7966), .ZN(n7806) );
  NAND2_X1 U9484 ( .A1(n7807), .A2(n7966), .ZN(n7808) );
  AOI21_X1 U9485 ( .B1(n8853), .B2(n7808), .A(n8854), .ZN(n7810) );
  AOI211_X1 U9486 ( .C1(n7819), .C2(n7811), .A(n7810), .B(n7809), .ZN(n8982)
         );
  INV_X1 U9487 ( .A(n7872), .ZN(n7812) );
  INV_X1 U9488 ( .A(n8980), .ZN(n7813) );
  AOI211_X1 U9489 ( .C1(n8980), .C2(n7812), .A(n10248), .B(n8862), .ZN(n8979)
         );
  NOR2_X1 U9490 ( .A1(n7813), .A2(n8869), .ZN(n7817) );
  OAI22_X1 U9491 ( .A1(n8881), .A2(n7815), .B1(n7814), .B2(n8888), .ZN(n7816)
         );
  AOI211_X1 U9492 ( .C1(n8979), .C2(n10171), .A(n7817), .B(n7816), .ZN(n7821)
         );
  NAND2_X1 U9493 ( .A1(n7819), .A2(n7818), .ZN(n7820) );
  OAI211_X1 U9494 ( .C1(n8982), .C2(n4392), .A(n7821), .B(n7820), .ZN(P2_U3280) );
  INV_X1 U9495 ( .A(n7822), .ZN(n7825) );
  OAI222_X1 U9496 ( .A1(P2_U3152), .A2(n7825), .B1(n9021), .B2(n7824), .C1(
        n7823), .C2(n9018), .ZN(P2_U3332) );
  NOR2_X1 U9497 ( .A1(n7827), .A2(n7828), .ZN(n7888) );
  AOI211_X1 U9498 ( .C1(n7828), .C2(n7827), .A(n7888), .B(n8377), .ZN(n7838)
         );
  NOR2_X1 U9499 ( .A1(n7829), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7831) );
  NOR2_X1 U9500 ( .A1(n7831), .A2(n7830), .ZN(n7892) );
  XNOR2_X1 U9501 ( .A(n7892), .B(n7893), .ZN(n7832) );
  NOR2_X1 U9502 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7832), .ZN(n7894) );
  AOI21_X1 U9503 ( .B1(n7832), .B2(P2_REG2_REG_15__SCAN_IN), .A(n7894), .ZN(
        n7833) );
  NOR2_X1 U9504 ( .A1(n7833), .A2(n8368), .ZN(n7837) );
  NOR2_X1 U9505 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6179), .ZN(n7834) );
  AOI21_X1 U9506 ( .B1(n8350), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7834), .ZN(
        n7835) );
  OAI21_X1 U9507 ( .B1(n8376), .B2(n7887), .A(n7835), .ZN(n7836) );
  OR3_X1 U9508 ( .A1(n7838), .A2(n7837), .A3(n7836), .ZN(P2_U3260) );
  XNOR2_X1 U9509 ( .A(n7839), .B(n4578), .ZN(n7927) );
  INV_X1 U9510 ( .A(n7927), .ZN(n7851) );
  NAND2_X1 U9511 ( .A1(n7840), .A2(n9709), .ZN(n7841) );
  AOI21_X1 U9512 ( .B1(n7842), .B2(n7841), .A(n10020), .ZN(n7926) );
  OAI211_X1 U9513 ( .C1(n7843), .C2(n9171), .A(n10003), .B(n9722), .ZN(n7924)
         );
  OAI22_X1 U9514 ( .A1(n9629), .A2(n7649), .B1(n9163), .B2(n10008), .ZN(n7845)
         );
  NOR2_X1 U9515 ( .A1(n9720), .A2(n9699), .ZN(n7844) );
  AOI211_X1 U9516 ( .C1(n9718), .C2(n9817), .A(n7845), .B(n7844), .ZN(n7848)
         );
  NAND2_X1 U9517 ( .A1(n7846), .A2(n10028), .ZN(n7847) );
  OAI211_X1 U9518 ( .C1(n7924), .C2(n9724), .A(n7848), .B(n7847), .ZN(n7849)
         );
  AOI21_X1 U9519 ( .B1(n7926), .B2(n9629), .A(n7849), .ZN(n7850) );
  OAI21_X1 U9520 ( .B1(n7851), .B2(n9706), .A(n7850), .ZN(P1_U3276) );
  NOR2_X1 U9521 ( .A1(n4917), .A2(n7853), .ZN(n7854) );
  XNOR2_X1 U9522 ( .A(n7852), .B(n7854), .ZN(n7858) );
  INV_X1 U9523 ( .A(n8827), .ZN(n8795) );
  AOI22_X1 U9524 ( .A1(n8817), .A2(n8303), .B1(n10138), .B2(n8795), .ZN(n7855)
         );
  NAND2_X1 U9525 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8386) );
  OAI211_X1 U9526 ( .C1(n8859), .C2(n10095), .A(n7855), .B(n8386), .ZN(n7856)
         );
  AOI21_X1 U9527 ( .B1(n8966), .B2(n10136), .A(n7856), .ZN(n7857) );
  OAI21_X1 U9528 ( .B1(n7858), .B2(n10098), .A(n7857), .ZN(P2_U3221) );
  INV_X1 U9529 ( .A(n7859), .ZN(n7884) );
  OAI222_X1 U9530 ( .A1(n9878), .A2(n7884), .B1(n7861), .B2(P1_U3084), .C1(
        n7860), .C2(n9874), .ZN(P1_U3326) );
  INV_X1 U9531 ( .A(n9058), .ZN(n7870) );
  AOI22_X1 U9532 ( .A1(n9461), .A2(n9819), .B1(n9818), .B2(n9460), .ZN(n7863)
         );
  NAND3_X1 U9533 ( .A1(n7864), .A2(n7863), .A3(n7862), .ZN(n7865) );
  AOI21_X1 U9534 ( .B1(n7866), .B2(n10066), .A(n7865), .ZN(n7868) );
  MUX2_X1 U9535 ( .A(n5172), .B(n7868), .S(n10076), .Z(n7867) );
  OAI21_X1 U9536 ( .B1(n7870), .B2(n9864), .A(n7867), .ZN(P1_U3490) );
  MUX2_X1 U9537 ( .A(n5169), .B(n7868), .S(n10083), .Z(n7869) );
  OAI21_X1 U9538 ( .B1(n7870), .B2(n9815), .A(n7869), .ZN(P1_U3535) );
  XNOR2_X1 U9539 ( .A(n7871), .B(n8041), .ZN(n8988) );
  AOI21_X1 U9540 ( .B1(n8984), .B2(n7873), .A(n7872), .ZN(n8985) );
  INV_X1 U9541 ( .A(n7874), .ZN(n7875) );
  AOI22_X1 U9542 ( .A1(n4392), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7875), .B2(
        n10159), .ZN(n7876) );
  OAI21_X1 U9543 ( .B1(n7877), .B2(n8869), .A(n7876), .ZN(n7881) );
  XNOR2_X1 U9544 ( .A(n7878), .B(n7971), .ZN(n7879) );
  AOI222_X1 U9545 ( .A1(n10156), .A2(n7879), .B1(n8330), .B2(n8879), .C1(n8332), .C2(n8877), .ZN(n8987) );
  NOR2_X1 U9546 ( .A1(n8987), .A2(n4392), .ZN(n7880) );
  AOI211_X1 U9547 ( .C1(n8985), .C2(n6504), .A(n7881), .B(n7880), .ZN(n7882)
         );
  OAI21_X1 U9548 ( .B1(n8988), .B2(n8874), .A(n7882), .ZN(P2_U3281) );
  NOR2_X1 U9549 ( .A1(n7887), .A2(n7886), .ZN(n7889) );
  NOR2_X1 U9550 ( .A1(n7889), .A2(n7888), .ZN(n7891) );
  XOR2_X1 U9551 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8345), .Z(n7890) );
  NAND2_X1 U9552 ( .A1(n7890), .A2(n7891), .ZN(n8344) );
  OAI21_X1 U9553 ( .B1(n7891), .B2(n7890), .A(n8344), .ZN(n7905) );
  NOR2_X1 U9554 ( .A1(n7893), .A2(n7892), .ZN(n7895) );
  NOR2_X1 U9555 ( .A1(n7895), .A2(n7894), .ZN(n7898) );
  NAND2_X1 U9556 ( .A1(n8345), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8340) );
  INV_X1 U9557 ( .A(n8340), .ZN(n7896) );
  AOI21_X1 U9558 ( .B1(n7815), .B2(n7903), .A(n7896), .ZN(n7897) );
  NAND2_X1 U9559 ( .A1(n7897), .A2(n7898), .ZN(n8339) );
  OAI211_X1 U9560 ( .C1(n7898), .C2(n7897), .A(n8382), .B(n8339), .ZN(n7902)
         );
  NOR2_X1 U9561 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7899), .ZN(n7900) );
  AOI21_X1 U9562 ( .B1(n8350), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n7900), .ZN(
        n7901) );
  OAI211_X1 U9563 ( .C1(n8376), .C2(n7903), .A(n7902), .B(n7901), .ZN(n7904)
         );
  AOI21_X1 U9564 ( .B1(n8381), .B2(n7905), .A(n7904), .ZN(n7906) );
  INV_X1 U9565 ( .A(n7906), .ZN(P2_U3261) );
  NAND2_X1 U9566 ( .A1(n7911), .A2(n7907), .ZN(n7909) );
  OAI211_X1 U9567 ( .C1(n9874), .C2(n7910), .A(n7909), .B(n7908), .ZN(P1_U3325) );
  NAND2_X1 U9568 ( .A1(n7911), .A2(n9016), .ZN(n7913) );
  OAI211_X1 U9569 ( .C1(n9018), .C2(n7914), .A(n7913), .B(n7912), .ZN(P2_U3330) );
  INV_X1 U9570 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n7918) );
  AOI211_X1 U9571 ( .C1(n7917), .C2(n10066), .A(n7916), .B(n7915), .ZN(n7920)
         );
  MUX2_X1 U9572 ( .A(n7918), .B(n7920), .S(n10076), .Z(n7919) );
  OAI21_X1 U9573 ( .B1(n7922), .B2(n9864), .A(n7919), .ZN(P1_U3496) );
  MUX2_X1 U9574 ( .A(n7537), .B(n7920), .S(n10083), .Z(n7921) );
  OAI21_X1 U9575 ( .B1(n7922), .B2(n9815), .A(n7921), .ZN(P1_U3537) );
  INV_X1 U9576 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7928) );
  AOI22_X1 U9577 ( .A1(n9459), .A2(n9818), .B1(n9819), .B2(n9817), .ZN(n7923)
         );
  NAND2_X1 U9578 ( .A1(n7924), .A2(n7923), .ZN(n7925) );
  AOI211_X1 U9579 ( .C1(n7927), .C2(n10066), .A(n7926), .B(n7925), .ZN(n7930)
         );
  MUX2_X1 U9580 ( .A(n7928), .B(n7930), .S(n10076), .Z(n7929) );
  OAI21_X1 U9581 ( .B1(n9171), .B2(n9864), .A(n7929), .ZN(P1_U3499) );
  MUX2_X1 U9582 ( .A(n7931), .B(n7930), .S(n10083), .Z(n7932) );
  OAI21_X1 U9583 ( .B1(n9171), .B2(n9815), .A(n7932), .ZN(P1_U3538) );
  OAI222_X1 U9584 ( .A1(n7956), .A2(P2_U3152), .B1(n9021), .B2(n7934), .C1(
        n7933), .C2(n9018), .ZN(P2_U3336) );
  NOR2_X1 U9585 ( .A1(n7935), .A2(n7942), .ZN(n7937) );
  NAND2_X1 U9586 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9477), .ZN(n7938) );
  OAI21_X1 U9587 ( .B1(n9477), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7938), .ZN(
        n9473) );
  AOI21_X1 U9588 ( .B1(n9477), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9472), .ZN(
        n9486) );
  XNOR2_X1 U9589 ( .A(n9487), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n9485) );
  NOR2_X1 U9590 ( .A1(n9486), .A2(n9485), .ZN(n9484) );
  NAND2_X1 U9591 ( .A1(n9993), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7939) );
  OAI21_X1 U9592 ( .B1(n9993), .B2(P1_REG2_REG_18__SCAN_IN), .A(n7939), .ZN(
        n9988) );
  INV_X1 U9593 ( .A(n7949), .ZN(n7947) );
  AOI22_X1 U9594 ( .A1(n9993), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n9798), .B2(
        n7940), .ZN(n9996) );
  NOR2_X1 U9595 ( .A1(n7942), .A2(n7941), .ZN(n7944) );
  NOR2_X1 U9596 ( .A1(n7944), .A2(n7943), .ZN(n9476) );
  XNOR2_X1 U9597 ( .A(n9477), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9475) );
  NOR2_X1 U9598 ( .A1(n9476), .A2(n9475), .ZN(n9474) );
  AOI21_X1 U9599 ( .B1(n9477), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9474), .ZN(
        n9495) );
  XNOR2_X1 U9600 ( .A(n9487), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9494) );
  NOR2_X1 U9601 ( .A1(n9495), .A2(n9494), .ZN(n9493) );
  AOI21_X1 U9602 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9487), .A(n9493), .ZN(
        n9995) );
  NAND2_X1 U9603 ( .A1(n9996), .A2(n9995), .ZN(n9994) );
  OAI21_X1 U9604 ( .B1(n9993), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9994), .ZN(
        n7945) );
  XNOR2_X1 U9605 ( .A(n7945), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n7948) );
  OAI21_X1 U9606 ( .B1(n7948), .B2(n9492), .A(n9491), .ZN(n7946) );
  AOI21_X1 U9607 ( .B1(n7947), .B2(n9966), .A(n7946), .ZN(n7951) );
  AOI22_X1 U9608 ( .A1(n7949), .A2(n9966), .B1(n9998), .B2(n7948), .ZN(n7950)
         );
  MUX2_X1 U9609 ( .A(n7951), .B(n7950), .S(n4390), .Z(n7953) );
  NAND2_X1 U9610 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3084), .ZN(n7952) );
  OAI211_X1 U9611 ( .C1(n4954), .C2(n9984), .A(n7953), .B(n7952), .ZN(P1_U3260) );
  NAND2_X1 U9612 ( .A1(n8935), .A2(n8271), .ZN(n8062) );
  NAND2_X1 U9613 ( .A1(n8926), .A2(n8260), .ZN(n8127) );
  NAND2_X1 U9614 ( .A1(n8724), .A2(n8322), .ZN(n7954) );
  NAND2_X1 U9615 ( .A1(n8127), .A2(n7954), .ZN(n7958) );
  OR2_X1 U9616 ( .A1(n7958), .A2(n8124), .ZN(n7957) );
  NOR2_X1 U9617 ( .A1(n8104), .A2(n8865), .ZN(n7955) );
  MUX2_X1 U9618 ( .A(n8062), .B(n7957), .S(n8098), .Z(n8067) );
  INV_X1 U9619 ( .A(n8109), .ZN(n7962) );
  OR2_X1 U9620 ( .A1(n8966), .A2(n8293), .ZN(n8111) );
  AND2_X1 U9621 ( .A1(n8111), .A2(n8097), .ZN(n7959) );
  NAND2_X1 U9622 ( .A1(n8118), .A2(n7959), .ZN(n8051) );
  NAND2_X1 U9623 ( .A1(n8958), .A2(n8827), .ZN(n8114) );
  NAND2_X1 U9624 ( .A1(n8966), .A2(n8293), .ZN(n8801) );
  AND2_X1 U9625 ( .A1(n8801), .A2(n8098), .ZN(n7960) );
  NAND2_X1 U9626 ( .A1(n8114), .A2(n7960), .ZN(n8050) );
  NAND2_X1 U9627 ( .A1(n8969), .A2(n8859), .ZN(n8108) );
  INV_X1 U9628 ( .A(n8108), .ZN(n7961) );
  OAI22_X1 U9629 ( .A1(n7962), .A2(n8051), .B1(n8050), .B2(n7961), .ZN(n8049)
         );
  NAND2_X1 U9630 ( .A1(n8975), .A2(n7963), .ZN(n7965) );
  AND2_X1 U9631 ( .A1(n8108), .A2(n7965), .ZN(n7964) );
  MUX2_X1 U9632 ( .A(n8107), .B(n7964), .S(n8097), .Z(n8047) );
  NAND2_X1 U9633 ( .A1(n8107), .A2(n7965), .ZN(n8848) );
  INV_X1 U9634 ( .A(n8848), .ZN(n8851) );
  MUX2_X1 U9635 ( .A(n7968), .B(n7967), .S(n8097), .Z(n8043) );
  NAND2_X1 U9636 ( .A1(n8037), .A2(n7573), .ZN(n7970) );
  NOR2_X1 U9637 ( .A1(n7971), .A2(n7970), .ZN(n8158) );
  AND2_X1 U9638 ( .A1(n7973), .A2(n7972), .ZN(n8016) );
  INV_X1 U9639 ( .A(n8016), .ZN(n7974) );
  NAND2_X1 U9640 ( .A1(n7974), .A2(n8015), .ZN(n7975) );
  AND2_X1 U9641 ( .A1(n8022), .A2(n7975), .ZN(n8013) );
  AND2_X1 U9642 ( .A1(n7987), .A2(n8171), .ZN(n7976) );
  OAI211_X1 U9643 ( .C1(n6906), .C2(n7976), .A(n7991), .B(n7988), .ZN(n7977)
         );
  NAND3_X1 U9644 ( .A1(n7977), .A2(n8098), .A3(n7989), .ZN(n7980) );
  AOI21_X1 U9645 ( .B1(n7981), .B2(n7978), .A(n8097), .ZN(n7979) );
  AOI21_X1 U9646 ( .B1(n7980), .B2(n6907), .A(n7979), .ZN(n7986) );
  NAND2_X1 U9647 ( .A1(n7984), .A2(n7981), .ZN(n7983) );
  NAND2_X1 U9648 ( .A1(n7995), .A2(n7997), .ZN(n7982) );
  AND2_X1 U9649 ( .A1(n7984), .A2(n7999), .ZN(n7985) );
  NAND2_X1 U9650 ( .A1(n7988), .A2(n7987), .ZN(n8144) );
  NAND3_X1 U9651 ( .A1(n8144), .A2(n7990), .A3(n7989), .ZN(n7992) );
  NAND3_X1 U9652 ( .A1(n7992), .A2(n8097), .A3(n7991), .ZN(n7993) );
  AND2_X1 U9653 ( .A1(n7995), .A2(n7994), .ZN(n7998) );
  OAI21_X1 U9654 ( .B1(n8098), .B2(n7999), .A(n8151), .ZN(n8000) );
  MUX2_X1 U9655 ( .A(n8002), .B(n8001), .S(n8098), .Z(n8003) );
  NAND2_X1 U9656 ( .A1(n8150), .A2(n8003), .ZN(n8004) );
  OR2_X1 U9657 ( .A1(n8005), .A2(n8004), .ZN(n8010) );
  MUX2_X1 U9658 ( .A(n8007), .B(n8006), .S(n8098), .Z(n8008) );
  AND2_X1 U9659 ( .A1(n8014), .A2(n8008), .ZN(n8009) );
  NAND2_X1 U9660 ( .A1(n8010), .A2(n8009), .ZN(n8017) );
  NAND2_X1 U9661 ( .A1(n8020), .A2(n8015), .ZN(n8011) );
  AOI21_X1 U9662 ( .B1(n8017), .B2(n8016), .A(n8011), .ZN(n8012) );
  MUX2_X1 U9663 ( .A(n8013), .B(n8012), .S(n8097), .Z(n8019) );
  NAND4_X1 U9664 ( .A1(n8017), .A2(n8016), .A3(n8015), .A4(n8014), .ZN(n8018)
         );
  NAND2_X1 U9665 ( .A1(n8019), .A2(n8018), .ZN(n8023) );
  NAND3_X1 U9666 ( .A1(n8023), .A2(n8020), .A3(n8026), .ZN(n8021) );
  NAND2_X1 U9667 ( .A1(n8021), .A2(n8024), .ZN(n8029) );
  NAND2_X1 U9668 ( .A1(n8023), .A2(n8022), .ZN(n8027) );
  INV_X1 U9669 ( .A(n8024), .ZN(n8025) );
  AOI21_X1 U9670 ( .B1(n8027), .B2(n8026), .A(n8025), .ZN(n8028) );
  MUX2_X1 U9671 ( .A(n8031), .B(n8030), .S(n8098), .Z(n8039) );
  NOR2_X1 U9672 ( .A1(n8032), .A2(n8097), .ZN(n8035) );
  AND2_X1 U9673 ( .A1(n8032), .A2(n8097), .ZN(n8034) );
  MUX2_X1 U9674 ( .A(n8035), .B(n8034), .S(n8033), .Z(n8036) );
  NAND2_X1 U9675 ( .A1(n8037), .A2(n8036), .ZN(n8038) );
  NAND2_X1 U9676 ( .A1(n8039), .A2(n8038), .ZN(n8040) );
  NAND2_X1 U9677 ( .A1(n8041), .A2(n8040), .ZN(n8042) );
  MUX2_X1 U9678 ( .A(n8044), .B(n8852), .S(n8098), .Z(n8045) );
  NAND3_X1 U9679 ( .A1(n8047), .A2(n8109), .A3(n8046), .ZN(n8048) );
  NAND2_X1 U9680 ( .A1(n8049), .A2(n8048), .ZN(n8054) );
  OAI22_X1 U9681 ( .A1(n8801), .A2(n8051), .B1(n8050), .B2(n8111), .ZN(n8052)
         );
  INV_X1 U9682 ( .A(n8052), .ZN(n8053) );
  NAND2_X1 U9683 ( .A1(n8054), .A2(n8053), .ZN(n8057) );
  INV_X1 U9684 ( .A(n8804), .ZN(n8292) );
  AND2_X1 U9685 ( .A1(n8952), .A2(n8292), .ZN(n8121) );
  INV_X1 U9686 ( .A(n8114), .ZN(n8055) );
  OR2_X1 U9687 ( .A1(n8952), .A2(n8292), .ZN(n8058) );
  AND2_X1 U9688 ( .A1(n8120), .A2(n8058), .ZN(n8056) );
  NAND2_X1 U9689 ( .A1(n8946), .A2(n8251), .ZN(n8119) );
  INV_X1 U9690 ( .A(n8121), .ZN(n8775) );
  OAI21_X1 U9691 ( .B1(n8057), .B2(n4773), .A(n8775), .ZN(n8059) );
  NAND2_X1 U9692 ( .A1(n8059), .A2(n8058), .ZN(n8060) );
  INV_X1 U9693 ( .A(n8120), .ZN(n8122) );
  AOI21_X1 U9694 ( .B1(n8060), .B2(n8119), .A(n8122), .ZN(n8061) );
  OR2_X1 U9695 ( .A1(n8940), .A2(n8236), .ZN(n8063) );
  NAND2_X1 U9696 ( .A1(n8940), .A2(n8236), .ZN(n8746) );
  NAND2_X1 U9697 ( .A1(n8063), .A2(n8746), .ZN(n8757) );
  INV_X1 U9698 ( .A(n8757), .ZN(n8758) );
  MUX2_X1 U9699 ( .A(n8063), .B(n8746), .S(n8098), .Z(n8064) );
  NAND3_X1 U9700 ( .A1(n8065), .A2(n8212), .A3(n8064), .ZN(n8066) );
  XNOR2_X1 U9701 ( .A(n8724), .B(n8322), .ZN(n8725) );
  INV_X1 U9702 ( .A(n8725), .ZN(n8163) );
  NAND3_X1 U9703 ( .A1(n4428), .A2(n4747), .A3(n8126), .ZN(n8072) );
  NOR2_X1 U9704 ( .A1(n8701), .A2(n4749), .ZN(n8069) );
  OR2_X1 U9705 ( .A1(n8920), .A2(n8681), .ZN(n8128) );
  NAND2_X1 U9706 ( .A1(n8130), .A2(n8128), .ZN(n8068) );
  AOI21_X1 U9707 ( .B1(n8070), .B2(n8069), .A(n8068), .ZN(n8071) );
  MUX2_X1 U9708 ( .A(n8072), .B(n8071), .S(n8097), .Z(n8075) );
  NAND2_X1 U9709 ( .A1(n8685), .A2(n8204), .ZN(n8129) );
  NAND3_X1 U9710 ( .A1(n8920), .A2(n8681), .A3(n8098), .ZN(n8073) );
  AND2_X1 U9711 ( .A1(n8129), .A2(n8073), .ZN(n8074) );
  NAND2_X1 U9712 ( .A1(n8075), .A2(n8074), .ZN(n8081) );
  NAND2_X1 U9713 ( .A1(n8081), .A2(n8204), .ZN(n8078) );
  NAND2_X1 U9714 ( .A1(n8202), .A2(n6164), .ZN(n8077) );
  NAND2_X1 U9715 ( .A1(n8905), .A2(n8682), .ZN(n8132) );
  NAND2_X1 U9716 ( .A1(n8078), .A2(n8222), .ZN(n8080) );
  NAND2_X1 U9717 ( .A1(n8084), .A2(n8097), .ZN(n8079) );
  NAND2_X1 U9718 ( .A1(n8080), .A2(n8079), .ZN(n8083) );
  OAI211_X1 U9719 ( .C1(n8097), .C2(n8685), .A(n8081), .B(n8129), .ZN(n8082)
         );
  MUX2_X1 U9720 ( .A(n8132), .B(n8084), .S(n8098), .Z(n8092) );
  NAND2_X1 U9721 ( .A1(n8234), .A2(n6164), .ZN(n8086) );
  INV_X1 U9722 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8235) );
  INV_X1 U9723 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8670) );
  NAND2_X1 U9724 ( .A1(n8087), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8089) );
  NAND2_X1 U9725 ( .A1(n5901), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8088) );
  OAI211_X1 U9726 ( .C1(n4396), .C2(n8670), .A(n8089), .B(n8088), .ZN(n8328)
         );
  INV_X1 U9727 ( .A(n8328), .ZN(n8090) );
  NAND2_X1 U9728 ( .A1(n8134), .A2(n8090), .ZN(n8096) );
  NAND2_X1 U9729 ( .A1(n8137), .A2(n8096), .ZN(n8091) );
  NAND2_X1 U9730 ( .A1(n9868), .A2(n6164), .ZN(n8094) );
  INV_X1 U9731 ( .A(n8392), .ZN(n8095) );
  MUX2_X1 U9732 ( .A(n8167), .B(n8168), .S(n8097), .Z(n8102) );
  MUX2_X1 U9733 ( .A(n8100), .B(n8099), .S(n8098), .Z(n8101) );
  INV_X1 U9734 ( .A(n6494), .ZN(n8103) );
  NOR3_X1 U9735 ( .A1(n8173), .A2(n4779), .A3(n8103), .ZN(n8177) );
  INV_X1 U9736 ( .A(n8852), .ZN(n8105) );
  NOR2_X1 U9737 ( .A1(n8848), .A2(n8105), .ZN(n8106) );
  NAND2_X1 U9738 ( .A1(n8840), .A2(n8832), .ZN(n8110) );
  NAND2_X1 U9739 ( .A1(n8110), .A2(n8109), .ZN(n8822) );
  INV_X1 U9740 ( .A(n8822), .ZN(n8113) );
  NAND2_X1 U9741 ( .A1(n8111), .A2(n8801), .ZN(n8825) );
  INV_X1 U9742 ( .A(n8805), .ZN(n8116) );
  INV_X1 U9743 ( .A(n8801), .ZN(n8115) );
  NOR2_X1 U9744 ( .A1(n8116), .A2(n8115), .ZN(n8117) );
  XNOR2_X1 U9745 ( .A(n8952), .B(n8292), .ZN(n8160) );
  INV_X1 U9746 ( .A(n8776), .ZN(n8773) );
  NOR2_X1 U9747 ( .A1(n8773), .A2(n8121), .ZN(n8123) );
  NAND2_X1 U9748 ( .A1(n8212), .A2(n8746), .ZN(n8125) );
  OAI21_X2 U9749 ( .B1(n8761), .B2(n8125), .A(n8124), .ZN(n8726) );
  NAND2_X1 U9750 ( .A1(n8126), .A2(n8127), .ZN(n8708) );
  INV_X1 U9751 ( .A(n8708), .ZN(n8713) );
  NAND2_X1 U9752 ( .A1(n8130), .A2(n8129), .ZN(n8675) );
  INV_X1 U9753 ( .A(n8675), .ZN(n8678) );
  INV_X1 U9754 ( .A(n8130), .ZN(n8131) );
  AOI21_X1 U9755 ( .B1(n8679), .B2(n8678), .A(n8131), .ZN(n8221) );
  NAND2_X1 U9756 ( .A1(n8221), .A2(n8222), .ZN(n8220) );
  NAND2_X1 U9757 ( .A1(n8220), .A2(n8135), .ZN(n8136) );
  OAI21_X1 U9758 ( .B1(n4467), .B2(n8137), .A(n8136), .ZN(n8140) );
  INV_X1 U9759 ( .A(n8222), .ZN(n8166) );
  INV_X1 U9760 ( .A(n8832), .ZN(n8839) );
  OR4_X1 U9761 ( .A1(n8146), .A2(n6906), .A3(n8145), .A4(n8144), .ZN(n8148) );
  NOR4_X1 U9762 ( .A1(n8149), .A2(n8148), .A3(n8147), .A4(n6905), .ZN(n8152)
         );
  NAND4_X1 U9763 ( .A1(n8152), .A2(n8151), .A3(n8150), .A4(n8893), .ZN(n8153)
         );
  NOR4_X1 U9764 ( .A1(n8156), .A2(n8155), .A3(n8154), .A4(n8153), .ZN(n8157)
         );
  NAND4_X1 U9765 ( .A1(n7806), .A2(n8158), .A3(n10154), .A4(n8157), .ZN(n8159)
         );
  NOR4_X1 U9766 ( .A1(n8825), .A2(n8839), .A3(n8848), .A4(n8159), .ZN(n8161)
         );
  INV_X1 U9767 ( .A(n8160), .ZN(n8794) );
  NAND4_X1 U9768 ( .A1(n8776), .A2(n8805), .A3(n8161), .A4(n8794), .ZN(n8162)
         );
  NOR4_X1 U9769 ( .A1(n8708), .A2(n8757), .A3(n8748), .A4(n8162), .ZN(n8164)
         );
  NAND4_X1 U9770 ( .A1(n8678), .A2(n8164), .A3(n8163), .A4(n4747), .ZN(n8165)
         );
  XNOR2_X1 U9771 ( .A(n8169), .B(n8734), .ZN(n8172) );
  OAI22_X1 U9772 ( .A1(n8172), .A2(n8171), .B1(n8170), .B2(n6494), .ZN(n8174)
         );
  NAND2_X1 U9773 ( .A1(n8174), .A2(n8173), .ZN(n8175) );
  NOR2_X1 U9774 ( .A1(n8177), .A2(n8176), .ZN(n8183) );
  NOR4_X1 U9775 ( .A1(n10176), .A2(n8856), .A3(n8223), .A4(n8178), .ZN(n8181)
         );
  OAI21_X1 U9776 ( .B1(n8182), .B2(n8179), .A(P2_B_REG_SCAN_IN), .ZN(n8180) );
  OAI22_X1 U9777 ( .A1(n8183), .A2(n8182), .B1(n8181), .B2(n8180), .ZN(
        P2_U3244) );
  OAI21_X1 U9778 ( .B1(n9287), .B2(n9864), .A(n8186), .ZN(P1_U3522) );
  NOR2_X1 U9779 ( .A1(n10024), .A2(n9731), .ZN(n9503) );
  NOR2_X1 U9780 ( .A1(n9287), .A2(n9623), .ZN(n8187) );
  AOI211_X1 U9781 ( .C1(n10024), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9503), .B(
        n8187), .ZN(n8188) );
  OAI21_X1 U9782 ( .B1(n9724), .B2(n8189), .A(n8188), .ZN(P1_U3261) );
  AOI21_X1 U9783 ( .B1(n8190), .B2(n8191), .A(n10098), .ZN(n8194) );
  NOR3_X1 U9784 ( .A1(n8192), .A2(n8260), .A3(n8315), .ZN(n8193) );
  NOR2_X1 U9785 ( .A1(n8194), .A2(n8193), .ZN(n8201) );
  OAI22_X1 U9786 ( .A1(n10130), .A2(n8204), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8195), .ZN(n8198) );
  INV_X1 U9787 ( .A(n8698), .ZN(n8196) );
  OAI22_X1 U9788 ( .A1(n10095), .A2(n8260), .B1(n10152), .B2(n8196), .ZN(n8197) );
  AOI211_X1 U9789 ( .C1(n8920), .C2(n10136), .A(n8198), .B(n8197), .ZN(n8199)
         );
  OAI21_X1 U9790 ( .B1(n8201), .B2(n8200), .A(n8199), .ZN(P2_U3216) );
  INV_X1 U9791 ( .A(n8202), .ZN(n9020) );
  OAI222_X1 U9792 ( .A1(n9878), .A2(n9020), .B1(n8203), .B2(P1_U3084), .C1(
        n8607), .C2(n9874), .ZN(P1_U3324) );
  INV_X1 U9793 ( .A(n8940), .ZN(n8211) );
  NOR2_X2 U9794 ( .A1(n8206), .A2(n8205), .ZN(n8849) );
  INV_X1 U9795 ( .A(n8293), .ZN(n8842) );
  AOI21_X2 U9796 ( .B1(n8795), .B2(n8958), .A(n8963), .ZN(n8788) );
  NOR2_X1 U9797 ( .A1(n8952), .A2(n8804), .ZN(n8210) );
  INV_X1 U9798 ( .A(n8952), .ZN(n8792) );
  INV_X1 U9799 ( .A(n8251), .ZN(n8796) );
  OAI22_X1 U9800 ( .A1(n8740), .A2(n8212), .B1(n8729), .B2(n8935), .ZN(n8723)
         );
  NAND2_X1 U9801 ( .A1(n8723), .A2(n8725), .ZN(n8722) );
  NAND2_X1 U9802 ( .A1(n8722), .A2(n8213), .ZN(n8709) );
  NAND2_X1 U9803 ( .A1(n8676), .A2(n8675), .ZN(n8674) );
  INV_X1 U9804 ( .A(n8935), .ZN(n8745) );
  INV_X1 U9805 ( .A(n8975), .ZN(n8870) );
  NAND2_X1 U9806 ( .A1(n8745), .A2(n8768), .ZN(n8730) );
  INV_X1 U9807 ( .A(n8217), .ZN(n8218) );
  AOI22_X1 U9808 ( .A1(n4392), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8218), .B2(
        n10159), .ZN(n8219) );
  OAI21_X1 U9809 ( .B1(n4548), .B2(n8869), .A(n8219), .ZN(n8231) );
  OAI21_X1 U9810 ( .B1(n8222), .B2(n8221), .A(n8220), .ZN(n8229) );
  INV_X1 U9811 ( .A(n8223), .ZN(n8224) );
  AND2_X1 U9812 ( .A1(n8224), .A2(P2_B_REG_SCAN_IN), .ZN(n8225) );
  NOR2_X1 U9813 ( .A1(n8858), .A2(n8225), .ZN(n8391) );
  NAND2_X1 U9814 ( .A1(n8391), .A2(n8328), .ZN(n8226) );
  AOI211_X1 U9815 ( .C1(n6504), .C2(n8906), .A(n8231), .B(n8230), .ZN(n8232)
         );
  OAI21_X1 U9816 ( .B1(n8909), .B2(n8874), .A(n8232), .ZN(P2_U3267) );
  INV_X1 U9817 ( .A(n8234), .ZN(n9877) );
  OAI222_X1 U9818 ( .A1(P2_U3152), .A2(n8233), .B1(n9021), .B2(n9877), .C1(
        n8235), .C2(n9018), .ZN(P2_U3328) );
  AOI22_X1 U9819 ( .A1(n8238), .A2(n10145), .B1(n10118), .B2(n8779), .ZN(n8245) );
  OR2_X1 U9820 ( .A1(n8271), .A2(n8858), .ZN(n8240) );
  NAND2_X1 U9821 ( .A1(n8796), .A2(n8877), .ZN(n8239) );
  NAND2_X1 U9822 ( .A1(n8240), .A2(n8239), .ZN(n8762) );
  AOI22_X1 U9823 ( .A1(n8241), .A2(n8762), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8242) );
  OAI21_X1 U9824 ( .B1(n10152), .B2(n8764), .A(n8242), .ZN(n8243) );
  AOI21_X1 U9825 ( .B1(n8940), .B2(n10136), .A(n8243), .ZN(n8244) );
  OAI21_X1 U9826 ( .B1(n8245), .B2(n8268), .A(n8244), .ZN(P2_U3218) );
  AOI21_X1 U9827 ( .B1(n8246), .B2(n4464), .A(n10098), .ZN(n8250) );
  NOR3_X1 U9828 ( .A1(n8247), .A2(n8827), .A3(n8315), .ZN(n8249) );
  OAI21_X1 U9829 ( .B1(n8250), .B2(n8249), .A(n8248), .ZN(n8255) );
  OAI22_X1 U9830 ( .A1(n10130), .A2(n8251), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8606), .ZN(n8253) );
  OAI22_X1 U9831 ( .A1(n10095), .A2(n8827), .B1(n10152), .B2(n8789), .ZN(n8252) );
  AOI211_X1 U9832 ( .C1(n8952), .C2(n10136), .A(n8253), .B(n8252), .ZN(n8254)
         );
  NAND2_X1 U9833 ( .A1(n8255), .A2(n8254), .ZN(P2_U3225) );
  AOI21_X1 U9834 ( .B1(n8258), .B2(n8257), .A(n8256), .ZN(n8266) );
  NAND2_X1 U9835 ( .A1(n8724), .A2(n10213), .ZN(n8932) );
  INV_X1 U9836 ( .A(n8932), .ZN(n8264) );
  OAI22_X1 U9837 ( .A1(n10130), .A2(n8260), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8259), .ZN(n8262) );
  OAI22_X1 U9838 ( .A1(n10095), .A2(n8271), .B1(n10152), .B2(n8733), .ZN(n8261) );
  AOI211_X1 U9839 ( .C1(n8264), .C2(n8263), .A(n8262), .B(n8261), .ZN(n8265)
         );
  OAI21_X1 U9840 ( .B1(n8266), .B2(n10098), .A(n8265), .ZN(P2_U3227) );
  NOR2_X1 U9841 ( .A1(n8268), .A2(n8267), .ZN(n8270) );
  XNOR2_X1 U9842 ( .A(n8270), .B(n8269), .ZN(n8274) );
  OAI22_X1 U9843 ( .A1(n8274), .A2(n10098), .B1(n8271), .B2(n8315), .ZN(n8272)
         );
  OAI21_X1 U9844 ( .B1(n8274), .B2(n8273), .A(n8272), .ZN(n8278) );
  AOI22_X1 U9845 ( .A1(n10138), .A2(n8751), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n8277) );
  AOI22_X1 U9846 ( .A1(n8743), .A2(n8303), .B1(n10140), .B2(n8779), .ZN(n8276)
         );
  NAND2_X1 U9847 ( .A1(n8935), .A2(n10136), .ZN(n8275) );
  NAND4_X1 U9848 ( .A1(n8278), .A2(n8277), .A3(n8276), .A4(n8275), .ZN(
        P2_U3231) );
  OAI22_X1 U9849 ( .A1(n8327), .A2(n10202), .B1(n10152), .B2(n8279), .ZN(n8280) );
  AOI211_X1 U9850 ( .C1(n10138), .C2(n8878), .A(n8281), .B(n8280), .ZN(n8290)
         );
  OAI21_X1 U9851 ( .B1(n8285), .B2(n8282), .A(n8283), .ZN(n8284) );
  NAND2_X1 U9852 ( .A1(n10145), .A2(n8284), .ZN(n8289) );
  NOR3_X1 U9853 ( .A1(n8315), .A2(n8286), .A3(n8285), .ZN(n8287) );
  OAI21_X1 U9854 ( .B1(n8287), .B2(n10140), .A(n8337), .ZN(n8288) );
  NAND3_X1 U9855 ( .A1(n8290), .A2(n8289), .A3(n8288), .ZN(P2_U3232) );
  INV_X1 U9856 ( .A(n8958), .ZN(n8810) );
  OAI211_X1 U9857 ( .C1(n8291), .C2(n4460), .A(n8246), .B(n10145), .ZN(n8297)
         );
  NOR2_X1 U9858 ( .A1(n10130), .A2(n8292), .ZN(n8295) );
  OAI22_X1 U9859 ( .A1(n10095), .A2(n8293), .B1(n10152), .B2(n8811), .ZN(n8294) );
  AOI211_X1 U9860 ( .C1(P2_REG3_REG_20__SCAN_IN), .C2(P2_U3152), .A(n8295), 
        .B(n8294), .ZN(n8296) );
  OAI211_X1 U9861 ( .C1(n8810), .C2(n8327), .A(n8297), .B(n8296), .ZN(P2_U3235) );
  NAND2_X1 U9862 ( .A1(n10118), .A2(n8796), .ZN(n8301) );
  NAND2_X1 U9863 ( .A1(n10145), .A2(n8298), .ZN(n8300) );
  MUX2_X1 U9864 ( .A(n8301), .B(n8300), .S(n8299), .Z(n8307) );
  AOI22_X1 U9865 ( .A1(n10140), .A2(n8804), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8306) );
  INV_X1 U9866 ( .A(n8302), .ZN(n8782) );
  AOI22_X1 U9867 ( .A1(n8782), .A2(n8303), .B1(n10138), .B2(n8779), .ZN(n8305)
         );
  NAND2_X1 U9868 ( .A1(n8946), .A2(n10136), .ZN(n8304) );
  NAND4_X1 U9869 ( .A1(n8307), .A2(n8306), .A3(n8305), .A4(n8304), .ZN(
        P2_U3237) );
  INV_X1 U9870 ( .A(n10214), .ZN(n8308) );
  OAI22_X1 U9871 ( .A1(n8327), .A2(n8308), .B1(n10152), .B2(n8887), .ZN(n8309)
         );
  AOI211_X1 U9872 ( .C1(n10138), .C2(n10126), .A(n8310), .B(n8309), .ZN(n8319)
         );
  OAI21_X1 U9873 ( .B1(n8313), .B2(n10144), .A(n8311), .ZN(n8312) );
  NAND2_X1 U9874 ( .A1(n8312), .A2(n10145), .ZN(n8318) );
  NOR3_X1 U9875 ( .A1(n8315), .A2(n8314), .A3(n8313), .ZN(n8316) );
  OAI21_X1 U9876 ( .B1(n8316), .B2(n10140), .A(n8878), .ZN(n8317) );
  NAND3_X1 U9877 ( .A1(n8319), .A2(n8318), .A3(n8317), .ZN(P2_U3241) );
  OAI211_X1 U9878 ( .C1(n8321), .C2(n8320), .A(n8190), .B(n10145), .ZN(n8326)
         );
  NOR2_X1 U9879 ( .A1(n10130), .A2(n8681), .ZN(n8324) );
  OAI22_X1 U9880 ( .A1(n10095), .A2(n8322), .B1(n10152), .B2(n8718), .ZN(n8323) );
  AOI211_X1 U9881 ( .C1(P2_REG3_REG_26__SCAN_IN), .C2(P2_U3152), .A(n8324), 
        .B(n8323), .ZN(n8325) );
  OAI211_X1 U9882 ( .C1(n8214), .C2(n8327), .A(n8326), .B(n8325), .ZN(P2_U3242) );
  MUX2_X1 U9883 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8328), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9884 ( .A(n8329), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8338), .Z(
        P2_U3581) );
  MUX2_X1 U9885 ( .A(n8702), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8338), .Z(
        P2_U3580) );
  MUX2_X1 U9886 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8714), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9887 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8728), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U9888 ( .A(n8751), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8338), .Z(
        P2_U3577) );
  MUX2_X1 U9889 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8729), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U9890 ( .A(n8779), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8338), .Z(
        P2_U3575) );
  MUX2_X1 U9891 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8796), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9892 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8804), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U9893 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8795), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9894 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8842), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9895 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n4866), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9896 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8841), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9897 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8330), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9898 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8331), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9899 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8332), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9900 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8333), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9901 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8334), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9902 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n10093), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U9903 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8335), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U9904 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8336), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U9905 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n10084), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U9906 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n10126), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U9907 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n10137), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U9908 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8878), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U9909 ( .A(n10139), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8338), .Z(
        P2_U3556) );
  MUX2_X1 U9910 ( .A(n8337), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8338), .Z(
        P2_U3555) );
  MUX2_X1 U9911 ( .A(n10111), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8338), .Z(
        P2_U3554) );
  MUX2_X1 U9912 ( .A(n6491), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8338), .Z(
        P2_U3553) );
  MUX2_X1 U9913 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n6497), .S(P2_U3966), .Z(
        P2_U3552) );
  NAND2_X1 U9914 ( .A1(n8340), .A2(n8339), .ZN(n8343) );
  OR2_X1 U9915 ( .A1(n8358), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8341) );
  NAND2_X1 U9916 ( .A1(n8358), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8355) );
  AND2_X1 U9917 ( .A1(n8341), .A2(n8355), .ZN(n8342) );
  NAND2_X1 U9918 ( .A1(n8342), .A2(n8343), .ZN(n8354) );
  OAI211_X1 U9919 ( .C1(n8343), .C2(n8342), .A(n8382), .B(n8354), .ZN(n8352)
         );
  NOR2_X1 U9920 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8652), .ZN(n8349) );
  OAI21_X1 U9921 ( .B1(n8345), .B2(P2_REG1_REG_16__SCAN_IN), .A(n8344), .ZN(
        n8347) );
  XNOR2_X1 U9922 ( .A(n8358), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8346) );
  NOR2_X1 U9923 ( .A1(n8346), .A2(n8347), .ZN(n8357) );
  AOI211_X1 U9924 ( .C1(n8347), .C2(n8346), .A(n8357), .B(n8377), .ZN(n8348)
         );
  AOI211_X1 U9925 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n8350), .A(n8349), .B(
        n8348), .ZN(n8351) );
  OAI211_X1 U9926 ( .C1(n8376), .C2(n8353), .A(n8352), .B(n8351), .ZN(P2_U3262) );
  NAND2_X1 U9927 ( .A1(n8355), .A2(n8354), .ZN(n8370) );
  XOR2_X1 U9928 ( .A(n8362), .B(n8370), .Z(n8356) );
  NOR2_X1 U9929 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8356), .ZN(n8372) );
  AOI21_X1 U9930 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8356), .A(n8372), .ZN(
        n8369) );
  AOI22_X1 U9931 ( .A1(n8375), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n8359), .B2(
        n8362), .ZN(n8360) );
  OAI21_X1 U9932 ( .B1(n8361), .B2(n8360), .A(n8374), .ZN(n8366) );
  NOR2_X1 U9933 ( .A1(n8376), .A2(n8362), .ZN(n8365) );
  INV_X1 U9934 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10315) );
  OAI21_X1 U9935 ( .B1(n8389), .B2(n10315), .A(n8363), .ZN(n8364) );
  AOI211_X1 U9936 ( .C1(n8366), .C2(n8381), .A(n8365), .B(n8364), .ZN(n8367)
         );
  OAI21_X1 U9937 ( .B1(n8369), .B2(n8368), .A(n8367), .ZN(P2_U3263) );
  NOR2_X1 U9938 ( .A1(n8375), .A2(n8370), .ZN(n8371) );
  NOR2_X1 U9939 ( .A1(n8372), .A2(n8371), .ZN(n8373) );
  XOR2_X1 U9940 ( .A(n8373), .B(P2_REG2_REG_19__SCAN_IN), .Z(n8383) );
  INV_X1 U9941 ( .A(n8383), .ZN(n8379) );
  OAI21_X1 U9942 ( .B1(n8380), .B2(n8377), .A(n8376), .ZN(n8378) );
  AOI21_X1 U9943 ( .B1(n8379), .B2(n8382), .A(n8378), .ZN(n8385) );
  AOI22_X1 U9944 ( .A1(n8383), .A2(n8382), .B1(n8381), .B2(n8380), .ZN(n8384)
         );
  MUX2_X1 U9945 ( .A(n8385), .B(n8384), .S(n8865), .Z(n8387) );
  OAI211_X1 U9946 ( .C1(n8389), .C2(n8388), .A(n8387), .B(n8386), .ZN(P2_U3264) );
  NAND2_X1 U9947 ( .A1(n8904), .A2(n8668), .ZN(n8899) );
  INV_X1 U9948 ( .A(n8898), .ZN(n8396) );
  NAND2_X1 U9949 ( .A1(n8390), .A2(n10161), .ZN(n8393) );
  AND2_X1 U9950 ( .A1(n8392), .A2(n8391), .ZN(n8901) );
  NAND2_X1 U9951 ( .A1(n8881), .A2(n8901), .ZN(n8669) );
  OAI211_X1 U9952 ( .C1(n8881), .C2(n8394), .A(n8393), .B(n8669), .ZN(n8395)
         );
  AOI21_X1 U9953 ( .B1(n8396), .B2(n6504), .A(n8395), .ZN(n8667) );
  NOR4_X1 U9954 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_17__SCAN_IN), 
        .A3(P2_REG0_REG_17__SCAN_IN), .A4(P2_REG1_REG_16__SCAN_IN), .ZN(n8397)
         );
  NAND3_X1 U9955 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .A3(n8397), .ZN(n8403) );
  NOR4_X1 U9956 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG1_REG_23__SCAN_IN), 
        .A3(P1_REG0_REG_9__SCAN_IN), .A4(P1_REG1_REG_8__SCAN_IN), .ZN(n8401)
         );
  NOR4_X1 U9957 ( .A1(P1_REG1_REG_26__SCAN_IN), .A2(P2_REG1_REG_10__SCAN_IN), 
        .A3(P2_REG1_REG_8__SCAN_IN), .A4(P2_REG2_REG_5__SCAN_IN), .ZN(n8400)
         );
  NOR4_X1 U9958 ( .A1(P1_REG2_REG_23__SCAN_IN), .A2(P1_REG1_REG_21__SCAN_IN), 
        .A3(P1_REG1_REG_20__SCAN_IN), .A4(P1_REG2_REG_20__SCAN_IN), .ZN(n8399)
         );
  NOR4_X1 U9959 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG2_REG_8__SCAN_IN), .A4(P1_REG3_REG_0__SCAN_IN), .ZN(n8398) );
  NAND4_X1 U9960 ( .A1(n8401), .A2(n8400), .A3(n8399), .A4(n8398), .ZN(n8402)
         );
  OR4_X1 U9961 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(P2_REG2_REG_26__SCAN_IN), 
        .A3(n8403), .A4(n8402), .ZN(n8447) );
  NAND4_X1 U9962 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG0_REG_17__SCAN_IN), 
        .A3(P1_REG1_REG_17__SCAN_IN), .A4(P1_REG0_REG_11__SCAN_IN), .ZN(n8407)
         );
  NAND4_X1 U9963 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG1_REG_10__SCAN_IN), 
        .A3(P1_REG2_REG_6__SCAN_IN), .A4(P1_REG1_REG_4__SCAN_IN), .ZN(n8406)
         );
  NAND4_X1 U9964 ( .A1(P1_REG2_REG_27__SCAN_IN), .A2(P2_REG2_REG_20__SCAN_IN), 
        .A3(P2_REG0_REG_18__SCAN_IN), .A4(P2_REG2_REG_30__SCAN_IN), .ZN(n8405)
         );
  NAND4_X1 U9965 ( .A1(P1_REG2_REG_28__SCAN_IN), .A2(P1_REG0_REG_19__SCAN_IN), 
        .A3(P1_REG1_REG_18__SCAN_IN), .A4(P2_REG0_REG_16__SCAN_IN), .ZN(n8404)
         );
  NOR4_X1 U9966 ( .A1(n8407), .A2(n8406), .A3(n8405), .A4(n8404), .ZN(n8413)
         );
  NAND4_X1 U9967 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .A3(P2_REG0_REG_12__SCAN_IN), .A4(P2_REG2_REG_1__SCAN_IN), .ZN(n8411)
         );
  NAND4_X1 U9968 ( .A1(P2_REG0_REG_26__SCAN_IN), .A2(P2_REG1_REG_21__SCAN_IN), 
        .A3(P2_REG0_REG_7__SCAN_IN), .A4(P2_REG0_REG_24__SCAN_IN), .ZN(n8410)
         );
  NAND4_X1 U9969 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_REG1_REG_24__SCAN_IN), 
        .A3(P2_REG1_REG_7__SCAN_IN), .A4(P2_REG3_REG_0__SCAN_IN), .ZN(n8409)
         );
  NAND4_X1 U9970 ( .A1(P2_REG1_REG_19__SCAN_IN), .A2(P2_REG2_REG_9__SCAN_IN), 
        .A3(P2_REG2_REG_2__SCAN_IN), .A4(P2_REG1_REG_2__SCAN_IN), .ZN(n8408)
         );
  NOR4_X1 U9971 ( .A1(n8411), .A2(n8410), .A3(n8409), .A4(n8408), .ZN(n8412)
         );
  NAND2_X1 U9972 ( .A1(n8413), .A2(n8412), .ZN(n8446) );
  NOR4_X1 U9973 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P2_REG3_REG_13__SCAN_IN), .A4(P2_WR_REG_SCAN_IN), .ZN(n8435) );
  INV_X1 U9974 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n8415) );
  INV_X1 U9975 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8414) );
  NAND4_X1 U9976 ( .A1(n8415), .A2(n8414), .A3(n10312), .A4(n10315), .ZN(n8417) );
  NAND4_X1 U9977 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_D_REG_1__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n8416) );
  NOR2_X1 U9978 ( .A1(n8417), .A2(n8416), .ZN(n8434) );
  NAND4_X1 U9979 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .A3(P2_REG2_REG_25__SCAN_IN), .A4(P2_REG0_REG_28__SCAN_IN), .ZN(n8418)
         );
  INV_X1 U9980 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8647) );
  NOR2_X1 U9981 ( .A1(n8418), .A2(n8647), .ZN(n8423) );
  NOR4_X1 U9982 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .A3(
        P1_IR_REG_8__SCAN_IN), .A4(P1_REG3_REG_6__SCAN_IN), .ZN(n8420) );
  NOR4_X1 U9983 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG0_REG_22__SCAN_IN), 
        .A3(P2_REG1_REG_23__SCAN_IN), .A4(P2_REG0_REG_29__SCAN_IN), .ZN(n8419)
         );
  AND2_X1 U9984 ( .A1(n8420), .A2(n8419), .ZN(n8422) );
  NOR4_X1 U9985 ( .A1(SI_27_), .A2(P2_RD_REG_SCAN_IN), .A3(SI_28_), .A4(
        P2_DATAO_REG_29__SCAN_IN), .ZN(n8421) );
  INV_X1 U9986 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8500) );
  NAND4_X1 U9987 ( .A1(n8423), .A2(n8422), .A3(n8421), .A4(
        P2_IR_REG_20__SCAN_IN), .ZN(n8424) );
  NOR2_X1 U9988 ( .A1(SI_1_), .A2(n8424), .ZN(n8425) );
  NAND3_X1 U9989 ( .A1(n5933), .A2(P1_ADDR_REG_12__SCAN_IN), .A3(n8425), .ZN(
        n8429) );
  INV_X1 U9990 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8426) );
  NAND4_X1 U9991 ( .A1(n5873), .A2(n4798), .A3(n8426), .A4(
        P2_DATAO_REG_1__SCAN_IN), .ZN(n8428) );
  INV_X1 U9992 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9480) );
  NAND4_X1 U9993 ( .A1(n9480), .A2(n8483), .A3(n8606), .A4(
        P2_IR_REG_19__SCAN_IN), .ZN(n8427) );
  NOR3_X1 U9994 ( .A1(n8429), .A2(n8428), .A3(n8427), .ZN(n8433) );
  AND4_X1 U9995 ( .A1(n8431), .A2(n8430), .A3(P2_ADDR_REG_4__SCAN_IN), .A4(
        P2_ADDR_REG_1__SCAN_IN), .ZN(n8432) );
  AND4_X1 U9996 ( .A1(n8435), .A2(n8434), .A3(n8433), .A4(n8432), .ZN(n8444)
         );
  NAND4_X1 U9997 ( .A1(SI_12_), .A2(n8464), .A3(n8557), .A4(n8436), .ZN(n8440)
         );
  INV_X1 U9998 ( .A(SI_18_), .ZN(n8526) );
  NAND4_X1 U9999 ( .A1(SI_20_), .A2(n8552), .A3(n8526), .A4(n8634), .ZN(n8439)
         );
  INV_X1 U10000 ( .A(SI_4_), .ZN(n8532) );
  NAND4_X1 U10001 ( .A1(SI_3_), .A2(P2_DATAO_REG_2__SCAN_IN), .A3(
        P2_DATAO_REG_0__SCAN_IN), .A4(n8532), .ZN(n8438) );
  NAND4_X1 U10002 ( .A1(SI_11_), .A2(P1_DATAO_REG_9__SCAN_IN), .A3(
        P1_DATAO_REG_8__SCAN_IN), .A4(SI_7_), .ZN(n8437) );
  NOR4_X1 U10003 ( .A1(n8440), .A2(n8439), .A3(n8438), .A4(n8437), .ZN(n8443)
         );
  NOR4_X1 U10004 ( .A1(P2_D_REG_0__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_U3152), .A4(n8639), .ZN(n8442) );
  INV_X1 U10005 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10182) );
  INV_X1 U10006 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10180) );
  INV_X1 U10007 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n10177) );
  INV_X1 U10008 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n10183) );
  NOR4_X1 U10009 ( .A1(n10182), .A2(n10180), .A3(n10177), .A4(n10183), .ZN(
        n8441) );
  NAND4_X1 U10010 ( .A1(n8444), .A2(n8443), .A3(n8442), .A4(n8441), .ZN(n8445)
         );
  NOR3_X1 U10011 ( .A1(n8447), .A2(n8446), .A3(n8445), .ZN(n8665) );
  AOI22_X1 U10012 ( .A1(n9853), .A2(keyinput34), .B1(n8449), .B2(keyinput84), 
        .ZN(n8448) );
  OAI221_X1 U10013 ( .B1(n9853), .B2(keyinput34), .C1(n8449), .C2(keyinput84), 
        .A(n8448), .ZN(n8458) );
  AOI22_X1 U10014 ( .A1(n10315), .A2(keyinput18), .B1(n10180), .B2(keyinput53), 
        .ZN(n8450) );
  OAI221_X1 U10015 ( .B1(n10315), .B2(keyinput18), .C1(n10180), .C2(keyinput53), .A(n8450), .ZN(n8457) );
  INV_X1 U10016 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n10178) );
  AOI22_X1 U10017 ( .A1(n10178), .A2(keyinput90), .B1(keyinput36), .B2(n6642), 
        .ZN(n8451) );
  OAI221_X1 U10018 ( .B1(n10178), .B2(keyinput90), .C1(n6642), .C2(keyinput36), 
        .A(n8451), .ZN(n8456) );
  INV_X1 U10019 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8453) );
  AOI22_X1 U10020 ( .A1(n8454), .A2(keyinput64), .B1(keyinput24), .B2(n8453), 
        .ZN(n8452) );
  OAI221_X1 U10021 ( .B1(n8454), .B2(keyinput64), .C1(n8453), .C2(keyinput24), 
        .A(n8452), .ZN(n8455) );
  NOR4_X1 U10022 ( .A1(n8458), .A2(n8457), .A3(n8456), .A4(n8455), .ZN(n8568)
         );
  AOI22_X1 U10023 ( .A1(n5986), .A2(keyinput21), .B1(n10182), .B2(keyinput79), 
        .ZN(n8459) );
  OAI221_X1 U10024 ( .B1(n5986), .B2(keyinput21), .C1(n10182), .C2(keyinput79), 
        .A(n8459), .ZN(n8468) );
  AOI22_X1 U10025 ( .A1(n8462), .A2(keyinput4), .B1(n8461), .B2(keyinput0), 
        .ZN(n8460) );
  OAI221_X1 U10026 ( .B1(n8462), .B2(keyinput4), .C1(n8461), .C2(keyinput0), 
        .A(n8460), .ZN(n8467) );
  AOI22_X1 U10027 ( .A1(n8465), .A2(keyinput122), .B1(n8464), .B2(keyinput33), 
        .ZN(n8463) );
  OAI221_X1 U10028 ( .B1(n8465), .B2(keyinput122), .C1(n8464), .C2(keyinput33), 
        .A(n8463), .ZN(n8466) );
  NOR3_X1 U10029 ( .A1(n8468), .A2(n8467), .A3(n8466), .ZN(n8498) );
  AOI22_X1 U10030 ( .A1(n8470), .A2(keyinput117), .B1(n5467), .B2(keyinput47), 
        .ZN(n8469) );
  OAI221_X1 U10031 ( .B1(n8470), .B2(keyinput117), .C1(n5467), .C2(keyinput47), 
        .A(n8469), .ZN(n8476) );
  XNOR2_X1 U10032 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput102), .ZN(n8474) );
  XNOR2_X1 U10033 ( .A(P2_IR_REG_0__SCAN_IN), .B(keyinput69), .ZN(n8473) );
  XNOR2_X1 U10034 ( .A(P2_REG0_REG_28__SCAN_IN), .B(keyinput22), .ZN(n8472) );
  XNOR2_X1 U10035 ( .A(keyinput94), .B(SI_1_), .ZN(n8471) );
  NAND4_X1 U10036 ( .A1(n8474), .A2(n8473), .A3(n8472), .A4(n8471), .ZN(n8475)
         );
  NOR2_X1 U10037 ( .A1(n8476), .A2(n8475), .ZN(n8497) );
  INV_X1 U10038 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10041) );
  AOI22_X1 U10039 ( .A1(n6335), .A2(keyinput49), .B1(n10041), .B2(keyinput98), 
        .ZN(n8477) );
  OAI221_X1 U10040 ( .B1(n6335), .B2(keyinput49), .C1(n10041), .C2(keyinput98), 
        .A(n8477), .ZN(n8481) );
  INV_X1 U10041 ( .A(P2_RD_REG_SCAN_IN), .ZN(n8479) );
  AOI22_X1 U10042 ( .A1(n8479), .A2(keyinput118), .B1(n4931), .B2(keyinput8), 
        .ZN(n8478) );
  OAI221_X1 U10043 ( .B1(n8479), .B2(keyinput118), .C1(n4931), .C2(keyinput8), 
        .A(n8478), .ZN(n8480) );
  NOR2_X1 U10044 ( .A1(n8481), .A2(n8480), .ZN(n8496) );
  AOI22_X1 U10045 ( .A1(n8484), .A2(keyinput40), .B1(n8483), .B2(keyinput99), 
        .ZN(n8482) );
  OAI221_X1 U10046 ( .B1(n8484), .B2(keyinput40), .C1(n8483), .C2(keyinput99), 
        .A(n8482), .ZN(n8485) );
  INV_X1 U10047 ( .A(n8485), .ZN(n8489) );
  XNOR2_X1 U10048 ( .A(keyinput95), .B(n7278), .ZN(n8487) );
  XNOR2_X1 U10049 ( .A(keyinput37), .B(n9593), .ZN(n8486) );
  NOR2_X1 U10050 ( .A1(n8487), .A2(n8486), .ZN(n8488) );
  NAND2_X1 U10051 ( .A1(n8489), .A2(n8488), .ZN(n8494) );
  INV_X1 U10052 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8491) );
  AOI22_X1 U10053 ( .A1(n8492), .A2(keyinput61), .B1(keyinput42), .B2(n8491), 
        .ZN(n8490) );
  OAI221_X1 U10054 ( .B1(n8492), .B2(keyinput61), .C1(n8491), .C2(keyinput42), 
        .A(n8490), .ZN(n8493) );
  NOR2_X1 U10055 ( .A1(n8494), .A2(n8493), .ZN(n8495) );
  NAND4_X1 U10056 ( .A1(n8498), .A2(n8497), .A3(n8496), .A4(n8495), .ZN(n8523)
         );
  AOI22_X1 U10057 ( .A1(n8500), .A2(keyinput85), .B1(n9151), .B2(keyinput91), 
        .ZN(n8499) );
  OAI221_X1 U10058 ( .B1(n8500), .B2(keyinput85), .C1(n9151), .C2(keyinput91), 
        .A(n8499), .ZN(n8506) );
  XNOR2_X1 U10059 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(keyinput78), .ZN(n8504) );
  XNOR2_X1 U10060 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput93), .ZN(n8503) );
  XNOR2_X1 U10061 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput114), .ZN(n8502)
         );
  XNOR2_X1 U10062 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput65), .ZN(n8501) );
  NAND4_X1 U10063 ( .A1(n8504), .A2(n8503), .A3(n8502), .A4(n8501), .ZN(n8505)
         );
  NOR2_X1 U10064 ( .A1(n8506), .A2(n8505), .ZN(n8521) );
  INV_X1 U10065 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n10181) );
  XNOR2_X1 U10066 ( .A(n10181), .B(keyinput43), .ZN(n8508) );
  XNOR2_X1 U10067 ( .A(n10177), .B(keyinput125), .ZN(n8507) );
  NOR2_X1 U10068 ( .A1(n8508), .A2(n8507), .ZN(n8520) );
  XNOR2_X1 U10069 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput14), .ZN(n8512) );
  XNOR2_X1 U10070 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput116), .ZN(n8511)
         );
  XNOR2_X1 U10071 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput68), .ZN(n8510) );
  XNOR2_X1 U10072 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput81), .ZN(n8509) );
  NAND4_X1 U10073 ( .A1(n8512), .A2(n8511), .A3(n8510), .A4(n8509), .ZN(n8518)
         );
  XNOR2_X1 U10074 ( .A(P2_REG1_REG_19__SCAN_IN), .B(keyinput5), .ZN(n8516) );
  XNOR2_X1 U10075 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput121), .ZN(n8515)
         );
  XNOR2_X1 U10076 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput57), .ZN(n8514) );
  XNOR2_X1 U10077 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput70), .ZN(n8513) );
  NAND4_X1 U10078 ( .A1(n8516), .A2(n8515), .A3(n8514), .A4(n8513), .ZN(n8517)
         );
  NOR2_X1 U10079 ( .A1(n8518), .A2(n8517), .ZN(n8519) );
  NAND3_X1 U10080 ( .A1(n8521), .A2(n8520), .A3(n8519), .ZN(n8522) );
  NOR2_X1 U10081 ( .A1(n8523), .A2(n8522), .ZN(n8567) );
  AOI22_X1 U10082 ( .A1(n8526), .A2(keyinput73), .B1(n8525), .B2(keyinput62), 
        .ZN(n8524) );
  OAI221_X1 U10083 ( .B1(n8526), .B2(keyinput73), .C1(n8525), .C2(keyinput62), 
        .A(n8524), .ZN(n8536) );
  INV_X1 U10084 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9784) );
  AOI22_X1 U10085 ( .A1(n6670), .A2(keyinput10), .B1(n9784), .B2(keyinput97), 
        .ZN(n8527) );
  OAI221_X1 U10086 ( .B1(n6670), .B2(keyinput10), .C1(n9784), .C2(keyinput97), 
        .A(n8527), .ZN(n8535) );
  AOI22_X1 U10087 ( .A1(n6123), .A2(keyinput106), .B1(n8529), .B2(keyinput52), 
        .ZN(n8528) );
  OAI221_X1 U10088 ( .B1(n6123), .B2(keyinput106), .C1(n8529), .C2(keyinput52), 
        .A(n8528), .ZN(n8534) );
  AOI22_X1 U10089 ( .A1(n8532), .A2(keyinput110), .B1(keyinput46), .B2(n8531), 
        .ZN(n8530) );
  OAI221_X1 U10090 ( .B1(n8532), .B2(keyinput110), .C1(n8531), .C2(keyinput46), 
        .A(n8530), .ZN(n8533) );
  NOR4_X1 U10091 ( .A1(n8536), .A2(n8535), .A3(n8534), .A4(n8533), .ZN(n8566)
         );
  AOI22_X1 U10092 ( .A1(n6861), .A2(keyinput16), .B1(keyinput17), .B2(n6985), 
        .ZN(n8537) );
  OAI221_X1 U10093 ( .B1(n6861), .B2(keyinput16), .C1(n6985), .C2(keyinput17), 
        .A(n8537), .ZN(n8545) );
  INV_X1 U10094 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10045) );
  AOI22_X1 U10095 ( .A1(n10045), .A2(keyinput103), .B1(keyinput120), .B2(n8539), .ZN(n8538) );
  OAI221_X1 U10096 ( .B1(n10045), .B2(keyinput103), .C1(n8539), .C2(
        keyinput120), .A(n8538), .ZN(n8544) );
  AOI22_X1 U10097 ( .A1(n8542), .A2(keyinput86), .B1(n8541), .B2(keyinput60), 
        .ZN(n8540) );
  OAI221_X1 U10098 ( .B1(n8542), .B2(keyinput86), .C1(n8541), .C2(keyinput60), 
        .A(n8540), .ZN(n8543) );
  NOR3_X1 U10099 ( .A1(n8545), .A2(n8544), .A3(n8543), .ZN(n8564) );
  AOI22_X1 U10100 ( .A1(n8547), .A2(keyinput28), .B1(n6775), .B2(keyinput6), 
        .ZN(n8546) );
  OAI221_X1 U10101 ( .B1(n8547), .B2(keyinput28), .C1(n6775), .C2(keyinput6), 
        .A(n8546), .ZN(n8550) );
  AOI22_X1 U10102 ( .A1(n6643), .A2(keyinput89), .B1(keyinput67), .B2(n9480), 
        .ZN(n8548) );
  OAI221_X1 U10103 ( .B1(n6643), .B2(keyinput89), .C1(n9480), .C2(keyinput67), 
        .A(n8548), .ZN(n8549) );
  NOR2_X1 U10104 ( .A1(n8550), .A2(n8549), .ZN(n8563) );
  AOI22_X1 U10105 ( .A1(n8552), .A2(keyinput38), .B1(keyinput59), .B2(n6039), 
        .ZN(n8551) );
  OAI221_X1 U10106 ( .B1(n8552), .B2(keyinput38), .C1(n6039), .C2(keyinput59), 
        .A(n8551), .ZN(n8555) );
  INV_X1 U10107 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10312) );
  AOI22_X1 U10108 ( .A1(n10312), .A2(keyinput72), .B1(n6749), .B2(keyinput30), 
        .ZN(n8553) );
  OAI221_X1 U10109 ( .B1(n10312), .B2(keyinput72), .C1(n6749), .C2(keyinput30), 
        .A(n8553), .ZN(n8554) );
  NOR2_X1 U10110 ( .A1(n8555), .A2(n8554), .ZN(n8562) );
  AOI22_X1 U10111 ( .A1(n8557), .A2(keyinput7), .B1(keyinput104), .B2(n6598), 
        .ZN(n8556) );
  OAI221_X1 U10112 ( .B1(n8557), .B2(keyinput7), .C1(n6598), .C2(keyinput104), 
        .A(n8556), .ZN(n8560) );
  INV_X1 U10113 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9649) );
  INV_X1 U10114 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9885) );
  AOI22_X1 U10115 ( .A1(n9649), .A2(keyinput80), .B1(keyinput44), .B2(n9885), 
        .ZN(n8558) );
  OAI221_X1 U10116 ( .B1(n9649), .B2(keyinput80), .C1(n9885), .C2(keyinput44), 
        .A(n8558), .ZN(n8559) );
  NOR2_X1 U10117 ( .A1(n8560), .A2(n8559), .ZN(n8561) );
  AND4_X1 U10118 ( .A1(n8564), .A2(n8563), .A3(n8562), .A4(n8561), .ZN(n8565)
         );
  NAND4_X1 U10119 ( .A1(n8568), .A2(n8567), .A3(n8566), .A4(n8565), .ZN(n8663)
         );
  AOI22_X1 U10120 ( .A1(n10185), .A2(keyinput92), .B1(keyinput55), .B2(n8570), 
        .ZN(n8569) );
  OAI221_X1 U10121 ( .B1(n10185), .B2(keyinput92), .C1(n8570), .C2(keyinput55), 
        .A(n8569), .ZN(n8577) );
  INV_X1 U10122 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10050) );
  AOI22_X1 U10123 ( .A1(n6631), .A2(keyinput19), .B1(n10050), .B2(keyinput107), 
        .ZN(n8571) );
  OAI221_X1 U10124 ( .B1(n6631), .B2(keyinput19), .C1(n10050), .C2(keyinput107), .A(n8571), .ZN(n8576) );
  AOI22_X1 U10125 ( .A1(n5119), .A2(keyinput2), .B1(keyinput87), .B2(n5084), 
        .ZN(n8572) );
  OAI221_X1 U10126 ( .B1(n5119), .B2(keyinput2), .C1(n5084), .C2(keyinput87), 
        .A(n8572), .ZN(n8575) );
  AOI22_X1 U10127 ( .A1(n5918), .A2(keyinput83), .B1(n6308), .B2(keyinput11), 
        .ZN(n8573) );
  OAI221_X1 U10128 ( .B1(n5918), .B2(keyinput83), .C1(n6308), .C2(keyinput11), 
        .A(n8573), .ZN(n8574) );
  NOR4_X1 U10129 ( .A1(n8577), .A2(n8576), .A3(n8575), .A4(n8574), .ZN(n8617)
         );
  INV_X1 U10130 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9916) );
  AOI22_X1 U10131 ( .A1(n9128), .A2(keyinput56), .B1(keyinput9), .B2(n9916), 
        .ZN(n8578) );
  OAI221_X1 U10132 ( .B1(n9128), .B2(keyinput56), .C1(n9916), .C2(keyinput9), 
        .A(n8578), .ZN(n8587) );
  AOI22_X1 U10133 ( .A1(n4715), .A2(keyinput35), .B1(keyinput101), .B2(n4798), 
        .ZN(n8579) );
  OAI221_X1 U10134 ( .B1(n4715), .B2(keyinput35), .C1(n4798), .C2(keyinput101), 
        .A(n8579), .ZN(n8586) );
  AOI22_X1 U10135 ( .A1(n9745), .A2(keyinput109), .B1(keyinput88), .B2(n9884), 
        .ZN(n8580) );
  OAI221_X1 U10136 ( .B1(n9745), .B2(keyinput109), .C1(n9884), .C2(keyinput88), 
        .A(n8580), .ZN(n8585) );
  AOI22_X1 U10137 ( .A1(n8583), .A2(keyinput31), .B1(n8582), .B2(keyinput51), 
        .ZN(n8581) );
  OAI221_X1 U10138 ( .B1(n8583), .B2(keyinput31), .C1(n8582), .C2(keyinput51), 
        .A(n8581), .ZN(n8584) );
  NOR4_X1 U10139 ( .A1(n8587), .A2(n8586), .A3(n8585), .A4(n8584), .ZN(n8616)
         );
  AOI22_X1 U10140 ( .A1(n8590), .A2(keyinput96), .B1(keyinput66), .B2(n8589), 
        .ZN(n8588) );
  OAI221_X1 U10141 ( .B1(n8590), .B2(keyinput96), .C1(n8589), .C2(keyinput66), 
        .A(n8588), .ZN(n8600) );
  INV_X1 U10142 ( .A(P2_WR_REG_SCAN_IN), .ZN(n8592) );
  AOI22_X1 U10143 ( .A1(n8593), .A2(keyinput105), .B1(keyinput48), .B2(n8592), 
        .ZN(n8591) );
  OAI221_X1 U10144 ( .B1(n8593), .B2(keyinput105), .C1(n8592), .C2(keyinput48), 
        .A(n8591), .ZN(n8599) );
  AOI22_X1 U10145 ( .A1(n5459), .A2(keyinput32), .B1(keyinput23), .B2(n8670), 
        .ZN(n8594) );
  OAI221_X1 U10146 ( .B1(n5459), .B2(keyinput32), .C1(n8670), .C2(keyinput23), 
        .A(n8594), .ZN(n8598) );
  AOI22_X1 U10147 ( .A1(n8596), .A2(keyinput124), .B1(n5439), .B2(keyinput100), 
        .ZN(n8595) );
  OAI221_X1 U10148 ( .B1(n8596), .B2(keyinput124), .C1(n5439), .C2(keyinput100), .A(n8595), .ZN(n8597) );
  NOR4_X1 U10149 ( .A1(n8600), .A2(n8599), .A3(n8598), .A4(n8597), .ZN(n8615)
         );
  AOI22_X1 U10150 ( .A1(n8414), .A2(keyinput39), .B1(n9798), .B2(keyinput3), 
        .ZN(n8601) );
  OAI221_X1 U10151 ( .B1(n8414), .B2(keyinput39), .C1(n9798), .C2(keyinput3), 
        .A(n8601), .ZN(n8613) );
  INV_X1 U10152 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8603) );
  AOI22_X1 U10153 ( .A1(n8604), .A2(keyinput71), .B1(n8603), .B2(keyinput127), 
        .ZN(n8602) );
  OAI221_X1 U10154 ( .B1(n8604), .B2(keyinput71), .C1(n8603), .C2(keyinput127), 
        .A(n8602), .ZN(n8612) );
  AOI22_X1 U10155 ( .A1(n8607), .A2(keyinput13), .B1(n8606), .B2(keyinput29), 
        .ZN(n8605) );
  OAI221_X1 U10156 ( .B1(n8607), .B2(keyinput13), .C1(n8606), .C2(keyinput29), 
        .A(n8605), .ZN(n8611) );
  INV_X1 U10157 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10179) );
  AOI22_X1 U10158 ( .A1(n10179), .A2(keyinput111), .B1(n8609), .B2(keyinput77), 
        .ZN(n8608) );
  OAI221_X1 U10159 ( .B1(n10179), .B2(keyinput111), .C1(n8609), .C2(keyinput77), .A(n8608), .ZN(n8610) );
  NOR4_X1 U10160 ( .A1(n8613), .A2(n8612), .A3(n8611), .A4(n8610), .ZN(n8614)
         );
  NAND4_X1 U10161 ( .A1(n8617), .A2(n8616), .A3(n8615), .A4(n8614), .ZN(n8662)
         );
  AOI22_X1 U10162 ( .A1(n8620), .A2(keyinput41), .B1(keyinput54), .B2(n8619), 
        .ZN(n8618) );
  OAI221_X1 U10163 ( .B1(n8620), .B2(keyinput41), .C1(n8619), .C2(keyinput54), 
        .A(n8618), .ZN(n8630) );
  AOI22_X1 U10164 ( .A1(n8623), .A2(keyinput27), .B1(n8622), .B2(keyinput82), 
        .ZN(n8621) );
  OAI221_X1 U10165 ( .B1(n8623), .B2(keyinput27), .C1(n8622), .C2(keyinput82), 
        .A(n8621), .ZN(n8629) );
  INV_X1 U10166 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n8625) );
  INV_X1 U10167 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10043) );
  AOI22_X1 U10168 ( .A1(n8625), .A2(keyinput126), .B1(n10043), .B2(keyinput15), 
        .ZN(n8624) );
  OAI221_X1 U10169 ( .B1(n8625), .B2(keyinput126), .C1(n10043), .C2(keyinput15), .A(n8624), .ZN(n8628) );
  AOI22_X1 U10170 ( .A1(P2_U3152), .A2(keyinput74), .B1(keyinput58), .B2(
        n10183), .ZN(n8626) );
  OAI221_X1 U10171 ( .B1(P2_U3152), .B2(keyinput74), .C1(n10183), .C2(
        keyinput58), .A(n8626), .ZN(n8627) );
  NOR4_X1 U10172 ( .A1(n8630), .A2(n8629), .A3(n8628), .A4(n8627), .ZN(n8660)
         );
  INV_X1 U10173 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10046) );
  AOI22_X1 U10174 ( .A1(n8632), .A2(keyinput123), .B1(n10046), .B2(keyinput119), .ZN(n8631) );
  OAI221_X1 U10175 ( .B1(n8632), .B2(keyinput123), .C1(n10046), .C2(
        keyinput119), .A(n8631), .ZN(n8643) );
  INV_X1 U10176 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10044) );
  AOI22_X1 U10177 ( .A1(n10044), .A2(keyinput50), .B1(keyinput20), .B2(n8634), 
        .ZN(n8633) );
  OAI221_X1 U10178 ( .B1(n10044), .B2(keyinput50), .C1(n8634), .C2(keyinput20), 
        .A(n8633), .ZN(n8642) );
  AOI22_X1 U10179 ( .A1(n5085), .A2(keyinput112), .B1(n8636), .B2(keyinput113), 
        .ZN(n8635) );
  OAI221_X1 U10180 ( .B1(n5085), .B2(keyinput112), .C1(n8636), .C2(keyinput113), .A(n8635), .ZN(n8641) );
  AOI22_X1 U10181 ( .A1(n8639), .A2(keyinput108), .B1(keyinput76), .B2(n8638), 
        .ZN(n8637) );
  OAI221_X1 U10182 ( .B1(n8639), .B2(keyinput108), .C1(n8638), .C2(keyinput76), 
        .A(n8637), .ZN(n8640) );
  NOR4_X1 U10183 ( .A1(n8643), .A2(n8642), .A3(n8641), .A4(n8640), .ZN(n8659)
         );
  INV_X1 U10184 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8645) );
  AOI22_X1 U10185 ( .A1(n8415), .A2(keyinput25), .B1(n8645), .B2(keyinput75), 
        .ZN(n8644) );
  OAI221_X1 U10186 ( .B1(n8415), .B2(keyinput25), .C1(n8645), .C2(keyinput75), 
        .A(n8644), .ZN(n8657) );
  INV_X1 U10187 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10042) );
  AOI22_X1 U10188 ( .A1(n10042), .A2(keyinput1), .B1(keyinput63), .B2(n8647), 
        .ZN(n8646) );
  OAI221_X1 U10189 ( .B1(n10042), .B2(keyinput1), .C1(n8647), .C2(keyinput63), 
        .A(n8646), .ZN(n8656) );
  AOI22_X1 U10190 ( .A1(n8650), .A2(keyinput12), .B1(keyinput45), .B2(n8649), 
        .ZN(n8648) );
  OAI221_X1 U10191 ( .B1(n8650), .B2(keyinput12), .C1(n8649), .C2(keyinput45), 
        .A(n8648), .ZN(n8655) );
  AOI22_X1 U10192 ( .A1(n8653), .A2(keyinput115), .B1(keyinput26), .B2(n8652), 
        .ZN(n8651) );
  OAI221_X1 U10193 ( .B1(n8653), .B2(keyinput115), .C1(n8652), .C2(keyinput26), 
        .A(n8651), .ZN(n8654) );
  NOR4_X1 U10194 ( .A1(n8657), .A2(n8656), .A3(n8655), .A4(n8654), .ZN(n8658)
         );
  NAND3_X1 U10195 ( .A1(n8660), .A2(n8659), .A3(n8658), .ZN(n8661) );
  OR3_X1 U10196 ( .A1(n8663), .A2(n8662), .A3(n8661), .ZN(n8664) );
  XNOR2_X1 U10197 ( .A(n8665), .B(n8664), .ZN(n8666) );
  XNOR2_X1 U10198 ( .A(n8667), .B(n8666), .ZN(P2_U3265) );
  NAND2_X1 U10199 ( .A1(n8134), .A2(n4550), .ZN(n8900) );
  NAND3_X1 U10200 ( .A1(n8900), .A2(n6504), .A3(n8899), .ZN(n8673) );
  OAI21_X1 U10201 ( .B1(n8881), .B2(n8670), .A(n8669), .ZN(n8671) );
  AOI21_X1 U10202 ( .B1(n8134), .B2(n10161), .A(n8671), .ZN(n8672) );
  NAND2_X1 U10203 ( .A1(n8673), .A2(n8672), .ZN(P2_U3266) );
  OAI21_X1 U10204 ( .B1(n8676), .B2(n8675), .A(n8674), .ZN(n8677) );
  INV_X1 U10205 ( .A(n8677), .ZN(n8919) );
  XNOR2_X1 U10206 ( .A(n8679), .B(n8678), .ZN(n8680) );
  OAI222_X1 U10207 ( .A1(n8858), .A2(n8682), .B1(n8856), .B2(n8681), .C1(n8854), .C2(n8680), .ZN(n8910) );
  INV_X1 U10208 ( .A(n8683), .ZN(n8684) );
  AOI21_X1 U10209 ( .B1(n8685), .B2(n8695), .A(n8684), .ZN(n8911) );
  NAND2_X1 U10210 ( .A1(n8911), .A2(n6504), .ZN(n8688) );
  AOI22_X1 U10211 ( .A1(P2_REG2_REG_28__SCAN_IN), .A2(n4392), .B1(n8686), .B2(
        n10159), .ZN(n8687) );
  OAI211_X1 U10212 ( .C1(n8689), .C2(n8869), .A(n8688), .B(n8687), .ZN(n8690)
         );
  AOI21_X1 U10213 ( .B1(n8910), .B2(n8881), .A(n8690), .ZN(n8691) );
  OAI21_X1 U10214 ( .B1(n8919), .B2(n8874), .A(n8691), .ZN(P2_U3268) );
  OAI21_X1 U10215 ( .B1(n8693), .B2(n8701), .A(n8692), .ZN(n8694) );
  INV_X1 U10216 ( .A(n8694), .ZN(n8924) );
  INV_X1 U10217 ( .A(n8716), .ZN(n8697) );
  INV_X1 U10218 ( .A(n8695), .ZN(n8696) );
  AOI21_X1 U10219 ( .B1(n8920), .B2(n8697), .A(n8696), .ZN(n8921) );
  AOI22_X1 U10220 ( .A1(n4392), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8698), .B2(
        n10159), .ZN(n8699) );
  OAI21_X1 U10221 ( .B1(n8216), .B2(n8869), .A(n8699), .ZN(n8705) );
  XOR2_X1 U10222 ( .A(n8701), .B(n8700), .Z(n8703) );
  AOI222_X1 U10223 ( .A1(n10156), .A2(n8703), .B1(n8702), .B2(n8879), .C1(
        n8728), .C2(n8877), .ZN(n8923) );
  NOR2_X1 U10224 ( .A1(n8923), .A2(n4392), .ZN(n8704) );
  AOI211_X1 U10225 ( .C1(n8921), .C2(n6504), .A(n8705), .B(n8704), .ZN(n8706)
         );
  OAI21_X1 U10226 ( .B1(n8924), .B2(n8874), .A(n8706), .ZN(P2_U3269) );
  OAI21_X1 U10227 ( .B1(n8709), .B2(n8708), .A(n8707), .ZN(n8710) );
  INV_X1 U10228 ( .A(n8710), .ZN(n8929) );
  AOI22_X1 U10229 ( .A1(n8926), .A2(n10161), .B1(n4392), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8721) );
  OAI21_X1 U10230 ( .B1(n8713), .B2(n8712), .A(n8711), .ZN(n8715) );
  AOI222_X1 U10231 ( .A1(n10156), .A2(n8715), .B1(n8714), .B2(n8879), .C1(
        n8751), .C2(n8877), .ZN(n8928) );
  AOI211_X1 U10232 ( .C1(n8926), .C2(n8731), .A(n10248), .B(n8716), .ZN(n8925)
         );
  NAND2_X1 U10233 ( .A1(n8925), .A2(n8865), .ZN(n8717) );
  OAI211_X1 U10234 ( .C1(n8888), .C2(n8718), .A(n8928), .B(n8717), .ZN(n8719)
         );
  NAND2_X1 U10235 ( .A1(n8719), .A2(n8881), .ZN(n8720) );
  OAI211_X1 U10236 ( .C1(n8929), .C2(n8874), .A(n8721), .B(n8720), .ZN(
        P2_U3270) );
  OAI21_X1 U10237 ( .B1(n8723), .B2(n8725), .A(n8722), .ZN(n8930) );
  INV_X1 U10238 ( .A(n8930), .ZN(n8739) );
  AOI22_X1 U10239 ( .A1(n8724), .A2(n10161), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n4392), .ZN(n8738) );
  XNOR2_X1 U10240 ( .A(n8726), .B(n8725), .ZN(n8727) );
  AOI222_X1 U10241 ( .A1(n8729), .A2(n8877), .B1(n8728), .B2(n8879), .C1(
        n10156), .C2(n8727), .ZN(n8933) );
  INV_X1 U10242 ( .A(n8933), .ZN(n8736) );
  INV_X1 U10243 ( .A(n8730), .ZN(n8741) );
  OAI211_X1 U10244 ( .C1(n8732), .C2(n8741), .A(n10215), .B(n8731), .ZN(n8931)
         );
  OAI22_X1 U10245 ( .A1(n8931), .A2(n8734), .B1(n8888), .B2(n8733), .ZN(n8735)
         );
  OAI21_X1 U10246 ( .B1(n8736), .B2(n8735), .A(n8881), .ZN(n8737) );
  OAI211_X1 U10247 ( .C1(n8739), .C2(n8874), .A(n8738), .B(n8737), .ZN(
        P2_U3271) );
  XNOR2_X1 U10248 ( .A(n8740), .B(n8748), .ZN(n8939) );
  INV_X1 U10249 ( .A(n8768), .ZN(n8742) );
  AOI21_X1 U10250 ( .B1(n8935), .B2(n8742), .A(n8741), .ZN(n8936) );
  AOI22_X1 U10251 ( .A1(n4392), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8743), .B2(
        n10159), .ZN(n8744) );
  OAI21_X1 U10252 ( .B1(n8745), .B2(n8869), .A(n8744), .ZN(n8753) );
  INV_X1 U10253 ( .A(n8746), .ZN(n8747) );
  NOR2_X1 U10254 ( .A1(n8761), .A2(n8747), .ZN(n8749) );
  XNOR2_X1 U10255 ( .A(n8749), .B(n8748), .ZN(n8750) );
  AOI222_X1 U10256 ( .A1(n8779), .A2(n8877), .B1(n8751), .B2(n8879), .C1(
        n10156), .C2(n8750), .ZN(n8938) );
  NOR2_X1 U10257 ( .A1(n8938), .A2(n4392), .ZN(n8752) );
  AOI211_X1 U10258 ( .C1(n8936), .C2(n6504), .A(n8753), .B(n8752), .ZN(n8754)
         );
  OAI21_X1 U10259 ( .B1(n8939), .B2(n8874), .A(n8754), .ZN(P2_U3272) );
  OAI21_X1 U10260 ( .B1(n8755), .B2(n8757), .A(n8756), .ZN(n8944) );
  NOR2_X1 U10261 ( .A1(n8759), .A2(n8758), .ZN(n8760) );
  OR2_X1 U10262 ( .A1(n8761), .A2(n8760), .ZN(n8763) );
  AOI21_X1 U10263 ( .B1(n8763), .B2(n10156), .A(n8762), .ZN(n8943) );
  INV_X1 U10264 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8765) );
  OAI22_X1 U10265 ( .A1(n8881), .A2(n8765), .B1(n8764), .B2(n8888), .ZN(n8766)
         );
  AOI21_X1 U10266 ( .B1(n8940), .B2(n10161), .A(n8766), .ZN(n8770) );
  AND2_X1 U10267 ( .A1(n8940), .A2(n8947), .ZN(n8767) );
  NOR2_X1 U10268 ( .A1(n8768), .A2(n8767), .ZN(n8941) );
  NAND2_X1 U10269 ( .A1(n8941), .A2(n6504), .ZN(n8769) );
  OAI211_X1 U10270 ( .C1(n8943), .C2(n4392), .A(n8770), .B(n8769), .ZN(n8771)
         );
  INV_X1 U10271 ( .A(n8771), .ZN(n8772) );
  OAI21_X1 U10272 ( .B1(n8944), .B2(n8874), .A(n8772), .ZN(P2_U3273) );
  XNOR2_X1 U10273 ( .A(n8774), .B(n8773), .ZN(n8951) );
  NAND2_X1 U10274 ( .A1(n8793), .A2(n8775), .ZN(n8777) );
  XNOR2_X1 U10275 ( .A(n8777), .B(n8776), .ZN(n8778) );
  AOI222_X1 U10276 ( .A1(n8804), .A2(n8877), .B1(n8779), .B2(n8879), .C1(
        n10156), .C2(n8778), .ZN(n8950) );
  INV_X1 U10277 ( .A(n8950), .ZN(n8786) );
  NOR2_X1 U10278 ( .A1(n4541), .A2(n4405), .ZN(n8945) );
  INV_X1 U10279 ( .A(n8947), .ZN(n8781) );
  NOR3_X1 U10280 ( .A1(n8945), .A2(n8781), .A3(n8780), .ZN(n8785) );
  AOI22_X1 U10281 ( .A1(n4392), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8782), .B2(
        n10159), .ZN(n8783) );
  OAI21_X1 U10282 ( .B1(n4541), .B2(n8869), .A(n8783), .ZN(n8784) );
  AOI211_X1 U10283 ( .C1(n8786), .C2(n8881), .A(n8785), .B(n8784), .ZN(n8787)
         );
  OAI21_X1 U10284 ( .B1(n8951), .B2(n8874), .A(n8787), .ZN(P2_U3274) );
  XNOR2_X1 U10285 ( .A(n8788), .B(n8794), .ZN(n8956) );
  AOI21_X1 U10286 ( .B1(n8952), .B2(n4545), .A(n4405), .ZN(n8953) );
  INV_X1 U10287 ( .A(n8789), .ZN(n8790) );
  AOI22_X1 U10288 ( .A1(n4392), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8790), .B2(
        n10159), .ZN(n8791) );
  OAI21_X1 U10289 ( .B1(n8792), .B2(n8869), .A(n8791), .ZN(n8799) );
  OAI21_X1 U10290 ( .B1(n4419), .B2(n8794), .A(n8793), .ZN(n8797) );
  AOI222_X1 U10291 ( .A1(n10156), .A2(n8797), .B1(n8796), .B2(n8879), .C1(
        n8795), .C2(n8877), .ZN(n8955) );
  NOR2_X1 U10292 ( .A1(n8955), .A2(n4392), .ZN(n8798) );
  AOI211_X1 U10293 ( .C1(n8953), .C2(n6504), .A(n8799), .B(n8798), .ZN(n8800)
         );
  OAI21_X1 U10294 ( .B1(n8956), .B2(n8874), .A(n8800), .ZN(P2_U3275) );
  NAND2_X1 U10295 ( .A1(n8823), .A2(n8801), .ZN(n8802) );
  XNOR2_X1 U10296 ( .A(n8802), .B(n8805), .ZN(n8803) );
  AOI222_X1 U10297 ( .A1(n8842), .A2(n8877), .B1(n8804), .B2(n8879), .C1(
        n10156), .C2(n8803), .ZN(n8961) );
  INV_X1 U10298 ( .A(n8963), .ZN(n8807) );
  NAND2_X1 U10299 ( .A1(n8806), .A2(n8805), .ZN(n8957) );
  NAND3_X1 U10300 ( .A1(n8807), .A2(n10172), .A3(n8957), .ZN(n8815) );
  AOI21_X1 U10301 ( .B1(n8958), .B2(n8809), .A(n8808), .ZN(n8959) );
  NOR2_X1 U10302 ( .A1(n8810), .A2(n8869), .ZN(n8813) );
  OAI22_X1 U10303 ( .A1(n8881), .A2(n8491), .B1(n8811), .B2(n8888), .ZN(n8812)
         );
  AOI211_X1 U10304 ( .C1(n8959), .C2(n6504), .A(n8813), .B(n8812), .ZN(n8814)
         );
  OAI211_X1 U10305 ( .C1(n4392), .C2(n8961), .A(n8815), .B(n8814), .ZN(
        P2_U3276) );
  XOR2_X1 U10306 ( .A(n8816), .B(n8825), .Z(n8968) );
  INV_X1 U10307 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8819) );
  INV_X1 U10308 ( .A(n8817), .ZN(n8818) );
  OAI22_X1 U10309 ( .A1(n8881), .A2(n8819), .B1(n8818), .B2(n8888), .ZN(n8830)
         );
  XNOR2_X1 U10310 ( .A(n8820), .B(n8834), .ZN(n8821) );
  NOR2_X1 U10311 ( .A1(n8821), .A2(n10248), .ZN(n8965) );
  INV_X1 U10312 ( .A(n8823), .ZN(n8824) );
  AOI21_X1 U10313 ( .B1(n8822), .B2(n8825), .A(n8824), .ZN(n8826) );
  OAI222_X1 U10314 ( .A1(n8858), .A2(n8827), .B1(n8856), .B2(n8859), .C1(n8854), .C2(n8826), .ZN(n8964) );
  AOI21_X1 U10315 ( .B1(n8965), .B2(n8865), .A(n8964), .ZN(n8828) );
  NOR2_X1 U10316 ( .A1(n8828), .A2(n4392), .ZN(n8829) );
  AOI211_X1 U10317 ( .C1(n10161), .C2(n8966), .A(n8830), .B(n8829), .ZN(n8831)
         );
  OAI21_X1 U10318 ( .B1(n8968), .B2(n8874), .A(n8831), .ZN(P2_U3277) );
  XNOR2_X1 U10319 ( .A(n8833), .B(n8832), .ZN(n8973) );
  INV_X1 U10320 ( .A(n8863), .ZN(n8835) );
  AOI21_X1 U10321 ( .B1(n8969), .B2(n8835), .A(n8834), .ZN(n8970) );
  AOI22_X1 U10322 ( .A1(n4392), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8836), .B2(
        n10159), .ZN(n8837) );
  OAI21_X1 U10323 ( .B1(n8838), .B2(n8869), .A(n8837), .ZN(n8845) );
  XNOR2_X1 U10324 ( .A(n8840), .B(n8839), .ZN(n8843) );
  AOI222_X1 U10325 ( .A1(n10156), .A2(n8843), .B1(n8842), .B2(n8879), .C1(
        n8841), .C2(n8877), .ZN(n8972) );
  NOR2_X1 U10326 ( .A1(n8972), .A2(n4392), .ZN(n8844) );
  AOI211_X1 U10327 ( .C1(n8970), .C2(n6504), .A(n8845), .B(n8844), .ZN(n8846)
         );
  OAI21_X1 U10328 ( .B1(n8973), .B2(n8874), .A(n8846), .ZN(P2_U3278) );
  OAI21_X1 U10329 ( .B1(n8849), .B2(n8848), .A(n8847), .ZN(n8850) );
  INV_X1 U10330 ( .A(n8850), .ZN(n8978) );
  AOI21_X1 U10331 ( .B1(n8853), .B2(n8852), .A(n8851), .ZN(n8855) );
  NOR3_X1 U10332 ( .A1(n4453), .A2(n8855), .A3(n8854), .ZN(n8861) );
  OAI22_X1 U10333 ( .A1(n8859), .A2(n8858), .B1(n8857), .B2(n8856), .ZN(n8860)
         );
  NOR2_X1 U10334 ( .A1(n8861), .A2(n8860), .ZN(n8977) );
  INV_X1 U10335 ( .A(n8862), .ZN(n8864) );
  AOI211_X1 U10336 ( .C1(n8975), .C2(n8864), .A(n10248), .B(n8863), .ZN(n8974)
         );
  NAND2_X1 U10337 ( .A1(n8974), .A2(n8865), .ZN(n8866) );
  OAI211_X1 U10338 ( .C1(n8888), .C2(n8867), .A(n8977), .B(n8866), .ZN(n8872)
         );
  OAI22_X1 U10339 ( .A1(n8870), .A2(n8869), .B1(n8868), .B2(n8881), .ZN(n8871)
         );
  AOI21_X1 U10340 ( .B1(n8872), .B2(n8881), .A(n8871), .ZN(n8873) );
  OAI21_X1 U10341 ( .B1(n8978), .B2(n8874), .A(n8873), .ZN(P2_U3279) );
  OAI21_X1 U10342 ( .B1(n8893), .B2(n8876), .A(n8875), .ZN(n8880) );
  AOI222_X1 U10343 ( .A1(n10156), .A2(n8880), .B1(n10126), .B2(n8879), .C1(
        n8878), .C2(n8877), .ZN(n10220) );
  MUX2_X1 U10344 ( .A(n8882), .B(n10220), .S(n8881), .Z(n8896) );
  AND2_X1 U10345 ( .A1(n8883), .A2(n10214), .ZN(n8884) );
  NOR2_X1 U10346 ( .A1(n8885), .A2(n8884), .ZN(n10216) );
  NAND2_X1 U10347 ( .A1(n6504), .A2(n10216), .ZN(n8886) );
  OAI21_X1 U10348 ( .B1(n8888), .B2(n8887), .A(n8886), .ZN(n8889) );
  AOI21_X1 U10349 ( .B1(n10161), .B2(n10214), .A(n8889), .ZN(n8895) );
  NAND2_X1 U10350 ( .A1(n8892), .A2(n8893), .ZN(n10217) );
  NAND3_X1 U10351 ( .A1(n8891), .A2(n10217), .A3(n10172), .ZN(n8894) );
  NAND3_X1 U10352 ( .A1(n8896), .A2(n8895), .A3(n8894), .ZN(P2_U3290) );
  AOI21_X1 U10353 ( .B1(n8390), .B2(n10213), .A(n8901), .ZN(n8897) );
  OAI21_X1 U10354 ( .B1(n8898), .B2(n10248), .A(n8897), .ZN(n8995) );
  MUX2_X1 U10355 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8995), .S(n10275), .Z(
        P2_U3551) );
  NAND3_X1 U10356 ( .A1(n8900), .A2(n10215), .A3(n8899), .ZN(n8903) );
  INV_X1 U10357 ( .A(n8901), .ZN(n8902) );
  OAI211_X1 U10358 ( .C1(n8904), .C2(n10255), .A(n8903), .B(n8902), .ZN(n8996)
         );
  INV_X2 U10359 ( .A(n10273), .ZN(n10275) );
  MUX2_X1 U10360 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8996), .S(n10275), .Z(
        P2_U3550) );
  MUX2_X1 U10361 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8997), .S(n10275), .Z(
        P2_U3549) );
  INV_X1 U10362 ( .A(n8910), .ZN(n8917) );
  INV_X1 U10363 ( .A(n8911), .ZN(n8912) );
  INV_X1 U10364 ( .A(n8913), .ZN(n8914) );
  AND2_X1 U10365 ( .A1(n8915), .A2(n8914), .ZN(n8916) );
  OAI21_X1 U10366 ( .B1(n8919), .B2(n8993), .A(n8918), .ZN(n8998) );
  MUX2_X1 U10367 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8998), .S(n10275), .Z(
        P2_U3548) );
  AOI22_X1 U10368 ( .A1(n8921), .A2(n10215), .B1(n8920), .B2(n10213), .ZN(
        n8922) );
  OAI211_X1 U10369 ( .C1(n8924), .C2(n8993), .A(n8923), .B(n8922), .ZN(n8999)
         );
  MUX2_X1 U10370 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8999), .S(n10275), .Z(
        P2_U3547) );
  AOI21_X1 U10371 ( .B1(n8926), .B2(n10213), .A(n8925), .ZN(n8927) );
  OAI211_X1 U10372 ( .C1(n8929), .C2(n8993), .A(n8928), .B(n8927), .ZN(n9000)
         );
  MUX2_X1 U10373 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9000), .S(n10275), .Z(
        P2_U3546) );
  NAND2_X1 U10374 ( .A1(n8930), .A2(n10259), .ZN(n8934) );
  NAND4_X1 U10375 ( .A1(n8934), .A2(n8933), .A3(n8932), .A4(n8931), .ZN(n9001)
         );
  MUX2_X1 U10376 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9001), .S(n10275), .Z(
        P2_U3545) );
  AOI22_X1 U10377 ( .A1(n8936), .A2(n10215), .B1(n8935), .B2(n10213), .ZN(
        n8937) );
  OAI211_X1 U10378 ( .C1(n8939), .C2(n8993), .A(n8938), .B(n8937), .ZN(n9002)
         );
  MUX2_X1 U10379 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9002), .S(n10275), .Z(
        P2_U3544) );
  AOI22_X1 U10380 ( .A1(n8941), .A2(n10215), .B1(n8940), .B2(n10213), .ZN(
        n8942) );
  OAI211_X1 U10381 ( .C1(n8944), .C2(n8993), .A(n8943), .B(n8942), .ZN(n9003)
         );
  MUX2_X1 U10382 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9003), .S(n10275), .Z(
        P2_U3543) );
  NOR2_X1 U10383 ( .A1(n8945), .A2(n10248), .ZN(n8948) );
  AOI22_X1 U10384 ( .A1(n8948), .A2(n8947), .B1(n8946), .B2(n10213), .ZN(n8949) );
  OAI211_X1 U10385 ( .C1(n8951), .C2(n8993), .A(n8950), .B(n8949), .ZN(n9004)
         );
  MUX2_X1 U10386 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9004), .S(n10275), .Z(
        P2_U3542) );
  AOI22_X1 U10387 ( .A1(n8953), .A2(n10215), .B1(n8952), .B2(n10213), .ZN(
        n8954) );
  OAI211_X1 U10388 ( .C1(n8956), .C2(n8993), .A(n8955), .B(n8954), .ZN(n9005)
         );
  MUX2_X1 U10389 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9005), .S(n10275), .Z(
        P2_U3541) );
  NAND2_X1 U10390 ( .A1(n8957), .A2(n10259), .ZN(n8962) );
  AOI22_X1 U10391 ( .A1(n8959), .A2(n10215), .B1(n8958), .B2(n10213), .ZN(
        n8960) );
  OAI211_X1 U10392 ( .C1(n8963), .C2(n8962), .A(n8961), .B(n8960), .ZN(n9006)
         );
  MUX2_X1 U10393 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9006), .S(n10275), .Z(
        P2_U3540) );
  AOI211_X1 U10394 ( .C1(n8966), .C2(n10213), .A(n8965), .B(n8964), .ZN(n8967)
         );
  OAI21_X1 U10395 ( .B1(n8968), .B2(n8993), .A(n8967), .ZN(n9007) );
  MUX2_X1 U10396 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9007), .S(n10275), .Z(
        P2_U3539) );
  AOI22_X1 U10397 ( .A1(n8970), .A2(n10215), .B1(n8969), .B2(n10213), .ZN(
        n8971) );
  OAI211_X1 U10398 ( .C1(n8973), .C2(n8993), .A(n8972), .B(n8971), .ZN(n9008)
         );
  MUX2_X1 U10399 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9008), .S(n10275), .Z(
        P2_U3538) );
  AOI21_X1 U10400 ( .B1(n8975), .B2(n10213), .A(n8974), .ZN(n8976) );
  OAI211_X1 U10401 ( .C1(n8978), .C2(n8993), .A(n8977), .B(n8976), .ZN(n9009)
         );
  MUX2_X1 U10402 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9009), .S(n10275), .Z(
        P2_U3537) );
  AOI21_X1 U10403 ( .B1(n8980), .B2(n10213), .A(n8979), .ZN(n8981) );
  OAI211_X1 U10404 ( .C1(n10228), .C2(n8983), .A(n8982), .B(n8981), .ZN(n9010)
         );
  MUX2_X1 U10405 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9010), .S(n10275), .Z(
        P2_U3536) );
  AOI22_X1 U10406 ( .A1(n8985), .A2(n10215), .B1(n8984), .B2(n10213), .ZN(
        n8986) );
  OAI211_X1 U10407 ( .C1(n8988), .C2(n8993), .A(n8987), .B(n8986), .ZN(n9011)
         );
  MUX2_X1 U10408 ( .A(n9011), .B(P2_REG1_REG_15__SCAN_IN), .S(n10273), .Z(
        P2_U3535) );
  AOI22_X1 U10409 ( .A1(n8990), .A2(n10215), .B1(n8989), .B2(n10213), .ZN(
        n8991) );
  OAI211_X1 U10410 ( .C1(n8994), .C2(n8993), .A(n8992), .B(n8991), .ZN(n9012)
         );
  MUX2_X1 U10411 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n9012), .S(n10275), .Z(
        P2_U3534) );
  MUX2_X1 U10412 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8995), .S(n4393), .Z(
        P2_U3519) );
  MUX2_X1 U10413 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8996), .S(n4393), .Z(
        P2_U3518) );
  MUX2_X1 U10414 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8998), .S(n4393), .Z(
        P2_U3516) );
  MUX2_X1 U10415 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8999), .S(n4393), .Z(
        P2_U3515) );
  MUX2_X1 U10416 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9000), .S(n4393), .Z(
        P2_U3514) );
  MUX2_X1 U10417 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9001), .S(n4393), .Z(
        P2_U3513) );
  MUX2_X1 U10418 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9002), .S(n4393), .Z(
        P2_U3512) );
  MUX2_X1 U10419 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9003), .S(n4393), .Z(
        P2_U3511) );
  MUX2_X1 U10420 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9004), .S(n4393), .Z(
        P2_U3510) );
  MUX2_X1 U10421 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9005), .S(n4393), .Z(
        P2_U3509) );
  MUX2_X1 U10422 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9006), .S(n4393), .Z(
        P2_U3508) );
  MUX2_X1 U10423 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9007), .S(n4393), .Z(
        P2_U3507) );
  MUX2_X1 U10424 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9008), .S(n4393), .Z(
        P2_U3505) );
  MUX2_X1 U10425 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9009), .S(n4393), .Z(
        P2_U3502) );
  MUX2_X1 U10426 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9010), .S(n4393), .Z(
        P2_U3499) );
  MUX2_X1 U10427 ( .A(n9011), .B(P2_REG0_REG_15__SCAN_IN), .S(n10260), .Z(
        P2_U3496) );
  MUX2_X1 U10428 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n9012), .S(n4393), .Z(
        P2_U3493) );
  NAND3_X1 U10429 ( .A1(n4506), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n9014) );
  OAI22_X1 U10430 ( .A1(n9013), .A2(n9014), .B1(n6574), .B2(n9018), .ZN(n9015)
         );
  AOI21_X1 U10431 ( .B1(n9868), .B2(n9016), .A(n9015), .ZN(n9017) );
  INV_X1 U10432 ( .A(n9017), .ZN(P2_U3327) );
  OAI222_X1 U10433 ( .A1(P2_U3152), .A2(n9022), .B1(n9021), .B2(n9020), .C1(
        n9019), .C2(n9018), .ZN(P2_U3329) );
  MUX2_X1 U10434 ( .A(n9023), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10435 ( .A1(n9024), .A2(n5709), .ZN(n9025) );
  XOR2_X1 U10436 ( .A(n9026), .B(n9025), .Z(n9033) );
  OAI22_X1 U10437 ( .A1(n9164), .A2(n9027), .B1(n9162), .B2(n9074), .ZN(n9028)
         );
  AOI211_X1 U10438 ( .C1(n9167), .C2(n9460), .A(n9029), .B(n9028), .ZN(n9032)
         );
  NAND2_X1 U10439 ( .A1(n9030), .A2(n9142), .ZN(n9031) );
  OAI211_X1 U10440 ( .C1(n9033), .C2(n9144), .A(n9032), .B(n9031), .ZN(
        P1_U3213) );
  XOR2_X1 U10441 ( .A(n9035), .B(n9034), .Z(n9040) );
  OAI22_X1 U10442 ( .A1(n9162), .A2(n9769), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9036), .ZN(n9038) );
  OAI22_X1 U10443 ( .A1(n9139), .A2(n9700), .B1(n9164), .B2(n9663), .ZN(n9037)
         );
  AOI211_X1 U10444 ( .C1(n9670), .C2(n9142), .A(n9038), .B(n9037), .ZN(n9039)
         );
  OAI21_X1 U10445 ( .B1(n9040), .B2(n9144), .A(n9039), .ZN(P1_U3217) );
  NAND2_X1 U10446 ( .A1(n9041), .A2(n9102), .ZN(n9042) );
  XOR2_X1 U10447 ( .A(n9043), .B(n9042), .Z(n9049) );
  OAI22_X1 U10448 ( .A1(n9603), .A2(n9162), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9044), .ZN(n9047) );
  INV_X1 U10449 ( .A(n9640), .ZN(n9045) );
  OAI22_X1 U10450 ( .A1(n9139), .A2(n9769), .B1(n9164), .B2(n9045), .ZN(n9046)
         );
  AOI211_X1 U10451 ( .C1(n9772), .C2(n9142), .A(n9047), .B(n9046), .ZN(n9048)
         );
  OAI21_X1 U10452 ( .B1(n9049), .B2(n9144), .A(n9048), .ZN(P1_U3221) );
  INV_X1 U10453 ( .A(n9051), .ZN(n9052) );
  AOI21_X1 U10454 ( .B1(n9053), .B2(n9050), .A(n9052), .ZN(n9061) );
  NOR2_X1 U10455 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9054), .ZN(n9975) );
  OAI22_X1 U10456 ( .A1(n9164), .A2(n9056), .B1(n9162), .B2(n9055), .ZN(n9057)
         );
  AOI211_X1 U10457 ( .C1(n9167), .C2(n9461), .A(n9975), .B(n9057), .ZN(n9060)
         );
  NAND2_X1 U10458 ( .A1(n9058), .A2(n9142), .ZN(n9059) );
  OAI211_X1 U10459 ( .C1(n9061), .C2(n9144), .A(n9060), .B(n9059), .ZN(
        P1_U3222) );
  INV_X1 U10460 ( .A(n9563), .ZN(n9840) );
  OAI21_X1 U10461 ( .B1(n9063), .B2(n9062), .A(n9147), .ZN(n9064) );
  NAND2_X1 U10462 ( .A1(n9064), .A2(n9160), .ZN(n9068) );
  AOI22_X1 U10463 ( .A1(n9600), .A2(n9167), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9065) );
  OAI21_X1 U10464 ( .B1(n9164), .B2(n9564), .A(n9065), .ZN(n9066) );
  AOI21_X1 U10465 ( .B1(n9116), .B2(n9560), .A(n9066), .ZN(n9067) );
  OAI211_X1 U10466 ( .C1(n9840), .C2(n9170), .A(n9068), .B(n9067), .ZN(
        P1_U3223) );
  INV_X1 U10467 ( .A(n9080), .ZN(n9070) );
  AOI21_X1 U10468 ( .B1(n9072), .B2(n9071), .A(n9070), .ZN(n9078) );
  OAI22_X1 U10469 ( .A1(n9162), .A2(n9721), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9073), .ZN(n9076) );
  OAI22_X1 U10470 ( .A1(n9139), .A2(n9074), .B1(n9164), .B2(n9715), .ZN(n9075)
         );
  AOI211_X1 U10471 ( .C1(n9727), .C2(n9142), .A(n9076), .B(n9075), .ZN(n9077)
         );
  OAI21_X1 U10472 ( .B1(n9078), .B2(n9144), .A(n9077), .ZN(P1_U3224) );
  NAND2_X1 U10473 ( .A1(n9080), .A2(n9079), .ZN(n9081) );
  XOR2_X1 U10474 ( .A(n9082), .B(n9081), .Z(n9087) );
  OAI22_X1 U10475 ( .A1(n9162), .A2(n9700), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9083), .ZN(n9085) );
  OAI22_X1 U10476 ( .A1(n9139), .A2(n9699), .B1(n9164), .B2(n9693), .ZN(n9084)
         );
  AOI211_X1 U10477 ( .C1(n9802), .C2(n9142), .A(n9085), .B(n9084), .ZN(n9086)
         );
  OAI21_X1 U10478 ( .B1(n9087), .B2(n9144), .A(n9086), .ZN(P1_U3226) );
  INV_X1 U10479 ( .A(n9756), .ZN(n9099) );
  INV_X1 U10480 ( .A(n9088), .ZN(n9091) );
  AOI21_X1 U10481 ( .B1(n6515), .B2(n6516), .A(n9089), .ZN(n9090) );
  OAI21_X1 U10482 ( .B1(n9091), .B2(n9090), .A(n9160), .ZN(n9098) );
  NAND2_X1 U10483 ( .A1(n9614), .A2(n9167), .ZN(n9094) );
  NAND2_X1 U10484 ( .A1(n9574), .A2(n9092), .ZN(n9093) );
  OAI211_X1 U10485 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9095), .A(n9094), .B(
        n9093), .ZN(n9096) );
  AOI21_X1 U10486 ( .B1(n9578), .B2(n9116), .A(n9096), .ZN(n9097) );
  OAI211_X1 U10487 ( .C1(n9099), .C2(n9170), .A(n9098), .B(n9097), .ZN(
        P1_U3227) );
  NAND2_X1 U10488 ( .A1(n9102), .A2(n9101), .ZN(n9103) );
  XNOR2_X1 U10489 ( .A(n9100), .B(n9103), .ZN(n9108) );
  OAI22_X1 U10490 ( .A1(n9777), .A2(n9162), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9104), .ZN(n9106) );
  OAI22_X1 U10491 ( .A1(n9139), .A2(n9776), .B1(n9164), .B2(n9648), .ZN(n9105)
         );
  AOI211_X1 U10492 ( .C1(n9657), .C2(n9142), .A(n9106), .B(n9105), .ZN(n9107)
         );
  OAI21_X1 U10493 ( .B1(n9108), .B2(n9144), .A(n9107), .ZN(P1_U3231) );
  NAND2_X1 U10494 ( .A1(n9110), .A2(n9109), .ZN(n9111) );
  XOR2_X1 U10495 ( .A(n4451), .B(n9111), .Z(n9119) );
  OAI22_X1 U10496 ( .A1(n9139), .A2(n9113), .B1(n9164), .B2(n9112), .ZN(n9114)
         );
  AOI211_X1 U10497 ( .C1(n9116), .C2(n9817), .A(n9115), .B(n9114), .ZN(n9118)
         );
  NAND2_X1 U10498 ( .A1(n9816), .A2(n9142), .ZN(n9117) );
  OAI211_X1 U10499 ( .C1(n9119), .C2(n9144), .A(n9118), .B(n9117), .ZN(
        P1_U3232) );
  AND2_X1 U10500 ( .A1(n9122), .A2(n9121), .ZN(n9124) );
  AOI21_X1 U10501 ( .B1(n9124), .B2(n9126), .A(n9123), .ZN(n9125) );
  AOI21_X1 U10502 ( .B1(n9127), .B2(n9126), .A(n9125), .ZN(n9132) );
  OAI22_X1 U10503 ( .A1(n9139), .A2(n9777), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9128), .ZN(n9130) );
  OAI22_X1 U10504 ( .A1(n9581), .A2(n9162), .B1(n9164), .B2(n9619), .ZN(n9129)
         );
  AOI211_X1 U10505 ( .C1(n9618), .C2(n9142), .A(n9130), .B(n9129), .ZN(n9131)
         );
  OAI21_X1 U10506 ( .B1(n9132), .B2(n9144), .A(n9131), .ZN(P1_U3233) );
  AND2_X1 U10507 ( .A1(n9135), .A2(n9134), .ZN(n9136) );
  NAND2_X1 U10508 ( .A1(n9133), .A2(n9136), .ZN(n9137) );
  XOR2_X1 U10509 ( .A(n9138), .B(n9137), .Z(n9145) );
  NAND2_X1 U10510 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9985) );
  OAI21_X1 U10511 ( .B1(n9162), .B2(n9776), .A(n9985), .ZN(n9141) );
  OAI22_X1 U10512 ( .A1(n9139), .A2(n9721), .B1(n9164), .B2(n9682), .ZN(n9140)
         );
  AOI211_X1 U10513 ( .C1(n9685), .C2(n9142), .A(n9141), .B(n9140), .ZN(n9143)
         );
  OAI21_X1 U10514 ( .B1(n9145), .B2(n9144), .A(n9143), .ZN(P1_U3236) );
  AND2_X1 U10515 ( .A1(n9147), .A2(n9146), .ZN(n9150) );
  OAI211_X1 U10516 ( .C1(n9150), .C2(n9149), .A(n9160), .B(n9148), .ZN(n9155)
         );
  OAI22_X1 U10517 ( .A1(n9549), .A2(n9164), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9151), .ZN(n9153) );
  NOR2_X1 U10518 ( .A1(n9546), .A2(n9162), .ZN(n9152) );
  AOI211_X1 U10519 ( .C1(n9167), .C2(n9578), .A(n9153), .B(n9152), .ZN(n9154)
         );
  OAI211_X1 U10520 ( .C1(n9836), .C2(n9170), .A(n9155), .B(n9154), .ZN(
        P1_U3238) );
  NAND2_X1 U10521 ( .A1(n9157), .A2(n9156), .ZN(n9159) );
  XNOR2_X1 U10522 ( .A(n9159), .B(n9158), .ZN(n9161) );
  NAND2_X1 U10523 ( .A1(n9161), .A2(n9160), .ZN(n9169) );
  OAI22_X1 U10524 ( .A1(n9164), .A2(n9163), .B1(n9162), .B2(n9699), .ZN(n9165)
         );
  AOI211_X1 U10525 ( .C1(n9167), .C2(n9817), .A(n9166), .B(n9165), .ZN(n9168)
         );
  OAI211_X1 U10526 ( .C1(n9171), .C2(n9170), .A(n9169), .B(n9168), .ZN(
        P1_U3239) );
  INV_X1 U10527 ( .A(n9176), .ZN(n9303) );
  AND2_X1 U10528 ( .A1(n9174), .A2(n9379), .ZN(n9376) );
  AOI21_X1 U10529 ( .B1(n9180), .B2(n9376), .A(n9175), .ZN(n9182) );
  AND2_X1 U10530 ( .A1(n9177), .A2(n9176), .ZN(n9179) );
  AOI21_X1 U10531 ( .B1(n9180), .B2(n9179), .A(n9178), .ZN(n9181) );
  MUX2_X1 U10532 ( .A(n9182), .B(n9181), .S(n9284), .Z(n9185) );
  INV_X1 U10533 ( .A(n9183), .ZN(n9184) );
  NAND2_X1 U10534 ( .A1(n9185), .A2(n9184), .ZN(n9191) );
  AND2_X1 U10535 ( .A1(n9300), .A2(n9418), .ZN(n9375) );
  NAND2_X1 U10536 ( .A1(n9192), .A2(n9187), .ZN(n9365) );
  INV_X1 U10537 ( .A(n9347), .ZN(n9186) );
  AND2_X1 U10538 ( .A1(n9188), .A2(n9187), .ZN(n9190) );
  NAND2_X1 U10539 ( .A1(n10011), .A2(n9418), .ZN(n9189) );
  NAND2_X1 U10540 ( .A1(n9307), .A2(n9192), .ZN(n9194) );
  AND2_X1 U10541 ( .A1(n9346), .A2(n9308), .ZN(n9193) );
  INV_X1 U10542 ( .A(n9195), .ZN(n9197) );
  NAND2_X1 U10543 ( .A1(n9203), .A2(n9346), .ZN(n9196) );
  MUX2_X1 U10544 ( .A(n9197), .B(n9196), .S(n4588), .Z(n9200) );
  INV_X1 U10545 ( .A(n9314), .ZN(n9198) );
  NAND2_X1 U10546 ( .A1(n9198), .A2(n9210), .ZN(n9199) );
  NOR2_X1 U10547 ( .A1(n9200), .A2(n9199), .ZN(n9201) );
  AND2_X1 U10548 ( .A1(n9210), .A2(n9202), .ZN(n9342) );
  INV_X1 U10549 ( .A(n9342), .ZN(n9204) );
  NAND2_X1 U10550 ( .A1(n9204), .A2(n9203), .ZN(n9205) );
  NAND3_X1 U10551 ( .A1(n9216), .A2(n9343), .A3(n9205), .ZN(n9209) );
  NAND2_X1 U10552 ( .A1(n9218), .A2(n9206), .ZN(n9214) );
  INV_X1 U10553 ( .A(n9214), .ZN(n9208) );
  INV_X1 U10554 ( .A(n9352), .ZN(n9207) );
  INV_X1 U10555 ( .A(n9210), .ZN(n9211) );
  NOR2_X1 U10556 ( .A1(n9212), .A2(n9211), .ZN(n9213) );
  OR2_X1 U10557 ( .A1(n9214), .A2(n9213), .ZN(n9351) );
  INV_X1 U10558 ( .A(n9351), .ZN(n9215) );
  NAND2_X1 U10559 ( .A1(n9216), .A2(n9215), .ZN(n9219) );
  NAND2_X1 U10560 ( .A1(n9218), .A2(n9217), .ZN(n9350) );
  NAND3_X1 U10561 ( .A1(n9219), .A2(n9352), .A3(n9350), .ZN(n9220) );
  MUX2_X1 U10562 ( .A(n9355), .B(n9353), .S(n4588), .Z(n9221) );
  INV_X1 U10563 ( .A(n9676), .ZN(n9222) );
  INV_X1 U10564 ( .A(n9697), .ZN(n9224) );
  MUX2_X1 U10565 ( .A(n9354), .B(n9369), .S(n9284), .Z(n9223) );
  NAND2_X1 U10566 ( .A1(n9233), .A2(n5273), .ZN(n9371) );
  INV_X1 U10567 ( .A(n9371), .ZN(n9226) );
  MUX2_X1 U10568 ( .A(n9335), .B(n9226), .S(n4588), .Z(n9227) );
  NAND2_X1 U10569 ( .A1(n9228), .A2(n9227), .ZN(n9235) );
  NAND3_X1 U10570 ( .A1(n9235), .A2(n9229), .A3(n9333), .ZN(n9231) );
  NOR2_X1 U10571 ( .A1(n9298), .A2(n9284), .ZN(n9230) );
  INV_X1 U10572 ( .A(n9234), .ZN(n9340) );
  NAND2_X1 U10573 ( .A1(n9333), .A2(n9284), .ZN(n9232) );
  NAND2_X1 U10574 ( .A1(n9234), .A2(n9233), .ZN(n9334) );
  INV_X1 U10575 ( .A(n9334), .ZN(n9236) );
  NAND3_X1 U10576 ( .A1(n9237), .A2(n9236), .A3(n9235), .ZN(n9241) );
  INV_X1 U10577 ( .A(n9299), .ZN(n9632) );
  NAND3_X1 U10578 ( .A1(n9297), .A2(n9244), .A3(n9632), .ZN(n9239) );
  NAND2_X1 U10579 ( .A1(n9244), .A2(n9298), .ZN(n9238) );
  AND2_X1 U10580 ( .A1(n9243), .A2(n9238), .ZN(n9339) );
  INV_X1 U10581 ( .A(n9339), .ZN(n9341) );
  MUX2_X1 U10582 ( .A(n9239), .B(n9341), .S(n9284), .Z(n9240) );
  INV_X1 U10583 ( .A(n9297), .ZN(n9242) );
  NOR2_X1 U10584 ( .A1(n9243), .A2(n9242), .ZN(n9247) );
  OR2_X1 U10585 ( .A1(n9341), .A2(n9244), .ZN(n9245) );
  AND2_X1 U10586 ( .A1(n9245), .A2(n9297), .ZN(n9362) );
  INV_X1 U10587 ( .A(n9362), .ZN(n9246) );
  NAND2_X1 U10588 ( .A1(n9583), .A2(n9598), .ZN(n9323) );
  INV_X1 U10589 ( .A(n9249), .ZN(n9250) );
  NAND2_X1 U10590 ( .A1(n9361), .A2(n9250), .ZN(n9251) );
  AND2_X1 U10591 ( .A1(n9251), .A2(n9253), .ZN(n9252) );
  AND2_X1 U10592 ( .A1(n9252), .A2(n9262), .ZN(n9427) );
  INV_X1 U10593 ( .A(n9427), .ZN(n9257) );
  NAND2_X1 U10594 ( .A1(n9361), .A2(n9336), .ZN(n9254) );
  NAND2_X1 U10595 ( .A1(n9254), .A2(n9253), .ZN(n9255) );
  NAND2_X1 U10596 ( .A1(n9541), .A2(n9255), .ZN(n9256) );
  MUX2_X1 U10597 ( .A(n9257), .B(n9256), .S(n9284), .Z(n9258) );
  INV_X1 U10598 ( .A(n9258), .ZN(n9259) );
  NAND2_X1 U10599 ( .A1(n9260), .A2(n9259), .ZN(n9264) );
  NAND2_X1 U10600 ( .A1(n9261), .A2(n4588), .ZN(n9267) );
  INV_X1 U10601 ( .A(n9262), .ZN(n9263) );
  XNOR2_X1 U10602 ( .A(n9265), .B(n9560), .ZN(n9543) );
  NAND2_X1 U10603 ( .A1(n9385), .A2(n9284), .ZN(n9266) );
  NAND3_X1 U10604 ( .A1(n9275), .A2(n9390), .A3(n9391), .ZN(n9268) );
  NAND2_X1 U10605 ( .A1(n9268), .A2(n9272), .ZN(n9270) );
  INV_X1 U10606 ( .A(n9437), .ZN(n9269) );
  INV_X1 U10607 ( .A(n9390), .ZN(n9274) );
  NAND2_X1 U10608 ( .A1(n9272), .A2(n9271), .ZN(n9388) );
  INV_X1 U10609 ( .A(n9388), .ZN(n9273) );
  OAI21_X1 U10610 ( .B1(n9275), .B2(n9274), .A(n9273), .ZN(n9276) );
  NAND2_X1 U10611 ( .A1(n9276), .A2(n9391), .ZN(n9277) );
  INV_X1 U10612 ( .A(n9392), .ZN(n9278) );
  NAND2_X1 U10613 ( .A1(n9288), .A2(n9456), .ZN(n9279) );
  NAND2_X1 U10614 ( .A1(n9501), .A2(n9279), .ZN(n9396) );
  INV_X1 U10615 ( .A(n9456), .ZN(n9294) );
  NOR2_X1 U10616 ( .A1(n9501), .A2(n9294), .ZN(n9328) );
  INV_X1 U10617 ( .A(n9328), .ZN(n9280) );
  NAND2_X1 U10618 ( .A1(n9280), .A2(n9288), .ZN(n9281) );
  INV_X1 U10619 ( .A(n9287), .ZN(n9290) );
  NAND2_X1 U10620 ( .A1(n9281), .A2(n9290), .ZN(n9400) );
  NAND2_X1 U10621 ( .A1(n9282), .A2(n9400), .ZN(n9286) );
  INV_X1 U10622 ( .A(n9400), .ZN(n9283) );
  NAND2_X1 U10623 ( .A1(n9284), .A2(n9283), .ZN(n9285) );
  AND2_X1 U10624 ( .A1(n9287), .A2(n9288), .ZN(n9439) );
  INV_X1 U10625 ( .A(n9439), .ZN(n9404) );
  OAI21_X1 U10626 ( .B1(n4588), .B2(n9396), .A(n9404), .ZN(n9292) );
  INV_X1 U10627 ( .A(n9288), .ZN(n9289) );
  AND2_X1 U10628 ( .A1(n9290), .A2(n9289), .ZN(n9329) );
  INV_X1 U10629 ( .A(n9329), .ZN(n9291) );
  NAND2_X1 U10630 ( .A1(n9292), .A2(n9291), .ZN(n9293) );
  AND2_X1 U10631 ( .A1(n9501), .A2(n9294), .ZN(n9408) );
  INV_X1 U10632 ( .A(n9295), .ZN(n9325) );
  NAND2_X1 U10633 ( .A1(n9297), .A2(n9296), .ZN(n9609) );
  NOR2_X1 U10634 ( .A1(n9299), .A2(n9298), .ZN(n9646) );
  NAND4_X1 U10635 ( .A1(n9376), .A2(n9302), .A3(n9301), .A4(n9300), .ZN(n9306)
         );
  OR2_X1 U10636 ( .A1(n9377), .A2(n9303), .ZN(n9420) );
  NOR4_X1 U10637 ( .A1(n9306), .A2(n9420), .A3(n9305), .A4(n9304), .ZN(n9312)
         );
  AND2_X1 U10638 ( .A1(n9308), .A2(n9307), .ZN(n10013) );
  INV_X1 U10639 ( .A(n9309), .ZN(n9310) );
  NAND4_X1 U10640 ( .A1(n9312), .A2(n10013), .A3(n9311), .A4(n9310), .ZN(n9316) );
  NOR4_X1 U10641 ( .A1(n9316), .A2(n9315), .A3(n9314), .A4(n9313), .ZN(n9317)
         );
  NAND4_X1 U10642 ( .A1(n4578), .A2(n9319), .A3(n9318), .A4(n9317), .ZN(n9320)
         );
  NOR4_X1 U10643 ( .A1(n9680), .A2(n9708), .A3(n9697), .A4(n9320), .ZN(n9321)
         );
  NAND4_X1 U10644 ( .A1(n9634), .A2(n9646), .A3(n9661), .A4(n9321), .ZN(n9322)
         );
  NOR4_X1 U10645 ( .A1(n9558), .A2(n9323), .A3(n9609), .A4(n9322), .ZN(n9324)
         );
  NAND4_X1 U10646 ( .A1(n9325), .A2(n9431), .A3(n9324), .A4(n9543), .ZN(n9326)
         );
  NOR4_X1 U10647 ( .A1(n9439), .A2(n9408), .A3(n9327), .A4(n9326), .ZN(n9330)
         );
  NOR2_X1 U10648 ( .A1(n9329), .A2(n9328), .ZN(n9441) );
  AOI21_X1 U10649 ( .B1(n9330), .B2(n9441), .A(n9411), .ZN(n9402) );
  INV_X1 U10650 ( .A(n9402), .ZN(n9331) );
  OAI211_X1 U10651 ( .C1(n9335), .C2(n9334), .A(n9632), .B(n9333), .ZN(n9338)
         );
  INV_X1 U10652 ( .A(n9336), .ZN(n9337) );
  AOI21_X1 U10653 ( .B1(n9339), .B2(n9338), .A(n9337), .ZN(n9363) );
  OR2_X1 U10654 ( .A1(n9341), .A2(n9340), .ZN(n9372) );
  INV_X1 U10655 ( .A(n9346), .ZN(n9345) );
  OAI211_X1 U10656 ( .C1(n9345), .C2(n9344), .A(n9343), .B(n9342), .ZN(n9366)
         );
  AND2_X1 U10657 ( .A1(n9347), .A2(n9346), .ZN(n9348) );
  NOR2_X1 U10658 ( .A1(n9366), .A2(n9348), .ZN(n9349) );
  AOI21_X1 U10659 ( .B1(n9351), .B2(n9350), .A(n9349), .ZN(n9356) );
  NAND2_X1 U10660 ( .A1(n9353), .A2(n9352), .ZN(n9364) );
  OAI211_X1 U10661 ( .C1(n9356), .C2(n9364), .A(n9355), .B(n9354), .ZN(n9357)
         );
  NAND2_X1 U10662 ( .A1(n9357), .A2(n9369), .ZN(n9358) );
  OR2_X1 U10663 ( .A1(n9371), .A2(n9358), .ZN(n9359) );
  OR2_X1 U10664 ( .A1(n9372), .A2(n9359), .ZN(n9360) );
  NAND4_X1 U10665 ( .A1(n9363), .A2(n9362), .A3(n9361), .A4(n9360), .ZN(n9429)
         );
  INV_X1 U10666 ( .A(n9364), .ZN(n9368) );
  NOR2_X1 U10667 ( .A1(n9366), .A2(n9365), .ZN(n9367) );
  NAND3_X1 U10668 ( .A1(n9369), .A2(n9368), .A3(n9367), .ZN(n9370) );
  OR3_X1 U10669 ( .A1(n9372), .A2(n9371), .A3(n9370), .ZN(n9426) );
  INV_X1 U10670 ( .A(n9373), .ZN(n9374) );
  NOR2_X1 U10671 ( .A1(n9420), .A2(n9374), .ZN(n9424) );
  OAI21_X1 U10672 ( .B1(n9377), .B2(n9376), .A(n9375), .ZN(n9382) );
  NAND2_X1 U10673 ( .A1(n9469), .A2(n10057), .ZN(n9378) );
  AND3_X1 U10674 ( .A1(n9418), .A2(n9379), .A3(n9378), .ZN(n9380) );
  AND2_X1 U10675 ( .A1(n9419), .A2(n9380), .ZN(n9417) );
  NAND2_X1 U10676 ( .A1(n7309), .A2(n9417), .ZN(n9381) );
  OAI21_X1 U10677 ( .B1(n9424), .B2(n9382), .A(n9381), .ZN(n9383) );
  NOR2_X1 U10678 ( .A1(n9426), .A2(n9383), .ZN(n9384) );
  OAI21_X1 U10679 ( .B1(n9429), .B2(n9384), .A(n9427), .ZN(n9389) );
  INV_X1 U10680 ( .A(n9385), .ZN(n9386) );
  AND2_X1 U10681 ( .A1(n9390), .A2(n9386), .ZN(n9387) );
  OR2_X1 U10682 ( .A1(n9388), .A2(n9387), .ZN(n9434) );
  AOI21_X1 U10683 ( .B1(n9390), .B2(n9389), .A(n9434), .ZN(n9397) );
  AND2_X1 U10684 ( .A1(n9392), .A2(n9391), .ZN(n9395) );
  OR2_X1 U10685 ( .A1(n9434), .A2(n9393), .ZN(n9394) );
  NAND2_X1 U10686 ( .A1(n9395), .A2(n9394), .ZN(n9432) );
  OAI211_X1 U10687 ( .C1(n9397), .C2(n9432), .A(n9396), .B(n9437), .ZN(n9399)
         );
  AOI211_X1 U10688 ( .C1(n9400), .C2(n9399), .A(n9398), .B(n9439), .ZN(n9401)
         );
  NOR2_X1 U10689 ( .A1(n9402), .A2(n9401), .ZN(n9403) );
  AND4_X1 U10690 ( .A1(n9406), .A2(n9411), .A3(n9405), .A4(n9404), .ZN(n9407)
         );
  INV_X1 U10691 ( .A(n9408), .ZN(n9438) );
  INV_X1 U10692 ( .A(n9409), .ZN(n9412) );
  NAND2_X1 U10693 ( .A1(n5597), .A2(n10053), .ZN(n9410) );
  NAND3_X1 U10694 ( .A1(n9412), .A2(n9411), .A3(n9410), .ZN(n9413) );
  NAND2_X1 U10695 ( .A1(n9414), .A2(n9413), .ZN(n9416) );
  OAI21_X1 U10696 ( .B1(n7003), .B2(n9416), .A(n9415), .ZN(n9423) );
  INV_X1 U10697 ( .A(n9417), .ZN(n9422) );
  NAND3_X1 U10698 ( .A1(n9420), .A2(n9419), .A3(n9418), .ZN(n9421) );
  AOI22_X1 U10699 ( .A1(n9424), .A2(n9423), .B1(n9422), .B2(n9421), .ZN(n9425)
         );
  NOR2_X1 U10700 ( .A1(n9426), .A2(n9425), .ZN(n9428) );
  OAI21_X1 U10701 ( .B1(n9429), .B2(n9428), .A(n9427), .ZN(n9430) );
  AND2_X1 U10702 ( .A1(n9431), .A2(n9430), .ZN(n9435) );
  INV_X1 U10703 ( .A(n9432), .ZN(n9433) );
  OAI21_X1 U10704 ( .B1(n9435), .B2(n9434), .A(n9433), .ZN(n9436) );
  NAND3_X1 U10705 ( .A1(n9438), .A2(n9437), .A3(n9436), .ZN(n9440) );
  AOI21_X1 U10706 ( .B1(n9441), .B2(n9440), .A(n9439), .ZN(n9442) );
  XNOR2_X1 U10707 ( .A(n9442), .B(n4390), .ZN(n9444) );
  NAND4_X1 U10708 ( .A1(n9450), .A2(n10051), .A3(n9449), .A4(n9448), .ZN(n9451) );
  OAI211_X1 U10709 ( .C1(n9452), .C2(n9454), .A(n9451), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9453) );
  OAI21_X1 U10710 ( .B1(n9455), .B2(n9454), .A(n9453), .ZN(P1_U3240) );
  MUX2_X1 U10711 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9456), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10712 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9457), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10713 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9458), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10714 ( .A(n9560), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9471), .Z(
        P1_U3581) );
  MUX2_X1 U10715 ( .A(n9578), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9471), .Z(
        P1_U3580) );
  MUX2_X1 U10716 ( .A(n9600), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9471), .Z(
        P1_U3579) );
  MUX2_X1 U10717 ( .A(n9614), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9471), .Z(
        P1_U3578) );
  MUX2_X1 U10718 ( .A(n9636), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9471), .Z(
        P1_U3577) );
  MUX2_X1 U10719 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9613), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10720 ( .A(n9787), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9471), .Z(
        P1_U3575) );
  MUX2_X1 U10721 ( .A(n9651), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9471), .Z(
        P1_U3574) );
  MUX2_X1 U10722 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9786), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10723 ( .A(n9806), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9471), .Z(
        P1_U3572) );
  MUX2_X1 U10724 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9459), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10725 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9807), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10726 ( .A(n9817), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9471), .Z(
        P1_U3569) );
  MUX2_X1 U10727 ( .A(n9460), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9471), .Z(
        P1_U3568) );
  MUX2_X1 U10728 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9820), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10729 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9461), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10730 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9462), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10731 ( .A(n9463), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9471), .Z(
        P1_U3564) );
  MUX2_X1 U10732 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9464), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10733 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9465), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10734 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9466), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10735 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9467), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10736 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9468), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10737 ( .A(n9469), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9471), .Z(
        P1_U3558) );
  MUX2_X1 U10738 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9470), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10739 ( .A(n5597), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9471), .Z(
        P1_U3556) );
  AOI211_X1 U10740 ( .C1(n4455), .C2(n9473), .A(n9472), .B(n9986), .ZN(n9483)
         );
  AOI211_X1 U10741 ( .C1(n9476), .C2(n9475), .A(n9474), .B(n9492), .ZN(n9482)
         );
  NAND2_X1 U10742 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n9479) );
  NAND2_X1 U10743 ( .A1(n9992), .A2(n9477), .ZN(n9478) );
  OAI211_X1 U10744 ( .C1(n9984), .C2(n9480), .A(n9479), .B(n9478), .ZN(n9481)
         );
  OR3_X1 U10745 ( .A1(n9483), .A2(n9482), .A3(n9481), .ZN(P1_U3257) );
  AOI211_X1 U10746 ( .C1(n9486), .C2(n9485), .A(n9484), .B(n9986), .ZN(n9498)
         );
  INV_X1 U10747 ( .A(n9487), .ZN(n9490) );
  NAND2_X1 U10748 ( .A1(n9997), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9489) );
  NAND2_X1 U10749 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n9488) );
  OAI211_X1 U10750 ( .C1(n9491), .C2(n9490), .A(n9489), .B(n9488), .ZN(n9497)
         );
  AOI211_X1 U10751 ( .C1(n9495), .C2(n9494), .A(n9493), .B(n9492), .ZN(n9496)
         );
  OR3_X1 U10752 ( .A1(n9498), .A2(n9497), .A3(n9496), .ZN(P1_U3258) );
  INV_X1 U10753 ( .A(n9499), .ZN(n9500) );
  XNOR2_X1 U10754 ( .A(n9501), .B(n9500), .ZN(n9502) );
  NAND2_X1 U10755 ( .A1(n9733), .A2(n10006), .ZN(n9505) );
  AOI21_X1 U10756 ( .B1(n10024), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9503), .ZN(
        n9504) );
  OAI211_X1 U10757 ( .C1(n6431), .C2(n9623), .A(n9505), .B(n9504), .ZN(
        P1_U3262) );
  INV_X1 U10758 ( .A(n9506), .ZN(n9514) );
  NAND2_X1 U10759 ( .A1(n9507), .A2(n10006), .ZN(n9510) );
  AOI22_X1 U10760 ( .A1(n9508), .A2(n10035), .B1(P1_REG2_REG_29__SCAN_IN), 
        .B2(n10024), .ZN(n9509) );
  OAI211_X1 U10761 ( .C1(n4625), .C2(n9623), .A(n9510), .B(n9509), .ZN(n9511)
         );
  AOI21_X1 U10762 ( .B1(n9512), .B2(n9629), .A(n9511), .ZN(n9513) );
  OAI21_X1 U10763 ( .B1(n9514), .B2(n9706), .A(n9513), .ZN(P1_U3355) );
  INV_X1 U10764 ( .A(n9515), .ZN(n9521) );
  NOR2_X1 U10765 ( .A1(n9516), .A2(n9724), .ZN(n9520) );
  AOI22_X1 U10766 ( .A1(n9517), .A2(n10035), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10024), .ZN(n9518) );
  OAI21_X1 U10767 ( .B1(n5486), .B2(n9623), .A(n9518), .ZN(n9519) );
  AOI211_X1 U10768 ( .C1(n9521), .C2(n9629), .A(n9520), .B(n9519), .ZN(n9522)
         );
  OAI21_X1 U10769 ( .B1(n9523), .B2(n9706), .A(n9522), .ZN(P1_U3263) );
  XNOR2_X1 U10770 ( .A(n9524), .B(n9530), .ZN(n9740) );
  AOI211_X1 U10771 ( .C1(n9737), .C2(n9525), .A(n9695), .B(n5487), .ZN(n9736)
         );
  AOI22_X1 U10772 ( .A1(n9527), .A2(n10035), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10024), .ZN(n9528) );
  OAI21_X1 U10773 ( .B1(n9529), .B2(n9623), .A(n9528), .ZN(n9538) );
  AOI21_X1 U10774 ( .B1(n9531), .B2(n9530), .A(n10020), .ZN(n9536) );
  OAI22_X1 U10775 ( .A1(n9534), .A2(n10062), .B1(n9533), .B2(n10015), .ZN(
        n9535) );
  AOI21_X1 U10776 ( .B1(n9536), .B2(n9532), .A(n9535), .ZN(n9739) );
  NOR2_X1 U10777 ( .A1(n9739), .A2(n10024), .ZN(n9537) );
  OAI21_X1 U10778 ( .B1(n9740), .B2(n9706), .A(n9539), .ZN(P1_U3264) );
  XNOR2_X1 U10779 ( .A(n9540), .B(n9543), .ZN(n9743) );
  NAND2_X1 U10780 ( .A1(n9542), .A2(n9541), .ZN(n9544) );
  XNOR2_X1 U10781 ( .A(n9544), .B(n4584), .ZN(n9548) );
  OAI22_X1 U10782 ( .A1(n9546), .A2(n10062), .B1(n9545), .B2(n10015), .ZN(
        n9547) );
  AOI21_X1 U10783 ( .B1(n9548), .B2(n9637), .A(n9547), .ZN(n9742) );
  INV_X1 U10784 ( .A(n9742), .ZN(n9554) );
  OAI211_X1 U10785 ( .C1(n4449), .C2(n9836), .A(n10003), .B(n9525), .ZN(n9741)
         );
  NOR2_X1 U10786 ( .A1(n9741), .A2(n9724), .ZN(n9553) );
  INV_X1 U10787 ( .A(n9549), .ZN(n9550) );
  AOI22_X1 U10788 ( .A1(n9550), .A2(n10035), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10024), .ZN(n9551) );
  OAI21_X1 U10789 ( .B1(n9836), .B2(n9623), .A(n9551), .ZN(n9552) );
  AOI211_X1 U10790 ( .C1(n9554), .C2(n9629), .A(n9553), .B(n9552), .ZN(n9555)
         );
  OAI21_X1 U10791 ( .B1(n9743), .B2(n9706), .A(n9555), .ZN(P1_U3265) );
  OAI21_X1 U10792 ( .B1(n4440), .B2(n9558), .A(n9556), .ZN(n9749) );
  INV_X1 U10793 ( .A(n9749), .ZN(n9570) );
  XNOR2_X1 U10794 ( .A(n9557), .B(n9558), .ZN(n9559) );
  NAND2_X1 U10795 ( .A1(n9559), .A2(n9637), .ZN(n9562) );
  AOI22_X1 U10796 ( .A1(n9560), .A2(n9818), .B1(n9819), .B2(n9600), .ZN(n9561)
         );
  NAND2_X1 U10797 ( .A1(n9562), .A2(n9561), .ZN(n9747) );
  AOI211_X1 U10798 ( .C1(n9563), .C2(n9572), .A(n9695), .B(n4449), .ZN(n9748)
         );
  NAND2_X1 U10799 ( .A1(n9748), .A2(n10006), .ZN(n9567) );
  INV_X1 U10800 ( .A(n9564), .ZN(n9565) );
  AOI22_X1 U10801 ( .A1(n9565), .A2(n10035), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10024), .ZN(n9566) );
  OAI211_X1 U10802 ( .C1(n9840), .C2(n9623), .A(n9567), .B(n9566), .ZN(n9568)
         );
  AOI21_X1 U10803 ( .B1(n9747), .B2(n9629), .A(n9568), .ZN(n9569) );
  OAI21_X1 U10804 ( .B1(n9570), .B2(n9706), .A(n9569), .ZN(P1_U3266) );
  INV_X1 U10805 ( .A(n9572), .ZN(n9573) );
  AOI211_X1 U10806 ( .C1(n9756), .C2(n9571), .A(n9695), .B(n9573), .ZN(n9755)
         );
  INV_X1 U10807 ( .A(n9574), .ZN(n9575) );
  NOR2_X1 U10808 ( .A1(n9575), .A2(n10008), .ZN(n9582) );
  OAI211_X1 U10809 ( .C1(n9577), .C2(n9583), .A(n9576), .B(n9637), .ZN(n9580)
         );
  NAND2_X1 U10810 ( .A1(n9578), .A2(n9818), .ZN(n9579) );
  OAI211_X1 U10811 ( .C1(n9581), .C2(n10015), .A(n9580), .B(n9579), .ZN(n9754)
         );
  AOI211_X1 U10812 ( .C1(n9755), .C2(n4390), .A(n9582), .B(n9754), .ZN(n9587)
         );
  NAND2_X1 U10813 ( .A1(n9584), .A2(n9583), .ZN(n9752) );
  NAND3_X1 U10814 ( .A1(n9753), .A2(n9752), .A3(n9714), .ZN(n9586) );
  AOI22_X1 U10815 ( .A1(n9756), .A2(n10028), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10024), .ZN(n9585) );
  OAI211_X1 U10816 ( .C1(n10024), .C2(n9587), .A(n9586), .B(n9585), .ZN(
        P1_U3267) );
  XOR2_X1 U10817 ( .A(n9588), .B(n9598), .Z(n9763) );
  INV_X1 U10818 ( .A(n9589), .ZN(n9591) );
  INV_X1 U10819 ( .A(n9571), .ZN(n9590) );
  AOI211_X1 U10820 ( .C1(n9761), .C2(n9591), .A(n9695), .B(n9590), .ZN(n9760)
         );
  NOR2_X1 U10821 ( .A1(n9592), .A2(n9623), .ZN(n9596) );
  OAI22_X1 U10822 ( .A1(n9594), .A2(n10008), .B1(n9593), .B2(n9629), .ZN(n9595) );
  AOI211_X1 U10823 ( .C1(n9760), .C2(n10006), .A(n9596), .B(n9595), .ZN(n9605)
         );
  OAI211_X1 U10824 ( .C1(n9599), .C2(n9598), .A(n9597), .B(n9637), .ZN(n9602)
         );
  NAND2_X1 U10825 ( .A1(n9600), .A2(n9818), .ZN(n9601) );
  OAI211_X1 U10826 ( .C1(n9603), .C2(n10015), .A(n9602), .B(n9601), .ZN(n9759)
         );
  NAND2_X1 U10827 ( .A1(n9759), .A2(n9629), .ZN(n9604) );
  OAI211_X1 U10828 ( .C1(n9763), .C2(n9706), .A(n9605), .B(n9604), .ZN(
        P1_U3268) );
  XOR2_X1 U10829 ( .A(n9606), .B(n9609), .Z(n9766) );
  INV_X1 U10830 ( .A(n9766), .ZN(n9626) );
  NAND2_X1 U10831 ( .A1(n9607), .A2(n9608), .ZN(n9611) );
  INV_X1 U10832 ( .A(n9609), .ZN(n9610) );
  XNOR2_X1 U10833 ( .A(n9611), .B(n9610), .ZN(n9612) );
  NAND2_X1 U10834 ( .A1(n9612), .A2(n9637), .ZN(n9616) );
  AOI22_X1 U10835 ( .A1(n9818), .A2(n9614), .B1(n9613), .B2(n9819), .ZN(n9615)
         );
  NAND2_X1 U10836 ( .A1(n9616), .A2(n9615), .ZN(n9764) );
  INV_X1 U10837 ( .A(n9639), .ZN(n9617) );
  AOI211_X1 U10838 ( .C1(n9618), .C2(n9617), .A(n9695), .B(n9589), .ZN(n9765)
         );
  NAND2_X1 U10839 ( .A1(n9765), .A2(n10006), .ZN(n9622) );
  INV_X1 U10840 ( .A(n9619), .ZN(n9620) );
  AOI22_X1 U10841 ( .A1(n9620), .A2(n10035), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10024), .ZN(n9621) );
  OAI211_X1 U10842 ( .C1(n9846), .C2(n9623), .A(n9622), .B(n9621), .ZN(n9624)
         );
  AOI21_X1 U10843 ( .B1(n9764), .B2(n9629), .A(n9624), .ZN(n9625) );
  OAI21_X1 U10844 ( .B1(n9626), .B2(n9706), .A(n9625), .ZN(P1_U3269) );
  OAI21_X1 U10845 ( .B1(n4401), .B2(n9628), .A(n9627), .ZN(n9775) );
  INV_X1 U10846 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9630) );
  OAI22_X1 U10847 ( .A1(n9769), .A2(n9631), .B1(n9630), .B2(n9629), .ZN(n9643)
         );
  AND2_X1 U10848 ( .A1(n9633), .A2(n9632), .ZN(n9635) );
  OAI21_X1 U10849 ( .B1(n9635), .B2(n9634), .A(n9607), .ZN(n9638) );
  AOI22_X1 U10850 ( .A1(n9638), .A2(n9637), .B1(n9818), .B2(n9636), .ZN(n9774)
         );
  AOI211_X1 U10851 ( .C1(n9772), .C2(n9653), .A(n9695), .B(n9639), .ZN(n9770)
         );
  AOI22_X1 U10852 ( .A1(n9770), .A2(n4390), .B1(n10035), .B2(n9640), .ZN(n9641) );
  AOI21_X1 U10853 ( .B1(n9774), .B2(n9641), .A(n10024), .ZN(n9642) );
  AOI211_X1 U10854 ( .C1(n10028), .C2(n9772), .A(n9643), .B(n9642), .ZN(n9644)
         );
  OAI21_X1 U10855 ( .B1(n9775), .B2(n9706), .A(n9644), .ZN(P1_U3270) );
  XOR2_X1 U10856 ( .A(n9645), .B(n9646), .Z(n9781) );
  XNOR2_X1 U10857 ( .A(n9647), .B(n9646), .ZN(n9783) );
  NAND2_X1 U10858 ( .A1(n9783), .A2(n9714), .ZN(n9659) );
  OAI22_X1 U10859 ( .A1(n9629), .A2(n9649), .B1(n9648), .B2(n10008), .ZN(n9650) );
  AOI21_X1 U10860 ( .B1(n9718), .B2(n9651), .A(n9650), .ZN(n9652) );
  OAI21_X1 U10861 ( .B1(n9777), .B2(n9720), .A(n9652), .ZN(n9656) );
  NAND2_X1 U10862 ( .A1(n9674), .A2(n9855), .ZN(n9667) );
  AOI21_X1 U10863 ( .B1(n9667), .B2(n9657), .A(n9695), .ZN(n9654) );
  NAND2_X1 U10864 ( .A1(n9654), .A2(n9653), .ZN(n9779) );
  NOR2_X1 U10865 ( .A1(n9779), .A2(n9724), .ZN(n9655) );
  AOI211_X1 U10866 ( .C1(n10028), .C2(n9657), .A(n9656), .B(n9655), .ZN(n9658)
         );
  OAI211_X1 U10867 ( .C1(n9781), .C2(n9730), .A(n9659), .B(n9658), .ZN(
        P1_U3271) );
  XOR2_X1 U10868 ( .A(n9660), .B(n9661), .Z(n9790) );
  XNOR2_X1 U10869 ( .A(n9662), .B(n9661), .ZN(n9792) );
  NAND2_X1 U10870 ( .A1(n9792), .A2(n9714), .ZN(n9672) );
  INV_X1 U10871 ( .A(n9663), .ZN(n9664) );
  AOI22_X1 U10872 ( .A1(n10024), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9664), 
        .B2(n10035), .ZN(n9666) );
  NAND2_X1 U10873 ( .A1(n9718), .A2(n9786), .ZN(n9665) );
  OAI211_X1 U10874 ( .C1(n9769), .C2(n9720), .A(n9666), .B(n9665), .ZN(n9669)
         );
  OAI211_X1 U10875 ( .C1(n9674), .C2(n9855), .A(n10003), .B(n9667), .ZN(n9788)
         );
  NOR2_X1 U10876 ( .A1(n9788), .A2(n9724), .ZN(n9668) );
  AOI211_X1 U10877 ( .C1(n10028), .C2(n9670), .A(n9669), .B(n9668), .ZN(n9671)
         );
  OAI211_X1 U10878 ( .C1(n9730), .C2(n9790), .A(n9672), .B(n9671), .ZN(
        P1_U3272) );
  INV_X1 U10879 ( .A(n9673), .ZN(n9675) );
  AOI211_X1 U10880 ( .C1(n9685), .C2(n9675), .A(n9695), .B(n9674), .ZN(n9796)
         );
  NAND2_X1 U10881 ( .A1(n9677), .A2(n9676), .ZN(n9678) );
  XOR2_X1 U10882 ( .A(n9680), .B(n9678), .Z(n9679) );
  OAI222_X1 U10883 ( .A1(n10062), .A2(n9776), .B1(n10015), .B2(n9721), .C1(
        n10020), .C2(n9679), .ZN(n9795) );
  AOI21_X1 U10884 ( .B1(n9796), .B2(n4390), .A(n9795), .ZN(n9688) );
  XOR2_X1 U10885 ( .A(n9681), .B(n9680), .Z(n9797) );
  NAND2_X1 U10886 ( .A1(n9797), .A2(n9714), .ZN(n9687) );
  OAI22_X1 U10887 ( .A1(n9629), .A2(n9683), .B1(n9682), .B2(n10008), .ZN(n9684) );
  AOI21_X1 U10888 ( .B1(n9685), .B2(n10028), .A(n9684), .ZN(n9686) );
  OAI211_X1 U10889 ( .C1(n10024), .C2(n9688), .A(n9687), .B(n9686), .ZN(
        P1_U3273) );
  NAND2_X1 U10890 ( .A1(n7839), .A2(n9689), .ZN(n9691) );
  NAND2_X1 U10891 ( .A1(n9691), .A2(n9690), .ZN(n9692) );
  XNOR2_X1 U10892 ( .A(n9692), .B(n9697), .ZN(n9805) );
  INV_X1 U10893 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9694) );
  OAI22_X1 U10894 ( .A1(n9629), .A2(n9694), .B1(n9693), .B2(n10008), .ZN(n9704) );
  AOI211_X1 U10895 ( .C1(n9802), .C2(n4454), .A(n9695), .B(n9673), .ZN(n9801)
         );
  XNOR2_X1 U10896 ( .A(n9696), .B(n9697), .ZN(n9698) );
  OAI222_X1 U10897 ( .A1(n10062), .A2(n9700), .B1(n10015), .B2(n9699), .C1(
        n9698), .C2(n10020), .ZN(n9800) );
  AOI21_X1 U10898 ( .B1(n9801), .B2(n4390), .A(n9800), .ZN(n9702) );
  NOR2_X1 U10899 ( .A1(n9702), .A2(n10024), .ZN(n9703) );
  AOI211_X1 U10900 ( .C1(n10028), .C2(n9802), .A(n9704), .B(n9703), .ZN(n9705)
         );
  OAI21_X1 U10901 ( .B1(n9706), .B2(n9805), .A(n9705), .ZN(P1_U3274) );
  XNOR2_X1 U10902 ( .A(n9707), .B(n9708), .ZN(n9810) );
  NAND2_X1 U10903 ( .A1(n7839), .A2(n9709), .ZN(n9711) );
  NAND2_X1 U10904 ( .A1(n9711), .A2(n9710), .ZN(n9713) );
  XNOR2_X1 U10905 ( .A(n9713), .B(n9712), .ZN(n9812) );
  NAND2_X1 U10906 ( .A1(n9812), .A2(n9714), .ZN(n9729) );
  OAI22_X1 U10907 ( .A1(n9629), .A2(n9716), .B1(n9715), .B2(n10008), .ZN(n9717) );
  AOI21_X1 U10908 ( .B1(n9718), .B2(n9807), .A(n9717), .ZN(n9719) );
  OAI21_X1 U10909 ( .B1(n9721), .B2(n9720), .A(n9719), .ZN(n9726) );
  INV_X1 U10910 ( .A(n9722), .ZN(n9723) );
  INV_X1 U10911 ( .A(n9727), .ZN(n9865) );
  OAI211_X1 U10912 ( .C1(n9723), .C2(n9865), .A(n10003), .B(n4454), .ZN(n9808)
         );
  NOR2_X1 U10913 ( .A1(n9808), .A2(n9724), .ZN(n9725) );
  AOI211_X1 U10914 ( .C1(n10028), .C2(n9727), .A(n9726), .B(n9725), .ZN(n9728)
         );
  OAI211_X1 U10915 ( .C1(n9810), .C2(n9730), .A(n9729), .B(n9728), .ZN(
        P1_U3275) );
  INV_X1 U10916 ( .A(n9731), .ZN(n9732) );
  NOR2_X1 U10917 ( .A1(n9733), .A2(n9732), .ZN(n9829) );
  MUX2_X1 U10918 ( .A(n9734), .B(n9829), .S(n10083), .Z(n9735) );
  OAI21_X1 U10919 ( .B1(n6431), .B2(n9815), .A(n9735), .ZN(P1_U3553) );
  AOI21_X1 U10920 ( .B1(n9803), .B2(n9737), .A(n9736), .ZN(n9738) );
  OAI211_X1 U10921 ( .C1(n9740), .C2(n7672), .A(n9739), .B(n9738), .ZN(n9832)
         );
  MUX2_X1 U10922 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9832), .S(n10083), .Z(
        P1_U3550) );
  OAI211_X1 U10923 ( .C1(n9743), .C2(n7672), .A(n9742), .B(n9741), .ZN(n9744)
         );
  INV_X1 U10924 ( .A(n9744), .ZN(n9833) );
  MUX2_X1 U10925 ( .A(n9745), .B(n9833), .S(n10083), .Z(n9746) );
  OAI21_X1 U10926 ( .B1(n9836), .B2(n9815), .A(n9746), .ZN(P1_U3549) );
  AOI211_X1 U10927 ( .C1(n9749), .C2(n10066), .A(n9748), .B(n9747), .ZN(n9837)
         );
  MUX2_X1 U10928 ( .A(n9750), .B(n9837), .S(n10083), .Z(n9751) );
  OAI21_X1 U10929 ( .B1(n9840), .B2(n9815), .A(n9751), .ZN(P1_U3548) );
  NAND3_X1 U10930 ( .A1(n9753), .A2(n10066), .A3(n9752), .ZN(n9758) );
  AOI211_X1 U10931 ( .C1(n9803), .C2(n9756), .A(n9755), .B(n9754), .ZN(n9757)
         );
  NAND2_X1 U10932 ( .A1(n9758), .A2(n9757), .ZN(n9841) );
  MUX2_X1 U10933 ( .A(n9841), .B(P1_REG1_REG_24__SCAN_IN), .S(n10081), .Z(
        P1_U3547) );
  AOI211_X1 U10934 ( .C1(n9803), .C2(n9761), .A(n9760), .B(n9759), .ZN(n9762)
         );
  OAI21_X1 U10935 ( .B1(n9763), .B2(n7672), .A(n9762), .ZN(n9842) );
  MUX2_X1 U10936 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9842), .S(n10083), .Z(
        P1_U3546) );
  AOI211_X1 U10937 ( .C1(n9766), .C2(n10066), .A(n9765), .B(n9764), .ZN(n9843)
         );
  MUX2_X1 U10938 ( .A(n9767), .B(n9843), .S(n10083), .Z(n9768) );
  OAI21_X1 U10939 ( .B1(n9846), .B2(n9815), .A(n9768), .ZN(P1_U3545) );
  NOR2_X1 U10940 ( .A1(n9769), .A2(n10015), .ZN(n9771) );
  AOI211_X1 U10941 ( .C1(n9803), .C2(n9772), .A(n9771), .B(n9770), .ZN(n9773)
         );
  OAI211_X1 U10942 ( .C1(n9775), .C2(n7672), .A(n9774), .B(n9773), .ZN(n9847)
         );
  MUX2_X1 U10943 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9847), .S(n10083), .Z(
        P1_U3544) );
  OAI22_X1 U10944 ( .A1(n9777), .A2(n10062), .B1(n9776), .B2(n10015), .ZN(
        n9778) );
  INV_X1 U10945 ( .A(n9778), .ZN(n9780) );
  OAI211_X1 U10946 ( .C1(n9781), .C2(n10020), .A(n9780), .B(n9779), .ZN(n9782)
         );
  AOI21_X1 U10947 ( .B1(n9783), .B2(n10066), .A(n9782), .ZN(n9848) );
  MUX2_X1 U10948 ( .A(n9784), .B(n9848), .S(n10083), .Z(n9785) );
  OAI21_X1 U10949 ( .B1(n9851), .B2(n9815), .A(n9785), .ZN(P1_U3543) );
  AOI22_X1 U10950 ( .A1(n9818), .A2(n9787), .B1(n9786), .B2(n9819), .ZN(n9789)
         );
  OAI211_X1 U10951 ( .C1(n9790), .C2(n10020), .A(n9789), .B(n9788), .ZN(n9791)
         );
  AOI21_X1 U10952 ( .B1(n9792), .B2(n10066), .A(n9791), .ZN(n9852) );
  MUX2_X1 U10953 ( .A(n9793), .B(n9852), .S(n10083), .Z(n9794) );
  OAI21_X1 U10954 ( .B1(n9855), .B2(n9815), .A(n9794), .ZN(P1_U3542) );
  AOI211_X1 U10955 ( .C1(n9797), .C2(n10066), .A(n9796), .B(n9795), .ZN(n9856)
         );
  MUX2_X1 U10956 ( .A(n9798), .B(n9856), .S(n10083), .Z(n9799) );
  OAI21_X1 U10957 ( .B1(n9859), .B2(n9815), .A(n9799), .ZN(P1_U3541) );
  AOI211_X1 U10958 ( .C1(n9803), .C2(n9802), .A(n9801), .B(n9800), .ZN(n9804)
         );
  OAI21_X1 U10959 ( .B1(n9805), .B2(n7672), .A(n9804), .ZN(n9860) );
  MUX2_X1 U10960 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9860), .S(n10083), .Z(
        P1_U3540) );
  AOI22_X1 U10961 ( .A1(n9807), .A2(n9819), .B1(n9818), .B2(n9806), .ZN(n9809)
         );
  OAI211_X1 U10962 ( .C1(n9810), .C2(n10020), .A(n9809), .B(n9808), .ZN(n9811)
         );
  AOI21_X1 U10963 ( .B1(n9812), .B2(n10066), .A(n9811), .ZN(n9861) );
  MUX2_X1 U10964 ( .A(n9813), .B(n9861), .S(n10083), .Z(n9814) );
  OAI21_X1 U10965 ( .B1(n9865), .B2(n9815), .A(n9814), .ZN(P1_U3539) );
  INV_X1 U10966 ( .A(n9816), .ZN(n9823) );
  AOI22_X1 U10967 ( .A1(n9820), .A2(n9819), .B1(n9818), .B2(n9817), .ZN(n9821)
         );
  OAI211_X1 U10968 ( .C1(n9823), .C2(n10071), .A(n9822), .B(n9821), .ZN(n9824)
         );
  AOI211_X1 U10969 ( .C1(n9826), .C2(n10066), .A(n9825), .B(n9824), .ZN(n9827)
         );
  INV_X1 U10970 ( .A(n9827), .ZN(n9866) );
  MUX2_X1 U10971 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9866), .S(n10083), .Z(
        P1_U3536) );
  MUX2_X1 U10972 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9828), .S(n10083), .Z(
        P1_U3523) );
  INV_X1 U10973 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9830) );
  MUX2_X1 U10974 ( .A(n9830), .B(n9829), .S(n10076), .Z(n9831) );
  OAI21_X1 U10975 ( .B1(n6431), .B2(n9864), .A(n9831), .ZN(P1_U3521) );
  MUX2_X1 U10976 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9832), .S(n10076), .Z(
        P1_U3518) );
  INV_X1 U10977 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9834) );
  MUX2_X1 U10978 ( .A(n9834), .B(n9833), .S(n10076), .Z(n9835) );
  OAI21_X1 U10979 ( .B1(n9836), .B2(n9864), .A(n9835), .ZN(P1_U3517) );
  INV_X1 U10980 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9838) );
  MUX2_X1 U10981 ( .A(n9838), .B(n9837), .S(n10076), .Z(n9839) );
  OAI21_X1 U10982 ( .B1(n9840), .B2(n9864), .A(n9839), .ZN(P1_U3516) );
  MUX2_X1 U10983 ( .A(n9841), .B(P1_REG0_REG_24__SCAN_IN), .S(n10075), .Z(
        P1_U3515) );
  MUX2_X1 U10984 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9842), .S(n10076), .Z(
        P1_U3514) );
  INV_X1 U10985 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9844) );
  MUX2_X1 U10986 ( .A(n9844), .B(n9843), .S(n10076), .Z(n9845) );
  OAI21_X1 U10987 ( .B1(n9846), .B2(n9864), .A(n9845), .ZN(P1_U3513) );
  MUX2_X1 U10988 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9847), .S(n10076), .Z(
        P1_U3512) );
  MUX2_X1 U10989 ( .A(n9849), .B(n9848), .S(n10076), .Z(n9850) );
  OAI21_X1 U10990 ( .B1(n9851), .B2(n9864), .A(n9850), .ZN(P1_U3511) );
  MUX2_X1 U10991 ( .A(n9853), .B(n9852), .S(n10076), .Z(n9854) );
  OAI21_X1 U10992 ( .B1(n9855), .B2(n9864), .A(n9854), .ZN(P1_U3510) );
  INV_X1 U10993 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9857) );
  MUX2_X1 U10994 ( .A(n9857), .B(n9856), .S(n10076), .Z(n9858) );
  OAI21_X1 U10995 ( .B1(n9859), .B2(n9864), .A(n9858), .ZN(P1_U3508) );
  MUX2_X1 U10996 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9860), .S(n10076), .Z(
        P1_U3505) );
  INV_X1 U10997 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9862) );
  MUX2_X1 U10998 ( .A(n9862), .B(n9861), .S(n10076), .Z(n9863) );
  OAI21_X1 U10999 ( .B1(n9865), .B2(n9864), .A(n9863), .ZN(P1_U3502) );
  MUX2_X1 U11000 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9866), .S(n10076), .Z(
        P1_U3493) );
  MUX2_X1 U11001 ( .A(P1_D_REG_0__SCAN_IN), .B(n9867), .S(n10051), .Z(P1_U3440) );
  INV_X1 U11002 ( .A(n9868), .ZN(n9873) );
  NOR4_X1 U11003 ( .A1(n9869), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n5187), .ZN(n9870) );
  AOI21_X1 U11004 ( .B1(n9871), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9870), .ZN(
        n9872) );
  OAI21_X1 U11005 ( .B1(n9873), .B2(n9878), .A(n9872), .ZN(P1_U3322) );
  OAI222_X1 U11006 ( .A1(n9878), .A2(n9877), .B1(n9876), .B2(P1_U3084), .C1(
        n9875), .C2(n9874), .ZN(P1_U3323) );
  NOR2_X1 U11007 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9879) );
  AOI21_X1 U11008 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9879), .ZN(n10282) );
  NOR2_X1 U11009 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_16__SCAN_IN), 
        .ZN(n9880) );
  AOI21_X1 U11010 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9880), .ZN(n10285) );
  NOR2_X1 U11011 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9881) );
  AOI21_X1 U11012 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9881), .ZN(n10288) );
  NOR2_X1 U11013 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9882) );
  AOI21_X1 U11014 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9882), .ZN(n10291) );
  NOR2_X1 U11015 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9883) );
  AOI21_X1 U11016 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9883), .ZN(n10294) );
  NOR2_X1 U11017 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(P1_ADDR_REG_4__SCAN_IN), 
        .ZN(n9891) );
  INV_X1 U11018 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9931) );
  AOI22_X1 U11019 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n9931), .B1(
        P1_ADDR_REG_4__SCAN_IN), .B2(n9884), .ZN(n10325) );
  NAND2_X1 U11020 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9889) );
  XOR2_X1 U11021 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10323) );
  NAND2_X1 U11022 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9887) );
  XOR2_X1 U11023 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10321) );
  AOI21_X1 U11024 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10276) );
  NAND3_X1 U11025 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10278) );
  OAI21_X1 U11026 ( .B1(n10276), .B2(n9885), .A(n10278), .ZN(n10320) );
  NAND2_X1 U11027 ( .A1(n10321), .A2(n10320), .ZN(n9886) );
  NAND2_X1 U11028 ( .A1(n9887), .A2(n9886), .ZN(n10322) );
  NAND2_X1 U11029 ( .A1(n10323), .A2(n10322), .ZN(n9888) );
  NAND2_X1 U11030 ( .A1(n9889), .A2(n9888), .ZN(n10324) );
  NOR2_X1 U11031 ( .A1(n10325), .A2(n10324), .ZN(n9890) );
  NOR2_X1 U11032 ( .A1(n9891), .A2(n9890), .ZN(n9892) );
  NOR2_X1 U11033 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9892), .ZN(n10308) );
  AND2_X1 U11034 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9892), .ZN(n10307) );
  NOR2_X1 U11035 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10307), .ZN(n9893) );
  NOR2_X1 U11036 ( .A1(n10308), .A2(n9893), .ZN(n9894) );
  NAND2_X1 U11037 ( .A1(n9894), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9896) );
  XOR2_X1 U11038 ( .A(n9894), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10306) );
  NAND2_X1 U11039 ( .A1(n10306), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9895) );
  NAND2_X1 U11040 ( .A1(n9896), .A2(n9895), .ZN(n9897) );
  AND2_X1 U11041 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9897), .ZN(n9898) );
  XNOR2_X1 U11042 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9897), .ZN(n10311) );
  INV_X1 U11043 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n9900) );
  NOR2_X1 U11044 ( .A1(n9899), .A2(n9900), .ZN(n9901) );
  XNOR2_X1 U11045 ( .A(n9900), .B(n9899), .ZN(n10305) );
  INV_X1 U11046 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n9903) );
  NOR2_X1 U11047 ( .A1(n9902), .A2(n9903), .ZN(n9904) );
  INV_X1 U11048 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10319) );
  XNOR2_X1 U11049 ( .A(n9903), .B(n9902), .ZN(n10318) );
  NAND2_X1 U11050 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9905) );
  OAI21_X1 U11051 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9905), .ZN(n10302) );
  NAND2_X1 U11052 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9906) );
  OAI21_X1 U11053 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9906), .ZN(n10299) );
  AOI21_X1 U11054 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10298), .ZN(n10297) );
  NOR2_X1 U11055 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(P2_ADDR_REG_12__SCAN_IN), 
        .ZN(n9907) );
  AOI21_X1 U11056 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9907), .ZN(n10296) );
  NAND2_X1 U11057 ( .A1(n10297), .A2(n10296), .ZN(n10295) );
  OAI21_X1 U11058 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10295), .ZN(n10293) );
  NAND2_X1 U11059 ( .A1(n10294), .A2(n10293), .ZN(n10292) );
  OAI21_X1 U11060 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10292), .ZN(n10290) );
  NAND2_X1 U11061 ( .A1(n10291), .A2(n10290), .ZN(n10289) );
  OAI21_X1 U11062 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10289), .ZN(n10287) );
  NAND2_X1 U11063 ( .A1(n10288), .A2(n10287), .ZN(n10286) );
  OAI21_X1 U11064 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10286), .ZN(n10284) );
  NAND2_X1 U11065 ( .A1(n10285), .A2(n10284), .ZN(n10283) );
  OAI21_X1 U11066 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10283), .ZN(n10281) );
  NAND2_X1 U11067 ( .A1(n10282), .A2(n10281), .ZN(n10280) );
  OAI21_X1 U11068 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10280), .ZN(n10314) );
  NOR2_X1 U11069 ( .A1(n10315), .A2(n10314), .ZN(n9908) );
  NAND2_X1 U11070 ( .A1(n10315), .A2(n10314), .ZN(n10313) );
  OAI21_X1 U11071 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9908), .A(n10313), .ZN(
        n9910) );
  XOR2_X1 U11072 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n9909) );
  XNOR2_X1 U11073 ( .A(n9910), .B(n9909), .ZN(ADD_1071_U4) );
  OAI21_X1 U11074 ( .B1(n9912), .B2(n10071), .A(n9911), .ZN(n9914) );
  NOR2_X1 U11075 ( .A1(n9914), .A2(n9913), .ZN(n9917) );
  AOI22_X1 U11076 ( .A1(n10083), .A2(n9917), .B1(n9915), .B2(n10081), .ZN(
        P1_U3534) );
  AOI22_X1 U11077 ( .A1(n10076), .A2(n9917), .B1(n9916), .B2(n10075), .ZN(
        P1_U3487) );
  XNOR2_X1 U11078 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11079 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  OAI21_X1 U11080 ( .B1(n9920), .B2(n9919), .A(n9918), .ZN(n9925) );
  OAI21_X1 U11081 ( .B1(n9923), .B2(n9922), .A(n9921), .ZN(n9924) );
  AOI22_X1 U11082 ( .A1(n9998), .A2(n9925), .B1(n9966), .B2(n9924), .ZN(n9930)
         );
  AOI211_X1 U11083 ( .C1(n9992), .C2(n9928), .A(n9927), .B(n9926), .ZN(n9929)
         );
  OAI211_X1 U11084 ( .C1(n9984), .C2(n9931), .A(n9930), .B(n9929), .ZN(
        P1_U3245) );
  INV_X1 U11085 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9944) );
  AOI21_X1 U11086 ( .B1(n9992), .B2(n9933), .A(n9932), .ZN(n9943) );
  OAI21_X1 U11087 ( .B1(n9936), .B2(n9935), .A(n9934), .ZN(n9941) );
  OAI21_X1 U11088 ( .B1(n9939), .B2(n9938), .A(n9937), .ZN(n9940) );
  AOI22_X1 U11089 ( .A1(n9998), .A2(n9941), .B1(n9966), .B2(n9940), .ZN(n9942)
         );
  OAI211_X1 U11090 ( .C1(n9984), .C2(n9944), .A(n9943), .B(n9942), .ZN(
        P1_U3248) );
  AOI21_X1 U11091 ( .B1(n9992), .B2(n9946), .A(n9945), .ZN(n9956) );
  OAI21_X1 U11092 ( .B1(n9949), .B2(n9948), .A(n9947), .ZN(n9954) );
  OAI21_X1 U11093 ( .B1(n9952), .B2(n9951), .A(n9950), .ZN(n9953) );
  AOI22_X1 U11094 ( .A1(n9966), .A2(n9954), .B1(n9998), .B2(n9953), .ZN(n9955)
         );
  OAI211_X1 U11095 ( .C1(n8415), .C2(n9984), .A(n9956), .B(n9955), .ZN(
        P1_U3249) );
  INV_X1 U11096 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9970) );
  AOI21_X1 U11097 ( .B1(n9992), .B2(n9958), .A(n9957), .ZN(n9969) );
  OAI21_X1 U11098 ( .B1(n9961), .B2(n9960), .A(n9959), .ZN(n9967) );
  OAI21_X1 U11099 ( .B1(n9964), .B2(n9963), .A(n9962), .ZN(n9965) );
  AOI22_X1 U11100 ( .A1(n9998), .A2(n9967), .B1(n9966), .B2(n9965), .ZN(n9968)
         );
  OAI211_X1 U11101 ( .C1(n9984), .C2(n9970), .A(n9969), .B(n9968), .ZN(
        P1_U3252) );
  INV_X1 U11102 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9983) );
  AOI211_X1 U11103 ( .C1(n9973), .C2(n9972), .A(n9971), .B(n9986), .ZN(n9974)
         );
  AOI211_X1 U11104 ( .C1(n9992), .C2(n9976), .A(n9975), .B(n9974), .ZN(n9982)
         );
  OAI21_X1 U11105 ( .B1(n9979), .B2(n9978), .A(n9977), .ZN(n9980) );
  NAND2_X1 U11106 ( .A1(n9980), .A2(n9998), .ZN(n9981) );
  OAI211_X1 U11107 ( .C1(n9984), .C2(n9983), .A(n9982), .B(n9981), .ZN(
        P1_U3253) );
  INV_X1 U11108 ( .A(n9985), .ZN(n9991) );
  AOI211_X1 U11109 ( .C1(n9989), .C2(n9988), .A(n9987), .B(n9986), .ZN(n9990)
         );
  AOI211_X1 U11110 ( .C1(n9993), .C2(n9992), .A(n9991), .B(n9990), .ZN(n10001)
         );
  OAI21_X1 U11111 ( .B1(n9996), .B2(n9995), .A(n9994), .ZN(n9999) );
  AOI22_X1 U11112 ( .A1(n9999), .A2(n9998), .B1(n9997), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n10000) );
  NAND2_X1 U11113 ( .A1(n10001), .A2(n10000), .ZN(P1_U3259) );
  NAND2_X1 U11114 ( .A1(n10002), .A2(n10027), .ZN(n10004) );
  NAND2_X1 U11115 ( .A1(n10004), .A2(n10003), .ZN(n10005) );
  OR2_X1 U11116 ( .A1(n4462), .A2(n10005), .ZN(n10070) );
  INV_X1 U11117 ( .A(n10070), .ZN(n10007) );
  NAND2_X1 U11118 ( .A1(n10007), .A2(n10006), .ZN(n10030) );
  OAI22_X1 U11119 ( .A1(n9629), .A2(n4736), .B1(n10009), .B2(n10008), .ZN(
        n10026) );
  XNOR2_X1 U11120 ( .A(n10010), .B(n10013), .ZN(n10023) );
  NAND2_X1 U11121 ( .A1(n10012), .A2(n10011), .ZN(n10014) );
  XNOR2_X1 U11122 ( .A(n10014), .B(n10013), .ZN(n10021) );
  OAI22_X1 U11123 ( .A1(n10017), .A2(n10062), .B1(n10016), .B2(n10015), .ZN(
        n10018) );
  INV_X1 U11124 ( .A(n10018), .ZN(n10019) );
  OAI21_X1 U11125 ( .B1(n10021), .B2(n10020), .A(n10019), .ZN(n10022) );
  AOI21_X1 U11126 ( .B1(n10023), .B2(n10066), .A(n10022), .ZN(n10074) );
  NOR2_X1 U11127 ( .A1(n10074), .A2(n10024), .ZN(n10025) );
  AOI211_X1 U11128 ( .C1(n10028), .C2(n10027), .A(n10026), .B(n10025), .ZN(
        n10029) );
  NAND2_X1 U11129 ( .A1(n10030), .A2(n10029), .ZN(P1_U3282) );
  OAI21_X1 U11130 ( .B1(n4509), .B2(n10032), .A(n10031), .ZN(n10033) );
  AOI22_X1 U11131 ( .A1(n10035), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n10034), 
        .B2(n10033), .ZN(n10036) );
  AND2_X1 U11132 ( .A1(n10037), .A2(n10036), .ZN(n10038) );
  AOI22_X1 U11133 ( .A1(n10024), .A2(n10039), .B1(n10038), .B2(n9629), .ZN(
        P1_U3291) );
  AND2_X1 U11134 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10048), .ZN(P1_U3292) );
  AND2_X1 U11135 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10048), .ZN(P1_U3293) );
  AND2_X1 U11136 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10048), .ZN(P1_U3294) );
  NOR2_X1 U11137 ( .A1(n10047), .A2(n10041), .ZN(P1_U3295) );
  AND2_X1 U11138 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10048), .ZN(P1_U3296) );
  AND2_X1 U11139 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10048), .ZN(P1_U3297) );
  NOR2_X1 U11140 ( .A1(n10047), .A2(n10042), .ZN(P1_U3298) );
  AND2_X1 U11141 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10048), .ZN(P1_U3299) );
  NOR2_X1 U11142 ( .A1(n10047), .A2(n10043), .ZN(P1_U3300) );
  AND2_X1 U11143 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10048), .ZN(P1_U3301) );
  AND2_X1 U11144 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10048), .ZN(P1_U3302) );
  AND2_X1 U11145 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10048), .ZN(P1_U3303) );
  AND2_X1 U11146 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10048), .ZN(P1_U3304) );
  AND2_X1 U11147 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10048), .ZN(P1_U3305) );
  AND2_X1 U11148 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10048), .ZN(P1_U3306) );
  AND2_X1 U11149 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10048), .ZN(P1_U3307) );
  NOR2_X1 U11150 ( .A1(n10047), .A2(n10044), .ZN(P1_U3308) );
  AND2_X1 U11151 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10048), .ZN(P1_U3309) );
  AND2_X1 U11152 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10048), .ZN(P1_U3310) );
  AND2_X1 U11153 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10048), .ZN(P1_U3311) );
  NOR2_X1 U11154 ( .A1(n10047), .A2(n10045), .ZN(P1_U3312) );
  AND2_X1 U11155 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10048), .ZN(P1_U3313) );
  AND2_X1 U11156 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10048), .ZN(P1_U3314) );
  NOR2_X1 U11157 ( .A1(n10047), .A2(n10046), .ZN(P1_U3315) );
  AND2_X1 U11158 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10048), .ZN(P1_U3316) );
  AND2_X1 U11159 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10048), .ZN(P1_U3317) );
  AND2_X1 U11160 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10048), .ZN(P1_U3318) );
  AND2_X1 U11161 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10048), .ZN(P1_U3319) );
  AND2_X1 U11162 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10048), .ZN(P1_U3320) );
  AND2_X1 U11163 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10048), .ZN(P1_U3321) );
  OAI21_X1 U11164 ( .B1(n10051), .B2(n10050), .A(n10049), .ZN(P1_U3441) );
  OAI21_X1 U11165 ( .B1(n10053), .B2(n10071), .A(n10052), .ZN(n10055) );
  NOR2_X1 U11166 ( .A1(n10055), .A2(n10054), .ZN(n10078) );
  AOI22_X1 U11167 ( .A1(n10076), .A2(n10078), .B1(n4943), .B2(n10075), .ZN(
        P1_U3457) );
  OAI21_X1 U11168 ( .B1(n10057), .B2(n10071), .A(n10056), .ZN(n10058) );
  INV_X1 U11169 ( .A(n10058), .ZN(n10059) );
  AND2_X1 U11170 ( .A1(n10060), .A2(n10059), .ZN(n10079) );
  AOI22_X1 U11171 ( .A1(n10076), .A2(n10079), .B1(n4991), .B2(n10075), .ZN(
        P1_U3463) );
  OAI22_X1 U11172 ( .A1(n10063), .A2(n10062), .B1(n10061), .B2(n10071), .ZN(
        n10064) );
  AOI211_X1 U11173 ( .C1(n10067), .C2(n10066), .A(n10065), .B(n10064), .ZN(
        n10069) );
  AND2_X1 U11174 ( .A1(n10069), .A2(n10068), .ZN(n10080) );
  AOI22_X1 U11175 ( .A1(n10076), .A2(n10080), .B1(n5052), .B2(n10075), .ZN(
        P1_U3469) );
  OAI21_X1 U11176 ( .B1(n4629), .B2(n10071), .A(n10070), .ZN(n10072) );
  INV_X1 U11177 ( .A(n10072), .ZN(n10073) );
  AND2_X1 U11178 ( .A1(n10074), .A2(n10073), .ZN(n10082) );
  AOI22_X1 U11179 ( .A1(n10076), .A2(n10082), .B1(n5119), .B2(n10075), .ZN(
        P1_U3481) );
  AOI22_X1 U11180 ( .A1(n10083), .A2(n10078), .B1(n10077), .B2(n10081), .ZN(
        P1_U3524) );
  AOI22_X1 U11181 ( .A1(n10083), .A2(n10079), .B1(n4992), .B2(n10081), .ZN(
        P1_U3526) );
  AOI22_X1 U11182 ( .A1(n10083), .A2(n10080), .B1(n5046), .B2(n10081), .ZN(
        P1_U3528) );
  AOI22_X1 U11183 ( .A1(n10083), .A2(n10082), .B1(n6862), .B2(n10081), .ZN(
        P1_U3532) );
  AOI22_X1 U11184 ( .A1(n10138), .A2(n10084), .B1(n10140), .B2(n10137), .ZN(
        n10090) );
  AOI22_X1 U11185 ( .A1(n10136), .A2(n10085), .B1(P2_REG3_REG_7__SCAN_IN), 
        .B2(P2_U3152), .ZN(n10089) );
  OAI211_X1 U11186 ( .C1(n10087), .C2(n10086), .A(n10119), .B(n10145), .ZN(
        n10088) );
  AND3_X1 U11187 ( .A1(n10090), .A2(n10089), .A3(n10088), .ZN(n10091) );
  OAI21_X1 U11188 ( .B1(n10152), .B2(n10092), .A(n10091), .ZN(P2_U3215) );
  AOI22_X1 U11189 ( .A1(n10138), .A2(n10093), .B1(P2_REG3_REG_10__SCAN_IN), 
        .B2(P2_U3152), .ZN(n10094) );
  OAI21_X1 U11190 ( .B1(n10129), .B2(n10095), .A(n10094), .ZN(n10102) );
  INV_X1 U11191 ( .A(n10096), .ZN(n10097) );
  AOI211_X1 U11192 ( .C1(n10100), .C2(n10099), .A(n10098), .B(n10097), .ZN(
        n10101) );
  AOI211_X1 U11193 ( .C1(n10136), .C2(n7345), .A(n10102), .B(n10101), .ZN(
        n10103) );
  OAI21_X1 U11194 ( .B1(n10152), .B2(n10104), .A(n10103), .ZN(P2_U3219) );
  INV_X1 U11195 ( .A(n10105), .ZN(n10106) );
  NAND3_X1 U11196 ( .A1(n10118), .A2(n10111), .A3(n10106), .ZN(n10110) );
  INV_X1 U11197 ( .A(n6817), .ZN(n10108) );
  OAI21_X1 U11198 ( .B1(n10108), .B2(n10107), .A(n10145), .ZN(n10109) );
  NAND2_X1 U11199 ( .A1(n10110), .A2(n10109), .ZN(n10115) );
  AOI22_X1 U11200 ( .A1(n10140), .A2(n10111), .B1(n10138), .B2(n10139), .ZN(
        n10113) );
  NAND2_X1 U11201 ( .A1(n10136), .A2(n6902), .ZN(n10112) );
  OAI211_X1 U11202 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n5966), .A(n10113), .B(
        n10112), .ZN(n10114) );
  AOI21_X1 U11203 ( .B1(n8282), .B2(n10115), .A(n10114), .ZN(n10116) );
  OAI21_X1 U11204 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n10152), .A(n10116), .ZN(
        P2_U3220) );
  NAND3_X1 U11205 ( .A1(n10118), .A2(n10126), .A3(n10117), .ZN(n10124) );
  INV_X1 U11206 ( .A(n10119), .ZN(n10121) );
  OAI21_X1 U11207 ( .B1(n10121), .B2(n10120), .A(n10145), .ZN(n10123) );
  AOI21_X1 U11208 ( .B1(n10124), .B2(n10123), .A(n10122), .ZN(n10132) );
  AOI22_X1 U11209 ( .A1(n10140), .A2(n10126), .B1(n10136), .B2(n10125), .ZN(
        n10128) );
  OAI211_X1 U11210 ( .C1(n10130), .C2(n10129), .A(n10128), .B(n10127), .ZN(
        n10131) );
  NOR2_X1 U11211 ( .A1(n10132), .A2(n10131), .ZN(n10133) );
  OAI21_X1 U11212 ( .B1(n10152), .B2(n10134), .A(n10133), .ZN(P2_U3223) );
  AOI22_X1 U11213 ( .A1(n10136), .A2(n10135), .B1(P2_REG3_REG_5__SCAN_IN), 
        .B2(P2_U3152), .ZN(n10149) );
  NAND2_X1 U11214 ( .A1(n10138), .A2(n10137), .ZN(n10148) );
  NAND2_X1 U11215 ( .A1(n10140), .A2(n10139), .ZN(n10147) );
  NAND2_X1 U11216 ( .A1(n10142), .A2(n10141), .ZN(n10143) );
  NAND3_X1 U11217 ( .A1(n10145), .A2(n10144), .A3(n10143), .ZN(n10146) );
  AND4_X1 U11218 ( .A1(n10149), .A2(n10148), .A3(n10147), .A4(n10146), .ZN(
        n10150) );
  OAI21_X1 U11219 ( .B1(n10152), .B2(n10151), .A(n10150), .ZN(P2_U3229) );
  XOR2_X1 U11220 ( .A(n10153), .B(n10154), .Z(n10157) );
  AOI21_X1 U11221 ( .B1(n10157), .B2(n10156), .A(n10155), .ZN(n10254) );
  INV_X1 U11222 ( .A(n10158), .ZN(n10160) );
  AOI222_X1 U11223 ( .A1(n10162), .A2(n10161), .B1(n10160), .B2(n10159), .C1(
        P2_REG2_REG_12__SCAN_IN), .C2(n4392), .ZN(n10174) );
  AND2_X1 U11224 ( .A1(n10164), .A2(n10163), .ZN(n10167) );
  NAND2_X1 U11225 ( .A1(n10167), .A2(n10166), .ZN(n10165) );
  OAI21_X1 U11226 ( .B1(n10167), .B2(n10166), .A(n10165), .ZN(n10258) );
  OAI211_X1 U11227 ( .C1(n10169), .C2(n10256), .A(n10215), .B(n10168), .ZN(
        n10253) );
  INV_X1 U11228 ( .A(n10253), .ZN(n10170) );
  AOI22_X1 U11229 ( .A1(n10258), .A2(n10172), .B1(n10171), .B2(n10170), .ZN(
        n10173) );
  OAI211_X1 U11230 ( .C1(n4392), .C2(n10254), .A(n10174), .B(n10173), .ZN(
        P2_U3284) );
  AND2_X1 U11231 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10187), .ZN(P2_U3297) );
  AND2_X1 U11232 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10187), .ZN(P2_U3298) );
  AND2_X1 U11233 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10187), .ZN(P2_U3299) );
  AND2_X1 U11234 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10187), .ZN(P2_U3300) );
  AND2_X1 U11235 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10187), .ZN(P2_U3301) );
  AND2_X1 U11236 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10187), .ZN(P2_U3302) );
  AND2_X1 U11237 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10187), .ZN(P2_U3303) );
  NOR2_X1 U11238 ( .A1(n10184), .A2(n10177), .ZN(P2_U3304) );
  AND2_X1 U11239 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10187), .ZN(P2_U3305) );
  AND2_X1 U11240 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10187), .ZN(P2_U3306) );
  AND2_X1 U11241 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10187), .ZN(P2_U3307) );
  AND2_X1 U11242 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10187), .ZN(P2_U3308) );
  AND2_X1 U11243 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10187), .ZN(P2_U3309) );
  AND2_X1 U11244 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10187), .ZN(P2_U3310) );
  NOR2_X1 U11245 ( .A1(n10184), .A2(n10178), .ZN(P2_U3311) );
  AND2_X1 U11246 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10187), .ZN(P2_U3312) );
  AND2_X1 U11247 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10187), .ZN(P2_U3313) );
  AND2_X1 U11248 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10187), .ZN(P2_U3314) );
  AND2_X1 U11249 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10187), .ZN(P2_U3315) );
  AND2_X1 U11250 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10187), .ZN(P2_U3316) );
  NOR2_X1 U11251 ( .A1(n10184), .A2(n10179), .ZN(P2_U3317) );
  NOR2_X1 U11252 ( .A1(n10184), .A2(n10180), .ZN(P2_U3318) );
  AND2_X1 U11253 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10187), .ZN(P2_U3319) );
  NOR2_X1 U11254 ( .A1(n10184), .A2(n10181), .ZN(P2_U3320) );
  NOR2_X1 U11255 ( .A1(n10184), .A2(n10182), .ZN(P2_U3321) );
  NOR2_X1 U11256 ( .A1(n10184), .A2(n10183), .ZN(P2_U3322) );
  AND2_X1 U11257 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10187), .ZN(P2_U3323) );
  AND2_X1 U11258 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10187), .ZN(P2_U3324) );
  AND2_X1 U11259 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10187), .ZN(P2_U3325) );
  AND2_X1 U11260 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10187), .ZN(P2_U3326) );
  AOI22_X1 U11261 ( .A1(n10190), .A2(n10186), .B1(n10185), .B2(n10187), .ZN(
        P2_U3437) );
  AOI22_X1 U11262 ( .A1(n10190), .A2(n10189), .B1(n10188), .B2(n10187), .ZN(
        P2_U3438) );
  AOI22_X1 U11263 ( .A1(n10192), .A2(n10259), .B1(n10191), .B2(n4779), .ZN(
        n10193) );
  AND2_X1 U11264 ( .A1(n10194), .A2(n10193), .ZN(n10262) );
  AOI22_X1 U11265 ( .A1(n4393), .A2(n10262), .B1(n5919), .B2(n10260), .ZN(
        P2_U3451) );
  OAI22_X1 U11266 ( .A1(n10196), .A2(n10248), .B1(n10195), .B2(n10255), .ZN(
        n10199) );
  INV_X1 U11267 ( .A(n10197), .ZN(n10198) );
  AOI211_X1 U11268 ( .C1(n10259), .C2(n10200), .A(n10199), .B(n10198), .ZN(
        n10263) );
  AOI22_X1 U11269 ( .A1(n4393), .A2(n10263), .B1(n5952), .B2(n10260), .ZN(
        P2_U3457) );
  INV_X1 U11270 ( .A(n10201), .ZN(n10203) );
  OAI22_X1 U11271 ( .A1(n10203), .A2(n10248), .B1(n10202), .B2(n10255), .ZN(
        n10206) );
  INV_X1 U11272 ( .A(n10204), .ZN(n10205) );
  AOI211_X1 U11273 ( .C1(n10259), .C2(n10207), .A(n10206), .B(n10205), .ZN(
        n10264) );
  AOI22_X1 U11274 ( .A1(n4393), .A2(n10264), .B1(n5985), .B2(n10260), .ZN(
        P2_U3463) );
  OAI21_X1 U11275 ( .B1(n10209), .B2(n10255), .A(n10208), .ZN(n10211) );
  AOI211_X1 U11276 ( .C1(n10259), .C2(n10212), .A(n10211), .B(n10210), .ZN(
        n10265) );
  AOI22_X1 U11277 ( .A1(n4393), .A2(n10265), .B1(n6001), .B2(n10260), .ZN(
        P2_U3466) );
  AOI22_X1 U11278 ( .A1(n10216), .A2(n10215), .B1(n10214), .B2(n10213), .ZN(
        n10219) );
  NAND3_X1 U11279 ( .A1(n8891), .A2(n10217), .A3(n10259), .ZN(n10218) );
  AND3_X1 U11280 ( .A1(n10220), .A2(n10219), .A3(n10218), .ZN(n10267) );
  AOI22_X1 U11281 ( .A1(n4393), .A2(n10267), .B1(n6020), .B2(n10260), .ZN(
        P2_U3469) );
  INV_X1 U11282 ( .A(n10221), .ZN(n10227) );
  OAI22_X1 U11283 ( .A1(n10223), .A2(n10248), .B1(n10222), .B2(n10255), .ZN(
        n10226) );
  INV_X1 U11284 ( .A(n10224), .ZN(n10225) );
  AOI211_X1 U11285 ( .C1(n10259), .C2(n10227), .A(n10226), .B(n10225), .ZN(
        n10268) );
  AOI22_X1 U11286 ( .A1(n4393), .A2(n10268), .B1(n6039), .B2(n10260), .ZN(
        P2_U3472) );
  INV_X1 U11287 ( .A(n10228), .ZN(n10246) );
  OAI22_X1 U11288 ( .A1(n10230), .A2(n10248), .B1(n10229), .B2(n10255), .ZN(
        n10232) );
  AOI211_X1 U11289 ( .C1(n10246), .C2(n10233), .A(n10232), .B(n10231), .ZN(
        n10269) );
  AOI22_X1 U11290 ( .A1(n4393), .A2(n10269), .B1(n6055), .B2(n10260), .ZN(
        P2_U3475) );
  OAI22_X1 U11291 ( .A1(n10235), .A2(n10248), .B1(n10234), .B2(n10255), .ZN(
        n10238) );
  INV_X1 U11292 ( .A(n10236), .ZN(n10237) );
  AOI211_X1 U11293 ( .C1(n10246), .C2(n10239), .A(n10238), .B(n10237), .ZN(
        n10270) );
  AOI22_X1 U11294 ( .A1(n4393), .A2(n10270), .B1(n6069), .B2(n10260), .ZN(
        P2_U3478) );
  INV_X1 U11295 ( .A(n10240), .ZN(n10245) );
  INV_X1 U11296 ( .A(n7345), .ZN(n10241) );
  OAI22_X1 U11297 ( .A1(n10242), .A2(n10248), .B1(n10241), .B2(n10255), .ZN(
        n10244) );
  AOI211_X1 U11298 ( .C1(n10246), .C2(n10245), .A(n10244), .B(n10243), .ZN(
        n10271) );
  AOI22_X1 U11299 ( .A1(n4393), .A2(n10271), .B1(n6087), .B2(n10260), .ZN(
        P2_U3481) );
  OAI22_X1 U11300 ( .A1(n10249), .A2(n10248), .B1(n10247), .B2(n10255), .ZN(
        n10251) );
  AOI211_X1 U11301 ( .C1(n10252), .C2(n10259), .A(n10251), .B(n10250), .ZN(
        n10272) );
  AOI22_X1 U11302 ( .A1(n4393), .A2(n10272), .B1(n6104), .B2(n10260), .ZN(
        P2_U3484) );
  OAI211_X1 U11303 ( .C1(n10256), .C2(n10255), .A(n10254), .B(n10253), .ZN(
        n10257) );
  AOI21_X1 U11304 ( .B1(n10259), .B2(n10258), .A(n10257), .ZN(n10274) );
  AOI22_X1 U11305 ( .A1(n4393), .A2(n10274), .B1(n6123), .B2(n10260), .ZN(
        P2_U3487) );
  INV_X1 U11306 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10261) );
  AOI22_X1 U11307 ( .A1(n10275), .A2(n10262), .B1(n10261), .B2(n10273), .ZN(
        P2_U3520) );
  AOI22_X1 U11308 ( .A1(n10275), .A2(n10263), .B1(n6631), .B2(n10273), .ZN(
        P2_U3522) );
  AOI22_X1 U11309 ( .A1(n10275), .A2(n10264), .B1(n6633), .B2(n10273), .ZN(
        P2_U3524) );
  AOI22_X1 U11310 ( .A1(n10275), .A2(n10265), .B1(n5999), .B2(n10273), .ZN(
        P2_U3525) );
  INV_X1 U11311 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10266) );
  AOI22_X1 U11312 ( .A1(n10275), .A2(n10267), .B1(n10266), .B2(n10273), .ZN(
        P2_U3526) );
  AOI22_X1 U11313 ( .A1(n10275), .A2(n10268), .B1(n6670), .B2(n10273), .ZN(
        P2_U3527) );
  AOI22_X1 U11314 ( .A1(n10275), .A2(n10269), .B1(n6749), .B2(n10273), .ZN(
        P2_U3528) );
  AOI22_X1 U11315 ( .A1(n10275), .A2(n10270), .B1(n6929), .B2(n10273), .ZN(
        P2_U3529) );
  AOI22_X1 U11316 ( .A1(n10275), .A2(n10271), .B1(n6985), .B2(n10273), .ZN(
        P2_U3530) );
  AOI22_X1 U11317 ( .A1(n10275), .A2(n10272), .B1(n7069), .B2(n10273), .ZN(
        P2_U3531) );
  AOI22_X1 U11318 ( .A1(n10275), .A2(n10274), .B1(n7254), .B2(n10273), .ZN(
        P2_U3532) );
  INV_X1 U11319 ( .A(n10276), .ZN(n10277) );
  NAND2_X1 U11320 ( .A1(n10278), .A2(n10277), .ZN(n10279) );
  XNOR2_X1 U11321 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10279), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11322 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11323 ( .B1(n10282), .B2(n10281), .A(n10280), .ZN(ADD_1071_U56) );
  OAI21_X1 U11324 ( .B1(n10285), .B2(n10284), .A(n10283), .ZN(ADD_1071_U57) );
  OAI21_X1 U11325 ( .B1(n10288), .B2(n10287), .A(n10286), .ZN(ADD_1071_U58) );
  OAI21_X1 U11326 ( .B1(n10291), .B2(n10290), .A(n10289), .ZN(ADD_1071_U59) );
  OAI21_X1 U11327 ( .B1(n10294), .B2(n10293), .A(n10292), .ZN(ADD_1071_U60) );
  OAI21_X1 U11328 ( .B1(n10297), .B2(n10296), .A(n10295), .ZN(ADD_1071_U61) );
  AOI21_X1 U11329 ( .B1(n10300), .B2(n10299), .A(n10298), .ZN(ADD_1071_U62) );
  AOI21_X1 U11330 ( .B1(n10303), .B2(n10302), .A(n10301), .ZN(ADD_1071_U63) );
  AOI21_X1 U11331 ( .B1(n8415), .B2(n10305), .A(n10304), .ZN(ADD_1071_U48) );
  XOR2_X1 U11332 ( .A(n10306), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11333 ( .A1(n10308), .A2(n10307), .ZN(n10309) );
  XOR2_X1 U11334 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10309), .Z(ADD_1071_U51) );
  AOI21_X1 U11335 ( .B1(n10312), .B2(n10311), .A(n10310), .ZN(ADD_1071_U49) );
  OAI21_X1 U11336 ( .B1(n10315), .B2(n10314), .A(n10313), .ZN(n10316) );
  XNOR2_X1 U11337 ( .A(n10316), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11338 ( .B1(n10319), .B2(n10318), .A(n10317), .ZN(ADD_1071_U47) );
  XOR2_X1 U11339 ( .A(n10321), .B(n10320), .Z(ADD_1071_U54) );
  XOR2_X1 U11340 ( .A(n10323), .B(n10322), .Z(ADD_1071_U53) );
  XNOR2_X1 U11341 ( .A(n10325), .B(n10324), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4919 ( .A(n5598), .Z(n4388) );
endmodule

