

module b22_C_gen_AntiSAT_k_256_9 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, 
        keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, 
        keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, 
        keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, 
        keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, 
        keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, 
        keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, 
        keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, 
        keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104, 
        keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108, 
        keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112, 
        keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116, 
        keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120, 
        keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124, 
        keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, 
        keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, 
        keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, 
        keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, 
        keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, 
        keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, 
        keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, 
        keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0,
         keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5,
         keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10,
         keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15,
         keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20,
         keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25,
         keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30,
         keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35,
         keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40,
         keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45,
         keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50,
         keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55,
         keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60,
         keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65,
         keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70,
         keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75,
         keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80,
         keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85,
         keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90,
         keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95,
         keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100,
         keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104,
         keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108,
         keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112,
         keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116,
         keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120,
         keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124,
         keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66,
         keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71,
         keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76,
         keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81,
         keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86,
         keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91,
         keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96,
         keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100,
         keyinput_g101, keyinput_g102, keyinput_g103, keyinput_g104,
         keyinput_g105, keyinput_g106, keyinput_g107, keyinput_g108,
         keyinput_g109, keyinput_g110, keyinput_g111, keyinput_g112,
         keyinput_g113, keyinput_g114, keyinput_g115, keyinput_g116,
         keyinput_g117, keyinput_g118, keyinput_g119, keyinput_g120,
         keyinput_g121, keyinput_g122, keyinput_g123, keyinput_g124,
         keyinput_g125, keyinput_g126, keyinput_g127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6667, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871;

  INV_X4 U7415 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NAND2_X1 U7416 ( .A1(n7465), .A2(n7464), .ZN(n14134) );
  CLKBUF_X1 U7418 ( .A(n7966), .Z(n11717) );
  INV_X2 U7419 ( .A(n12862), .ZN(n9838) );
  CLKBUF_X2 U7420 ( .A(n6669), .Z(n13044) );
  INV_X1 U7421 ( .A(n13228), .ZN(n13221) );
  NAND4_X1 U7422 ( .A1(n7879), .A2(n7877), .A3(n7878), .A4(n7880), .ZN(n11400)
         );
  OR2_X2 U7423 ( .A1(n10511), .A2(n9931), .ZN(n15061) );
  XNOR2_X1 U7424 ( .A(n9212), .B(n9211), .ZN(n9263) );
  NAND2_X1 U7425 ( .A1(n9210), .A2(n9209), .ZN(n9212) );
  BUF_X1 U7426 ( .A(n8535), .Z(n6680) );
  XOR2_X1 U7427 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n9553), .Z(n9264) );
  AND2_X1 U7428 ( .A1(n8417), .A2(n8416), .ZN(n8464) );
  XNOR2_X1 U7429 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n6878) );
  AND2_X2 U7430 ( .A1(n8387), .A2(n7747), .ZN(n9748) );
  INV_X1 U7431 ( .A(n9162), .ZN(n14272) );
  MUX2_X1 U7432 ( .A(n7693), .B(n15107), .S(n9963), .Z(n11506) );
  INV_X2 U7433 ( .A(n10024), .ZN(n9951) );
  NOR2_X1 U7436 ( .A1(n14090), .A2(n14292), .ZN(n14077) );
  INV_X1 U7437 ( .A(n10760), .ZN(n8884) );
  AND2_X1 U7439 ( .A1(n10760), .A2(n10717), .ZN(n8535) );
  INV_X1 U7440 ( .A(n6681), .ZN(n8510) );
  NAND2_X1 U7441 ( .A1(n10175), .A2(n10174), .ZN(n15386) );
  OR2_X1 U7442 ( .A1(n14863), .A2(n14859), .ZN(n7758) );
  OAI21_X1 U7443 ( .B1(n9079), .B2(n7671), .A(n7670), .ZN(n9100) );
  NAND2_X1 U7444 ( .A1(n7235), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7234) );
  AOI21_X1 U7445 ( .B1(n11975), .B2(n11974), .A(n7751), .ZN(n12026) );
  CLKBUF_X3 U7446 ( .A(n7993), .Z(n6669) );
  XNOR2_X1 U7447 ( .A(n7848), .B(P3_IR_REG_29__SCAN_IN), .ZN(n7849) );
  NAND2_X1 U7448 ( .A1(n7594), .A2(n7589), .ZN(n9178) );
  NAND2_X1 U7449 ( .A1(n8886), .A2(n8885), .ZN(n14345) );
  AND2_X1 U7450 ( .A1(n8373), .A2(n7439), .ZN(n9747) );
  NAND2_X1 U7451 ( .A1(n10210), .A2(n10209), .ZN(n15064) );
  AND2_X1 U7452 ( .A1(n14989), .A2(n14773), .ZN(n14727) );
  NAND2_X1 U7453 ( .A1(n10487), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7568) );
  INV_X1 U7454 ( .A(n14922), .ZN(n15509) );
  AND2_X1 U7455 ( .A1(n12952), .A2(n6740), .ZN(n6667) );
  INV_X2 U7456 ( .A(n15731), .ZN(n15729) );
  NOR2_X2 U7457 ( .A1(n7585), .A2(n10185), .ZN(n7584) );
  NOR2_X2 U7458 ( .A1(n15855), .A2(n9273), .ZN(n9275) );
  OAI21_X2 U7459 ( .B1(n6692), .B2(n13234), .A(n13233), .ZN(n13235) );
  NAND3_X2 U7460 ( .A1(n9946), .A2(n9945), .A3(n9944), .ZN(n11443) );
  AND2_X2 U7461 ( .A1(n9943), .A2(n9942), .ZN(n9945) );
  INV_X2 U7462 ( .A(n7043), .ZN(n11110) );
  AND2_X2 U7463 ( .A1(n8276), .A2(n8279), .ZN(n12496) );
  OAI21_X2 U7464 ( .B1(n8764), .B2(n8763), .A(n8762), .ZN(n8765) );
  NOR2_X1 U7465 ( .A1(n11736), .A2(n7764), .ZN(n11793) );
  OAI21_X2 U7466 ( .B1(n14195), .B2(n6783), .A(n9672), .ZN(n14180) );
  XNOR2_X1 U7467 ( .A(n13944), .B(n11125), .ZN(n11093) );
  NAND2_X2 U7468 ( .A1(n8512), .A2(n7531), .ZN(n11125) );
  XNOR2_X2 U7469 ( .A(n9215), .B(n9407), .ZN(n9262) );
  NOR3_X2 U7470 ( .A1(n9979), .A2(n10185), .A3(n6893), .ZN(n6892) );
  NAND4_X2 U7471 ( .A1(n9961), .A2(n7693), .A3(n9948), .A4(n9887), .ZN(n9979)
         );
  NAND2_X2 U7472 ( .A1(n6872), .A2(n9214), .ZN(n9215) );
  INV_X1 U7473 ( .A(n9906), .ZN(n12706) );
  INV_X1 U7474 ( .A(n9178), .ZN(n15698) );
  INV_X4 U7475 ( .A(n10512), .ZN(n12846) );
  NAND2_X2 U7476 ( .A1(n15085), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9900) );
  XNOR2_X2 U7477 ( .A(n7568), .B(P1_IR_REG_22__SCAN_IN), .ZN(n10412) );
  NAND4_X2 U7479 ( .A1(n8518), .A2(n8517), .A3(n8516), .A4(n8515), .ZN(n13944)
         );
  AOI211_X1 U7480 ( .C1(n14067), .C2(n15269), .A(n14066), .B(n14065), .ZN(
        n14068) );
  NOR2_X2 U7481 ( .A1(n14941), .A2(n15052), .ZN(n14905) );
  NAND2_X2 U7482 ( .A1(n10258), .A2(n10257), .ZN(n15052) );
  AOI211_X2 U7483 ( .C1(n14958), .C2(n14997), .A(n14784), .B(n14783), .ZN(
        n14785) );
  XNOR2_X2 U7484 ( .A(n9100), .B(n9099), .ZN(n14415) );
  XNOR2_X2 U7485 ( .A(n13783), .B(n13945), .ZN(n11568) );
  AOI21_X2 U7486 ( .B1(n12910), .B2(n7394), .A(n7395), .ZN(n13022) );
  OAI21_X2 U7487 ( .B1(n13536), .B2(n13192), .A(n13191), .ZN(n13522) );
  NAND2_X2 U7488 ( .A1(n7845), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7832) );
  OAI21_X2 U7489 ( .B1(n9778), .B2(n13238), .A(n9779), .ZN(n6679) );
  XNOR2_X1 U7490 ( .A(n7834), .B(n7833), .ZN(n6670) );
  XNOR2_X1 U7491 ( .A(n7834), .B(n7833), .ZN(n6671) );
  INV_X1 U7492 ( .A(n10612), .ZN(n6672) );
  XNOR2_X1 U7493 ( .A(n7834), .B(n7833), .ZN(n8267) );
  OR2_X1 U7494 ( .A1(n15808), .A2(n9789), .ZN(n13108) );
  OAI21_X2 U7495 ( .B1(n8087), .B2(n7642), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n7834) );
  OAI22_X1 U7496 ( .A1(n13770), .A2(n13769), .B1(n6811), .B2(n13752), .ZN(
        n13853) );
  NAND2_X1 U7497 ( .A1(n7372), .A2(n9844), .ZN(n9846) );
  NAND2_X1 U7498 ( .A1(n14125), .A2(n14385), .ZN(n14104) );
  NAND2_X1 U7499 ( .A1(n12483), .A2(n7529), .ZN(n14363) );
  NAND2_X1 U7500 ( .A1(n12099), .A2(n12098), .ZN(n12183) );
  NAND2_X1 U7501 ( .A1(n12265), .A2(n6957), .ZN(n12450) );
  NAND2_X2 U7502 ( .A1(n15061), .A2(n12846), .ZN(n12788) );
  INV_X1 U7503 ( .A(n13804), .ZN(n14078) );
  INV_X4 U7504 ( .A(n8469), .ZN(n9124) );
  INV_X8 U7505 ( .A(n8582), .ZN(n6673) );
  NAND2_X2 U7506 ( .A1(n9748), .A2(n12707), .ZN(n10957) );
  NAND2_X4 U7507 ( .A1(n8266), .A2(n6670), .ZN(n8268) );
  INV_X1 U7508 ( .A(n10404), .ZN(n10417) );
  NAND2_X4 U7509 ( .A1(n10501), .A2(n15094), .ZN(n9963) );
  XNOR2_X1 U7510 ( .A(n14726), .B(n14725), .ZN(n14992) );
  AOI21_X1 U7511 ( .B1(n15003), .B2(n15549), .A(n15002), .ZN(n15004) );
  AND2_X1 U7512 ( .A1(n6920), .A2(n6919), .ZN(n14379) );
  NAND2_X1 U7513 ( .A1(n14540), .A2(n14541), .ZN(n14539) );
  AND2_X1 U7514 ( .A1(n14298), .A2(n6921), .ZN(n6920) );
  OR2_X1 U7515 ( .A1(n9015), .A2(n9014), .ZN(n9055) );
  NOR2_X1 U7516 ( .A1(n14051), .A2(n15263), .ZN(n14280) );
  AOI21_X1 U7517 ( .B1(n14087), .B2(n15256), .A(n14086), .ZN(n14298) );
  AND2_X1 U7518 ( .A1(n7445), .A2(n6732), .ZN(n13904) );
  NAND2_X1 U7519 ( .A1(n6667), .A2(n9847), .ZN(n12922) );
  NAND2_X1 U7520 ( .A1(n7443), .A2(n7448), .ZN(n7446) );
  NAND2_X1 U7521 ( .A1(n14085), .A2(n14088), .ZN(n14084) );
  AND2_X1 U7522 ( .A1(n12921), .A2(n12923), .ZN(n9849) );
  OR2_X1 U7523 ( .A1(n9846), .A2(n9845), .ZN(n9847) );
  AOI21_X1 U7524 ( .B1(n6867), .B2(n6866), .A(n13231), .ZN(n6865) );
  AND2_X1 U7525 ( .A1(n14832), .A2(n7286), .ZN(n14773) );
  AND2_X1 U7526 ( .A1(n7161), .A2(n6990), .ZN(n6989) );
  OR2_X1 U7527 ( .A1(n14292), .A2(n13763), .ZN(n9736) );
  NAND2_X2 U7528 ( .A1(n9064), .A2(n9063), .ZN(n14292) );
  AOI21_X1 U7529 ( .B1(n6704), .B2(n7251), .A(n7247), .ZN(n7246) );
  NAND2_X1 U7530 ( .A1(n9082), .A2(n9081), .ZN(n14091) );
  NOR2_X1 U7531 ( .A1(n15140), .A2(n15139), .ZN(n15138) );
  NAND2_X1 U7532 ( .A1(n14888), .A2(n14713), .ZN(n14876) );
  NAND2_X1 U7533 ( .A1(n7036), .A2(n7034), .ZN(n13815) );
  OAI21_X1 U7534 ( .B1(n6907), .B2(n7317), .A(n6905), .ZN(n8207) );
  NAND2_X1 U7535 ( .A1(n12890), .A2(n9833), .ZN(n12967) );
  NAND2_X1 U7536 ( .A1(n6877), .A2(n15435), .ZN(n15440) );
  NAND2_X1 U7537 ( .A1(n9003), .A2(n9002), .ZN(n14316) );
  AOI21_X1 U7538 ( .B1(n14864), .B2(n7704), .A(n7703), .ZN(n7702) );
  OR2_X1 U7539 ( .A1(n14215), .A2(n9720), .ZN(n14212) );
  NAND2_X1 U7540 ( .A1(n6931), .A2(n7528), .ZN(n6930) );
  NAND2_X1 U7541 ( .A1(n7264), .A2(n6741), .ZN(n7413) );
  NAND2_X1 U7542 ( .A1(n7478), .A2(n7477), .ZN(n12742) );
  XNOR2_X1 U7543 ( .A(n9017), .B(SI_24_), .ZN(n9020) );
  AND2_X1 U7544 ( .A1(n7607), .A2(n7611), .ZN(n15254) );
  NAND2_X1 U7545 ( .A1(n9001), .A2(n9000), .ZN(n9017) );
  AND2_X1 U7546 ( .A1(n9711), .A2(n13934), .ZN(n6684) );
  AND2_X1 U7547 ( .A1(n10271), .A2(n10270), .ZN(n14911) );
  OAI22_X1 U7548 ( .A1(n7047), .A2(n7048), .B1(n12183), .B2(n7054), .ZN(n13719) );
  NAND2_X1 U7549 ( .A1(n15213), .A2(n13162), .ZN(n15203) );
  NAND2_X1 U7550 ( .A1(n11900), .A2(n7456), .ZN(n12099) );
  NAND2_X1 U7551 ( .A1(n7016), .A2(n11765), .ZN(n11900) );
  OAI21_X1 U7552 ( .B1(n11648), .B2(n7587), .A(n7106), .ZN(n7105) );
  NAND2_X1 U7553 ( .A1(n12151), .A2(n9799), .ZN(n12267) );
  NAND2_X1 U7554 ( .A1(n7107), .A2(n9699), .ZN(n11648) );
  NAND2_X1 U7555 ( .A1(n11745), .A2(n7017), .ZN(n11763) );
  NAND2_X1 U7556 ( .A1(n6841), .A2(n7320), .ZN(n12318) );
  NAND2_X1 U7557 ( .A1(n11485), .A2(n11484), .ZN(n11745) );
  NAND2_X1 U7558 ( .A1(n8769), .A2(n8768), .ZN(n15280) );
  NAND2_X1 U7559 ( .A1(n11959), .A2(n13137), .ZN(n12282) );
  NAND2_X1 U7560 ( .A1(n10629), .A2(n10628), .ZN(n12424) );
  OR2_X1 U7561 ( .A1(n11808), .A2(n11879), .ZN(n11856) );
  NAND2_X1 U7562 ( .A1(n10093), .A2(n10092), .ZN(n12554) );
  NAND2_X1 U7563 ( .A1(n8642), .A2(n8641), .ZN(n11879) );
  NAND2_X1 U7564 ( .A1(n15862), .A2(n9286), .ZN(n9288) );
  OAI211_X1 U7565 ( .C1(n7241), .C2(n12849), .A(n7237), .B(n7236), .ZN(n11668)
         );
  NAND2_X1 U7566 ( .A1(n7646), .A2(n7644), .ZN(n8665) );
  AND2_X1 U7567 ( .A1(n7470), .A2(n11563), .ZN(n11386) );
  OR2_X1 U7568 ( .A1(n8186), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8199) );
  AOI21_X1 U7569 ( .B1(n11417), .B2(n11416), .A(n11415), .ZN(n11707) );
  XNOR2_X1 U7570 ( .A(n9281), .B(n9280), .ZN(n15126) );
  INV_X1 U7571 ( .A(n11696), .ZN(n12083) );
  OR2_X1 U7572 ( .A1(n10536), .A2(n15513), .ZN(n11913) );
  NAND2_X1 U7573 ( .A1(n8541), .A2(n8540), .ZN(n11590) );
  NAND2_X1 U7574 ( .A1(n15858), .A2(n9277), .ZN(n9281) );
  NAND2_X2 U7575 ( .A1(n8454), .A2(n8453), .ZN(n13783) );
  INV_X1 U7576 ( .A(n8214), .ZN(n15785) );
  INV_X2 U7577 ( .A(n9850), .ZN(n12862) );
  OAI211_X1 U7578 ( .C1(n8469), .C2(n8440), .A(n8478), .B(n7755), .ZN(n11109)
         );
  INV_X4 U7579 ( .A(n10689), .ZN(P3_U3897) );
  CLKBUF_X3 U7580 ( .A(n11110), .Z(n13806) );
  INV_X4 U7581 ( .A(n6673), .ZN(n9114) );
  NAND2_X1 U7582 ( .A1(n8446), .A2(n8447), .ZN(n8503) );
  NAND4_X1 U7583 ( .A1(n7902), .A2(n7901), .A3(n7900), .A4(n7899), .ZN(n11796)
         );
  NAND4_X1 U7584 ( .A1(n8429), .A2(n8428), .A3(n8427), .A4(n8426), .ZN(n13947)
         );
  NAND4_X1 U7585 ( .A1(n8468), .A2(n8467), .A3(n8466), .A4(n8465), .ZN(n13946)
         );
  OR2_X2 U7586 ( .A1(n10509), .A2(n10508), .ZN(n12787) );
  NAND2_X1 U7587 ( .A1(n10429), .A2(n9929), .ZN(n10024) );
  BUF_X2 U7588 ( .A(n8535), .Z(n6681) );
  BUF_X2 U7589 ( .A(n7898), .Z(n8346) );
  INV_X2 U7590 ( .A(n10110), .ZN(n10423) );
  NAND4_X1 U7591 ( .A1(n9937), .A2(n9936), .A3(n9935), .A4(n9934), .ZN(n14563)
         );
  INV_X2 U7592 ( .A(n13050), .ZN(n6677) );
  NAND2_X1 U7593 ( .A1(n8439), .A2(SI_2_), .ZN(n8444) );
  NAND2_X2 U7594 ( .A1(n9963), .A2(n10717), .ZN(n10424) );
  NAND2_X2 U7595 ( .A1(n15690), .A2(n12707), .ZN(n15263) );
  INV_X2 U7596 ( .A(n8464), .ZN(n9130) );
  NOR2_X1 U7597 ( .A1(n10764), .A2(P2_U3088), .ZN(P2_U3947) );
  NAND2_X1 U7598 ( .A1(n8268), .A2(n10717), .ZN(n7993) );
  CLKBUF_X2 U7599 ( .A(n10380), .Z(n6674) );
  AND2_X1 U7600 ( .A1(n8417), .A2(n14412), .ZN(n8542) );
  CLKBUF_X2 U7601 ( .A(n10380), .Z(n6675) );
  INV_X1 U7602 ( .A(n11788), .ZN(n13105) );
  XNOR2_X1 U7603 ( .A(n8280), .B(P3_IR_REG_26__SCAN_IN), .ZN(n13707) );
  XNOR2_X1 U7604 ( .A(n8277), .B(P3_IR_REG_25__SCAN_IN), .ZN(n8282) );
  XNOR2_X1 U7605 ( .A(n6913), .B(P3_IR_REG_30__SCAN_IN), .ZN(n7850) );
  NAND2_X1 U7606 ( .A1(n6970), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8280) );
  NAND2_X1 U7607 ( .A1(n8279), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8277) );
  XNOR2_X1 U7608 ( .A(n7114), .B(n7113), .ZN(n14412) );
  XNOR2_X1 U7609 ( .A(n8413), .B(n8412), .ZN(n8415) );
  XNOR2_X1 U7610 ( .A(n8378), .B(n8377), .ZN(n9162) );
  INV_X2 U7611 ( .A(n15090), .ZN(n15104) );
  NAND2_X1 U7612 ( .A1(n13689), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6913) );
  XNOR2_X1 U7613 ( .A(n8382), .B(n8381), .ZN(n12707) );
  NAND2_X1 U7614 ( .A1(n8397), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U7615 ( .A1(n8211), .A2(n6688), .ZN(n11788) );
  NAND2_X1 U7616 ( .A1(n8399), .A2(n8400), .ZN(n10767) );
  XNOR2_X1 U7617 ( .A(n7782), .B(n7781), .ZN(n13393) );
  NAND2_X1 U7618 ( .A1(n8414), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7114) );
  OR2_X1 U7619 ( .A1(n14405), .A2(n14406), .ZN(n8413) );
  OR2_X1 U7620 ( .A1(n8396), .A2(n7738), .ZN(n8400) );
  XNOR2_X1 U7621 ( .A(n9903), .B(n9902), .ZN(n9904) );
  NAND2_X1 U7622 ( .A1(n7501), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9918) );
  MUX2_X1 U7623 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7776), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n7779) );
  OR2_X1 U7624 ( .A1(n9926), .A2(n10013), .ZN(n7233) );
  INV_X4 U7625 ( .A(n9919), .ZN(n10717) );
  OAI21_X1 U7626 ( .B1(n6972), .B2(n6776), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n7776) );
  OR2_X1 U7627 ( .A1(n6972), .A2(n7400), .ZN(n7780) );
  NOR2_X1 U7628 ( .A1(n7642), .A2(P3_IR_REG_27__SCAN_IN), .ZN(n7640) );
  CLKBUF_X1 U7629 ( .A(n8087), .Z(n6972) );
  NAND2_X1 U7630 ( .A1(n7431), .A2(n7883), .ZN(n11023) );
  NOR2_X1 U7631 ( .A1(n8087), .A2(P3_IR_REG_28__SCAN_IN), .ZN(n7332) );
  NOR2_X1 U7632 ( .A1(n7368), .A2(n6777), .ZN(n9901) );
  NAND2_X1 U7633 ( .A1(n8009), .A2(n7775), .ZN(n8087) );
  INV_X1 U7634 ( .A(n7778), .ZN(n7338) );
  INV_X1 U7635 ( .A(n7585), .ZN(n6891) );
  AND2_X1 U7636 ( .A1(n7775), .A2(n7918), .ZN(n6966) );
  NAND2_X1 U7637 ( .A1(n7367), .A2(n6894), .ZN(n6893) );
  AND3_X1 U7638 ( .A1(n6898), .A2(n6897), .A3(n6899), .ZN(n7771) );
  AND4_X1 U7639 ( .A1(n7774), .A2(n7773), .A3(n8022), .A4(n7772), .ZN(n7775)
         );
  AND3_X1 U7640 ( .A1(n7403), .A2(n8118), .A3(n7781), .ZN(n7757) );
  AND4_X1 U7641 ( .A1(n9896), .A2(n9895), .A3(n9894), .A4(n9893), .ZN(n9897)
         );
  NAND2_X1 U7642 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n6978), .ZN(n6977) );
  INV_X1 U7643 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9961) );
  INV_X4 U7644 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X2 U7645 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U7646 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n6898) );
  NOR2_X1 U7647 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_5__SCAN_IN), .ZN(
        n6897) );
  NOR2_X1 U7648 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n7370) );
  INV_X1 U7649 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7369) );
  INV_X1 U7650 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7770) );
  INV_X1 U7651 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n9553) );
  INV_X1 U7652 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7403) );
  NOR2_X1 U7653 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n7067) );
  INV_X1 U7654 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8393) );
  NOR2_X1 U7655 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n9892) );
  INV_X1 U7656 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7781) );
  NOR2_X1 U7657 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n7060) );
  NOR2_X1 U7658 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n7061) );
  NOR2_X1 U7659 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n7062) );
  INV_X1 U7660 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n7367) );
  INV_X1 U7661 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6894) );
  NOR2_X1 U7662 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n7773) );
  NOR2_X1 U7663 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n7774) );
  INV_X1 U7664 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8412) );
  NOR2_X1 U7665 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n9888) );
  XNOR2_X2 U7666 ( .A(n12658), .B(n12547), .ZN(n12663) );
  OAI21_X2 U7667 ( .B1(n12054), .B2(n7349), .A(n7346), .ZN(n12298) );
  NAND2_X1 U7668 ( .A1(n7345), .A2(n9906), .ZN(n10380) );
  INV_X1 U7669 ( .A(n13050), .ZN(n6676) );
  OAI21_X2 U7670 ( .B1(n14103), .B2(n9680), .A(n7513), .ZN(n14089) );
  CLKBUF_X1 U7671 ( .A(n15094), .Z(n6678) );
  XNOR2_X1 U7672 ( .A(n9918), .B(n9917), .ZN(n15094) );
  OAI21_X2 U7673 ( .B1(n12988), .B2(n12991), .A(n12989), .ZN(n12910) );
  NOR2_X2 U7674 ( .A1(n9810), .A2(n9809), .ZN(n12988) );
  NOR2_X2 U7675 ( .A1(n14258), .A2(n14353), .ZN(n7467) );
  NAND2_X1 U7676 ( .A1(n10713), .A2(n8535), .ZN(n8478) );
  XNOR2_X2 U7677 ( .A(n8394), .B(n8410), .ZN(n9203) );
  OAI21_X2 U7678 ( .B1(n9778), .B2(n13238), .A(n9779), .ZN(n9850) );
  INV_X2 U7679 ( .A(n11109), .ZN(n6915) );
  NOR2_X1 U7680 ( .A1(n7134), .A2(n7141), .ZN(n7131) );
  NAND2_X1 U7681 ( .A1(n8900), .A2(n8899), .ZN(n8907) );
  OAI21_X1 U7682 ( .B1(n13522), .B2(n6903), .A(n6778), .ZN(n13477) );
  OR2_X1 U7683 ( .A1(n6903), .A2(n7322), .ZN(n6902) );
  NAND2_X1 U7684 ( .A1(n6904), .A2(n13202), .ZN(n6903) );
  NAND2_X1 U7685 ( .A1(n7428), .A2(n7427), .ZN(n13247) );
  INV_X1 U7686 ( .A(n12415), .ZN(n7427) );
  NAND2_X1 U7687 ( .A1(n7413), .A2(n13284), .ZN(n13318) );
  OR2_X1 U7688 ( .A1(n13050), .A2(n7761), .ZN(n7886) );
  NAND2_X1 U7689 ( .A1(n10499), .A2(n10558), .ZN(n10543) );
  AND2_X1 U7690 ( .A1(n10561), .A2(n10559), .ZN(n10499) );
  NAND2_X1 U7691 ( .A1(n14840), .A2(n14721), .ZN(n14808) );
  AND2_X1 U7692 ( .A1(n8423), .A2(n8422), .ZN(n8485) );
  NAND2_X1 U7693 ( .A1(n7742), .A2(n6739), .ZN(n7741) );
  INV_X1 U7694 ( .A(n8921), .ZN(n7085) );
  INV_X1 U7695 ( .A(n7087), .ZN(n7086) );
  OAI21_X1 U7696 ( .B1(n7088), .B2(n8876), .A(n7739), .ZN(n7087) );
  NAND2_X1 U7697 ( .A1(n8896), .A2(n7740), .ZN(n7739) );
  INV_X1 U7698 ( .A(n6739), .ZN(n7740) );
  INV_X1 U7699 ( .A(n8854), .ZN(n7730) );
  INV_X1 U7700 ( .A(n7601), .ZN(n7600) );
  OAI21_X1 U7701 ( .B1(n12486), .B2(n7602), .A(n9716), .ZN(n7601) );
  NAND2_X1 U7702 ( .A1(n12517), .A2(n9808), .ZN(n9810) );
  NAND2_X1 U7703 ( .A1(n11146), .A2(n10595), .ZN(n11025) );
  NAND2_X1 U7704 ( .A1(n7423), .A2(n7422), .ZN(n11203) );
  INV_X1 U7705 ( .A(n10597), .ZN(n7423) );
  NAND2_X1 U7706 ( .A1(n10596), .A2(n11209), .ZN(n7422) );
  AND2_X1 U7707 ( .A1(n7282), .A2(n7281), .ZN(n10596) );
  AND2_X1 U7708 ( .A1(n12411), .A2(n12410), .ZN(n12412) );
  OAI21_X1 U7709 ( .B1(n13258), .B2(n13257), .A(n13256), .ZN(n13259) );
  AND2_X1 U7710 ( .A1(n7269), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7268) );
  NAND3_X1 U7711 ( .A1(n7151), .A2(n6703), .A3(n7150), .ZN(n7421) );
  INV_X1 U7712 ( .A(n13083), .ZN(n7319) );
  NAND2_X1 U7713 ( .A1(n13659), .A2(n13466), .ZN(n13460) );
  AOI21_X1 U7714 ( .B1(n13525), .B2(n13197), .A(n6754), .ZN(n7325) );
  INV_X1 U7715 ( .A(n7321), .ZN(n7320) );
  NAND2_X1 U7716 ( .A1(n12282), .A2(n6912), .ZN(n6841) );
  OAI21_X1 U7717 ( .B1(n7985), .B2(n6712), .A(n8000), .ZN(n7321) );
  INV_X1 U7718 ( .A(n7230), .ZN(n7823) );
  OAI21_X1 U7719 ( .B1(n8173), .B2(n8172), .A(n6830), .ZN(n7230) );
  INV_X1 U7720 ( .A(n7547), .ZN(n7546) );
  OAI21_X1 U7721 ( .B1(n8069), .B2(n7548), .A(n8084), .ZN(n7547) );
  NAND2_X1 U7722 ( .A1(n7218), .A2(n7217), .ZN(n7809) );
  NAND2_X1 U7723 ( .A1(n6698), .A2(n7221), .ZN(n7217) );
  OR2_X1 U7724 ( .A1(n8021), .A2(n7219), .ZN(n7218) );
  INV_X1 U7725 ( .A(n14412), .ZN(n8416) );
  INV_X1 U7726 ( .A(n7527), .ZN(n6929) );
  INV_X1 U7727 ( .A(n9710), .ZN(n7612) );
  NOR4_X1 U7728 ( .A1(n10447), .A2(n14982), .A3(n14690), .A4(n10446), .ZN(
        n10448) );
  NOR2_X1 U7729 ( .A1(n14802), .A2(n14762), .ZN(n7288) );
  NAND2_X1 U7730 ( .A1(n7681), .A2(n7680), .ZN(n14932) );
  AOI21_X1 U7731 ( .B1(n6682), .B2(n7687), .A(n7682), .ZN(n7681) );
  INV_X1 U7732 ( .A(n14744), .ZN(n7682) );
  AOI21_X1 U7733 ( .B1(n9126), .B2(n9125), .A(n9102), .ZN(n9116) );
  AND2_X1 U7734 ( .A1(n7174), .A2(n7170), .ZN(n7169) );
  AND2_X1 U7735 ( .A1(n7179), .A2(n8977), .ZN(n7174) );
  NAND2_X1 U7736 ( .A1(n8907), .A2(n8906), .ZN(n8959) );
  AND2_X1 U7737 ( .A1(n8831), .A2(n8811), .ZN(n8829) );
  AND2_X1 U7738 ( .A1(n8807), .A2(n8785), .ZN(n8805) );
  NAND2_X2 U7739 ( .A1(n7840), .A2(n7839), .ZN(n8405) );
  NAND2_X1 U7740 ( .A1(n12967), .A2(n7392), .ZN(n12901) );
  NOR2_X1 U7741 ( .A1(n12904), .A2(n7393), .ZN(n7392) );
  INV_X1 U7742 ( .A(n9835), .ZN(n7393) );
  OAI21_X1 U7743 ( .B1(n13235), .B2(n13236), .A(n6849), .ZN(n6848) );
  OR2_X1 U7744 ( .A1(n13237), .A2(n13238), .ZN(n6849) );
  NOR3_X1 U7745 ( .A1(n13234), .A2(n13080), .A3(n13079), .ZN(n13082) );
  XNOR2_X1 U7746 ( .A(n6843), .B(n13081), .ZN(n6842) );
  NAND2_X1 U7747 ( .A1(n6911), .A2(n6975), .ZN(n6843) );
  INV_X1 U7748 ( .A(n6976), .ZN(n6975) );
  OAI211_X1 U7749 ( .C1(n13056), .C2(n13232), .A(n13055), .B(n13054), .ZN(
        n6911) );
  NAND2_X1 U7750 ( .A1(n7149), .A2(n7148), .ZN(n7147) );
  INV_X1 U7751 ( .A(n11286), .ZN(n7148) );
  OR2_X1 U7752 ( .A1(n11306), .A2(n11307), .ZN(n7144) );
  NAND2_X1 U7753 ( .A1(n7405), .A2(n7404), .ZN(n11411) );
  INV_X1 U7754 ( .A(n11408), .ZN(n7404) );
  INV_X1 U7755 ( .A(n11405), .ZN(n7418) );
  NOR2_X1 U7756 ( .A1(n11703), .A2(n10675), .ZN(n11702) );
  OR2_X1 U7757 ( .A1(n15743), .A2(n8015), .ZN(n7263) );
  XNOR2_X1 U7758 ( .A(n12412), .B(n12425), .ZN(n15743) );
  NOR2_X1 U7759 ( .A1(n13260), .A2(n15190), .ZN(n13277) );
  INV_X1 U7760 ( .A(n6988), .ZN(n13267) );
  NAND2_X1 U7761 ( .A1(n7421), .A2(n7420), .ZN(n13364) );
  NAND2_X1 U7762 ( .A1(n13362), .A2(n13361), .ZN(n7420) );
  NAND2_X1 U7763 ( .A1(n13335), .A2(n13334), .ZN(n13362) );
  NOR2_X1 U7764 ( .A1(n8261), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n15162) );
  AND2_X1 U7765 ( .A1(n7624), .A2(n6973), .ZN(n13410) );
  NOR2_X1 U7766 ( .A1(n13407), .A2(n6735), .ZN(n6973) );
  NAND2_X1 U7767 ( .A1(n6946), .A2(n6949), .ZN(n7628) );
  XNOR2_X1 U7768 ( .A(n13224), .B(n12868), .ZN(n13223) );
  AOI21_X1 U7769 ( .B1(n13577), .B2(n6901), .A(n13182), .ZN(n6900) );
  INV_X1 U7770 ( .A(n13185), .ZN(n6901) );
  NAND2_X1 U7771 ( .A1(n12321), .A2(n13221), .ZN(n15789) );
  INV_X1 U7772 ( .A(n15211), .ZN(n15811) );
  CLKBUF_X1 U7773 ( .A(n8268), .Z(n10611) );
  AND2_X1 U7774 ( .A1(n13036), .A2(n7224), .ZN(n7223) );
  OR2_X1 U7775 ( .A1(n8325), .A2(n6833), .ZN(n7224) );
  NAND2_X1 U7776 ( .A1(n7829), .A2(n7828), .ZN(n8324) );
  NAND2_X1 U7777 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n14425), .ZN(n7828) );
  AND2_X1 U7778 ( .A1(n7783), .A2(n7785), .ZN(n6965) );
  INV_X1 U7779 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7785) );
  NAND2_X1 U7780 ( .A1(n7540), .A2(n6829), .ZN(n7206) );
  OR2_X1 U7781 ( .A1(n7538), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7205) );
  OAI21_X1 U7782 ( .B1(P2_DATAO_REG_17__SCAN_IN), .B2(n12066), .A(n7815), .ZN(
        n8117) );
  NAND2_X1 U7783 ( .A1(n7960), .A2(n7959), .ZN(n7801) );
  NAND2_X1 U7784 ( .A1(n7790), .A2(n7215), .ZN(n7214) );
  AND2_X1 U7785 ( .A1(n7792), .A2(n6700), .ZN(n7215) );
  NAND2_X1 U7786 ( .A1(n7541), .A2(n7794), .ZN(n7216) );
  OAI21_X1 U7787 ( .B1(n7903), .B2(n7543), .A(n7914), .ZN(n7541) );
  NAND2_X1 U7788 ( .A1(n12403), .A2(n12399), .ZN(n7451) );
  NOR2_X1 U7789 ( .A1(n10957), .A2(n9747), .ZN(n9684) );
  NAND2_X1 U7790 ( .A1(n6787), .A2(n7440), .ZN(n8384) );
  AND2_X1 U7791 ( .A1(n8415), .A2(n14412), .ZN(n8513) );
  NAND2_X1 U7792 ( .A1(n7009), .A2(n7008), .ZN(n14147) );
  NAND2_X1 U7793 ( .A1(n14363), .A2(n9668), .ZN(n14249) );
  NAND2_X1 U7794 ( .A1(n11648), .A2(n7517), .ZN(n7586) );
  NAND2_X1 U7795 ( .A1(n6916), .A2(n9647), .ZN(n10888) );
  NAND2_X1 U7796 ( .A1(n11842), .A2(n11841), .ZN(n6916) );
  NOR2_X1 U7797 ( .A1(n9748), .A2(n9747), .ZN(n15690) );
  NOR2_X1 U7798 ( .A1(n9759), .A2(n14424), .ZN(n15682) );
  NOR2_X1 U7799 ( .A1(n8836), .A2(n6924), .ZN(n6922) );
  INV_X1 U7800 ( .A(n8392), .ZN(n6923) );
  NAND2_X1 U7801 ( .A1(n6925), .A2(n8393), .ZN(n6924) );
  OAI211_X1 U7802 ( .C1(n11683), .C2(n11682), .A(n11681), .B(n11680), .ZN(
        n14507) );
  AOI22_X1 U7803 ( .A1(n11672), .A2(n11671), .B1(n11670), .B2(n11669), .ZN(
        n11681) );
  NAND2_X1 U7804 ( .A1(n15510), .A2(n10557), .ZN(n11438) );
  XNOR2_X1 U7806 ( .A(n14729), .B(n14549), .ZN(n14765) );
  NAND2_X1 U7807 ( .A1(n15026), .A2(n7366), .ZN(n14843) );
  AND2_X1 U7808 ( .A1(n14848), .A2(n14718), .ZN(n7366) );
  AOI21_X1 U7809 ( .B1(n14919), .B2(n14928), .A(n6761), .ZN(n14914) );
  AOI21_X1 U7810 ( .B1(n14961), .B2(n7686), .A(n6755), .ZN(n7685) );
  NOR2_X1 U7811 ( .A1(n12695), .A2(n7689), .ZN(n7686) );
  AOI21_X1 U7812 ( .B1(n12526), .B2(n7352), .A(n6760), .ZN(n7351) );
  NAND2_X1 U7813 ( .A1(n12024), .A2(n9797), .ZN(n12153) );
  OAI22_X1 U7814 ( .A1(n13331), .A2(n7273), .B1(n7274), .B2(n13354), .ZN(
        n13377) );
  OR2_X1 U7815 ( .A1(n13354), .A2(n13332), .ZN(n7273) );
  AND2_X1 U7816 ( .A1(n7157), .A2(n7160), .ZN(n6990) );
  INV_X1 U7817 ( .A(n13394), .ZN(n7160) );
  NAND2_X1 U7818 ( .A1(n7158), .A2(n12430), .ZN(n7157) );
  NAND2_X1 U7819 ( .A1(n14419), .A2(n6680), .ZN(n9082) );
  AND2_X1 U7820 ( .A1(n9744), .A2(n9743), .ZN(n14069) );
  XNOR2_X1 U7821 ( .A(n14089), .B(n14088), .ZN(n14300) );
  NAND2_X1 U7822 ( .A1(n10345), .A2(n10344), .ZN(n15014) );
  AND2_X1 U7823 ( .A1(n9989), .A2(n9988), .ZN(n9990) );
  AND2_X1 U7824 ( .A1(n8463), .A2(n8462), .ZN(n8495) );
  NAND2_X1 U7825 ( .A1(n13945), .A2(n6673), .ZN(n8463) );
  NAND2_X1 U7826 ( .A1(n13783), .A2(n8582), .ZN(n8462) );
  NAND2_X1 U7827 ( .A1(n8461), .A2(n8460), .ZN(n8498) );
  OAI21_X1 U7828 ( .B1(n7720), .B2(n7722), .A(n7721), .ZN(n8605) );
  NOR2_X1 U7829 ( .A1(n8585), .A2(n6744), .ZN(n7720) );
  NAND2_X1 U7830 ( .A1(n6714), .A2(n8557), .ZN(n7722) );
  NAND2_X1 U7831 ( .A1(n7734), .A2(n7733), .ZN(n7732) );
  INV_X1 U7832 ( .A(n6773), .ZN(n7734) );
  NAND2_X1 U7833 ( .A1(n7571), .A2(n10116), .ZN(n7570) );
  INV_X1 U7834 ( .A(n7101), .ZN(n7099) );
  AOI21_X1 U7835 ( .B1(n7101), .B2(n8729), .A(n6775), .ZN(n7100) );
  AND2_X1 U7836 ( .A1(n8707), .A2(n8708), .ZN(n7743) );
  NAND2_X1 U7837 ( .A1(n7098), .A2(n7096), .ZN(n7095) );
  INV_X1 U7838 ( .A(n7100), .ZN(n7096) );
  NAND2_X1 U7839 ( .A1(n7100), .A2(n7102), .ZN(n7093) );
  NAND2_X1 U7840 ( .A1(n7103), .A2(n8729), .ZN(n7102) );
  INV_X1 U7841 ( .A(n7743), .ZN(n7103) );
  INV_X1 U7842 ( .A(n7557), .ZN(n7556) );
  OAI211_X1 U7843 ( .C1(n7561), .C2(n7559), .A(n14918), .B(n7558), .ZN(n7557)
         );
  NAND2_X1 U7844 ( .A1(n14708), .A2(n7562), .ZN(n7558) );
  INV_X1 U7845 ( .A(n10255), .ZN(n7559) );
  NOR2_X1 U7846 ( .A1(n14708), .A2(n10255), .ZN(n7560) );
  INV_X1 U7847 ( .A(n13169), .ZN(n6853) );
  INV_X1 U7848 ( .A(n8779), .ZN(n7726) );
  NAND2_X1 U7849 ( .A1(n7741), .A2(n7091), .ZN(n7090) );
  NAND2_X1 U7850 ( .A1(n13196), .A2(n6861), .ZN(n6860) );
  NAND2_X1 U7851 ( .A1(n8877), .A2(n6756), .ZN(n7084) );
  NAND2_X1 U7852 ( .A1(n8973), .A2(n7081), .ZN(n7080) );
  INV_X1 U7853 ( .A(n8993), .ZN(n7731) );
  NAND2_X1 U7854 ( .A1(n13211), .A2(n13459), .ZN(n6984) );
  NAND2_X1 U7855 ( .A1(n13212), .A2(n13213), .ZN(n6983) );
  NAND2_X1 U7856 ( .A1(n10374), .A2(n7583), .ZN(n7582) );
  OAI21_X1 U7857 ( .B1(n7284), .B2(n7283), .A(n10703), .ZN(n7280) );
  NAND2_X1 U7858 ( .A1(n11146), .A2(n7281), .ZN(n7277) );
  INV_X1 U7859 ( .A(n13334), .ZN(n7156) );
  NOR2_X1 U7860 ( .A1(n7156), .A2(n13361), .ZN(n7155) );
  OR2_X1 U7861 ( .A1(n13550), .A2(n12897), .ZN(n13088) );
  INV_X1 U7862 ( .A(n8231), .ZN(n6942) );
  INV_X1 U7863 ( .A(n7814), .ZN(n7548) );
  NAND2_X1 U7864 ( .A1(n7611), .A2(n7606), .ZN(n7605) );
  INV_X1 U7865 ( .A(n9706), .ZN(n7606) );
  OAI21_X1 U7866 ( .B1(n6685), .B2(n7610), .A(n15280), .ZN(n7609) );
  INV_X1 U7867 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8365) );
  NOR2_X1 U7868 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n7066) );
  NOR2_X1 U7869 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n7068) );
  INV_X1 U7870 ( .A(n12053), .ZN(n7348) );
  NAND2_X1 U7871 ( .A1(n7671), .A2(n7670), .ZN(n7666) );
  NOR2_X1 U7872 ( .A1(n9099), .A2(n7669), .ZN(n7668) );
  INV_X1 U7873 ( .A(n7670), .ZN(n7669) );
  NAND2_X1 U7874 ( .A1(n7177), .A2(n7171), .ZN(n7170) );
  INV_X1 U7875 ( .A(n7182), .ZN(n7171) );
  AOI21_X1 U7876 ( .B1(n7194), .B2(n7196), .A(n7192), .ZN(n7191) );
  INV_X1 U7877 ( .A(n8731), .ZN(n7192) );
  NOR2_X1 U7878 ( .A1(n8712), .A2(n7198), .ZN(n7197) );
  INV_X1 U7879 ( .A(n8689), .ZN(n7198) );
  NAND2_X1 U7880 ( .A1(n9263), .A2(n9213), .ZN(n6872) );
  INV_X1 U7881 ( .A(n9855), .ZN(n7385) );
  NAND2_X1 U7882 ( .A1(n11260), .A2(n13098), .ZN(n9787) );
  OR2_X1 U7883 ( .A1(n10618), .A2(n11200), .ZN(n7425) );
  OR2_X1 U7884 ( .A1(n11289), .A2(n10599), .ZN(n7262) );
  OR2_X1 U7885 ( .A1(n13415), .A2(n9880), .ZN(n13225) );
  INV_X1 U7886 ( .A(n8251), .ZN(n6951) );
  INV_X1 U7887 ( .A(n6950), .ZN(n6949) );
  OAI21_X1 U7888 ( .B1(n13445), .B2(n6951), .A(n8252), .ZN(n6950) );
  OR2_X1 U7889 ( .A1(n8193), .A2(n7319), .ZN(n7318) );
  AND2_X1 U7890 ( .A1(n13218), .A2(n13215), .ZN(n13214) );
  XNOR2_X1 U7891 ( .A(n12951), .B(n13483), .ZN(n13459) );
  NAND2_X1 U7892 ( .A1(n13479), .A2(n8193), .ZN(n13458) );
  NAND2_X1 U7893 ( .A1(n13477), .A2(n13476), .ZN(n13479) );
  OR2_X1 U7894 ( .A1(n13499), .A2(n13507), .ZN(n13205) );
  AND2_X1 U7895 ( .A1(n13121), .A2(n13126), .ZN(n13124) );
  NAND2_X1 U7896 ( .A1(n13115), .A2(n13112), .ZN(n8215) );
  OAI21_X1 U7897 ( .B1(n8295), .B2(n8294), .A(n8293), .ZN(n8314) );
  INV_X1 U7898 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7783) );
  NAND2_X1 U7899 ( .A1(n7757), .A2(n7756), .ZN(n7778) );
  AND2_X1 U7900 ( .A1(n8103), .A2(n7777), .ZN(n7756) );
  NAND2_X1 U7901 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n12388), .ZN(n7817) );
  NOR2_X1 U7902 ( .A1(n9775), .A2(n14292), .ZN(n7472) );
  NOR2_X1 U7903 ( .A1(n6738), .A2(n14088), .ZN(n7512) );
  OR2_X1 U7904 ( .A1(n9677), .A2(n9728), .ZN(n7112) );
  NAND2_X1 U7905 ( .A1(n7476), .A2(n11994), .ZN(n6886) );
  INV_X1 U7906 ( .A(n9700), .ZN(n7587) );
  OAI21_X1 U7907 ( .B1(n7517), .B2(n7587), .A(n11806), .ZN(n7344) );
  INV_X1 U7908 ( .A(n9653), .ZN(n6934) );
  INV_X1 U7909 ( .A(n9746), .ZN(n14090) );
  INV_X1 U7910 ( .A(n14316), .ZN(n7464) );
  NOR2_X1 U7911 ( .A1(n7616), .A2(n7331), .ZN(n7330) );
  INV_X1 U7912 ( .A(n9723), .ZN(n7331) );
  INV_X1 U7913 ( .A(n7617), .ZN(n7616) );
  AOI21_X1 U7914 ( .B1(n7617), .B2(n7615), .A(n6764), .ZN(n7614) );
  INV_X1 U7915 ( .A(n9724), .ZN(n7615) );
  NOR2_X1 U7916 ( .A1(n14223), .A2(n14341), .ZN(n14204) );
  AND2_X1 U7917 ( .A1(n7314), .A2(n9719), .ZN(n7313) );
  NOR2_X1 U7918 ( .A1(n14269), .A2(n14364), .ZN(n14255) );
  NAND2_X1 U7919 ( .A1(n8884), .A2(n13964), .ZN(n7533) );
  AOI21_X1 U7920 ( .B1(n7479), .B2(n7481), .A(n6762), .ZN(n7477) );
  INV_X1 U7921 ( .A(n9904), .ZN(n7345) );
  NOR2_X1 U7922 ( .A1(n14794), .A2(n7356), .ZN(n7355) );
  INV_X1 U7923 ( .A(n14722), .ZN(n7356) );
  NAND2_X1 U7924 ( .A1(n12695), .A2(n14701), .ZN(n7361) );
  NAND2_X1 U7925 ( .A1(n14965), .A2(n7360), .ZN(n7362) );
  INV_X1 U7926 ( .A(n14701), .ZN(n7360) );
  OR2_X1 U7927 ( .A1(n15386), .A2(n15362), .ZN(n12693) );
  AND2_X1 U7928 ( .A1(n12615), .A2(n7678), .ZN(n7677) );
  OR2_X1 U7929 ( .A1(n12531), .A2(n7679), .ZN(n7678) );
  INV_X1 U7930 ( .A(n12532), .ZN(n7679) );
  NAND2_X1 U7931 ( .A1(n12251), .A2(n12250), .ZN(n12304) );
  OR2_X1 U7932 ( .A1(n11443), .A2(n11920), .ZN(n9953) );
  NAND2_X1 U7933 ( .A1(n7292), .A2(n15513), .ZN(n15502) );
  INV_X1 U7934 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9898) );
  INV_X1 U7935 ( .A(n9036), .ZN(n7651) );
  AND2_X1 U7936 ( .A1(n7261), .A2(n9921), .ZN(n7260) );
  INV_X1 U7937 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9889) );
  XNOR2_X1 U7938 ( .A(n8710), .B(SI_11_), .ZN(n8712) );
  AND2_X1 U7939 ( .A1(n8558), .A2(n8531), .ZN(n8532) );
  NAND2_X1 U7940 ( .A1(n6888), .A2(n6887), .ZN(n8404) );
  NAND2_X1 U7941 ( .A1(n8405), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6888) );
  OAI21_X1 U7942 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n9582), .A(n9228), .ZN(
        n9257) );
  NOR2_X1 U7943 ( .A1(n7389), .A2(n7385), .ZN(n7382) );
  OR2_X1 U7944 ( .A1(n9858), .A2(n9857), .ZN(n7389) );
  AOI21_X1 U7945 ( .B1(n7390), .B2(n9857), .A(n6770), .ZN(n7387) );
  OR2_X1 U7946 ( .A1(n13012), .A2(n9857), .ZN(n7388) );
  NAND2_X1 U7947 ( .A1(n7390), .A2(n7385), .ZN(n7384) );
  AND2_X1 U7948 ( .A1(n9858), .A2(n7391), .ZN(n7390) );
  OR2_X1 U7949 ( .A1(n13012), .A2(n9857), .ZN(n7391) );
  AND2_X1 U7950 ( .A1(n9855), .A2(n9853), .ZN(n12924) );
  NOR2_X1 U7951 ( .A1(n12453), .A2(n6958), .ZN(n6957) );
  INV_X1 U7952 ( .A(n9801), .ZN(n6958) );
  INV_X1 U7953 ( .A(n15209), .ZN(n12994) );
  INV_X1 U7954 ( .A(n9817), .ZN(n7397) );
  XNOR2_X1 U7955 ( .A(n11069), .B(P3_REG1_REG_2__SCAN_IN), .ZN(n11057) );
  NAND2_X1 U7956 ( .A1(n11051), .A2(n7145), .ZN(n7412) );
  NOR2_X1 U7957 ( .A1(n7146), .A2(n11030), .ZN(n7145) );
  INV_X1 U7958 ( .A(n10616), .ZN(n7146) );
  NAND2_X1 U7959 ( .A1(n7411), .A2(n7412), .ZN(n11142) );
  OAI21_X1 U7960 ( .B1(n7409), .B2(n7408), .A(n7407), .ZN(n7411) );
  NAND2_X1 U7961 ( .A1(n10648), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7407) );
  NAND2_X1 U7962 ( .A1(n10616), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7408) );
  AOI21_X1 U7963 ( .B1(n11051), .B2(n10616), .A(n10648), .ZN(n7410) );
  NAND2_X1 U7964 ( .A1(n7285), .A2(n7284), .ZN(n7282) );
  OR2_X1 U7965 ( .A1(n11025), .A2(n10646), .ZN(n11148) );
  NOR2_X1 U7966 ( .A1(n7425), .A2(n10619), .ZN(n11199) );
  NAND2_X1 U7967 ( .A1(n7424), .A2(n7425), .ZN(n7149) );
  XNOR2_X1 U7968 ( .A(n7262), .B(n10733), .ZN(n11314) );
  NOR2_X1 U7969 ( .A1(n11314), .A2(n10666), .ZN(n11313) );
  NAND2_X1 U7970 ( .A1(n7144), .A2(n6742), .ZN(n7405) );
  INV_X1 U7971 ( .A(n7406), .ZN(n10621) );
  OR2_X1 U7972 ( .A1(n11702), .A2(n10604), .ZN(n7430) );
  OR2_X1 U7973 ( .A1(n11699), .A2(n10626), .ZN(n10629) );
  AND2_X1 U7974 ( .A1(n12423), .A2(n12425), .ZN(n7415) );
  NAND2_X1 U7975 ( .A1(n7263), .A2(n6717), .ZN(n7428) );
  NOR2_X1 U7976 ( .A1(n13277), .A2(n13276), .ZN(n13278) );
  OR2_X1 U7977 ( .A1(n13278), .A2(n13283), .ZN(n7143) );
  AND2_X1 U7978 ( .A1(n7272), .A2(n6734), .ZN(n13322) );
  NAND2_X1 U7979 ( .A1(n13318), .A2(n13319), .ZN(n13320) );
  OR2_X1 U7980 ( .A1(n13322), .A2(n13321), .ZN(n13330) );
  NAND2_X1 U7981 ( .A1(n13364), .A2(n13363), .ZN(n13388) );
  OAI21_X1 U7982 ( .B1(n6721), .B2(n13226), .A(n13225), .ZN(n13056) );
  INV_X1 U7983 ( .A(n7626), .ZN(n7625) );
  NAND2_X1 U7984 ( .A1(n13446), .A2(n6949), .ZN(n6948) );
  AOI21_X1 U7985 ( .B1(n6949), .B2(n6951), .A(n6743), .ZN(n6947) );
  AOI21_X1 U7986 ( .B1(n6710), .B2(n7319), .A(n7316), .ZN(n7315) );
  INV_X1 U7987 ( .A(n13215), .ZN(n7316) );
  AND2_X1 U7988 ( .A1(n13216), .A2(n13219), .ZN(n13432) );
  NAND2_X1 U7989 ( .A1(n13479), .A2(n6710), .ZN(n7317) );
  AND2_X1 U7990 ( .A1(n7867), .A2(n7866), .ZN(n13448) );
  NAND2_X1 U7991 ( .A1(n8248), .A2(n7631), .ZN(n7630) );
  NOR2_X1 U7992 ( .A1(n6767), .A2(n7632), .ZN(n7631) );
  INV_X1 U7993 ( .A(n8247), .ZN(n7632) );
  INV_X1 U7994 ( .A(n7325), .ZN(n7324) );
  AOI21_X1 U7995 ( .B1(n7325), .B2(n7323), .A(n6766), .ZN(n7322) );
  INV_X1 U7996 ( .A(n13197), .ZN(n7323) );
  NAND2_X1 U7997 ( .A1(n13531), .A2(n8244), .ZN(n13517) );
  OAI21_X1 U7998 ( .B1(n13565), .B2(n7335), .A(n7333), .ZN(n13536) );
  INV_X1 U7999 ( .A(n7336), .ZN(n7335) );
  AOI21_X1 U8000 ( .B1(n7336), .B2(n13558), .A(n7334), .ZN(n7333) );
  NOR2_X1 U8001 ( .A1(n13094), .A2(n7337), .ZN(n7336) );
  NAND2_X1 U8002 ( .A1(n13542), .A2(n6956), .ZN(n13531) );
  AND2_X1 U8003 ( .A1(n13535), .A2(n8243), .ZN(n6956) );
  NAND2_X1 U8004 ( .A1(n13565), .A2(n13564), .ZN(n13563) );
  INV_X1 U8005 ( .A(n13176), .ZN(n12636) );
  AND2_X1 U8006 ( .A1(n6731), .A2(n8235), .ZN(n6944) );
  NAND2_X1 U8007 ( .A1(n15182), .A2(n8231), .ZN(n6945) );
  NAND2_X1 U8008 ( .A1(n15203), .A2(n15202), .ZN(n6910) );
  AND2_X1 U8009 ( .A1(n6792), .A2(n13166), .ZN(n15202) );
  NOR2_X1 U8010 ( .A1(n13066), .A2(n7639), .ZN(n7638) );
  INV_X1 U8011 ( .A(n8224), .ZN(n7639) );
  NAND2_X1 U8012 ( .A1(n12283), .A2(n8224), .ZN(n12119) );
  NAND2_X1 U8013 ( .A1(n12282), .A2(n6953), .ZN(n12281) );
  AND2_X1 U8014 ( .A1(n11961), .A2(n8223), .ZN(n12284) );
  NAND2_X1 U8015 ( .A1(n12284), .A2(n13144), .ZN(n12283) );
  OR2_X1 U8016 ( .A1(n13239), .A2(n8312), .ZN(n15211) );
  INV_X1 U8017 ( .A(n11260), .ZN(n15803) );
  INV_X1 U8018 ( .A(n15787), .ZN(n15809) );
  OR2_X1 U8019 ( .A1(n15161), .A2(n15160), .ZN(n15222) );
  NAND2_X1 U8020 ( .A1(n8327), .A2(n8326), .ZN(n13053) );
  NAND2_X1 U8021 ( .A1(n7842), .A2(n7841), .ZN(n13224) );
  NAND2_X1 U8022 ( .A1(n7859), .A2(n7858), .ZN(n13010) );
  OR2_X1 U8023 ( .A1(n12321), .A2(n13228), .ZN(n15787) );
  AND2_X1 U8024 ( .A1(n7332), .A2(n7640), .ZN(n7847) );
  OAI22_X1 U8025 ( .A1(n8324), .A2(n8323), .B1(P2_DATAO_REG_27__SCAN_IN), .B2(
        n9080), .ZN(n8336) );
  AOI21_X1 U8026 ( .B1(n8195), .B2(n7827), .A(n7826), .ZN(n7857) );
  AND2_X1 U8027 ( .A1(n15098), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7826) );
  NOR2_X1 U8028 ( .A1(P3_IR_REG_23__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), .ZN(
        n6969) );
  AOI21_X1 U8029 ( .B1(n7232), .B2(n7231), .A(n6831), .ZN(n8173) );
  INV_X1 U8030 ( .A(n8161), .ZN(n7231) );
  INV_X1 U8031 ( .A(n8162), .ZN(n7232) );
  NAND2_X1 U8032 ( .A1(n7554), .A2(n7821), .ZN(n8162) );
  NAND2_X1 U8033 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n12511), .ZN(n7821) );
  NAND2_X1 U8034 ( .A1(n8151), .A2(n8149), .ZN(n7554) );
  OAI21_X1 U8035 ( .B1(P2_DATAO_REG_18__SCAN_IN), .B2(n12317), .A(n7816), .ZN(
        n8131) );
  NAND2_X1 U8036 ( .A1(n7210), .A2(n7208), .ZN(n8101) );
  AOI21_X1 U8037 ( .B1(n7212), .B2(n7213), .A(n7209), .ZN(n7208) );
  AND2_X1 U8038 ( .A1(n7546), .A2(n6820), .ZN(n7212) );
  NAND2_X1 U8039 ( .A1(n7211), .A2(n7813), .ZN(n8070) );
  NAND2_X1 U8040 ( .A1(n8055), .A2(n7812), .ZN(n7211) );
  NAND2_X1 U8041 ( .A1(n7806), .A2(n7805), .ZN(n8021) );
  NAND2_X1 U8042 ( .A1(n7201), .A2(n7199), .ZN(n7806) );
  AOI21_X1 U8043 ( .B1(n7202), .B2(n7552), .A(n7200), .ZN(n7199) );
  INV_X1 U8044 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7802) );
  XNOR2_X1 U8045 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n7973) );
  NAND2_X1 U8046 ( .A1(n7801), .A2(n7800), .ZN(n7975) );
  OR2_X1 U8047 ( .A1(n7961), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n7976) );
  OAI21_X1 U8048 ( .B1(n7946), .B2(n7798), .A(n7799), .ZN(n7960) );
  XNOR2_X1 U8049 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n7930) );
  XNOR2_X1 U8050 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n7914) );
  INV_X1 U8051 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7791) );
  XNOR2_X1 U8052 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n7903) );
  NAND2_X1 U8053 ( .A1(n7790), .A2(n7789), .ZN(n7905) );
  NAND2_X1 U8054 ( .A1(n8010), .A2(n7434), .ZN(n7433) );
  NAND2_X1 U8055 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n7435) );
  OR3_X1 U8056 ( .A1(n14431), .A2(n14427), .A3(n14424), .ZN(n10507) );
  AOI21_X1 U8057 ( .B1(n7441), .B2(n7033), .A(n13762), .ZN(n7032) );
  NAND2_X1 U8058 ( .A1(n11177), .A2(n11115), .ZN(n13779) );
  NAND2_X1 U8059 ( .A1(n7506), .A2(n10717), .ZN(n7591) );
  INV_X1 U8060 ( .A(n7458), .ZN(n7040) );
  INV_X1 U8061 ( .A(n7039), .ZN(n7038) );
  OAI21_X1 U8062 ( .B1(n7041), .B2(n7040), .A(n13864), .ZN(n7039) );
  OR2_X1 U8063 ( .A1(n13875), .A2(n13750), .ZN(n7744) );
  OR2_X1 U8064 ( .A1(n7460), .A2(n7459), .ZN(n7458) );
  INV_X1 U8065 ( .A(n13741), .ZN(n7459) );
  AND2_X1 U8066 ( .A1(n7453), .A2(n12401), .ZN(n7452) );
  NAND2_X1 U8067 ( .A1(n12399), .A2(n7454), .ZN(n7453) );
  INV_X1 U8068 ( .A(n12184), .ZN(n7454) );
  NAND2_X1 U8069 ( .A1(n12183), .A2(n12182), .ZN(n12185) );
  INV_X1 U8070 ( .A(n7447), .ZN(n7033) );
  AND2_X1 U8071 ( .A1(n7444), .A2(n7442), .ZN(n7441) );
  AND2_X1 U8072 ( .A1(n6732), .A2(n13903), .ZN(n7444) );
  NAND2_X1 U8073 ( .A1(n7447), .A2(n13854), .ZN(n7442) );
  OAI21_X1 U8074 ( .B1(n6709), .B2(n7052), .A(n7049), .ZN(n7048) );
  AOI21_X1 U8075 ( .B1(n9161), .B2(n9160), .A(n9159), .ZN(n9172) );
  OR2_X1 U8076 ( .A1(n10870), .A2(n10869), .ZN(n12352) );
  OR2_X1 U8077 ( .A1(n7119), .A2(n14099), .ZN(n7118) );
  AOI21_X1 U8078 ( .B1(n7510), .B2(n7511), .A(n14072), .ZN(n7508) );
  NAND2_X1 U8079 ( .A1(n7329), .A2(n7327), .ZN(n14150) );
  NOR2_X1 U8080 ( .A1(n7008), .A2(n7328), .ZN(n7327) );
  INV_X1 U8081 ( .A(n7614), .ZN(n7328) );
  NAND2_X1 U8082 ( .A1(n7619), .A2(n9726), .ZN(n14167) );
  NAND2_X1 U8083 ( .A1(n14182), .A2(n9724), .ZN(n7619) );
  NOR2_X1 U8084 ( .A1(n14166), .A2(n7618), .ZN(n7617) );
  INV_X1 U8085 ( .A(n9726), .ZN(n7618) );
  INV_X1 U8086 ( .A(n9674), .ZN(n14166) );
  NAND2_X1 U8087 ( .A1(n14196), .A2(n9723), .ZN(n14182) );
  AOI21_X1 U8088 ( .B1(n7528), .B2(n14244), .A(n6763), .ZN(n7527) );
  NAND2_X1 U8089 ( .A1(n7467), .A2(n7466), .ZN(n14223) );
  AND2_X1 U8090 ( .A1(n14238), .A2(n9669), .ZN(n7528) );
  NAND2_X1 U8091 ( .A1(n14255), .A2(n14256), .ZN(n14258) );
  NAND2_X1 U8092 ( .A1(n14249), .A2(n7136), .ZN(n14250) );
  NAND2_X1 U8093 ( .A1(n7137), .A2(n7138), .ZN(n14245) );
  AOI21_X1 U8094 ( .B1(n6684), .B2(n7140), .A(n7139), .ZN(n7138) );
  NAND2_X1 U8095 ( .A1(n15254), .A2(n7132), .ZN(n7137) );
  NAND2_X1 U8096 ( .A1(n14245), .A2(n14244), .ZN(n14243) );
  AOI21_X1 U8097 ( .B1(n15254), .B2(n9712), .A(n6684), .ZN(n12487) );
  NAND2_X1 U8098 ( .A1(n9662), .A2(n9661), .ZN(n11893) );
  AOI21_X1 U8099 ( .B1(n11647), .B2(n7516), .A(n6722), .ZN(n7515) );
  NAND2_X1 U8100 ( .A1(n11527), .A2(n6939), .ZN(n7107) );
  NAND2_X1 U8101 ( .A1(n11092), .A2(n9652), .ZN(n6935) );
  NOR2_X1 U8102 ( .A1(n11590), .A2(n11125), .ZN(n7470) );
  NAND2_X1 U8103 ( .A1(n10888), .A2(n10889), .ZN(n6914) );
  NAND2_X1 U8104 ( .A1(n10890), .A2(n10887), .ZN(n9689) );
  INV_X1 U8105 ( .A(n10889), .ZN(n10887) );
  OAI21_X1 U8106 ( .B1(n9684), .B2(n6836), .A(n9162), .ZN(n15711) );
  INV_X1 U8107 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8410) );
  NOR2_X1 U8108 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n8398) );
  NAND2_X1 U8109 ( .A1(n6787), .A2(n7437), .ZN(n9194) );
  NOR2_X1 U8110 ( .A1(n8379), .A2(n6774), .ZN(n7437) );
  INV_X1 U8111 ( .A(n8388), .ZN(n7438) );
  OR2_X1 U8112 ( .A1(n8570), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n8615) );
  NAND2_X1 U8113 ( .A1(n11378), .A2(n11379), .ZN(n11683) );
  NAND2_X1 U8114 ( .A1(n7243), .A2(n12849), .ZN(n7236) );
  NAND2_X1 U8115 ( .A1(n7239), .A2(n10510), .ZN(n7241) );
  NAND2_X1 U8116 ( .A1(n7244), .A2(n7238), .ZN(n7237) );
  INV_X1 U8117 ( .A(n14750), .ZN(n14710) );
  AOI21_X1 U8118 ( .B1(n14436), .B2(n12836), .A(n12845), .ZN(n7491) );
  INV_X1 U8119 ( .A(n7491), .ZN(n7489) );
  NOR2_X1 U8120 ( .A1(n12236), .A2(n7494), .ZN(n7493) );
  INV_X1 U8121 ( .A(n12233), .ZN(n7494) );
  INV_X1 U8122 ( .A(n10520), .ZN(n10521) );
  NOR2_X1 U8123 ( .A1(n14465), .A2(n7497), .ZN(n7496) );
  NAND2_X1 U8124 ( .A1(n14514), .A2(n7250), .ZN(n7249) );
  INV_X1 U8125 ( .A(n12777), .ZN(n7497) );
  INV_X1 U8126 ( .A(n14525), .ZN(n7247) );
  INV_X1 U8127 ( .A(n14514), .ZN(n7251) );
  XNOR2_X1 U8128 ( .A(n10518), .B(n12672), .ZN(n10533) );
  NAND2_X1 U8129 ( .A1(n10517), .A2(n10516), .ZN(n10518) );
  OR2_X1 U8130 ( .A1(n12785), .A2(n11920), .ZN(n10516) );
  INV_X1 U8131 ( .A(n11691), .ZN(n7483) );
  OR2_X1 U8132 ( .A1(n10178), .A2(n10177), .ZN(n10193) );
  NAND2_X1 U8133 ( .A1(n10190), .A2(n10189), .ZN(n14700) );
  AOI211_X1 U8134 ( .C1(n10451), .C2(n10450), .A(n10449), .B(n10448), .ZN(
        n10456) );
  NAND2_X1 U8135 ( .A1(n10411), .A2(n10410), .ZN(n10445) );
  NOR2_X1 U8136 ( .A1(n7287), .A2(n14779), .ZN(n7286) );
  INV_X1 U8137 ( .A(n7288), .ZN(n7287) );
  INV_X1 U8138 ( .A(n7015), .ZN(n14796) );
  NAND2_X1 U8139 ( .A1(n14912), .A2(n7357), .ZN(n14888) );
  NOR2_X1 U8140 ( .A1(n14891), .A2(n7358), .ZN(n7357) );
  INV_X1 U8141 ( .A(n14711), .ZN(n7358) );
  NOR2_X1 U8142 ( .A1(n14928), .A2(n7698), .ZN(n7697) );
  INV_X1 U8143 ( .A(n14747), .ZN(n7698) );
  INV_X1 U8144 ( .A(n14918), .ZN(n14928) );
  AND2_X1 U8145 ( .A1(n10264), .A2(n14749), .ZN(n14918) );
  OR2_X1 U8146 ( .A1(n14949), .A2(n6733), .ZN(n6895) );
  NAND2_X1 U8147 ( .A1(n12696), .A2(n12695), .ZN(n14742) );
  NAND2_X1 U8148 ( .A1(n12529), .A2(n10465), .ZN(n12526) );
  NAND2_X1 U8149 ( .A1(n15503), .A2(n14814), .ZN(n11436) );
  INV_X1 U8150 ( .A(n14559), .ZN(n12006) );
  OAI21_X1 U8151 ( .B1(n15500), .B2(n15491), .A(n11913), .ZN(n12138) );
  AND2_X1 U8152 ( .A1(n11438), .A2(n10577), .ZN(n14735) );
  NAND2_X1 U8153 ( .A1(n7506), .A2(n9919), .ZN(n7505) );
  NAND2_X1 U8154 ( .A1(n10717), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7507) );
  NAND2_X1 U8155 ( .A1(n12672), .A2(n11440), .ZN(n15529) );
  XNOR2_X1 U8156 ( .A(n9103), .B(n9115), .ZN(n12705) );
  XNOR2_X1 U8157 ( .A(n9079), .B(n9078), .ZN(n14419) );
  NAND2_X1 U8158 ( .A1(n7167), .A2(n7175), .ZN(n7173) );
  INV_X1 U8159 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7567) );
  XNOR2_X1 U8160 ( .A(n8930), .B(n8929), .ZN(n12463) );
  NAND2_X1 U8161 ( .A1(n8665), .A2(n8664), .ZN(n8690) );
  INV_X1 U8162 ( .A(n7648), .ZN(n7647) );
  OAI21_X1 U8163 ( .B1(n8612), .B2(n7649), .A(n8636), .ZN(n7648) );
  INV_X1 U8164 ( .A(n8632), .ZN(n7649) );
  NAND2_X1 U8165 ( .A1(n8609), .A2(n8608), .ZN(n8613) );
  AND2_X1 U8166 ( .A1(n8472), .A2(n8473), .ZN(n10713) );
  NAND2_X1 U8167 ( .A1(n7662), .A2(n8444), .ZN(n8470) );
  INV_X1 U8168 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n7188) );
  INV_X1 U8169 ( .A(n9266), .ZN(n7305) );
  XNOR2_X1 U8170 ( .A(n9262), .B(n15475), .ZN(n9272) );
  NAND2_X1 U8171 ( .A1(n15131), .A2(n9292), .ZN(n6995) );
  OAI21_X1 U8172 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n15736), .A(n9233), .ZN(
        n9253) );
  OAI22_X1 U8173 ( .A1(n9238), .A2(P1_ADDR_REG_13__SCAN_IN), .B1(n9298), .B2(
        n9237), .ZN(n9250) );
  INV_X1 U8174 ( .A(n13659), .ZN(n12713) );
  NAND2_X1 U8175 ( .A1(n8153), .A2(n8152), .ZN(n13086) );
  AND3_X1 U8176 ( .A1(n8160), .A2(n8159), .A3(n8158), .ZN(n13496) );
  INV_X1 U8177 ( .A(n13018), .ZN(n7012) );
  NAND2_X1 U8178 ( .A1(n9863), .A2(n11465), .ZN(n13035) );
  AND2_X1 U8179 ( .A1(n9861), .A2(n9860), .ZN(n13023) );
  NAND2_X1 U8180 ( .A1(n6842), .A2(n13239), .ZN(n6850) );
  NAND2_X1 U8181 ( .A1(n13235), .A2(n15798), .ZN(n6846) );
  INV_X1 U8182 ( .A(n6848), .ZN(n6847) );
  AND2_X1 U8183 ( .A1(n11723), .A2(n8333), .ZN(n13411) );
  NAND2_X1 U8184 ( .A1(n7855), .A2(n7854), .ZN(n12868) );
  NAND2_X1 U8185 ( .A1(n8182), .A2(n8181), .ZN(n13466) );
  XNOR2_X1 U8186 ( .A(n7406), .B(n10733), .ZN(n11306) );
  NOR2_X1 U8187 ( .A1(n13377), .A2(n13376), .ZN(n13379) );
  OR2_X1 U8188 ( .A1(n10688), .A2(n6672), .ZN(n15744) );
  NAND2_X1 U8189 ( .A1(n13046), .A2(n13045), .ZN(n13057) );
  OAI21_X1 U8190 ( .B1(n8354), .B2(n15811), .A(n8353), .ZN(n13398) );
  INV_X1 U8191 ( .A(n11475), .ZN(n11467) );
  NAND2_X1 U8192 ( .A1(n15854), .A2(n15796), .ZN(n13626) );
  INV_X1 U8193 ( .A(n13053), .ZN(n13400) );
  NOR2_X1 U8194 ( .A1(n13398), .A2(n8355), .ZN(n8364) );
  AND2_X1 U8195 ( .A1(n15241), .A2(n13402), .ZN(n8355) );
  INV_X1 U8196 ( .A(n13010), .ZN(n13647) );
  NAND2_X1 U8197 ( .A1(n8092), .A2(n8091), .ZN(n13681) );
  OAI211_X1 U8198 ( .C1(n13044), .C2(SI_9_), .A(n7999), .B(n7998), .ZN(n13147)
         );
  AND3_X1 U8199 ( .A1(n7951), .A2(n7950), .A3(n7949), .ZN(n12030) );
  NAND2_X1 U8200 ( .A1(n15846), .A2(n15796), .ZN(n13676) );
  INV_X1 U8201 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7831) );
  AND2_X1 U8202 ( .A1(n7786), .A2(n8272), .ZN(n13243) );
  INV_X1 U8203 ( .A(n7401), .ZN(n7400) );
  XNOR2_X1 U8204 ( .A(n13752), .B(n6811), .ZN(n13770) );
  AND2_X1 U8205 ( .A1(n13789), .A2(n13737), .ZN(n7460) );
  NAND2_X1 U8206 ( .A1(n7461), .A2(n13736), .ZN(n13893) );
  INV_X1 U8207 ( .A(n13892), .ZN(n7461) );
  NAND2_X1 U8208 ( .A1(n10966), .A2(n15676), .ZN(n13914) );
  OR2_X1 U8209 ( .A1(n9130), .A2(n11591), .ZN(n8547) );
  NAND2_X1 U8210 ( .A1(n8542), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8418) );
  NAND2_X1 U8211 ( .A1(n9025), .A2(n9024), .ZN(n14310) );
  AND2_X1 U8212 ( .A1(n9677), .A2(n9676), .ZN(n7534) );
  NOR2_X1 U8213 ( .A1(n14274), .A2(n7530), .ZN(n7529) );
  INV_X1 U8214 ( .A(n9667), .ZN(n7530) );
  NAND2_X1 U8215 ( .A1(n14067), .A2(n15722), .ZN(n7190) );
  NAND2_X1 U8216 ( .A1(n14300), .A2(n15722), .ZN(n6919) );
  INV_X1 U8217 ( .A(n14299), .ZN(n6921) );
  NAND2_X1 U8218 ( .A1(n9767), .A2(n9766), .ZN(n15685) );
  NAND2_X1 U8219 ( .A1(n11610), .A2(n11612), .ZN(n11611) );
  AND4_X1 U8220 ( .A1(n10199), .A2(n10198), .A3(n10197), .A4(n10196), .ZN(
        n15326) );
  NAND2_X1 U8221 ( .A1(n10163), .A2(n10162), .ZN(n15342) );
  INV_X1 U8222 ( .A(n15513), .ZN(n11936) );
  AOI21_X1 U8223 ( .B1(n12860), .B2(n10423), .A(n9920), .ZN(n14989) );
  AOI21_X1 U8224 ( .B1(n14770), .B2(n7713), .A(n6779), .ZN(n7712) );
  AND2_X1 U8225 ( .A1(n14838), .A2(n14719), .ZN(n7365) );
  NAND2_X1 U8226 ( .A1(n10219), .A2(n10218), .ZN(n15371) );
  INV_X1 U8227 ( .A(n14973), .ZN(n14814) );
  NAND2_X1 U8228 ( .A1(n10080), .A2(n10079), .ZN(n12302) );
  INV_X1 U8229 ( .A(n15505), .ZN(n14873) );
  NAND2_X1 U8230 ( .A1(n15133), .A2(n15132), .ZN(n15131) );
  NOR2_X1 U8231 ( .A1(n15424), .A2(n15425), .ZN(n15423) );
  OAI21_X1 U8232 ( .B1(n15437), .B2(n15436), .A(n7301), .ZN(n6877) );
  INV_X1 U8233 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7301) );
  NAND2_X1 U8234 ( .A1(n15111), .A2(n15110), .ZN(n15109) );
  OAI21_X1 U8235 ( .B1(n15111), .B2(n15110), .A(n7310), .ZN(n7309) );
  INV_X1 U8236 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n7310) );
  AND2_X1 U8237 ( .A1(n8487), .A2(n8486), .ZN(n8488) );
  NAND2_X1 U8238 ( .A1(n8436), .A2(n8435), .ZN(n8490) );
  NAND2_X1 U8239 ( .A1(n8433), .A2(n15691), .ZN(n8436) );
  NAND2_X1 U8240 ( .A1(n13947), .A2(n7746), .ZN(n8435) );
  NAND2_X1 U8241 ( .A1(n8498), .A2(n8495), .ZN(n8489) );
  INV_X1 U8242 ( .A(n8495), .ZN(n8496) );
  NAND2_X1 U8243 ( .A1(n10048), .A2(n10050), .ZN(n7566) );
  OR2_X1 U8244 ( .A1(n7580), .A2(n10082), .ZN(n7579) );
  INV_X1 U8245 ( .A(n10081), .ZN(n7580) );
  NAND2_X1 U8246 ( .A1(n9114), .A2(n13942), .ZN(n7063) );
  INV_X1 U8247 ( .A(n8631), .ZN(n7733) );
  NAND2_X1 U8248 ( .A1(n6773), .A2(n8631), .ZN(n7735) );
  OAI21_X1 U8249 ( .B1(n8605), .B2(n7071), .A(n6711), .ZN(n7069) );
  NOR2_X1 U8250 ( .A1(n8607), .A2(n6790), .ZN(n7071) );
  NOR2_X1 U8251 ( .A1(n8708), .A2(n8707), .ZN(n7101) );
  NAND2_X1 U8252 ( .A1(n10149), .A2(n10151), .ZN(n7564) );
  NOR2_X1 U8253 ( .A1(n14707), .A2(n7562), .ZN(n7561) );
  NAND2_X1 U8254 ( .A1(n7097), .A2(n7743), .ZN(n7094) );
  NAND2_X1 U8255 ( .A1(n7556), .A2(n7560), .ZN(n6987) );
  NAND2_X1 U8256 ( .A1(n6852), .A2(n13168), .ZN(n6851) );
  INV_X1 U8257 ( .A(n8801), .ZN(n7076) );
  NOR2_X1 U8258 ( .A1(n8801), .A2(n8804), .ZN(n7077) );
  NAND2_X1 U8259 ( .A1(n7728), .A2(n7725), .ZN(n8802) );
  NAND2_X1 U8260 ( .A1(n7727), .A2(n7726), .ZN(n7725) );
  INV_X1 U8261 ( .A(n8780), .ZN(n7727) );
  NOR2_X1 U8262 ( .A1(n6719), .A2(n7074), .ZN(n7073) );
  INV_X1 U8263 ( .A(n8826), .ZN(n7074) );
  INV_X1 U8264 ( .A(n7077), .ZN(n7075) );
  NAND2_X1 U8265 ( .A1(n7741), .A2(n7089), .ZN(n7088) );
  INV_X1 U8266 ( .A(n8875), .ZN(n7089) );
  NAND2_X1 U8267 ( .A1(n7574), .A2(n10318), .ZN(n7573) );
  OAI21_X1 U8268 ( .B1(n10306), .B2(n10305), .A(n6772), .ZN(n7572) );
  NAND2_X1 U8269 ( .A1(n13199), .A2(n13200), .ZN(n6858) );
  NAND2_X1 U8270 ( .A1(n7084), .A2(n6746), .ZN(n8924) );
  NAND2_X1 U8271 ( .A1(n7577), .A2(n10346), .ZN(n7576) );
  OR2_X1 U8272 ( .A1(n9928), .A2(n12393), .ZN(n9929) );
  AND2_X1 U8273 ( .A1(n13432), .A2(n13215), .ZN(n6863) );
  NAND2_X1 U8274 ( .A1(n13216), .A2(n13228), .ZN(n6862) );
  NAND2_X1 U8275 ( .A1(n7079), .A2(n7078), .ZN(n9013) );
  AOI21_X1 U8276 ( .B1(n6689), .B2(n7082), .A(n6784), .ZN(n7078) );
  AND2_X1 U8277 ( .A1(n8972), .A2(n8975), .ZN(n7082) );
  NAND2_X1 U8278 ( .A1(n7322), .A2(n7324), .ZN(n6904) );
  NAND2_X1 U8279 ( .A1(n11178), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7221) );
  NAND2_X1 U8280 ( .A1(n7220), .A2(n7221), .ZN(n7219) );
  INV_X1 U8281 ( .A(n7807), .ZN(n7220) );
  AOI21_X1 U8282 ( .B1(n9735), .B2(n7597), .A(n7596), .ZN(n7595) );
  INV_X1 U8283 ( .A(n14088), .ZN(n7597) );
  INV_X1 U8284 ( .A(n9736), .ZN(n7596) );
  NAND2_X1 U8285 ( .A1(n7142), .A2(n7599), .ZN(n7133) );
  OR2_X1 U8286 ( .A1(n6716), .A2(n9718), .ZN(n7314) );
  AND2_X1 U8287 ( .A1(n7479), .A2(n7254), .ZN(n7253) );
  NAND2_X1 U8288 ( .A1(n12681), .A2(n7255), .ZN(n7254) );
  NOR2_X1 U8289 ( .A1(n15347), .A2(n7750), .ZN(n7255) );
  INV_X1 U8290 ( .A(n7257), .ZN(n7256) );
  AND2_X1 U8291 ( .A1(n7480), .A2(n15303), .ZN(n7479) );
  OR2_X1 U8292 ( .A1(n12726), .A2(n7481), .ZN(n7480) );
  INV_X1 U8293 ( .A(n12731), .ZN(n7481) );
  INV_X1 U8294 ( .A(n9951), .ZN(n10025) );
  AND2_X1 U8295 ( .A1(n9018), .A2(n7655), .ZN(n7654) );
  INV_X1 U8296 ( .A(n9037), .ZN(n7655) );
  NOR2_X1 U8297 ( .A1(n9037), .A2(n9016), .ZN(n7652) );
  AND2_X1 U8298 ( .A1(n6823), .A2(n8906), .ZN(n7182) );
  NAND2_X1 U8299 ( .A1(n8783), .A2(n10864), .ZN(n8807) );
  OAI21_X1 U8300 ( .B1(n8405), .B2(n6986), .A(n6985), .ZN(n8442) );
  NAND2_X1 U8301 ( .A1(n8405), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6985) );
  NAND2_X1 U8302 ( .A1(n6880), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n7840) );
  NAND2_X1 U8303 ( .A1(n6881), .A2(n7838), .ZN(n7839) );
  INV_X1 U8304 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7838) );
  INV_X1 U8305 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n9407) );
  INV_X1 U8306 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n9517) );
  INV_X1 U8307 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7772) );
  AOI21_X1 U8308 ( .B1(n13230), .B2(n7535), .A(n13229), .ZN(n6868) );
  OR2_X1 U8309 ( .A1(n13224), .A2(n13434), .ZN(n7535) );
  INV_X1 U8310 ( .A(n13232), .ZN(n6981) );
  OAI21_X1 U8311 ( .B1(n6725), .B2(n13058), .A(n13233), .ZN(n6976) );
  INV_X1 U8312 ( .A(n11051), .ZN(n7409) );
  OAI21_X1 U8313 ( .B1(n7278), .B2(n11025), .A(n7276), .ZN(n10597) );
  NAND2_X1 U8314 ( .A1(n7279), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7278) );
  NAND2_X1 U8315 ( .A1(n7279), .A2(n7277), .ZN(n7276) );
  AND2_X1 U8316 ( .A1(n11403), .A2(n10602), .ZN(n10603) );
  AOI21_X1 U8317 ( .B1(n13303), .B2(n7155), .A(n6834), .ZN(n7152) );
  OR2_X1 U8318 ( .A1(n13302), .A2(n7153), .ZN(n7151) );
  NAND2_X1 U8319 ( .A1(n13361), .A2(n7154), .ZN(n7153) );
  NOR2_X1 U8320 ( .A1(n13223), .A2(n6743), .ZN(n7627) );
  OR2_X1 U8321 ( .A1(n13446), .A2(n6951), .ZN(n6946) );
  NOR2_X1 U8322 ( .A1(n6735), .A2(n7623), .ZN(n7622) );
  INV_X1 U8323 ( .A(n8252), .ZN(n7623) );
  OAI21_X1 U8324 ( .B1(n7627), .B2(n6735), .A(n13407), .ZN(n7626) );
  NOR2_X1 U8325 ( .A1(n8199), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8198) );
  OR2_X1 U8326 ( .A1(n8176), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8186) );
  AND2_X1 U8327 ( .A1(n8155), .A2(n8154), .ZN(n8165) );
  INV_X1 U8328 ( .A(n13093), .ZN(n7337) );
  INV_X1 U8329 ( .A(n13088), .ZN(n7334) );
  OAI21_X1 U8330 ( .B1(n15182), .B2(n6943), .A(n6941), .ZN(n7636) );
  INV_X1 U8331 ( .A(n6944), .ZN(n6943) );
  AOI21_X1 U8332 ( .B1(n6944), .B2(n6942), .A(n6781), .ZN(n6941) );
  INV_X1 U8333 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n12431) );
  INV_X1 U8334 ( .A(n8284), .ZN(n8293) );
  NAND2_X1 U8335 ( .A1(n6971), .A2(n11788), .ZN(n13238) );
  INV_X1 U8336 ( .A(n13243), .ZN(n8258) );
  INV_X1 U8337 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n6899) );
  NAND2_X1 U8338 ( .A1(n7540), .A2(n7817), .ZN(n7819) );
  NAND2_X1 U8339 ( .A1(n7403), .A2(n8103), .ZN(n7402) );
  INV_X1 U8340 ( .A(n7813), .ZN(n7213) );
  INV_X1 U8341 ( .A(n7544), .ZN(n7209) );
  AOI21_X1 U8342 ( .B1(n7546), .B2(n7548), .A(n6817), .ZN(n7544) );
  INV_X1 U8343 ( .A(n8007), .ZN(n7200) );
  INV_X1 U8344 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7804) );
  INV_X1 U8345 ( .A(n7803), .ZN(n7553) );
  AND2_X1 U8346 ( .A1(n8816), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8843) );
  AND2_X1 U8347 ( .A1(n9026), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n9041) );
  INV_X1 U8348 ( .A(n7451), .ZN(n7050) );
  INV_X1 U8349 ( .A(n9733), .ZN(n7123) );
  AND2_X1 U8350 ( .A1(n9738), .A2(n9734), .ZN(n7116) );
  INV_X1 U8351 ( .A(n7595), .ZN(n7125) );
  INV_X1 U8352 ( .A(n7609), .ZN(n7608) );
  NOR2_X1 U8353 ( .A1(n8719), .A2(n8718), .ZN(n8743) );
  NOR2_X1 U8354 ( .A1(n12191), .A2(n6886), .ZN(n7474) );
  NOR2_X1 U8355 ( .A1(n8645), .A2(n8644), .ZN(n8669) );
  NOR2_X1 U8356 ( .A1(n7517), .A2(n6939), .ZN(n6938) );
  INV_X1 U8357 ( .A(n9658), .ZN(n7516) );
  NAND2_X1 U8358 ( .A1(n9698), .A2(n9697), .ZN(n11527) );
  AND2_X1 U8359 ( .A1(n7068), .A2(n7066), .ZN(n7065) );
  AND2_X1 U8360 ( .A1(n8365), .A2(n8366), .ZN(n7064) );
  INV_X1 U8361 ( .A(n10510), .ZN(n7240) );
  AND2_X1 U8362 ( .A1(n12672), .A2(n14561), .ZN(n7243) );
  AND2_X1 U8363 ( .A1(n11676), .A2(n11675), .ZN(n11677) );
  INV_X1 U8364 ( .A(n12773), .ZN(n7250) );
  AND2_X1 U8365 ( .A1(n10436), .A2(n10437), .ZN(n10442) );
  INV_X1 U8366 ( .A(n14756), .ZN(n7704) );
  INV_X1 U8367 ( .A(n14847), .ZN(n7703) );
  NOR2_X1 U8368 ( .A1(n7705), .A2(n7701), .ZN(n7700) );
  INV_X1 U8369 ( .A(n7707), .ZN(n7701) );
  NOR2_X1 U8370 ( .A1(n14878), .A2(n7708), .ZN(n7707) );
  INV_X1 U8371 ( .A(n14753), .ZN(n7708) );
  AND2_X1 U8372 ( .A1(n7300), .A2(n14884), .ZN(n7299) );
  NOR2_X1 U8373 ( .A1(n15041), .A2(n15046), .ZN(n7300) );
  NOR2_X1 U8374 ( .A1(n12697), .A2(n14700), .ZN(n14687) );
  INV_X1 U8375 ( .A(n12468), .ZN(n7352) );
  AND3_X1 U8376 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n10038) );
  NOR2_X1 U8377 ( .A1(n14563), .A2(n11506), .ZN(n11912) );
  NAND2_X1 U8378 ( .A1(n6890), .A2(n14715), .ZN(n14865) );
  AND2_X1 U8379 ( .A1(n7347), .A2(n12244), .ZN(n7346) );
  NAND2_X1 U8380 ( .A1(n7667), .A2(n7664), .ZN(n9126) );
  INV_X1 U8381 ( .A(n7665), .ZN(n7664) );
  OAI21_X1 U8382 ( .B1(n9099), .B2(n7666), .A(n9098), .ZN(n7665) );
  NAND2_X1 U8383 ( .A1(n9898), .A2(n7718), .ZN(n7717) );
  INV_X1 U8384 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7718) );
  NAND2_X1 U8385 ( .A1(n9017), .A2(SI_24_), .ZN(n9018) );
  OR2_X1 U8386 ( .A1(n8958), .A2(n7180), .ZN(n7179) );
  NAND2_X1 U8387 ( .A1(n8907), .A2(n7172), .ZN(n7175) );
  AND2_X1 U8388 ( .A1(n7182), .A2(SI_22_), .ZN(n7172) );
  NAND2_X1 U8389 ( .A1(n8860), .A2(n8859), .ZN(n8900) );
  XNOR2_X1 U8390 ( .A(n8733), .B(n10742), .ZN(n8731) );
  AOI21_X1 U8391 ( .B1(n7195), .B2(n7197), .A(n6780), .ZN(n7194) );
  INV_X1 U8392 ( .A(n7197), .ZN(n7196) );
  OR2_X1 U8393 ( .A1(n10051), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n10077) );
  NOR2_X1 U8394 ( .A1(n7184), .A2(n7185), .ZN(n6885) );
  INV_X1 U8395 ( .A(n8527), .ZN(n7184) );
  NAND2_X1 U8396 ( .A1(n6896), .A2(n8444), .ZN(n8473) );
  INV_X1 U8397 ( .A(n7661), .ZN(n6896) );
  NAND2_X1 U8398 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n9208), .ZN(n9209) );
  INV_X1 U8399 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n9211) );
  OAI21_X1 U8400 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n9222), .A(n9221), .ZN(
        n9223) );
  OAI21_X1 U8401 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n9565), .A(n9227), .ZN(
        n9259) );
  INV_X1 U8402 ( .A(n9790), .ZN(n7378) );
  INV_X1 U8403 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n11407) );
  NOR2_X1 U8404 ( .A1(n9848), .A2(n6964), .ZN(n6963) );
  INV_X1 U8405 ( .A(n9845), .ZN(n6964) );
  NAND2_X1 U8406 ( .A1(n7987), .A2(n7986), .ZN(n8001) );
  NOR2_X1 U8407 ( .A1(n12893), .A2(n6962), .ZN(n6961) );
  INV_X1 U8408 ( .A(n9829), .ZN(n6962) );
  NAND2_X1 U8409 ( .A1(n7399), .A2(n7398), .ZN(n12911) );
  INV_X1 U8410 ( .A(n12913), .ZN(n7398) );
  INV_X1 U8411 ( .A(n12910), .ZN(n7399) );
  NOR2_X1 U8412 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), .ZN(
        n6839) );
  NOR2_X1 U8413 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n6838) );
  NAND2_X1 U8414 ( .A1(n7147), .A2(n10620), .ZN(n7406) );
  OR2_X1 U8415 ( .A1(n11313), .A2(n10601), .ZN(n7419) );
  INV_X1 U8416 ( .A(n7262), .ZN(n10600) );
  NAND2_X1 U8417 ( .A1(n11411), .A2(n10622), .ZN(n10624) );
  XNOR2_X1 U8418 ( .A(n10603), .B(n10677), .ZN(n11703) );
  NOR2_X1 U8419 ( .A1(n15733), .A2(n12427), .ZN(n13258) );
  NAND2_X1 U8420 ( .A1(n13247), .A2(n13246), .ZN(n6988) );
  OR2_X1 U8421 ( .A1(n13248), .A2(n8048), .ZN(n7264) );
  XNOR2_X1 U8422 ( .A(n13259), .B(n15124), .ZN(n13260) );
  OR2_X1 U8423 ( .A1(n13318), .A2(n13308), .ZN(n7267) );
  NAND2_X1 U8424 ( .A1(n13318), .A2(n6835), .ZN(n7271) );
  INV_X1 U8425 ( .A(n13319), .ZN(n7270) );
  NAND2_X1 U8426 ( .A1(n7143), .A2(n13304), .ZN(n13299) );
  INV_X1 U8427 ( .A(n7421), .ZN(n13360) );
  NAND2_X1 U8428 ( .A1(n13330), .A2(n13329), .ZN(n13353) );
  AOI21_X1 U8429 ( .B1(n13356), .B2(n13361), .A(n13355), .ZN(n13383) );
  XNOR2_X1 U8430 ( .A(n13390), .B(n7159), .ZN(n7158) );
  INV_X1 U8431 ( .A(n13389), .ZN(n7159) );
  OR2_X1 U8432 ( .A1(n8262), .A2(n15162), .ZN(n13416) );
  INV_X1 U8433 ( .A(n6906), .ZN(n6905) );
  OAI21_X1 U8434 ( .B1(n7315), .B2(n6907), .A(n13219), .ZN(n6906) );
  INV_X1 U8435 ( .A(n13216), .ZN(n6907) );
  NAND2_X1 U8436 ( .A1(n13444), .A2(n8251), .ZN(n13430) );
  AND2_X1 U8437 ( .A1(n8206), .A2(n8205), .ZN(n13433) );
  NAND2_X1 U8438 ( .A1(n13446), .A2(n13445), .ZN(n13444) );
  NAND2_X1 U8439 ( .A1(n13458), .A2(n13083), .ZN(n13443) );
  NAND2_X1 U8440 ( .A1(n13480), .A2(n8249), .ZN(n13465) );
  NAND2_X1 U8441 ( .A1(n13465), .A2(n13464), .ZN(n13463) );
  NAND2_X1 U8442 ( .A1(n7630), .A2(n7629), .ZN(n13480) );
  AND2_X1 U8443 ( .A1(n13481), .A2(n6718), .ZN(n7629) );
  NAND2_X1 U8444 ( .A1(n13460), .A2(n13207), .ZN(n13481) );
  OR2_X1 U8445 ( .A1(n8135), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8144) );
  NAND2_X1 U8446 ( .A1(n7326), .A2(n13196), .ZN(n13523) );
  NAND2_X1 U8447 ( .A1(n7620), .A2(n13094), .ZN(n13542) );
  AND2_X1 U8448 ( .A1(n8109), .A2(n12944), .ZN(n8123) );
  INV_X1 U8449 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n12944) );
  NAND2_X1 U8450 ( .A1(n13557), .A2(n13558), .ZN(n13556) );
  NAND2_X1 U8451 ( .A1(n7636), .A2(n8238), .ZN(n13571) );
  NAND2_X1 U8452 ( .A1(n7636), .A2(n7634), .ZN(n13573) );
  NOR2_X1 U8453 ( .A1(n13577), .A2(n7635), .ZN(n7634) );
  INV_X1 U8454 ( .A(n8238), .ZN(n7635) );
  NAND2_X1 U8455 ( .A1(n8063), .A2(n12883), .ZN(n8077) );
  NAND2_X1 U8456 ( .A1(n6840), .A2(n13170), .ZN(n15177) );
  NAND2_X1 U8457 ( .A1(n6910), .A2(n6908), .ZN(n6840) );
  NOR2_X1 U8458 ( .A1(n8053), .A2(n6909), .ZN(n6908) );
  INV_X1 U8459 ( .A(n13166), .ZN(n6909) );
  NOR2_X1 U8460 ( .A1(n8047), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8063) );
  OAI21_X1 U8461 ( .B1(n12284), .B2(n6954), .A(n6952), .ZN(n12320) );
  INV_X1 U8462 ( .A(n7638), .ZN(n6954) );
  AOI21_X1 U8463 ( .B1(n7638), .B2(n6953), .A(n6726), .ZN(n6952) );
  NAND2_X1 U8464 ( .A1(n12320), .A2(n13151), .ZN(n12319) );
  AND2_X1 U8465 ( .A1(n8268), .A2(n10632), .ZN(n12321) );
  NAND2_X1 U8466 ( .A1(n11778), .A2(n8220), .ZN(n11625) );
  NAND2_X1 U8467 ( .A1(n7633), .A2(n11778), .ZN(n11627) );
  AND2_X1 U8468 ( .A1(n8221), .A2(n8220), .ZN(n7633) );
  NAND2_X1 U8469 ( .A1(n6837), .A2(n13121), .ZN(n11631) );
  AND2_X1 U8470 ( .A1(n13127), .A2(n13133), .ZN(n13062) );
  NAND2_X1 U8471 ( .A1(n11540), .A2(n6955), .ZN(n11778) );
  AND2_X1 U8472 ( .A1(n11779), .A2(n8218), .ZN(n6955) );
  AND2_X1 U8473 ( .A1(n11540), .A2(n8218), .ZN(n11780) );
  NAND2_X1 U8474 ( .A1(n11537), .A2(n13123), .ZN(n11777) );
  AND2_X1 U8475 ( .A1(n8215), .A2(n11424), .ZN(n6974) );
  NOR2_X1 U8476 ( .A1(n10608), .A2(n15815), .ZN(n11465) );
  NAND2_X1 U8477 ( .A1(n8213), .A2(n8212), .ZN(n15783) );
  INV_X1 U8478 ( .A(n13393), .ZN(n13081) );
  NAND2_X1 U8479 ( .A1(n11464), .A2(n11463), .ZN(n11466) );
  NAND2_X1 U8480 ( .A1(n8197), .A2(n8196), .ZN(n12920) );
  NAND2_X1 U8481 ( .A1(n8185), .A2(n8184), .ZN(n12951) );
  NAND2_X1 U8482 ( .A1(n12495), .A2(n6676), .ZN(n8185) );
  INV_X1 U8483 ( .A(n15831), .ZN(n15842) );
  INV_X1 U8484 ( .A(n15815), .ZN(n15796) );
  OR2_X1 U8485 ( .A1(n8316), .A2(n8315), .ZN(n9876) );
  NOR2_X1 U8486 ( .A1(n7226), .A2(n7228), .ZN(n7225) );
  INV_X1 U8487 ( .A(n13047), .ZN(n7226) );
  NAND2_X1 U8488 ( .A1(n7825), .A2(n7824), .ZN(n8195) );
  XNOR2_X1 U8489 ( .A(n7823), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n8183) );
  INV_X1 U8490 ( .A(n7817), .ZN(n7539) );
  NAND2_X1 U8491 ( .A1(n8131), .A2(n8129), .ZN(n7540) );
  NOR2_X1 U8492 ( .A1(n7402), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n7401) );
  NAND2_X1 U8493 ( .A1(n7641), .A2(n7403), .ZN(n8102) );
  NAND2_X1 U8494 ( .A1(n7811), .A2(n7810), .ZN(n8055) );
  OR2_X1 U8495 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n7809), .ZN(n7810) );
  XNOR2_X1 U8496 ( .A(n7809), .B(n11258), .ZN(n8042) );
  OR2_X1 U8497 ( .A1(n8028), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n8029) );
  AND2_X1 U8498 ( .A1(n7549), .A2(n7203), .ZN(n7202) );
  NAND2_X1 U8499 ( .A1(n7551), .A2(n7204), .ZN(n7203) );
  AOI21_X1 U8500 ( .B1(n7551), .B2(n7553), .A(n6782), .ZN(n7549) );
  INV_X1 U8501 ( .A(n7800), .ZN(n7204) );
  INV_X1 U8502 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n7979) );
  XNOR2_X1 U8503 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n7959) );
  NAND2_X1 U8504 ( .A1(n7797), .A2(n7796), .ZN(n7946) );
  INV_X1 U8505 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7795) );
  NOR2_X1 U8506 ( .A1(n8010), .A2(n7165), .ZN(n7164) );
  NAND2_X1 U8507 ( .A1(n7906), .A2(n7163), .ZN(n7162) );
  NAND2_X1 U8508 ( .A1(n8010), .A2(n7165), .ZN(n7163) );
  XNOR2_X1 U8509 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7882) );
  NOR2_X1 U8510 ( .A1(n8406), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7881) );
  INV_X1 U8511 ( .A(n12447), .ZN(n7052) );
  AND2_X1 U8512 ( .A1(n7449), .A2(n12439), .ZN(n7053) );
  OR2_X1 U8513 ( .A1(n10761), .A2(n10765), .ZN(n13855) );
  INV_X1 U8514 ( .A(n13808), .ZN(n7023) );
  AOI21_X1 U8515 ( .B1(n7029), .B2(n7032), .A(n7028), .ZN(n7027) );
  NOR2_X1 U8516 ( .A1(n13801), .A2(n13800), .ZN(n7028) );
  NOR2_X1 U8517 ( .A1(n7441), .A2(n13802), .ZN(n7029) );
  NAND2_X1 U8518 ( .A1(n7032), .A2(n7031), .ZN(n7030) );
  INV_X1 U8519 ( .A(n13802), .ZN(n7031) );
  OR2_X1 U8520 ( .A1(n8597), .A2(n11489), .ZN(n8621) );
  NAND2_X1 U8521 ( .A1(n10957), .A2(n14272), .ZN(n7044) );
  NAND2_X1 U8522 ( .A1(n10957), .A2(n7046), .ZN(n7045) );
  INV_X1 U8523 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8644) );
  NOR2_X1 U8524 ( .A1(n6769), .A2(n7042), .ZN(n7041) );
  INV_X1 U8525 ( .A(n13731), .ZN(n7042) );
  NAND2_X1 U8526 ( .A1(n12403), .A2(n7450), .ZN(n7449) );
  INV_X1 U8527 ( .A(n7452), .ZN(n7450) );
  NAND2_X1 U8528 ( .A1(n8843), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8865) );
  NAND2_X1 U8529 ( .A1(n13851), .A2(n13731), .ZN(n13892) );
  INV_X1 U8530 ( .A(n13855), .ZN(n13907) );
  INV_X1 U8531 ( .A(n12707), .ZN(n10963) );
  AND4_X1 U8532 ( .A1(n9136), .A2(n9135), .A3(n9134), .A4(n9133), .ZN(n13809)
         );
  INV_X1 U8533 ( .A(n8514), .ZN(n9112) );
  AND2_X1 U8534 ( .A1(n12352), .A2(n12351), .ZN(n14038) );
  OR2_X1 U8535 ( .A1(n10877), .A2(n10876), .ZN(n14043) );
  INV_X1 U8536 ( .A(n7472), .ZN(n7471) );
  AND2_X1 U8537 ( .A1(n7124), .A2(n7122), .ZN(n7121) );
  NAND2_X1 U8538 ( .A1(n9735), .A2(n7115), .ZN(n7122) );
  NAND2_X1 U8539 ( .A1(n7125), .A2(n9738), .ZN(n7124) );
  AND2_X1 U8540 ( .A1(n7116), .A2(n7123), .ZN(n7115) );
  AND2_X1 U8541 ( .A1(n10955), .A2(n10765), .ZN(n13906) );
  AOI21_X1 U8542 ( .B1(n7512), .B2(n7514), .A(n6693), .ZN(n7510) );
  INV_X1 U8543 ( .A(n7512), .ZN(n7511) );
  XNOR2_X1 U8544 ( .A(n14091), .B(n13921), .ZN(n14088) );
  NAND2_X1 U8545 ( .A1(n9732), .A2(n9731), .ZN(n14099) );
  AOI21_X1 U8546 ( .B1(n7110), .B2(n9677), .A(n14117), .ZN(n7109) );
  AND2_X1 U8547 ( .A1(n14315), .A2(n9678), .ZN(n14118) );
  NAND2_X1 U8548 ( .A1(n14118), .A2(n14117), .ZN(n14116) );
  NAND2_X1 U8549 ( .A1(n6932), .A2(n9671), .ZN(n14195) );
  NAND2_X1 U8550 ( .A1(n6930), .A2(n6928), .ZN(n6932) );
  NOR2_X1 U8551 ( .A1(n6929), .A2(n9670), .ZN(n6928) );
  NAND2_X1 U8552 ( .A1(n12485), .A2(n9714), .ZN(n14264) );
  NAND2_X1 U8553 ( .A1(n12487), .A2(n12486), .ZN(n12485) );
  OR2_X1 U8554 ( .A1(n8771), .A2(n8770), .ZN(n8792) );
  NAND2_X1 U8555 ( .A1(n7613), .A2(n6685), .ZN(n7607) );
  NAND2_X1 U8556 ( .A1(n11807), .A2(n7474), .ZN(n12197) );
  OR2_X1 U8557 ( .A1(n8699), .A2(n8698), .ZN(n8719) );
  INV_X1 U8558 ( .A(n6886), .ZN(n7475) );
  NAND2_X1 U8559 ( .A1(n7105), .A2(n9701), .ZN(n11849) );
  INV_X1 U8560 ( .A(n7344), .ZN(n7106) );
  NAND2_X1 U8561 ( .A1(n6940), .A2(n9660), .ZN(n11860) );
  NAND2_X1 U8562 ( .A1(n11807), .A2(n11994), .ZN(n11888) );
  NAND2_X1 U8563 ( .A1(n6936), .A2(n9655), .ZN(n11385) );
  NAND2_X1 U8564 ( .A1(n6935), .A2(n6933), .ZN(n6936) );
  NAND2_X1 U8565 ( .A1(n11386), .A2(n11580), .ZN(n11524) );
  NAND2_X1 U8566 ( .A1(n11563), .A2(n15662), .ZN(n11326) );
  OAI21_X1 U8567 ( .B1(n11842), .B2(n11833), .A(n9687), .ZN(n10890) );
  NAND2_X1 U8568 ( .A1(n7588), .A2(n15691), .ZN(n11833) );
  INV_X1 U8569 ( .A(n13947), .ZN(n7588) );
  NAND2_X1 U8570 ( .A1(n14150), .A2(n9728), .ZN(n14130) );
  INV_X1 U8571 ( .A(n7465), .ZN(n14133) );
  NAND2_X1 U8572 ( .A1(n7329), .A2(n7614), .ZN(n14148) );
  AND3_X1 U8573 ( .A1(n14186), .A2(n14293), .A3(n14185), .ZN(n14336) );
  NAND2_X1 U8574 ( .A1(n7521), .A2(n7523), .ZN(n15266) );
  NAND2_X1 U8575 ( .A1(n7526), .A2(n6687), .ZN(n7521) );
  INV_X1 U8576 ( .A(n7532), .ZN(n7531) );
  OAI21_X1 U8577 ( .B1(n8469), .B2(n7793), .A(n7533), .ZN(n7532) );
  INV_X1 U8578 ( .A(n15722), .ZN(n15285) );
  OR2_X1 U8579 ( .A1(n9685), .A2(n10963), .ZN(n15710) );
  NOR2_X1 U8580 ( .A1(n15686), .A2(n9770), .ZN(n11556) );
  NOR2_X1 U8581 ( .A1(n8392), .A2(n8836), .ZN(n6926) );
  CLKBUF_X1 U8582 ( .A(n8374), .Z(n8837) );
  NAND2_X1 U8583 ( .A1(n8474), .A2(n8366), .ZN(n8511) );
  NAND2_X1 U8584 ( .A1(n6705), .A2(n12759), .ZN(n7498) );
  AND2_X1 U8585 ( .A1(n12681), .A2(n7259), .ZN(n7257) );
  NAND2_X1 U8586 ( .A1(n15346), .A2(n15347), .ZN(n7258) );
  AND2_X1 U8587 ( .A1(n12828), .A2(n12826), .ZN(n14474) );
  INV_X1 U8588 ( .A(n14828), .ZN(n14761) );
  OAI21_X1 U8589 ( .B1(n11688), .B2(n11687), .A(n11686), .ZN(n11689) );
  NAND2_X1 U8590 ( .A1(n10222), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10246) );
  AND2_X1 U8591 ( .A1(n14495), .A2(n12805), .ZN(n14448) );
  AND2_X1 U8592 ( .A1(n14472), .A2(n12815), .ZN(n14497) );
  NAND2_X1 U8593 ( .A1(n10527), .A2(n10526), .ZN(n11373) );
  INV_X1 U8594 ( .A(n10524), .ZN(n10527) );
  NOR2_X1 U8595 ( .A1(n10259), .A2(n14459), .ZN(n10266) );
  OR2_X1 U8596 ( .A1(n14457), .A2(n7251), .ZN(n7245) );
  INV_X1 U8597 ( .A(n10278), .ZN(n10296) );
  NAND2_X1 U8598 ( .A1(n10296), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n10295) );
  INV_X1 U8599 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10119) );
  OR2_X1 U8600 ( .A1(n14485), .A2(n12759), .ZN(n7500) );
  NOR3_X1 U8601 ( .A1(n10480), .A2(n10479), .A3(n10478), .ZN(n10481) );
  AND4_X1 U8602 ( .A1(n9913), .A2(n9912), .A3(n9911), .A4(n9910), .ZN(n12853)
         );
  CLKBUF_X1 U8603 ( .A(n6674), .Z(n10297) );
  OR2_X1 U8604 ( .A1(n6674), .A2(n9933), .ZN(n9936) );
  INV_X1 U8605 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9208) );
  AND2_X1 U8606 ( .A1(n7584), .A2(n10012), .ZN(n10216) );
  NOR2_X1 U8607 ( .A1(n7714), .A2(n7711), .ZN(n7710) );
  INV_X1 U8608 ( .A(n7753), .ZN(n7713) );
  NAND2_X1 U8609 ( .A1(n7015), .A2(n6695), .ZN(n14781) );
  INV_X1 U8610 ( .A(n7752), .ZN(n7354) );
  NAND2_X1 U8611 ( .A1(n14832), .A2(n7288), .ZN(n14797) );
  NAND2_X1 U8612 ( .A1(n14832), .A2(n15008), .ZN(n14812) );
  AND2_X1 U8613 ( .A1(n15026), .A2(n14718), .ZN(n14844) );
  NAND2_X1 U8614 ( .A1(n14905), .A2(n7297), .ZN(n14863) );
  NOR2_X1 U8615 ( .A1(n15024), .A2(n7298), .ZN(n7297) );
  INV_X1 U8616 ( .A(n7299), .ZN(n7298) );
  NAND2_X1 U8617 ( .A1(n7706), .A2(n14756), .ZN(n14862) );
  NAND2_X1 U8618 ( .A1(n14754), .A2(n7707), .ZN(n7706) );
  NAND2_X1 U8619 ( .A1(n14862), .A2(n14864), .ZN(n14861) );
  NAND2_X1 U8620 ( .A1(n14905), .A2(n7300), .ZN(n14893) );
  NAND2_X1 U8621 ( .A1(n14905), .A2(n14911), .ZN(n14906) );
  NOR2_X1 U8622 ( .A1(n14913), .A2(n7696), .ZN(n7694) );
  NAND2_X1 U8623 ( .A1(n14687), .A2(n15324), .ZN(n14970) );
  NOR2_X1 U8624 ( .A1(n14970), .A2(n15064), .ZN(n14952) );
  AND2_X1 U8625 ( .A1(n7362), .A2(n14704), .ZN(n7359) );
  NAND2_X1 U8626 ( .A1(n7361), .A2(n14965), .ZN(n7363) );
  NAND2_X1 U8627 ( .A1(n7364), .A2(n12692), .ZN(n14702) );
  NAND2_X1 U8628 ( .A1(n7676), .A2(n7675), .ZN(n12643) );
  AOI21_X1 U8629 ( .B1(n7677), .B2(n7679), .A(n6765), .ZN(n7675) );
  OR2_X1 U8630 ( .A1(n12644), .A2(n15342), .ZN(n12645) );
  OR2_X1 U8631 ( .A1(n10120), .A2(n10119), .ZN(n10139) );
  NOR2_X1 U8632 ( .A1(n10139), .A2(n12683), .ZN(n10153) );
  OAI21_X1 U8633 ( .B1(n12598), .B2(n7679), .A(n7677), .ZN(n12607) );
  NAND2_X1 U8634 ( .A1(n12602), .A2(n12532), .ZN(n12533) );
  NAND2_X1 U8635 ( .A1(n12598), .A2(n12531), .ZN(n12602) );
  NAND2_X1 U8636 ( .A1(n12310), .A2(n6686), .ZN(n12592) );
  NAND2_X1 U8637 ( .A1(n12310), .A2(n15537), .ZN(n12475) );
  AND2_X1 U8638 ( .A1(n12301), .A2(n12303), .ZN(n7719) );
  NAND2_X1 U8639 ( .A1(n12304), .A2(n12303), .ZN(n12305) );
  NOR2_X1 U8640 ( .A1(n10071), .A2(n10070), .ZN(n10085) );
  NAND2_X1 U8641 ( .A1(n12057), .A2(n12056), .ZN(n12246) );
  NOR2_X1 U8642 ( .A1(n12048), .A2(n12248), .ZN(n12258) );
  NAND2_X1 U8643 ( .A1(n12002), .A2(n12049), .ZN(n12057) );
  OR2_X1 U8644 ( .A1(n11998), .A2(n12055), .ZN(n12048) );
  AND2_X1 U8645 ( .A1(n10467), .A2(n12000), .ZN(n12003) );
  OR2_X1 U8646 ( .A1(n10578), .A2(n10931), .ZN(n14967) );
  NAND2_X1 U8647 ( .A1(n10783), .A2(n10931), .ZN(n14966) );
  NAND2_X1 U8648 ( .A1(n12170), .A2(n12083), .ZN(n11998) );
  NOR2_X1 U8649 ( .A1(n15502), .A2(n12131), .ZN(n12169) );
  AND2_X1 U8650 ( .A1(n12169), .A2(n15528), .ZN(n12170) );
  INV_X1 U8651 ( .A(n14966), .ZN(n14825) );
  INV_X1 U8652 ( .A(n14967), .ZN(n14827) );
  INV_X1 U8653 ( .A(n15534), .ZN(n15393) );
  AND2_X1 U8654 ( .A1(n11438), .A2(n11437), .ZN(n11503) );
  INV_X1 U8655 ( .A(n15529), .ZN(n15549) );
  INV_X1 U8656 ( .A(n15061), .ZN(n15503) );
  NAND2_X1 U8657 ( .A1(n10563), .A2(n10565), .ZN(n15545) );
  INV_X1 U8658 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9902) );
  XNOR2_X1 U8659 ( .A(n9126), .B(n9125), .ZN(n12860) );
  NOR2_X1 U8660 ( .A1(n7717), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n7716) );
  NOR2_X1 U8661 ( .A1(n9076), .A2(SI_27_), .ZN(n7671) );
  NAND2_X1 U8662 ( .A1(n9076), .A2(SI_27_), .ZN(n7670) );
  INV_X1 U8663 ( .A(n7717), .ZN(n7715) );
  XNOR2_X1 U8664 ( .A(n10498), .B(P1_IR_REG_26__SCAN_IN), .ZN(n10558) );
  XNOR2_X1 U8665 ( .A(n10489), .B(n10488), .ZN(n10782) );
  OAI21_X1 U8666 ( .B1(n10487), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10489) );
  INV_X1 U8667 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9927) );
  INV_X1 U8668 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9922) );
  INV_X1 U8669 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9921) );
  NAND2_X1 U8670 ( .A1(n8690), .A2(n8689), .ZN(n8713) );
  AOI21_X1 U8671 ( .B1(n7647), .B2(n7649), .A(n7645), .ZN(n7644) );
  NAND2_X1 U8672 ( .A1(n8613), .A2(n7647), .ZN(n7646) );
  INV_X1 U8673 ( .A(n8659), .ZN(n7645) );
  OAI21_X1 U8674 ( .B1(n10187), .B2(P1_IR_REG_8__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10160) );
  OR2_X1 U8675 ( .A1(n10077), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n10187) );
  CLKBUF_X1 U8676 ( .A(n9979), .Z(n9980) );
  NOR2_X1 U8677 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n9960) );
  AND2_X1 U8678 ( .A1(n7306), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n9266) );
  INV_X1 U8679 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7306) );
  INV_X1 U8680 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n9574) );
  NAND2_X1 U8681 ( .A1(n6993), .A2(n6991), .ZN(n9265) );
  NAND2_X1 U8682 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n6992), .ZN(n6991) );
  NAND2_X1 U8683 ( .A1(n6878), .A2(n9266), .ZN(n6993) );
  INV_X1 U8684 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6992) );
  NOR2_X1 U8685 ( .A1(n15125), .A2(n9282), .ZN(n9283) );
  NOR2_X1 U8686 ( .A1(n15128), .A2(n9289), .ZN(n9290) );
  AND2_X1 U8687 ( .A1(n15135), .A2(n15134), .ZN(n9296) );
  OAI21_X1 U8688 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n9240), .A(n9239), .ZN(
        n9249) );
  NAND2_X1 U8689 ( .A1(n12153), .A2(n12152), .ZN(n12151) );
  INV_X1 U8690 ( .A(n7390), .ZN(n7386) );
  AND2_X1 U8691 ( .A1(n7387), .A2(n7384), .ZN(n7383) );
  NAND2_X1 U8692 ( .A1(n9847), .A2(n12952), .ZN(n12709) );
  NAND2_X1 U8693 ( .A1(n12450), .A2(n6815), .ZN(n12517) );
  NAND2_X1 U8694 ( .A1(n12450), .A2(n9805), .ZN(n12516) );
  OR2_X1 U8695 ( .A1(n9879), .A2(n12321), .ZN(n13016) );
  NAND2_X1 U8696 ( .A1(n7374), .A2(n7376), .ZN(n11735) );
  NAND2_X1 U8697 ( .A1(n9830), .A2(n9829), .ZN(n12892) );
  AND2_X1 U8698 ( .A1(n12870), .A2(n7004), .ZN(n7003) );
  AND2_X1 U8699 ( .A1(n12865), .A2(n13023), .ZN(n7004) );
  NAND2_X1 U8700 ( .A1(n8338), .A2(n8337), .ZN(n13415) );
  NAND2_X1 U8701 ( .A1(n9788), .A2(n9786), .ZN(n11263) );
  NAND2_X1 U8702 ( .A1(n12967), .A2(n9835), .ZN(n12903) );
  XNOR2_X1 U8703 ( .A(n9820), .B(n13559), .ZN(n12935) );
  NAND2_X1 U8704 ( .A1(n12265), .A2(n9801), .ZN(n12452) );
  INV_X1 U8705 ( .A(n13518), .ZN(n13547) );
  INV_X1 U8706 ( .A(n7372), .ZN(n7371) );
  NAND2_X1 U8707 ( .A1(n8164), .A2(n8163), .ZN(n13499) );
  XNOR2_X1 U8708 ( .A(n9827), .B(n13560), .ZN(n13001) );
  NAND2_X1 U8709 ( .A1(n8122), .A2(n8121), .ZN(n13550) );
  INV_X1 U8710 ( .A(n13023), .ZN(n13008) );
  NAND2_X1 U8711 ( .A1(n12026), .A2(n12025), .ZN(n12024) );
  OR2_X1 U8712 ( .A1(n9879), .A2(n12285), .ZN(n13028) );
  AND2_X1 U8713 ( .A1(n7397), .A2(n9813), .ZN(n7394) );
  NAND2_X1 U8714 ( .A1(n12913), .A2(n9813), .ZN(n7396) );
  AND2_X1 U8715 ( .A1(n11723), .A2(n11722), .ZN(n15161) );
  INV_X1 U8716 ( .A(n13448), .ZN(n11520) );
  INV_X1 U8717 ( .A(n13433), .ZN(n13467) );
  NAND2_X1 U8718 ( .A1(n8192), .A2(n8191), .ZN(n13483) );
  NAND2_X1 U8719 ( .A1(n8010), .A2(n7770), .ZN(n7265) );
  NAND2_X1 U8720 ( .A1(n7894), .A2(P3_IR_REG_2__SCAN_IN), .ZN(n7266) );
  AND2_X1 U8721 ( .A1(n11140), .A2(n7412), .ZN(n11024) );
  INV_X1 U8722 ( .A(n7282), .ZN(n11151) );
  AND2_X1 U8723 ( .A1(n7920), .A2(n7919), .ZN(n11162) );
  NAND2_X1 U8724 ( .A1(n7424), .A2(n7426), .ZN(n11201) );
  INV_X1 U8725 ( .A(n7149), .ZN(n11287) );
  INV_X1 U8726 ( .A(n7147), .ZN(n11285) );
  INV_X1 U8727 ( .A(n7144), .ZN(n11305) );
  INV_X1 U8728 ( .A(n7405), .ZN(n11409) );
  INV_X1 U8729 ( .A(n7419), .ZN(n11406) );
  XNOR2_X1 U8730 ( .A(n10624), .B(n10623), .ZN(n11700) );
  NAND2_X1 U8731 ( .A1(n7430), .A2(n7429), .ZN(n12411) );
  INV_X1 U8732 ( .A(n10606), .ZN(n7429) );
  INV_X1 U8733 ( .A(n7430), .ZN(n10607) );
  NAND2_X1 U8734 ( .A1(n7417), .A2(n12426), .ZN(n7416) );
  INV_X1 U8735 ( .A(n12423), .ZN(n7417) );
  NOR2_X1 U8736 ( .A1(n15734), .A2(n15735), .ZN(n15733) );
  INV_X1 U8737 ( .A(n7263), .ZN(n15742) );
  INV_X1 U8738 ( .A(n7428), .ZN(n12416) );
  XNOR2_X1 U8739 ( .A(n6988), .B(n15124), .ZN(n13248) );
  INV_X1 U8740 ( .A(n7264), .ZN(n13268) );
  INV_X1 U8741 ( .A(n7413), .ZN(n13274) );
  INV_X1 U8742 ( .A(n7143), .ZN(n13298) );
  NOR2_X1 U8743 ( .A1(n15143), .A2(n15144), .ZN(n15142) );
  XNOR2_X1 U8744 ( .A(n13353), .B(n13361), .ZN(n13331) );
  INV_X1 U8745 ( .A(n13364), .ZN(n13366) );
  NAND2_X1 U8746 ( .A1(n8209), .A2(n13405), .ZN(n13406) );
  OR2_X1 U8747 ( .A1(n13410), .A2(n13409), .ZN(n13414) );
  NAND2_X1 U8748 ( .A1(n6948), .A2(n6947), .ZN(n8339) );
  NAND2_X1 U8749 ( .A1(n7317), .A2(n7315), .ZN(n13431) );
  NAND2_X1 U8750 ( .A1(n8248), .A2(n8247), .ZN(n13493) );
  OAI21_X1 U8751 ( .B1(n13522), .B2(n7324), .A(n7322), .ZN(n13498) );
  AOI21_X1 U8752 ( .B1(n11660), .B2(n6677), .A(n8143), .ZN(n13528) );
  NAND2_X1 U8753 ( .A1(n13563), .A2(n13093), .ZN(n13549) );
  NAND2_X1 U8754 ( .A1(n8108), .A2(n8107), .ZN(n13568) );
  NAND2_X1 U8755 ( .A1(n13578), .A2(n13577), .ZN(n13580) );
  NAND2_X1 U8756 ( .A1(n8083), .A2(n13185), .ZN(n13578) );
  NAND2_X1 U8757 ( .A1(n8076), .A2(n8075), .ZN(n13179) );
  NAND2_X1 U8758 ( .A1(n6945), .A2(n6944), .ZN(n8237) );
  AND2_X1 U8759 ( .A1(n6945), .A2(n6731), .ZN(n15171) );
  NAND2_X1 U8760 ( .A1(n6910), .A2(n13166), .ZN(n15192) );
  NAND2_X1 U8761 ( .A1(n12283), .A2(n7638), .ZN(n12121) );
  NAND2_X1 U8762 ( .A1(n12281), .A2(n7985), .ZN(n12124) );
  NOR2_X1 U8763 ( .A1(n11466), .A2(n15798), .ZN(n15217) );
  AND2_X1 U8764 ( .A1(n15801), .A2(n15754), .ZN(n15218) );
  AND2_X1 U8765 ( .A1(n15801), .A2(n15795), .ZN(n15819) );
  AOI21_X1 U8766 ( .B1(n13586), .B2(n15241), .A(n13587), .ZN(n13641) );
  INV_X1 U8767 ( .A(n12920), .ZN(n13651) );
  INV_X1 U8768 ( .A(n12951), .ZN(n13655) );
  AND2_X1 U8769 ( .A1(n8175), .A2(n8174), .ZN(n13659) );
  NAND2_X1 U8770 ( .A1(n8134), .A2(n8133), .ZN(n13671) );
  AND3_X1 U8771 ( .A1(n7984), .A2(n7983), .A3(n7982), .ZN(n15759) );
  OR2_X1 U8772 ( .A1(n6669), .A2(n9388), .ZN(n7875) );
  AND2_X1 U8773 ( .A1(n9874), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13685) );
  NAND2_X1 U8774 ( .A1(n7227), .A2(n7225), .ZN(n13039) );
  AND2_X1 U8775 ( .A1(n7227), .A2(n7229), .ZN(n13048) );
  AOI21_X1 U8776 ( .B1(n8336), .B2(n8325), .A(n6833), .ZN(n13037) );
  INV_X1 U8777 ( .A(n7849), .ZN(n13697) );
  AND2_X1 U8778 ( .A1(n6969), .A2(n6968), .ZN(n6967) );
  XNOR2_X1 U8779 ( .A(n8183), .B(n15102), .ZN(n12495) );
  INV_X1 U8780 ( .A(SI_16_), .ZN(n10975) );
  NAND2_X1 U8781 ( .A1(n7545), .A2(n7814), .ZN(n8086) );
  NAND2_X1 U8782 ( .A1(n8070), .A2(n8069), .ZN(n7545) );
  INV_X1 U8783 ( .A(SI_15_), .ZN(n10864) );
  NAND2_X1 U8784 ( .A1(n7222), .A2(n7808), .ZN(n8027) );
  OR2_X1 U8785 ( .A1(n8021), .A2(n7807), .ZN(n7222) );
  INV_X1 U8786 ( .A(SI_11_), .ZN(n10724) );
  INV_X1 U8787 ( .A(SI_10_), .ZN(n10720) );
  NAND2_X1 U8788 ( .A1(n7550), .A2(n7803), .ZN(n7995) );
  NAND2_X1 U8789 ( .A1(n7975), .A2(n7973), .ZN(n7550) );
  INV_X1 U8790 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7962) );
  INV_X1 U8791 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7947) );
  AND2_X1 U8792 ( .A1(n7214), .A2(n7216), .ZN(n7932) );
  INV_X1 U8793 ( .A(n11162), .ZN(n10706) );
  NAND2_X1 U8794 ( .A1(n7542), .A2(n7792), .ZN(n7916) );
  NAND2_X1 U8795 ( .A1(n7905), .A2(n7903), .ZN(n7542) );
  INV_X1 U8796 ( .A(n7432), .ZN(n7431) );
  OAI21_X1 U8797 ( .B1(n7435), .B2(n8010), .A(n7433), .ZN(n7432) );
  OR2_X1 U8798 ( .A1(n10507), .A2(n10762), .ZN(n10764) );
  NAND2_X1 U8799 ( .A1(n7026), .A2(n7032), .ZN(n13803) );
  NAND2_X1 U8800 ( .A1(n12183), .A2(n7057), .ZN(n7056) );
  NOR2_X1 U8801 ( .A1(n11902), .A2(n7457), .ZN(n7456) );
  INV_X1 U8802 ( .A(n11899), .ZN(n7457) );
  NAND2_X1 U8803 ( .A1(n11900), .A2(n11899), .ZN(n11901) );
  NAND2_X1 U8804 ( .A1(n7018), .A2(n11120), .ZN(n13780) );
  INV_X1 U8805 ( .A(n13778), .ZN(n11120) );
  OAI21_X1 U8806 ( .B1(n7027), .B2(n13808), .A(n7021), .ZN(n7020) );
  NAND2_X1 U8807 ( .A1(n7027), .A2(n7022), .ZN(n7021) );
  NAND2_X1 U8808 ( .A1(n7030), .A2(n7023), .ZN(n7022) );
  NAND2_X1 U8809 ( .A1(n7025), .A2(n13808), .ZN(n7024) );
  INV_X1 U8810 ( .A(n7030), .ZN(n7025) );
  AND2_X1 U8811 ( .A1(n11750), .A2(n11742), .ZN(n7017) );
  NAND2_X1 U8812 ( .A1(n10760), .A2(n7593), .ZN(n7594) );
  AND2_X1 U8813 ( .A1(n9919), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7593) );
  AOI21_X1 U8814 ( .B1(n7038), .B2(n7040), .A(n7035), .ZN(n7034) );
  INV_X1 U8815 ( .A(n13863), .ZN(n7035) );
  NAND2_X1 U8816 ( .A1(n8932), .A2(n8931), .ZN(n14337) );
  NAND2_X1 U8817 ( .A1(n12185), .A2(n12184), .ZN(n12400) );
  NAND2_X1 U8818 ( .A1(n13723), .A2(n13722), .ZN(n13832) );
  AND2_X1 U8819 ( .A1(n13722), .A2(n13724), .ZN(n7463) );
  NAND2_X1 U8820 ( .A1(n7037), .A2(n7458), .ZN(n13865) );
  NAND2_X1 U8821 ( .A1(n13851), .A2(n7041), .ZN(n7037) );
  NAND2_X1 U8822 ( .A1(n8909), .A2(n8908), .ZN(n14341) );
  OAI21_X1 U8823 ( .B1(n12185), .B2(n7455), .A(n7452), .ZN(n12402) );
  AND2_X1 U8824 ( .A1(n11347), .A2(n11339), .ZN(n7462) );
  INV_X1 U8825 ( .A(n11346), .ZN(n11347) );
  NAND2_X1 U8826 ( .A1(n11340), .A2(n11339), .ZN(n11345) );
  NAND2_X1 U8827 ( .A1(n11123), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13912) );
  NAND2_X1 U8828 ( .A1(n7446), .A2(n7447), .ZN(n7445) );
  AOI21_X1 U8829 ( .B1(n9172), .B2(n12707), .A(n7754), .ZN(n9192) );
  AND2_X1 U8830 ( .A1(n9194), .A2(n8372), .ZN(n7439) );
  NAND4_X1 U8831 ( .A1(n8459), .A2(n8458), .A3(n8457), .A4(n8456), .ZN(n13945)
         );
  NAND2_X1 U8832 ( .A1(n8464), .A2(n8455), .ZN(n8459) );
  NAND2_X1 U8833 ( .A1(n8542), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8466) );
  INV_X1 U8834 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7836) );
  NAND2_X1 U8835 ( .A1(n9040), .A2(n9039), .ZN(n14108) );
  OAI21_X1 U8836 ( .B1(n14150), .B2(n9677), .A(n7110), .ZN(n14113) );
  NAND2_X1 U8837 ( .A1(n14147), .A2(n9676), .ZN(n14140) );
  NAND2_X1 U8838 ( .A1(n8982), .A2(n8981), .ZN(n14159) );
  NAND2_X1 U8839 ( .A1(n7619), .A2(n7617), .ZN(n14169) );
  NAND2_X1 U8840 ( .A1(n6930), .A2(n7527), .ZN(n14221) );
  NAND2_X1 U8841 ( .A1(n14250), .A2(n7528), .ZN(n14237) );
  NAND2_X1 U8842 ( .A1(n14243), .A2(n9718), .ZN(n14229) );
  NAND2_X1 U8843 ( .A1(n8842), .A2(n8841), .ZN(n14359) );
  NAND2_X1 U8844 ( .A1(n12483), .A2(n9667), .ZN(n14275) );
  NAND2_X1 U8845 ( .A1(n8815), .A2(n8814), .ZN(n14364) );
  NAND2_X1 U8846 ( .A1(n8791), .A2(n8790), .ZN(n12570) );
  OR2_X1 U8847 ( .A1(n15652), .A2(n15672), .ZN(n15663) );
  NAND2_X1 U8848 ( .A1(n7613), .A2(n9708), .ZN(n12194) );
  INV_X1 U8849 ( .A(n7762), .ZN(n7524) );
  NAND2_X1 U8850 ( .A1(n7526), .A2(n7763), .ZN(n7525) );
  NAND2_X1 U8851 ( .A1(n7586), .A2(n9700), .ZN(n11810) );
  NAND2_X1 U8852 ( .A1(n9659), .A2(n9658), .ZN(n11646) );
  NAND2_X1 U8853 ( .A1(n11523), .A2(n11526), .ZN(n9659) );
  NAND2_X1 U8854 ( .A1(n6935), .A2(n9653), .ZN(n11325) );
  OR2_X1 U8855 ( .A1(n10760), .A2(n8450), .ZN(n8452) );
  OR2_X1 U8856 ( .A1(n11561), .A2(n14272), .ZN(n15654) );
  INV_X1 U8857 ( .A(n14261), .ZN(n15269) );
  OAI21_X1 U8858 ( .B1(n10884), .B2(n8510), .A(n8668), .ZN(n11991) );
  AND2_X1 U8859 ( .A1(n9105), .A2(n9104), .ZN(n14377) );
  INV_X1 U8860 ( .A(n14159), .ZN(n14391) );
  NAND2_X1 U8861 ( .A1(n8961), .A2(n8960), .ZN(n14394) );
  INV_X1 U8862 ( .A(n15686), .ZN(n15689) );
  OR2_X1 U8863 ( .A1(n8395), .A2(n7736), .ZN(n8414) );
  NAND2_X1 U8864 ( .A1(n7738), .A2(n8410), .ZN(n7736) );
  XNOR2_X1 U8865 ( .A(n9196), .B(n9195), .ZN(n14431) );
  OAI21_X1 U8866 ( .B1(n9194), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9196) );
  INV_X1 U8867 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12559) );
  INV_X1 U8868 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n12066) );
  INV_X1 U8869 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11987) );
  INV_X1 U8870 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11820) );
  INV_X1 U8871 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10750) );
  AND2_X1 U8872 ( .A1(n8571), .A2(n8615), .ZN(n13995) );
  CLKBUF_X1 U8873 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n15565) );
  NAND2_X1 U8874 ( .A1(n12071), .A2(n12070), .ZN(n12075) );
  XNOR2_X1 U8875 ( .A(n7252), .B(n14436), .ZN(n14437) );
  NAND2_X1 U8876 ( .A1(n14539), .A2(n12837), .ZN(n7252) );
  NOR2_X1 U8877 ( .A1(n10568), .A2(n10569), .ZN(n11688) );
  NOR2_X1 U8878 ( .A1(n7489), .A2(n12852), .ZN(n7486) );
  OAI22_X1 U8879 ( .A1(n7489), .A2(n7488), .B1(n12852), .B2(n7491), .ZN(n7487)
         );
  NOR2_X1 U8880 ( .A1(n14436), .A2(n12852), .ZN(n7488) );
  INV_X1 U8881 ( .A(n12852), .ZN(n7490) );
  NAND2_X1 U8882 ( .A1(n10387), .A2(n10386), .ZN(n14779) );
  INV_X1 U8883 ( .A(n7495), .ZN(n12545) );
  NAND2_X1 U8884 ( .A1(n12234), .A2(n12233), .ZN(n12235) );
  INV_X1 U8885 ( .A(n14563), .ZN(n11616) );
  NAND2_X1 U8886 ( .A1(n12778), .A2(n12777), .ZN(n14466) );
  NAND2_X1 U8887 ( .A1(n14515), .A2(n14514), .ZN(n12778) );
  AND2_X1 U8888 ( .A1(n7258), .A2(n7259), .ZN(n12682) );
  AND4_X1 U8889 ( .A1(n10215), .A2(n10214), .A3(n10213), .A4(n10212), .ZN(
        n15325) );
  NAND2_X1 U8890 ( .A1(n11689), .A2(n14505), .ZN(n11690) );
  NAND2_X1 U8891 ( .A1(n14457), .A2(n12773), .ZN(n14515) );
  NAND2_X1 U8892 ( .A1(n12727), .A2(n12726), .ZN(n15338) );
  NAND2_X1 U8893 ( .A1(n7248), .A2(n7246), .ZN(n12796) );
  NAND2_X1 U8894 ( .A1(n10532), .A2(n10534), .ZN(n10535) );
  AND2_X1 U8895 ( .A1(n14735), .A2(n14732), .ZN(n15348) );
  NAND2_X1 U8896 ( .A1(n7500), .A2(n12758), .ZN(n14530) );
  NAND2_X1 U8897 ( .A1(n10244), .A2(n10243), .ZN(n15057) );
  NAND2_X1 U8898 ( .A1(n7484), .A2(n7482), .ZN(n12071) );
  AND2_X1 U8899 ( .A1(n6690), .A2(n11947), .ZN(n7482) );
  AND2_X1 U8900 ( .A1(n7484), .A2(n6690), .ZN(n11948) );
  AND4_X1 U8901 ( .A1(n10183), .A2(n10182), .A3(n10181), .A4(n10180), .ZN(
        n15362) );
  NAND2_X1 U8902 ( .A1(n11374), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15369) );
  INV_X1 U8903 ( .A(n15337), .ZN(n15365) );
  OR3_X1 U8904 ( .A1(n10408), .A2(n10407), .A3(n10406), .ZN(n14690) );
  INV_X1 U8905 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n12317) );
  AND4_X1 U8906 ( .A1(n10254), .A2(n10253), .A3(n10252), .A4(n10251), .ZN(
        n14489) );
  NAND3_X2 U8907 ( .A1(n6715), .A2(n9959), .A3(n7673), .ZN(n10536) );
  OR2_X1 U8908 ( .A1(n6675), .A2(n14576), .ZN(n9959) );
  INV_X1 U8909 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7835) );
  AND2_X1 U8910 ( .A1(n10426), .A2(n10425), .ZN(n14985) );
  NAND2_X1 U8911 ( .A1(n14771), .A2(n14770), .ZN(n14769) );
  NAND2_X1 U8912 ( .A1(n14788), .A2(n7753), .ZN(n14771) );
  NAND2_X1 U8913 ( .A1(n10373), .A2(n10372), .ZN(n14802) );
  AOI21_X1 U8914 ( .B1(n14806), .B2(n14722), .A(n7711), .ZN(n14795) );
  AND2_X1 U8915 ( .A1(n14843), .A2(n14719), .ZN(n14839) );
  NAND2_X1 U8916 ( .A1(n10328), .A2(n10327), .ZN(n14859) );
  NAND2_X1 U8917 ( .A1(n14754), .A2(n14753), .ZN(n14879) );
  NAND2_X1 U8918 ( .A1(n14912), .A2(n14711), .ZN(n14890) );
  NAND2_X1 U8919 ( .A1(n14748), .A2(n14747), .ZN(n14929) );
  INV_X1 U8920 ( .A(n15057), .ZN(n14944) );
  NAND2_X1 U8921 ( .A1(n7683), .A2(n7685), .ZN(n14951) );
  NAND2_X1 U8922 ( .A1(n7684), .A2(n7688), .ZN(n7683) );
  NAND2_X1 U8923 ( .A1(n14742), .A2(n14741), .ZN(n14962) );
  NAND2_X1 U8924 ( .A1(n12622), .A2(n12621), .ZN(n12624) );
  NAND2_X1 U8925 ( .A1(n12467), .A2(n12466), .ZN(n7353) );
  NAND2_X1 U8926 ( .A1(n10115), .A2(n10114), .ZN(n15543) );
  OR2_X1 U8927 ( .A1(n10884), .A2(n10110), .ZN(n10115) );
  NAND2_X1 U8928 ( .A1(n10582), .A2(n10780), .ZN(n14975) );
  INV_X1 U8929 ( .A(n11436), .ZN(n10582) );
  OR2_X1 U8930 ( .A1(n10424), .A2(n10718), .ZN(n7291) );
  OR2_X1 U8931 ( .A1(n9964), .A2(n10110), .ZN(n7290) );
  INV_X1 U8932 ( .A(n14960), .ZN(n15506) );
  AND2_X1 U8933 ( .A1(n14735), .A2(n11829), .ZN(n15505) );
  NAND2_X1 U8934 ( .A1(n9963), .A2(n7503), .ZN(n7502) );
  AND2_X1 U8935 ( .A1(n7505), .A2(n7507), .ZN(n7503) );
  OR2_X1 U8936 ( .A1(n15509), .A2(n11826), .ZN(n15497) );
  AND2_X2 U8937 ( .A1(n11503), .A2(n14732), .ZN(n15559) );
  INV_X1 U8938 ( .A(n14986), .ZN(n7294) );
  AOI21_X1 U8939 ( .B1(n14991), .B2(n15534), .A(n14990), .ZN(n7293) );
  NAND2_X2 U8940 ( .A1(n10780), .A2(n10571), .ZN(n15510) );
  XNOR2_X1 U8941 ( .A(n9123), .B(n9122), .ZN(n10409) );
  INV_X1 U8942 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n15098) );
  INV_X1 U8943 ( .A(n9931), .ZN(n12513) );
  INV_X1 U8944 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n12296) );
  INV_X1 U8945 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n12037) );
  INV_X1 U8946 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11973) );
  INV_X1 U8947 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11804) );
  INV_X1 U8948 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n11609) );
  INV_X1 U8949 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n11178) );
  INV_X1 U8950 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10883) );
  NAND2_X1 U8951 ( .A1(n8690), .A2(n6882), .ZN(n10884) );
  NAND2_X1 U8952 ( .A1(n6883), .A2(n7195), .ZN(n6882) );
  INV_X1 U8953 ( .A(n8665), .ZN(n6883) );
  NAND2_X1 U8954 ( .A1(n8633), .A2(n8632), .ZN(n8637) );
  NAND2_X1 U8955 ( .A1(n8614), .A2(n8633), .ZN(n10793) );
  INV_X1 U8956 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10751) );
  INV_X1 U8957 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10747) );
  NAND2_X1 U8958 ( .A1(n7657), .A2(n8437), .ZN(n8408) );
  NOR2_X1 U8959 ( .A1(n15869), .A2(n9270), .ZN(n15116) );
  NAND2_X1 U8960 ( .A1(n15115), .A2(n7311), .ZN(n15866) );
  OAI21_X1 U8961 ( .B1(n15116), .B2(n15117), .A(n7312), .ZN(n7311) );
  NOR2_X1 U8962 ( .A1(n15866), .A2(n15867), .ZN(n15865) );
  XNOR2_X1 U8963 ( .A(n9272), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15856) );
  XNOR2_X1 U8964 ( .A(n6875), .B(n9275), .ZN(n15860) );
  INV_X1 U8965 ( .A(n9276), .ZN(n6875) );
  NAND2_X1 U8966 ( .A1(n15860), .A2(n15859), .ZN(n15858) );
  XNOR2_X1 U8967 ( .A(n9283), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15864) );
  NAND2_X1 U8968 ( .A1(n15864), .A2(n15863), .ZN(n15862) );
  XNOR2_X1 U8969 ( .A(n9288), .B(n9287), .ZN(n15130) );
  NOR2_X1 U8970 ( .A1(n15130), .A2(n15129), .ZN(n15128) );
  XNOR2_X1 U8971 ( .A(n9290), .B(n7304), .ZN(n15133) );
  INV_X1 U8972 ( .A(n9291), .ZN(n7304) );
  INV_X1 U8973 ( .A(n6995), .ZN(n9294) );
  INV_X1 U8974 ( .A(n9293), .ZN(n6994) );
  NOR2_X1 U8975 ( .A1(n9296), .A2(n9295), .ZN(n15419) );
  AND2_X1 U8976 ( .A1(n6874), .A2(n6873), .ZN(n15428) );
  NAND2_X1 U8977 ( .A1(n9297), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6873) );
  NAND2_X1 U8978 ( .A1(n15427), .A2(n7000), .ZN(n15432) );
  OAI21_X1 U8979 ( .B1(n15428), .B2(n15429), .A(n7001), .ZN(n7000) );
  INV_X1 U8980 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7001) );
  NAND2_X1 U8981 ( .A1(n15432), .A2(n15433), .ZN(n15431) );
  NAND2_X1 U8982 ( .A1(n7302), .A2(n15431), .ZN(n15437) );
  OAI21_X1 U8983 ( .B1(n15432), .B2(n15433), .A(n7303), .ZN(n7302) );
  INV_X1 U8984 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7303) );
  OAI21_X1 U8985 ( .B1(n15440), .B2(n15441), .A(n6999), .ZN(n6876) );
  INV_X1 U8986 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n6999) );
  NOR2_X1 U8987 ( .A1(n7012), .A2(n7011), .ZN(n7010) );
  NOR2_X1 U8988 ( .A1(n13647), .A2(n13035), .ZN(n7011) );
  NAND2_X1 U8989 ( .A1(n6844), .A2(n13244), .ZN(P3_U3296) );
  NAND2_X1 U8990 ( .A1(n6845), .A2(n9875), .ZN(n6844) );
  OAI21_X1 U8991 ( .B1(n13397), .B2(n15744), .A(n6989), .ZN(P3_U3201) );
  OAI21_X1 U8992 ( .B1(n13400), .B2(n13626), .A(n8361), .ZN(n8362) );
  OAI21_X1 U8993 ( .B1(n13641), .B2(n15851), .A(n7342), .ZN(P3_U3487) );
  INV_X1 U8994 ( .A(n7343), .ZN(n7342) );
  OAI22_X1 U8995 ( .A1(n13643), .A2(n13626), .B1(n15854), .B2(n13588), .ZN(
        n7343) );
  OAI21_X1 U8996 ( .B1(n13400), .B2(n13676), .A(n8357), .ZN(n8358) );
  OAI21_X1 U8997 ( .B1(n13641), .B2(n15844), .A(n7005), .ZN(P3_U3455) );
  INV_X1 U8998 ( .A(n7006), .ZN(n7005) );
  OAI21_X1 U8999 ( .B1(n13643), .B2(n13676), .A(n7007), .ZN(n7006) );
  OR2_X1 U9000 ( .A1(n15846), .A2(n13642), .ZN(n7007) );
  NAND2_X1 U9001 ( .A1(n13893), .A2(n7460), .ZN(n13798) );
  OAI21_X1 U9002 ( .B1(n14379), .B2(n15729), .A(n6917), .ZN(P2_U3526) );
  INV_X1 U9003 ( .A(n6918), .ZN(n6917) );
  OAI22_X1 U9004 ( .A1(n14381), .A2(n14351), .B1(n15731), .B2(n14301), .ZN(
        n6918) );
  NAND2_X1 U9005 ( .A1(n14050), .A2(n9774), .ZN(n6879) );
  OAI21_X1 U9006 ( .B1(n14287), .B2(n9771), .A(n9772), .ZN(n9777) );
  NAND2_X1 U9007 ( .A1(n7341), .A2(n7339), .ZN(P2_U3494) );
  INV_X1 U9008 ( .A(n7340), .ZN(n7339) );
  OAI22_X1 U9009 ( .A1(n14381), .A2(n14401), .B1(n15724), .B2(n14380), .ZN(
        n7340) );
  XNOR2_X1 U9010 ( .A(n7308), .B(n7307), .ZN(SUB_1596_U4) );
  XNOR2_X1 U9011 ( .A(n9645), .B(n9309), .ZN(n7307) );
  NAND2_X1 U9012 ( .A1(n7309), .A2(n15109), .ZN(n7308) );
  INV_X1 U9013 ( .A(n14244), .ZN(n7136) );
  INV_X2 U9014 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8010) );
  INV_X1 U9015 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n14406) );
  INV_X1 U9016 ( .A(n11526), .ZN(n6939) );
  AND2_X1 U9017 ( .A1(n7685), .A2(n14743), .ZN(n6682) );
  OR2_X1 U9018 ( .A1(n12394), .A2(n13935), .ZN(n6683) );
  INV_X1 U9019 ( .A(n12672), .ZN(n7239) );
  INV_X1 U9020 ( .A(n13854), .ZN(n7448) );
  AND2_X1 U9021 ( .A1(n9709), .A2(n9708), .ZN(n6685) );
  AND2_X1 U9022 ( .A1(n15537), .A2(n7296), .ZN(n6686) );
  INV_X1 U9023 ( .A(n14770), .ZN(n7714) );
  AND2_X1 U9024 ( .A1(n13822), .A2(n13755), .ZN(n7447) );
  AND2_X1 U9025 ( .A1(n6683), .A2(n7763), .ZN(n6687) );
  NAND3_X1 U9026 ( .A1(n6966), .A2(n7338), .A3(n6796), .ZN(n6688) );
  AND2_X1 U9027 ( .A1(n6759), .A2(n7080), .ZN(n6689) );
  NAND2_X1 U9028 ( .A1(n9843), .A2(n9844), .ZN(n12982) );
  NAND2_X1 U9029 ( .A1(n11941), .A2(n11940), .ZN(n6690) );
  AND2_X1 U9030 ( .A1(n7595), .A2(n9737), .ZN(n6691) );
  AND2_X1 U9031 ( .A1(n6864), .A2(n6758), .ZN(n6692) );
  AND2_X1 U9032 ( .A1(n14091), .A2(n13921), .ZN(n6693) );
  OR2_X1 U9033 ( .A1(n8827), .A2(n8826), .ZN(n6694) );
  AND2_X1 U9034 ( .A1(n7714), .A2(n7354), .ZN(n6695) );
  AND2_X1 U9035 ( .A1(n7014), .A2(n12621), .ZN(n6696) );
  INV_X1 U9036 ( .A(n7599), .ZN(n7140) );
  NAND2_X1 U9037 ( .A1(n7603), .A2(n9714), .ZN(n7599) );
  INV_X1 U9038 ( .A(n10703), .ZN(n11209) );
  OR2_X1 U9039 ( .A1(n7936), .A2(n7935), .ZN(n10703) );
  AND2_X1 U9040 ( .A1(n8689), .A2(n8663), .ZN(n8664) );
  INV_X1 U9041 ( .A(n8664), .ZN(n7195) );
  INV_X1 U9042 ( .A(n7280), .ZN(n7279) );
  AND2_X1 U9043 ( .A1(n6686), .A2(n7295), .ZN(n6697) );
  NAND2_X1 U9044 ( .A1(n6813), .A2(n7808), .ZN(n6698) );
  OR2_X1 U9045 ( .A1(n7073), .A2(n8824), .ZN(n6699) );
  AND2_X1 U9046 ( .A1(n7789), .A2(n7794), .ZN(n6700) );
  AOI22_X1 U9047 ( .A1(n10409), .A2(n6680), .B1(n9124), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n14373) );
  INV_X1 U9048 ( .A(n14373), .ZN(n14050) );
  OR2_X1 U9049 ( .A1(n6972), .A2(n7402), .ZN(n6701) );
  NOR2_X1 U9050 ( .A1(n14965), .A2(n7689), .ZN(n7688) );
  AND2_X1 U9051 ( .A1(n8129), .A2(n7818), .ZN(n6702) );
  INV_X1 U9052 ( .A(n12242), .ZN(n7349) );
  AND2_X1 U9053 ( .A1(n7152), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n6703) );
  OR2_X2 U9054 ( .A1(n9108), .A2(n10957), .ZN(n8582) );
  INV_X1 U9055 ( .A(n14864), .ZN(n7705) );
  INV_X2 U9056 ( .A(n8405), .ZN(n9919) );
  AND4_X1 U9057 ( .A1(n7370), .A2(n7770), .A3(n7434), .A4(n7369), .ZN(n7918)
         );
  INV_X1 U9058 ( .A(n10920), .ZN(n7504) );
  INV_X1 U9059 ( .A(n15562), .ZN(n7592) );
  INV_X2 U9060 ( .A(n8643), .ZN(n8596) );
  AND2_X1 U9061 ( .A1(n7496), .A2(n7249), .ZN(n6704) );
  AND2_X1 U9062 ( .A1(n12763), .A2(n12758), .ZN(n6705) );
  NOR2_X1 U9063 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n10614) );
  NAND2_X1 U9064 ( .A1(n14843), .A2(n7365), .ZN(n14840) );
  NAND2_X1 U9065 ( .A1(n7245), .A2(n6704), .ZN(n14463) );
  OR2_X1 U9066 ( .A1(n14186), .A2(n14394), .ZN(n6706) );
  AND2_X1 U9067 ( .A1(n7500), .A2(n6705), .ZN(n6707) );
  AND2_X1 U9068 ( .A1(n14905), .A2(n7299), .ZN(n6708) );
  XNOR2_X1 U9069 ( .A(n14802), .B(n14764), .ZN(n14794) );
  INV_X1 U9070 ( .A(n14794), .ZN(n7711) );
  AND2_X1 U9071 ( .A1(n12561), .A2(n12560), .ZN(n6709) );
  INV_X1 U9072 ( .A(n13094), .ZN(n13548) );
  AND2_X1 U9073 ( .A1(n13214), .A2(n7318), .ZN(n6710) );
  AOI21_X1 U9074 ( .B1(n7895), .B2(n7164), .A(n7162), .ZN(n10648) );
  AND2_X1 U9075 ( .A1(n7732), .A2(n7070), .ZN(n6711) );
  XNOR2_X1 U9076 ( .A(n11754), .B(n11759), .ZN(n11647) );
  INV_X1 U9077 ( .A(n11647), .ZN(n7517) );
  AND2_X1 U9078 ( .A1(n7918), .A2(n7771), .ZN(n8009) );
  AND2_X1 U9079 ( .A1(n13148), .A2(n13147), .ZN(n6712) );
  OR2_X1 U9080 ( .A1(n9963), .A2(n7504), .ZN(n6713) );
  OR2_X1 U9081 ( .A1(n8553), .A2(n8552), .ZN(n6714) );
  OR2_X1 U9082 ( .A1(n10404), .A2(n7674), .ZN(n6715) );
  AND2_X1 U9083 ( .A1(n14353), .A2(n13840), .ZN(n6716) );
  OR2_X1 U9084 ( .A1(n12425), .A2(n12412), .ZN(n6717) );
  OR2_X1 U9085 ( .A1(n13499), .A2(n13482), .ZN(n6718) );
  INV_X1 U9086 ( .A(n7552), .ZN(n7551) );
  OAI21_X1 U9087 ( .B1(n7973), .B2(n7553), .A(n7994), .ZN(n7552) );
  OR2_X1 U9088 ( .A1(n7076), .A2(n8803), .ZN(n6719) );
  INV_X1 U9089 ( .A(n9737), .ZN(n9738) );
  OR2_X1 U9090 ( .A1(n8087), .A2(n7778), .ZN(n6720) );
  NAND2_X2 U9091 ( .A1(n10760), .A2(n9919), .ZN(n8469) );
  AND2_X1 U9092 ( .A1(n8207), .A2(n13223), .ZN(n6721) );
  AND2_X1 U9093 ( .A1(n11754), .A2(n13940), .ZN(n6722) );
  INV_X1 U9094 ( .A(n14072), .ZN(n14070) );
  AND2_X1 U9095 ( .A1(n9736), .A2(n9174), .ZN(n14072) );
  INV_X1 U9096 ( .A(n9735), .ZN(n7598) );
  AND2_X1 U9097 ( .A1(n14072), .A2(n14073), .ZN(n9735) );
  INV_X1 U9098 ( .A(n14436), .ZN(n7492) );
  OR2_X1 U9099 ( .A1(n13019), .A2(n13020), .ZN(n6723) );
  NAND2_X1 U9100 ( .A1(n8781), .A2(SI_14_), .ZN(n6724) );
  OR2_X1 U9101 ( .A1(n15167), .A2(n13051), .ZN(n6725) );
  AND2_X1 U9102 ( .A1(n13148), .A2(n12458), .ZN(n6726) );
  NAND2_X1 U9103 ( .A1(n10355), .A2(n10354), .ZN(n14762) );
  INV_X1 U9104 ( .A(n10722), .ZN(n7506) );
  OR3_X1 U9105 ( .A1(n9190), .A2(n9153), .A3(n9152), .ZN(n6727) );
  INV_X1 U9106 ( .A(n12301), .ZN(n12466) );
  AND2_X1 U9107 ( .A1(n7371), .A2(n9844), .ZN(n6728) );
  NOR2_X1 U9108 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n8391) );
  INV_X1 U9109 ( .A(n10375), .ZN(n7583) );
  NAND2_X1 U9110 ( .A1(n10216), .A2(n9897), .ZN(n10495) );
  AND2_X1 U9111 ( .A1(n12394), .A2(n13935), .ZN(n6729) );
  AND2_X1 U9112 ( .A1(n6995), .A2(n6994), .ZN(n6730) );
  OR2_X1 U9113 ( .A1(n8230), .A2(n15183), .ZN(n6731) );
  NAND2_X1 U9114 ( .A1(n13759), .A2(n13758), .ZN(n6732) );
  INV_X1 U9115 ( .A(n14911), .ZN(n15046) );
  NOR2_X1 U9116 ( .A1(n15064), .A2(n14705), .ZN(n6733) );
  NAND2_X1 U9117 ( .A1(n15146), .A2(n13320), .ZN(n6734) );
  NOR2_X1 U9118 ( .A1(n13224), .A2(n12868), .ZN(n6735) );
  AND2_X1 U9119 ( .A1(n7373), .A2(n7376), .ZN(n6736) );
  NAND2_X1 U9120 ( .A1(n8717), .A2(n8716), .ZN(n12191) );
  NAND2_X1 U9121 ( .A1(n10317), .A2(n10316), .ZN(n15024) );
  NAND2_X1 U9122 ( .A1(n9960), .A2(n9961), .ZN(n9977) );
  NAND2_X1 U9123 ( .A1(n10492), .A2(n9898), .ZN(n10497) );
  AND2_X1 U9124 ( .A1(n12526), .A2(n12466), .ZN(n6737) );
  AND2_X1 U9125 ( .A1(n7513), .A2(n9680), .ZN(n6738) );
  AND2_X1 U9126 ( .A1(n8895), .A2(n8894), .ZN(n6739) );
  NOR2_X1 U9127 ( .A1(n13466), .A2(n9848), .ZN(n6740) );
  INV_X1 U9128 ( .A(n11125), .ZN(n15662) );
  INV_X1 U9129 ( .A(n7514), .ZN(n7513) );
  NOR2_X1 U9130 ( .A1(n14385), .A2(n13764), .ZN(n7514) );
  OR2_X1 U9131 ( .A1(n13281), .A2(n13267), .ZN(n6741) );
  INV_X1 U9132 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7738) );
  INV_X1 U9133 ( .A(n12399), .ZN(n7455) );
  INV_X1 U9134 ( .A(n7186), .ZN(n8407) );
  OAI211_X1 U9135 ( .C1(n8405), .C2(P2_DATAO_REG_0__SCAN_IN), .A(SI_0_), .B(
        n7187), .ZN(n7186) );
  OR2_X1 U9136 ( .A1(n11315), .A2(n10621), .ZN(n6742) );
  AND2_X1 U9137 ( .A1(n13010), .A2(n11520), .ZN(n6743) );
  AND2_X1 U9138 ( .A1(n7063), .A2(n8583), .ZN(n6744) );
  AND2_X1 U9139 ( .A1(n14084), .A2(n9735), .ZN(n6745) );
  AND2_X1 U9140 ( .A1(n7083), .A2(n8920), .ZN(n6746) );
  INV_X1 U9141 ( .A(n9714), .ZN(n7602) );
  AND2_X1 U9142 ( .A1(n7498), .A2(n12768), .ZN(n6747) );
  AND2_X1 U9143 ( .A1(n12424), .A2(n12423), .ZN(n6748) );
  INV_X1 U9144 ( .A(n10319), .ZN(n7574) );
  AND2_X1 U9145 ( .A1(n13214), .A2(n6983), .ZN(n6749) );
  INV_X1 U9146 ( .A(n10117), .ZN(n7571) );
  INV_X1 U9147 ( .A(n10347), .ZN(n7577) );
  AND2_X1 U9148 ( .A1(n7088), .A2(n7090), .ZN(n6750) );
  AND2_X1 U9149 ( .A1(n9144), .A2(n9094), .ZN(n6751) );
  NAND2_X1 U9150 ( .A1(n12544), .A2(n12543), .ZN(n6752) );
  OR2_X1 U9151 ( .A1(n8657), .A2(n8656), .ZN(n6753) );
  INV_X1 U9152 ( .A(n7688), .ZN(n7687) );
  AND2_X1 U9153 ( .A1(n9128), .A2(n9127), .ZN(n14291) );
  INV_X1 U9154 ( .A(n14291), .ZN(n9775) );
  AND2_X1 U9155 ( .A1(n13086), .A2(n13496), .ZN(n6754) );
  AND2_X1 U9156 ( .A1(n15371), .A2(n15359), .ZN(n6755) );
  AND2_X1 U9157 ( .A1(n7086), .A2(n7085), .ZN(n6756) );
  INV_X1 U9158 ( .A(n7135), .ZN(n7134) );
  NOR2_X1 U9159 ( .A1(n6716), .A2(n7136), .ZN(n7135) );
  AND2_X1 U9160 ( .A1(n13187), .A2(n13186), .ZN(n13577) );
  INV_X1 U9161 ( .A(n13577), .ZN(n8240) );
  INV_X1 U9162 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8103) );
  INV_X1 U9163 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9915) );
  OR2_X1 U9164 ( .A1(n8499), .A2(n8498), .ZN(n6757) );
  AND2_X1 U9165 ( .A1(n6725), .A2(n6981), .ZN(n6758) );
  OR2_X1 U9166 ( .A1(n8993), .A2(n8995), .ZN(n6759) );
  NOR2_X1 U9167 ( .A1(n15543), .A2(n14554), .ZN(n6760) );
  NOR2_X1 U9168 ( .A1(n15052), .A2(n14709), .ZN(n6761) );
  NOR2_X1 U9169 ( .A1(n12736), .A2(n12735), .ZN(n6762) );
  NOR2_X1 U9170 ( .A1(n14353), .A2(n13930), .ZN(n6763) );
  NOR2_X1 U9171 ( .A1(n14394), .A2(n9727), .ZN(n6764) );
  NOR2_X1 U9172 ( .A1(n12687), .A2(n15333), .ZN(n6765) );
  AND2_X1 U9173 ( .A1(n13225), .A2(n8340), .ZN(n13407) );
  AND2_X1 U9174 ( .A1(n13667), .A2(n13519), .ZN(n6766) );
  AND2_X1 U9175 ( .A1(n13499), .A2(n13482), .ZN(n6767) );
  AND3_X1 U9176 ( .A1(n7871), .A2(n7869), .A3(n7868), .ZN(n6768) );
  NOR2_X1 U9177 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8474) );
  NOR2_X1 U9178 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n8388) );
  NAND2_X1 U9179 ( .A1(n13736), .A2(n13741), .ZN(n6769) );
  NOR2_X1 U9180 ( .A1(n9858), .A2(n7388), .ZN(n6770) );
  AND4_X1 U9181 ( .A1(n6839), .A2(n6838), .A3(n7783), .A4(n6968), .ZN(n6771)
         );
  OR2_X1 U9182 ( .A1(n10318), .A2(n7574), .ZN(n6772) );
  AND2_X1 U9183 ( .A1(n8628), .A2(n8627), .ZN(n6773) );
  INV_X1 U9184 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n6978) );
  INV_X1 U9185 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8118) );
  INV_X1 U9186 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7833) );
  INV_X1 U9187 ( .A(n7141), .ZN(n7132) );
  OR2_X1 U9188 ( .A1(n7599), .A2(n15280), .ZN(n7141) );
  OR2_X1 U9189 ( .A1(n7438), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n6774) );
  AND2_X1 U9190 ( .A1(n8728), .A2(n8727), .ZN(n6775) );
  NAND2_X1 U9191 ( .A1(n7401), .A2(n7781), .ZN(n6776) );
  INV_X1 U9192 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9917) );
  NAND2_X1 U9193 ( .A1(n7716), .A2(n9915), .ZN(n6777) );
  AND2_X1 U9194 ( .A1(n6902), .A2(n13205), .ZN(n6778) );
  NOR2_X1 U9195 ( .A1(n14995), .A2(n14789), .ZN(n6779) );
  AND2_X1 U9196 ( .A1(n8711), .A2(n10724), .ZN(n6780) );
  AND2_X1 U9197 ( .A1(n12693), .A2(n10200), .ZN(n12623) );
  INV_X1 U9198 ( .A(n12623), .ZN(n7014) );
  INV_X1 U9199 ( .A(n7283), .ZN(n7281) );
  AND2_X1 U9200 ( .A1(n10706), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7283) );
  OR2_X1 U9201 ( .A1(n8239), .A2(n7637), .ZN(n6781) );
  AND2_X1 U9202 ( .A1(n7804), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n6782) );
  AND2_X1 U9203 ( .A1(n14341), .A2(n13928), .ZN(n6783) );
  INV_X1 U9204 ( .A(n14749), .ZN(n7696) );
  NOR2_X1 U9205 ( .A1(n7731), .A2(n8994), .ZN(n6784) );
  OR2_X1 U9206 ( .A1(n7762), .A2(n6729), .ZN(n6785) );
  INV_X1 U9207 ( .A(n7142), .ZN(n7139) );
  INV_X1 U9208 ( .A(n7611), .ZN(n7610) );
  NAND2_X1 U9209 ( .A1(n9709), .A2(n7612), .ZN(n7611) );
  INV_X1 U9210 ( .A(n7098), .ZN(n7097) );
  NAND2_X1 U9211 ( .A1(n7099), .A2(n8730), .ZN(n7098) );
  OR2_X1 U9212 ( .A1(n14700), .A2(n15326), .ZN(n14741) );
  INV_X1 U9213 ( .A(n14741), .ZN(n7689) );
  AND2_X1 U9214 ( .A1(n7027), .A2(n7023), .ZN(n6786) );
  INV_X1 U9215 ( .A(n9677), .ZN(n14139) );
  AND2_X1 U9216 ( .A1(n6927), .A2(n8377), .ZN(n6787) );
  INV_X2 U9217 ( .A(n10069), .ZN(n9970) );
  OAI21_X1 U9218 ( .B1(n8665), .B2(n7196), .A(n7194), .ZN(n8732) );
  AND2_X1 U9219 ( .A1(n12245), .A2(n14557), .ZN(n6788) );
  AND2_X1 U9220 ( .A1(n7293), .A2(n7294), .ZN(n6789) );
  INV_X1 U9221 ( .A(n14884), .ZN(n15033) );
  NAND2_X1 U9222 ( .A1(n15106), .A2(n9963), .ZN(n14884) );
  AND2_X1 U9223 ( .A1(n8604), .A2(n8603), .ZN(n6790) );
  AND2_X1 U9224 ( .A1(n7472), .A2(n14377), .ZN(n6791) );
  INV_X1 U9225 ( .A(n9734), .ZN(n7126) );
  NAND2_X1 U9226 ( .A1(n15204), .A2(n15209), .ZN(n6792) );
  AND2_X1 U9227 ( .A1(n8437), .A2(n7663), .ZN(n6793) );
  INV_X1 U9228 ( .A(n12182), .ZN(n7058) );
  AND2_X1 U9229 ( .A1(n7075), .A2(n8826), .ZN(n6794) );
  AND2_X1 U9230 ( .A1(n7275), .A2(n7274), .ZN(n6795) );
  AND2_X1 U9231 ( .A1(n7771), .A2(n7783), .ZN(n6796) );
  AND2_X1 U9232 ( .A1(n9927), .A2(n7567), .ZN(n6797) );
  OR2_X1 U9233 ( .A1(n7577), .A2(n10346), .ZN(n6798) );
  OR2_X1 U9234 ( .A1(n10151), .A2(n10149), .ZN(n6799) );
  AND2_X1 U9235 ( .A1(n12923), .A2(n9782), .ZN(n12953) );
  OR2_X1 U9236 ( .A1(n10083), .A2(n10081), .ZN(n6800) );
  OR2_X1 U9237 ( .A1(n7583), .A2(n10374), .ZN(n6801) );
  OR2_X1 U9238 ( .A1(n10048), .A2(n10050), .ZN(n6802) );
  OR2_X1 U9239 ( .A1(n8854), .A2(n8856), .ZN(n6803) );
  AND2_X1 U9240 ( .A1(n8805), .A2(n6724), .ZN(n6804) );
  NAND2_X1 U9241 ( .A1(n8780), .A2(n8779), .ZN(n6805) );
  AND2_X1 U9242 ( .A1(n7630), .A2(n6718), .ZN(n6806) );
  OAI21_X1 U9243 ( .B1(n9817), .B2(n7396), .A(n9816), .ZN(n7395) );
  AND2_X1 U9244 ( .A1(n7094), .A2(n7093), .ZN(n6807) );
  NAND2_X1 U9245 ( .A1(n10614), .A2(n7770), .ZN(n7895) );
  INV_X1 U9246 ( .A(n7523), .ZN(n7522) );
  NAND2_X1 U9247 ( .A1(n6785), .A2(n6683), .ZN(n7523) );
  NAND2_X1 U9248 ( .A1(n10148), .A2(n10147), .ZN(n12687) );
  OR2_X1 U9249 ( .A1(n7598), .A2(n7126), .ZN(n6808) );
  INV_X1 U9250 ( .A(n7111), .ZN(n7110) );
  NAND2_X1 U9251 ( .A1(n7112), .A2(n9730), .ZN(n7111) );
  INV_X1 U9252 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7113) );
  INV_X1 U9253 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n6968) );
  INV_X1 U9254 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7434) );
  OR2_X1 U9255 ( .A1(n7571), .A2(n10116), .ZN(n6809) );
  OR2_X1 U9256 ( .A1(n7492), .A2(n7490), .ZN(n6810) );
  INV_X1 U9257 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7165) );
  INV_X1 U9258 ( .A(n14144), .ZN(n7008) );
  INV_X1 U9259 ( .A(n10528), .ZN(n12819) );
  XOR2_X1 U9260 ( .A(n14159), .B(n13806), .Z(n6811) );
  INV_X1 U9261 ( .A(n12043), .ZN(n7526) );
  INV_X1 U9262 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n8440) );
  INV_X1 U9263 ( .A(n9747), .ZN(n7046) );
  NAND2_X1 U9264 ( .A1(n12911), .A2(n9813), .ZN(n12876) );
  NAND2_X1 U9265 ( .A1(n6895), .A2(n14706), .ZN(n14933) );
  NAND2_X1 U9266 ( .A1(n7258), .A2(n7257), .ZN(n12727) );
  AND2_X1 U9267 ( .A1(n7056), .A2(n7449), .ZN(n6812) );
  INV_X1 U9268 ( .A(n7289), .ZN(n12697) );
  NOR2_X1 U9269 ( .A1(n12645), .A2(n15386), .ZN(n7289) );
  INV_X1 U9270 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6986) );
  NAND2_X1 U9271 ( .A1(n14702), .A2(n14701), .ZN(n14964) );
  NAND2_X1 U9272 ( .A1(n15338), .A2(n12731), .ZN(n15302) );
  XOR2_X1 U9273 ( .A(n11178), .B(P1_DATAO_REG_12__SCAN_IN), .Z(n6813) );
  INV_X1 U9274 ( .A(n8975), .ZN(n7081) );
  NAND3_X1 U9275 ( .A1(n6926), .A2(n6927), .A3(n6925), .ZN(n6814) );
  INV_X1 U9276 ( .A(n7467), .ZN(n14232) );
  AND2_X1 U9277 ( .A1(n9806), .A2(n9805), .ZN(n6815) );
  INV_X1 U9278 ( .A(n13196), .ZN(n13525) );
  AND2_X1 U9279 ( .A1(n13197), .A2(n13198), .ZN(n13196) );
  NAND2_X1 U9280 ( .A1(n7695), .A2(n14749), .ZN(n6816) );
  NAND2_X1 U9281 ( .A1(n15389), .A2(n12690), .ZN(n12691) );
  INV_X1 U9282 ( .A(n12691), .ZN(n7364) );
  AND2_X1 U9283 ( .A1(n11973), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n6817) );
  INV_X1 U9284 ( .A(n8087), .ZN(n7641) );
  INV_X1 U9285 ( .A(n13182), .ZN(n13186) );
  AND2_X1 U9286 ( .A1(n13681), .A2(n12947), .ZN(n13182) );
  AND2_X1 U9287 ( .A1(n7525), .A2(n7524), .ZN(n6818) );
  OR2_X1 U9288 ( .A1(n8781), .A2(SI_14_), .ZN(n6819) );
  OR2_X1 U9289 ( .A1(n7812), .A2(n7213), .ZN(n6820) );
  AND2_X1 U9290 ( .A1(n13542), .A2(n8243), .ZN(n6821) );
  OR2_X1 U9291 ( .A1(n7730), .A2(n8855), .ZN(n6822) );
  AND2_X1 U9292 ( .A1(n7759), .A2(n7765), .ZN(n6823) );
  AND2_X1 U9293 ( .A1(n14250), .A2(n9669), .ZN(n6824) );
  INV_X1 U9294 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10698) );
  INV_X1 U9295 ( .A(n7178), .ZN(n7177) );
  NAND2_X1 U9296 ( .A1(n8958), .A2(n7180), .ZN(n7178) );
  INV_X2 U9297 ( .A(n15801), .ZN(n15822) );
  AND2_X1 U9298 ( .A1(n11825), .A2(n14975), .ZN(n15495) );
  INV_X1 U9299 ( .A(n13144), .ZN(n6953) );
  INV_X1 U9300 ( .A(n12486), .ZN(n9666) );
  INV_X1 U9301 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7261) );
  NAND2_X1 U9302 ( .A1(n8742), .A2(n8741), .ZN(n12394) );
  INV_X1 U9303 ( .A(n12394), .ZN(n7473) );
  NAND2_X1 U9304 ( .A1(n8281), .A2(n13707), .ZN(n8284) );
  INV_X1 U9305 ( .A(n14345), .ZN(n7466) );
  NAND2_X1 U9306 ( .A1(n8697), .A2(n8696), .ZN(n12105) );
  INV_X1 U9307 ( .A(n12105), .ZN(n7476) );
  OAI22_X1 U9308 ( .A1(n8284), .A2(P3_D_REG_0__SCAN_IN), .B1(n13707), .B2(
        n12496), .ZN(n9778) );
  AND2_X1 U9309 ( .A1(n11807), .A2(n7475), .ZN(n6825) );
  AND2_X1 U9310 ( .A1(n6697), .A2(n12310), .ZN(n6826) );
  NAND2_X1 U9311 ( .A1(n6937), .A2(n7515), .ZN(n11805) );
  NAND2_X1 U9312 ( .A1(n6889), .A2(n12528), .ZN(n12617) );
  NAND2_X1 U9313 ( .A1(n12054), .A2(n12053), .ZN(n12243) );
  NAND2_X1 U9314 ( .A1(n7353), .A2(n12468), .ZN(n12527) );
  AND2_X1 U9315 ( .A1(n7817), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6827) );
  NAND3_X1 U9316 ( .A1(n7584), .A2(n10012), .A3(n7260), .ZN(n6828) );
  INV_X1 U9317 ( .A(n15124), .ZN(n13281) );
  INV_X1 U9318 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7059) );
  AND2_X1 U9319 ( .A1(n6827), .A2(n12392), .ZN(n6829) );
  NAND2_X1 U9320 ( .A1(n12628), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6830) );
  AND2_X1 U9321 ( .A1(n12559), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6831) );
  INV_X1 U9322 ( .A(n8542), .ZN(n8643) );
  AND2_X1 U9323 ( .A1(n7539), .A2(n7818), .ZN(n6832) );
  INV_X1 U9324 ( .A(n11534), .ZN(n7469) );
  XNOR2_X1 U9325 ( .A(n8073), .B(n8072), .ZN(n15146) );
  NAND4_X1 U9326 ( .A1(n7890), .A2(n7889), .A3(n7888), .A4(n7887), .ZN(n15808)
         );
  INV_X1 U9327 ( .A(n15808), .ZN(n7377) );
  AND2_X1 U9328 ( .A1(n12716), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6833) );
  NAND2_X1 U9329 ( .A1(n9784), .A2(n15790), .ZN(n9788) );
  AND2_X2 U9330 ( .A1(n10896), .A2(n10895), .ZN(n15731) );
  NAND2_X1 U9331 ( .A1(n11611), .A2(n10535), .ZN(n11378) );
  INV_X1 U9332 ( .A(n15543), .ZN(n7296) );
  NAND2_X1 U9333 ( .A1(n10130), .A2(n10129), .ZN(n15403) );
  INV_X1 U9334 ( .A(n15403), .ZN(n7295) );
  NAND2_X1 U9335 ( .A1(n7779), .A2(n6720), .ZN(n11663) );
  INV_X1 U9336 ( .A(n11663), .ZN(n6971) );
  XNOR2_X1 U9337 ( .A(n10533), .B(n10532), .ZN(n11610) );
  INV_X1 U9338 ( .A(n15501), .ZN(n7292) );
  AND2_X1 U9339 ( .A1(n7156), .A2(n13361), .ZN(n6834) );
  AND2_X1 U9340 ( .A1(n13319), .A2(n13308), .ZN(n6835) );
  AND2_X1 U9341 ( .A1(n10957), .A2(n9747), .ZN(n6836) );
  INV_X1 U9342 ( .A(SI_22_), .ZN(n7180) );
  INV_X1 U9343 ( .A(n7229), .ZN(n7228) );
  NAND2_X1 U9344 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n12861), .ZN(n7229) );
  NAND2_X1 U9345 ( .A1(n9901), .A2(n9902), .ZN(n15085) );
  NOR2_X1 U9346 ( .A1(n8395), .A2(n7737), .ZN(n14405) );
  INV_X1 U9347 ( .A(SI_2_), .ZN(n7663) );
  INV_X1 U9348 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n11008) );
  INV_X1 U9349 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7312) );
  XNOR2_X1 U9350 ( .A(n13299), .B(n15146), .ZN(n15143) );
  NAND2_X1 U9351 ( .A1(n7270), .A2(n15146), .ZN(n7269) );
  NOR2_X1 U9352 ( .A1(n11475), .A2(n15807), .ZN(n11260) );
  NAND2_X1 U9353 ( .A1(n6768), .A2(n7870), .ZN(n15807) );
  AND3_X2 U9354 ( .A1(n7876), .A2(n7874), .A3(n7875), .ZN(n11475) );
  NAND2_X1 U9355 ( .A1(n11631), .A2(n13062), .ZN(n11633) );
  NAND2_X1 U9356 ( .A1(n11777), .A2(n13124), .ZN(n6837) );
  NAND2_X2 U9357 ( .A1(n8268), .A2(n9919), .ZN(n13050) );
  XNOR2_X2 U9358 ( .A(n7832), .B(n7831), .ZN(n8266) );
  NAND2_X1 U9359 ( .A1(n11960), .A2(n13060), .ZN(n11959) );
  OAI21_X2 U9360 ( .B1(n8083), .B2(n8240), .A(n6900), .ZN(n13565) );
  NAND3_X1 U9361 ( .A1(n6850), .A2(n6847), .A3(n6846), .ZN(n6845) );
  AOI21_X1 U9362 ( .B1(n6851), .B2(n13172), .A(n15176), .ZN(n13178) );
  NAND2_X1 U9363 ( .A1(n6854), .A2(n6853), .ZN(n6852) );
  NAND2_X1 U9364 ( .A1(n6855), .A2(n6792), .ZN(n6854) );
  NAND2_X1 U9365 ( .A1(n6856), .A2(n13164), .ZN(n6855) );
  OAI21_X1 U9366 ( .B1(n13161), .B2(n13160), .A(n13159), .ZN(n6856) );
  NAND2_X1 U9367 ( .A1(n6857), .A2(n13201), .ZN(n13206) );
  OR2_X1 U9368 ( .A1(n6859), .A2(n6858), .ZN(n6857) );
  AOI21_X1 U9369 ( .B1(n6982), .B2(n13195), .A(n6860), .ZN(n6859) );
  INV_X1 U9370 ( .A(n13194), .ZN(n6861) );
  AOI21_X1 U9371 ( .B1(n13217), .B2(n6863), .A(n6862), .ZN(n6980) );
  NAND2_X1 U9372 ( .A1(n6984), .A2(n6749), .ZN(n13217) );
  OAI21_X1 U9373 ( .B1(n6868), .B2(n13227), .A(n6865), .ZN(n6864) );
  NOR2_X1 U9374 ( .A1(n13229), .A2(n13228), .ZN(n6866) );
  INV_X1 U9375 ( .A(n13230), .ZN(n6867) );
  NAND2_X1 U9376 ( .A1(n6869), .A2(n13114), .ZN(n13119) );
  NAND2_X1 U9377 ( .A1(n6870), .A2(n13112), .ZN(n6869) );
  NAND2_X1 U9378 ( .A1(n6871), .A2(n13110), .ZN(n6870) );
  NAND3_X1 U9379 ( .A1(n13106), .A2(n13107), .A3(n15785), .ZN(n6871) );
  INV_X1 U9380 ( .A(n15423), .ZN(n6874) );
  NAND2_X1 U9381 ( .A1(n15420), .A2(n15418), .ZN(n15424) );
  NAND2_X1 U9382 ( .A1(n6876), .A2(n15439), .ZN(n15139) );
  NAND2_X1 U9383 ( .A1(n15440), .A2(n15441), .ZN(n15439) );
  NAND2_X1 U9384 ( .A1(n15437), .A2(n15436), .ZN(n15435) );
  XNOR2_X1 U9385 ( .A(n7305), .B(n6878), .ZN(n9268) );
  NAND2_X1 U9386 ( .A1(n14372), .A2(n6879), .ZN(P2_U3498) );
  NOR2_X2 U9388 ( .A1(n6706), .A2(n14159), .ZN(n7465) );
  NAND3_X1 U9389 ( .A1(n7836), .A2(n7835), .A3(n7643), .ZN(n6880) );
  NAND3_X1 U9390 ( .A1(n7837), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n6881) );
  NAND2_X1 U9391 ( .A1(n8559), .A2(n8558), .ZN(n8564) );
  OAI211_X1 U9392 ( .C1(n8507), .C2(n7184), .A(n8532), .B(n6884), .ZN(n8559)
         );
  NAND2_X1 U9393 ( .A1(n8503), .A2(n6885), .ZN(n6884) );
  NAND2_X1 U9394 ( .A1(n9746), .A2(n6791), .ZN(n14056) );
  NOR2_X2 U9395 ( .A1(n14104), .A2(n14091), .ZN(n9746) );
  NAND3_X1 U9396 ( .A1(n7840), .A2(n7839), .A3(P2_DATAO_REG_1__SCAN_IN), .ZN(
        n6887) );
  NAND2_X1 U9397 ( .A1(n8404), .A2(SI_1_), .ZN(n8437) );
  NAND2_X1 U9398 ( .A1(n12617), .A2(n12616), .ZN(n12619) );
  NAND2_X1 U9399 ( .A1(n12591), .A2(n12599), .ZN(n6889) );
  NAND2_X1 U9400 ( .A1(n7350), .A2(n7351), .ZN(n12591) );
  INV_X1 U9401 ( .A(n14865), .ZN(n14716) );
  NAND2_X1 U9402 ( .A1(n14876), .A2(n14878), .ZN(n6890) );
  NOR2_X2 U9403 ( .A1(n9979), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n10012) );
  NAND3_X1 U9404 ( .A1(n6892), .A2(n9897), .A3(n6891), .ZN(n7368) );
  OAI21_X2 U9405 ( .B1(n14933), .B2(n14708), .A(n14707), .ZN(n14919) );
  NAND2_X2 U9406 ( .A1(n12622), .A2(n6696), .ZN(n15389) );
  NAND2_X2 U9407 ( .A1(n14808), .A2(n14807), .ZN(n14806) );
  OAI21_X1 U9408 ( .B1(n15177), .B2(n13175), .A(n13173), .ZN(n12635) );
  NOR2_X1 U9409 ( .A1(n13144), .A2(n6712), .ZN(n6912) );
  NAND2_X1 U9410 ( .A1(n11633), .A2(n13127), .ZN(n11960) );
  NAND3_X1 U9411 ( .A1(n7332), .A2(n7640), .A3(n7846), .ZN(n13689) );
  NAND2_X1 U9412 ( .A1(n6914), .A2(n9648), .ZN(n11559) );
  XNOR2_X2 U9413 ( .A(n6915), .B(n13946), .ZN(n10889) );
  NAND2_X2 U9414 ( .A1(n14116), .A2(n9679), .ZN(n14103) );
  NAND3_X1 U9415 ( .A1(n6922), .A2(n6923), .A3(n6927), .ZN(n8395) );
  NAND2_X1 U9416 ( .A1(n6926), .A2(n6927), .ZN(n9197) );
  INV_X1 U9417 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6925) );
  INV_X1 U9418 ( .A(n8374), .ZN(n6927) );
  INV_X1 U9419 ( .A(n14249), .ZN(n6931) );
  NOR2_X1 U9420 ( .A1(n9654), .A2(n6934), .ZN(n6933) );
  NAND2_X1 U9421 ( .A1(n11385), .A2(n11388), .ZN(n9657) );
  NAND2_X1 U9422 ( .A1(n6938), .A2(n11523), .ZN(n6937) );
  NAND2_X1 U9423 ( .A1(n11805), .A2(n11809), .ZN(n6940) );
  NAND2_X2 U9424 ( .A1(n9203), .A2(n10767), .ZN(n10760) );
  NAND2_X1 U9425 ( .A1(n11539), .A2(n13116), .ZN(n11540) );
  NAND2_X1 U9426 ( .A1(n11792), .A2(n9793), .ZN(n11975) );
  NAND2_X1 U9427 ( .A1(n11793), .A2(n11794), .ZN(n11792) );
  AND2_X1 U9428 ( .A1(n7374), .A2(n6736), .ZN(n11736) );
  NAND3_X1 U9429 ( .A1(n9788), .A2(n9786), .A3(n6959), .ZN(n7375) );
  NAND2_X1 U9430 ( .A1(n9787), .A2(n6960), .ZN(n6959) );
  NAND2_X1 U9431 ( .A1(n12862), .A2(n15805), .ZN(n6960) );
  NAND2_X1 U9432 ( .A1(n9830), .A2(n6961), .ZN(n12890) );
  NAND2_X1 U9433 ( .A1(n9846), .A2(n9845), .ZN(n12952) );
  NAND2_X1 U9434 ( .A1(n9846), .A2(n6963), .ZN(n12921) );
  NAND4_X1 U9435 ( .A1(n6966), .A2(n7338), .A3(n7771), .A4(n6965), .ZN(n8272)
         );
  NAND2_X1 U9436 ( .A1(n8273), .A2(n8297), .ZN(n8275) );
  NAND2_X1 U9437 ( .A1(n8273), .A2(n6969), .ZN(n8279) );
  NAND2_X1 U9438 ( .A1(n8273), .A2(n6967), .ZN(n6970) );
  NAND2_X1 U9439 ( .A1(n12926), .A2(n9855), .ZN(n13011) );
  NAND2_X1 U9440 ( .A1(n9840), .A2(n9839), .ZN(n9843) );
  NAND2_X1 U9441 ( .A1(n9849), .A2(n12922), .ZN(n9854) );
  NAND2_X1 U9442 ( .A1(n7375), .A2(n9788), .ZN(n7380) );
  NAND2_X1 U9443 ( .A1(n9843), .A2(n13507), .ZN(n7372) );
  NAND2_X1 U9444 ( .A1(n11627), .A2(n8222), .ZN(n11962) );
  NAND2_X1 U9445 ( .A1(n12319), .A2(n8226), .ZN(n15207) );
  INV_X1 U9446 ( .A(n11737), .ZN(n7373) );
  NAND2_X1 U9447 ( .A1(n7380), .A2(n7379), .ZN(n7374) );
  NAND2_X1 U9448 ( .A1(n13505), .A2(n8246), .ZN(n8248) );
  NAND2_X1 U9449 ( .A1(n11962), .A2(n13134), .ZN(n11961) );
  NAND2_X1 U9450 ( .A1(n11425), .A2(n6974), .ZN(n11429) );
  NAND2_X1 U9451 ( .A1(n12901), .A2(n9837), .ZN(n9842) );
  XNOR2_X1 U9452 ( .A(n13011), .B(n13012), .ZN(n13013) );
  NAND2_X1 U9453 ( .A1(n6979), .A2(n6977), .ZN(n8276) );
  NAND2_X1 U9454 ( .A1(n8274), .A2(P3_IR_REG_24__SCAN_IN), .ZN(n6979) );
  NAND2_X1 U9455 ( .A1(n13517), .A2(n13525), .ZN(n13516) );
  NAND2_X1 U9456 ( .A1(n8591), .A2(n8590), .ZN(n8609) );
  NAND2_X1 U9457 ( .A1(n8832), .A2(n8831), .ZN(n8858) );
  NAND2_X1 U9458 ( .A1(n8736), .A2(n8735), .ZN(n8764) );
  NAND2_X1 U9459 ( .A1(n7662), .A2(n8441), .ZN(n7661) );
  XNOR2_X1 U9460 ( .A(n8883), .B(n8882), .ZN(n12387) );
  NOR2_X1 U9461 ( .A1(n13410), .A2(n8341), .ZN(n8343) );
  OAI21_X1 U9462 ( .B1(n9061), .B2(n13710), .A(n9060), .ZN(n7166) );
  NAND2_X1 U9463 ( .A1(n9079), .A2(n7668), .ZN(n7667) );
  NAND2_X1 U9464 ( .A1(n8979), .A2(n7173), .ZN(n8998) );
  NAND2_X1 U9465 ( .A1(n7181), .A2(n8958), .ZN(n8978) );
  NAND3_X1 U9466 ( .A1(n7190), .A2(n14061), .A3(n14069), .ZN(n14287) );
  INV_X1 U9467 ( .A(n6980), .ZN(n7536) );
  MUX2_X1 U9468 ( .A(n13132), .B(n13131), .S(n13228), .Z(n13142) );
  NAND2_X1 U9469 ( .A1(n7338), .A2(n6771), .ZN(n7642) );
  OR2_X1 U9470 ( .A1(n11427), .A2(n12109), .ZN(n13123) );
  NAND3_X1 U9471 ( .A1(n13190), .A2(n13548), .A3(n13564), .ZN(n6982) );
  NAND2_X1 U9472 ( .A1(n13108), .A2(n13111), .ZN(n8214) );
  OR2_X1 U9473 ( .A1(n7847), .A2(n8010), .ZN(n7848) );
  INV_X1 U9474 ( .A(n11496), .ZN(n7379) );
  NAND3_X1 U9475 ( .A1(n7657), .A2(n8437), .A3(n8407), .ZN(n8438) );
  NAND2_X1 U9476 ( .A1(n7189), .A2(n10728), .ZN(n7657) );
  NAND2_X1 U9477 ( .A1(n14806), .A2(n7355), .ZN(n7015) );
  NAND3_X1 U9478 ( .A1(n7555), .A2(n6987), .A3(n10265), .ZN(n10274) );
  OAI21_X1 U9479 ( .B1(n14992), .B2(n15529), .A(n6789), .ZN(n15072) );
  NAND2_X1 U9480 ( .A1(n7419), .A2(n7418), .ZN(n11403) );
  NOR2_X1 U9481 ( .A1(n11203), .A2(n10657), .ZN(n11202) );
  NAND2_X1 U9482 ( .A1(n11056), .A2(n11057), .ZN(n11055) );
  NOR2_X1 U9483 ( .A1(n11291), .A2(n11290), .ZN(n11289) );
  INV_X1 U9484 ( .A(n14145), .ZN(n7009) );
  NAND2_X1 U9485 ( .A1(n7166), .A2(n9062), .ZN(n9079) );
  NAND2_X1 U9486 ( .A1(n6691), .A2(n6808), .ZN(n7120) );
  INV_X1 U9487 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7643) );
  NAND2_X1 U9488 ( .A1(n8978), .A2(SI_22_), .ZN(n8979) );
  NAND2_X1 U9489 ( .A1(n8998), .A2(n8997), .ZN(n9001) );
  NAND2_X1 U9490 ( .A1(n7193), .A2(n7191), .ZN(n8736) );
  NAND2_X1 U9491 ( .A1(n7653), .A2(n7650), .ZN(n9061) );
  NAND2_X1 U9492 ( .A1(n8765), .A2(n6819), .ZN(n7672) );
  NAND2_X1 U9493 ( .A1(n15109), .A2(n6996), .ZN(n15112) );
  NAND2_X1 U9494 ( .A1(n6998), .A2(n6997), .ZN(n6996) );
  INV_X1 U9495 ( .A(n15110), .ZN(n6997) );
  INV_X1 U9496 ( .A(n15111), .ZN(n6998) );
  OAI211_X1 U9497 ( .C1(n12874), .C2(n12875), .A(n7002), .B(n12873), .ZN(
        P3_U3160) );
  NAND2_X1 U9498 ( .A1(n12874), .A2(n7003), .ZN(n7002) );
  NAND2_X2 U9499 ( .A1(n9854), .A2(n12924), .ZN(n12926) );
  OR2_X1 U9500 ( .A1(n11009), .A2(n11239), .ZN(n11061) );
  NOR2_X2 U9501 ( .A1(n15151), .A2(n15152), .ZN(n15150) );
  NOR2_X2 U9502 ( .A1(n15741), .A2(n15740), .ZN(n15739) );
  NAND2_X1 U9503 ( .A1(n13396), .A2(n13395), .ZN(n7161) );
  AOI21_X1 U9504 ( .B1(n11157), .B2(n11156), .A(n11155), .ZN(n11212) );
  NAND2_X1 U9505 ( .A1(n7628), .A2(n7627), .ZN(n7624) );
  AOI21_X1 U9506 ( .B1(n14180), .B2(n14181), .A(n9673), .ZN(n14163) );
  NAND2_X1 U9507 ( .A1(n7013), .A2(n7010), .ZN(P3_U3180) );
  NAND2_X1 U9508 ( .A1(n13013), .A2(n13023), .ZN(n7013) );
  AND3_X2 U9509 ( .A1(n7290), .A2(n9965), .A3(n7291), .ZN(n15513) );
  NAND2_X1 U9510 ( .A1(n15499), .A2(n15500), .ZN(n11925) );
  NAND2_X2 U9511 ( .A1(n11913), .A2(n9986), .ZN(n15500) );
  NAND2_X1 U9512 ( .A1(n10492), .A2(n7715), .ZN(n7501) );
  NAND2_X1 U9513 ( .A1(n11763), .A2(n11758), .ZN(n7016) );
  INV_X1 U9514 ( .A(n13779), .ZN(n7018) );
  NAND2_X1 U9515 ( .A1(n11111), .A2(n11171), .ZN(n11177) );
  NAND2_X1 U9516 ( .A1(n7443), .A2(n6786), .ZN(n7019) );
  OAI211_X1 U9517 ( .C1(n7443), .C2(n7024), .A(n7019), .B(n7020), .ZN(n13814)
         );
  NAND2_X1 U9518 ( .A1(n7443), .A2(n7441), .ZN(n7026) );
  OAI21_X1 U9519 ( .B1(n7443), .B2(n7033), .A(n7441), .ZN(n13902) );
  NAND2_X1 U9520 ( .A1(n13851), .A2(n7038), .ZN(n7036) );
  OAI21_X2 U9521 ( .B1(n9684), .B2(n7045), .A(n7044), .ZN(n7043) );
  NOR2_X1 U9522 ( .A1(n7053), .A2(n6709), .ZN(n7047) );
  NOR2_X1 U9523 ( .A1(n7451), .A2(n7058), .ZN(n7057) );
  INV_X1 U9524 ( .A(n7054), .ZN(n7055) );
  NAND2_X1 U9525 ( .A1(n7053), .A2(n7052), .ZN(n7054) );
  NAND3_X1 U9526 ( .A1(n7051), .A2(n7050), .A3(n12182), .ZN(n7049) );
  INV_X1 U9527 ( .A(n6709), .ZN(n7051) );
  NAND2_X1 U9528 ( .A1(n7056), .A2(n7055), .ZN(n12562) );
  NAND4_X1 U9529 ( .A1(n7062), .A2(n7061), .A3(n7060), .A4(n7059), .ZN(n8836)
         );
  NAND4_X1 U9530 ( .A1(n7065), .A2(n8474), .A3(n7067), .A4(n7064), .ZN(n8374)
         );
  NAND2_X1 U9531 ( .A1(n8607), .A2(n6790), .ZN(n7070) );
  NAND2_X1 U9532 ( .A1(n7069), .A2(n7735), .ZN(n8657) );
  INV_X1 U9533 ( .A(n8802), .ZN(n7072) );
  AOI21_X1 U9534 ( .B1(n7072), .B2(n6794), .A(n6699), .ZN(n8825) );
  OAI21_X1 U9535 ( .B1(n8802), .B2(n7077), .A(n6719), .ZN(n8827) );
  NAND2_X1 U9536 ( .A1(n8974), .A2(n6689), .ZN(n7079) );
  OAI21_X1 U9537 ( .B1(n8877), .B2(n6750), .A(n7086), .ZN(n8922) );
  NAND3_X1 U9538 ( .A1(n7086), .A2(n6750), .A3(n7085), .ZN(n7083) );
  INV_X1 U9539 ( .A(n8876), .ZN(n7091) );
  NAND2_X1 U9540 ( .A1(n8709), .A2(n7095), .ZN(n7092) );
  NAND2_X1 U9541 ( .A1(n7092), .A2(n6807), .ZN(n8755) );
  NAND2_X1 U9542 ( .A1(n11094), .A2(n11093), .ZN(n9693) );
  NAND2_X1 U9543 ( .A1(n7104), .A2(n9690), .ZN(n11094) );
  NAND2_X1 U9544 ( .A1(n11567), .A2(n11568), .ZN(n7104) );
  NAND2_X1 U9545 ( .A1(n9689), .A2(n9688), .ZN(n11567) );
  INV_X1 U9546 ( .A(n14150), .ZN(n7108) );
  OAI21_X1 U9547 ( .B1(n7108), .B2(n7111), .A(n7109), .ZN(n9732) );
  NAND2_X1 U9548 ( .A1(n9735), .A2(n7116), .ZN(n7119) );
  NAND2_X1 U9549 ( .A1(n14099), .A2(n9733), .ZN(n7127) );
  NAND4_X1 U9550 ( .A1(n7121), .A2(n7120), .A3(n7118), .A4(n7117), .ZN(n9741)
         );
  NAND3_X1 U9551 ( .A1(n6691), .A2(n14099), .A3(n9733), .ZN(n7117) );
  NAND2_X1 U9552 ( .A1(n7127), .A2(n9734), .ZN(n14085) );
  NAND2_X1 U9553 ( .A1(n7131), .A2(n15254), .ZN(n7130) );
  NAND4_X1 U9554 ( .A1(n7130), .A2(n7313), .A3(n7129), .A4(n7128), .ZN(n14215)
         );
  NAND3_X1 U9555 ( .A1(n7135), .A2(n7133), .A3(n7139), .ZN(n7128) );
  NAND3_X1 U9556 ( .A1(n7135), .A2(n7133), .A3(n6684), .ZN(n7129) );
  OR2_X1 U9557 ( .A1(n7600), .A2(n9715), .ZN(n7142) );
  NAND2_X1 U9558 ( .A1(n13302), .A2(n7155), .ZN(n7150) );
  NAND3_X1 U9559 ( .A1(n7151), .A2(n7152), .A3(n7150), .ZN(n13337) );
  OR2_X1 U9560 ( .A1(n13302), .A2(n13303), .ZN(n13335) );
  INV_X1 U9561 ( .A(n13303), .ZN(n7154) );
  NAND2_X1 U9562 ( .A1(n7181), .A2(n7177), .ZN(n7176) );
  NAND2_X1 U9563 ( .A1(n8907), .A2(n7182), .ZN(n7181) );
  INV_X1 U9564 ( .A(n7168), .ZN(n7167) );
  OAI21_X1 U9565 ( .B1(n8907), .B2(n7178), .A(n7169), .ZN(n7168) );
  NAND3_X1 U9566 ( .A1(n7176), .A2(n7175), .A3(n7179), .ZN(n8976) );
  OAI21_X1 U9567 ( .B1(n8503), .B2(n8506), .A(n7183), .ZN(n8533) );
  AOI21_X1 U9568 ( .B1(n8507), .B2(n7185), .A(n7184), .ZN(n7183) );
  INV_X1 U9569 ( .A(n8502), .ZN(n7185) );
  NAND2_X1 U9570 ( .A1(n8508), .A2(n8507), .ZN(n8528) );
  NAND2_X1 U9571 ( .A1(n8503), .A2(n8502), .ZN(n8508) );
  NAND2_X1 U9572 ( .A1(n8438), .A2(n8437), .ZN(n8439) );
  NAND2_X1 U9573 ( .A1(n8405), .A2(n7188), .ZN(n7187) );
  INV_X1 U9574 ( .A(n8404), .ZN(n7189) );
  NAND2_X1 U9575 ( .A1(n8665), .A2(n7194), .ZN(n7193) );
  NAND2_X1 U9576 ( .A1(n7801), .A2(n7202), .ZN(n7201) );
  OAI21_X1 U9577 ( .B1(n7801), .B2(n7552), .A(n7202), .ZN(n8008) );
  NAND3_X1 U9578 ( .A1(n7206), .A2(n7820), .A3(n7205), .ZN(n8151) );
  NAND2_X1 U9579 ( .A1(n7538), .A2(n7207), .ZN(n8142) );
  NAND2_X1 U9580 ( .A1(n7540), .A2(n6827), .ZN(n7207) );
  NAND2_X1 U9581 ( .A1(n8055), .A2(n7212), .ZN(n7210) );
  NAND3_X1 U9582 ( .A1(n7214), .A2(n7216), .A3(n7930), .ZN(n7797) );
  OAI21_X1 U9583 ( .B1(n8336), .B2(n6833), .A(n7223), .ZN(n7227) );
  NAND2_X2 U9584 ( .A1(n9931), .A2(n12393), .ZN(n10509) );
  XNOR2_X2 U9585 ( .A(n7233), .B(n9927), .ZN(n12393) );
  NAND2_X1 U9586 ( .A1(n9926), .A2(n9927), .ZN(n7235) );
  OR2_X1 U9587 ( .A1(n12672), .A2(n14561), .ZN(n7242) );
  NAND2_X1 U9588 ( .A1(n11667), .A2(n11668), .ZN(n11685) );
  NAND2_X1 U9589 ( .A1(n7240), .A2(n7239), .ZN(n7238) );
  NAND2_X1 U9590 ( .A1(n10510), .A2(n7242), .ZN(n7244) );
  NAND2_X1 U9591 ( .A1(n14457), .A2(n6704), .ZN(n7248) );
  OAI22_X2 U9592 ( .A1(n15315), .A2(n15314), .B1(n12669), .B2(n12668), .ZN(
        n15346) );
  OAI21_X1 U9593 ( .B1(n15346), .B2(n7256), .A(n7253), .ZN(n7478) );
  INV_X1 U9594 ( .A(n7750), .ZN(n7259) );
  NAND4_X1 U9595 ( .A1(n7584), .A2(n10012), .A3(n7260), .A4(n9922), .ZN(n9923)
         );
  NAND3_X1 U9596 ( .A1(n7584), .A2(n10012), .A3(n9921), .ZN(n10206) );
  NAND3_X1 U9597 ( .A1(n14505), .A2(n7483), .A3(n11689), .ZN(n7484) );
  AND3_X2 U9598 ( .A1(n7895), .A2(n7266), .A3(n7265), .ZN(n11069) );
  NAND3_X1 U9599 ( .A1(n7271), .A2(n7269), .A3(n7267), .ZN(n15148) );
  NAND3_X1 U9600 ( .A1(n7271), .A2(n7268), .A3(n7267), .ZN(n7272) );
  INV_X1 U9601 ( .A(n7272), .ZN(n15147) );
  OR2_X1 U9602 ( .A1(n13331), .A2(n13332), .ZN(n7275) );
  INV_X1 U9603 ( .A(n7275), .ZN(n13352) );
  NAND2_X1 U9604 ( .A1(n13353), .A2(n13361), .ZN(n7274) );
  NAND2_X1 U9605 ( .A1(n11148), .A2(n11146), .ZN(n7285) );
  INV_X1 U9606 ( .A(n11147), .ZN(n7284) );
  NAND3_X1 U9607 ( .A1(n12653), .A2(n6697), .A3(n12310), .ZN(n12644) );
  NAND2_X1 U9608 ( .A1(n13523), .A2(n13197), .ZN(n13509) );
  INV_X1 U9609 ( .A(n13522), .ZN(n7326) );
  NAND2_X1 U9610 ( .A1(n8438), .A2(n6793), .ZN(n7662) );
  NAND2_X1 U9611 ( .A1(n14196), .A2(n7330), .ZN(n7329) );
  NAND2_X1 U9612 ( .A1(n7640), .A2(n7641), .ZN(n7845) );
  OAI21_X2 U9613 ( .B1(n10793), .B2(n8510), .A(n8619), .ZN(n11754) );
  OR2_X2 U9614 ( .A1(n14379), .A2(n9771), .ZN(n7341) );
  NOR2_X2 U9615 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n10126) );
  NAND2_X2 U9616 ( .A1(n12706), .A2(n7345), .ZN(n9956) );
  NAND2_X1 U9617 ( .A1(n12242), .A2(n7348), .ZN(n7347) );
  NAND2_X1 U9618 ( .A1(n12298), .A2(n12297), .ZN(n12300) );
  NAND2_X1 U9619 ( .A1(n12467), .A2(n6737), .ZN(n7350) );
  NOR2_X1 U9620 ( .A1(n14796), .A2(n7752), .ZN(n14782) );
  OAI21_X2 U9621 ( .B1(n12691), .B2(n7363), .A(n7359), .ZN(n14949) );
  INV_X1 U9622 ( .A(n7368), .ZN(n10492) );
  INV_X1 U9623 ( .A(n7375), .ZN(n11261) );
  INV_X1 U9624 ( .A(n7380), .ZN(n11497) );
  NAND2_X1 U9625 ( .A1(n7378), .A2(n7377), .ZN(n7376) );
  NAND2_X1 U9626 ( .A1(n12926), .A2(n7382), .ZN(n7381) );
  OAI211_X1 U9627 ( .C1(n12926), .C2(n7386), .A(n7383), .B(n7381), .ZN(n9862)
         );
  OAI21_X2 U9628 ( .B1(n13011), .B2(n9857), .A(n7390), .ZN(n12874) );
  NAND2_X1 U9629 ( .A1(n11931), .A2(n11930), .ZN(n12005) );
  NAND2_X1 U9630 ( .A1(n10126), .A2(n9888), .ZN(n10185) );
  INV_X1 U9631 ( .A(n7410), .ZN(n11140) );
  NAND2_X1 U9632 ( .A1(n12424), .A2(n7415), .ZN(n7414) );
  OAI211_X1 U9633 ( .C1(n12424), .C2(n12425), .A(n7416), .B(n7414), .ZN(n15734) );
  INV_X1 U9634 ( .A(n13259), .ZN(n13275) );
  INV_X1 U9635 ( .A(n10619), .ZN(n7424) );
  INV_X1 U9636 ( .A(n10618), .ZN(n7426) );
  OAI21_X1 U9637 ( .B1(n10959), .B2(n7436), .A(n11172), .ZN(n10962) );
  NAND2_X1 U9638 ( .A1(n10959), .A2(n7436), .ZN(n11172) );
  XNOR2_X1 U9639 ( .A(n11107), .B(n11106), .ZN(n7436) );
  NOR2_X1 U9640 ( .A1(n8379), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n7440) );
  INV_X1 U9641 ( .A(n13853), .ZN(n7443) );
  INV_X1 U9642 ( .A(n7446), .ZN(n13852) );
  NOR2_X1 U9643 ( .A1(n13852), .A2(n13756), .ZN(n13823) );
  NAND2_X1 U9644 ( .A1(n11340), .A2(n7462), .ZN(n11483) );
  NAND2_X1 U9645 ( .A1(n11221), .A2(n11228), .ZN(n11340) );
  NAND2_X1 U9646 ( .A1(n13723), .A2(n7463), .ZN(n13830) );
  NAND2_X1 U9647 ( .A1(n13830), .A2(n13726), .ZN(n13727) );
  OR2_X2 U9648 ( .A1(n15263), .A2(n14272), .ZN(n13804) );
  INV_X1 U9649 ( .A(n11524), .ZN(n7468) );
  NAND2_X1 U9650 ( .A1(n7468), .A2(n7469), .ZN(n11654) );
  NOR2_X2 U9651 ( .A1(n14090), .A2(n7471), .ZN(n14057) );
  INV_X1 U9652 ( .A(n14057), .ZN(n14049) );
  NAND3_X1 U9653 ( .A1(n11807), .A2(n7474), .A3(n7473), .ZN(n15264) );
  INV_X1 U9654 ( .A(n7484), .ZN(n11942) );
  OAI211_X1 U9655 ( .C1(n14539), .C2(n6810), .A(n7487), .B(n7485), .ZN(n12859)
         );
  NAND2_X1 U9656 ( .A1(n14539), .A2(n7486), .ZN(n7485) );
  NAND2_X1 U9657 ( .A1(n12234), .A2(n7493), .ZN(n7495) );
  INV_X1 U9658 ( .A(n12658), .ZN(n12660) );
  NAND2_X2 U9659 ( .A1(n7495), .A2(n6752), .ZN(n12658) );
  NAND2_X1 U9660 ( .A1(n14485), .A2(n6705), .ZN(n7499) );
  NAND2_X2 U9661 ( .A1(n7499), .A2(n6747), .ZN(n14457) );
  NAND2_X2 U9662 ( .A1(n6713), .A2(n7502), .ZN(n11920) );
  NAND2_X2 U9663 ( .A1(n9963), .A2(n9919), .ZN(n10110) );
  OAI21_X1 U9664 ( .B1(n14103), .B2(n7511), .A(n7510), .ZN(n14071) );
  NAND2_X1 U9665 ( .A1(n7509), .A2(n7508), .ZN(n9682) );
  NAND2_X1 U9666 ( .A1(n14103), .A2(n7510), .ZN(n7509) );
  INV_X1 U9667 ( .A(n7518), .ZN(n7519) );
  OAI21_X1 U9668 ( .B1(n7522), .B2(n6687), .A(n15267), .ZN(n7518) );
  NAND2_X1 U9669 ( .A1(n12043), .A2(n7523), .ZN(n7520) );
  NAND2_X1 U9670 ( .A1(n7520), .A2(n7519), .ZN(n15265) );
  NAND2_X2 U9671 ( .A1(n12484), .A2(n9666), .ZN(n12483) );
  NAND2_X1 U9672 ( .A1(n14147), .A2(n7534), .ZN(n14315) );
  NAND3_X1 U9673 ( .A1(n7537), .A2(n7536), .A3(n13223), .ZN(n13230) );
  OR2_X1 U9674 ( .A1(n13222), .A2(n13228), .ZN(n7537) );
  AOI21_X1 U9675 ( .B1(n8131), .B2(n6702), .A(n6832), .ZN(n7538) );
  INV_X1 U9676 ( .A(n7792), .ZN(n7543) );
  NAND2_X1 U9677 ( .A1(n10241), .A2(n7556), .ZN(n7555) );
  INV_X1 U9678 ( .A(n10240), .ZN(n7562) );
  NAND3_X1 U9679 ( .A1(n10138), .A2(n10137), .A3(n6799), .ZN(n7563) );
  NAND2_X1 U9680 ( .A1(n7563), .A2(n7564), .ZN(n10166) );
  NAND3_X1 U9681 ( .A1(n10033), .A2(n10032), .A3(n6802), .ZN(n7565) );
  NAND2_X1 U9682 ( .A1(n7565), .A2(n7566), .ZN(n10063) );
  NAND2_X1 U9683 ( .A1(n9926), .A2(n6797), .ZN(n10487) );
  NAND2_X1 U9684 ( .A1(n7569), .A2(n7570), .ZN(n10133) );
  NAND3_X1 U9685 ( .A1(n10101), .A2(n10100), .A3(n6809), .ZN(n7569) );
  OAI21_X1 U9686 ( .B1(n7572), .B2(n10307), .A(n7573), .ZN(n10331) );
  NAND3_X1 U9687 ( .A1(n10336), .A2(n10335), .A3(n6798), .ZN(n7575) );
  NAND2_X1 U9688 ( .A1(n7575), .A2(n7576), .ZN(n10358) );
  NAND3_X1 U9689 ( .A1(n10068), .A2(n10067), .A3(n6800), .ZN(n7578) );
  NAND2_X1 U9690 ( .A1(n7578), .A2(n7579), .ZN(n10096) );
  NAND3_X1 U9691 ( .A1(n10363), .A2(n10362), .A3(n6801), .ZN(n7581) );
  NAND2_X1 U9692 ( .A1(n7581), .A2(n7582), .ZN(n10390) );
  NAND4_X1 U9693 ( .A1(n9890), .A2(n9891), .A3(n9892), .A4(n9889), .ZN(n7585)
         );
  XNOR2_X2 U9694 ( .A(n15698), .B(n9686), .ZN(n11842) );
  OAI21_X1 U9695 ( .B1(n10760), .B2(n7592), .A(n7590), .ZN(n7589) );
  NAND2_X1 U9696 ( .A1(n10760), .A2(n7591), .ZN(n7590) );
  INV_X1 U9697 ( .A(n9715), .ZN(n7603) );
  OAI21_X1 U9698 ( .B1(n14287), .B2(n15729), .A(n14289), .ZN(n14290) );
  OR2_X1 U9699 ( .A1(n12038), .A2(n7605), .ZN(n7604) );
  OR2_X1 U9700 ( .A1(n12038), .A2(n9706), .ZN(n7613) );
  NAND2_X1 U9701 ( .A1(n7604), .A2(n7608), .ZN(n9711) );
  INV_X1 U9702 ( .A(n13544), .ZN(n7620) );
  NAND2_X1 U9703 ( .A1(n7621), .A2(n7625), .ZN(n13408) );
  NAND2_X1 U9704 ( .A1(n13430), .A2(n7622), .ZN(n7621) );
  NAND2_X1 U9705 ( .A1(n8237), .A2(n8236), .ZN(n12633) );
  INV_X1 U9706 ( .A(n8236), .ZN(n7637) );
  NAND3_X1 U9707 ( .A1(n7165), .A2(n10614), .A3(n7770), .ZN(n7906) );
  NAND2_X1 U9708 ( .A1(n8613), .A2(n8612), .ZN(n8633) );
  OAI21_X1 U9709 ( .B1(n8613), .B2(n7649), .A(n7647), .ZN(n8660) );
  OAI21_X1 U9710 ( .B1(n9020), .B2(n9019), .A(n9018), .ZN(n7656) );
  AOI21_X1 U9711 ( .B1(n9018), .B2(n7652), .A(n7651), .ZN(n7650) );
  NAND2_X1 U9712 ( .A1(n9020), .A2(n7654), .ZN(n7653) );
  XNOR2_X1 U9713 ( .A(n7656), .B(n9037), .ZN(n14426) );
  NAND2_X1 U9714 ( .A1(n7658), .A2(n10491), .ZN(n10506) );
  NAND4_X1 U9715 ( .A1(n7659), .A2(n10486), .A3(n10485), .A4(n10484), .ZN(
        n7658) );
  NAND2_X1 U9716 ( .A1(n7660), .A2(n10434), .ZN(n7659) );
  INV_X1 U9717 ( .A(n10441), .ZN(n7660) );
  NAND2_X1 U9718 ( .A1(n7661), .A2(n8444), .ZN(n8447) );
  AND2_X1 U9719 ( .A1(n7672), .A2(n6724), .ZN(n8806) );
  NAND2_X1 U9720 ( .A1(n7672), .A2(n6804), .ZN(n8808) );
  XNOR2_X1 U9721 ( .A(n8765), .B(SI_14_), .ZN(n8782) );
  AND2_X1 U9722 ( .A1(n9957), .A2(n9958), .ZN(n7673) );
  INV_X1 U9723 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7674) );
  NAND2_X1 U9724 ( .A1(n12598), .A2(n7677), .ZN(n7676) );
  INV_X1 U9725 ( .A(n12696), .ZN(n7684) );
  NAND2_X1 U9726 ( .A1(n6682), .A2(n12696), .ZN(n7680) );
  OAI21_X1 U9727 ( .B1(n12002), .B2(n7692), .A(n7690), .ZN(n7691) );
  AOI21_X1 U9728 ( .B1(n12050), .B2(n12056), .A(n6788), .ZN(n7690) );
  NAND2_X1 U9729 ( .A1(n7691), .A2(n12249), .ZN(n12253) );
  INV_X1 U9730 ( .A(n12056), .ZN(n7692) );
  INV_X2 U9731 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7693) );
  NAND2_X1 U9732 ( .A1(n14748), .A2(n7697), .ZN(n7695) );
  NAND2_X1 U9733 ( .A1(n7695), .A2(n7694), .ZN(n14903) );
  NAND2_X1 U9734 ( .A1(n7699), .A2(n7702), .ZN(n14758) );
  NAND2_X1 U9735 ( .A1(n14754), .A2(n7700), .ZN(n7699) );
  NAND2_X1 U9736 ( .A1(n14786), .A2(n14794), .ZN(n14788) );
  NAND2_X1 U9737 ( .A1(n7709), .A2(n7712), .ZN(n14766) );
  NAND2_X1 U9738 ( .A1(n14786), .A2(n7710), .ZN(n7709) );
  NAND2_X1 U9739 ( .A1(n10492), .A2(n7716), .ZN(n9914) );
  NAND2_X1 U9740 ( .A1(n12304), .A2(n7719), .ZN(n12470) );
  NAND2_X1 U9741 ( .A1(n8585), .A2(n6744), .ZN(n7721) );
  NAND2_X1 U9742 ( .A1(n9056), .A2(n9095), .ZN(n7723) );
  NAND2_X1 U9743 ( .A1(n9052), .A2(n9095), .ZN(n7724) );
  NAND3_X1 U9744 ( .A1(n7724), .A2(n7723), .A3(n6751), .ZN(n9161) );
  NAND3_X1 U9745 ( .A1(n8760), .A2(n8759), .A3(n6805), .ZN(n7728) );
  NAND2_X1 U9746 ( .A1(n7729), .A2(n6822), .ZN(n8877) );
  NAND3_X1 U9747 ( .A1(n8828), .A2(n6803), .A3(n6694), .ZN(n7729) );
  NOR2_X1 U9748 ( .A1(n8395), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n8411) );
  NAND3_X1 U9749 ( .A1(n8410), .A2(n7738), .A3(n7113), .ZN(n7737) );
  INV_X1 U9750 ( .A(n8896), .ZN(n7742) );
  INV_X1 U9751 ( .A(n8384), .ZN(n8386) );
  NAND2_X1 U9752 ( .A1(n8209), .A2(n8208), .ZN(n13427) );
  NOR2_X2 U9753 ( .A1(n13783), .A2(n11562), .ZN(n11563) );
  AOI21_X1 U9754 ( .B1(n9950), .B2(n9949), .A(n11919), .ZN(n9968) );
  OR2_X1 U9755 ( .A1(n8183), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7825) );
  NAND2_X1 U9756 ( .A1(n9741), .A2(n15256), .ZN(n9744) );
  BUF_X8 U9757 ( .A(n10525), .Z(n12849) );
  NAND2_X1 U9758 ( .A1(n11443), .A2(n11920), .ZN(n11910) );
  NAND2_X1 U9759 ( .A1(n14563), .A2(n10525), .ZN(n10526) );
  OR2_X1 U9760 ( .A1(n9785), .A2(n9850), .ZN(n9786) );
  XNOR2_X1 U9761 ( .A(n9061), .B(n9038), .ZN(n14423) );
  INV_X1 U9762 ( .A(n7850), .ZN(n13695) );
  INV_X1 U9763 ( .A(n15500), .ZN(n9966) );
  NAND2_X1 U9764 ( .A1(n13751), .A2(n7744), .ZN(n13752) );
  INV_X1 U9765 ( .A(n12788), .ZN(n10519) );
  NOR2_X1 U9766 ( .A1(n9153), .A2(n9147), .ZN(n9160) );
  NAND2_X1 U9767 ( .A1(n9952), .A2(n9951), .ZN(n9955) );
  OR2_X1 U9768 ( .A1(n9901), .A2(n10013), .ZN(n9903) );
  INV_X1 U9769 ( .A(n10412), .ZN(n10563) );
  OR2_X1 U9770 ( .A1(n10412), .A2(n14973), .ZN(n9925) );
  INV_X1 U9771 ( .A(n10445), .ZN(n14982) );
  OR2_X1 U9772 ( .A1(n15263), .A2(n9162), .ZN(n10964) );
  OR2_X1 U9773 ( .A1(n9163), .A2(n9162), .ZN(n7745) );
  AND2_X1 U9774 ( .A1(n6673), .A2(n8434), .ZN(n7746) );
  AND2_X2 U9775 ( .A1(n11464), .A2(n8308), .ZN(n15854) );
  NAND2_X1 U9776 ( .A1(n8386), .A2(n8385), .ZN(n7747) );
  OR2_X1 U9777 ( .A1(n13425), .A2(n13676), .ZN(n7748) );
  OR2_X1 U9778 ( .A1(n13425), .A2(n13626), .ZN(n7749) );
  AND2_X1 U9779 ( .A1(n12676), .A2(n12675), .ZN(n7750) );
  AND2_X1 U9780 ( .A1(n9795), .A2(n12027), .ZN(n7751) );
  AND2_X1 U9781 ( .A1(n15001), .A2(n14723), .ZN(n7752) );
  OR2_X1 U9782 ( .A1(n15001), .A2(n14764), .ZN(n7753) );
  OR2_X1 U9783 ( .A1(n9166), .A2(n9748), .ZN(n7754) );
  OR2_X1 U9784 ( .A1(n10760), .A2(n8477), .ZN(n7755) );
  INV_X1 U9785 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10013) );
  AND2_X2 U9786 ( .A1(n8319), .A2(n9860), .ZN(n15846) );
  OR2_X1 U9787 ( .A1(n8954), .A2(SI_20_), .ZN(n7759) );
  AND2_X1 U9788 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7760) );
  INV_X1 U9789 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12390) );
  INV_X1 U9790 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n7924) );
  INV_X1 U9791 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9899) );
  INV_X1 U9792 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n7986) );
  NAND2_X1 U9793 ( .A1(n8367), .A2(n8391), .ZN(n8379) );
  INV_X1 U9794 ( .A(n12630), .ZN(n10491) );
  XOR2_X1 U9795 ( .A(n7882), .B(n7881), .Z(n7761) );
  INV_X1 U9796 ( .A(n15652), .ZN(n15659) );
  INV_X1 U9797 ( .A(n10677), .ZN(n10623) );
  INV_X1 U9798 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7818) );
  AND2_X1 U9799 ( .A1(n12191), .A2(n13936), .ZN(n7762) );
  OR2_X1 U9800 ( .A1(n12191), .A2(n13936), .ZN(n7763) );
  AND2_X1 U9801 ( .A1(n9791), .A2(n11796), .ZN(n7764) );
  INV_X1 U9802 ( .A(n12659), .ZN(n12547) );
  OR2_X1 U9803 ( .A1(n8956), .A2(SI_21_), .ZN(n7765) );
  INV_X1 U9804 ( .A(n9193), .ZN(n9166) );
  AND2_X2 U9805 ( .A1(n10896), .A2(n11556), .ZN(n15724) );
  AND2_X1 U9806 ( .A1(n9740), .A2(n9739), .ZN(n15668) );
  XOR2_X1 U9807 ( .A(n9191), .B(n14272), .Z(n7766) );
  AND2_X1 U9808 ( .A1(n10522), .A2(n10521), .ZN(n7767) );
  AND2_X1 U9809 ( .A1(n8047), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n7768) );
  INV_X1 U9810 ( .A(n13507), .ZN(n13482) );
  AND2_X1 U9811 ( .A1(n8171), .A2(n8170), .ZN(n13507) );
  NOR2_X1 U9812 ( .A1(n12709), .A2(n13466), .ZN(n7769) );
  INV_X1 U9813 ( .A(n12953), .ZN(n9848) );
  INV_X1 U9814 ( .A(n15691), .ZN(n8434) );
  NAND2_X1 U9815 ( .A1(n8482), .A2(n8481), .ZN(n8492) );
  AOI21_X1 U9816 ( .B1(n11125), .B2(n6673), .A(n8519), .ZN(n8523) );
  NAND2_X1 U9817 ( .A1(n9987), .A2(n9951), .ZN(n9988) );
  INV_X1 U9818 ( .A(n8554), .ZN(n8555) );
  NAND2_X1 U9819 ( .A1(n8556), .A2(n8555), .ZN(n8557) );
  INV_X1 U9820 ( .A(n8653), .ZN(n8654) );
  INV_X1 U9821 ( .A(n8752), .ZN(n8753) );
  INV_X1 U9822 ( .A(n10167), .ZN(n10168) );
  OAI21_X1 U9823 ( .B1(n6673), .B2(n9713), .A(n8800), .ZN(n8801) );
  OAI21_X1 U9824 ( .B1(n10232), .B2(n10231), .A(n10230), .ZN(n10241) );
  INV_X1 U9825 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7777) );
  CLKBUF_X3 U9826 ( .A(n10025), .Z(n10428) );
  INV_X1 U9827 ( .A(n12297), .ZN(n12250) );
  AND2_X1 U9828 ( .A1(n10617), .A2(n11209), .ZN(n10618) );
  NOR2_X1 U9829 ( .A1(n8093), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8109) );
  AOI22_X1 U9830 ( .A1(n9173), .A2(n9114), .B1(n6673), .B2(n13918), .ZN(n9150)
         );
  OR2_X1 U9831 ( .A1(n12730), .A2(n12729), .ZN(n12731) );
  OAI22_X1 U9832 ( .A1(n11506), .A2(n12787), .B1(n10543), .B2(n7693), .ZN(
        n10520) );
  MUX2_X1 U9833 ( .A(n12853), .B(n14989), .S(n10428), .Z(n10397) );
  INV_X1 U9834 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n8403) );
  INV_X1 U9835 ( .A(n13148), .ZN(n9803) );
  INV_X1 U9836 ( .A(n15816), .ZN(n9783) );
  INV_X1 U9837 ( .A(n10624), .ZN(n10625) );
  OR2_X1 U9838 ( .A1(n7862), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8261) );
  NAND2_X1 U9839 ( .A1(n8165), .A2(n9564), .ZN(n8176) );
  NAND2_X1 U9840 ( .A1(n8123), .A2(n13002), .ZN(n8135) );
  INV_X1 U9841 ( .A(n13062), .ZN(n8221) );
  AND2_X1 U9842 ( .A1(n13415), .A2(n11821), .ZN(n8341) );
  INV_X1 U9843 ( .A(n8272), .ZN(n8273) );
  INV_X1 U9844 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8022) );
  OR2_X1 U9845 ( .A1(n9190), .A2(n9146), .ZN(n9147) );
  AND2_X1 U9846 ( .A1(n9065), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n9066) );
  NOR2_X1 U9847 ( .A1(n8792), .A2(n12566), .ZN(n8816) );
  INV_X1 U9848 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8620) );
  INV_X1 U9849 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8366) );
  INV_X1 U9850 ( .A(n12819), .ZN(n10529) );
  NOR2_X1 U9851 ( .A1(n12660), .A2(n12547), .ZN(n12661) );
  NAND2_X1 U9852 ( .A1(n14563), .A2(n10519), .ZN(n10522) );
  INV_X1 U9853 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10070) );
  INV_X1 U9854 ( .A(n12526), .ZN(n12471) );
  INV_X1 U9855 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9887) );
  XNOR2_X1 U9856 ( .A(n9850), .B(n9783), .ZN(n9784) );
  AND2_X1 U9857 ( .A1(n12496), .A2(n8282), .ZN(n8296) );
  INV_X1 U9858 ( .A(n13365), .ZN(n13363) );
  INV_X1 U9859 ( .A(n13214), .ZN(n13445) );
  INV_X1 U9860 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n12883) );
  AND2_X1 U9861 ( .A1(n8283), .A2(n10985), .ZN(n11461) );
  INV_X1 U9862 ( .A(n13079), .ZN(n8342) );
  OR2_X1 U9863 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n11609), .ZN(n7812) );
  INV_X1 U9864 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7793) );
  INV_X1 U9865 ( .A(n13833), .ZN(n13724) );
  NOR2_X1 U9866 ( .A1(n8910), .A2(n13868), .ZN(n8933) );
  INV_X1 U9867 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8543) );
  OR2_X1 U9868 ( .A1(n8865), .A2(n12373), .ZN(n8888) );
  AND2_X1 U9869 ( .A1(n14045), .A2(n12341), .ZN(n15578) );
  OR2_X1 U9870 ( .A1(n8621), .A2(n8620), .ZN(n8645) );
  NAND2_X1 U9871 ( .A1(n14212), .A2(n14213), .ZN(n14198) );
  NAND2_X1 U9872 ( .A1(n9696), .A2(n9695), .ZN(n11389) );
  OR2_X1 U9873 ( .A1(n8766), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n8786) );
  INV_X1 U9874 ( .A(n12068), .ZN(n12069) );
  NAND2_X1 U9875 ( .A1(n10530), .A2(n10529), .ZN(n10531) );
  INV_X1 U9876 ( .A(n11685), .ZN(n11687) );
  INV_X1 U9877 ( .A(n12769), .ZN(n12772) );
  INV_X1 U9878 ( .A(n14531), .ZN(n12763) );
  INV_X1 U9879 ( .A(n10295), .ZN(n10310) );
  OR2_X1 U9880 ( .A1(n10246), .A2(n10245), .ZN(n10259) );
  INV_X1 U9881 ( .A(n10309), .ZN(n10322) );
  AND2_X1 U9882 ( .A1(n10038), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10055) );
  INV_X1 U9883 ( .A(n14687), .ZN(n14972) );
  NAND2_X1 U9884 ( .A1(n8809), .A2(n10975), .ZN(n8831) );
  NAND2_X1 U9885 ( .A1(n8661), .A2(SI_10_), .ZN(n8689) );
  INV_X1 U9886 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n9582) );
  OR2_X1 U9887 ( .A1(n9251), .A2(n9250), .ZN(n9239) );
  NAND2_X1 U9888 ( .A1(n9796), .A2(n11963), .ZN(n9797) );
  OR2_X1 U9889 ( .A1(n9792), .A2(n11427), .ZN(n9793) );
  NOR2_X1 U9890 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n7923) );
  NOR2_X1 U9891 ( .A1(n8144), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8155) );
  OR2_X1 U9892 ( .A1(n8077), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8093) );
  AOI21_X1 U9893 ( .B1(n13416), .B2(n8328), .A(n8265), .ZN(n9880) );
  INV_X1 U9894 ( .A(n10629), .ZN(n10631) );
  INV_X1 U9895 ( .A(n12425), .ZN(n12426) );
  INV_X1 U9896 ( .A(n13574), .ZN(n13546) );
  OR2_X1 U9897 ( .A1(n8036), .A2(n7843), .ZN(n8047) );
  OR2_X1 U9898 ( .A1(n8001), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8036) );
  AND2_X1 U9899 ( .A1(n7967), .A2(n11407), .ZN(n7987) );
  OR2_X1 U9900 ( .A1(n7939), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U9901 ( .A1(n15217), .A2(n15796), .ZN(n15760) );
  INV_X1 U9902 ( .A(n13224), .ZN(n13425) );
  AND2_X1 U9903 ( .A1(n13162), .A2(n13165), .ZN(n15214) );
  INV_X1 U9904 ( .A(n8215), .ZN(n13063) );
  NAND2_X1 U9905 ( .A1(n10588), .A2(n13685), .ZN(n10608) );
  INV_X1 U9906 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8297) );
  NOR2_X1 U9907 ( .A1(n8983), .A2(n13774), .ZN(n9004) );
  OR2_X1 U9908 ( .A1(n8962), .A2(n13883), .ZN(n8983) );
  INV_X1 U9909 ( .A(n13891), .ZN(n13736) );
  INV_X1 U9910 ( .A(n13910), .ZN(n13884) );
  OR2_X1 U9911 ( .A1(n8888), .A2(n8887), .ZN(n8910) );
  INV_X1 U9912 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n11489) );
  OR2_X1 U9913 ( .A1(n10836), .A2(n10835), .ZN(n10873) );
  OR2_X1 U9914 ( .A1(n10841), .A2(n10840), .ZN(n10866) );
  AND2_X1 U9915 ( .A1(n15578), .A2(n15577), .ZN(n15580) );
  NOR2_X1 U9916 ( .A1(n8411), .A2(n8398), .ZN(n8399) );
  XNOR2_X1 U9917 ( .A(n14056), .B(n14050), .ZN(n14051) );
  NAND2_X1 U9918 ( .A1(n9705), .A2(n9704), .ZN(n12038) );
  INV_X1 U9919 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n14288) );
  INV_X1 U9920 ( .A(n15724), .ZN(n9771) );
  NAND2_X1 U9921 ( .A1(n12707), .A2(n9162), .ZN(n9773) );
  AND2_X1 U9922 ( .A1(n14427), .A2(n9758), .ZN(n9759) );
  INV_X1 U9923 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8377) );
  INV_X1 U9924 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10102) );
  OR2_X1 U9925 ( .A1(n12232), .A2(n12231), .ZN(n12233) );
  NAND2_X1 U9926 ( .A1(n7767), .A2(n11373), .ZN(n11372) );
  INV_X1 U9927 ( .A(n14557), .ZN(n12247) );
  NAND2_X1 U9928 ( .A1(n10441), .A2(n10440), .ZN(n10486) );
  AND2_X1 U9929 ( .A1(n10266), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n10277) );
  INV_X1 U9930 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n12683) );
  INV_X1 U9931 ( .A(n10501), .ZN(n10931) );
  INV_X1 U9932 ( .A(n14720), .ZN(n14846) );
  INV_X1 U9933 ( .A(n14765), .ZN(n14725) );
  INV_X1 U9934 ( .A(n15545), .ZN(n15387) );
  AND3_X1 U9935 ( .A1(n11436), .A2(n11435), .A3(n11434), .ZN(n11437) );
  AND2_X1 U9936 ( .A1(n8859), .A2(n8835), .ZN(n8857) );
  AND2_X1 U9937 ( .A1(n8586), .A2(n8562), .ZN(n8563) );
  NAND2_X1 U9938 ( .A1(n8473), .A2(n8443), .ZN(n8448) );
  OAI21_X1 U9939 ( .B1(n9232), .B2(n9231), .A(n9230), .ZN(n9255) );
  OAI21_X1 U9940 ( .B1(n13425), .B2(n13035), .A(n9883), .ZN(n9884) );
  INV_X1 U9941 ( .A(n13016), .ZN(n13026) );
  INV_X1 U9942 ( .A(n13035), .ZN(n13006) );
  OR2_X1 U9943 ( .A1(n11267), .A2(n9875), .ZN(n13031) );
  OR2_X1 U9944 ( .A1(n10588), .A2(n11266), .ZN(n10689) );
  INV_X1 U9945 ( .A(n15738), .ZN(n13349) );
  INV_X1 U9946 ( .A(n15789), .ZN(n15806) );
  NOR2_X1 U9947 ( .A1(n7952), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7967) );
  INV_X1 U9948 ( .A(n13124), .ZN(n11779) );
  AND2_X1 U9949 ( .A1(n8301), .A2(n8316), .ZN(n11464) );
  OR2_X1 U9950 ( .A1(n15814), .A2(n15842), .ZN(n15241) );
  AND2_X1 U9951 ( .A1(n10764), .A2(n10763), .ZN(n10769) );
  AND2_X1 U9952 ( .A1(n10968), .A2(n10967), .ZN(n13910) );
  NOR2_X1 U9953 ( .A1(n11554), .A2(n10954), .ZN(n10968) );
  OR2_X1 U9954 ( .A1(n12367), .A2(n15642), .ZN(n15643) );
  INV_X1 U9955 ( .A(n15654), .ZN(n15270) );
  INV_X1 U9956 ( .A(n15663), .ZN(n15261) );
  INV_X1 U9957 ( .A(n15668), .ZN(n15256) );
  INV_X1 U9958 ( .A(n14351), .ZN(n14333) );
  INV_X1 U9959 ( .A(n14401), .ZN(n9774) );
  AND2_X1 U9960 ( .A1(n15690), .A2(n9773), .ZN(n15281) );
  NAND2_X1 U9961 ( .A1(n15711), .A2(n15710), .ZN(n15722) );
  INV_X1 U9962 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9195) );
  AND2_X1 U9963 ( .A1(n8695), .A2(n8714), .ZN(n14040) );
  OR2_X1 U9964 ( .A1(n10103), .A2(n10102), .ZN(n10120) );
  AND2_X1 U9965 ( .A1(n10220), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10222) );
  NAND2_X1 U9966 ( .A1(n10583), .A2(n14975), .ZN(n15351) );
  NOR2_X1 U9967 ( .A1(n10193), .A2(n10192), .ZN(n10220) );
  AND4_X1 U9968 ( .A1(n10302), .A2(n10301), .A3(n10300), .A4(n10299), .ZN(
        n14714) );
  INV_X1 U9969 ( .A(n15481), .ZN(n15462) );
  XNOR2_X1 U9970 ( .A(n15041), .B(n14712), .ZN(n14891) );
  INV_X1 U9971 ( .A(n14979), .ZN(n14958) );
  INV_X1 U9972 ( .A(n15497), .ZN(n14963) );
  AND2_X1 U9973 ( .A1(n10560), .A2(n10785), .ZN(n14732) );
  NAND2_X1 U9974 ( .A1(n11442), .A2(n11441), .ZN(n15534) );
  INV_X1 U9975 ( .A(n14732), .ZN(n11824) );
  NAND2_X1 U9976 ( .A1(n10546), .A2(n10558), .ZN(n10571) );
  AND2_X1 U9977 ( .A1(n8559), .A2(n8534), .ZN(n10743) );
  AND2_X1 U9978 ( .A1(n10692), .A2(n10691), .ZN(n15732) );
  INV_X1 U9979 ( .A(n9884), .ZN(n9885) );
  INV_X1 U9980 ( .A(n13031), .ZN(n12958) );
  INV_X1 U9981 ( .A(n13496), .ZN(n13519) );
  OR2_X1 U9982 ( .A1(n10688), .A2(n10632), .ZN(n15752) );
  AND2_X1 U9983 ( .A1(n13521), .A2(n13520), .ZN(n13616) );
  NAND2_X1 U9984 ( .A1(n11465), .A2(n15798), .ZN(n15782) );
  NAND2_X1 U9985 ( .A1(n11466), .A2(n15782), .ZN(n15801) );
  INV_X1 U9986 ( .A(n15854), .ZN(n15851) );
  INV_X1 U9987 ( .A(n8358), .ZN(n8359) );
  INV_X1 U9988 ( .A(n15846), .ZN(n15844) );
  NAND2_X1 U9989 ( .A1(n8284), .A2(n13685), .ZN(n10984) );
  INV_X1 U9990 ( .A(SI_20_), .ZN(n11661) );
  INV_X1 U9991 ( .A(SI_18_), .ZN(n11183) );
  INV_X1 U9992 ( .A(SI_12_), .ZN(n10742) );
  INV_X1 U9993 ( .A(SI_5_), .ZN(n10701) );
  INV_X1 U9994 ( .A(n10648), .ZN(n11030) );
  INV_X1 U9995 ( .A(n13914), .ZN(n13901) );
  INV_X1 U9996 ( .A(n13809), .ZN(n13919) );
  CLKBUF_X2 U9997 ( .A(P2_U3947), .Z(n15560) );
  INV_X1 U9998 ( .A(n15635), .ZN(n15592) );
  AND2_X1 U9999 ( .A1(n11561), .A2(n15676), .ZN(n15652) );
  INV_X1 U10000 ( .A(n15659), .ZN(n15678) );
  OR2_X1 U10001 ( .A1(n15652), .A2(n11558), .ZN(n14261) );
  INV_X1 U10002 ( .A(n14108), .ZN(n14385) );
  OR2_X1 U10003 ( .A1(n14369), .A2(n14368), .ZN(n14404) );
  OR2_X1 U10004 ( .A1(n15686), .A2(n15682), .ZN(n15683) );
  OR2_X1 U10005 ( .A1(n9765), .A2(P2_U3088), .ZN(n15686) );
  NAND2_X1 U10006 ( .A1(n9201), .A2(n8395), .ZN(n14424) );
  INV_X1 U10007 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12465) );
  INV_X1 U10008 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10981) );
  INV_X1 U10009 ( .A(n14802), .ZN(n15001) );
  INV_X1 U10010 ( .A(n11443), .ZN(n11508) );
  NAND2_X1 U10011 ( .A1(n11438), .A2(n10567), .ZN(n15337) );
  INV_X1 U10012 ( .A(n12853), .ZN(n14549) );
  INV_X1 U10013 ( .A(n15325), .ZN(n14705) );
  CLKBUF_X1 U10014 ( .A(n11443), .Z(n14562) );
  INV_X1 U10015 ( .A(n15460), .ZN(n15485) );
  AND2_X1 U10016 ( .A1(n14940), .A2(n14939), .ZN(n15059) );
  OR2_X1 U10017 ( .A1(n15509), .A2(n15393), .ZN(n14979) );
  OR2_X1 U10018 ( .A1(n15509), .A2(n15529), .ZN(n14960) );
  INV_X1 U10019 ( .A(n15559), .ZN(n15557) );
  NAND2_X1 U10020 ( .A1(n11503), .A2(n11824), .ZN(n15550) );
  AND2_X1 U10021 ( .A1(n10782), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10790) );
  XNOR2_X1 U10022 ( .A(n9924), .B(n9506), .ZN(n14973) );
  INV_X1 U10023 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n11258) );
  XNOR2_X1 U10024 ( .A(n9644), .B(n9643), .ZN(n9645) );
  INV_X1 U10025 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n8309) );
  NAND2_X1 U10026 ( .A1(n7780), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7782) );
  NAND2_X1 U10027 ( .A1(n11663), .A2(n13081), .ZN(n15817) );
  NAND2_X1 U10028 ( .A1(n6688), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7784) );
  MUX2_X1 U10029 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7784), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n7786) );
  OR2_X1 U10030 ( .A1(n15817), .A2(n13243), .ZN(n15831) );
  INV_X1 U10031 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n12628) );
  INV_X1 U10032 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n12388) );
  AOI22_X1 U10033 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n12390), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n12388), .ZN(n8129) );
  AOI22_X1 U10034 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n12317), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n12296), .ZN(n8115) );
  XNOR2_X1 U10035 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .ZN(n8100) );
  NAND2_X1 U10036 ( .A1(n7882), .A2(n7881), .ZN(n7788) );
  NAND2_X1 U10037 ( .A1(n10698), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7787) );
  NAND2_X1 U10038 ( .A1(n7788), .A2(n7787), .ZN(n7893) );
  XNOR2_X1 U10039 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n7891) );
  NAND2_X1 U10040 ( .A1(n7893), .A2(n7891), .ZN(n7790) );
  NAND2_X1 U10041 ( .A1(n8440), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7789) );
  NAND2_X1 U10042 ( .A1(n7791), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7792) );
  NAND2_X1 U10043 ( .A1(n7793), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7794) );
  NAND2_X1 U10044 ( .A1(n7795), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7796) );
  AND2_X1 U10045 ( .A1(n10750), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7798) );
  NAND2_X1 U10046 ( .A1(n10747), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7799) );
  NAND2_X1 U10047 ( .A1(n10751), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7800) );
  NAND2_X1 U10048 ( .A1(n7802), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7803) );
  XNOR2_X1 U10049 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n7994) );
  XNOR2_X1 U10050 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n8007) );
  NAND2_X1 U10051 ( .A1(n10883), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7805) );
  NOR2_X1 U10052 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n10981), .ZN(n7807) );
  NAND2_X1 U10053 ( .A1(n10981), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7808) );
  NAND2_X1 U10054 ( .A1(n8042), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7811) );
  NAND2_X1 U10055 ( .A1(n11609), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7813) );
  XNOR2_X1 U10056 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n8069) );
  NAND2_X1 U10057 ( .A1(n11804), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7814) );
  XNOR2_X1 U10058 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n8084) );
  NAND2_X1 U10059 ( .A1(n8100), .A2(n8101), .ZN(n7815) );
  NAND2_X1 U10060 ( .A1(n8115), .A2(n8117), .ZN(n7816) );
  NAND2_X1 U10061 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n7819), .ZN(n7820) );
  INV_X1 U10062 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n12392) );
  INV_X1 U10063 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12511) );
  AOI22_X1 U10064 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n12465), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n12511), .ZN(n8149) );
  INV_X1 U10065 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7822) );
  AOI22_X1 U10066 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(
        P1_DATAO_REG_22__SCAN_IN), .B1(n12559), .B2(n7822), .ZN(n8161) );
  INV_X1 U10067 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n12632) );
  AOI22_X1 U10068 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(
        P1_DATAO_REG_23__SCAN_IN), .B1(n12628), .B2(n12632), .ZN(n8172) );
  NAND2_X1 U10069 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n7823), .ZN(n7824) );
  INV_X1 U10070 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n14429) );
  NAND2_X1 U10071 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n14429), .ZN(n7827) );
  INV_X1 U10072 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14425) );
  INV_X1 U10073 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15095) );
  AOI22_X1 U10074 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n14425), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n15095), .ZN(n7856) );
  NAND2_X1 U10075 ( .A1(n7857), .A2(n7856), .ZN(n7829) );
  INV_X1 U10076 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9080) );
  INV_X1 U10077 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15092) );
  AOI22_X1 U10078 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n9080), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n15092), .ZN(n7830) );
  XNOR2_X1 U10079 ( .A(n8324), .B(n7830), .ZN(n13704) );
  INV_X1 U10080 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7837) );
  NAND2_X1 U10081 ( .A1(n13704), .A2(n6677), .ZN(n7842) );
  INV_X1 U10082 ( .A(SI_27_), .ZN(n13705) );
  OR2_X1 U10083 ( .A1(n13044), .A2(n13705), .ZN(n7841) );
  NAND2_X1 U10084 ( .A1(n7923), .A2(n7924), .ZN(n7939) );
  INV_X1 U10085 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n12993) );
  NAND2_X1 U10086 ( .A1(n12993), .A2(n12431), .ZN(n7843) );
  INV_X1 U10087 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n13002) );
  INV_X1 U10088 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8154) );
  INV_X1 U10089 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n9564) );
  INV_X1 U10090 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n7860) );
  NAND2_X1 U10091 ( .A1(n8198), .A2(n7860), .ZN(n7862) );
  NAND2_X1 U10092 ( .A1(n7862), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n7844) );
  NAND2_X1 U10093 ( .A1(n8261), .A2(n7844), .ZN(n13423) );
  INV_X1 U10094 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7846) );
  AND2_X2 U10095 ( .A1(n7850), .A2(n7849), .ZN(n8062) );
  NAND2_X1 U10096 ( .A1(n13423), .A2(n8328), .ZN(n7855) );
  NAND2_X2 U10097 ( .A1(n7849), .A2(n13695), .ZN(n7909) );
  AND2_X2 U10098 ( .A1(n7850), .A2(n13697), .ZN(n7966) );
  NAND2_X1 U10099 ( .A1(n11717), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n7852) );
  AND2_X2 U10100 ( .A1(n13695), .A2(n13697), .ZN(n7898) );
  NAND2_X1 U10101 ( .A1(n8346), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n7851) );
  OAI211_X1 U10102 ( .C1(n8331), .C2(n8309), .A(n7852), .B(n7851), .ZN(n7853)
         );
  INV_X1 U10103 ( .A(n7853), .ZN(n7854) );
  XNOR2_X1 U10104 ( .A(n7857), .B(n7856), .ZN(n13708) );
  NAND2_X1 U10105 ( .A1(n13708), .A2(n6676), .ZN(n7859) );
  INV_X1 U10106 ( .A(SI_26_), .ZN(n13710) );
  OR2_X1 U10107 ( .A1(n6669), .A2(n13710), .ZN(n7858) );
  OR2_X1 U10108 ( .A1(n8198), .A2(n7860), .ZN(n7861) );
  NAND2_X1 U10109 ( .A1(n7862), .A2(n7861), .ZN(n13438) );
  NAND2_X1 U10110 ( .A1(n13438), .A2(n8328), .ZN(n7867) );
  INV_X1 U10111 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13591) );
  NAND2_X1 U10112 ( .A1(n11717), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n7864) );
  NAND2_X1 U10113 ( .A1(n8346), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n7863) );
  OAI211_X1 U10114 ( .C1(n13591), .C2(n8331), .A(n7864), .B(n7863), .ZN(n7865)
         );
  INV_X1 U10115 ( .A(n7865), .ZN(n7866) );
  OR2_X1 U10116 ( .A1(n13010), .A2(n13448), .ZN(n13216) );
  NAND2_X1 U10117 ( .A1(n7966), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7871) );
  NAND2_X1 U10118 ( .A1(n8062), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7870) );
  NAND2_X1 U10119 ( .A1(n7898), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n7869) );
  INV_X1 U10120 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10639) );
  OR2_X1 U10121 ( .A1(n7909), .A2(n10639), .ZN(n7868) );
  INV_X1 U10122 ( .A(n7881), .ZN(n7873) );
  INV_X1 U10123 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8406) );
  NAND2_X1 U10124 ( .A1(n8406), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7872) );
  NAND2_X1 U10125 ( .A1(n7873), .A2(n7872), .ZN(n10707) );
  NAND2_X1 U10126 ( .A1(n6676), .A2(n10707), .ZN(n7876) );
  OR2_X1 U10127 ( .A1(n8268), .A2(n7369), .ZN(n7874) );
  NAND2_X1 U10128 ( .A1(n7966), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7880) );
  NAND2_X1 U10129 ( .A1(n8062), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7879) );
  NAND2_X1 U10130 ( .A1(n7898), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7878) );
  INV_X1 U10131 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10634) );
  OR2_X1 U10132 ( .A1(n7909), .A2(n10634), .ZN(n7877) );
  INV_X1 U10133 ( .A(SI_1_), .ZN(n10728) );
  OR2_X1 U10134 ( .A1(n6669), .A2(n10728), .ZN(n7885) );
  INV_X1 U10135 ( .A(n10614), .ZN(n7883) );
  OR2_X1 U10136 ( .A1(n8268), .A2(n11023), .ZN(n7884) );
  AND3_X2 U10137 ( .A1(n7886), .A2(n7885), .A3(n7884), .ZN(n15816) );
  NAND2_X1 U10138 ( .A1(n11400), .A2(n15816), .ZN(n13098) );
  OR2_X1 U10139 ( .A1(n11400), .A2(n15816), .ZN(n13100) );
  NAND2_X1 U10140 ( .A1(n9787), .A2(n13100), .ZN(n15786) );
  NAND2_X1 U10141 ( .A1(n7966), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7890) );
  NAND2_X1 U10142 ( .A1(n8062), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n7889) );
  NAND2_X1 U10143 ( .A1(n7898), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n7888) );
  INV_X1 U10144 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10640) );
  OR2_X1 U10145 ( .A1(n7909), .A2(n10640), .ZN(n7887) );
  INV_X1 U10146 ( .A(n7891), .ZN(n7892) );
  XNOR2_X1 U10147 ( .A(n7893), .B(n7892), .ZN(n10726) );
  NAND2_X1 U10148 ( .A1(n6677), .A2(n10726), .ZN(n7897) );
  NOR2_X1 U10149 ( .A1(n10614), .A2(n8010), .ZN(n7894) );
  OR2_X1 U10150 ( .A1(n8268), .A2(n11069), .ZN(n7896) );
  OAI211_X1 U10151 ( .C1(n6669), .C2(SI_2_), .A(n7897), .B(n7896), .ZN(n9789)
         );
  NAND2_X1 U10152 ( .A1(n15808), .A2(n9789), .ZN(n13111) );
  NAND2_X1 U10153 ( .A1(n15786), .A2(n15785), .ZN(n15784) );
  NAND2_X1 U10154 ( .A1(n15784), .A2(n13108), .ZN(n11423) );
  NAND2_X1 U10155 ( .A1(n7966), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7902) );
  INV_X1 U10156 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n11740) );
  NAND2_X1 U10157 ( .A1(n8062), .A2(n11740), .ZN(n7901) );
  NAND2_X1 U10158 ( .A1(n7898), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n7900) );
  INV_X1 U10159 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10646) );
  OR2_X1 U10160 ( .A1(n7909), .A2(n10646), .ZN(n7899) );
  INV_X1 U10161 ( .A(n7903), .ZN(n7904) );
  XNOR2_X1 U10162 ( .A(n7905), .B(n7904), .ZN(n10700) );
  NAND2_X1 U10163 ( .A1(n6676), .A2(n10700), .ZN(n7908) );
  OR2_X1 U10164 ( .A1(n8268), .A2(n10648), .ZN(n7907) );
  OAI211_X1 U10165 ( .C1(n6669), .C2(SI_3_), .A(n7908), .B(n7907), .ZN(n11547)
         );
  OR2_X1 U10166 ( .A1(n11796), .A2(n11547), .ZN(n13115) );
  NAND2_X1 U10167 ( .A1(n11796), .A2(n11547), .ZN(n13112) );
  NAND2_X1 U10168 ( .A1(n11423), .A2(n13063), .ZN(n11422) );
  NAND2_X1 U10169 ( .A1(n11422), .A2(n13115), .ZN(n11538) );
  NAND2_X1 U10170 ( .A1(n8346), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n7913) );
  NAND2_X1 U10171 ( .A1(n7966), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7912) );
  OR2_X1 U10172 ( .A1(n7760), .A2(n7923), .ZN(n11791) );
  NAND2_X1 U10173 ( .A1(n8062), .A2(n11791), .ZN(n7911) );
  INV_X1 U10174 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n11552) );
  OR2_X1 U10175 ( .A1(n7909), .A2(n11552), .ZN(n7910) );
  NAND4_X1 U10176 ( .A1(n7913), .A2(n7912), .A3(n7911), .A4(n7910), .ZN(n11427) );
  INV_X1 U10177 ( .A(n7914), .ZN(n7915) );
  XNOR2_X1 U10178 ( .A(n7916), .B(n7915), .ZN(n10705) );
  NAND2_X1 U10179 ( .A1(n6677), .A2(n10705), .ZN(n7922) );
  NAND2_X1 U10180 ( .A1(n7906), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7917) );
  MUX2_X1 U10181 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7917), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n7920) );
  INV_X1 U10182 ( .A(n7918), .ZN(n7919) );
  OR2_X1 U10183 ( .A1(n8268), .A2(n11162), .ZN(n7921) );
  OAI211_X1 U10184 ( .C1(n6669), .C2(SI_4_), .A(n7922), .B(n7921), .ZN(n12109)
         );
  NAND2_X1 U10185 ( .A1(n11427), .A2(n12109), .ZN(n13120) );
  NAND2_X1 U10186 ( .A1(n13123), .A2(n13120), .ZN(n13116) );
  INV_X1 U10187 ( .A(n13116), .ZN(n13059) );
  NAND2_X1 U10188 ( .A1(n11538), .A2(n13059), .ZN(n11537) );
  NAND2_X1 U10189 ( .A1(n8346), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n7929) );
  NAND2_X1 U10190 ( .A1(n7966), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7928) );
  OR2_X1 U10191 ( .A1(n7924), .A2(n7923), .ZN(n7925) );
  NAND2_X1 U10192 ( .A1(n7939), .A2(n7925), .ZN(n11982) );
  NAND2_X1 U10193 ( .A1(n8062), .A2(n11982), .ZN(n7927) );
  INV_X1 U10194 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10657) );
  OR2_X1 U10195 ( .A1(n7909), .A2(n10657), .ZN(n7926) );
  NAND4_X1 U10196 ( .A1(n7929), .A2(n7928), .A3(n7927), .A4(n7926), .ZN(n11628) );
  INV_X1 U10197 ( .A(n7930), .ZN(n7931) );
  XNOR2_X1 U10198 ( .A(n7932), .B(n7931), .ZN(n10702) );
  NAND2_X1 U10199 ( .A1(n6677), .A2(n10702), .ZN(n7938) );
  NOR2_X1 U10200 ( .A1(n7918), .A2(n8010), .ZN(n7933) );
  MUX2_X1 U10201 ( .A(n8010), .B(n7933), .S(P3_IR_REG_5__SCAN_IN), .Z(n7936)
         );
  INV_X1 U10202 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7934) );
  NAND2_X1 U10203 ( .A1(n7918), .A2(n7934), .ZN(n7961) );
  INV_X1 U10204 ( .A(n7961), .ZN(n7935) );
  OR2_X1 U10205 ( .A1(n8268), .A2(n11209), .ZN(n7937) );
  OAI211_X1 U10206 ( .C1(n13044), .C2(SI_5_), .A(n7938), .B(n7937), .ZN(n11979) );
  OR2_X1 U10207 ( .A1(n11628), .A2(n11979), .ZN(n13121) );
  NAND2_X1 U10208 ( .A1(n11628), .A2(n11979), .ZN(n13126) );
  NAND2_X1 U10209 ( .A1(n8346), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n7944) );
  NAND2_X1 U10210 ( .A1(n7966), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7943) );
  NAND2_X1 U10211 ( .A1(n7939), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7940) );
  NAND2_X1 U10212 ( .A1(n7952), .A2(n7940), .ZN(n12023) );
  NAND2_X1 U10213 ( .A1(n8062), .A2(n12023), .ZN(n7942) );
  INV_X1 U10214 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10661) );
  OR2_X1 U10215 ( .A1(n7909), .A2(n10661), .ZN(n7941) );
  NAND4_X1 U10216 ( .A1(n7944), .A2(n7943), .A3(n7942), .A4(n7941), .ZN(n11963) );
  XNOR2_X1 U10217 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n7945) );
  XNOR2_X1 U10218 ( .A(n7946), .B(n7945), .ZN(n10709) );
  NAND2_X1 U10219 ( .A1(n6677), .A2(n10709), .ZN(n7951) );
  INV_X1 U10220 ( .A(SI_6_), .ZN(n10710) );
  OR2_X1 U10221 ( .A1(n13044), .A2(n10710), .ZN(n7950) );
  NAND2_X1 U10222 ( .A1(n7961), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7948) );
  XNOR2_X1 U10223 ( .A(n7948), .B(n7947), .ZN(n10712) );
  OR2_X1 U10224 ( .A1(n8268), .A2(n10712), .ZN(n7949) );
  OR2_X1 U10225 ( .A1(n11963), .A2(n12030), .ZN(n13127) );
  NAND2_X1 U10226 ( .A1(n11963), .A2(n12030), .ZN(n13133) );
  NAND2_X1 U10227 ( .A1(n7966), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7958) );
  AND2_X1 U10228 ( .A1(n7952), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7953) );
  NOR2_X1 U10229 ( .A1(n7967), .A2(n7953), .ZN(n15772) );
  INV_X1 U10230 ( .A(n15772), .ZN(n7954) );
  NAND2_X1 U10231 ( .A1(n8328), .A2(n7954), .ZN(n7957) );
  NAND2_X1 U10232 ( .A1(n8346), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n7956) );
  INV_X1 U10233 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n10666) );
  OR2_X1 U10234 ( .A1(n7909), .A2(n10666), .ZN(n7955) );
  NAND4_X1 U10235 ( .A1(n7958), .A2(n7957), .A3(n7956), .A4(n7955), .ZN(n12286) );
  XNOR2_X1 U10236 ( .A(n7960), .B(n7959), .ZN(n10731) );
  NAND2_X1 U10237 ( .A1(n6676), .A2(n10731), .ZN(n7965) );
  NAND2_X1 U10238 ( .A1(n7976), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7963) );
  XNOR2_X1 U10239 ( .A(n7963), .B(n7962), .ZN(n10733) );
  INV_X1 U10240 ( .A(n10733), .ZN(n11315) );
  OR2_X1 U10241 ( .A1(n8268), .A2(n11315), .ZN(n7964) );
  OAI211_X1 U10242 ( .C1(n13044), .C2(SI_7_), .A(n7965), .B(n7964), .ZN(n12157) );
  OR2_X1 U10243 ( .A1(n12286), .A2(n12157), .ZN(n13137) );
  NAND2_X1 U10244 ( .A1(n12286), .A2(n12157), .ZN(n13136) );
  NAND2_X1 U10245 ( .A1(n13137), .A2(n13136), .ZN(n13134) );
  INV_X1 U10246 ( .A(n13134), .ZN(n13060) );
  NAND2_X1 U10247 ( .A1(n8346), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7972) );
  NAND2_X1 U10248 ( .A1(n7966), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7971) );
  NOR2_X1 U10249 ( .A1(n7967), .A2(n11407), .ZN(n7968) );
  OR2_X1 U10250 ( .A1(n7987), .A2(n7968), .ZN(n12264) );
  NAND2_X1 U10251 ( .A1(n8328), .A2(n12264), .ZN(n7970) );
  INV_X1 U10252 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n10670) );
  OR2_X1 U10253 ( .A1(n8331), .A2(n10670), .ZN(n7969) );
  NAND4_X1 U10254 ( .A1(n7972), .A2(n7971), .A3(n7970), .A4(n7969), .ZN(n13143) );
  INV_X1 U10255 ( .A(n7973), .ZN(n7974) );
  XNOR2_X1 U10256 ( .A(n7975), .B(n7974), .ZN(n10734) );
  NAND2_X1 U10257 ( .A1(n6676), .A2(n10734), .ZN(n7984) );
  NOR2_X1 U10258 ( .A1(n7976), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n7980) );
  INV_X1 U10259 ( .A(n7980), .ZN(n7977) );
  NAND2_X1 U10260 ( .A1(n7977), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7978) );
  MUX2_X1 U10261 ( .A(n7978), .B(P3_IR_REG_31__SCAN_IN), .S(n7979), .Z(n7981)
         );
  NAND2_X1 U10262 ( .A1(n7980), .A2(n7979), .ZN(n7996) );
  NAND2_X1 U10263 ( .A1(n7981), .A2(n7996), .ZN(n10737) );
  OR2_X1 U10264 ( .A1(n8268), .A2(n10737), .ZN(n7983) );
  INV_X1 U10265 ( .A(SI_8_), .ZN(n10736) );
  OR2_X1 U10266 ( .A1(n13044), .A2(n10736), .ZN(n7982) );
  XNOR2_X1 U10267 ( .A(n13143), .B(n15759), .ZN(n13144) );
  OR2_X1 U10268 ( .A1(n13143), .A2(n15759), .ZN(n7985) );
  NAND2_X1 U10269 ( .A1(n11717), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7992) );
  OR2_X1 U10270 ( .A1(n7987), .A2(n7986), .ZN(n7988) );
  NAND2_X1 U10271 ( .A1(n8001), .A2(n7988), .ZN(n12459) );
  NAND2_X1 U10272 ( .A1(n8062), .A2(n12459), .ZN(n7991) );
  NAND2_X1 U10273 ( .A1(n8346), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7990) );
  INV_X1 U10274 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n10675) );
  OR2_X1 U10275 ( .A1(n8331), .A2(n10675), .ZN(n7989) );
  NAND4_X1 U10276 ( .A1(n7992), .A2(n7991), .A3(n7990), .A4(n7989), .ZN(n13148) );
  XNOR2_X1 U10277 ( .A(n7995), .B(n7994), .ZN(n10738) );
  NAND2_X1 U10278 ( .A1(n6677), .A2(n10738), .ZN(n7999) );
  NAND2_X1 U10279 ( .A1(n7996), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7997) );
  XNOR2_X1 U10280 ( .A(n7997), .B(P3_IR_REG_9__SCAN_IN), .ZN(n10677) );
  OR2_X1 U10281 ( .A1(n8268), .A2(n10677), .ZN(n7998) );
  OR2_X1 U10282 ( .A1(n13148), .A2(n13147), .ZN(n8000) );
  NAND2_X1 U10283 ( .A1(n8346), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8006) );
  NAND2_X1 U10284 ( .A1(n11717), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8005) );
  NAND2_X1 U10285 ( .A1(n8001), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8002) );
  NAND2_X1 U10286 ( .A1(n8036), .A2(n8002), .ZN(n12514) );
  NAND2_X1 U10287 ( .A1(n8062), .A2(n12514), .ZN(n8004) );
  INV_X1 U10288 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15852) );
  OR2_X1 U10289 ( .A1(n8331), .A2(n15852), .ZN(n8003) );
  NAND4_X1 U10290 ( .A1(n8006), .A2(n8005), .A3(n8004), .A4(n8003), .ZN(n15208) );
  XNOR2_X1 U10291 ( .A(n8008), .B(n8007), .ZN(n10719) );
  NAND2_X1 U10292 ( .A1(n6677), .A2(n10719), .ZN(n8013) );
  OR2_X1 U10293 ( .A1(n8009), .A2(n8010), .ZN(n8011) );
  XNOR2_X1 U10294 ( .A(n8011), .B(P3_IR_REG_10__SCAN_IN), .ZN(n10681) );
  OR2_X1 U10295 ( .A1(n8268), .A2(n10681), .ZN(n8012) );
  OAI211_X1 U10296 ( .C1(n13044), .C2(SI_10_), .A(n8013), .B(n8012), .ZN(
        n12520) );
  NAND2_X1 U10297 ( .A1(n15208), .A2(n12520), .ZN(n13153) );
  NAND2_X1 U10298 ( .A1(n12318), .A2(n13153), .ZN(n8014) );
  OR2_X1 U10299 ( .A1(n15208), .A2(n12520), .ZN(n13154) );
  NAND2_X1 U10300 ( .A1(n8014), .A2(n13154), .ZN(n15215) );
  XNOR2_X1 U10301 ( .A(n8036), .B(P3_REG3_REG_11__SCAN_IN), .ZN(n15212) );
  NAND2_X1 U10302 ( .A1(n8062), .A2(n15212), .ZN(n8019) );
  NAND2_X1 U10303 ( .A1(n11717), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8018) );
  NAND2_X1 U10304 ( .A1(n8346), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8017) );
  INV_X1 U10305 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n8015) );
  OR2_X1 U10306 ( .A1(n8331), .A2(n8015), .ZN(n8016) );
  NAND4_X1 U10307 ( .A1(n8019), .A2(n8018), .A3(n8017), .A4(n8016), .ZN(n15198) );
  XNOR2_X1 U10308 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8020) );
  XNOR2_X1 U10309 ( .A(n8021), .B(n8020), .ZN(n10725) );
  NAND2_X1 U10310 ( .A1(n10725), .A2(n6677), .ZN(n8026) );
  NAND2_X1 U10311 ( .A1(n8009), .A2(n8022), .ZN(n8028) );
  NAND2_X1 U10312 ( .A1(n8028), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8023) );
  XNOR2_X1 U10313 ( .A(n8023), .B(P3_IR_REG_11__SCAN_IN), .ZN(n12425) );
  OAI22_X1 U10314 ( .A1(n13044), .A2(SI_11_), .B1(n12425), .B2(n10611), .ZN(
        n8024) );
  INV_X1 U10315 ( .A(n8024), .ZN(n8025) );
  NAND2_X1 U10316 ( .A1(n8026), .A2(n8025), .ZN(n15216) );
  OR2_X1 U10317 ( .A1(n15198), .A2(n15216), .ZN(n13162) );
  NAND2_X1 U10318 ( .A1(n15198), .A2(n15216), .ZN(n13165) );
  NAND2_X1 U10319 ( .A1(n15215), .A2(n15214), .ZN(n15213) );
  XNOR2_X1 U10320 ( .A(n8027), .B(n6813), .ZN(n10740) );
  NAND2_X1 U10321 ( .A1(n10740), .A2(n6676), .ZN(n8035) );
  NOR2_X1 U10322 ( .A1(n8029), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n8057) );
  INV_X1 U10323 ( .A(n8057), .ZN(n8032) );
  NAND2_X1 U10324 ( .A1(n8029), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8030) );
  MUX2_X1 U10325 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8030), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n8031) );
  NAND2_X1 U10326 ( .A1(n8032), .A2(n8031), .ZN(n13255) );
  OAI22_X1 U10327 ( .A1(n13044), .A2(n10742), .B1(n10611), .B2(n13255), .ZN(
        n8033) );
  INV_X1 U10328 ( .A(n8033), .ZN(n8034) );
  NAND2_X1 U10329 ( .A1(n8035), .A2(n8034), .ZN(n9811) );
  INV_X1 U10330 ( .A(n9811), .ZN(n15204) );
  OAI21_X1 U10331 ( .B1(n8036), .B2(P3_REG3_REG_11__SCAN_IN), .A(
        P3_REG3_REG_12__SCAN_IN), .ZN(n8037) );
  NAND2_X1 U10332 ( .A1(n8037), .A2(n8047), .ZN(n15201) );
  NAND2_X1 U10333 ( .A1(n8062), .A2(n15201), .ZN(n8041) );
  NAND2_X1 U10334 ( .A1(n8346), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8040) );
  NAND2_X1 U10335 ( .A1(n11717), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8039) );
  INV_X1 U10336 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n12413) );
  OR2_X1 U10337 ( .A1(n8331), .A2(n12413), .ZN(n8038) );
  NAND4_X1 U10338 ( .A1(n8041), .A2(n8040), .A3(n8039), .A4(n8038), .ZN(n15209) );
  NAND2_X1 U10339 ( .A1(n12994), .A2(n9811), .ZN(n13166) );
  XNOR2_X1 U10340 ( .A(n8042), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n15119) );
  NAND2_X1 U10341 ( .A1(n15119), .A2(n6677), .ZN(n8046) );
  OR2_X1 U10342 ( .A1(n8057), .A2(n8010), .ZN(n8043) );
  INV_X1 U10343 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8056) );
  XNOR2_X1 U10344 ( .A(n8043), .B(n8056), .ZN(n15124) );
  OAI22_X1 U10345 ( .A1(n13044), .A2(SI_13_), .B1(n13281), .B2(n10611), .ZN(
        n8044) );
  INV_X1 U10346 ( .A(n8044), .ZN(n8045) );
  NAND2_X1 U10347 ( .A1(n8046), .A2(n8045), .ZN(n15194) );
  NOR2_X1 U10348 ( .A1(n8063), .A2(n7768), .ZN(n15189) );
  INV_X1 U10349 ( .A(n15189), .ZN(n12979) );
  NAND2_X1 U10350 ( .A1(n8062), .A2(n12979), .ZN(n8052) );
  NAND2_X1 U10351 ( .A1(n8346), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8051) );
  NAND2_X1 U10352 ( .A1(n11717), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8050) );
  INV_X1 U10353 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n8048) );
  OR2_X1 U10354 ( .A1(n8331), .A2(n8048), .ZN(n8049) );
  NAND4_X1 U10355 ( .A1(n8052), .A2(n8051), .A3(n8050), .A4(n8049), .ZN(n15199) );
  OR2_X1 U10356 ( .A1(n15194), .A2(n15199), .ZN(n13171) );
  INV_X1 U10357 ( .A(n13171), .ZN(n8053) );
  NAND2_X1 U10358 ( .A1(n15194), .A2(n15199), .ZN(n13170) );
  XNOR2_X1 U10359 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8054) );
  XNOR2_X1 U10360 ( .A(n8055), .B(n8054), .ZN(n10848) );
  NAND2_X1 U10361 ( .A1(n10848), .A2(n6677), .ZN(n8061) );
  NAND2_X1 U10362 ( .A1(n8057), .A2(n8056), .ZN(n8071) );
  NAND2_X1 U10363 ( .A1(n8071), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8058) );
  XNOR2_X1 U10364 ( .A(n8058), .B(P3_IR_REG_14__SCAN_IN), .ZN(n13270) );
  OAI22_X1 U10365 ( .A1(n6669), .A2(SI_14_), .B1(n13270), .B2(n10611), .ZN(
        n8059) );
  INV_X1 U10366 ( .A(n8059), .ZN(n8060) );
  NAND2_X1 U10367 ( .A1(n8061), .A2(n8060), .ZN(n15178) );
  OR2_X1 U10368 ( .A1(n8063), .A2(n12883), .ZN(n8064) );
  NAND2_X1 U10369 ( .A1(n8077), .A2(n8064), .ZN(n15175) );
  NAND2_X1 U10370 ( .A1(n8328), .A2(n15175), .ZN(n8068) );
  NAND2_X1 U10371 ( .A1(n8346), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8067) );
  NAND2_X1 U10372 ( .A1(n11717), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8066) );
  INV_X1 U10373 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13269) );
  OR2_X1 U10374 ( .A1(n8331), .A2(n13269), .ZN(n8065) );
  NAND4_X1 U10375 ( .A1(n8068), .A2(n8067), .A3(n8066), .A4(n8065), .ZN(n15187) );
  NAND2_X1 U10376 ( .A1(n15178), .A2(n15187), .ZN(n8232) );
  INV_X1 U10377 ( .A(n8232), .ZN(n13175) );
  OR2_X1 U10378 ( .A1(n15178), .A2(n15187), .ZN(n13173) );
  XNOR2_X1 U10379 ( .A(n8070), .B(n8069), .ZN(n10863) );
  NAND2_X1 U10380 ( .A1(n10863), .A2(n6676), .ZN(n8076) );
  OAI21_X1 U10381 ( .B1(n8071), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8073) );
  INV_X1 U10382 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8072) );
  INV_X1 U10383 ( .A(n15146), .ZN(n13308) );
  OAI22_X1 U10384 ( .A1(n13044), .A2(SI_15_), .B1(n13308), .B2(n10611), .ZN(
        n8074) );
  INV_X1 U10385 ( .A(n8074), .ZN(n8075) );
  NAND2_X1 U10386 ( .A1(n7898), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8082) );
  NAND2_X1 U10387 ( .A1(n11717), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8081) );
  NAND2_X1 U10388 ( .A1(n8077), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8078) );
  NAND2_X1 U10389 ( .A1(n8093), .A2(n8078), .ZN(n13032) );
  NAND2_X1 U10390 ( .A1(n8328), .A2(n13032), .ZN(n8080) );
  INV_X1 U10391 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n15149) );
  OR2_X1 U10392 ( .A1(n8331), .A2(n15149), .ZN(n8079) );
  NAND4_X1 U10393 ( .A1(n8082), .A2(n8081), .A3(n8080), .A4(n8079), .ZN(n15173) );
  XNOR2_X1 U10394 ( .A(n13179), .B(n15173), .ZN(n13176) );
  NAND2_X1 U10395 ( .A1(n12635), .A2(n12636), .ZN(n8083) );
  OR2_X1 U10396 ( .A1(n13179), .A2(n15173), .ZN(n13185) );
  INV_X1 U10397 ( .A(n8084), .ZN(n8085) );
  XNOR2_X1 U10398 ( .A(n8086), .B(n8085), .ZN(n10973) );
  NAND2_X1 U10399 ( .A1(n10973), .A2(n6677), .ZN(n8092) );
  NAND2_X1 U10400 ( .A1(n6972), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8088) );
  MUX2_X1 U10401 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8088), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n8089) );
  NAND2_X1 U10402 ( .A1(n8089), .A2(n8102), .ZN(n13333) );
  OAI22_X1 U10403 ( .A1(n13044), .A2(n10975), .B1(n10611), .B2(n13333), .ZN(
        n8090) );
  INV_X1 U10404 ( .A(n8090), .ZN(n8091) );
  NAND2_X1 U10405 ( .A1(n7898), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8099) );
  NAND2_X1 U10406 ( .A1(n11717), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8098) );
  INV_X1 U10407 ( .A(n8109), .ZN(n8095) );
  NAND2_X1 U10408 ( .A1(n8093), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8094) );
  NAND2_X1 U10409 ( .A1(n8095), .A2(n8094), .ZN(n13581) );
  NAND2_X1 U10410 ( .A1(n8328), .A2(n13581), .ZN(n8097) );
  INV_X1 U10411 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13310) );
  OR2_X1 U10412 ( .A1(n8331), .A2(n13310), .ZN(n8096) );
  NAND4_X1 U10413 ( .A1(n8099), .A2(n8098), .A3(n8097), .A4(n8096), .ZN(n13559) );
  INV_X1 U10414 ( .A(n13559), .ZN(n12947) );
  OR2_X1 U10415 ( .A1(n13681), .A2(n12947), .ZN(n13187) );
  XNOR2_X1 U10416 ( .A(n8101), .B(n8100), .ZN(n10976) );
  NAND2_X1 U10417 ( .A1(n10976), .A2(n6676), .ZN(n8108) );
  NAND2_X1 U10418 ( .A1(n8102), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8104) );
  MUX2_X1 U10419 ( .A(n8104), .B(P3_IR_REG_31__SCAN_IN), .S(n8103), .Z(n8105)
         );
  NAND2_X1 U10420 ( .A1(n8105), .A2(n6701), .ZN(n13361) );
  INV_X1 U10421 ( .A(n13361), .ZN(n13348) );
  OAI22_X1 U10422 ( .A1(n13044), .A2(SI_17_), .B1(n13348), .B2(n10611), .ZN(
        n8106) );
  INV_X1 U10423 ( .A(n8106), .ZN(n8107) );
  NAND2_X1 U10424 ( .A1(n7898), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8114) );
  NAND2_X1 U10425 ( .A1(n11717), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8113) );
  NOR2_X1 U10426 ( .A1(n8109), .A2(n12944), .ZN(n8110) );
  OR2_X1 U10427 ( .A1(n8123), .A2(n8110), .ZN(n13566) );
  NAND2_X1 U10428 ( .A1(n8328), .A2(n13566), .ZN(n8112) );
  INV_X1 U10429 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13332) );
  OR2_X1 U10430 ( .A1(n8331), .A2(n13332), .ZN(n8111) );
  NAND4_X1 U10431 ( .A1(n8114), .A2(n8113), .A3(n8112), .A4(n8111), .ZN(n13574) );
  XNOR2_X1 U10432 ( .A(n13568), .B(n13546), .ZN(n13564) );
  OR2_X1 U10433 ( .A1(n13568), .A2(n13574), .ZN(n13093) );
  INV_X1 U10434 ( .A(n8115), .ZN(n8116) );
  XNOR2_X1 U10435 ( .A(n8117), .B(n8116), .ZN(n11181) );
  NAND2_X1 U10436 ( .A1(n11181), .A2(n6676), .ZN(n8122) );
  NAND2_X1 U10437 ( .A1(n6701), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8119) );
  XNOR2_X1 U10438 ( .A(n8119), .B(n8118), .ZN(n13380) );
  OAI22_X1 U10439 ( .A1(n13044), .A2(n11183), .B1(n10611), .B2(n13380), .ZN(
        n8120) );
  INV_X1 U10440 ( .A(n8120), .ZN(n8121) );
  NAND2_X1 U10441 ( .A1(n8346), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8128) );
  NAND2_X1 U10442 ( .A1(n11717), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8127) );
  OR2_X1 U10443 ( .A1(n8123), .A2(n13002), .ZN(n8124) );
  NAND2_X1 U10444 ( .A1(n8135), .A2(n8124), .ZN(n13551) );
  NAND2_X1 U10445 ( .A1(n8328), .A2(n13551), .ZN(n8126) );
  INV_X1 U10446 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13624) );
  OR2_X1 U10447 ( .A1(n8331), .A2(n13624), .ZN(n8125) );
  NAND4_X1 U10448 ( .A1(n8128), .A2(n8127), .A3(n8126), .A4(n8125), .ZN(n13560) );
  INV_X1 U10449 ( .A(n13560), .ZN(n12897) );
  NAND2_X1 U10450 ( .A1(n13550), .A2(n12897), .ZN(n13092) );
  NAND2_X1 U10451 ( .A1(n13088), .A2(n13092), .ZN(n13094) );
  INV_X1 U10452 ( .A(n8129), .ZN(n8130) );
  XNOR2_X1 U10453 ( .A(n8131), .B(n8130), .ZN(n11253) );
  NAND2_X1 U10454 ( .A1(n11253), .A2(n6677), .ZN(n8134) );
  INV_X1 U10455 ( .A(SI_19_), .ZN(n11254) );
  OAI22_X1 U10456 ( .A1(n13044), .A2(n11254), .B1(n10611), .B2(n13393), .ZN(
        n8132) );
  INV_X1 U10457 ( .A(n8132), .ZN(n8133) );
  NAND2_X1 U10458 ( .A1(n8135), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8136) );
  NAND2_X1 U10459 ( .A1(n8144), .A2(n8136), .ZN(n13537) );
  NAND2_X1 U10460 ( .A1(n13537), .A2(n8328), .ZN(n8141) );
  NAND2_X1 U10461 ( .A1(n8346), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8140) );
  NAND2_X1 U10462 ( .A1(n11717), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8139) );
  INV_X1 U10463 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n8137) );
  OR2_X1 U10464 ( .A1(n8331), .A2(n8137), .ZN(n8138) );
  NAND4_X1 U10465 ( .A1(n8141), .A2(n8140), .A3(n8139), .A4(n8138), .ZN(n13518) );
  OR2_X1 U10466 ( .A1(n13671), .A2(n13547), .ZN(n13091) );
  INV_X1 U10467 ( .A(n13091), .ZN(n13192) );
  NAND2_X1 U10468 ( .A1(n13671), .A2(n13547), .ZN(n13191) );
  XNOR2_X1 U10469 ( .A(n8142), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n11660) );
  NOR2_X1 U10470 ( .A1(n6669), .A2(n11661), .ZN(n8143) );
  INV_X1 U10471 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n8148) );
  AND2_X1 U10472 ( .A1(n8144), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8145) );
  OR2_X1 U10473 ( .A1(n8145), .A2(n8155), .ZN(n13526) );
  NAND2_X1 U10474 ( .A1(n13526), .A2(n8328), .ZN(n8147) );
  AOI22_X1 U10475 ( .A1(n11717), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n8346), 
        .B2(P3_REG0_REG_20__SCAN_IN), .ZN(n8146) );
  OAI211_X1 U10476 ( .C1(n8331), .C2(n8148), .A(n8147), .B(n8146), .ZN(n13532)
         );
  NAND2_X1 U10477 ( .A1(n13528), .A2(n13532), .ZN(n13197) );
  INV_X1 U10478 ( .A(n13528), .ZN(n13613) );
  INV_X1 U10479 ( .A(n13532), .ZN(n13508) );
  NAND2_X1 U10480 ( .A1(n13613), .A2(n13508), .ZN(n13198) );
  INV_X1 U10481 ( .A(n8149), .ZN(n8150) );
  XNOR2_X1 U10482 ( .A(n8151), .B(n8150), .ZN(n11787) );
  NAND2_X1 U10483 ( .A1(n11787), .A2(n6677), .ZN(n8153) );
  INV_X1 U10484 ( .A(SI_21_), .ZN(n11789) );
  OR2_X1 U10485 ( .A1(n13044), .A2(n11789), .ZN(n8152) );
  NOR2_X1 U10486 ( .A1(n8155), .A2(n8154), .ZN(n8156) );
  OR2_X1 U10487 ( .A1(n8165), .A2(n8156), .ZN(n13511) );
  NAND2_X1 U10488 ( .A1(n13511), .A2(n8328), .ZN(n8160) );
  INV_X1 U10489 ( .A(n8331), .ZN(n8157) );
  AOI22_X1 U10490 ( .A1(n8157), .A2(P3_REG1_REG_21__SCAN_IN), .B1(n11717), 
        .B2(P3_REG2_REG_21__SCAN_IN), .ZN(n8159) );
  NAND2_X1 U10491 ( .A1(n8346), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8158) );
  INV_X1 U10492 ( .A(n13086), .ZN(n13667) );
  XNOR2_X1 U10493 ( .A(n8162), .B(n8161), .ZN(n11956) );
  NAND2_X1 U10494 ( .A1(n11956), .A2(n6676), .ZN(n8164) );
  OR2_X1 U10495 ( .A1(n13044), .A2(n7180), .ZN(n8163) );
  OR2_X1 U10496 ( .A1(n8165), .A2(n9564), .ZN(n8166) );
  NAND2_X1 U10497 ( .A1(n8176), .A2(n8166), .ZN(n13500) );
  NAND2_X1 U10498 ( .A1(n13500), .A2(n8328), .ZN(n8171) );
  INV_X1 U10499 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13607) );
  NAND2_X1 U10500 ( .A1(n8346), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8168) );
  NAND2_X1 U10501 ( .A1(n11717), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8167) );
  OAI211_X1 U10502 ( .C1(n13607), .C2(n8331), .A(n8168), .B(n8167), .ZN(n8169)
         );
  INV_X1 U10503 ( .A(n8169), .ZN(n8170) );
  NAND2_X1 U10504 ( .A1(n13499), .A2(n13507), .ZN(n13202) );
  XNOR2_X1 U10505 ( .A(n8173), .B(n8172), .ZN(n12175) );
  NAND2_X1 U10506 ( .A1(n12175), .A2(n6677), .ZN(n8175) );
  INV_X1 U10507 ( .A(SI_23_), .ZN(n12177) );
  OR2_X1 U10508 ( .A1(n6669), .A2(n12177), .ZN(n8174) );
  NAND2_X1 U10509 ( .A1(n8176), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8177) );
  NAND2_X1 U10510 ( .A1(n8186), .A2(n8177), .ZN(n13488) );
  NAND2_X1 U10511 ( .A1(n13488), .A2(n8328), .ZN(n8182) );
  INV_X1 U10512 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13603) );
  NAND2_X1 U10513 ( .A1(n8346), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8179) );
  NAND2_X1 U10514 ( .A1(n11717), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8178) );
  OAI211_X1 U10515 ( .C1(n13603), .C2(n8331), .A(n8179), .B(n8178), .ZN(n8180)
         );
  INV_X1 U10516 ( .A(n8180), .ZN(n8181) );
  INV_X1 U10517 ( .A(n13466), .ZN(n13495) );
  NAND2_X1 U10518 ( .A1(n12713), .A2(n13495), .ZN(n13207) );
  INV_X1 U10519 ( .A(n13481), .ZN(n13476) );
  INV_X1 U10520 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n15102) );
  INV_X1 U10521 ( .A(SI_24_), .ZN(n12498) );
  OR2_X1 U10522 ( .A1(n13044), .A2(n12498), .ZN(n8184) );
  NAND2_X1 U10523 ( .A1(n8186), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8187) );
  NAND2_X1 U10524 ( .A1(n8199), .A2(n8187), .ZN(n13471) );
  NAND2_X1 U10525 ( .A1(n13471), .A2(n8328), .ZN(n8192) );
  INV_X1 U10526 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13599) );
  NAND2_X1 U10527 ( .A1(n11717), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8189) );
  NAND2_X1 U10528 ( .A1(n8346), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8188) );
  OAI211_X1 U10529 ( .C1(n8331), .C2(n13599), .A(n8189), .B(n8188), .ZN(n8190)
         );
  INV_X1 U10530 ( .A(n8190), .ZN(n8191) );
  NAND2_X1 U10531 ( .A1(n13459), .A2(n13460), .ZN(n13213) );
  INV_X1 U10532 ( .A(n13213), .ZN(n8193) );
  INV_X1 U10533 ( .A(n13483), .ZN(n13447) );
  NAND2_X1 U10534 ( .A1(n12951), .A2(n13447), .ZN(n13083) );
  AOI22_X1 U10535 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .B1(n14429), .B2(n15098), .ZN(n8194) );
  XNOR2_X1 U10536 ( .A(n8195), .B(n8194), .ZN(n13714) );
  NAND2_X1 U10537 ( .A1(n13714), .A2(n6676), .ZN(n8197) );
  INV_X1 U10538 ( .A(SI_25_), .ZN(n13716) );
  OR2_X1 U10539 ( .A1(n13044), .A2(n13716), .ZN(n8196) );
  INV_X1 U10540 ( .A(n8198), .ZN(n8201) );
  NAND2_X1 U10541 ( .A1(n8199), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8200) );
  NAND2_X1 U10542 ( .A1(n8201), .A2(n8200), .ZN(n13453) );
  NAND2_X1 U10543 ( .A1(n13453), .A2(n8328), .ZN(n8206) );
  INV_X1 U10544 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13595) );
  NAND2_X1 U10545 ( .A1(n8346), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8203) );
  NAND2_X1 U10546 ( .A1(n11717), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8202) );
  OAI211_X1 U10547 ( .C1(n13595), .C2(n8331), .A(n8203), .B(n8202), .ZN(n8204)
         );
  INV_X1 U10548 ( .A(n8204), .ZN(n8205) );
  OR2_X1 U10549 ( .A1(n12920), .A2(n13433), .ZN(n13218) );
  NAND2_X1 U10550 ( .A1(n12920), .A2(n13433), .ZN(n13215) );
  NAND2_X1 U10551 ( .A1(n13010), .A2(n13448), .ZN(n13219) );
  INV_X1 U10552 ( .A(n6721), .ZN(n8209) );
  OR2_X1 U10553 ( .A1(n8207), .A2(n13223), .ZN(n8208) );
  NAND2_X1 U10554 ( .A1(n6720), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8210) );
  MUX2_X1 U10555 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8210), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n8211) );
  NOR2_X1 U10556 ( .A1(n11663), .A2(n11788), .ZN(n13239) );
  NOR2_X1 U10557 ( .A1(n8258), .A2(n13393), .ZN(n8312) );
  NAND2_X1 U10558 ( .A1(n13100), .A2(n13098), .ZN(n11259) );
  NAND2_X1 U10559 ( .A1(n15807), .A2(n11467), .ZN(n15805) );
  NAND2_X1 U10560 ( .A1(n11259), .A2(n15805), .ZN(n8213) );
  OR2_X1 U10561 ( .A1(n11400), .A2(n9783), .ZN(n8212) );
  NAND2_X1 U10562 ( .A1(n15783), .A2(n8214), .ZN(n11425) );
  INV_X1 U10563 ( .A(n9789), .ZN(n15797) );
  OR2_X1 U10564 ( .A1(n15808), .A2(n15797), .ZN(n11424) );
  INV_X1 U10565 ( .A(n11547), .ZN(n15779) );
  NAND2_X1 U10566 ( .A1(n11796), .A2(n15779), .ZN(n8216) );
  NAND2_X1 U10567 ( .A1(n11429), .A2(n8216), .ZN(n11539) );
  INV_X1 U10568 ( .A(n12109), .ZN(n8217) );
  NAND2_X1 U10569 ( .A1(n11427), .A2(n8217), .ZN(n8218) );
  INV_X1 U10570 ( .A(n11979), .ZN(n8219) );
  OR2_X1 U10571 ( .A1(n11628), .A2(n8219), .ZN(n8220) );
  INV_X1 U10572 ( .A(n12030), .ZN(n11847) );
  NAND2_X1 U10573 ( .A1(n11963), .A2(n11847), .ZN(n8222) );
  INV_X1 U10574 ( .A(n12157), .ZN(n15770) );
  NAND2_X1 U10575 ( .A1(n12286), .A2(n15770), .ZN(n8223) );
  INV_X1 U10576 ( .A(n15759), .ZN(n12289) );
  OR2_X1 U10577 ( .A1(n13143), .A2(n12289), .ZN(n8224) );
  INV_X1 U10578 ( .A(n13147), .ZN(n12458) );
  XNOR2_X1 U10579 ( .A(n13148), .B(n12458), .ZN(n13066) );
  NAND2_X1 U10580 ( .A1(n13154), .A2(n13153), .ZN(n13151) );
  INV_X1 U10581 ( .A(n12520), .ZN(n8225) );
  NAND2_X1 U10582 ( .A1(n15208), .A2(n8225), .ZN(n8226) );
  INV_X1 U10583 ( .A(n15216), .ZN(n8228) );
  OR2_X1 U10584 ( .A1(n15198), .A2(n8228), .ZN(n8227) );
  NAND2_X1 U10585 ( .A1(n15207), .A2(n8227), .ZN(n15182) );
  NAND2_X1 U10586 ( .A1(n15198), .A2(n8228), .ZN(n15181) );
  NAND2_X1 U10587 ( .A1(n9811), .A2(n15209), .ZN(n15184) );
  INV_X1 U10588 ( .A(n15199), .ZN(n12885) );
  OR2_X1 U10589 ( .A1(n15194), .A2(n12885), .ZN(n8233) );
  AND2_X1 U10590 ( .A1(n15184), .A2(n8233), .ZN(n8229) );
  AND2_X1 U10591 ( .A1(n15181), .A2(n8229), .ZN(n8231) );
  INV_X1 U10592 ( .A(n8229), .ZN(n8230) );
  INV_X1 U10593 ( .A(n15202), .ZN(n15183) );
  NAND2_X1 U10594 ( .A1(n13173), .A2(n8232), .ZN(n15176) );
  INV_X1 U10595 ( .A(n8233), .ZN(n8234) );
  NAND2_X1 U10596 ( .A1(n13171), .A2(n13170), .ZN(n15193) );
  OR2_X1 U10597 ( .A1(n8234), .A2(n15193), .ZN(n15170) );
  AND2_X1 U10598 ( .A1(n15176), .A2(n15170), .ZN(n8235) );
  INV_X1 U10599 ( .A(n15187), .ZN(n13029) );
  OR2_X1 U10600 ( .A1(n15178), .A2(n13029), .ZN(n8236) );
  INV_X1 U10601 ( .A(n15173), .ZN(n13180) );
  NOR2_X1 U10602 ( .A1(n13179), .A2(n13180), .ZN(n8239) );
  NAND2_X1 U10603 ( .A1(n13179), .A2(n13180), .ZN(n8238) );
  NAND2_X1 U10604 ( .A1(n13681), .A2(n13559), .ZN(n8241) );
  NAND2_X1 U10605 ( .A1(n13573), .A2(n8241), .ZN(n13557) );
  INV_X1 U10606 ( .A(n13564), .ZN(n13558) );
  OR2_X1 U10607 ( .A1(n13568), .A2(n13546), .ZN(n8242) );
  NAND2_X1 U10608 ( .A1(n13556), .A2(n8242), .ZN(n13544) );
  OR2_X1 U10609 ( .A1(n13550), .A2(n13560), .ZN(n8243) );
  NAND2_X1 U10610 ( .A1(n13091), .A2(n13191), .ZN(n13535) );
  NAND2_X1 U10611 ( .A1(n13671), .A2(n13518), .ZN(n8244) );
  NAND2_X1 U10612 ( .A1(n13613), .A2(n13532), .ZN(n8245) );
  NAND2_X1 U10613 ( .A1(n13516), .A2(n8245), .ZN(n13505) );
  OR2_X1 U10614 ( .A1(n13086), .A2(n13519), .ZN(n8246) );
  NAND2_X1 U10615 ( .A1(n13086), .A2(n13519), .ZN(n8247) );
  NAND2_X1 U10616 ( .A1(n12713), .A2(n13466), .ZN(n8249) );
  INV_X1 U10617 ( .A(n13459), .ZN(n13464) );
  NAND2_X1 U10618 ( .A1(n12951), .A2(n13483), .ZN(n8250) );
  NAND2_X1 U10619 ( .A1(n13463), .A2(n8250), .ZN(n13446) );
  NAND2_X1 U10620 ( .A1(n12920), .A2(n13467), .ZN(n8251) );
  OR2_X1 U10621 ( .A1(n13010), .A2(n11520), .ZN(n8252) );
  INV_X1 U10622 ( .A(n13223), .ZN(n13077) );
  XNOR2_X1 U10623 ( .A(n8339), .B(n13077), .ZN(n8271) );
  NAND2_X1 U10624 ( .A1(n11663), .A2(n13243), .ZN(n8253) );
  NAND2_X1 U10625 ( .A1(n8253), .A2(n13081), .ZN(n8254) );
  NAND2_X1 U10626 ( .A1(n8254), .A2(n11788), .ZN(n8257) );
  NAND2_X1 U10627 ( .A1(n11663), .A2(n11788), .ZN(n8255) );
  NAND2_X1 U10628 ( .A1(n8255), .A2(n8258), .ZN(n8256) );
  NAND2_X1 U10629 ( .A1(n8257), .A2(n8256), .ZN(n9864) );
  NAND2_X1 U10630 ( .A1(n8258), .A2(n11788), .ZN(n15815) );
  NAND2_X1 U10631 ( .A1(n11663), .A2(n13393), .ZN(n13236) );
  NOR2_X1 U10632 ( .A1(n15796), .A2(n13236), .ZN(n8259) );
  NAND2_X1 U10633 ( .A1(n9864), .A2(n8259), .ZN(n8260) );
  NAND2_X1 U10634 ( .A1(n13393), .A2(n13243), .ZN(n8302) );
  OR2_X1 U10635 ( .A1(n8302), .A2(n11663), .ZN(n8304) );
  NAND2_X1 U10636 ( .A1(n8260), .A2(n8304), .ZN(n15814) );
  AND2_X1 U10637 ( .A1(n8261), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8262) );
  INV_X1 U10638 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13588) );
  NAND2_X1 U10639 ( .A1(n11717), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8264) );
  NAND2_X1 U10640 ( .A1(n8346), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8263) );
  OAI211_X1 U10641 ( .C1(n13588), .C2(n8331), .A(n8264), .B(n8263), .ZN(n8265)
         );
  OR2_X1 U10642 ( .A1(n8266), .A2(n10612), .ZN(n10632) );
  NAND2_X2 U10643 ( .A1(n13243), .A2(n13105), .ZN(n13228) );
  OAI22_X1 U10644 ( .A1(n9880), .A2(n15787), .B1(n13448), .B2(n15789), .ZN(
        n8269) );
  AOI21_X1 U10645 ( .B1(n13427), .B2(n15814), .A(n8269), .ZN(n8270) );
  OAI21_X1 U10646 ( .B1(n15811), .B2(n8271), .A(n8270), .ZN(n13422) );
  AOI21_X1 U10647 ( .B1(n15842), .B2(n13427), .A(n13422), .ZN(n8320) );
  NAND2_X1 U10648 ( .A1(n8275), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8274) );
  INV_X1 U10649 ( .A(P3_B_REG_SCAN_IN), .ZN(n8344) );
  XNOR2_X1 U10650 ( .A(n12496), .B(n8344), .ZN(n8278) );
  INV_X1 U10651 ( .A(n8282), .ZN(n13718) );
  NAND2_X1 U10652 ( .A1(n8278), .A2(n13718), .ZN(n8281) );
  INV_X1 U10653 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n10987) );
  NAND2_X1 U10654 ( .A1(n8293), .A2(n10987), .ZN(n8283) );
  OR2_X1 U10655 ( .A1(n13707), .A2(n8282), .ZN(n10985) );
  INV_X1 U10656 ( .A(n9778), .ZN(n13686) );
  AND2_X1 U10657 ( .A1(n11461), .A2(n13686), .ZN(n8311) );
  NOR2_X1 U10658 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n8288) );
  NOR4_X1 U10659 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8287) );
  NOR4_X1 U10660 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n8286) );
  NOR4_X1 U10661 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8285) );
  NAND4_X1 U10662 ( .A1(n8288), .A2(n8287), .A3(n8286), .A4(n8285), .ZN(n8295)
         );
  NOR4_X1 U10663 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n8292) );
  NOR4_X1 U10664 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n8291) );
  NOR4_X1 U10665 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8290) );
  NOR4_X1 U10666 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8289) );
  NAND4_X1 U10667 ( .A1(n8292), .A2(n8291), .A3(n8290), .A4(n8289), .ZN(n8294)
         );
  NAND2_X1 U10668 ( .A1(n8296), .A2(n13707), .ZN(n10588) );
  NAND2_X1 U10669 ( .A1(n8272), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8298) );
  XNOR2_X1 U10670 ( .A(n8298), .B(n8297), .ZN(n9874) );
  INV_X1 U10671 ( .A(n10608), .ZN(n9860) );
  NAND2_X1 U10672 ( .A1(n8314), .A2(n9860), .ZN(n8299) );
  NOR2_X1 U10673 ( .A1(n8311), .A2(n8299), .ZN(n8301) );
  INV_X1 U10674 ( .A(n11461), .ZN(n8300) );
  NAND2_X1 U10675 ( .A1(n9778), .A2(n8300), .ZN(n8316) );
  OAI21_X1 U10676 ( .B1(n6971), .B2(n15815), .A(n8302), .ZN(n8303) );
  AOI21_X1 U10677 ( .B1(n8303), .B2(n13236), .A(n13221), .ZN(n8306) );
  NAND2_X1 U10678 ( .A1(n8304), .A2(n13228), .ZN(n11458) );
  NAND2_X1 U10679 ( .A1(n13236), .A2(n13221), .ZN(n9868) );
  NAND2_X1 U10680 ( .A1(n11458), .A2(n9868), .ZN(n11457) );
  NAND2_X1 U10681 ( .A1(n11461), .A2(n11457), .ZN(n8305) );
  OAI21_X1 U10682 ( .B1(n11461), .B2(n8306), .A(n8305), .ZN(n8307) );
  INV_X1 U10683 ( .A(n8307), .ZN(n8308) );
  MUX2_X1 U10684 ( .A(n8309), .B(n8320), .S(n15854), .Z(n8310) );
  NAND2_X1 U10685 ( .A1(n8310), .A2(n7749), .ZN(P3_U3486) );
  INV_X1 U10686 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n8321) );
  NAND2_X1 U10687 ( .A1(n8311), .A2(n8314), .ZN(n9865) );
  INV_X1 U10688 ( .A(n13238), .ZN(n8313) );
  NAND2_X1 U10689 ( .A1(n8313), .A2(n8312), .ZN(n9866) );
  OR2_X1 U10690 ( .A1(n13236), .A2(n13228), .ZN(n11235) );
  AND2_X1 U10691 ( .A1(n9866), .A2(n11235), .ZN(n8318) );
  INV_X1 U10692 ( .A(n8314), .ZN(n8315) );
  INV_X1 U10693 ( .A(n9864), .ZN(n8317) );
  OAI22_X1 U10694 ( .A1(n9865), .A2(n8318), .B1(n9876), .B2(n8317), .ZN(n8319)
         );
  MUX2_X1 U10695 ( .A(n8321), .B(n8320), .S(n15846), .Z(n8322) );
  NAND2_X1 U10696 ( .A1(n8322), .A2(n7748), .ZN(P3_U3454) );
  INV_X1 U10697 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12716) );
  INV_X1 U10698 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14418) );
  NAND2_X1 U10699 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n14418), .ZN(n8325) );
  NOR2_X1 U10700 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n15092), .ZN(n8323) );
  INV_X1 U10701 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14411) );
  INV_X1 U10702 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n12861) );
  AOI22_X1 U10703 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n14411), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n12861), .ZN(n13036) );
  XNOR2_X1 U10704 ( .A(n13037), .B(n13036), .ZN(n13696) );
  NAND2_X1 U10705 ( .A1(n13696), .A2(n6677), .ZN(n8327) );
  INV_X1 U10706 ( .A(SI_29_), .ZN(n13699) );
  OR2_X1 U10707 ( .A1(n13044), .A2(n13699), .ZN(n8326) );
  NAND2_X1 U10708 ( .A1(n15162), .A2(n8328), .ZN(n11723) );
  INV_X1 U10709 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8360) );
  NAND2_X1 U10710 ( .A1(n7966), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8330) );
  NAND2_X1 U10711 ( .A1(n8346), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8329) );
  OAI211_X1 U10712 ( .C1(n8331), .C2(n8360), .A(n8330), .B(n8329), .ZN(n8332)
         );
  INV_X1 U10713 ( .A(n8332), .ZN(n8333) );
  XNOR2_X1 U10714 ( .A(n13053), .B(n13411), .ZN(n13079) );
  AOI22_X1 U10715 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n14418), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n12716), .ZN(n8334) );
  INV_X1 U10716 ( .A(n8334), .ZN(n8335) );
  XNOR2_X1 U10717 ( .A(n8336), .B(n8335), .ZN(n13700) );
  NAND2_X1 U10718 ( .A1(n13700), .A2(n6677), .ZN(n8338) );
  INV_X1 U10719 ( .A(SI_28_), .ZN(n13701) );
  OR2_X1 U10720 ( .A1(n13044), .A2(n13701), .ZN(n8337) );
  NAND2_X1 U10721 ( .A1(n13415), .A2(n9880), .ZN(n8340) );
  INV_X1 U10722 ( .A(n12868), .ZN(n13434) );
  NAND2_X1 U10723 ( .A1(n13224), .A2(n13434), .ZN(n13405) );
  NAND2_X1 U10724 ( .A1(n8340), .A2(n13405), .ZN(n13226) );
  XNOR2_X1 U10725 ( .A(n13079), .B(n13056), .ZN(n13402) );
  INV_X1 U10726 ( .A(n9880), .ZN(n11821) );
  XNOR2_X1 U10727 ( .A(n8343), .B(n8342), .ZN(n8354) );
  OR2_X1 U10728 ( .A1(n8266), .A2(n8344), .ZN(n8345) );
  NAND2_X1 U10729 ( .A1(n15809), .A2(n8345), .ZN(n15160) );
  INV_X1 U10730 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n8349) );
  NAND2_X1 U10731 ( .A1(n8346), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8348) );
  NAND2_X1 U10732 ( .A1(n11717), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8347) );
  OAI211_X1 U10733 ( .C1(n8349), .C2(n7909), .A(n8348), .B(n8347), .ZN(n8350)
         );
  INV_X1 U10734 ( .A(n8350), .ZN(n8351) );
  AND2_X1 U10735 ( .A1(n11723), .A2(n8351), .ZN(n13051) );
  OAI22_X1 U10736 ( .A1(n9880), .A2(n15789), .B1(n15160), .B2(n13051), .ZN(
        n8352) );
  INV_X1 U10737 ( .A(n8352), .ZN(n8353) );
  INV_X1 U10738 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8356) );
  OR2_X1 U10739 ( .A1(n15846), .A2(n8356), .ZN(n8357) );
  OAI21_X1 U10740 ( .B1(n8364), .B2(n15844), .A(n8359), .ZN(P3_U3456) );
  OR2_X1 U10741 ( .A1(n15854), .A2(n8360), .ZN(n8361) );
  INV_X1 U10742 ( .A(n8362), .ZN(n8363) );
  OAI21_X1 U10743 ( .B1(n8364), .B2(n15851), .A(n8363), .ZN(P3_U3488) );
  INV_X1 U10744 ( .A(n8836), .ZN(n8367) );
  AND2_X1 U10745 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n8368) );
  NAND2_X1 U10746 ( .A1(n8384), .A2(n8368), .ZN(n8373) );
  INV_X1 U10747 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8371) );
  NAND2_X1 U10748 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n8369) );
  NAND2_X1 U10749 ( .A1(n8369), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8370) );
  OAI21_X1 U10750 ( .B1(n8371), .B2(P2_IR_REG_31__SCAN_IN), .A(n8370), .ZN(
        n8372) );
  INV_X1 U10751 ( .A(n8379), .ZN(n8375) );
  NAND2_X1 U10752 ( .A1(n8375), .A2(n6927), .ZN(n8376) );
  NAND2_X1 U10753 ( .A1(n8376), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8378) );
  NAND2_X1 U10754 ( .A1(n9747), .A2(n14272), .ZN(n9739) );
  NAND2_X1 U10755 ( .A1(n8375), .A2(n6787), .ZN(n8380) );
  NAND2_X1 U10756 ( .A1(n8380), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8382) );
  INV_X1 U10757 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8381) );
  NAND2_X1 U10758 ( .A1(n8384), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8383) );
  MUX2_X1 U10759 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8383), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n8387) );
  INV_X1 U10760 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8385) );
  OAI211_X1 U10761 ( .C1(n9739), .C2(n10963), .A(n9748), .B(n9773), .ZN(n9108)
         );
  NOR2_X1 U10762 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n8390) );
  NOR2_X1 U10763 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n8389) );
  NAND4_X1 U10764 ( .A1(n8391), .A2(n8390), .A3(n8389), .A4(n8388), .ZN(n8392)
         );
  INV_X1 U10765 ( .A(n8411), .ZN(n8397) );
  NAND2_X1 U10766 ( .A1(n8395), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8396) );
  INV_X1 U10767 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n8402) );
  NAND2_X1 U10768 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n15565), .ZN(n8401) );
  XNOR2_X1 U10769 ( .A(n8402), .B(n8401), .ZN(n15562) );
  NAND2_X1 U10770 ( .A1(n8408), .A2(n7186), .ZN(n8409) );
  NAND2_X1 U10771 ( .A1(n8438), .A2(n8409), .ZN(n10722) );
  NAND2_X1 U10772 ( .A1(n8582), .A2(n9178), .ZN(n8423) );
  INV_X1 U10773 ( .A(n8415), .ZN(n8417) );
  NAND2_X1 U10774 ( .A1(n8464), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8421) );
  AND2_X4 U10775 ( .A1(n8415), .A2(n8416), .ZN(n8514) );
  NAND2_X1 U10776 ( .A1(n8514), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8420) );
  NAND2_X1 U10777 ( .A1(n8513), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8419) );
  NAND4_X2 U10778 ( .A1(n8421), .A2(n8420), .A3(n8419), .A4(n8418), .ZN(n9686)
         );
  NAND2_X1 U10779 ( .A1(n9686), .A2(n6673), .ZN(n8422) );
  NAND2_X1 U10780 ( .A1(n9686), .A2(n8582), .ZN(n8425) );
  NAND2_X1 U10781 ( .A1(n6673), .A2(n9178), .ZN(n8424) );
  NAND2_X1 U10782 ( .A1(n8425), .A2(n8424), .ZN(n8484) );
  NAND2_X1 U10783 ( .A1(n8464), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8429) );
  NAND2_X1 U10784 ( .A1(n8542), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8428) );
  NAND2_X1 U10785 ( .A1(n8513), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8427) );
  NAND2_X1 U10786 ( .A1(n8514), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8426) );
  NAND2_X1 U10787 ( .A1(n10717), .A2(SI_0_), .ZN(n8430) );
  XNOR2_X1 U10788 ( .A(n8430), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n14435) );
  MUX2_X1 U10789 ( .A(n15565), .B(n14435), .S(n10760), .Z(n15691) );
  NAND2_X1 U10790 ( .A1(n13947), .A2(n8434), .ZN(n8431) );
  INV_X1 U10791 ( .A(n10957), .ZN(n11557) );
  NAND2_X1 U10792 ( .A1(n7046), .A2(n14272), .ZN(n9685) );
  NAND3_X1 U10793 ( .A1(n8431), .A2(n11557), .A3(n9685), .ZN(n8432) );
  OAI21_X1 U10794 ( .B1(n8485), .B2(n8484), .A(n8432), .ZN(n8491) );
  NOR2_X1 U10795 ( .A1(n13947), .A2(n6673), .ZN(n8433) );
  INV_X1 U10796 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10718) );
  MUX2_X1 U10797 ( .A(n10718), .B(n8440), .S(n8405), .Z(n8471) );
  INV_X1 U10798 ( .A(n8471), .ZN(n8441) );
  NAND2_X1 U10799 ( .A1(n8442), .A2(SI_3_), .ZN(n8502) );
  OAI21_X1 U10800 ( .B1(n8442), .B2(SI_3_), .A(n8502), .ZN(n8445) );
  AND2_X1 U10801 ( .A1(n8444), .A2(n8445), .ZN(n8443) );
  INV_X1 U10802 ( .A(n8445), .ZN(n8446) );
  AND2_X1 U10803 ( .A1(n8503), .A2(n8448), .ZN(n10715) );
  NAND2_X1 U10804 ( .A1(n10715), .A2(n6680), .ZN(n8454) );
  NAND2_X1 U10805 ( .A1(n8511), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8449) );
  XNOR2_X1 U10806 ( .A(n8449), .B(P2_IR_REG_3__SCAN_IN), .ZN(n13950) );
  INV_X1 U10807 ( .A(n13950), .ZN(n8450) );
  NAND2_X1 U10808 ( .A1(n9124), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8451) );
  AND2_X1 U10809 ( .A1(n8452), .A2(n8451), .ZN(n8453) );
  NAND2_X1 U10810 ( .A1(n13783), .A2(n6673), .ZN(n8461) );
  INV_X1 U10811 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8455) );
  NAND2_X1 U10812 ( .A1(n8542), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8458) );
  NAND2_X1 U10813 ( .A1(n8513), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8457) );
  NAND2_X1 U10814 ( .A1(n8514), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8456) );
  NAND2_X1 U10815 ( .A1(n13945), .A2(n8582), .ZN(n8460) );
  NAND2_X1 U10816 ( .A1(n8513), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8468) );
  NAND2_X1 U10817 ( .A1(n8514), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8467) );
  NAND2_X1 U10818 ( .A1(n8464), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8465) );
  NAND2_X1 U10819 ( .A1(n13946), .A2(n6673), .ZN(n8480) );
  NAND2_X1 U10820 ( .A1(n8470), .A2(n8471), .ZN(n8472) );
  INV_X1 U10821 ( .A(n8474), .ZN(n8475) );
  NAND2_X1 U10822 ( .A1(n8475), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8476) );
  XNOR2_X1 U10823 ( .A(n8476), .B(P2_IR_REG_2__SCAN_IN), .ZN(n10812) );
  INV_X1 U10824 ( .A(n10812), .ZN(n8477) );
  NAND2_X1 U10825 ( .A1(n11109), .A2(n8582), .ZN(n8479) );
  NAND2_X1 U10826 ( .A1(n8480), .A2(n8479), .ZN(n8493) );
  INV_X1 U10827 ( .A(n8493), .ZN(n8483) );
  NAND2_X1 U10828 ( .A1(n6673), .A2(n11109), .ZN(n8482) );
  NAND2_X1 U10829 ( .A1(n13946), .A2(n8582), .ZN(n8481) );
  NAND2_X1 U10830 ( .A1(n8483), .A2(n8492), .ZN(n8487) );
  NAND2_X1 U10831 ( .A1(n8485), .A2(n8484), .ZN(n8486) );
  OAI211_X1 U10832 ( .C1(n8491), .C2(n8490), .A(n8489), .B(n8488), .ZN(n8501)
         );
  INV_X1 U10833 ( .A(n8492), .ZN(n8494) );
  NAND2_X1 U10834 ( .A1(n8494), .A2(n8493), .ZN(n8499) );
  NAND2_X1 U10835 ( .A1(n8499), .A2(n8498), .ZN(n8497) );
  NAND2_X1 U10836 ( .A1(n8497), .A2(n8496), .ZN(n8500) );
  NAND3_X1 U10837 ( .A1(n8501), .A2(n8500), .A3(n6757), .ZN(n8524) );
  INV_X1 U10838 ( .A(n8508), .ZN(n8505) );
  MUX2_X1 U10839 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n8405), .Z(n8504) );
  NAND2_X1 U10840 ( .A1(n8504), .A2(SI_4_), .ZN(n8527) );
  OAI21_X1 U10841 ( .B1(SI_4_), .B2(n8504), .A(n8527), .ZN(n8506) );
  NAND2_X1 U10842 ( .A1(n8505), .A2(n8506), .ZN(n8509) );
  INV_X1 U10843 ( .A(n8506), .ZN(n8507) );
  NAND2_X1 U10844 ( .A1(n8509), .A2(n8528), .ZN(n9996) );
  OR2_X1 U10845 ( .A1(n9996), .A2(n8510), .ZN(n8512) );
  OR2_X1 U10846 ( .A1(n8511), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n8566) );
  NAND2_X1 U10847 ( .A1(n8566), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8537) );
  XNOR2_X1 U10848 ( .A(n8537), .B(P2_IR_REG_4__SCAN_IN), .ZN(n13964) );
  NAND2_X1 U10849 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8544) );
  OAI21_X1 U10850 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n8544), .ZN(n15661) );
  OR2_X1 U10851 ( .A1(n9130), .A2(n15661), .ZN(n8518) );
  INV_X1 U10852 ( .A(n8513), .ZN(n9132) );
  NAND2_X1 U10853 ( .A1(n9109), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8517) );
  NAND2_X1 U10854 ( .A1(n8542), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8516) );
  NAND2_X1 U10855 ( .A1(n8514), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8515) );
  AND2_X1 U10856 ( .A1(n13944), .A2(n8582), .ZN(n8519) );
  NAND2_X1 U10857 ( .A1(n11125), .A2(n9114), .ZN(n8521) );
  NAND2_X1 U10858 ( .A1(n13944), .A2(n6673), .ZN(n8520) );
  NAND2_X1 U10859 ( .A1(n8521), .A2(n8520), .ZN(n8522) );
  OAI21_X1 U10860 ( .B1(n8524), .B2(n8523), .A(n8522), .ZN(n8526) );
  NAND2_X1 U10861 ( .A1(n8524), .A2(n8523), .ZN(n8525) );
  NAND2_X1 U10862 ( .A1(n8526), .A2(n8525), .ZN(n8553) );
  MUX2_X1 U10863 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n8405), .Z(n8529) );
  NAND2_X1 U10864 ( .A1(n8529), .A2(SI_5_), .ZN(n8558) );
  INV_X1 U10865 ( .A(n8529), .ZN(n8530) );
  NAND2_X1 U10866 ( .A1(n8530), .A2(n10701), .ZN(n8531) );
  OR2_X1 U10867 ( .A1(n8533), .A2(n8532), .ZN(n8534) );
  NAND2_X1 U10868 ( .A1(n10743), .A2(n6681), .ZN(n8541) );
  INV_X1 U10869 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8536) );
  NAND2_X1 U10870 ( .A1(n8537), .A2(n8536), .ZN(n8538) );
  NAND2_X1 U10871 ( .A1(n8538), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8539) );
  XNOR2_X1 U10872 ( .A(n8539), .B(P2_IR_REG_5__SCAN_IN), .ZN(n13980) );
  AOI22_X1 U10873 ( .A1(n9124), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8884), .B2(
        n13980), .ZN(n8540) );
  NAND2_X1 U10874 ( .A1(n11590), .A2(n9114), .ZN(n8551) );
  NAND2_X1 U10875 ( .A1(n8514), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8549) );
  NAND2_X1 U10876 ( .A1(n8596), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8548) );
  NOR2_X1 U10877 ( .A1(n8544), .A2(n8543), .ZN(n8574) );
  INV_X1 U10878 ( .A(n8574), .ZN(n8576) );
  NAND2_X1 U10879 ( .A1(n8544), .A2(n8543), .ZN(n8545) );
  NAND2_X1 U10880 ( .A1(n8576), .A2(n8545), .ZN(n11591) );
  NAND2_X1 U10881 ( .A1(n9109), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8546) );
  NAND4_X1 U10882 ( .A1(n8549), .A2(n8548), .A3(n8547), .A4(n8546), .ZN(n13943) );
  NAND2_X1 U10883 ( .A1(n6673), .A2(n13943), .ZN(n8550) );
  NAND2_X1 U10884 ( .A1(n8551), .A2(n8550), .ZN(n8552) );
  NAND2_X1 U10885 ( .A1(n8553), .A2(n8552), .ZN(n8556) );
  AOI22_X1 U10886 ( .A1(n11590), .A2(n6673), .B1(n9114), .B2(n13943), .ZN(
        n8554) );
  MUX2_X1 U10887 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n10717), .Z(n8560) );
  NAND2_X1 U10888 ( .A1(n8560), .A2(SI_6_), .ZN(n8586) );
  INV_X1 U10889 ( .A(n8560), .ZN(n8561) );
  NAND2_X1 U10890 ( .A1(n8561), .A2(n10710), .ZN(n8562) );
  NAND2_X1 U10891 ( .A1(n8564), .A2(n8563), .ZN(n8587) );
  OR2_X1 U10892 ( .A1(n8564), .A2(n8563), .ZN(n8565) );
  NAND2_X1 U10893 ( .A1(n8587), .A2(n8565), .ZN(n10748) );
  OR2_X1 U10894 ( .A1(n10748), .A2(n8510), .ZN(n8573) );
  INV_X1 U10895 ( .A(n8566), .ZN(n8568) );
  NOR2_X1 U10896 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n8567) );
  NAND2_X1 U10897 ( .A1(n8568), .A2(n8567), .ZN(n8570) );
  NAND2_X1 U10898 ( .A1(n8570), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8569) );
  MUX2_X1 U10899 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8569), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n8571) );
  AOI22_X1 U10900 ( .A1(n9124), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8884), .B2(
        n13995), .ZN(n8572) );
  NAND2_X1 U10901 ( .A1(n8573), .A2(n8572), .ZN(n11395) );
  NAND2_X1 U10902 ( .A1(n11395), .A2(n6673), .ZN(n8583) );
  NAND2_X1 U10903 ( .A1(n8514), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8581) );
  NAND2_X1 U10904 ( .A1(n8596), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8580) );
  NAND2_X1 U10905 ( .A1(n8574), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8597) );
  INV_X1 U10906 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8575) );
  NAND2_X1 U10907 ( .A1(n8576), .A2(n8575), .ZN(n8577) );
  NAND2_X1 U10908 ( .A1(n8597), .A2(n8577), .ZN(n11579) );
  OR2_X1 U10909 ( .A1(n9130), .A2(n11579), .ZN(n8579) );
  NAND2_X1 U10910 ( .A1(n9109), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8578) );
  NAND4_X1 U10911 ( .A1(n8581), .A2(n8580), .A3(n8579), .A4(n8578), .ZN(n13942) );
  AOI22_X1 U10912 ( .A1(n11395), .A2(n9114), .B1(n6673), .B2(n13942), .ZN(
        n8584) );
  INV_X1 U10913 ( .A(n8584), .ZN(n8585) );
  NAND2_X1 U10914 ( .A1(n8587), .A2(n8586), .ZN(n8591) );
  MUX2_X1 U10915 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n10717), .Z(n8588) );
  NAND2_X1 U10916 ( .A1(n8588), .A2(SI_7_), .ZN(n8608) );
  OAI21_X1 U10917 ( .B1(SI_7_), .B2(n8588), .A(n8608), .ZN(n8589) );
  INV_X1 U10918 ( .A(n8589), .ZN(n8590) );
  OR2_X1 U10919 ( .A1(n8591), .A2(n8590), .ZN(n8592) );
  NAND2_X1 U10920 ( .A1(n8609), .A2(n8592), .ZN(n10752) );
  OR2_X1 U10921 ( .A1(n10752), .A2(n8510), .ZN(n8595) );
  NAND2_X1 U10922 ( .A1(n8615), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8593) );
  XNOR2_X1 U10923 ( .A(n8593), .B(P2_IR_REG_7__SCAN_IN), .ZN(n14011) );
  AOI22_X1 U10924 ( .A1(n9124), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8884), .B2(
        n14011), .ZN(n8594) );
  NAND2_X1 U10925 ( .A1(n8595), .A2(n8594), .ZN(n11534) );
  NAND2_X1 U10926 ( .A1(n11534), .A2(n9114), .ZN(n8604) );
  NAND2_X1 U10927 ( .A1(n8596), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8602) );
  NAND2_X1 U10928 ( .A1(n8514), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8601) );
  NAND2_X1 U10929 ( .A1(n8597), .A2(n11489), .ZN(n8598) );
  NAND2_X1 U10930 ( .A1(n8621), .A2(n8598), .ZN(n11602) );
  OR2_X1 U10931 ( .A1(n9130), .A2(n11602), .ZN(n8600) );
  NAND2_X1 U10932 ( .A1(n9109), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8599) );
  NAND4_X1 U10933 ( .A1(n8602), .A2(n8601), .A3(n8600), .A4(n8599), .ZN(n13941) );
  NAND2_X1 U10934 ( .A1(n6673), .A2(n13941), .ZN(n8603) );
  AOI22_X1 U10935 ( .A1(n11534), .A2(n6673), .B1(n9114), .B2(n13941), .ZN(
        n8606) );
  INV_X1 U10936 ( .A(n8606), .ZN(n8607) );
  MUX2_X1 U10937 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10717), .Z(n8610) );
  NAND2_X1 U10938 ( .A1(n8610), .A2(SI_8_), .ZN(n8632) );
  OAI21_X1 U10939 ( .B1(SI_8_), .B2(n8610), .A(n8632), .ZN(n8611) );
  INV_X1 U10940 ( .A(n8611), .ZN(n8612) );
  OR2_X1 U10941 ( .A1(n8613), .A2(n8612), .ZN(n8614) );
  INV_X1 U10942 ( .A(n8615), .ZN(n8617) );
  INV_X1 U10943 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n8616) );
  NAND2_X1 U10944 ( .A1(n8617), .A2(n8616), .ZN(n8639) );
  NAND2_X1 U10945 ( .A1(n8639), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8618) );
  XNOR2_X1 U10946 ( .A(n8618), .B(P2_IR_REG_8__SCAN_IN), .ZN(n14026) );
  AOI22_X1 U10947 ( .A1(n9124), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8884), .B2(
        n14026), .ZN(n8619) );
  NAND2_X1 U10948 ( .A1(n11754), .A2(n6673), .ZN(n8628) );
  NAND2_X1 U10949 ( .A1(n8514), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8626) );
  NAND2_X1 U10950 ( .A1(n8596), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8625) );
  INV_X2 U10951 ( .A(n9132), .ZN(n9109) );
  NAND2_X1 U10952 ( .A1(n9109), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8624) );
  NAND2_X1 U10953 ( .A1(n8621), .A2(n8620), .ZN(n8622) );
  NAND2_X1 U10954 ( .A1(n8645), .A2(n8622), .ZN(n11866) );
  OR2_X1 U10955 ( .A1(n9130), .A2(n11866), .ZN(n8623) );
  NAND4_X1 U10956 ( .A1(n8626), .A2(n8625), .A3(n8624), .A4(n8623), .ZN(n13940) );
  NAND2_X1 U10957 ( .A1(n13940), .A2(n9114), .ZN(n8627) );
  NAND2_X1 U10958 ( .A1(n11754), .A2(n9114), .ZN(n8630) );
  NAND2_X1 U10959 ( .A1(n6673), .A2(n13940), .ZN(n8629) );
  NAND2_X1 U10960 ( .A1(n8630), .A2(n8629), .ZN(n8631) );
  MUX2_X1 U10961 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10717), .Z(n8634) );
  NAND2_X1 U10962 ( .A1(n8634), .A2(SI_9_), .ZN(n8659) );
  OAI21_X1 U10963 ( .B1(n8634), .B2(SI_9_), .A(n8659), .ZN(n8635) );
  INV_X1 U10964 ( .A(n8635), .ZN(n8636) );
  OR2_X1 U10965 ( .A1(n8637), .A2(n8636), .ZN(n8638) );
  NAND2_X1 U10966 ( .A1(n8660), .A2(n8638), .ZN(n10853) );
  OR2_X1 U10967 ( .A1(n10853), .A2(n8510), .ZN(n8642) );
  OAI21_X1 U10968 ( .B1(n8639), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8640) );
  XNOR2_X1 U10969 ( .A(n8640), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10871) );
  AOI22_X1 U10970 ( .A1(n9124), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8884), .B2(
        n10871), .ZN(n8641) );
  NAND2_X1 U10971 ( .A1(n11879), .A2(n9114), .ZN(n8652) );
  NAND2_X1 U10972 ( .A1(n8514), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8650) );
  NAND2_X1 U10973 ( .A1(n8596), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8649) );
  NAND2_X1 U10974 ( .A1(n9109), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8648) );
  INV_X1 U10975 ( .A(n8669), .ZN(n8671) );
  NAND2_X1 U10976 ( .A1(n8645), .A2(n8644), .ZN(n8646) );
  NAND2_X1 U10977 ( .A1(n8671), .A2(n8646), .ZN(n11877) );
  OR2_X1 U10978 ( .A1(n9130), .A2(n11877), .ZN(n8647) );
  NAND4_X1 U10979 ( .A1(n8650), .A2(n8649), .A3(n8648), .A4(n8647), .ZN(n13939) );
  NAND2_X1 U10980 ( .A1(n6673), .A2(n13939), .ZN(n8651) );
  NAND2_X1 U10981 ( .A1(n8652), .A2(n8651), .ZN(n8656) );
  NAND2_X1 U10982 ( .A1(n8657), .A2(n8656), .ZN(n8655) );
  AOI22_X1 U10983 ( .A1(n11879), .A2(n6673), .B1(n9114), .B2(n13939), .ZN(
        n8653) );
  NAND2_X1 U10984 ( .A1(n8655), .A2(n8654), .ZN(n8658) );
  NAND2_X1 U10985 ( .A1(n8658), .A2(n6753), .ZN(n8683) );
  MUX2_X1 U10986 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10717), .Z(n8661) );
  INV_X1 U10987 ( .A(n8661), .ZN(n8662) );
  NAND2_X1 U10988 ( .A1(n8662), .A2(n10720), .ZN(n8663) );
  NAND2_X1 U10989 ( .A1(n8837), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8666) );
  MUX2_X1 U10990 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8666), .S(
        P2_IR_REG_10__SCAN_IN), .Z(n8667) );
  NOR2_X1 U10991 ( .A1(n8837), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n8694) );
  INV_X1 U10992 ( .A(n8694), .ZN(n8691) );
  NAND2_X1 U10993 ( .A1(n8667), .A2(n8691), .ZN(n10885) );
  INV_X1 U10994 ( .A(n10885), .ZN(n12350) );
  AOI22_X1 U10995 ( .A1(n9124), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8884), 
        .B2(n12350), .ZN(n8668) );
  NAND2_X1 U10996 ( .A1(n11991), .A2(n6673), .ZN(n8678) );
  NAND2_X1 U10997 ( .A1(n8596), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8676) );
  NAND2_X1 U10998 ( .A1(n8514), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8675) );
  NAND2_X1 U10999 ( .A1(n9109), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8674) );
  NAND2_X1 U11000 ( .A1(n8669), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8699) );
  INV_X1 U11001 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8670) );
  NAND2_X1 U11002 ( .A1(n8671), .A2(n8670), .ZN(n8672) );
  NAND2_X1 U11003 ( .A1(n8699), .A2(n8672), .ZN(n11904) );
  OR2_X1 U11004 ( .A1(n9130), .A2(n11904), .ZN(n8673) );
  NAND4_X1 U11005 ( .A1(n8676), .A2(n8675), .A3(n8674), .A4(n8673), .ZN(n13938) );
  NAND2_X1 U11006 ( .A1(n13938), .A2(n9114), .ZN(n8677) );
  NAND2_X1 U11007 ( .A1(n8678), .A2(n8677), .ZN(n8684) );
  NAND2_X1 U11008 ( .A1(n8683), .A2(n8684), .ZN(n8682) );
  NAND2_X1 U11009 ( .A1(n11991), .A2(n9114), .ZN(n8680) );
  NAND2_X1 U11010 ( .A1(n6673), .A2(n13938), .ZN(n8679) );
  NAND2_X1 U11011 ( .A1(n8680), .A2(n8679), .ZN(n8681) );
  NAND2_X1 U11012 ( .A1(n8682), .A2(n8681), .ZN(n8688) );
  INV_X1 U11013 ( .A(n8683), .ZN(n8686) );
  INV_X1 U11014 ( .A(n8684), .ZN(n8685) );
  NAND2_X1 U11015 ( .A1(n8686), .A2(n8685), .ZN(n8687) );
  NAND2_X1 U11016 ( .A1(n8688), .A2(n8687), .ZN(n8709) );
  MUX2_X1 U11017 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n10717), .Z(n8710) );
  XNOR2_X1 U11018 ( .A(n8713), .B(n8712), .ZN(n10978) );
  NAND2_X1 U11019 ( .A1(n10978), .A2(n6681), .ZN(n8697) );
  NAND2_X1 U11020 ( .A1(n8691), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8692) );
  MUX2_X1 U11021 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8692), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n8695) );
  INV_X1 U11022 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n8693) );
  AND2_X1 U11023 ( .A1(n8694), .A2(n8693), .ZN(n8739) );
  INV_X1 U11024 ( .A(n8739), .ZN(n8714) );
  AOI22_X1 U11025 ( .A1(n9124), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8884), 
        .B2(n14040), .ZN(n8696) );
  NAND2_X1 U11026 ( .A1(n12105), .A2(n9114), .ZN(n8706) );
  NAND2_X1 U11027 ( .A1(n8514), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8704) );
  NAND2_X1 U11028 ( .A1(n8596), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8703) );
  INV_X1 U11029 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8698) );
  NAND2_X1 U11030 ( .A1(n8699), .A2(n8698), .ZN(n8700) );
  NAND2_X1 U11031 ( .A1(n8719), .A2(n8700), .ZN(n12103) );
  OR2_X1 U11032 ( .A1(n9130), .A2(n12103), .ZN(n8702) );
  NAND2_X1 U11033 ( .A1(n9109), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8701) );
  NAND4_X1 U11034 ( .A1(n8704), .A2(n8703), .A3(n8702), .A4(n8701), .ZN(n13937) );
  NAND2_X1 U11035 ( .A1(n6673), .A2(n13937), .ZN(n8705) );
  NAND2_X1 U11036 ( .A1(n8706), .A2(n8705), .ZN(n8708) );
  AOI22_X1 U11037 ( .A1(n12105), .A2(n6673), .B1(n9114), .B2(n13937), .ZN(
        n8707) );
  INV_X1 U11038 ( .A(n8710), .ZN(n8711) );
  MUX2_X1 U11039 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n10717), .Z(n8733) );
  XNOR2_X1 U11040 ( .A(n8732), .B(n8731), .ZN(n11104) );
  NAND2_X1 U11041 ( .A1(n11104), .A2(n6681), .ZN(n8717) );
  NAND2_X1 U11042 ( .A1(n8714), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8715) );
  XNOR2_X1 U11043 ( .A(n8715), .B(P2_IR_REG_12__SCAN_IN), .ZN(n15586) );
  AOI22_X1 U11044 ( .A1(n9124), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8884), 
        .B2(n15586), .ZN(n8716) );
  NAND2_X1 U11045 ( .A1(n12191), .A2(n6673), .ZN(n8726) );
  NAND2_X1 U11046 ( .A1(n8596), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8724) );
  INV_X1 U11047 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8718) );
  INV_X1 U11048 ( .A(n8743), .ZN(n8744) );
  NAND2_X1 U11049 ( .A1(n8719), .A2(n8718), .ZN(n8720) );
  NAND2_X1 U11050 ( .A1(n8744), .A2(n8720), .ZN(n12189) );
  OR2_X1 U11051 ( .A1(n9130), .A2(n12189), .ZN(n8723) );
  NAND2_X1 U11052 ( .A1(n9109), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8722) );
  NAND2_X1 U11053 ( .A1(n8514), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8721) );
  NAND4_X1 U11054 ( .A1(n8724), .A2(n8723), .A3(n8722), .A4(n8721), .ZN(n13936) );
  NAND2_X1 U11055 ( .A1(n13936), .A2(n9114), .ZN(n8725) );
  NAND2_X1 U11056 ( .A1(n8726), .A2(n8725), .ZN(n8729) );
  NAND2_X1 U11057 ( .A1(n12191), .A2(n9114), .ZN(n8728) );
  NAND2_X1 U11058 ( .A1(n13936), .A2(n6673), .ZN(n8727) );
  INV_X1 U11059 ( .A(n8729), .ZN(n8730) );
  INV_X1 U11060 ( .A(n8733), .ZN(n8734) );
  NAND2_X1 U11061 ( .A1(n8734), .A2(n10742), .ZN(n8735) );
  MUX2_X1 U11062 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n10717), .Z(n8761) );
  INV_X1 U11063 ( .A(SI_13_), .ZN(n8737) );
  XNOR2_X1 U11064 ( .A(n8761), .B(n8737), .ZN(n8738) );
  XNOR2_X1 U11065 ( .A(n8764), .B(n8738), .ZN(n11256) );
  NAND2_X1 U11066 ( .A1(n11256), .A2(n6680), .ZN(n8742) );
  NAND2_X1 U11067 ( .A1(n8739), .A2(n7059), .ZN(n8766) );
  NAND2_X1 U11068 ( .A1(n8766), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8740) );
  XNOR2_X1 U11069 ( .A(n8740), .B(P2_IR_REG_13__SCAN_IN), .ZN(n15594) );
  AOI22_X1 U11070 ( .A1(n9124), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8884), 
        .B2(n15594), .ZN(n8741) );
  NAND2_X1 U11071 ( .A1(n12394), .A2(n9114), .ZN(n8751) );
  NAND2_X1 U11072 ( .A1(n8514), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8749) );
  NAND2_X1 U11073 ( .A1(n8596), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8748) );
  NAND2_X1 U11074 ( .A1(n8743), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8771) );
  INV_X1 U11075 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n12404) );
  NAND2_X1 U11076 ( .A1(n8744), .A2(n12404), .ZN(n8745) );
  NAND2_X1 U11077 ( .A1(n8771), .A2(n8745), .ZN(n12199) );
  OR2_X1 U11078 ( .A1(n9130), .A2(n12199), .ZN(n8747) );
  NAND2_X1 U11079 ( .A1(n9109), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8746) );
  NAND4_X1 U11080 ( .A1(n8749), .A2(n8748), .A3(n8747), .A4(n8746), .ZN(n13935) );
  NAND2_X1 U11081 ( .A1(n13935), .A2(n6673), .ZN(n8750) );
  NAND2_X1 U11082 ( .A1(n8751), .A2(n8750), .ZN(n8756) );
  NAND2_X1 U11083 ( .A1(n8755), .A2(n8756), .ZN(n8754) );
  AOI22_X1 U11084 ( .A1(n12394), .A2(n6673), .B1(n9114), .B2(n13935), .ZN(
        n8752) );
  NAND2_X1 U11085 ( .A1(n8754), .A2(n8753), .ZN(n8760) );
  INV_X1 U11086 ( .A(n8755), .ZN(n8758) );
  INV_X1 U11087 ( .A(n8756), .ZN(n8757) );
  NAND2_X1 U11088 ( .A1(n8758), .A2(n8757), .ZN(n8759) );
  NOR2_X1 U11089 ( .A1(n8761), .A2(SI_13_), .ZN(n8763) );
  NAND2_X1 U11090 ( .A1(n8761), .A2(SI_13_), .ZN(n8762) );
  MUX2_X1 U11091 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n10717), .Z(n8781) );
  XNOR2_X1 U11092 ( .A(n8782), .B(n8781), .ZN(n11608) );
  NAND2_X1 U11093 ( .A1(n11608), .A2(n6680), .ZN(n8769) );
  NAND2_X1 U11094 ( .A1(n8786), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8767) );
  XNOR2_X1 U11095 ( .A(n8767), .B(P2_IR_REG_14__SCAN_IN), .ZN(n15605) );
  AOI22_X1 U11096 ( .A1(n9124), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8884), 
        .B2(n15605), .ZN(n8768) );
  NAND2_X1 U11097 ( .A1(n15280), .A2(n6673), .ZN(n8778) );
  NAND2_X1 U11098 ( .A1(n8514), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8776) );
  NAND2_X1 U11099 ( .A1(n8596), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8775) );
  NAND2_X1 U11100 ( .A1(n9109), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8774) );
  INV_X1 U11101 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8770) );
  NAND2_X1 U11102 ( .A1(n8771), .A2(n8770), .ZN(n8772) );
  NAND2_X1 U11103 ( .A1(n8792), .A2(n8772), .ZN(n15258) );
  OR2_X1 U11104 ( .A1(n9130), .A2(n15258), .ZN(n8773) );
  NAND4_X1 U11105 ( .A1(n8776), .A2(n8775), .A3(n8774), .A4(n8773), .ZN(n13934) );
  NAND2_X1 U11106 ( .A1(n13934), .A2(n9114), .ZN(n8777) );
  NAND2_X1 U11107 ( .A1(n8778), .A2(n8777), .ZN(n8780) );
  AOI22_X1 U11108 ( .A1(n15280), .A2(n9114), .B1(n6673), .B2(n13934), .ZN(
        n8779) );
  MUX2_X1 U11109 ( .A(n11804), .B(n11820), .S(n10717), .Z(n8783) );
  INV_X1 U11110 ( .A(n8783), .ZN(n8784) );
  NAND2_X1 U11111 ( .A1(n8784), .A2(SI_15_), .ZN(n8785) );
  XNOR2_X1 U11112 ( .A(n8806), .B(n8805), .ZN(n11803) );
  NAND2_X1 U11113 ( .A1(n11803), .A2(n6680), .ZN(n8791) );
  OAI21_X1 U11114 ( .B1(n8786), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8788) );
  INV_X1 U11115 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8787) );
  NAND2_X1 U11116 ( .A1(n8788), .A2(n8787), .ZN(n8812) );
  OR2_X1 U11117 ( .A1(n8788), .A2(n8787), .ZN(n8789) );
  AND2_X1 U11118 ( .A1(n8812), .A2(n8789), .ZN(n15615) );
  AOI22_X1 U11119 ( .A1(n9124), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n15615), 
        .B2(n8884), .ZN(n8790) );
  NAND2_X1 U11120 ( .A1(n12570), .A2(n9114), .ZN(n8799) );
  INV_X1 U11121 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n12566) );
  INV_X1 U11122 ( .A(n8816), .ZN(n8818) );
  NAND2_X1 U11123 ( .A1(n8792), .A2(n12566), .ZN(n8793) );
  NAND2_X1 U11124 ( .A1(n8818), .A2(n8793), .ZN(n12565) );
  OR2_X1 U11125 ( .A1(n12565), .A2(n9130), .ZN(n8797) );
  NAND2_X1 U11126 ( .A1(n8514), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8796) );
  NAND2_X1 U11127 ( .A1(n8596), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U11128 ( .A1(n9109), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8794) );
  NAND4_X1 U11129 ( .A1(n8797), .A2(n8796), .A3(n8795), .A4(n8794), .ZN(n13933) );
  NAND2_X1 U11130 ( .A1(n13933), .A2(n6673), .ZN(n8798) );
  NAND2_X1 U11131 ( .A1(n8799), .A2(n8798), .ZN(n8803) );
  INV_X1 U11132 ( .A(n13933), .ZN(n9713) );
  NAND2_X1 U11133 ( .A1(n12570), .A2(n6673), .ZN(n8800) );
  INV_X1 U11134 ( .A(n8803), .ZN(n8804) );
  NAND2_X1 U11135 ( .A1(n8808), .A2(n8807), .ZN(n8830) );
  MUX2_X1 U11136 ( .A(n11973), .B(n11987), .S(n10717), .Z(n8809) );
  INV_X1 U11137 ( .A(n8809), .ZN(n8810) );
  NAND2_X1 U11138 ( .A1(n8810), .A2(SI_16_), .ZN(n8811) );
  XNOR2_X1 U11139 ( .A(n8830), .B(n8829), .ZN(n11972) );
  NAND2_X1 U11140 ( .A1(n11972), .A2(n6680), .ZN(n8815) );
  NAND2_X1 U11141 ( .A1(n8812), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8813) );
  XNOR2_X1 U11142 ( .A(n8813), .B(P2_IR_REG_16__SCAN_IN), .ZN(n15627) );
  AOI22_X1 U11143 ( .A1(n15627), .A2(n8884), .B1(n9124), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n8814) );
  NAND2_X1 U11144 ( .A1(n14364), .A2(n6673), .ZN(n8823) );
  INV_X1 U11145 ( .A(n8843), .ZN(n8845) );
  INV_X1 U11146 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8817) );
  NAND2_X1 U11147 ( .A1(n8818), .A2(n8817), .ZN(n8819) );
  NAND2_X1 U11148 ( .A1(n8845), .A2(n8819), .ZN(n14271) );
  AOI22_X1 U11149 ( .A1(n8514), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n8596), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n8821) );
  NAND2_X1 U11150 ( .A1(n9109), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8820) );
  OAI211_X1 U11151 ( .C1(n14271), .C2(n9130), .A(n8821), .B(n8820), .ZN(n13932) );
  NAND2_X1 U11152 ( .A1(n13932), .A2(n9114), .ZN(n8822) );
  NAND2_X1 U11153 ( .A1(n8823), .A2(n8822), .ZN(n8826) );
  AOI22_X1 U11154 ( .A1(n14364), .A2(n9114), .B1(n6673), .B2(n13932), .ZN(
        n8824) );
  INV_X1 U11155 ( .A(n8825), .ZN(n8828) );
  NAND2_X1 U11156 ( .A1(n8830), .A2(n8829), .ZN(n8832) );
  MUX2_X1 U11157 ( .A(n12037), .B(n12066), .S(n10717), .Z(n8833) );
  INV_X1 U11158 ( .A(SI_17_), .ZN(n10977) );
  NAND2_X1 U11159 ( .A1(n8833), .A2(n10977), .ZN(n8859) );
  INV_X1 U11160 ( .A(n8833), .ZN(n8834) );
  NAND2_X1 U11161 ( .A1(n8834), .A2(SI_17_), .ZN(n8835) );
  XNOR2_X1 U11162 ( .A(n8858), .B(n8857), .ZN(n12036) );
  NAND2_X1 U11163 ( .A1(n12036), .A2(n6681), .ZN(n8842) );
  OR2_X1 U11164 ( .A1(n8837), .A2(n8836), .ZN(n8839) );
  NAND2_X1 U11165 ( .A1(n8839), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8838) );
  MUX2_X1 U11166 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8838), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n8840) );
  OR2_X1 U11167 ( .A1(n8839), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n8861) );
  AND2_X1 U11168 ( .A1(n8840), .A2(n8861), .ZN(n15640) );
  AOI22_X1 U11169 ( .A1(n9124), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8884), 
        .B2(n15640), .ZN(n8841) );
  NAND2_X1 U11170 ( .A1(n14359), .A2(n9114), .ZN(n8851) );
  INV_X1 U11171 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8849) );
  INV_X1 U11172 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8844) );
  NAND2_X1 U11173 ( .A1(n8845), .A2(n8844), .ZN(n8846) );
  NAND2_X1 U11174 ( .A1(n8865), .A2(n8846), .ZN(n14253) );
  OR2_X1 U11175 ( .A1(n14253), .A2(n9130), .ZN(n8848) );
  AOI22_X1 U11176 ( .A1(n8514), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n8596), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n8847) );
  OAI211_X1 U11177 ( .C1(n9132), .C2(n8849), .A(n8848), .B(n8847), .ZN(n13931)
         );
  NAND2_X1 U11178 ( .A1(n13931), .A2(n6673), .ZN(n8850) );
  NAND2_X1 U11179 ( .A1(n8851), .A2(n8850), .ZN(n8855) );
  NAND2_X1 U11180 ( .A1(n14359), .A2(n6673), .ZN(n8853) );
  NAND2_X1 U11181 ( .A1(n13931), .A2(n9114), .ZN(n8852) );
  NAND2_X1 U11182 ( .A1(n8853), .A2(n8852), .ZN(n8854) );
  INV_X1 U11183 ( .A(n8855), .ZN(n8856) );
  NAND2_X1 U11184 ( .A1(n8858), .A2(n8857), .ZN(n8860) );
  XNOR2_X1 U11185 ( .A(n8900), .B(SI_18_), .ZN(n8879) );
  MUX2_X1 U11186 ( .A(n12296), .B(n12317), .S(n10717), .Z(n8897) );
  XNOR2_X1 U11187 ( .A(n8879), .B(n8897), .ZN(n12295) );
  NAND2_X1 U11188 ( .A1(n12295), .A2(n6681), .ZN(n8864) );
  NAND2_X1 U11189 ( .A1(n8861), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8862) );
  XNOR2_X1 U11190 ( .A(n8862), .B(P2_IR_REG_18__SCAN_IN), .ZN(n12579) );
  AOI22_X1 U11191 ( .A1(n9124), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8884), 
        .B2(n12579), .ZN(n8863) );
  NAND2_X2 U11192 ( .A1(n8864), .A2(n8863), .ZN(n14353) );
  NAND2_X1 U11193 ( .A1(n14353), .A2(n6673), .ZN(n8874) );
  INV_X1 U11194 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n12373) );
  NAND2_X1 U11195 ( .A1(n8865), .A2(n12373), .ZN(n8866) );
  NAND2_X1 U11196 ( .A1(n8888), .A2(n8866), .ZN(n14233) );
  OR2_X1 U11197 ( .A1(n14233), .A2(n9130), .ZN(n8872) );
  INV_X1 U11198 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8869) );
  NAND2_X1 U11199 ( .A1(n8596), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8868) );
  NAND2_X1 U11200 ( .A1(n9109), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8867) );
  OAI211_X1 U11201 ( .C1(n8869), .C2(n9112), .A(n8868), .B(n8867), .ZN(n8870)
         );
  INV_X1 U11202 ( .A(n8870), .ZN(n8871) );
  NAND2_X1 U11203 ( .A1(n8872), .A2(n8871), .ZN(n13930) );
  NAND2_X1 U11204 ( .A1(n13930), .A2(n9114), .ZN(n8873) );
  NAND2_X1 U11205 ( .A1(n8874), .A2(n8873), .ZN(n8876) );
  AOI22_X1 U11206 ( .A1(n14353), .A2(n9114), .B1(n6673), .B2(n13930), .ZN(
        n8875) );
  INV_X1 U11207 ( .A(n8897), .ZN(n8901) );
  NOR2_X1 U11208 ( .A1(n8900), .A2(n11183), .ZN(n8878) );
  AOI21_X1 U11209 ( .B1(n8879), .B2(n8901), .A(n8878), .ZN(n8883) );
  MUX2_X1 U11210 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10717), .Z(n8880) );
  NAND2_X1 U11211 ( .A1(n8880), .A2(SI_19_), .ZN(n8904) );
  INV_X1 U11212 ( .A(n8880), .ZN(n8881) );
  NAND2_X1 U11213 ( .A1(n8881), .A2(n11254), .ZN(n8902) );
  AND2_X1 U11214 ( .A1(n8904), .A2(n8902), .ZN(n8882) );
  NAND2_X1 U11215 ( .A1(n12387), .A2(n6680), .ZN(n8886) );
  AOI22_X1 U11216 ( .A1(n9124), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n14272), 
        .B2(n8884), .ZN(n8885) );
  NAND2_X1 U11217 ( .A1(n14345), .A2(n9114), .ZN(n8895) );
  INV_X1 U11218 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8887) );
  NAND2_X1 U11219 ( .A1(n8888), .A2(n8887), .ZN(n8889) );
  NAND2_X1 U11220 ( .A1(n8910), .A2(n8889), .ZN(n14219) );
  INV_X1 U11221 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14349) );
  NAND2_X1 U11222 ( .A1(n9109), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8891) );
  NAND2_X1 U11223 ( .A1(n8596), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8890) );
  OAI211_X1 U11224 ( .C1(n9112), .C2(n14349), .A(n8891), .B(n8890), .ZN(n8892)
         );
  INV_X1 U11225 ( .A(n8892), .ZN(n8893) );
  OAI21_X1 U11226 ( .B1(n14219), .B2(n9130), .A(n8893), .ZN(n13929) );
  NAND2_X1 U11227 ( .A1(n13929), .A2(n6673), .ZN(n8894) );
  AOI22_X1 U11228 ( .A1(n14345), .A2(n6673), .B1(n9114), .B2(n13929), .ZN(
        n8896) );
  OAI21_X1 U11229 ( .B1(n11183), .B2(n8897), .A(n8904), .ZN(n8898) );
  INV_X1 U11230 ( .A(n8898), .ZN(n8899) );
  NOR2_X1 U11231 ( .A1(n8901), .A2(SI_18_), .ZN(n8905) );
  INV_X1 U11232 ( .A(n8902), .ZN(n8903) );
  AOI21_X1 U11233 ( .B1(n8905), .B2(n8904), .A(n8903), .ZN(n8906) );
  XNOR2_X1 U11234 ( .A(n8959), .B(n11661), .ZN(n8925) );
  MUX2_X1 U11235 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n10717), .Z(n8954) );
  XNOR2_X1 U11236 ( .A(n8925), .B(n8954), .ZN(n12391) );
  NAND2_X1 U11237 ( .A1(n12391), .A2(n6681), .ZN(n8909) );
  NAND2_X1 U11238 ( .A1(n9124), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8908) );
  INV_X1 U11239 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13868) );
  INV_X1 U11240 ( .A(n8933), .ZN(n8935) );
  NAND2_X1 U11241 ( .A1(n8910), .A2(n13868), .ZN(n8911) );
  AND2_X1 U11242 ( .A1(n8935), .A2(n8911), .ZN(n14205) );
  NAND2_X1 U11243 ( .A1(n14205), .A2(n8464), .ZN(n8917) );
  INV_X1 U11244 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8914) );
  NAND2_X1 U11245 ( .A1(n8596), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8913) );
  NAND2_X1 U11246 ( .A1(n9109), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8912) );
  OAI211_X1 U11247 ( .C1(n8914), .C2(n9112), .A(n8913), .B(n8912), .ZN(n8915)
         );
  INV_X1 U11248 ( .A(n8915), .ZN(n8916) );
  NAND2_X1 U11249 ( .A1(n8917), .A2(n8916), .ZN(n13928) );
  AND2_X1 U11250 ( .A1(n13928), .A2(n9114), .ZN(n8918) );
  AOI21_X1 U11251 ( .B1(n14341), .B2(n6673), .A(n8918), .ZN(n8921) );
  INV_X1 U11252 ( .A(n13928), .ZN(n9722) );
  NAND2_X1 U11253 ( .A1(n14341), .A2(n9114), .ZN(n8919) );
  OAI21_X1 U11254 ( .B1(n9722), .B2(n9114), .A(n8919), .ZN(n8920) );
  NAND2_X1 U11255 ( .A1(n8922), .A2(n8921), .ZN(n8923) );
  NAND2_X1 U11256 ( .A1(n8924), .A2(n8923), .ZN(n8949) );
  INV_X1 U11257 ( .A(n8925), .ZN(n8926) );
  NAND2_X1 U11258 ( .A1(n8926), .A2(n8954), .ZN(n8928) );
  OR2_X1 U11259 ( .A1(n8959), .A2(n11661), .ZN(n8927) );
  NAND2_X1 U11260 ( .A1(n8928), .A2(n8927), .ZN(n8930) );
  MUX2_X1 U11261 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n10717), .Z(n8956) );
  XNOR2_X1 U11262 ( .A(n8956), .B(SI_21_), .ZN(n8929) );
  NAND2_X1 U11263 ( .A1(n12463), .A2(n6680), .ZN(n8932) );
  OR2_X1 U11264 ( .A1(n8469), .A2(n12465), .ZN(n8931) );
  NAND2_X1 U11265 ( .A1(n8933), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8962) );
  INV_X1 U11266 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8934) );
  NAND2_X1 U11267 ( .A1(n8935), .A2(n8934), .ZN(n8936) );
  NAND2_X1 U11268 ( .A1(n8962), .A2(n8936), .ZN(n14187) );
  OR2_X1 U11269 ( .A1(n14187), .A2(n9130), .ZN(n8942) );
  INV_X1 U11270 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8939) );
  NAND2_X1 U11271 ( .A1(n9109), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8938) );
  NAND2_X1 U11272 ( .A1(n8596), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8937) );
  OAI211_X1 U11273 ( .C1(n9112), .C2(n8939), .A(n8938), .B(n8937), .ZN(n8940)
         );
  INV_X1 U11274 ( .A(n8940), .ZN(n8941) );
  NAND2_X1 U11275 ( .A1(n8942), .A2(n8941), .ZN(n13927) );
  AND2_X1 U11276 ( .A1(n13927), .A2(n6673), .ZN(n8943) );
  AOI21_X1 U11277 ( .B1(n14337), .B2(n9114), .A(n8943), .ZN(n8950) );
  INV_X1 U11278 ( .A(n8950), .ZN(n8944) );
  NAND2_X1 U11279 ( .A1(n8949), .A2(n8944), .ZN(n8948) );
  NAND2_X1 U11280 ( .A1(n14337), .A2(n6673), .ZN(n8946) );
  NAND2_X1 U11281 ( .A1(n13927), .A2(n9114), .ZN(n8945) );
  NAND2_X1 U11282 ( .A1(n8946), .A2(n8945), .ZN(n8947) );
  NAND2_X1 U11283 ( .A1(n8948), .A2(n8947), .ZN(n8953) );
  INV_X1 U11284 ( .A(n8949), .ZN(n8951) );
  NAND2_X1 U11285 ( .A1(n8951), .A2(n8950), .ZN(n8952) );
  NAND2_X1 U11286 ( .A1(n8953), .A2(n8952), .ZN(n8974) );
  INV_X1 U11287 ( .A(n8954), .ZN(n8955) );
  NOR2_X1 U11288 ( .A1(n8955), .A2(n11661), .ZN(n8957) );
  AOI22_X1 U11289 ( .A1(n8957), .A2(n7765), .B1(n8956), .B2(SI_21_), .ZN(n8958) );
  MUX2_X1 U11290 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n10717), .Z(n8977) );
  XNOR2_X1 U11291 ( .A(n8976), .B(n8977), .ZN(n12557) );
  NAND2_X1 U11292 ( .A1(n12557), .A2(n6681), .ZN(n8961) );
  OR2_X1 U11293 ( .A1(n8469), .A2(n12559), .ZN(n8960) );
  NAND2_X1 U11294 ( .A1(n14394), .A2(n6673), .ZN(n8971) );
  INV_X1 U11295 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13883) );
  NAND2_X1 U11296 ( .A1(n8962), .A2(n13883), .ZN(n8963) );
  AND2_X1 U11297 ( .A1(n8983), .A2(n8963), .ZN(n14173) );
  NAND2_X1 U11298 ( .A1(n14173), .A2(n8464), .ZN(n8969) );
  INV_X1 U11299 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8966) );
  NAND2_X1 U11300 ( .A1(n9109), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8965) );
  NAND2_X1 U11301 ( .A1(n8596), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8964) );
  OAI211_X1 U11302 ( .C1(n9112), .C2(n8966), .A(n8965), .B(n8964), .ZN(n8967)
         );
  INV_X1 U11303 ( .A(n8967), .ZN(n8968) );
  NAND2_X1 U11304 ( .A1(n8969), .A2(n8968), .ZN(n13926) );
  NAND2_X1 U11305 ( .A1(n13926), .A2(n9114), .ZN(n8970) );
  NAND2_X1 U11306 ( .A1(n8971), .A2(n8970), .ZN(n8975) );
  AOI22_X1 U11307 ( .A1(n14394), .A2(n9114), .B1(n6673), .B2(n13926), .ZN(
        n8972) );
  INV_X1 U11308 ( .A(n8972), .ZN(n8973) );
  MUX2_X1 U11309 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10717), .Z(n8999) );
  XNOR2_X1 U11310 ( .A(n8999), .B(SI_23_), .ZN(n8980) );
  XNOR2_X1 U11311 ( .A(n8998), .B(n8980), .ZN(n12629) );
  NAND2_X1 U11312 ( .A1(n12629), .A2(n6680), .ZN(n8982) );
  OR2_X1 U11313 ( .A1(n8469), .A2(n12628), .ZN(n8981) );
  NAND2_X1 U11314 ( .A1(n14159), .A2(n9114), .ZN(n8991) );
  INV_X1 U11315 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13774) );
  AOI21_X1 U11316 ( .B1(n8983), .B2(n13774), .A(n9004), .ZN(n14155) );
  NAND2_X1 U11317 ( .A1(n14155), .A2(n8464), .ZN(n8989) );
  INV_X1 U11318 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8986) );
  NAND2_X1 U11319 ( .A1(n9109), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8985) );
  NAND2_X1 U11320 ( .A1(n8596), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8984) );
  OAI211_X1 U11321 ( .C1(n9112), .C2(n8986), .A(n8985), .B(n8984), .ZN(n8987)
         );
  INV_X1 U11322 ( .A(n8987), .ZN(n8988) );
  NAND2_X1 U11323 ( .A1(n8989), .A2(n8988), .ZN(n13925) );
  NAND2_X1 U11324 ( .A1(n13925), .A2(n6673), .ZN(n8990) );
  NAND2_X1 U11325 ( .A1(n8991), .A2(n8990), .ZN(n8994) );
  INV_X1 U11326 ( .A(n13925), .ZN(n13858) );
  NAND2_X1 U11327 ( .A1(n14159), .A2(n6673), .ZN(n8992) );
  OAI21_X1 U11328 ( .B1(n6673), .B2(n13858), .A(n8992), .ZN(n8993) );
  INV_X1 U11329 ( .A(n8994), .ZN(n8995) );
  INV_X1 U11330 ( .A(n8999), .ZN(n8996) );
  NAND2_X1 U11331 ( .A1(n8996), .A2(n12177), .ZN(n8997) );
  NAND2_X1 U11332 ( .A1(n8999), .A2(SI_23_), .ZN(n9000) );
  MUX2_X1 U11333 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n10717), .Z(n9016) );
  XNOR2_X1 U11334 ( .A(n9020), .B(n9016), .ZN(n14430) );
  NAND2_X1 U11335 ( .A1(n14430), .A2(n6681), .ZN(n9003) );
  NAND2_X1 U11336 ( .A1(n9124), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9002) );
  NAND2_X1 U11337 ( .A1(n14316), .A2(n6673), .ZN(n9010) );
  NAND2_X1 U11338 ( .A1(n8596), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9008) );
  NAND2_X1 U11339 ( .A1(n8514), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n9007) );
  NAND2_X1 U11340 ( .A1(n9109), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9006) );
  NAND2_X1 U11341 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n9004), .ZN(n9028) );
  OAI21_X1 U11342 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n9004), .A(n9028), .ZN(
        n14136) );
  OR2_X1 U11343 ( .A1(n9130), .A2(n14136), .ZN(n9005) );
  NAND4_X1 U11344 ( .A1(n9008), .A2(n9007), .A3(n9006), .A4(n9005), .ZN(n13924) );
  NAND2_X1 U11345 ( .A1(n13924), .A2(n9114), .ZN(n9009) );
  NAND2_X1 U11346 ( .A1(n9010), .A2(n9009), .ZN(n9012) );
  AOI22_X1 U11347 ( .A1(n14316), .A2(n9114), .B1(n6673), .B2(n13924), .ZN(
        n9011) );
  AOI21_X1 U11348 ( .B1(n9013), .B2(n9012), .A(n9011), .ZN(n9015) );
  NOR2_X1 U11349 ( .A1(n9013), .A2(n9012), .ZN(n9014) );
  INV_X1 U11350 ( .A(n9016), .ZN(n9019) );
  MUX2_X1 U11351 ( .A(n15098), .B(n14429), .S(n10717), .Z(n9021) );
  NAND2_X1 U11352 ( .A1(n9021), .A2(n13716), .ZN(n9036) );
  INV_X1 U11353 ( .A(n9021), .ZN(n9022) );
  NAND2_X1 U11354 ( .A1(n9022), .A2(SI_25_), .ZN(n9023) );
  NAND2_X1 U11355 ( .A1(n9036), .A2(n9023), .ZN(n9037) );
  NAND2_X1 U11356 ( .A1(n14426), .A2(n6680), .ZN(n9025) );
  OR2_X1 U11357 ( .A1(n8469), .A2(n14429), .ZN(n9024) );
  NAND2_X1 U11358 ( .A1(n14310), .A2(n9114), .ZN(n9035) );
  NAND2_X1 U11359 ( .A1(n8596), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9033) );
  NAND2_X1 U11360 ( .A1(n8514), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n9032) );
  NAND2_X1 U11361 ( .A1(n9109), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9031) );
  INV_X1 U11362 ( .A(n9028), .ZN(n9026) );
  INV_X1 U11363 ( .A(n9041), .ZN(n9043) );
  INV_X1 U11364 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9027) );
  NAND2_X1 U11365 ( .A1(n9028), .A2(n9027), .ZN(n9029) );
  NAND2_X1 U11366 ( .A1(n9043), .A2(n9029), .ZN(n14121) );
  OR2_X1 U11367 ( .A1(n9130), .A2(n14121), .ZN(n9030) );
  NAND4_X1 U11368 ( .A1(n9033), .A2(n9032), .A3(n9031), .A4(n9030), .ZN(n13923) );
  NAND2_X1 U11369 ( .A1(n6673), .A2(n13923), .ZN(n9034) );
  NAND2_X1 U11370 ( .A1(n9035), .A2(n9034), .ZN(n9054) );
  MUX2_X1 U11371 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n10717), .Z(n9059) );
  XNOR2_X1 U11372 ( .A(n9059), .B(n13710), .ZN(n9038) );
  NAND2_X1 U11373 ( .A1(n14423), .A2(n6681), .ZN(n9040) );
  OR2_X1 U11374 ( .A1(n8469), .A2(n14425), .ZN(n9039) );
  NAND2_X1 U11375 ( .A1(n8514), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n9048) );
  NAND2_X1 U11376 ( .A1(n8596), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9047) );
  NAND2_X1 U11377 ( .A1(n9041), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n9084) );
  INV_X1 U11378 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9042) );
  NAND2_X1 U11379 ( .A1(n9043), .A2(n9042), .ZN(n9044) );
  NAND2_X1 U11380 ( .A1(n9084), .A2(n9044), .ZN(n14106) );
  OR2_X1 U11381 ( .A1(n9130), .A2(n14106), .ZN(n9046) );
  NAND2_X1 U11382 ( .A1(n9109), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9045) );
  NAND4_X1 U11383 ( .A1(n9048), .A2(n9047), .A3(n9046), .A4(n9045), .ZN(n13922) );
  AND2_X1 U11384 ( .A1(n13922), .A2(n9114), .ZN(n9049) );
  AOI21_X1 U11385 ( .B1(n14108), .B2(n6673), .A(n9049), .ZN(n9058) );
  NAND2_X1 U11386 ( .A1(n14108), .A2(n9114), .ZN(n9051) );
  NAND2_X1 U11387 ( .A1(n6673), .A2(n13922), .ZN(n9050) );
  NAND2_X1 U11388 ( .A1(n9051), .A2(n9050), .ZN(n9057) );
  OAI22_X1 U11389 ( .A1(n9055), .A2(n9054), .B1(n9058), .B2(n9057), .ZN(n9052)
         );
  AOI22_X1 U11390 ( .A1(n14310), .A2(n6673), .B1(n9114), .B2(n13923), .ZN(
        n9053) );
  AOI21_X1 U11391 ( .B1(n9055), .B2(n9054), .A(n9053), .ZN(n9056) );
  NAND2_X1 U11392 ( .A1(n9058), .A2(n9057), .ZN(n9095) );
  INV_X1 U11393 ( .A(n9059), .ZN(n9060) );
  NAND2_X1 U11394 ( .A1(n9061), .A2(n13710), .ZN(n9062) );
  MUX2_X1 U11395 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n10717), .Z(n9076) );
  MUX2_X1 U11396 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n10717), .Z(n9096) );
  XNOR2_X1 U11397 ( .A(n9096), .B(SI_28_), .ZN(n9099) );
  NAND2_X1 U11398 ( .A1(n14415), .A2(n6680), .ZN(n9064) );
  OR2_X1 U11399 ( .A1(n8469), .A2(n14418), .ZN(n9063) );
  NAND2_X1 U11400 ( .A1(n8514), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n9072) );
  NAND2_X1 U11401 ( .A1(n8596), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9071) );
  NAND2_X1 U11402 ( .A1(n9109), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9070) );
  INV_X1 U11403 ( .A(n9084), .ZN(n9065) );
  NAND2_X1 U11404 ( .A1(n9066), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n14062) );
  INV_X1 U11405 ( .A(n9066), .ZN(n9086) );
  INV_X1 U11406 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9067) );
  NAND2_X1 U11407 ( .A1(n9086), .A2(n9067), .ZN(n9068) );
  NAND2_X1 U11408 ( .A1(n14062), .A2(n9068), .ZN(n14080) );
  OR2_X1 U11409 ( .A1(n9130), .A2(n14080), .ZN(n9069) );
  NAND4_X1 U11410 ( .A1(n9072), .A2(n9071), .A3(n9070), .A4(n9069), .ZN(n13920) );
  AND2_X1 U11411 ( .A1(n13920), .A2(n6673), .ZN(n9073) );
  AOI21_X1 U11412 ( .B1(n14292), .B2(n9114), .A(n9073), .ZN(n9140) );
  NAND2_X1 U11413 ( .A1(n14292), .A2(n6673), .ZN(n9075) );
  NAND2_X1 U11414 ( .A1(n13920), .A2(n9114), .ZN(n9074) );
  NAND2_X1 U11415 ( .A1(n9075), .A2(n9074), .ZN(n9139) );
  NAND2_X1 U11416 ( .A1(n9140), .A2(n9139), .ZN(n9144) );
  INV_X1 U11417 ( .A(n9076), .ZN(n9077) );
  XNOR2_X1 U11418 ( .A(n9077), .B(SI_27_), .ZN(n9078) );
  OR2_X1 U11419 ( .A1(n8469), .A2(n9080), .ZN(n9081) );
  NAND2_X1 U11420 ( .A1(n8596), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9090) );
  NAND2_X1 U11421 ( .A1(n8514), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n9089) );
  NAND2_X1 U11422 ( .A1(n9109), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9088) );
  INV_X1 U11423 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9083) );
  NAND2_X1 U11424 ( .A1(n9084), .A2(n9083), .ZN(n9085) );
  NAND2_X1 U11425 ( .A1(n9086), .A2(n9085), .ZN(n14092) );
  OR2_X1 U11426 ( .A1(n9130), .A2(n14092), .ZN(n9087) );
  NAND4_X1 U11427 ( .A1(n9090), .A2(n9089), .A3(n9088), .A4(n9087), .ZN(n13921) );
  AND2_X1 U11428 ( .A1(n13921), .A2(n6673), .ZN(n9091) );
  AOI21_X1 U11429 ( .B1(n14091), .B2(n9114), .A(n9091), .ZN(n9138) );
  NAND2_X1 U11430 ( .A1(n14091), .A2(n6673), .ZN(n9093) );
  NAND2_X1 U11431 ( .A1(n13921), .A2(n9114), .ZN(n9092) );
  NAND2_X1 U11432 ( .A1(n9093), .A2(n9092), .ZN(n9137) );
  NAND2_X1 U11433 ( .A1(n9138), .A2(n9137), .ZN(n9094) );
  INV_X1 U11434 ( .A(n9096), .ZN(n9097) );
  NAND2_X1 U11435 ( .A1(n9097), .A2(n13701), .ZN(n9098) );
  MUX2_X1 U11436 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n10717), .Z(n9101) );
  XNOR2_X1 U11437 ( .A(n9101), .B(n13699), .ZN(n9125) );
  NOR2_X1 U11438 ( .A1(n9101), .A2(SI_29_), .ZN(n9102) );
  INV_X1 U11439 ( .A(n9116), .ZN(n9103) );
  INV_X1 U11440 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13040) );
  INV_X1 U11441 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13038) );
  MUX2_X1 U11442 ( .A(n13040), .B(n13038), .S(n10717), .Z(n9117) );
  XNOR2_X1 U11443 ( .A(n9117), .B(SI_30_), .ZN(n9115) );
  NAND2_X1 U11444 ( .A1(n12705), .A2(n6681), .ZN(n9105) );
  OR2_X1 U11445 ( .A1(n8469), .A2(n13038), .ZN(n9104) );
  INV_X1 U11446 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n14281) );
  NAND2_X1 U11447 ( .A1(n8542), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9107) );
  NAND2_X1 U11448 ( .A1(n9109), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9106) );
  OAI211_X1 U11449 ( .C1(n9112), .C2(n14281), .A(n9107), .B(n9106), .ZN(n14052) );
  AND2_X1 U11450 ( .A1(n14052), .A2(n9114), .ZN(n9154) );
  INV_X1 U11451 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n14285) );
  NAND2_X1 U11452 ( .A1(n8542), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9111) );
  NAND2_X1 U11453 ( .A1(n9109), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9110) );
  OAI211_X1 U11454 ( .C1(n9112), .C2(n14285), .A(n9111), .B(n9110), .ZN(n13918) );
  OAI21_X1 U11455 ( .B1(n9154), .B2(n9108), .A(n13918), .ZN(n9113) );
  OAI21_X1 U11456 ( .B1(n14377), .B2(n9114), .A(n9113), .ZN(n9151) );
  INV_X1 U11457 ( .A(n14377), .ZN(n9173) );
  NOR2_X1 U11458 ( .A1(n9151), .A2(n9150), .ZN(n9153) );
  NAND2_X1 U11459 ( .A1(n9116), .A2(n9115), .ZN(n9120) );
  INV_X1 U11460 ( .A(n9117), .ZN(n9118) );
  NAND2_X1 U11461 ( .A1(n9118), .A2(SI_30_), .ZN(n9119) );
  NAND2_X1 U11462 ( .A1(n9120), .A2(n9119), .ZN(n9123) );
  MUX2_X1 U11463 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10717), .Z(n9121) );
  XNOR2_X1 U11464 ( .A(n9121), .B(SI_31_), .ZN(n9122) );
  XNOR2_X1 U11465 ( .A(n14373), .B(n14052), .ZN(n9190) );
  NAND2_X1 U11466 ( .A1(n12860), .A2(n6681), .ZN(n9128) );
  OR2_X1 U11467 ( .A1(n8469), .A2(n14411), .ZN(n9127) );
  NAND2_X1 U11468 ( .A1(n8514), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n9136) );
  INV_X1 U11469 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n9129) );
  OR2_X1 U11470 ( .A1(n8643), .A2(n9129), .ZN(n9135) );
  OR2_X1 U11471 ( .A1(n9130), .A2(n14062), .ZN(n9134) );
  INV_X1 U11472 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n9131) );
  OR2_X1 U11473 ( .A1(n9132), .A2(n9131), .ZN(n9133) );
  OAI22_X1 U11474 ( .A1(n14291), .A2(n9114), .B1(n6673), .B2(n13809), .ZN(
        n9148) );
  AOI22_X1 U11475 ( .A1(n9775), .A2(n9114), .B1(n6673), .B2(n13919), .ZN(n9149) );
  NOR2_X1 U11476 ( .A1(n9138), .A2(n9137), .ZN(n9143) );
  INV_X1 U11477 ( .A(n9139), .ZN(n9142) );
  INV_X1 U11478 ( .A(n9140), .ZN(n9141) );
  AOI22_X1 U11479 ( .A1(n9144), .A2(n9143), .B1(n9142), .B2(n9141), .ZN(n9145)
         );
  OAI21_X1 U11480 ( .B1(n9148), .B2(n9149), .A(n9145), .ZN(n9146) );
  AOI22_X1 U11481 ( .A1(n9151), .A2(n9150), .B1(n9149), .B2(n9148), .ZN(n9152)
         );
  NOR2_X1 U11482 ( .A1(n9154), .A2(n6673), .ZN(n9156) );
  AND2_X1 U11483 ( .A1(n6673), .A2(n14052), .ZN(n9155) );
  MUX2_X1 U11484 ( .A(n9156), .B(n9155), .S(n14373), .Z(n9157) );
  INV_X1 U11485 ( .A(n9157), .ZN(n9158) );
  NAND2_X1 U11486 ( .A1(n6727), .A2(n9158), .ZN(n9159) );
  INV_X1 U11487 ( .A(n9172), .ZN(n9164) );
  INV_X1 U11488 ( .A(n9748), .ZN(n12464) );
  MUX2_X1 U11489 ( .A(n7046), .B(n12464), .S(n10963), .Z(n9163) );
  NAND2_X1 U11490 ( .A1(n9164), .A2(n7745), .ZN(n9171) );
  NAND2_X1 U11491 ( .A1(n9194), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9165) );
  XNOR2_X1 U11492 ( .A(n9165), .B(P2_IR_REG_23__SCAN_IN), .ZN(n10762) );
  AND2_X1 U11493 ( .A1(n10762), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9193) );
  INV_X1 U11494 ( .A(n9684), .ZN(n9167) );
  OAI211_X1 U11495 ( .C1(n14272), .C2(n12464), .A(n9773), .B(n9167), .ZN(n9168) );
  INV_X1 U11496 ( .A(n9168), .ZN(n9169) );
  NAND2_X1 U11497 ( .A1(n9172), .A2(n9169), .ZN(n9170) );
  NAND3_X1 U11498 ( .A1(n9171), .A2(n9193), .A3(n9170), .ZN(n9207) );
  XOR2_X1 U11499 ( .A(n13918), .B(n9173), .Z(n9189) );
  XNOR2_X1 U11500 ( .A(n9775), .B(n13919), .ZN(n9737) );
  INV_X1 U11501 ( .A(n13920), .ZN(n13763) );
  NAND2_X1 U11502 ( .A1(n14292), .A2(n13763), .ZN(n9174) );
  INV_X1 U11503 ( .A(n13922), .ZN(n13764) );
  OR2_X1 U11504 ( .A1(n14108), .A2(n13764), .ZN(n9733) );
  NAND2_X1 U11505 ( .A1(n14108), .A2(n13764), .ZN(n9734) );
  NAND2_X1 U11506 ( .A1(n9733), .A2(n9734), .ZN(n14102) );
  INV_X1 U11507 ( .A(n13923), .ZN(n13856) );
  XNOR2_X1 U11508 ( .A(n14310), .B(n13856), .ZN(n14117) );
  INV_X1 U11509 ( .A(n13924), .ZN(n9729) );
  XNOR2_X1 U11510 ( .A(n14316), .B(n9729), .ZN(n9677) );
  XNOR2_X1 U11511 ( .A(n14159), .B(n13925), .ZN(n14144) );
  XOR2_X1 U11512 ( .A(n14345), .B(n13929), .Z(n14222) );
  XNOR2_X1 U11513 ( .A(n14341), .B(n9722), .ZN(n14194) );
  INV_X1 U11514 ( .A(n13930), .ZN(n13840) );
  XNOR2_X1 U11515 ( .A(n14353), .B(n13840), .ZN(n14238) );
  XNOR2_X1 U11516 ( .A(n14359), .B(n13931), .ZN(n14244) );
  INV_X1 U11517 ( .A(n13934), .ZN(n9175) );
  XNOR2_X1 U11518 ( .A(n15280), .B(n9175), .ZN(n15267) );
  INV_X1 U11519 ( .A(n13936), .ZN(n9707) );
  XNOR2_X1 U11520 ( .A(n12191), .B(n9707), .ZN(n12042) );
  INV_X1 U11521 ( .A(n13935), .ZN(n9176) );
  OR2_X1 U11522 ( .A1(n12394), .A2(n9176), .ZN(n9709) );
  NAND2_X1 U11523 ( .A1(n12394), .A2(n9176), .ZN(n9710) );
  NAND2_X1 U11524 ( .A1(n9709), .A2(n9710), .ZN(n12196) );
  XNOR2_X1 U11525 ( .A(n11991), .B(n13938), .ZN(n11859) );
  INV_X1 U11526 ( .A(n13940), .ZN(n11759) );
  INV_X1 U11527 ( .A(n13941), .ZN(n11746) );
  XNOR2_X1 U11528 ( .A(n11534), .B(n11746), .ZN(n11526) );
  INV_X1 U11529 ( .A(n13942), .ZN(n11488) );
  XNOR2_X1 U11530 ( .A(n11395), .B(n11488), .ZN(n11388) );
  XNOR2_X1 U11531 ( .A(n11590), .B(n13943), .ZN(n11328) );
  OR2_X1 U11532 ( .A1(n13947), .A2(n15691), .ZN(n9177) );
  NAND2_X1 U11533 ( .A1(n13947), .A2(n15691), .ZN(n11841) );
  AND2_X1 U11534 ( .A1(n9177), .A2(n11841), .ZN(n15693) );
  NOR4_X1 U11535 ( .A1(n15693), .A2(n11842), .A3(n10889), .A4(n12707), .ZN(
        n9179) );
  NAND4_X1 U11536 ( .A1(n11328), .A2(n9179), .A3(n11093), .A4(n11568), .ZN(
        n9180) );
  NOR4_X1 U11537 ( .A1(n11647), .A2(n11526), .A3(n11388), .A4(n9180), .ZN(
        n9181) );
  XNOR2_X1 U11538 ( .A(n12105), .B(n13937), .ZN(n11892) );
  XNOR2_X1 U11539 ( .A(n11879), .B(n13939), .ZN(n11806) );
  NAND4_X1 U11540 ( .A1(n11859), .A2(n9181), .A3(n11892), .A4(n11806), .ZN(
        n9182) );
  NOR4_X1 U11541 ( .A1(n15267), .A2(n12042), .A3(n12196), .A4(n9182), .ZN(
        n9183) );
  XNOR2_X1 U11542 ( .A(n14364), .B(n13932), .ZN(n14274) );
  XNOR2_X1 U11543 ( .A(n12570), .B(n13933), .ZN(n12486) );
  NAND4_X1 U11544 ( .A1(n14244), .A2(n9183), .A3(n14274), .A4(n12486), .ZN(
        n9184) );
  NOR4_X1 U11545 ( .A1(n14222), .A2(n14194), .A3(n14238), .A4(n9184), .ZN(
        n9185) );
  XNOR2_X1 U11546 ( .A(n14394), .B(n13926), .ZN(n9674) );
  XNOR2_X1 U11547 ( .A(n14337), .B(n13927), .ZN(n14179) );
  NAND4_X1 U11548 ( .A1(n14144), .A2(n9185), .A3(n9674), .A4(n14179), .ZN(
        n9186) );
  NOR4_X1 U11549 ( .A1(n14102), .A2(n14117), .A3(n9677), .A4(n9186), .ZN(n9187) );
  NAND4_X1 U11550 ( .A1(n9737), .A2(n14072), .A3(n9187), .A4(n14088), .ZN(
        n9188) );
  NOR3_X1 U11551 ( .A1(n9190), .A2(n9189), .A3(n9188), .ZN(n9191) );
  NAND2_X1 U11552 ( .A1(n9192), .A2(n7766), .ZN(n9206) );
  NAND2_X1 U11553 ( .A1(n9197), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9198) );
  MUX2_X1 U11554 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9198), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9199) );
  NAND2_X1 U11555 ( .A1(n9199), .A2(n6814), .ZN(n14427) );
  NAND2_X1 U11556 ( .A1(n6814), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9200) );
  MUX2_X1 U11557 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9200), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n9201) );
  INV_X1 U11558 ( .A(n10762), .ZN(n9202) );
  NAND2_X1 U11559 ( .A1(n10507), .A2(n9202), .ZN(n9765) );
  NAND2_X1 U11560 ( .A1(n9748), .A2(n9747), .ZN(n10761) );
  INV_X1 U11561 ( .A(n9773), .ZN(n10967) );
  NOR2_X1 U11562 ( .A1(n10761), .A2(n10967), .ZN(n9768) );
  NOR2_X1 U11563 ( .A1(n9765), .A2(n9768), .ZN(n10960) );
  NOR2_X1 U11564 ( .A1(n10767), .A2(P2_U3088), .ZN(n14420) );
  INV_X1 U11565 ( .A(n10761), .ZN(n10955) );
  INV_X1 U11566 ( .A(n9203), .ZN(n10765) );
  NAND3_X1 U11567 ( .A1(n10960), .A2(n14420), .A3(n13906), .ZN(n9204) );
  OAI211_X1 U11568 ( .C1(n9747), .C2(n9166), .A(n9204), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9205) );
  NAND3_X1 U11569 ( .A1(n9207), .A2(n9206), .A3(n9205), .ZN(P2_U3328) );
  INV_X1 U11570 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9301) );
  INV_X1 U11571 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n15145) );
  INV_X1 U11572 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15490) );
  NOR2_X1 U11573 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n15490), .ZN(n9241) );
  INV_X1 U11574 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9240) );
  XOR2_X1 U11575 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .Z(n9251) );
  INV_X1 U11576 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n9238) );
  INV_X1 U11577 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n9235) );
  XNOR2_X1 U11578 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(P3_ADDR_REG_12__SCAN_IN), 
        .ZN(n9252) );
  INV_X1 U11579 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n15736) );
  XNOR2_X1 U11580 ( .A(P1_ADDR_REG_11__SCAN_IN), .B(P3_ADDR_REG_11__SCAN_IN), 
        .ZN(n9254) );
  INV_X1 U11581 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9229) );
  XOR2_X1 U11582 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n9582), .Z(n9258) );
  INV_X1 U11583 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n9565) );
  XNOR2_X1 U11584 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(P3_ADDR_REG_8__SCAN_IN), 
        .ZN(n9260) );
  INV_X1 U11585 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n9222) );
  XNOR2_X1 U11586 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n9278) );
  NAND2_X1 U11587 ( .A1(n9264), .A2(n9265), .ZN(n9210) );
  NAND2_X1 U11588 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n9212), .ZN(n9214) );
  INV_X1 U11589 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9213) );
  NAND2_X1 U11590 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n9215), .ZN(n9217) );
  INV_X1 U11591 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n15475) );
  NAND2_X1 U11592 ( .A1(n9262), .A2(n15475), .ZN(n9216) );
  NAND2_X1 U11593 ( .A1(n9217), .A2(n9216), .ZN(n9218) );
  NAND2_X1 U11594 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n9218), .ZN(n9220) );
  XNOR2_X1 U11595 ( .A(n9218), .B(n9517), .ZN(n9274) );
  INV_X1 U11596 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14608) );
  NAND2_X1 U11597 ( .A1(n9274), .A2(n14608), .ZN(n9219) );
  NAND2_X1 U11598 ( .A1(n9220), .A2(n9219), .ZN(n9279) );
  NAND2_X1 U11599 ( .A1(n9278), .A2(n9279), .ZN(n9221) );
  NAND2_X1 U11600 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n9223), .ZN(n9226) );
  XOR2_X1 U11601 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n9223), .Z(n9285) );
  INV_X1 U11602 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9224) );
  NAND2_X1 U11603 ( .A1(n9285), .A2(n9224), .ZN(n9225) );
  NAND2_X1 U11604 ( .A1(n9226), .A2(n9225), .ZN(n9261) );
  NAND2_X1 U11605 ( .A1(n9260), .A2(n9261), .ZN(n9227) );
  NAND2_X1 U11606 ( .A1(n9258), .A2(n9259), .ZN(n9228) );
  NOR2_X1 U11607 ( .A1(n9229), .A2(n9257), .ZN(n9232) );
  INV_X1 U11608 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n9231) );
  NAND2_X1 U11609 ( .A1(n9229), .A2(n9257), .ZN(n9230) );
  NAND2_X1 U11610 ( .A1(n9254), .A2(n9255), .ZN(n9233) );
  NAND2_X1 U11611 ( .A1(n9252), .A2(n9253), .ZN(n9234) );
  OAI21_X1 U11612 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n9235), .A(n9234), .ZN(
        n9236) );
  INV_X1 U11613 ( .A(n9236), .ZN(n9298) );
  AND2_X1 U11614 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n9238), .ZN(n9237) );
  OAI22_X1 U11615 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n15145), .B1(n9241), 
        .B2(n9249), .ZN(n9243) );
  INV_X1 U11616 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9242) );
  NOR2_X1 U11617 ( .A1(n9243), .A2(n9242), .ZN(n9245) );
  XOR2_X1 U11618 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n9243), .Z(n9246) );
  NOR2_X1 U11619 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n9246), .ZN(n9244) );
  NOR2_X1 U11620 ( .A1(n9245), .A2(n9244), .ZN(n9302) );
  XNOR2_X1 U11621 ( .A(n9301), .B(n9302), .ZN(n9303) );
  XNOR2_X1 U11622 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n9303), .ZN(n15140) );
  XNOR2_X1 U11623 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n9246), .ZN(n15441) );
  NOR2_X1 U11624 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n15145), .ZN(n9247) );
  AOI21_X1 U11625 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n15145), .A(n9247), .ZN(
        n9248) );
  XNOR2_X1 U11626 ( .A(n9249), .B(n9248), .ZN(n15436) );
  XNOR2_X1 U11627 ( .A(n9251), .B(n9250), .ZN(n15433) );
  XOR2_X1 U11628 ( .A(n9253), .B(n9252), .Z(n15425) );
  XNOR2_X1 U11629 ( .A(n9255), .B(n9254), .ZN(n9295) );
  XOR2_X1 U11630 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(P3_ADDR_REG_10__SCAN_IN), 
        .Z(n9256) );
  XOR2_X1 U11631 ( .A(n9257), .B(n9256), .Z(n9293) );
  XOR2_X1 U11632 ( .A(n9259), .B(n9258), .Z(n9291) );
  XOR2_X1 U11633 ( .A(n9261), .B(n9260), .Z(n9287) );
  AND2_X1 U11634 ( .A1(n9272), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n9273) );
  XNOR2_X1 U11635 ( .A(n9263), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n15867) );
  XOR2_X1 U11636 ( .A(n9265), .B(n9264), .Z(n15117) );
  INV_X1 U11637 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9269) );
  NOR2_X1 U11638 ( .A1(n9268), .A2(n9269), .ZN(n9270) );
  AOI21_X1 U11639 ( .B1(n9574), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n9266), .ZN(
        n15861) );
  INV_X1 U11640 ( .A(n15861), .ZN(n9267) );
  NAND2_X1 U11641 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n9267), .ZN(n15871) );
  XNOR2_X1 U11642 ( .A(n9269), .B(n9268), .ZN(n15870) );
  NOR2_X1 U11643 ( .A1(n15871), .A2(n15870), .ZN(n15869) );
  NAND2_X1 U11644 ( .A1(n15117), .A2(n15116), .ZN(n15115) );
  NAND2_X1 U11645 ( .A1(n15867), .A2(n15866), .ZN(n9271) );
  AOI21_X1 U11646 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n9271), .A(n15865), .ZN(
        n15857) );
  NOR2_X1 U11647 ( .A1(n15857), .A2(n15856), .ZN(n15855) );
  XNOR2_X1 U11648 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n9274), .ZN(n9276) );
  NAND2_X1 U11649 ( .A1(n9275), .A2(n9276), .ZN(n9277) );
  INV_X1 U11650 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15859) );
  INV_X1 U11651 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n9280) );
  NOR2_X1 U11652 ( .A1(n9281), .A2(n9280), .ZN(n9282) );
  XOR2_X1 U11653 ( .A(n9279), .B(n9278), .Z(n15127) );
  NOR2_X1 U11654 ( .A1(n15127), .A2(n15126), .ZN(n15125) );
  INV_X1 U11655 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9284) );
  NAND2_X1 U11656 ( .A1(n9283), .A2(n9284), .ZN(n9286) );
  XNOR2_X1 U11657 ( .A(n9285), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15863) );
  NOR2_X1 U11658 ( .A1(n9287), .A2(n9288), .ZN(n9289) );
  INV_X1 U11659 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n15129) );
  NAND2_X1 U11660 ( .A1(n9291), .A2(n9290), .ZN(n9292) );
  INV_X1 U11661 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n15132) );
  INV_X1 U11662 ( .A(n6730), .ZN(n15135) );
  INV_X1 U11663 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n15137) );
  NAND2_X1 U11664 ( .A1(n9294), .A2(n9293), .ZN(n15136) );
  NAND2_X1 U11665 ( .A1(n15137), .A2(n15136), .ZN(n15134) );
  INV_X1 U11666 ( .A(n15419), .ZN(n15420) );
  INV_X1 U11667 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n15422) );
  NAND2_X1 U11668 ( .A1(n9296), .A2(n9295), .ZN(n15421) );
  NAND2_X1 U11669 ( .A1(n15422), .A2(n15421), .ZN(n15418) );
  NAND2_X1 U11670 ( .A1(n15425), .A2(n15424), .ZN(n9297) );
  XNOR2_X1 U11671 ( .A(P1_ADDR_REG_13__SCAN_IN), .B(P3_ADDR_REG_13__SCAN_IN), 
        .ZN(n9299) );
  XNOR2_X1 U11672 ( .A(n9299), .B(n9298), .ZN(n15429) );
  NAND2_X1 U11673 ( .A1(n15428), .A2(n15429), .ZN(n15427) );
  NAND2_X1 U11674 ( .A1(n15140), .A2(n15139), .ZN(n9300) );
  AOI21_X2 U11675 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(n9300), .A(n15138), .ZN(
        n15111) );
  NAND2_X1 U11676 ( .A1(n9302), .A2(n9301), .ZN(n9306) );
  INV_X1 U11677 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n9304) );
  OR2_X1 U11678 ( .A1(n9304), .A2(n9303), .ZN(n9305) );
  NAND2_X1 U11679 ( .A1(n9306), .A2(n9305), .ZN(n9310) );
  INV_X1 U11680 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n9313) );
  NOR2_X1 U11681 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n9313), .ZN(n9307) );
  AOI21_X1 U11682 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9313), .A(n9307), .ZN(
        n9311) );
  XOR2_X1 U11683 ( .A(n9310), .B(n9311), .Z(n15110) );
  XNOR2_X1 U11684 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n9308) );
  XNOR2_X1 U11685 ( .A(n9308), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n9309) );
  NAND2_X1 U11686 ( .A1(n9311), .A2(n9310), .ZN(n9312) );
  OAI21_X1 U11687 ( .B1(n9313), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n9312), .ZN(
        n9644) );
  INV_X1 U11688 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n11280) );
  XOR2_X1 U11689 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(keyinput_g82), .Z(n9320)
         );
  AOI22_X1 U11690 ( .A1(SI_31_), .A2(keyinput_g1), .B1(P3_REG3_REG_8__SCAN_IN), 
        .B2(keyinput_g43), .ZN(n9314) );
  OAI221_X1 U11691 ( .B1(SI_31_), .B2(keyinput_g1), .C1(P3_REG3_REG_8__SCAN_IN), .C2(keyinput_g43), .A(n9314), .ZN(n9319) );
  AOI22_X1 U11692 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput_g116), .B1(SI_25_), 
        .B2(keyinput_g7), .ZN(n9315) );
  OAI221_X1 U11693 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput_g116), .C1(SI_25_), .C2(keyinput_g7), .A(n9315), .ZN(n9318) );
  AOI22_X1 U11694 ( .A1(SI_26_), .A2(keyinput_g6), .B1(P3_REG3_REG_5__SCAN_IN), 
        .B2(keyinput_g49), .ZN(n9316) );
  OAI221_X1 U11695 ( .B1(SI_26_), .B2(keyinput_g6), .C1(P3_REG3_REG_5__SCAN_IN), .C2(keyinput_g49), .A(n9316), .ZN(n9317) );
  NOR4_X1 U11696 ( .A1(n9320), .A2(n9319), .A3(n9318), .A4(n9317), .ZN(n9348)
         );
  AOI22_X1 U11697 ( .A1(P3_DATAO_REG_28__SCAN_IN), .A2(keyinput_g68), .B1(
        P3_RD_REG_SCAN_IN), .B2(keyinput_g33), .ZN(n9321) );
  OAI221_X1 U11698 ( .B1(P3_DATAO_REG_28__SCAN_IN), .B2(keyinput_g68), .C1(
        P3_RD_REG_SCAN_IN), .C2(keyinput_g33), .A(n9321), .ZN(n9328) );
  AOI22_X1 U11699 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(keyinput_g35), .B1(
        P3_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .ZN(n9322) );
  OAI221_X1 U11700 ( .B1(P3_REG3_REG_7__SCAN_IN), .B2(keyinput_g35), .C1(
        P3_REG3_REG_10__SCAN_IN), .C2(keyinput_g39), .A(n9322), .ZN(n9327) );
  AOI22_X1 U11701 ( .A1(P3_DATAO_REG_2__SCAN_IN), .A2(keyinput_g94), .B1(
        P3_DATAO_REG_25__SCAN_IN), .B2(keyinput_g71), .ZN(n9323) );
  OAI221_X1 U11702 ( .B1(P3_DATAO_REG_2__SCAN_IN), .B2(keyinput_g94), .C1(
        P3_DATAO_REG_25__SCAN_IN), .C2(keyinput_g71), .A(n9323), .ZN(n9326) );
  AOI22_X1 U11703 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput_g110), .B1(
        P3_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .ZN(n9324) );
  OAI221_X1 U11704 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput_g110), .C1(
        P3_REG3_REG_11__SCAN_IN), .C2(keyinput_g58), .A(n9324), .ZN(n9325) );
  NOR4_X1 U11705 ( .A1(n9328), .A2(n9327), .A3(n9326), .A4(n9325), .ZN(n9347)
         );
  AOI22_X1 U11706 ( .A1(P3_DATAO_REG_11__SCAN_IN), .A2(keyinput_g85), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .ZN(n9329) );
  OAI221_X1 U11707 ( .B1(P3_DATAO_REG_11__SCAN_IN), .B2(keyinput_g85), .C1(
        P3_REG3_REG_2__SCAN_IN), .C2(keyinput_g59), .A(n9329), .ZN(n9336) );
  AOI22_X1 U11708 ( .A1(P3_DATAO_REG_21__SCAN_IN), .A2(keyinput_g75), .B1(
        SI_15_), .B2(keyinput_g17), .ZN(n9330) );
  OAI221_X1 U11709 ( .B1(P3_DATAO_REG_21__SCAN_IN), .B2(keyinput_g75), .C1(
        SI_15_), .C2(keyinput_g17), .A(n9330), .ZN(n9335) );
  AOI22_X1 U11710 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput_g108), .B1(SI_17_), 
        .B2(keyinput_g15), .ZN(n9331) );
  OAI221_X1 U11711 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput_g108), .C1(SI_17_), .C2(keyinput_g15), .A(n9331), .ZN(n9334) );
  AOI22_X1 U11712 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput_g112), .B1(
        P3_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .ZN(n9332) );
  OAI221_X1 U11713 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput_g112), .C1(
        P3_REG3_REG_17__SCAN_IN), .C2(keyinput_g50), .A(n9332), .ZN(n9333) );
  NOR4_X1 U11714 ( .A1(n9336), .A2(n9335), .A3(n9334), .A4(n9333), .ZN(n9346)
         );
  AOI22_X1 U11715 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(keyinput_g100), .B1(SI_6_), .B2(keyinput_g26), .ZN(n9337) );
  OAI221_X1 U11716 ( .B1(P3_ADDR_REG_3__SCAN_IN), .B2(keyinput_g100), .C1(
        SI_6_), .C2(keyinput_g26), .A(n9337), .ZN(n9344) );
  AOI22_X1 U11717 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(keyinput_g122), .B1(SI_4_), 
        .B2(keyinput_g28), .ZN(n9338) );
  OAI221_X1 U11718 ( .B1(P1_IR_REG_15__SCAN_IN), .B2(keyinput_g122), .C1(SI_4_), .C2(keyinput_g28), .A(n9338), .ZN(n9343) );
  AOI22_X1 U11719 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput_g115), .B1(
        P1_IR_REG_7__SCAN_IN), .B2(keyinput_g114), .ZN(n9339) );
  OAI221_X1 U11720 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(keyinput_g115), .C1(
        P1_IR_REG_7__SCAN_IN), .C2(keyinput_g114), .A(n9339), .ZN(n9342) );
  AOI22_X1 U11721 ( .A1(SI_19_), .A2(keyinput_g13), .B1(
        P3_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .ZN(n9340) );
  OAI221_X1 U11722 ( .B1(SI_19_), .B2(keyinput_g13), .C1(
        P3_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(n9340), .ZN(n9341) );
  NOR4_X1 U11723 ( .A1(n9344), .A2(n9343), .A3(n9342), .A4(n9341), .ZN(n9345)
         );
  NAND4_X1 U11724 ( .A1(n9348), .A2(n9347), .A3(n9346), .A4(n9345), .ZN(n9469)
         );
  AOI22_X1 U11725 ( .A1(P3_DATAO_REG_13__SCAN_IN), .A2(keyinput_g83), .B1(
        SI_3_), .B2(keyinput_g29), .ZN(n9349) );
  OAI221_X1 U11726 ( .B1(P3_DATAO_REG_13__SCAN_IN), .B2(keyinput_g83), .C1(
        SI_3_), .C2(keyinput_g29), .A(n9349), .ZN(n9356) );
  AOI22_X1 U11727 ( .A1(P3_DATAO_REG_27__SCAN_IN), .A2(keyinput_g69), .B1(
        SI_30_), .B2(keyinput_g2), .ZN(n9350) );
  OAI221_X1 U11728 ( .B1(P3_DATAO_REG_27__SCAN_IN), .B2(keyinput_g69), .C1(
        SI_30_), .C2(keyinput_g2), .A(n9350), .ZN(n9355) );
  AOI22_X1 U11729 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(keyinput_g99), .B1(
        P3_ADDR_REG_6__SCAN_IN), .B2(keyinput_g103), .ZN(n9351) );
  OAI221_X1 U11730 ( .B1(P3_ADDR_REG_2__SCAN_IN), .B2(keyinput_g99), .C1(
        P3_ADDR_REG_6__SCAN_IN), .C2(keyinput_g103), .A(n9351), .ZN(n9354) );
  AOI22_X1 U11731 ( .A1(P3_DATAO_REG_22__SCAN_IN), .A2(keyinput_g74), .B1(
        P3_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .ZN(n9352) );
  OAI221_X1 U11732 ( .B1(P3_DATAO_REG_22__SCAN_IN), .B2(keyinput_g74), .C1(
        P3_REG3_REG_20__SCAN_IN), .C2(keyinput_g55), .A(n9352), .ZN(n9353) );
  NOR4_X1 U11733 ( .A1(n9356), .A2(n9355), .A3(n9354), .A4(n9353), .ZN(n9385)
         );
  AOI22_X1 U11734 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(keyinput_g104), .B1(SI_9_), .B2(keyinput_g23), .ZN(n9357) );
  OAI221_X1 U11735 ( .B1(P3_ADDR_REG_7__SCAN_IN), .B2(keyinput_g104), .C1(
        SI_9_), .C2(keyinput_g23), .A(n9357), .ZN(n9364) );
  AOI22_X1 U11736 ( .A1(SI_13_), .A2(keyinput_g19), .B1(SI_22_), .B2(
        keyinput_g10), .ZN(n9358) );
  OAI221_X1 U11737 ( .B1(SI_13_), .B2(keyinput_g19), .C1(SI_22_), .C2(
        keyinput_g10), .A(n9358), .ZN(n9363) );
  AOI22_X1 U11738 ( .A1(P3_DATAO_REG_16__SCAN_IN), .A2(keyinput_g80), .B1(
        SI_29_), .B2(keyinput_g3), .ZN(n9359) );
  OAI221_X1 U11739 ( .B1(P3_DATAO_REG_16__SCAN_IN), .B2(keyinput_g80), .C1(
        SI_29_), .C2(keyinput_g3), .A(n9359), .ZN(n9362) );
  AOI22_X1 U11740 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput_g126), .B1(
        P3_REG3_REG_21__SCAN_IN), .B2(keyinput_g45), .ZN(n9360) );
  OAI221_X1 U11741 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(keyinput_g126), .C1(
        P3_REG3_REG_21__SCAN_IN), .C2(keyinput_g45), .A(n9360), .ZN(n9361) );
  NOR4_X1 U11742 ( .A1(n9364), .A2(n9363), .A3(n9362), .A4(n9361), .ZN(n9384)
         );
  AOI22_X1 U11743 ( .A1(P3_DATAO_REG_9__SCAN_IN), .A2(keyinput_g87), .B1(
        P1_IR_REG_18__SCAN_IN), .B2(keyinput_g125), .ZN(n9365) );
  OAI221_X1 U11744 ( .B1(P3_DATAO_REG_9__SCAN_IN), .B2(keyinput_g87), .C1(
        P1_IR_REG_18__SCAN_IN), .C2(keyinput_g125), .A(n9365), .ZN(n9372) );
  AOI22_X1 U11745 ( .A1(P3_ADDR_REG_8__SCAN_IN), .A2(keyinput_g105), .B1(
        P1_IR_REG_14__SCAN_IN), .B2(keyinput_g121), .ZN(n9366) );
  OAI221_X1 U11746 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(keyinput_g105), .C1(
        P1_IR_REG_14__SCAN_IN), .C2(keyinput_g121), .A(n9366), .ZN(n9371) );
  AOI22_X1 U11747 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(keyinput_g109), .B1(
        P1_IR_REG_20__SCAN_IN), .B2(keyinput_g127), .ZN(n9367) );
  OAI221_X1 U11748 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(keyinput_g109), .C1(
        P1_IR_REG_20__SCAN_IN), .C2(keyinput_g127), .A(n9367), .ZN(n9370) );
  AOI22_X1 U11749 ( .A1(SI_10_), .A2(keyinput_g22), .B1(P3_REG3_REG_3__SCAN_IN), .B2(keyinput_g40), .ZN(n9368) );
  OAI221_X1 U11750 ( .B1(SI_10_), .B2(keyinput_g22), .C1(
        P3_REG3_REG_3__SCAN_IN), .C2(keyinput_g40), .A(n9368), .ZN(n9369) );
  NOR4_X1 U11751 ( .A1(n9372), .A2(n9371), .A3(n9370), .A4(n9369), .ZN(n9383)
         );
  AOI22_X1 U11752 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(keyinput_g44), .B1(
        P3_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .ZN(n9373) );
  OAI221_X1 U11753 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput_g60), .A(n9373), .ZN(n9381) );
  INV_X1 U11754 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n11454) );
  AOI22_X1 U11755 ( .A1(SI_21_), .A2(keyinput_g11), .B1(n11454), .B2(
        keyinput_g86), .ZN(n9374) );
  OAI221_X1 U11756 ( .B1(SI_21_), .B2(keyinput_g11), .C1(n11454), .C2(
        keyinput_g86), .A(n9374), .ZN(n9380) );
  INV_X1 U11757 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9539) );
  AOI22_X1 U11758 ( .A1(n12431), .A2(keyinput_g46), .B1(keyinput_g117), .B2(
        n9539), .ZN(n9375) );
  OAI221_X1 U11759 ( .B1(n12431), .B2(keyinput_g46), .C1(n9539), .C2(
        keyinput_g117), .A(n9375), .ZN(n9379) );
  INV_X1 U11760 ( .A(P3_WR_REG_SCAN_IN), .ZN(n9377) );
  AOI22_X1 U11761 ( .A1(n9377), .A2(keyinput_g0), .B1(n10728), .B2(
        keyinput_g31), .ZN(n9376) );
  OAI221_X1 U11762 ( .B1(n9377), .B2(keyinput_g0), .C1(n10728), .C2(
        keyinput_g31), .A(n9376), .ZN(n9378) );
  NOR4_X1 U11763 ( .A1(n9381), .A2(n9380), .A3(n9379), .A4(n9378), .ZN(n9382)
         );
  NAND4_X1 U11764 ( .A1(n9385), .A2(n9384), .A3(n9383), .A4(n9382), .ZN(n9468)
         );
  INV_X1 U11765 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9525) );
  AOI22_X1 U11766 ( .A1(n9525), .A2(keyinput_g47), .B1(keyinput_g102), .B2(
        n9517), .ZN(n9386) );
  OAI221_X1 U11767 ( .B1(n9525), .B2(keyinput_g47), .C1(n9517), .C2(
        keyinput_g102), .A(n9386), .ZN(n9395) );
  INV_X1 U11768 ( .A(SI_0_), .ZN(n9388) );
  AOI22_X1 U11769 ( .A1(n12498), .A2(keyinput_g8), .B1(keyinput_g32), .B2(
        n9388), .ZN(n9387) );
  OAI221_X1 U11770 ( .B1(n12498), .B2(keyinput_g8), .C1(n9388), .C2(
        keyinput_g32), .A(n9387), .ZN(n9394) );
  INV_X1 U11771 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n11359) );
  INV_X1 U11772 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n11726) );
  AOI22_X1 U11773 ( .A1(n11359), .A2(keyinput_g79), .B1(n11726), .B2(
        keyinput_g65), .ZN(n9389) );
  OAI221_X1 U11774 ( .B1(n11359), .B2(keyinput_g79), .C1(n11726), .C2(
        keyinput_g65), .A(n9389), .ZN(n9393) );
  XOR2_X1 U11775 ( .A(n9574), .B(keyinput_g97), .Z(n9391) );
  XNOR2_X1 U11776 ( .A(SI_2_), .B(keyinput_g30), .ZN(n9390) );
  NAND2_X1 U11777 ( .A1(n9391), .A2(n9390), .ZN(n9392) );
  NOR4_X1 U11778 ( .A1(n9395), .A2(n9394), .A3(n9393), .A4(n9392), .ZN(n9427)
         );
  INV_X1 U11779 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9397) );
  INV_X1 U11780 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n11361) );
  AOI22_X1 U11781 ( .A1(n9397), .A2(keyinput_g120), .B1(keyinput_g91), .B2(
        n11361), .ZN(n9396) );
  OAI221_X1 U11782 ( .B1(n9397), .B2(keyinput_g120), .C1(n11361), .C2(
        keyinput_g91), .A(n9396), .ZN(n9405) );
  INV_X1 U11783 ( .A(P3_DATAO_REG_6__SCAN_IN), .ZN(n11363) );
  AOI22_X1 U11784 ( .A1(n8344), .A2(keyinput_g64), .B1(keyinput_g90), .B2(
        n11363), .ZN(n9398) );
  OAI221_X1 U11785 ( .B1(n8344), .B2(keyinput_g64), .C1(n11363), .C2(
        keyinput_g90), .A(n9398), .ZN(n9404) );
  INV_X1 U11786 ( .A(SI_14_), .ZN(n10849) );
  AOI22_X1 U11787 ( .A1(n10849), .A2(keyinput_g18), .B1(n7860), .B2(
        keyinput_g62), .ZN(n9399) );
  OAI221_X1 U11788 ( .B1(n10849), .B2(keyinput_g18), .C1(n7860), .C2(
        keyinput_g62), .A(n9399), .ZN(n9403) );
  XOR2_X1 U11789 ( .A(n10128), .B(keyinput_g118), .Z(n9401) );
  XNOR2_X1 U11790 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_g107), .ZN(n9400) );
  NAND2_X1 U11791 ( .A1(n9401), .A2(n9400), .ZN(n9402) );
  NOR4_X1 U11792 ( .A1(n9405), .A2(n9404), .A3(n9403), .A4(n9402), .ZN(n9426)
         );
  INV_X1 U11793 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n11288) );
  AOI22_X1 U11794 ( .A1(n9407), .A2(keyinput_g101), .B1(n11288), .B2(
        keyinput_g61), .ZN(n9406) );
  OAI221_X1 U11795 ( .B1(n9407), .B2(keyinput_g101), .C1(n11288), .C2(
        keyinput_g61), .A(n9406), .ZN(n9414) );
  INV_X1 U11796 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n11731) );
  AOI22_X1 U11797 ( .A1(n11731), .A2(keyinput_g67), .B1(n7261), .B2(
        keyinput_g124), .ZN(n9408) );
  OAI221_X1 U11798 ( .B1(n11731), .B2(keyinput_g67), .C1(n7261), .C2(
        keyinput_g124), .A(n9408), .ZN(n9413) );
  INV_X1 U11799 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n11402) );
  AOI22_X1 U11800 ( .A1(n7986), .A2(keyinput_g53), .B1(keyinput_g95), .B2(
        n11402), .ZN(n9409) );
  OAI221_X1 U11801 ( .B1(n7986), .B2(keyinput_g53), .C1(n11402), .C2(
        keyinput_g95), .A(n9409), .ZN(n9412) );
  INV_X1 U11802 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n11278) );
  INV_X1 U11803 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n11165) );
  AOI22_X1 U11804 ( .A1(n11278), .A2(keyinput_g76), .B1(keyinput_g73), .B2(
        n11165), .ZN(n9410) );
  OAI221_X1 U11805 ( .B1(n11278), .B2(keyinput_g76), .C1(n11165), .C2(
        keyinput_g73), .A(n9410), .ZN(n9411) );
  NOR4_X1 U11806 ( .A1(n9414), .A2(n9413), .A3(n9412), .A4(n9411), .ZN(n9425)
         );
  INV_X1 U11807 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n12975) );
  AOI22_X1 U11808 ( .A1(P3_U3151), .A2(keyinput_g34), .B1(keyinput_g56), .B2(
        n12975), .ZN(n9415) );
  OAI221_X1 U11809 ( .B1(P3_U3151), .B2(keyinput_g34), .C1(n12975), .C2(
        keyinput_g56), .A(n9415), .ZN(n9423) );
  INV_X1 U11810 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n11728) );
  INV_X1 U11811 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n11276) );
  AOI22_X1 U11812 ( .A1(n11728), .A2(keyinput_g66), .B1(keyinput_g78), .B2(
        n11276), .ZN(n9416) );
  OAI221_X1 U11813 ( .B1(n11728), .B2(keyinput_g66), .C1(n11276), .C2(
        keyinput_g78), .A(n9416), .ZN(n9422) );
  INV_X1 U11814 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n9586) );
  AOI22_X1 U11815 ( .A1(n11661), .A2(keyinput_g12), .B1(n9586), .B2(
        keyinput_g38), .ZN(n9417) );
  OAI221_X1 U11816 ( .B1(n11661), .B2(keyinput_g12), .C1(n9586), .C2(
        keyinput_g38), .A(n9417), .ZN(n9421) );
  XNOR2_X1 U11817 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_g111), .ZN(n9419) );
  XNOR2_X1 U11818 ( .A(SI_23_), .B(keyinput_g9), .ZN(n9418) );
  NAND2_X1 U11819 ( .A1(n9419), .A2(n9418), .ZN(n9420) );
  NOR4_X1 U11820 ( .A1(n9423), .A2(n9422), .A3(n9421), .A4(n9420), .ZN(n9424)
         );
  NAND4_X1 U11821 ( .A1(n9427), .A2(n9426), .A3(n9425), .A4(n9424), .ZN(n9467)
         );
  INV_X1 U11822 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n11399) );
  AOI22_X1 U11823 ( .A1(n11399), .A2(keyinput_g93), .B1(n13701), .B2(
        keyinput_g4), .ZN(n9428) );
  OAI221_X1 U11824 ( .B1(n11399), .B2(keyinput_g93), .C1(n13701), .C2(
        keyinput_g4), .A(n9428), .ZN(n9435) );
  AOI22_X1 U11825 ( .A1(n10701), .A2(keyinput_g27), .B1(keyinput_g106), .B2(
        n9582), .ZN(n9429) );
  OAI221_X1 U11826 ( .B1(n10701), .B2(keyinput_g27), .C1(n9582), .C2(
        keyinput_g106), .A(n9429), .ZN(n9434) );
  INV_X1 U11827 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n11371) );
  INV_X1 U11828 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9878) );
  AOI22_X1 U11829 ( .A1(n11371), .A2(keyinput_g89), .B1(n9878), .B2(
        keyinput_g36), .ZN(n9430) );
  OAI221_X1 U11830 ( .B1(n11371), .B2(keyinput_g89), .C1(n9878), .C2(
        keyinput_g36), .A(n9430), .ZN(n9433) );
  INV_X1 U11831 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n11324) );
  AOI22_X1 U11832 ( .A1(n10975), .A2(keyinput_g16), .B1(keyinput_g72), .B2(
        n11324), .ZN(n9431) );
  OAI221_X1 U11833 ( .B1(n10975), .B2(keyinput_g16), .C1(n11324), .C2(
        keyinput_g72), .A(n9431), .ZN(n9432) );
  NOR4_X1 U11834 ( .A1(n9435), .A2(n9434), .A3(n9433), .A4(n9432), .ZN(n9465)
         );
  INV_X1 U11835 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n10983) );
  AOI22_X1 U11836 ( .A1(n11183), .A2(keyinput_g14), .B1(keyinput_g77), .B2(
        n10983), .ZN(n9436) );
  OAI221_X1 U11837 ( .B1(n11183), .B2(keyinput_g14), .C1(n10983), .C2(
        keyinput_g77), .A(n9436), .ZN(n9444) );
  INV_X1 U11838 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9562) );
  INV_X1 U11839 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n13025) );
  AOI22_X1 U11840 ( .A1(n9562), .A2(keyinput_g119), .B1(n13025), .B2(
        keyinput_g63), .ZN(n9437) );
  OAI221_X1 U11841 ( .B1(n9562), .B2(keyinput_g119), .C1(n13025), .C2(
        keyinput_g63), .A(n9437), .ZN(n9443) );
  INV_X1 U11842 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n12894) );
  AOI22_X1 U11843 ( .A1(n10742), .A2(keyinput_g20), .B1(n12894), .B2(
        keyinput_g41), .ZN(n9438) );
  OAI221_X1 U11844 ( .B1(n10742), .B2(keyinput_g20), .C1(n12894), .C2(
        keyinput_g41), .A(n9438), .ZN(n9442) );
  XNOR2_X1 U11845 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_g113), .ZN(n9440) );
  XNOR2_X1 U11846 ( .A(P3_REG3_REG_4__SCAN_IN), .B(keyinput_g52), .ZN(n9439)
         );
  NAND2_X1 U11847 ( .A1(n9440), .A2(n9439), .ZN(n9441) );
  NOR4_X1 U11848 ( .A1(n9444), .A2(n9443), .A3(n9442), .A4(n9441), .ZN(n9464)
         );
  INV_X1 U11849 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n12959) );
  AOI22_X1 U11850 ( .A1(n12959), .A2(keyinput_g51), .B1(keyinput_g24), .B2(
        n10736), .ZN(n9445) );
  OAI221_X1 U11851 ( .B1(n12959), .B2(keyinput_g51), .C1(n10736), .C2(
        keyinput_g24), .A(n9445), .ZN(n9449) );
  AOI22_X1 U11852 ( .A1(n10724), .A2(keyinput_g21), .B1(n13705), .B2(
        keyinput_g5), .ZN(n9446) );
  OAI221_X1 U11853 ( .B1(n10724), .B2(keyinput_g21), .C1(n13705), .C2(
        keyinput_g5), .A(n9446), .ZN(n9448) );
  XNOR2_X1 U11854 ( .A(n9921), .B(keyinput_g123), .ZN(n9447) );
  OR3_X1 U11855 ( .A1(n9449), .A2(n9448), .A3(n9447), .ZN(n9453) );
  INV_X1 U11856 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n11522) );
  INV_X1 U11857 ( .A(P3_DATAO_REG_8__SCAN_IN), .ZN(n11456) );
  AOI22_X1 U11858 ( .A1(n11522), .A2(keyinput_g70), .B1(keyinput_g88), .B2(
        n11456), .ZN(n9450) );
  OAI221_X1 U11859 ( .B1(n11522), .B2(keyinput_g70), .C1(n11456), .C2(
        keyinput_g88), .A(n9450), .ZN(n9452) );
  XNOR2_X1 U11860 ( .A(n11008), .B(keyinput_g98), .ZN(n9451) );
  NOR3_X1 U11861 ( .A1(n9453), .A2(n9452), .A3(n9451), .ZN(n9463) );
  INV_X1 U11862 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n11241) );
  AOI22_X1 U11863 ( .A1(n11241), .A2(keyinput_g54), .B1(n9564), .B2(
        keyinput_g57), .ZN(n9454) );
  OAI221_X1 U11864 ( .B1(n11241), .B2(keyinput_g54), .C1(n9564), .C2(
        keyinput_g57), .A(n9454), .ZN(n9461) );
  INV_X1 U11865 ( .A(SI_7_), .ZN(n10732) );
  INV_X1 U11866 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n11365) );
  AOI22_X1 U11867 ( .A1(n10732), .A2(keyinput_g25), .B1(keyinput_g81), .B2(
        n11365), .ZN(n9455) );
  OAI221_X1 U11868 ( .B1(n10732), .B2(keyinput_g25), .C1(n11365), .C2(
        keyinput_g81), .A(n9455), .ZN(n9460) );
  INV_X1 U11869 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U11870 ( .A1(n11353), .A2(keyinput_g96), .B1(n12883), .B2(
        keyinput_g37), .ZN(n9456) );
  OAI221_X1 U11871 ( .B1(n11353), .B2(keyinput_g96), .C1(n12883), .C2(
        keyinput_g37), .A(n9456), .ZN(n9459) );
  INV_X1 U11872 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n12936) );
  INV_X1 U11873 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n11450) );
  AOI22_X1 U11874 ( .A1(n12936), .A2(keyinput_g48), .B1(keyinput_g84), .B2(
        n11450), .ZN(n9457) );
  OAI221_X1 U11875 ( .B1(n12936), .B2(keyinput_g48), .C1(n11450), .C2(
        keyinput_g84), .A(n9457), .ZN(n9458) );
  NOR4_X1 U11876 ( .A1(n9461), .A2(n9460), .A3(n9459), .A4(n9458), .ZN(n9462)
         );
  NAND4_X1 U11877 ( .A1(n9465), .A2(n9464), .A3(n9463), .A4(n9462), .ZN(n9466)
         );
  NOR4_X1 U11878 ( .A1(n9469), .A2(n9468), .A3(n9467), .A4(n9466), .ZN(n9642)
         );
  OAI22_X1 U11879 ( .A1(SI_23_), .A2(keyinput_f9), .B1(
        P3_DATAO_REG_15__SCAN_IN), .B2(keyinput_f81), .ZN(n9470) );
  AOI221_X1 U11880 ( .B1(SI_23_), .B2(keyinput_f9), .C1(keyinput_f81), .C2(
        P3_DATAO_REG_15__SCAN_IN), .A(n9470), .ZN(n9477) );
  OAI22_X1 U11881 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(keyinput_f61), .B1(
        keyinput_f1), .B2(SI_31_), .ZN(n9471) );
  AOI221_X1 U11882 ( .B1(P3_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .C1(
        SI_31_), .C2(keyinput_f1), .A(n9471), .ZN(n9476) );
  OAI22_X1 U11883 ( .A1(P3_REG3_REG_0__SCAN_IN), .A2(keyinput_f54), .B1(
        keyinput_f89), .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n9472) );
  AOI221_X1 U11884 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput_f54), .C1(
        P3_DATAO_REG_7__SCAN_IN), .C2(keyinput_f89), .A(n9472), .ZN(n9475) );
  OAI22_X1 U11885 ( .A1(SI_2_), .A2(keyinput_f30), .B1(
        P3_DATAO_REG_29__SCAN_IN), .B2(keyinput_f67), .ZN(n9473) );
  AOI221_X1 U11886 ( .B1(SI_2_), .B2(keyinput_f30), .C1(keyinput_f67), .C2(
        P3_DATAO_REG_29__SCAN_IN), .A(n9473), .ZN(n9474) );
  NAND4_X1 U11887 ( .A1(n9477), .A2(n9476), .A3(n9475), .A4(n9474), .ZN(n9600)
         );
  OAI22_X1 U11888 ( .A1(P3_B_REG_SCAN_IN), .A2(keyinput_f64), .B1(SI_9_), .B2(
        keyinput_f23), .ZN(n9478) );
  AOI221_X1 U11889 ( .B1(P3_B_REG_SCAN_IN), .B2(keyinput_f64), .C1(
        keyinput_f23), .C2(SI_9_), .A(n9478), .ZN(n9503) );
  OAI22_X1 U11890 ( .A1(SI_0_), .A2(keyinput_f32), .B1(P3_RD_REG_SCAN_IN), 
        .B2(keyinput_f33), .ZN(n9479) );
  AOI221_X1 U11891 ( .B1(SI_0_), .B2(keyinput_f32), .C1(keyinput_f33), .C2(
        P3_RD_REG_SCAN_IN), .A(n9479), .ZN(n9482) );
  OAI22_X1 U11892 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(keyinput_f123), .B1(
        P3_DATAO_REG_13__SCAN_IN), .B2(keyinput_f83), .ZN(n9480) );
  AOI221_X1 U11893 ( .B1(P1_IR_REG_16__SCAN_IN), .B2(keyinput_f123), .C1(
        keyinput_f83), .C2(P3_DATAO_REG_13__SCAN_IN), .A(n9480), .ZN(n9481) );
  OAI211_X1 U11894 ( .C1(n11183), .C2(keyinput_f14), .A(n9482), .B(n9481), 
        .ZN(n9483) );
  AOI21_X1 U11895 ( .B1(n11183), .B2(keyinput_f14), .A(n9483), .ZN(n9502) );
  AOI22_X1 U11896 ( .A1(SI_5_), .A2(keyinput_f27), .B1(P3_REG3_REG_13__SCAN_IN), .B2(keyinput_f56), .ZN(n9484) );
  OAI221_X1 U11897 ( .B1(SI_5_), .B2(keyinput_f27), .C1(
        P3_REG3_REG_13__SCAN_IN), .C2(keyinput_f56), .A(n9484), .ZN(n9491) );
  AOI22_X1 U11898 ( .A1(SI_20_), .A2(keyinput_f12), .B1(
        P3_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .ZN(n9485) );
  OAI221_X1 U11899 ( .B1(SI_20_), .B2(keyinput_f12), .C1(
        P3_REG3_REG_10__SCAN_IN), .C2(keyinput_f39), .A(n9485), .ZN(n9490) );
  AOI22_X1 U11900 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput_f110), .B1(
        P3_REG3_REG_4__SCAN_IN), .B2(keyinput_f52), .ZN(n9486) );
  OAI221_X1 U11901 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput_f110), .C1(
        P3_REG3_REG_4__SCAN_IN), .C2(keyinput_f52), .A(n9486), .ZN(n9489) );
  AOI22_X1 U11902 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(keyinput_f103), .B1(
        P3_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .ZN(n9487) );
  OAI221_X1 U11903 ( .B1(P3_ADDR_REG_6__SCAN_IN), .B2(keyinput_f103), .C1(
        P3_REG3_REG_26__SCAN_IN), .C2(keyinput_f62), .A(n9487), .ZN(n9488) );
  NOR4_X1 U11904 ( .A1(n9491), .A2(n9490), .A3(n9489), .A4(n9488), .ZN(n9501)
         );
  AOI22_X1 U11905 ( .A1(keyinput_f71), .A2(P3_DATAO_REG_25__SCAN_IN), .B1(
        SI_19_), .B2(keyinput_f13), .ZN(n9492) );
  OAI221_X1 U11906 ( .B1(keyinput_f71), .B2(P3_DATAO_REG_25__SCAN_IN), .C1(
        SI_19_), .C2(keyinput_f13), .A(n9492), .ZN(n9499) );
  AOI22_X1 U11907 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(keyinput_f111), .B1(
        P3_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .ZN(n9493) );
  OAI221_X1 U11908 ( .B1(P1_IR_REG_4__SCAN_IN), .B2(keyinput_f111), .C1(
        P3_REG3_REG_8__SCAN_IN), .C2(keyinput_f43), .A(n9493), .ZN(n9498) );
  AOI22_X1 U11909 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput_f116), .B1(SI_14_), 
        .B2(keyinput_f18), .ZN(n9494) );
  OAI221_X1 U11910 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput_f116), .C1(SI_14_), .C2(keyinput_f18), .A(n9494), .ZN(n9497) );
  AOI22_X1 U11911 ( .A1(keyinput_f75), .A2(P3_DATAO_REG_21__SCAN_IN), .B1(
        P3_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .ZN(n9495) );
  OAI221_X1 U11912 ( .B1(keyinput_f75), .B2(P3_DATAO_REG_21__SCAN_IN), .C1(
        P3_REG3_REG_21__SCAN_IN), .C2(keyinput_f45), .A(n9495), .ZN(n9496) );
  NOR4_X1 U11913 ( .A1(n9499), .A2(n9498), .A3(n9497), .A4(n9496), .ZN(n9500)
         );
  NAND4_X1 U11914 ( .A1(n9503), .A2(n9502), .A3(n9501), .A4(n9500), .ZN(n9599)
         );
  INV_X1 U11915 ( .A(SI_4_), .ZN(n10704) );
  AOI22_X1 U11916 ( .A1(n10736), .A2(keyinput_f24), .B1(keyinput_f28), .B2(
        n10704), .ZN(n9504) );
  OAI221_X1 U11917 ( .B1(n10736), .B2(keyinput_f24), .C1(n10704), .C2(
        keyinput_f28), .A(n9504), .ZN(n9513) );
  INV_X1 U11918 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9506) );
  AOI22_X1 U11919 ( .A1(n9506), .A2(keyinput_f126), .B1(n12883), .B2(
        keyinput_f37), .ZN(n9505) );
  OAI221_X1 U11920 ( .B1(n9506), .B2(keyinput_f126), .C1(n12883), .C2(
        keyinput_f37), .A(n9505), .ZN(n9512) );
  AOI22_X1 U11921 ( .A1(n10728), .A2(keyinput_f31), .B1(keyinput_f88), .B2(
        n11456), .ZN(n9507) );
  OAI221_X1 U11922 ( .B1(n10728), .B2(keyinput_f31), .C1(n11456), .C2(
        keyinput_f88), .A(n9507), .ZN(n9511) );
  INV_X1 U11923 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9509) );
  AOI22_X1 U11924 ( .A1(n9509), .A2(keyinput_f112), .B1(keyinput_f78), .B2(
        n11276), .ZN(n9508) );
  OAI221_X1 U11925 ( .B1(n9509), .B2(keyinput_f112), .C1(n11276), .C2(
        keyinput_f78), .A(n9508), .ZN(n9510) );
  NOR4_X1 U11926 ( .A1(n9513), .A2(n9512), .A3(n9511), .A4(n9510), .ZN(n9549)
         );
  INV_X1 U11927 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n11367) );
  AOI22_X1 U11928 ( .A1(n11367), .A2(keyinput_f82), .B1(n12944), .B2(
        keyinput_f50), .ZN(n9514) );
  OAI221_X1 U11929 ( .B1(n11367), .B2(keyinput_f82), .C1(n12944), .C2(
        keyinput_f50), .A(n9514), .ZN(n9523) );
  INV_X1 U11930 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n11355) );
  AOI22_X1 U11931 ( .A1(n11355), .A2(keyinput_f87), .B1(n13710), .B2(
        keyinput_f6), .ZN(n9515) );
  OAI221_X1 U11932 ( .B1(n11355), .B2(keyinput_f87), .C1(n13710), .C2(
        keyinput_f6), .A(n9515), .ZN(n9522) );
  AOI22_X1 U11933 ( .A1(n10732), .A2(keyinput_f25), .B1(n13705), .B2(
        keyinput_f5), .ZN(n9516) );
  OAI221_X1 U11934 ( .B1(n10732), .B2(keyinput_f25), .C1(n13705), .C2(
        keyinput_f5), .A(n9516), .ZN(n9521) );
  XOR2_X1 U11935 ( .A(n9517), .B(keyinput_f102), .Z(n9519) );
  XNOR2_X1 U11936 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_f107), .ZN(n9518) );
  NAND2_X1 U11937 ( .A1(n9519), .A2(n9518), .ZN(n9520) );
  NOR4_X1 U11938 ( .A1(n9523), .A2(n9522), .A3(n9521), .A4(n9520), .ZN(n9548)
         );
  AOI22_X1 U11939 ( .A1(n9525), .A2(keyinput_f47), .B1(n9878), .B2(
        keyinput_f36), .ZN(n9524) );
  OAI221_X1 U11940 ( .B1(n9525), .B2(keyinput_f47), .C1(n9878), .C2(
        keyinput_f36), .A(n9524), .ZN(n9533) );
  INV_X1 U11941 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9527) );
  AOI22_X1 U11942 ( .A1(n9527), .A2(keyinput_f115), .B1(keyinput_f91), .B2(
        n11361), .ZN(n9526) );
  OAI221_X1 U11943 ( .B1(n9527), .B2(keyinput_f115), .C1(n11361), .C2(
        keyinput_f91), .A(n9526), .ZN(n9532) );
  AOI22_X1 U11944 ( .A1(n11324), .A2(keyinput_f72), .B1(n10128), .B2(
        keyinput_f118), .ZN(n9528) );
  OAI221_X1 U11945 ( .B1(n11324), .B2(keyinput_f72), .C1(n10128), .C2(
        keyinput_f118), .A(n9528), .ZN(n9531) );
  AOI22_X1 U11946 ( .A1(n11450), .A2(keyinput_f84), .B1(n9211), .B2(
        keyinput_f100), .ZN(n9529) );
  OAI221_X1 U11947 ( .B1(n11450), .B2(keyinput_f84), .C1(n9211), .C2(
        keyinput_f100), .A(n9529), .ZN(n9530) );
  NOR4_X1 U11948 ( .A1(n9533), .A2(n9532), .A3(n9531), .A4(n9530), .ZN(n9547)
         );
  INV_X1 U11949 ( .A(keyinput_f0), .ZN(n9535) );
  AOI22_X1 U11950 ( .A1(n11359), .A2(keyinput_f79), .B1(P3_WR_REG_SCAN_IN), 
        .B2(n9535), .ZN(n9534) );
  OAI221_X1 U11951 ( .B1(n11359), .B2(keyinput_f79), .C1(n9535), .C2(
        P3_WR_REG_SCAN_IN), .A(n9534), .ZN(n9545) );
  INV_X1 U11952 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n9537) );
  AOI22_X1 U11953 ( .A1(n10983), .A2(keyinput_f77), .B1(n9537), .B2(
        keyinput_f55), .ZN(n9536) );
  OAI221_X1 U11954 ( .B1(n10983), .B2(keyinput_f77), .C1(n9537), .C2(
        keyinput_f55), .A(n9536), .ZN(n9544) );
  AOI22_X1 U11955 ( .A1(n13701), .A2(keyinput_f4), .B1(n12431), .B2(
        keyinput_f46), .ZN(n9538) );
  OAI221_X1 U11956 ( .B1(n13701), .B2(keyinput_f4), .C1(n12431), .C2(
        keyinput_f46), .A(n9538), .ZN(n9543) );
  XOR2_X1 U11957 ( .A(n9539), .B(keyinput_f117), .Z(n9541) );
  XNOR2_X1 U11958 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_f125), .ZN(n9540)
         );
  NAND2_X1 U11959 ( .A1(n9541), .A2(n9540), .ZN(n9542) );
  NOR4_X1 U11960 ( .A1(n9545), .A2(n9544), .A3(n9543), .A4(n9542), .ZN(n9546)
         );
  NAND4_X1 U11961 ( .A1(n9549), .A2(n9548), .A3(n9547), .A4(n9546), .ZN(n9598)
         );
  AOI22_X1 U11962 ( .A1(n11454), .A2(keyinput_f86), .B1(n12894), .B2(
        keyinput_f41), .ZN(n9550) );
  OAI221_X1 U11963 ( .B1(n11454), .B2(keyinput_f86), .C1(n12894), .C2(
        keyinput_f41), .A(n9550), .ZN(n9558) );
  AOI22_X1 U11964 ( .A1(n10720), .A2(keyinput_f22), .B1(n13025), .B2(
        keyinput_f63), .ZN(n9551) );
  OAI221_X1 U11965 ( .B1(n10720), .B2(keyinput_f22), .C1(n13025), .C2(
        keyinput_f63), .A(n9551), .ZN(n9557) );
  INV_X1 U11966 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n11823) );
  AOI22_X1 U11967 ( .A1(n11823), .A2(keyinput_f68), .B1(n9553), .B2(
        keyinput_f99), .ZN(n9552) );
  OAI221_X1 U11968 ( .B1(n11823), .B2(keyinput_f68), .C1(n9553), .C2(
        keyinput_f99), .A(n9552), .ZN(n9556) );
  INV_X1 U11969 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11014) );
  AOI22_X1 U11970 ( .A1(n12936), .A2(keyinput_f48), .B1(keyinput_f44), .B2(
        n11014), .ZN(n9554) );
  OAI221_X1 U11971 ( .B1(n12936), .B2(keyinput_f48), .C1(n11014), .C2(
        keyinput_f44), .A(n9554), .ZN(n9555) );
  NOR4_X1 U11972 ( .A1(n9558), .A2(n9557), .A3(n9556), .A4(n9555), .ZN(n9596)
         );
  INV_X1 U11973 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n9560) );
  AOI22_X1 U11974 ( .A1(n10864), .A2(keyinput_f17), .B1(n9560), .B2(
        keyinput_f42), .ZN(n9559) );
  OAI221_X1 U11975 ( .B1(n10864), .B2(keyinput_f17), .C1(n9560), .C2(
        keyinput_f42), .A(n9559), .ZN(n9571) );
  AOI22_X1 U11976 ( .A1(n9562), .A2(keyinput_f119), .B1(n12498), .B2(
        keyinput_f8), .ZN(n9561) );
  OAI221_X1 U11977 ( .B1(n9562), .B2(keyinput_f119), .C1(n12498), .C2(
        keyinput_f8), .A(n9561), .ZN(n9570) );
  AOI22_X1 U11978 ( .A1(n11789), .A2(keyinput_f11), .B1(n9564), .B2(
        keyinput_f57), .ZN(n9563) );
  OAI221_X1 U11979 ( .B1(n11789), .B2(keyinput_f11), .C1(n9564), .C2(
        keyinput_f57), .A(n9563), .ZN(n9569) );
  XOR2_X1 U11980 ( .A(n9565), .B(keyinput_f105), .Z(n9567) );
  XNOR2_X1 U11981 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_f113), .ZN(n9566) );
  NAND2_X1 U11982 ( .A1(n9567), .A2(n9566), .ZN(n9568) );
  NOR4_X1 U11983 ( .A1(n9571), .A2(n9570), .A3(n9569), .A4(n9568), .ZN(n9595)
         );
  AOI22_X1 U11984 ( .A1(n11740), .A2(keyinput_f40), .B1(keyinput_f93), .B2(
        n11399), .ZN(n9572) );
  OAI221_X1 U11985 ( .B1(n11740), .B2(keyinput_f40), .C1(n11399), .C2(
        keyinput_f93), .A(n9572), .ZN(n9580) );
  INV_X1 U11986 ( .A(SI_30_), .ZN(n13693) );
  AOI22_X1 U11987 ( .A1(n9574), .A2(keyinput_f97), .B1(n13693), .B2(
        keyinput_f2), .ZN(n9573) );
  OAI221_X1 U11988 ( .B1(n9574), .B2(keyinput_f97), .C1(n13693), .C2(
        keyinput_f2), .A(n9573), .ZN(n9579) );
  AOI22_X1 U11989 ( .A1(n11278), .A2(keyinput_f76), .B1(keyinput_f73), .B2(
        n11165), .ZN(n9575) );
  OAI221_X1 U11990 ( .B1(n11278), .B2(keyinput_f76), .C1(n11165), .C2(
        keyinput_f73), .A(n9575), .ZN(n9578) );
  INV_X1 U11991 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U11992 ( .A1(n11622), .A2(keyinput_f69), .B1(n7924), .B2(
        keyinput_f49), .ZN(n9576) );
  OAI221_X1 U11993 ( .B1(n11622), .B2(keyinput_f69), .C1(n7924), .C2(
        keyinput_f49), .A(n9576), .ZN(n9577) );
  NOR4_X1 U11994 ( .A1(n9580), .A2(n9579), .A3(n9578), .A4(n9577), .ZN(n9594)
         );
  INV_X1 U11995 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n11282) );
  AOI22_X1 U11996 ( .A1(n11282), .A2(keyinput_f94), .B1(n9582), .B2(
        keyinput_f106), .ZN(n9581) );
  OAI221_X1 U11997 ( .B1(n11282), .B2(keyinput_f94), .C1(n9582), .C2(
        keyinput_f106), .A(n9581), .ZN(n9592) );
  INV_X1 U11998 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9584) );
  AOI22_X1 U11999 ( .A1(n9584), .A2(keyinput_f121), .B1(keyinput_f98), .B2(
        n11008), .ZN(n9583) );
  OAI221_X1 U12000 ( .B1(n9584), .B2(keyinput_f121), .C1(n11008), .C2(
        keyinput_f98), .A(n9583), .ZN(n9591) );
  INV_X1 U12001 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U12002 ( .A1(n13002), .A2(keyinput_f60), .B1(keyinput_f80), .B2(
        n11357), .ZN(n9585) );
  OAI221_X1 U12003 ( .B1(n13002), .B2(keyinput_f60), .C1(n11357), .C2(
        keyinput_f80), .A(n9585), .ZN(n9590) );
  XOR2_X1 U12004 ( .A(n9586), .B(keyinput_f38), .Z(n9588) );
  XNOR2_X1 U12005 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_f127), .ZN(n9587)
         );
  NAND2_X1 U12006 ( .A1(n9588), .A2(n9587), .ZN(n9589) );
  NOR4_X1 U12007 ( .A1(n9592), .A2(n9591), .A3(n9590), .A4(n9589), .ZN(n9593)
         );
  NAND4_X1 U12008 ( .A1(n9596), .A2(n9595), .A3(n9594), .A4(n9593), .ZN(n9597)
         );
  NOR4_X1 U12009 ( .A1(n9600), .A2(n9599), .A3(n9598), .A4(n9597), .ZN(n9638)
         );
  OAI22_X1 U12010 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(keyinput_f53), .B1(
        keyinput_f101), .B2(P3_ADDR_REG_4__SCAN_IN), .ZN(n9601) );
  AOI221_X1 U12011 ( .B1(P3_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .C1(
        P3_ADDR_REG_4__SCAN_IN), .C2(keyinput_f101), .A(n9601), .ZN(n9608) );
  OAI22_X1 U12012 ( .A1(SI_25_), .A2(keyinput_f7), .B1(P3_DATAO_REG_6__SCAN_IN), .B2(keyinput_f90), .ZN(n9602) );
  AOI221_X1 U12013 ( .B1(SI_25_), .B2(keyinput_f7), .C1(keyinput_f90), .C2(
        P3_DATAO_REG_6__SCAN_IN), .A(n9602), .ZN(n9607) );
  OAI22_X1 U12014 ( .A1(P3_STATE_REG_SCAN_IN), .A2(keyinput_f34), .B1(
        keyinput_f58), .B2(P3_REG3_REG_11__SCAN_IN), .ZN(n9603) );
  AOI221_X1 U12015 ( .B1(P3_STATE_REG_SCAN_IN), .B2(keyinput_f34), .C1(
        P3_REG3_REG_11__SCAN_IN), .C2(keyinput_f58), .A(n9603), .ZN(n9606) );
  OAI22_X1 U12016 ( .A1(SI_29_), .A2(keyinput_f3), .B1(keyinput_f95), .B2(
        P3_DATAO_REG_1__SCAN_IN), .ZN(n9604) );
  AOI221_X1 U12017 ( .B1(SI_29_), .B2(keyinput_f3), .C1(
        P3_DATAO_REG_1__SCAN_IN), .C2(keyinput_f95), .A(n9604), .ZN(n9605) );
  NAND4_X1 U12018 ( .A1(n9608), .A2(n9607), .A3(n9606), .A4(n9605), .ZN(n9636)
         );
  OAI22_X1 U12019 ( .A1(SI_22_), .A2(keyinput_f10), .B1(SI_12_), .B2(
        keyinput_f20), .ZN(n9609) );
  AOI221_X1 U12020 ( .B1(SI_22_), .B2(keyinput_f10), .C1(keyinput_f20), .C2(
        SI_12_), .A(n9609), .ZN(n9616) );
  OAI22_X1 U12021 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput_f108), .B1(
        P3_DATAO_REG_0__SCAN_IN), .B2(keyinput_f96), .ZN(n9610) );
  AOI221_X1 U12022 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput_f108), .C1(
        keyinput_f96), .C2(P3_DATAO_REG_0__SCAN_IN), .A(n9610), .ZN(n9615) );
  OAI22_X1 U12023 ( .A1(P3_REG3_REG_2__SCAN_IN), .A2(keyinput_f59), .B1(
        keyinput_f70), .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n9611) );
  AOI221_X1 U12024 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(keyinput_f59), .C1(
        P3_DATAO_REG_26__SCAN_IN), .C2(keyinput_f70), .A(n9611), .ZN(n9614) );
  OAI22_X1 U12025 ( .A1(SI_16_), .A2(keyinput_f16), .B1(P1_IR_REG_13__SCAN_IN), 
        .B2(keyinput_f120), .ZN(n9612) );
  AOI221_X1 U12026 ( .B1(SI_16_), .B2(keyinput_f16), .C1(keyinput_f120), .C2(
        P1_IR_REG_13__SCAN_IN), .A(n9612), .ZN(n9613) );
  NAND4_X1 U12027 ( .A1(n9616), .A2(n9615), .A3(n9614), .A4(n9613), .ZN(n9635)
         );
  OAI22_X1 U12028 ( .A1(SI_13_), .A2(keyinput_f19), .B1(P1_IR_REG_2__SCAN_IN), 
        .B2(keyinput_f109), .ZN(n9617) );
  AOI221_X1 U12029 ( .B1(SI_13_), .B2(keyinput_f19), .C1(keyinput_f109), .C2(
        P1_IR_REG_2__SCAN_IN), .A(n9617), .ZN(n9624) );
  OAI22_X1 U12030 ( .A1(SI_11_), .A2(keyinput_f21), .B1(
        P3_DATAO_REG_22__SCAN_IN), .B2(keyinput_f74), .ZN(n9618) );
  AOI221_X1 U12031 ( .B1(SI_11_), .B2(keyinput_f21), .C1(keyinput_f74), .C2(
        P3_DATAO_REG_22__SCAN_IN), .A(n9618), .ZN(n9623) );
  OAI22_X1 U12032 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(keyinput_f51), .B1(
        keyinput_f104), .B2(P3_ADDR_REG_7__SCAN_IN), .ZN(n9619) );
  AOI221_X1 U12033 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .C1(
        P3_ADDR_REG_7__SCAN_IN), .C2(keyinput_f104), .A(n9619), .ZN(n9622) );
  OAI22_X1 U12034 ( .A1(SI_3_), .A2(keyinput_f29), .B1(keyinput_f122), .B2(
        P1_IR_REG_15__SCAN_IN), .ZN(n9620) );
  AOI221_X1 U12035 ( .B1(SI_3_), .B2(keyinput_f29), .C1(P1_IR_REG_15__SCAN_IN), 
        .C2(keyinput_f122), .A(n9620), .ZN(n9621) );
  NAND4_X1 U12036 ( .A1(n9624), .A2(n9623), .A3(n9622), .A4(n9621), .ZN(n9634)
         );
  OAI22_X1 U12037 ( .A1(SI_6_), .A2(keyinput_f26), .B1(keyinput_f114), .B2(
        P1_IR_REG_7__SCAN_IN), .ZN(n9625) );
  AOI221_X1 U12038 ( .B1(SI_6_), .B2(keyinput_f26), .C1(P1_IR_REG_7__SCAN_IN), 
        .C2(keyinput_f114), .A(n9625), .ZN(n9632) );
  OAI22_X1 U12039 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(keyinput_f35), .B1(SI_17_), .B2(keyinput_f15), .ZN(n9626) );
  AOI221_X1 U12040 ( .B1(P3_REG3_REG_7__SCAN_IN), .B2(keyinput_f35), .C1(
        keyinput_f15), .C2(SI_17_), .A(n9626), .ZN(n9631) );
  OAI22_X1 U12041 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput_f124), .B1(
        P3_DATAO_REG_11__SCAN_IN), .B2(keyinput_f85), .ZN(n9627) );
  AOI221_X1 U12042 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput_f124), .C1(
        keyinput_f85), .C2(P3_DATAO_REG_11__SCAN_IN), .A(n9627), .ZN(n9630) );
  OAI22_X1 U12043 ( .A1(n11728), .A2(keyinput_f66), .B1(keyinput_f65), .B2(
        P3_DATAO_REG_31__SCAN_IN), .ZN(n9628) );
  AOI221_X1 U12044 ( .B1(n11728), .B2(keyinput_f66), .C1(
        P3_DATAO_REG_31__SCAN_IN), .C2(keyinput_f65), .A(n9628), .ZN(n9629) );
  NAND4_X1 U12045 ( .A1(n9632), .A2(n9631), .A3(n9630), .A4(n9629), .ZN(n9633)
         );
  NOR4_X1 U12046 ( .A1(n9636), .A2(n9635), .A3(n9634), .A4(n9633), .ZN(n9637)
         );
  AOI22_X1 U12047 ( .A1(n9638), .A2(n9637), .B1(keyinput_f92), .B2(
        P3_DATAO_REG_4__SCAN_IN), .ZN(n9639) );
  OAI21_X1 U12048 ( .B1(keyinput_f92), .B2(P3_DATAO_REG_4__SCAN_IN), .A(n9639), 
        .ZN(n9640) );
  OAI21_X1 U12049 ( .B1(n11280), .B2(keyinput_g92), .A(n9640), .ZN(n9641) );
  AOI211_X1 U12050 ( .C1(n11280), .C2(keyinput_g92), .A(n9642), .B(n9641), 
        .ZN(n9643) );
  OR2_X1 U12051 ( .A1(n9686), .A2(n9178), .ZN(n9647) );
  OR2_X1 U12052 ( .A1(n13946), .A2(n11109), .ZN(n9648) );
  INV_X1 U12053 ( .A(n11568), .ZN(n9649) );
  NAND2_X1 U12054 ( .A1(n11559), .A2(n9649), .ZN(n9651) );
  INV_X1 U12055 ( .A(n13783), .ZN(n15708) );
  INV_X1 U12056 ( .A(n13945), .ZN(n11130) );
  NAND2_X1 U12057 ( .A1(n15708), .A2(n11130), .ZN(n9650) );
  NAND2_X1 U12058 ( .A1(n9651), .A2(n9650), .ZN(n11092) );
  INV_X1 U12059 ( .A(n11093), .ZN(n9652) );
  INV_X1 U12060 ( .A(n13944), .ZN(n9691) );
  NAND2_X1 U12061 ( .A1(n15662), .A2(n9691), .ZN(n9653) );
  NOR2_X1 U12062 ( .A1(n11590), .A2(n13943), .ZN(n9654) );
  NAND2_X1 U12063 ( .A1(n11590), .A2(n13943), .ZN(n9655) );
  NAND2_X1 U12064 ( .A1(n11395), .A2(n13942), .ZN(n9656) );
  NAND2_X1 U12065 ( .A1(n9657), .A2(n9656), .ZN(n11523) );
  NAND2_X1 U12066 ( .A1(n11534), .A2(n13941), .ZN(n9658) );
  INV_X1 U12067 ( .A(n11806), .ZN(n11809) );
  NAND2_X1 U12068 ( .A1(n11879), .A2(n13939), .ZN(n9660) );
  INV_X1 U12069 ( .A(n11859), .ZN(n11850) );
  NAND2_X1 U12070 ( .A1(n11860), .A2(n11850), .ZN(n9662) );
  NAND2_X1 U12071 ( .A1(n11991), .A2(n13938), .ZN(n9661) );
  AND2_X1 U12072 ( .A1(n12105), .A2(n13937), .ZN(n9664) );
  OR2_X1 U12073 ( .A1(n12105), .A2(n13937), .ZN(n9663) );
  OAI21_X2 U12074 ( .B1(n11893), .B2(n9664), .A(n9663), .ZN(n12043) );
  NAND2_X1 U12075 ( .A1(n15280), .A2(n13934), .ZN(n9665) );
  AND2_X2 U12076 ( .A1(n15265), .A2(n9665), .ZN(n12484) );
  OR2_X1 U12077 ( .A1(n12570), .A2(n13933), .ZN(n9667) );
  NAND2_X1 U12078 ( .A1(n14364), .A2(n13932), .ZN(n9668) );
  NAND2_X1 U12079 ( .A1(n14359), .A2(n13931), .ZN(n9669) );
  NOR2_X1 U12080 ( .A1(n14345), .A2(n13929), .ZN(n9670) );
  NAND2_X1 U12081 ( .A1(n14345), .A2(n13929), .ZN(n9671) );
  OR2_X1 U12082 ( .A1(n14341), .A2(n13928), .ZN(n9672) );
  INV_X1 U12083 ( .A(n14179), .ZN(n14181) );
  NOR2_X1 U12084 ( .A1(n14337), .A2(n13927), .ZN(n9673) );
  NAND2_X1 U12085 ( .A1(n14163), .A2(n14166), .ZN(n14165) );
  NAND2_X1 U12086 ( .A1(n14394), .A2(n13926), .ZN(n9675) );
  NAND2_X1 U12087 ( .A1(n14165), .A2(n9675), .ZN(n14145) );
  OR2_X1 U12088 ( .A1(n14159), .A2(n13925), .ZN(n9676) );
  NAND2_X1 U12089 ( .A1(n14316), .A2(n13924), .ZN(n9678) );
  OR2_X1 U12090 ( .A1(n14310), .A2(n13923), .ZN(n9679) );
  NOR2_X1 U12091 ( .A1(n14108), .A2(n13922), .ZN(n9680) );
  NAND2_X1 U12092 ( .A1(n14292), .A2(n13920), .ZN(n9681) );
  NAND2_X1 U12093 ( .A1(n9682), .A2(n9681), .ZN(n9683) );
  XNOR2_X1 U12094 ( .A(n9683), .B(n9737), .ZN(n14067) );
  INV_X1 U12095 ( .A(n14194), .ZN(n14197) );
  INV_X1 U12096 ( .A(n13929), .ZN(n9721) );
  NOR2_X1 U12097 ( .A1(n14345), .A2(n9721), .ZN(n9720) );
  OR2_X1 U12098 ( .A1(n9686), .A2(n15698), .ZN(n9687) );
  OR2_X1 U12099 ( .A1(n6915), .A2(n13946), .ZN(n9688) );
  NAND2_X1 U12100 ( .A1(n13783), .A2(n11130), .ZN(n9690) );
  NAND2_X1 U12101 ( .A1(n11125), .A2(n9691), .ZN(n9692) );
  NAND2_X1 U12102 ( .A1(n9693), .A2(n9692), .ZN(n11327) );
  NAND2_X1 U12103 ( .A1(n11327), .A2(n11328), .ZN(n9696) );
  INV_X1 U12104 ( .A(n13943), .ZN(n9694) );
  NAND2_X1 U12105 ( .A1(n11590), .A2(n9694), .ZN(n9695) );
  INV_X1 U12106 ( .A(n11388), .ZN(n11384) );
  NAND2_X1 U12107 ( .A1(n11389), .A2(n11384), .ZN(n9698) );
  NAND2_X1 U12108 ( .A1(n11395), .A2(n11488), .ZN(n9697) );
  NAND2_X1 U12109 ( .A1(n11534), .A2(n11746), .ZN(n9699) );
  NAND2_X1 U12110 ( .A1(n11754), .A2(n11759), .ZN(n9700) );
  INV_X1 U12111 ( .A(n13939), .ZN(n11851) );
  NAND2_X1 U12112 ( .A1(n11879), .A2(n11851), .ZN(n9701) );
  NAND2_X1 U12113 ( .A1(n11849), .A2(n11859), .ZN(n9703) );
  INV_X1 U12114 ( .A(n13938), .ZN(n11760) );
  NAND2_X1 U12115 ( .A1(n11991), .A2(n11760), .ZN(n9702) );
  NAND2_X1 U12116 ( .A1(n9703), .A2(n9702), .ZN(n11884) );
  NAND2_X1 U12117 ( .A1(n11884), .A2(n11892), .ZN(n9705) );
  INV_X1 U12118 ( .A(n13937), .ZN(n11852) );
  NAND2_X1 U12119 ( .A1(n12105), .A2(n11852), .ZN(n9704) );
  AND2_X1 U12120 ( .A1(n12191), .A2(n9707), .ZN(n9706) );
  OR2_X1 U12121 ( .A1(n12191), .A2(n9707), .ZN(n9708) );
  INV_X1 U12122 ( .A(n15280), .ZN(n9712) );
  NAND2_X1 U12123 ( .A1(n12570), .A2(n9713), .ZN(n9714) );
  INV_X1 U12124 ( .A(n13932), .ZN(n13845) );
  OR2_X1 U12125 ( .A1(n14364), .A2(n13845), .ZN(n9716) );
  AND2_X1 U12126 ( .A1(n14364), .A2(n13845), .ZN(n9715) );
  INV_X1 U12127 ( .A(n13931), .ZN(n9717) );
  OR2_X1 U12128 ( .A1(n14359), .A2(n9717), .ZN(n9718) );
  OR2_X1 U12129 ( .A1(n14353), .A2(n13840), .ZN(n9719) );
  NAND2_X1 U12130 ( .A1(n14345), .A2(n9721), .ZN(n14213) );
  NAND2_X1 U12131 ( .A1(n14197), .A2(n14198), .ZN(n14196) );
  NAND2_X1 U12132 ( .A1(n14341), .A2(n9722), .ZN(n9723) );
  INV_X1 U12133 ( .A(n13927), .ZN(n9725) );
  OR2_X1 U12134 ( .A1(n14337), .A2(n9725), .ZN(n9724) );
  NAND2_X1 U12135 ( .A1(n14337), .A2(n9725), .ZN(n9726) );
  INV_X1 U12136 ( .A(n13926), .ZN(n9727) );
  NAND2_X1 U12137 ( .A1(n14159), .A2(n13858), .ZN(n9728) );
  NAND2_X1 U12138 ( .A1(n14316), .A2(n9729), .ZN(n9730) );
  INV_X1 U12139 ( .A(n14117), .ZN(n14112) );
  NAND2_X1 U12140 ( .A1(n14310), .A2(n13856), .ZN(n9731) );
  INV_X1 U12141 ( .A(n13921), .ZN(n13810) );
  NAND2_X1 U12142 ( .A1(n14091), .A2(n13810), .ZN(n14073) );
  NAND2_X1 U12143 ( .A1(n9748), .A2(n10963), .ZN(n9740) );
  INV_X1 U12144 ( .A(n10767), .ZN(n10773) );
  NAND2_X1 U12145 ( .A1(n10773), .A2(P2_B_REG_SCAN_IN), .ZN(n9742) );
  AND2_X1 U12146 ( .A1(n13907), .A2(n9742), .ZN(n14053) );
  AOI22_X1 U12147 ( .A1(n14053), .A2(n13918), .B1(n13920), .B2(n13906), .ZN(
        n9743) );
  INV_X1 U12148 ( .A(n14359), .ZN(n14256) );
  INV_X1 U12149 ( .A(n12191), .ZN(n15289) );
  INV_X1 U12150 ( .A(n11991), .ZN(n11994) );
  INV_X1 U12151 ( .A(n11754), .ZN(n11865) );
  INV_X1 U12152 ( .A(n11395), .ZN(n11580) );
  NOR2_X1 U12153 ( .A1(n9178), .A2(n15691), .ZN(n11836) );
  NAND2_X1 U12154 ( .A1(n6915), .A2(n11836), .ZN(n11562) );
  INV_X1 U12155 ( .A(n11654), .ZN(n9745) );
  NAND2_X1 U12156 ( .A1(n11865), .A2(n9745), .ZN(n11808) );
  INV_X2 U12157 ( .A(n11856), .ZN(n11807) );
  OR2_X2 U12158 ( .A1(n15280), .A2(n15264), .ZN(n12490) );
  OR2_X2 U12159 ( .A1(n12570), .A2(n12490), .ZN(n14269) );
  INV_X1 U12160 ( .A(n14337), .ZN(n14191) );
  NAND2_X1 U12161 ( .A1(n14204), .A2(n14191), .ZN(n14186) );
  INV_X1 U12162 ( .A(n15263), .ZN(n14293) );
  OAI211_X1 U12163 ( .C1(n14291), .C2(n14077), .A(n14293), .B(n14049), .ZN(
        n14061) );
  NOR4_X1 U12164 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n9752) );
  NOR4_X1 U12165 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n9751) );
  NOR4_X1 U12166 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9750) );
  NOR4_X1 U12167 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n9749) );
  NAND4_X1 U12168 ( .A1(n9752), .A2(n9751), .A3(n9750), .A4(n9749), .ZN(n9761)
         );
  NOR2_X1 U12169 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n9756) );
  NOR4_X1 U12170 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9755) );
  NOR4_X1 U12171 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n9754) );
  NOR4_X1 U12172 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n9753) );
  NAND4_X1 U12173 ( .A1(n9756), .A2(n9755), .A3(n9754), .A4(n9753), .ZN(n9760)
         );
  INV_X1 U12174 ( .A(P2_B_REG_SCAN_IN), .ZN(n9757) );
  XOR2_X1 U12175 ( .A(n14431), .B(n9757), .Z(n9758) );
  OAI21_X1 U12176 ( .B1(n9761), .B2(n9760), .A(n15682), .ZN(n10952) );
  INV_X1 U12177 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15687) );
  NAND2_X1 U12178 ( .A1(n15682), .A2(n15687), .ZN(n9763) );
  NAND2_X1 U12179 ( .A1(n14424), .A2(n14427), .ZN(n9762) );
  NAND2_X1 U12180 ( .A1(n9763), .A2(n9762), .ZN(n15688) );
  AND2_X1 U12181 ( .A1(n10964), .A2(n15688), .ZN(n9764) );
  AND2_X1 U12182 ( .A1(n10952), .A2(n9764), .ZN(n10896) );
  NAND2_X1 U12183 ( .A1(n14431), .A2(n14424), .ZN(n9767) );
  INV_X1 U12184 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15684) );
  NAND2_X1 U12185 ( .A1(n15682), .A2(n15684), .ZN(n9766) );
  INV_X1 U12186 ( .A(n9768), .ZN(n9769) );
  NAND2_X1 U12187 ( .A1(n15685), .A2(n9769), .ZN(n9770) );
  OR2_X1 U12188 ( .A1(n15724), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9772) );
  NAND2_X1 U12189 ( .A1(n15724), .A2(n15281), .ZN(n14401) );
  NAND2_X1 U12190 ( .A1(n9775), .A2(n9774), .ZN(n9776) );
  NAND2_X1 U12191 ( .A1(n9777), .A2(n9776), .ZN(P2_U3496) );
  OAI21_X1 U12192 ( .B1(n13105), .B2(n13393), .A(n11663), .ZN(n9779) );
  XNOR2_X1 U12193 ( .A(n13224), .B(n12862), .ZN(n12869) );
  NOR2_X1 U12194 ( .A1(n12869), .A2(n12868), .ZN(n12864) );
  AOI21_X1 U12195 ( .B1(n12869), .B2(n12868), .A(n12864), .ZN(n9858) );
  XNOR2_X1 U12196 ( .A(n12951), .B(n9838), .ZN(n9780) );
  NAND2_X1 U12197 ( .A1(n9780), .A2(n13447), .ZN(n12923) );
  INV_X1 U12198 ( .A(n9780), .ZN(n9781) );
  NAND2_X1 U12199 ( .A1(n9781), .A2(n13483), .ZN(n9782) );
  INV_X1 U12200 ( .A(n11400), .ZN(n15790) );
  NAND2_X1 U12201 ( .A1(n11400), .A2(n9783), .ZN(n9785) );
  XNOR2_X1 U12202 ( .A(n6679), .B(n9789), .ZN(n9790) );
  XNOR2_X1 U12203 ( .A(n9790), .B(n15808), .ZN(n11496) );
  XNOR2_X1 U12204 ( .A(n6679), .B(n11547), .ZN(n9791) );
  XNOR2_X1 U12205 ( .A(n9791), .B(n11796), .ZN(n11737) );
  XNOR2_X1 U12206 ( .A(n9850), .B(n12109), .ZN(n9792) );
  XOR2_X1 U12207 ( .A(n11427), .B(n9792), .Z(n11794) );
  XNOR2_X1 U12208 ( .A(n9838), .B(n11979), .ZN(n9794) );
  XOR2_X1 U12209 ( .A(n11628), .B(n9794), .Z(n11974) );
  INV_X1 U12210 ( .A(n9794), .ZN(n9795) );
  INV_X1 U12211 ( .A(n11628), .ZN(n12027) );
  XNOR2_X1 U12212 ( .A(n9838), .B(n12030), .ZN(n9796) );
  XOR2_X1 U12213 ( .A(n11963), .B(n9796), .Z(n12025) );
  INV_X1 U12214 ( .A(n11963), .ZN(n12154) );
  XNOR2_X1 U12215 ( .A(n13134), .B(n12862), .ZN(n12152) );
  INV_X1 U12216 ( .A(n12152), .ZN(n9798) );
  NAND2_X1 U12217 ( .A1(n9798), .A2(n12286), .ZN(n9799) );
  XNOR2_X1 U12218 ( .A(n9838), .B(n15759), .ZN(n9800) );
  XOR2_X1 U12219 ( .A(n13143), .B(n9800), .Z(n12266) );
  NAND2_X1 U12220 ( .A1(n12267), .A2(n12266), .ZN(n12265) );
  NAND2_X1 U12221 ( .A1(n9800), .A2(n13143), .ZN(n9801) );
  XNOR2_X1 U12222 ( .A(n9838), .B(n13147), .ZN(n9802) );
  XNOR2_X1 U12223 ( .A(n9802), .B(n13148), .ZN(n12453) );
  INV_X1 U12224 ( .A(n9802), .ZN(n9804) );
  NAND2_X1 U12225 ( .A1(n9804), .A2(n9803), .ZN(n9805) );
  XNOR2_X1 U12226 ( .A(n9838), .B(n12520), .ZN(n9807) );
  XNOR2_X1 U12227 ( .A(n9807), .B(n15208), .ZN(n12515) );
  INV_X1 U12228 ( .A(n12515), .ZN(n9806) );
  NAND2_X1 U12229 ( .A1(n9807), .A2(n15208), .ZN(n9808) );
  XNOR2_X1 U12230 ( .A(n9838), .B(n15216), .ZN(n9809) );
  INV_X1 U12231 ( .A(n15198), .ZN(n12991) );
  NAND2_X1 U12232 ( .A1(n9810), .A2(n9809), .ZN(n12989) );
  XNOR2_X1 U12233 ( .A(n9838), .B(n9811), .ZN(n9812) );
  XNOR2_X1 U12234 ( .A(n9812), .B(n12994), .ZN(n12913) );
  NAND2_X1 U12235 ( .A1(n9812), .A2(n12994), .ZN(n9813) );
  XNOR2_X1 U12236 ( .A(n15194), .B(n9838), .ZN(n12973) );
  NOR2_X1 U12237 ( .A1(n12973), .A2(n15199), .ZN(n12877) );
  XNOR2_X1 U12238 ( .A(n13179), .B(n9838), .ZN(n9818) );
  XNOR2_X1 U12239 ( .A(n9818), .B(n15173), .ZN(n13019) );
  XNOR2_X1 U12240 ( .A(n15178), .B(n9838), .ZN(n9814) );
  NOR2_X1 U12241 ( .A1(n9814), .A2(n15187), .ZN(n13020) );
  OR2_X1 U12242 ( .A1(n12877), .A2(n6723), .ZN(n9817) );
  XNOR2_X1 U12243 ( .A(n9814), .B(n15187), .ZN(n12882) );
  INV_X1 U12244 ( .A(n12882), .ZN(n9815) );
  NAND2_X1 U12245 ( .A1(n12973), .A2(n15199), .ZN(n12878) );
  AND2_X1 U12246 ( .A1(n9815), .A2(n12878), .ZN(n12879) );
  OR2_X1 U12247 ( .A1(n6723), .A2(n12879), .ZN(n9816) );
  NAND2_X1 U12248 ( .A1(n9818), .A2(n15173), .ZN(n9819) );
  NAND2_X1 U12249 ( .A1(n13022), .A2(n9819), .ZN(n12934) );
  XNOR2_X1 U12250 ( .A(n13681), .B(n9838), .ZN(n9820) );
  NAND2_X1 U12251 ( .A1(n12934), .A2(n12935), .ZN(n9823) );
  INV_X1 U12252 ( .A(n9820), .ZN(n9821) );
  NAND2_X1 U12253 ( .A1(n9821), .A2(n13559), .ZN(n9822) );
  NAND2_X1 U12254 ( .A1(n9823), .A2(n9822), .ZN(n12942) );
  XNOR2_X1 U12255 ( .A(n13568), .B(n9838), .ZN(n9824) );
  XNOR2_X1 U12256 ( .A(n9824), .B(n13546), .ZN(n12943) );
  NAND2_X1 U12257 ( .A1(n12942), .A2(n12943), .ZN(n9826) );
  NAND2_X1 U12258 ( .A1(n9824), .A2(n13574), .ZN(n9825) );
  NAND2_X1 U12259 ( .A1(n9826), .A2(n9825), .ZN(n13000) );
  XNOR2_X1 U12260 ( .A(n13550), .B(n9838), .ZN(n9827) );
  NAND2_X1 U12261 ( .A1(n13000), .A2(n13001), .ZN(n9830) );
  INV_X1 U12262 ( .A(n9827), .ZN(n9828) );
  NAND2_X1 U12263 ( .A1(n9828), .A2(n13560), .ZN(n9829) );
  XNOR2_X1 U12264 ( .A(n13671), .B(n9838), .ZN(n9831) );
  XNOR2_X1 U12265 ( .A(n9831), .B(n13547), .ZN(n12893) );
  XNOR2_X1 U12266 ( .A(n13528), .B(n9838), .ZN(n9834) );
  XNOR2_X1 U12267 ( .A(n9834), .B(n13532), .ZN(n12965) );
  INV_X1 U12268 ( .A(n12965), .ZN(n9832) );
  NAND2_X1 U12269 ( .A1(n9831), .A2(n13547), .ZN(n12964) );
  AND2_X1 U12270 ( .A1(n9832), .A2(n12964), .ZN(n9833) );
  NAND2_X1 U12271 ( .A1(n9834), .A2(n13532), .ZN(n9835) );
  XNOR2_X1 U12272 ( .A(n13086), .B(n6679), .ZN(n9836) );
  XNOR2_X1 U12273 ( .A(n9836), .B(n13496), .ZN(n12904) );
  NAND2_X1 U12274 ( .A1(n9836), .A2(n13496), .ZN(n9837) );
  INV_X1 U12275 ( .A(n9842), .ZN(n9840) );
  XNOR2_X1 U12276 ( .A(n13499), .B(n9838), .ZN(n9841) );
  INV_X1 U12277 ( .A(n9841), .ZN(n9839) );
  NAND2_X1 U12278 ( .A1(n9842), .A2(n9841), .ZN(n9844) );
  XNOR2_X1 U12279 ( .A(n12713), .B(n9838), .ZN(n9845) );
  XNOR2_X1 U12280 ( .A(n12920), .B(n9838), .ZN(n9851) );
  NAND2_X1 U12281 ( .A1(n9851), .A2(n13433), .ZN(n9855) );
  INV_X1 U12282 ( .A(n9851), .ZN(n9852) );
  NAND2_X1 U12283 ( .A1(n9852), .A2(n13467), .ZN(n9853) );
  XNOR2_X1 U12284 ( .A(n13010), .B(n12862), .ZN(n9856) );
  NOR2_X1 U12285 ( .A1(n9856), .A2(n11520), .ZN(n9857) );
  AOI21_X1 U12286 ( .B1(n9856), .B2(n11520), .A(n9857), .ZN(n13012) );
  NAND2_X1 U12287 ( .A1(n9864), .A2(n15815), .ZN(n9859) );
  OAI22_X1 U12288 ( .A1(n9865), .A2(n9859), .B1(n9876), .B2(n9866), .ZN(n9861)
         );
  NAND2_X1 U12289 ( .A1(n9862), .A2(n13023), .ZN(n9886) );
  NAND2_X1 U12290 ( .A1(n9865), .A2(n15817), .ZN(n9863) );
  NAND2_X1 U12291 ( .A1(n9865), .A2(n9864), .ZN(n9870) );
  INV_X1 U12292 ( .A(n9866), .ZN(n9867) );
  NAND2_X1 U12293 ( .A1(n9876), .A2(n9867), .ZN(n9869) );
  NAND4_X1 U12294 ( .A1(n9870), .A2(n10588), .A3(n9869), .A4(n9868), .ZN(n9871) );
  NAND2_X1 U12295 ( .A1(n9871), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9873) );
  NOR2_X1 U12296 ( .A1(n10608), .A2(n11235), .ZN(n13241) );
  NAND2_X1 U12297 ( .A1(n9876), .A2(n13241), .ZN(n9872) );
  NAND2_X1 U12298 ( .A1(n9873), .A2(n9872), .ZN(n11267) );
  INV_X1 U12299 ( .A(n9874), .ZN(n10609) );
  NAND2_X1 U12300 ( .A1(n10609), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13245) );
  INV_X1 U12301 ( .A(n13245), .ZN(n9875) );
  INV_X1 U12302 ( .A(n9876), .ZN(n9877) );
  NAND2_X1 U12303 ( .A1(n9877), .A2(n13241), .ZN(n9879) );
  INV_X1 U12304 ( .A(n12321), .ZN(n12285) );
  OAI22_X1 U12305 ( .A1(n13448), .A2(n13028), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9878), .ZN(n9882) );
  NOR2_X1 U12306 ( .A1(n9880), .A2(n13016), .ZN(n9881) );
  AOI211_X1 U12307 ( .C1(n13423), .C2(n13031), .A(n9882), .B(n9881), .ZN(n9883) );
  NAND2_X1 U12308 ( .A1(n9886), .A2(n9885), .ZN(P3_U3154) );
  NOR2_X1 U12309 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), 
        .ZN(n9891) );
  NOR2_X1 U12310 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n9890) );
  NOR2_X1 U12311 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n9896) );
  NOR2_X1 U12312 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), 
        .ZN(n9895) );
  NOR2_X1 U12313 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), 
        .ZN(n9894) );
  NOR2_X1 U12314 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n9893) );
  XNOR2_X2 U12315 ( .A(n9900), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9906) );
  NAND2_X2 U12316 ( .A1(n9906), .A2(n9904), .ZN(n10404) );
  NAND2_X1 U12317 ( .A1(n10417), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9913) );
  INV_X2 U12318 ( .A(n9956), .ZN(n9971) );
  INV_X4 U12319 ( .A(n9971), .ZN(n10422) );
  INV_X1 U12320 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9905) );
  OR2_X1 U12321 ( .A1(n10422), .A2(n9905), .ZN(n9912) );
  NAND2_X1 U12322 ( .A1(n10055), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10071) );
  NAND2_X1 U12323 ( .A1(n10085), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10103) );
  NAND2_X1 U12324 ( .A1(n10153), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10178) );
  INV_X1 U12325 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n10177) );
  INV_X1 U12326 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n10192) );
  INV_X1 U12327 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n10245) );
  INV_X1 U12328 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n14459) );
  NAND2_X1 U12329 ( .A1(n10277), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n10278) );
  NAND2_X1 U12330 ( .A1(n10310), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n10309) );
  NAND2_X1 U12331 ( .A1(n10322), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n10321) );
  INV_X1 U12332 ( .A(n10321), .ZN(n10339) );
  NAND2_X1 U12333 ( .A1(n10339), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n10338) );
  INV_X1 U12334 ( .A(n10338), .ZN(n10348) );
  NAND2_X1 U12335 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n10348), .ZN(n10365) );
  INV_X1 U12336 ( .A(n10365), .ZN(n9907) );
  NAND2_X1 U12337 ( .A1(n9907), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n10378) );
  INV_X1 U12338 ( .A(n10378), .ZN(n9908) );
  NAND2_X1 U12339 ( .A1(n9908), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n14733) );
  OR2_X1 U12340 ( .A1(n10297), .A2(n14733), .ZN(n9911) );
  AND2_X2 U12341 ( .A1(n9904), .A2(n12706), .ZN(n10069) );
  INV_X1 U12342 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9909) );
  OR2_X1 U12343 ( .A1(n9970), .A2(n9909), .ZN(n9910) );
  NAND2_X1 U12344 ( .A1(n9914), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9916) );
  XNOR2_X2 U12345 ( .A(n9916), .B(n9915), .ZN(n10501) );
  NOR2_X1 U12346 ( .A1(n10424), .A2(n12861), .ZN(n9920) );
  NOR2_X2 U12347 ( .A1(n9923), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n9926) );
  NAND2_X1 U12348 ( .A1(n9923), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9924) );
  NAND2_X1 U12349 ( .A1(n10412), .A2(n14973), .ZN(n11439) );
  NAND2_X1 U12350 ( .A1(n11439), .A2(n9925), .ZN(n9928) );
  NAND2_X1 U12351 ( .A1(n9928), .A2(n12513), .ZN(n10429) );
  INV_X1 U12352 ( .A(n10397), .ZN(n10401) );
  NOR2_X1 U12353 ( .A1(n10717), .A2(n9388), .ZN(n9930) );
  XNOR2_X1 U12354 ( .A(n9930), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n15107) );
  INV_X1 U12355 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9932) );
  OR2_X1 U12356 ( .A1(n10404), .A2(n9932), .ZN(n9937) );
  INV_X1 U12357 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9933) );
  INV_X1 U12358 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10523) );
  OR2_X1 U12359 ( .A1(n9956), .A2(n10523), .ZN(n9935) );
  NAND2_X1 U12360 ( .A1(n10069), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9934) );
  OAI21_X1 U12361 ( .B1(n11506), .B2(n10509), .A(n14563), .ZN(n9939) );
  NAND2_X1 U12362 ( .A1(n11506), .A2(n10509), .ZN(n9938) );
  NAND2_X1 U12363 ( .A1(n9939), .A2(n9938), .ZN(n9940) );
  NAND2_X1 U12364 ( .A1(n9940), .A2(n9951), .ZN(n9950) );
  NAND2_X1 U12365 ( .A1(n11912), .A2(n10024), .ZN(n9949) );
  INV_X1 U12366 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n11827) );
  OR2_X1 U12367 ( .A1(n10404), .A2(n11827), .ZN(n9946) );
  INV_X1 U12368 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9941) );
  OR2_X1 U12369 ( .A1(n9956), .A2(n9941), .ZN(n9943) );
  NAND2_X1 U12370 ( .A1(n10069), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9942) );
  INV_X1 U12371 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n11613) );
  OR2_X1 U12372 ( .A1(n10380), .A2(n11613), .ZN(n9944) );
  INV_X1 U12373 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U12374 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9947) );
  XNOR2_X1 U12375 ( .A(n9948), .B(n9947), .ZN(n10920) );
  NAND2_X2 U12376 ( .A1(n9953), .A2(n11910), .ZN(n11919) );
  INV_X1 U12377 ( .A(n11910), .ZN(n9952) );
  INV_X1 U12378 ( .A(n9953), .ZN(n11911) );
  NAND2_X1 U12379 ( .A1(n11911), .A2(n10024), .ZN(n9954) );
  NAND2_X1 U12380 ( .A1(n9955), .A2(n9954), .ZN(n9967) );
  INV_X1 U12381 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10921) );
  OR2_X1 U12382 ( .A1(n9956), .A2(n10921), .ZN(n9958) );
  NAND2_X1 U12383 ( .A1(n10069), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9957) );
  INV_X1 U12384 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14576) );
  OR2_X1 U12385 ( .A1(n9960), .A2(n10013), .ZN(n9962) );
  XNOR2_X1 U12386 ( .A(n9962), .B(n9961), .ZN(n14584) );
  OR2_X1 U12387 ( .A1(n9963), .A2(n14584), .ZN(n9965) );
  INV_X1 U12388 ( .A(n10713), .ZN(n9964) );
  NAND2_X1 U12389 ( .A1(n10536), .A2(n15513), .ZN(n9986) );
  OAI21_X1 U12390 ( .B1(n9968), .B2(n9967), .A(n9966), .ZN(n9991) );
  INV_X1 U12391 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9969) );
  OR2_X1 U12392 ( .A1(n9970), .A2(n9969), .ZN(n9975) );
  OR2_X1 U12393 ( .A1(n6674), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9974) );
  NAND2_X1 U12394 ( .A1(n9971), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9973) );
  INV_X1 U12395 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10901) );
  OR2_X1 U12396 ( .A1(n10404), .A2(n10901), .ZN(n9972) );
  NAND4_X2 U12397 ( .A1(n9975), .A2(n9974), .A3(n9973), .A4(n9972), .ZN(n14561) );
  INV_X1 U12398 ( .A(n10715), .ZN(n9976) );
  OR2_X1 U12399 ( .A1(n9976), .A2(n10110), .ZN(n9984) );
  NAND2_X1 U12400 ( .A1(n9977), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9978) );
  MUX2_X1 U12401 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9978), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n9981) );
  NAND2_X1 U12402 ( .A1(n9981), .A2(n9980), .ZN(n14598) );
  OR2_X1 U12403 ( .A1(n9963), .A2(n14598), .ZN(n9983) );
  OR2_X1 U12404 ( .A1(n10424), .A2(n6986), .ZN(n9982) );
  AND3_X2 U12405 ( .A1(n9984), .A2(n9983), .A3(n9982), .ZN(n15518) );
  XNOR2_X1 U12406 ( .A(n14561), .B(n15518), .ZN(n12130) );
  INV_X1 U12407 ( .A(n12130), .ZN(n12137) );
  INV_X1 U12408 ( .A(n11913), .ZN(n9985) );
  NAND2_X1 U12409 ( .A1(n9985), .A2(n10024), .ZN(n9989) );
  INV_X1 U12410 ( .A(n9986), .ZN(n9987) );
  NAND3_X1 U12411 ( .A1(n9991), .A2(n12137), .A3(n9990), .ZN(n9995) );
  INV_X1 U12412 ( .A(n15518), .ZN(n12131) );
  NAND2_X1 U12413 ( .A1(n9951), .A2(n12131), .ZN(n9993) );
  NAND2_X1 U12414 ( .A1(n15518), .A2(n10024), .ZN(n9992) );
  MUX2_X1 U12415 ( .A(n9993), .B(n9992), .S(n14561), .Z(n9994) );
  NAND2_X1 U12416 ( .A1(n9995), .A2(n9994), .ZN(n10009) );
  OR2_X1 U12417 ( .A1(n9996), .A2(n10110), .ZN(n9999) );
  INV_X2 U12418 ( .A(n10424), .ZN(n10256) );
  INV_X2 U12419 ( .A(n9963), .ZN(n10781) );
  NAND2_X1 U12420 ( .A1(n9980), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9997) );
  XNOR2_X1 U12421 ( .A(n9997), .B(P1_IR_REG_4__SCAN_IN), .ZN(n15459) );
  AOI22_X1 U12422 ( .A1(n10256), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n10781), 
        .B2(n15459), .ZN(n9998) );
  NAND2_X1 U12423 ( .A1(n9999), .A2(n9998), .ZN(n14508) );
  NAND2_X1 U12424 ( .A1(n10417), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10005) );
  INV_X1 U12425 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10000) );
  OR2_X1 U12426 ( .A1(n10422), .A2(n10000), .ZN(n10004) );
  XNOR2_X1 U12427 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n14509) );
  OR2_X1 U12428 ( .A1(n6674), .A2(n14509), .ZN(n10003) );
  INV_X1 U12429 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10001) );
  OR2_X1 U12430 ( .A1(n9970), .A2(n10001), .ZN(n10002) );
  NAND4_X1 U12431 ( .A1(n10005), .A2(n10004), .A3(n10003), .A4(n10002), .ZN(
        n14560) );
  MUX2_X1 U12432 ( .A(n14508), .B(n14560), .S(n9951), .Z(n10006) );
  INV_X1 U12433 ( .A(n10006), .ZN(n10008) );
  MUX2_X1 U12434 ( .A(n14508), .B(n14560), .S(n10025), .Z(n10007) );
  OAI21_X1 U12435 ( .B1(n10009), .B2(n10008), .A(n10007), .ZN(n10011) );
  NAND2_X1 U12436 ( .A1(n10009), .A2(n10008), .ZN(n10010) );
  NAND2_X1 U12437 ( .A1(n10011), .A2(n10010), .ZN(n10028) );
  NAND2_X1 U12438 ( .A1(n10743), .A2(n10423), .ZN(n10016) );
  OR2_X1 U12439 ( .A1(n10012), .A2(n10013), .ZN(n10014) );
  XNOR2_X1 U12440 ( .A(n10014), .B(P1_IR_REG_5__SCAN_IN), .ZN(n14610) );
  AOI22_X1 U12441 ( .A1(n10256), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n10781), 
        .B2(n14610), .ZN(n10015) );
  NAND2_X1 U12442 ( .A1(n10016), .A2(n10015), .ZN(n11696) );
  INV_X1 U12443 ( .A(n6675), .ZN(n10280) );
  AOI21_X1 U12444 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10017) );
  NOR2_X1 U12445 ( .A1(n10017), .A2(n10038), .ZN(n11692) );
  NAND2_X1 U12446 ( .A1(n10280), .A2(n11692), .ZN(n10023) );
  INV_X1 U12447 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10907) );
  OR2_X1 U12448 ( .A1(n10404), .A2(n10907), .ZN(n10022) );
  INV_X1 U12449 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10018) );
  OR2_X1 U12450 ( .A1(n10422), .A2(n10018), .ZN(n10021) );
  INV_X1 U12451 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10019) );
  OR2_X1 U12452 ( .A1(n9970), .A2(n10019), .ZN(n10020) );
  NAND4_X1 U12453 ( .A1(n10023), .A2(n10022), .A3(n10021), .A4(n10020), .ZN(
        n14559) );
  MUX2_X1 U12454 ( .A(n11696), .B(n14559), .S(n10025), .Z(n10029) );
  NAND2_X1 U12455 ( .A1(n10028), .A2(n10029), .ZN(n10027) );
  MUX2_X1 U12456 ( .A(n11696), .B(n14559), .S(n9951), .Z(n10026) );
  NAND2_X1 U12457 ( .A1(n10027), .A2(n10026), .ZN(n10033) );
  INV_X1 U12458 ( .A(n10028), .ZN(n10031) );
  INV_X1 U12459 ( .A(n10029), .ZN(n10030) );
  NAND2_X1 U12460 ( .A1(n10031), .A2(n10030), .ZN(n10032) );
  OR2_X1 U12461 ( .A1(n10748), .A2(n10110), .ZN(n10036) );
  NAND2_X1 U12462 ( .A1(n10012), .A2(n9509), .ZN(n10051) );
  NAND2_X1 U12463 ( .A1(n10051), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10034) );
  XNOR2_X1 U12464 ( .A(n10034), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10923) );
  AOI22_X1 U12465 ( .A1(n10256), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n10781), 
        .B2(n10923), .ZN(n10035) );
  NAND2_X1 U12466 ( .A1(n10036), .A2(n10035), .ZN(n12055) );
  NAND2_X1 U12467 ( .A1(n10417), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10047) );
  INV_X1 U12468 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10037) );
  OR2_X1 U12469 ( .A1(n10422), .A2(n10037), .ZN(n10046) );
  INV_X1 U12470 ( .A(n10055), .ZN(n10042) );
  INV_X1 U12471 ( .A(n10038), .ZN(n10040) );
  INV_X1 U12472 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n10039) );
  NAND2_X1 U12473 ( .A1(n10040), .A2(n10039), .ZN(n10041) );
  NAND2_X1 U12474 ( .A1(n10042), .A2(n10041), .ZN(n12014) );
  OR2_X1 U12475 ( .A1(n10297), .A2(n12014), .ZN(n10045) );
  INV_X1 U12476 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10043) );
  OR2_X1 U12477 ( .A1(n9970), .A2(n10043), .ZN(n10044) );
  NAND4_X1 U12478 ( .A1(n10047), .A2(n10046), .A3(n10045), .A4(n10044), .ZN(
        n14558) );
  MUX2_X1 U12479 ( .A(n12055), .B(n14558), .S(n9951), .Z(n10049) );
  MUX2_X1 U12480 ( .A(n12055), .B(n14558), .S(n10025), .Z(n10048) );
  INV_X1 U12481 ( .A(n10049), .ZN(n10050) );
  OR2_X1 U12482 ( .A1(n10752), .A2(n10110), .ZN(n10054) );
  NAND2_X1 U12483 ( .A1(n10077), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10052) );
  XNOR2_X1 U12484 ( .A(n10052), .B(P1_IR_REG_7__SCAN_IN), .ZN(n14627) );
  AOI22_X1 U12485 ( .A1(n10256), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n10781), 
        .B2(n14627), .ZN(n10053) );
  NAND2_X1 U12486 ( .A1(n10054), .A2(n10053), .ZN(n12248) );
  NAND2_X1 U12487 ( .A1(n10417), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10060) );
  INV_X1 U12488 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10924) );
  OR2_X1 U12489 ( .A1(n10422), .A2(n10924), .ZN(n10059) );
  OAI21_X1 U12490 ( .B1(n10055), .B2(P1_REG3_REG_7__SCAN_IN), .A(n10071), .ZN(
        n12145) );
  OR2_X1 U12491 ( .A1(n6674), .A2(n12145), .ZN(n10058) );
  INV_X1 U12492 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10056) );
  OR2_X1 U12493 ( .A1(n9970), .A2(n10056), .ZN(n10057) );
  NAND4_X1 U12494 ( .A1(n10060), .A2(n10059), .A3(n10058), .A4(n10057), .ZN(
        n14557) );
  MUX2_X1 U12495 ( .A(n12248), .B(n14557), .S(n10025), .Z(n10064) );
  NAND2_X1 U12496 ( .A1(n10063), .A2(n10064), .ZN(n10062) );
  MUX2_X1 U12497 ( .A(n14557), .B(n12248), .S(n10025), .Z(n10061) );
  NAND2_X1 U12498 ( .A1(n10062), .A2(n10061), .ZN(n10068) );
  INV_X1 U12499 ( .A(n10063), .ZN(n10066) );
  INV_X1 U12500 ( .A(n10064), .ZN(n10065) );
  NAND2_X1 U12501 ( .A1(n10066), .A2(n10065), .ZN(n10067) );
  NAND2_X1 U12502 ( .A1(n10418), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10076) );
  INV_X1 U12503 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10926) );
  OR2_X1 U12504 ( .A1(n10422), .A2(n10926), .ZN(n10075) );
  AND2_X1 U12505 ( .A1(n10071), .A2(n10070), .ZN(n10072) );
  OR2_X1 U12506 ( .A1(n10072), .A2(n10085), .ZN(n12259) );
  OR2_X1 U12507 ( .A1(n10297), .A2(n12259), .ZN(n10074) );
  INV_X1 U12508 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10910) );
  OR2_X1 U12509 ( .A1(n10404), .A2(n10910), .ZN(n10073) );
  NAND4_X1 U12510 ( .A1(n10076), .A2(n10075), .A3(n10074), .A4(n10073), .ZN(
        n14556) );
  OR2_X1 U12511 ( .A1(n10793), .A2(n10110), .ZN(n10080) );
  NAND2_X1 U12512 ( .A1(n10187), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10078) );
  XNOR2_X1 U12513 ( .A(n10078), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U12514 ( .A1(n10256), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n10781), 
        .B2(n10942), .ZN(n10079) );
  MUX2_X1 U12515 ( .A(n14556), .B(n12302), .S(n10025), .Z(n10082) );
  MUX2_X1 U12516 ( .A(n12302), .B(n14556), .S(n10428), .Z(n10081) );
  INV_X1 U12517 ( .A(n10082), .ZN(n10083) );
  NAND2_X1 U12518 ( .A1(n10417), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10091) );
  INV_X1 U12519 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10084) );
  OR2_X1 U12520 ( .A1(n10422), .A2(n10084), .ZN(n10090) );
  OR2_X1 U12521 ( .A1(n10085), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10086) );
  NAND2_X1 U12522 ( .A1(n10103), .A2(n10086), .ZN(n12550) );
  OR2_X1 U12523 ( .A1(n10297), .A2(n12550), .ZN(n10089) );
  INV_X1 U12524 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10087) );
  OR2_X1 U12525 ( .A1(n9970), .A2(n10087), .ZN(n10088) );
  NAND4_X1 U12526 ( .A1(n10091), .A2(n10090), .A3(n10089), .A4(n10088), .ZN(
        n14555) );
  OR2_X1 U12527 ( .A1(n10853), .A2(n10110), .ZN(n10093) );
  XNOR2_X1 U12528 ( .A(n10160), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10993) );
  AOI22_X1 U12529 ( .A1(n10256), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n10781), 
        .B2(n10993), .ZN(n10092) );
  MUX2_X1 U12530 ( .A(n14555), .B(n12554), .S(n9951), .Z(n10097) );
  NAND2_X1 U12531 ( .A1(n10096), .A2(n10097), .ZN(n10095) );
  MUX2_X1 U12532 ( .A(n14555), .B(n12554), .S(n10428), .Z(n10094) );
  NAND2_X1 U12533 ( .A1(n10095), .A2(n10094), .ZN(n10101) );
  INV_X1 U12534 ( .A(n10096), .ZN(n10099) );
  INV_X1 U12535 ( .A(n10097), .ZN(n10098) );
  NAND2_X1 U12536 ( .A1(n10099), .A2(n10098), .ZN(n10100) );
  NAND2_X1 U12537 ( .A1(n10418), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n10109) );
  NAND2_X1 U12538 ( .A1(n10103), .A2(n10102), .ZN(n10104) );
  NAND2_X1 U12539 ( .A1(n10120), .A2(n10104), .ZN(n15321) );
  OR2_X1 U12540 ( .A1(n6675), .A2(n15321), .ZN(n10108) );
  INV_X1 U12541 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n12479) );
  OR2_X1 U12542 ( .A1(n10404), .A2(n12479), .ZN(n10107) );
  INV_X1 U12543 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10105) );
  OR2_X1 U12544 ( .A1(n10422), .A2(n10105), .ZN(n10106) );
  NAND4_X1 U12545 ( .A1(n10109), .A2(n10108), .A3(n10107), .A4(n10106), .ZN(
        n14554) );
  INV_X1 U12546 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n10111) );
  NAND2_X1 U12547 ( .A1(n10160), .A2(n10111), .ZN(n10112) );
  NAND2_X1 U12548 ( .A1(n10112), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10113) );
  XNOR2_X1 U12549 ( .A(n10113), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U12550 ( .A1(n10256), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n10781), 
        .B2(n10994), .ZN(n10114) );
  MUX2_X1 U12551 ( .A(n14554), .B(n15543), .S(n10428), .Z(n10117) );
  MUX2_X1 U12552 ( .A(n14554), .B(n15543), .S(n9951), .Z(n10116) );
  NAND2_X1 U12553 ( .A1(n10418), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n10125) );
  INV_X1 U12554 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10118) );
  OR2_X1 U12555 ( .A1(n10422), .A2(n10118), .ZN(n10124) );
  NAND2_X1 U12556 ( .A1(n10120), .A2(n10119), .ZN(n10121) );
  NAND2_X1 U12557 ( .A1(n10139), .A2(n10121), .ZN(n15354) );
  OR2_X1 U12558 ( .A1(n6674), .A2(n15354), .ZN(n10123) );
  INV_X1 U12559 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10989) );
  OR2_X1 U12560 ( .A1(n10404), .A2(n10989), .ZN(n10122) );
  NAND4_X1 U12561 ( .A1(n10125), .A2(n10124), .A3(n10123), .A4(n10122), .ZN(
        n14553) );
  NAND2_X1 U12562 ( .A1(n10978), .A2(n10423), .ZN(n10130) );
  OR2_X1 U12563 ( .A1(n10126), .A2(n10013), .ZN(n10127) );
  NAND2_X1 U12564 ( .A1(n10160), .A2(n10127), .ZN(n10145) );
  INV_X1 U12565 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n10128) );
  XNOR2_X1 U12566 ( .A(n10145), .B(n10128), .ZN(n14648) );
  AOI22_X1 U12567 ( .A1(n10256), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n10781), 
        .B2(n14648), .ZN(n10129) );
  MUX2_X1 U12568 ( .A(n14553), .B(n15403), .S(n9951), .Z(n10134) );
  NAND2_X1 U12569 ( .A1(n10133), .A2(n10134), .ZN(n10132) );
  MUX2_X1 U12570 ( .A(n14553), .B(n15403), .S(n10428), .Z(n10131) );
  NAND2_X1 U12571 ( .A1(n10132), .A2(n10131), .ZN(n10138) );
  INV_X1 U12572 ( .A(n10133), .ZN(n10136) );
  INV_X1 U12573 ( .A(n10134), .ZN(n10135) );
  NAND2_X1 U12574 ( .A1(n10136), .A2(n10135), .ZN(n10137) );
  NAND2_X1 U12575 ( .A1(n10418), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10144) );
  INV_X1 U12576 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n12538) );
  OR2_X1 U12577 ( .A1(n10404), .A2(n12538), .ZN(n10143) );
  INV_X1 U12578 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10996) );
  OR2_X1 U12579 ( .A1(n10422), .A2(n10996), .ZN(n10142) );
  AND2_X1 U12580 ( .A1(n10139), .A2(n12683), .ZN(n10140) );
  OR2_X1 U12581 ( .A1(n10140), .A2(n10153), .ZN(n12684) );
  OR2_X1 U12582 ( .A1(n10297), .A2(n12684), .ZN(n10141) );
  NAND4_X1 U12583 ( .A1(n10144), .A2(n10143), .A3(n10142), .A4(n10141), .ZN(
        n14552) );
  NAND2_X1 U12584 ( .A1(n11104), .A2(n10423), .ZN(n10148) );
  OAI21_X1 U12585 ( .B1(n10145), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10146) );
  XNOR2_X1 U12586 ( .A(n10146), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11000) );
  AOI22_X1 U12587 ( .A1(n10256), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n10781), 
        .B2(n11000), .ZN(n10147) );
  MUX2_X1 U12588 ( .A(n14552), .B(n12687), .S(n10428), .Z(n10150) );
  MUX2_X1 U12589 ( .A(n14552), .B(n12687), .S(n9951), .Z(n10149) );
  INV_X1 U12590 ( .A(n10150), .ZN(n10151) );
  NAND2_X1 U12591 ( .A1(n10418), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n10158) );
  INV_X1 U12592 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10152) );
  OR2_X1 U12593 ( .A1(n10422), .A2(n10152), .ZN(n10157) );
  OR2_X1 U12594 ( .A1(n10153), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10154) );
  NAND2_X1 U12595 ( .A1(n10178), .A2(n10154), .ZN(n15345) );
  OR2_X1 U12596 ( .A1(n6674), .A2(n15345), .ZN(n10156) );
  INV_X1 U12597 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11084) );
  OR2_X1 U12598 ( .A1(n10404), .A2(n11084), .ZN(n10155) );
  NAND4_X1 U12599 ( .A1(n10158), .A2(n10157), .A3(n10156), .A4(n10155), .ZN(
        n14551) );
  NAND2_X1 U12600 ( .A1(n11256), .A2(n10423), .ZN(n10163) );
  NAND2_X1 U12601 ( .A1(n10185), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10159) );
  NAND2_X1 U12602 ( .A1(n10160), .A2(n10159), .ZN(n10172) );
  XNOR2_X1 U12603 ( .A(n10172), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11257) );
  INV_X1 U12604 ( .A(n11257), .ZN(n10161) );
  AOI22_X1 U12605 ( .A1(n10256), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n10781), 
        .B2(n10161), .ZN(n10162) );
  MUX2_X1 U12606 ( .A(n14551), .B(n15342), .S(n9951), .Z(n10167) );
  NAND2_X1 U12607 ( .A1(n10166), .A2(n10167), .ZN(n10165) );
  MUX2_X1 U12608 ( .A(n14551), .B(n15342), .S(n10428), .Z(n10164) );
  NAND2_X1 U12609 ( .A1(n10165), .A2(n10164), .ZN(n10171) );
  INV_X1 U12610 ( .A(n10166), .ZN(n10169) );
  NAND2_X1 U12611 ( .A1(n10169), .A2(n10168), .ZN(n10170) );
  NAND2_X1 U12612 ( .A1(n10171), .A2(n10170), .ZN(n10204) );
  NAND2_X1 U12613 ( .A1(n11608), .A2(n10423), .ZN(n10175) );
  OAI21_X1 U12614 ( .B1(n10172), .B2(P1_IR_REG_13__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10173) );
  XNOR2_X1 U12615 ( .A(n10173), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11195) );
  AOI22_X1 U12616 ( .A1(n10256), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n10781), 
        .B2(n11195), .ZN(n10174) );
  NAND2_X1 U12617 ( .A1(n10418), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n10183) );
  INV_X1 U12618 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10176) );
  OR2_X1 U12619 ( .A1(n10422), .A2(n10176), .ZN(n10182) );
  NAND2_X1 U12620 ( .A1(n10178), .A2(n10177), .ZN(n10179) );
  NAND2_X1 U12621 ( .A1(n10193), .A2(n10179), .ZN(n15311) );
  OR2_X1 U12622 ( .A1(n6675), .A2(n15311), .ZN(n10181) );
  INV_X1 U12623 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n12613) );
  OR2_X1 U12624 ( .A1(n10404), .A2(n12613), .ZN(n10180) );
  NAND2_X1 U12625 ( .A1(n15386), .A2(n15362), .ZN(n10200) );
  NAND2_X1 U12626 ( .A1(n11803), .A2(n10423), .ZN(n10190) );
  NAND3_X1 U12627 ( .A1(n9397), .A2(n9527), .A3(n9584), .ZN(n10184) );
  OR2_X1 U12628 ( .A1(n10185), .A2(n10184), .ZN(n10186) );
  OAI21_X1 U12629 ( .B1(n10187), .B2(n10186), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n10188) );
  XNOR2_X1 U12630 ( .A(n10188), .B(P1_IR_REG_15__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U12631 ( .A1(n10256), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n10781), 
        .B2(n12218), .ZN(n10189) );
  NAND2_X1 U12632 ( .A1(n10418), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n10199) );
  INV_X1 U12633 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10191) );
  OR2_X1 U12634 ( .A1(n10422), .A2(n10191), .ZN(n10198) );
  AND2_X1 U12635 ( .A1(n10193), .A2(n10192), .ZN(n10194) );
  OR2_X1 U12636 ( .A1(n10194), .A2(n10220), .ZN(n15368) );
  OR2_X1 U12637 ( .A1(n6675), .A2(n15368), .ZN(n10197) );
  INV_X1 U12638 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10195) );
  OR2_X1 U12639 ( .A1(n10404), .A2(n10195), .ZN(n10196) );
  NAND2_X1 U12640 ( .A1(n14741), .A2(n12693), .ZN(n10202) );
  NAND2_X1 U12641 ( .A1(n14700), .A2(n15326), .ZN(n10464) );
  NAND2_X1 U12642 ( .A1(n10464), .A2(n10200), .ZN(n10201) );
  MUX2_X1 U12643 ( .A(n10202), .B(n10201), .S(n10428), .Z(n10203) );
  AOI21_X1 U12644 ( .B1(n10204), .B2(n12623), .A(n10203), .ZN(n10232) );
  INV_X1 U12645 ( .A(n10464), .ZN(n10205) );
  MUX2_X1 U12646 ( .A(n10205), .B(n7689), .S(n10428), .Z(n10231) );
  NAND2_X1 U12647 ( .A1(n12036), .A2(n10423), .ZN(n10210) );
  NAND2_X1 U12648 ( .A1(n10206), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10207) );
  XNOR2_X1 U12649 ( .A(n10207), .B(n7261), .ZN(n12503) );
  INV_X1 U12650 ( .A(n12503), .ZN(n10208) );
  AOI22_X1 U12651 ( .A1(n10256), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n10781), 
        .B2(n10208), .ZN(n10209) );
  NAND2_X1 U12652 ( .A1(n10418), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n10215) );
  INV_X1 U12653 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n12205) );
  OR2_X1 U12654 ( .A1(n10404), .A2(n12205), .ZN(n10214) );
  INV_X1 U12655 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n12504) );
  OR2_X1 U12656 ( .A1(n10422), .A2(n12504), .ZN(n10213) );
  OR2_X1 U12657 ( .A1(n10222), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10211) );
  NAND2_X1 U12658 ( .A1(n10246), .A2(n10211), .ZN(n14953) );
  OR2_X1 U12659 ( .A1(n6674), .A2(n14953), .ZN(n10212) );
  XNOR2_X1 U12660 ( .A(n15064), .B(n15325), .ZN(n10463) );
  NAND2_X1 U12661 ( .A1(n11972), .A2(n10423), .ZN(n10219) );
  OR2_X1 U12662 ( .A1(n10216), .A2(n10013), .ZN(n10217) );
  XNOR2_X1 U12663 ( .A(n10217), .B(P1_IR_REG_16__SCAN_IN), .ZN(n14661) );
  AOI22_X1 U12664 ( .A1(n10256), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n10781), 
        .B2(n14661), .ZN(n10218) );
  INV_X1 U12665 ( .A(n15371), .ZN(n15324) );
  NAND2_X1 U12666 ( .A1(n10418), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n10227) );
  INV_X1 U12667 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n12214) );
  OR2_X1 U12668 ( .A1(n10422), .A2(n12214), .ZN(n10226) );
  NOR2_X1 U12669 ( .A1(n10220), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10221) );
  OR2_X1 U12670 ( .A1(n10222), .A2(n10221), .ZN(n15332) );
  OR2_X1 U12671 ( .A1(n10297), .A2(n15332), .ZN(n10225) );
  INV_X1 U12672 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10223) );
  OR2_X1 U12673 ( .A1(n10404), .A2(n10223), .ZN(n10224) );
  NAND4_X1 U12674 ( .A1(n10227), .A2(n10226), .A3(n10225), .A4(n10224), .ZN(
        n14703) );
  INV_X1 U12675 ( .A(n14703), .ZN(n15359) );
  MUX2_X1 U12676 ( .A(n15324), .B(n15359), .S(n10428), .Z(n10234) );
  OR2_X1 U12677 ( .A1(n15064), .A2(n15325), .ZN(n14744) );
  NAND2_X1 U12678 ( .A1(n15064), .A2(n15325), .ZN(n14743) );
  AND2_X1 U12679 ( .A1(n14703), .A2(n9951), .ZN(n10228) );
  AOI21_X1 U12680 ( .B1(n15371), .B2(n10428), .A(n10228), .ZN(n10229) );
  NAND3_X1 U12681 ( .A1(n14744), .A2(n14743), .A3(n10229), .ZN(n10233) );
  OAI21_X1 U12682 ( .B1(n10463), .B2(n10234), .A(n10233), .ZN(n10230) );
  INV_X1 U12683 ( .A(n10233), .ZN(n10239) );
  INV_X1 U12684 ( .A(n10234), .ZN(n10238) );
  OAI21_X1 U12685 ( .B1(n14705), .B2(n10428), .A(n15064), .ZN(n10237) );
  INV_X1 U12686 ( .A(n15064), .ZN(n10235) );
  OAI21_X1 U12687 ( .B1(n15325), .B2(n9951), .A(n10235), .ZN(n10236) );
  AOI22_X1 U12688 ( .A1(n10239), .A2(n10238), .B1(n10237), .B2(n10236), .ZN(
        n10240) );
  NAND2_X1 U12689 ( .A1(n12295), .A2(n10423), .ZN(n10244) );
  NAND2_X1 U12690 ( .A1(n6828), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10242) );
  XNOR2_X1 U12691 ( .A(n10242), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14674) );
  AOI22_X1 U12692 ( .A1(n10256), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n10781), 
        .B2(n14674), .ZN(n10243) );
  NAND2_X1 U12693 ( .A1(n10246), .A2(n10245), .ZN(n10247) );
  AND2_X1 U12694 ( .A1(n10259), .A2(n10247), .ZN(n14942) );
  NAND2_X1 U12695 ( .A1(n10280), .A2(n14942), .ZN(n10254) );
  INV_X1 U12696 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10248) );
  OR2_X1 U12697 ( .A1(n10422), .A2(n10248), .ZN(n10253) );
  INV_X1 U12698 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10249) );
  OR2_X1 U12699 ( .A1(n10404), .A2(n10249), .ZN(n10252) );
  INV_X1 U12700 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10250) );
  OR2_X1 U12701 ( .A1(n9970), .A2(n10250), .ZN(n10251) );
  INV_X1 U12702 ( .A(n14489), .ZN(n14746) );
  OR2_X1 U12703 ( .A1(n15057), .A2(n14746), .ZN(n14707) );
  MUX2_X1 U12704 ( .A(n14489), .B(n14944), .S(n10428), .Z(n10255) );
  AND2_X1 U12705 ( .A1(n15057), .A2(n14746), .ZN(n14708) );
  NAND2_X1 U12706 ( .A1(n12387), .A2(n10423), .ZN(n10258) );
  AOI22_X1 U12707 ( .A1(n10256), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14814), 
        .B2(n10781), .ZN(n10257) );
  AND2_X1 U12708 ( .A1(n10259), .A2(n14459), .ZN(n10260) );
  OR2_X1 U12709 ( .A1(n10260), .A2(n10266), .ZN(n14921) );
  AOI22_X1 U12710 ( .A1(n9971), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n10417), 
        .B2(P1_REG2_REG_19__SCAN_IN), .ZN(n10262) );
  NAND2_X1 U12711 ( .A1(n10418), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n10261) );
  OAI211_X1 U12712 ( .C1(n14921), .C2(n6675), .A(n10262), .B(n10261), .ZN(
        n14709) );
  INV_X1 U12713 ( .A(n14709), .ZN(n10263) );
  OR2_X1 U12714 ( .A1(n15052), .A2(n10263), .ZN(n10264) );
  NAND2_X1 U12715 ( .A1(n15052), .A2(n10263), .ZN(n14749) );
  MUX2_X1 U12716 ( .A(n14749), .B(n10264), .S(n9951), .Z(n10265) );
  NOR2_X1 U12717 ( .A1(n10266), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n10267) );
  OR2_X1 U12718 ( .A1(n10277), .A2(n10267), .ZN(n14908) );
  AOI22_X1 U12719 ( .A1(n9971), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n10417), 
        .B2(P1_REG2_REG_20__SCAN_IN), .ZN(n10269) );
  NAND2_X1 U12720 ( .A1(n10418), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n10268) );
  OAI211_X1 U12721 ( .C1(n14908), .C2(n10297), .A(n10269), .B(n10268), .ZN(
        n14750) );
  NAND2_X1 U12722 ( .A1(n12391), .A2(n10423), .ZN(n10271) );
  OR2_X1 U12723 ( .A1(n10424), .A2(n12392), .ZN(n10270) );
  MUX2_X1 U12724 ( .A(n14710), .B(n14911), .S(n9951), .Z(n10273) );
  MUX2_X1 U12725 ( .A(n14750), .B(n15046), .S(n10428), .Z(n10272) );
  OAI21_X1 U12726 ( .B1(n10274), .B2(n10273), .A(n10272), .ZN(n10288) );
  NAND2_X1 U12727 ( .A1(n10274), .A2(n10273), .ZN(n10287) );
  NAND2_X1 U12728 ( .A1(n12463), .A2(n10423), .ZN(n10276) );
  OR2_X1 U12729 ( .A1(n10424), .A2(n12511), .ZN(n10275) );
  NAND2_X2 U12730 ( .A1(n10276), .A2(n10275), .ZN(n15041) );
  OR2_X1 U12731 ( .A1(n10277), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n10279) );
  AND2_X1 U12732 ( .A1(n10279), .A2(n10278), .ZN(n14895) );
  NAND2_X1 U12733 ( .A1(n14895), .A2(n10280), .ZN(n10286) );
  INV_X1 U12734 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10283) );
  NAND2_X1 U12735 ( .A1(n10417), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n10282) );
  NAND2_X1 U12736 ( .A1(n10418), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n10281) );
  OAI211_X1 U12737 ( .C1(n10422), .C2(n10283), .A(n10282), .B(n10281), .ZN(
        n10284) );
  INV_X1 U12738 ( .A(n10284), .ZN(n10285) );
  NAND2_X1 U12739 ( .A1(n10286), .A2(n10285), .ZN(n14712) );
  NAND3_X1 U12740 ( .A1(n10288), .A2(n10287), .A3(n14891), .ZN(n10292) );
  AND2_X1 U12741 ( .A1(n14712), .A2(n10428), .ZN(n10290) );
  OAI21_X1 U12742 ( .B1(n14712), .B2(n10428), .A(n15041), .ZN(n10289) );
  OAI21_X1 U12743 ( .B1(n10290), .B2(n15041), .A(n10289), .ZN(n10291) );
  NAND2_X1 U12744 ( .A1(n10292), .A2(n10291), .ZN(n10306) );
  OR2_X1 U12745 ( .A1(n8976), .A2(n10717), .ZN(n10293) );
  XNOR2_X1 U12746 ( .A(n10293), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15106) );
  NAND2_X1 U12747 ( .A1(n10417), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n10302) );
  INV_X1 U12748 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10294) );
  OR2_X1 U12749 ( .A1(n10422), .A2(n10294), .ZN(n10301) );
  OAI21_X1 U12750 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n10296), .A(n10295), 
        .ZN(n14880) );
  OR2_X1 U12751 ( .A1(n10297), .A2(n14880), .ZN(n10300) );
  INV_X1 U12752 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10298) );
  OR2_X1 U12753 ( .A1(n9970), .A2(n10298), .ZN(n10299) );
  MUX2_X1 U12754 ( .A(n14884), .B(n14714), .S(n10428), .Z(n10303) );
  INV_X1 U12755 ( .A(n10303), .ZN(n10305) );
  MUX2_X1 U12756 ( .A(n14714), .B(n14884), .S(n10428), .Z(n10304) );
  AOI21_X1 U12757 ( .B1(n10306), .B2(n10305), .A(n10304), .ZN(n10307) );
  NAND2_X1 U12758 ( .A1(n10417), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n10315) );
  INV_X1 U12759 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10308) );
  OR2_X1 U12760 ( .A1(n10422), .A2(n10308), .ZN(n10314) );
  OAI21_X1 U12761 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n10310), .A(n10309), 
        .ZN(n14866) );
  OR2_X1 U12762 ( .A1(n6674), .A2(n14866), .ZN(n10313) );
  INV_X1 U12763 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10311) );
  OR2_X1 U12764 ( .A1(n9970), .A2(n10311), .ZN(n10312) );
  NAND4_X1 U12765 ( .A1(n10315), .A2(n10314), .A3(n10313), .A4(n10312), .ZN(
        n14717) );
  NAND2_X1 U12766 ( .A1(n12629), .A2(n10423), .ZN(n10317) );
  OR2_X1 U12767 ( .A1(n10424), .A2(n12632), .ZN(n10316) );
  MUX2_X1 U12768 ( .A(n14717), .B(n15024), .S(n10428), .Z(n10319) );
  MUX2_X1 U12769 ( .A(n14717), .B(n15024), .S(n9951), .Z(n10318) );
  NAND2_X1 U12770 ( .A1(n9971), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n10326) );
  INV_X1 U12771 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10320) );
  OR2_X1 U12772 ( .A1(n9970), .A2(n10320), .ZN(n10325) );
  OAI21_X1 U12773 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n10322), .A(n10321), 
        .ZN(n14854) );
  OR2_X1 U12774 ( .A1(n6675), .A2(n14854), .ZN(n10324) );
  INV_X1 U12775 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n14855) );
  OR2_X1 U12776 ( .A1(n10404), .A2(n14855), .ZN(n10323) );
  NAND4_X1 U12777 ( .A1(n10326), .A2(n10325), .A3(n10324), .A4(n10323), .ZN(
        n14826) );
  NAND2_X1 U12778 ( .A1(n14430), .A2(n10423), .ZN(n10328) );
  OR2_X1 U12779 ( .A1(n10424), .A2(n15102), .ZN(n10327) );
  MUX2_X1 U12780 ( .A(n14826), .B(n14859), .S(n9951), .Z(n10332) );
  NAND2_X1 U12781 ( .A1(n10331), .A2(n10332), .ZN(n10330) );
  MUX2_X1 U12782 ( .A(n14826), .B(n14859), .S(n10428), .Z(n10329) );
  NAND2_X1 U12783 ( .A1(n10330), .A2(n10329), .ZN(n10336) );
  INV_X1 U12784 ( .A(n10331), .ZN(n10334) );
  INV_X1 U12785 ( .A(n10332), .ZN(n10333) );
  NAND2_X1 U12786 ( .A1(n10334), .A2(n10333), .ZN(n10335) );
  NAND2_X1 U12787 ( .A1(n9971), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n10343) );
  INV_X1 U12788 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10337) );
  OR2_X1 U12789 ( .A1(n9970), .A2(n10337), .ZN(n10342) );
  OAI21_X1 U12790 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n10339), .A(n10338), 
        .ZN(n14833) );
  OR2_X1 U12791 ( .A1(n10297), .A2(n14833), .ZN(n10341) );
  INV_X1 U12792 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n14834) );
  OR2_X1 U12793 ( .A1(n10404), .A2(n14834), .ZN(n10340) );
  NAND4_X1 U12794 ( .A1(n10343), .A2(n10342), .A3(n10341), .A4(n10340), .ZN(
        n14720) );
  NAND2_X1 U12795 ( .A1(n14426), .A2(n10423), .ZN(n10345) );
  OR2_X1 U12796 ( .A1(n10424), .A2(n15098), .ZN(n10344) );
  MUX2_X1 U12797 ( .A(n14720), .B(n15014), .S(n10428), .Z(n10347) );
  MUX2_X1 U12798 ( .A(n15014), .B(n14720), .S(n10428), .Z(n10346) );
  NAND2_X1 U12799 ( .A1(n9971), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n10353) );
  INV_X1 U12800 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n14816) );
  OR2_X1 U12801 ( .A1(n10404), .A2(n14816), .ZN(n10352) );
  OAI21_X1 U12802 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n10348), .A(n10365), 
        .ZN(n14815) );
  OR2_X1 U12803 ( .A1(n6674), .A2(n14815), .ZN(n10351) );
  INV_X1 U12804 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10349) );
  OR2_X1 U12805 ( .A1(n9970), .A2(n10349), .ZN(n10350) );
  NAND4_X1 U12806 ( .A1(n10353), .A2(n10352), .A3(n10351), .A4(n10350), .ZN(
        n14828) );
  NAND2_X1 U12807 ( .A1(n14423), .A2(n10423), .ZN(n10355) );
  OR2_X1 U12808 ( .A1(n10424), .A2(n15095), .ZN(n10354) );
  MUX2_X1 U12809 ( .A(n14828), .B(n14762), .S(n9951), .Z(n10359) );
  NAND2_X1 U12810 ( .A1(n10358), .A2(n10359), .ZN(n10357) );
  MUX2_X1 U12811 ( .A(n14828), .B(n14762), .S(n10428), .Z(n10356) );
  NAND2_X1 U12812 ( .A1(n10357), .A2(n10356), .ZN(n10363) );
  INV_X1 U12813 ( .A(n10358), .ZN(n10361) );
  INV_X1 U12814 ( .A(n10359), .ZN(n10360) );
  NAND2_X1 U12815 ( .A1(n10361), .A2(n10360), .ZN(n10362) );
  NAND2_X1 U12816 ( .A1(n9971), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n10371) );
  INV_X1 U12817 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n14800) );
  OR2_X1 U12818 ( .A1(n10404), .A2(n14800), .ZN(n10370) );
  INV_X1 U12819 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n10364) );
  NAND2_X1 U12820 ( .A1(n10365), .A2(n10364), .ZN(n10366) );
  NAND2_X1 U12821 ( .A1(n10378), .A2(n10366), .ZN(n14799) );
  OR2_X1 U12822 ( .A1(n6675), .A2(n14799), .ZN(n10369) );
  INV_X1 U12823 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10367) );
  OR2_X1 U12824 ( .A1(n9970), .A2(n10367), .ZN(n10368) );
  NAND4_X1 U12825 ( .A1(n10371), .A2(n10370), .A3(n10369), .A4(n10368), .ZN(
        n14764) );
  NAND2_X1 U12826 ( .A1(n14419), .A2(n10423), .ZN(n10373) );
  OR2_X1 U12827 ( .A1(n10424), .A2(n15092), .ZN(n10372) );
  MUX2_X1 U12828 ( .A(n14764), .B(n14802), .S(n10428), .Z(n10375) );
  MUX2_X1 U12829 ( .A(n14764), .B(n14802), .S(n9951), .Z(n10374) );
  NAND2_X1 U12830 ( .A1(n10417), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n10385) );
  INV_X1 U12831 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n10376) );
  OR2_X1 U12832 ( .A1(n10422), .A2(n10376), .ZN(n10384) );
  INV_X1 U12833 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n10377) );
  NAND2_X1 U12834 ( .A1(n10378), .A2(n10377), .ZN(n10379) );
  NAND2_X1 U12835 ( .A1(n14733), .A2(n10379), .ZN(n14775) );
  OR2_X1 U12836 ( .A1(n6674), .A2(n14775), .ZN(n10383) );
  INV_X1 U12837 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n10381) );
  OR2_X1 U12838 ( .A1(n9970), .A2(n10381), .ZN(n10382) );
  NAND4_X1 U12839 ( .A1(n10385), .A2(n10384), .A3(n10383), .A4(n10382), .ZN(
        n14789) );
  NAND2_X1 U12840 ( .A1(n14415), .A2(n10423), .ZN(n10387) );
  OR2_X1 U12841 ( .A1(n10424), .A2(n12716), .ZN(n10386) );
  MUX2_X1 U12842 ( .A(n14789), .B(n14779), .S(n9951), .Z(n10391) );
  NAND2_X1 U12843 ( .A1(n10390), .A2(n10391), .ZN(n10389) );
  MUX2_X1 U12844 ( .A(n14789), .B(n14779), .S(n10428), .Z(n10388) );
  NAND2_X1 U12845 ( .A1(n10389), .A2(n10388), .ZN(n10395) );
  INV_X1 U12846 ( .A(n10390), .ZN(n10393) );
  INV_X1 U12847 ( .A(n10391), .ZN(n10392) );
  NAND2_X1 U12848 ( .A1(n10393), .A2(n10392), .ZN(n10394) );
  NAND2_X1 U12849 ( .A1(n10395), .A2(n10394), .ZN(n10400) );
  INV_X1 U12850 ( .A(n10400), .ZN(n10398) );
  INV_X1 U12851 ( .A(n14989), .ZN(n14729) );
  MUX2_X1 U12852 ( .A(n14729), .B(n14549), .S(n10428), .Z(n10396) );
  OAI21_X1 U12853 ( .B1(n10398), .B2(n10397), .A(n10396), .ZN(n10399) );
  OAI21_X1 U12854 ( .B1(n10401), .B2(n10400), .A(n10399), .ZN(n10441) );
  INV_X1 U12855 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10402) );
  NOR2_X1 U12856 ( .A1(n10422), .A2(n10402), .ZN(n10408) );
  INV_X1 U12857 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n10403) );
  NOR2_X1 U12858 ( .A1(n10404), .A2(n10403), .ZN(n10407) );
  INV_X1 U12859 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10405) );
  NOR2_X1 U12860 ( .A1(n9970), .A2(n10405), .ZN(n10406) );
  NAND2_X1 U12861 ( .A1(n10409), .A2(n10423), .ZN(n10411) );
  INV_X1 U12862 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n15087) );
  OR2_X1 U12863 ( .A1(n10424), .A2(n15087), .ZN(n10410) );
  NAND2_X1 U12864 ( .A1(n10445), .A2(n10428), .ZN(n10444) );
  NOR2_X1 U12865 ( .A1(n10445), .A2(n10428), .ZN(n10452) );
  NAND2_X1 U12866 ( .A1(n10412), .A2(n9931), .ZN(n10578) );
  NAND2_X1 U12867 ( .A1(n10563), .A2(n12393), .ZN(n10511) );
  NAND2_X1 U12868 ( .A1(n10578), .A2(n10511), .ZN(n10414) );
  OR2_X1 U12869 ( .A1(n10509), .A2(n14973), .ZN(n10413) );
  NAND2_X1 U12870 ( .A1(n10414), .A2(n10413), .ZN(n10453) );
  INV_X1 U12871 ( .A(n12393), .ZN(n10415) );
  NAND2_X1 U12872 ( .A1(n12513), .A2(n10415), .ZN(n10482) );
  NAND2_X1 U12873 ( .A1(n10453), .A2(n10482), .ZN(n10446) );
  AOI21_X1 U12874 ( .B1(n10452), .B2(n14690), .A(n10446), .ZN(n10416) );
  OAI21_X1 U12875 ( .B1(n14690), .B2(n10444), .A(n10416), .ZN(n10443) );
  INV_X1 U12876 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10421) );
  NAND2_X1 U12877 ( .A1(n10417), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n10420) );
  NAND2_X1 U12878 ( .A1(n10418), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n10419) );
  OAI211_X1 U12879 ( .C1(n10422), .C2(n10421), .A(n10420), .B(n10419), .ZN(
        n14731) );
  OAI21_X1 U12880 ( .B1(n14690), .B2(n12393), .A(n14731), .ZN(n10427) );
  NAND2_X1 U12881 ( .A1(n12705), .A2(n10423), .ZN(n10426) );
  OR2_X1 U12882 ( .A1(n10424), .A2(n13040), .ZN(n10425) );
  MUX2_X1 U12883 ( .A(n10427), .B(n14985), .S(n10428), .Z(n10436) );
  INV_X1 U12884 ( .A(n14985), .ZN(n10461) );
  NAND2_X1 U12885 ( .A1(n10461), .A2(n9951), .ZN(n10433) );
  NAND2_X1 U12886 ( .A1(n14690), .A2(n10428), .ZN(n10430) );
  NAND2_X1 U12887 ( .A1(n10430), .A2(n10429), .ZN(n10431) );
  NAND2_X1 U12888 ( .A1(n10431), .A2(n14731), .ZN(n10432) );
  NAND2_X1 U12889 ( .A1(n10433), .A2(n10432), .ZN(n10437) );
  NOR2_X1 U12890 ( .A1(n10443), .A2(n10442), .ZN(n10434) );
  XNOR2_X1 U12891 ( .A(n10445), .B(n14690), .ZN(n10460) );
  INV_X1 U12892 ( .A(n10453), .ZN(n10435) );
  NAND2_X1 U12893 ( .A1(n10460), .A2(n10435), .ZN(n10457) );
  INV_X1 U12894 ( .A(n10436), .ZN(n10439) );
  INV_X1 U12895 ( .A(n10437), .ZN(n10438) );
  AND2_X1 U12896 ( .A1(n10439), .A2(n10438), .ZN(n10450) );
  NOR2_X1 U12897 ( .A1(n10457), .A2(n10450), .ZN(n10440) );
  INV_X1 U12898 ( .A(n10442), .ZN(n10458) );
  INV_X1 U12899 ( .A(n10443), .ZN(n10451) );
  NOR3_X1 U12900 ( .A1(n10444), .A2(n14690), .A3(n10453), .ZN(n10449) );
  INV_X1 U12901 ( .A(n10444), .ZN(n10447) );
  XOR2_X1 U12902 ( .A(n10453), .B(n10452), .Z(n10454) );
  NAND4_X1 U12903 ( .A1(n10454), .A2(n14982), .A3(n10482), .A4(n14690), .ZN(
        n10455) );
  OAI211_X1 U12904 ( .C1(n10458), .C2(n10457), .A(n10456), .B(n10455), .ZN(
        n10459) );
  INV_X1 U12905 ( .A(n10459), .ZN(n10485) );
  INV_X1 U12906 ( .A(n10460), .ZN(n10480) );
  XOR2_X1 U12907 ( .A(n14731), .B(n10461), .Z(n10479) );
  XNOR2_X1 U12908 ( .A(n14762), .B(n14761), .ZN(n14807) );
  XNOR2_X1 U12909 ( .A(n15014), .B(n14846), .ZN(n14838) );
  INV_X1 U12910 ( .A(n14826), .ZN(n14480) );
  NAND2_X1 U12911 ( .A1(n14859), .A2(n14480), .ZN(n14759) );
  OR2_X1 U12912 ( .A1(n14859), .A2(n14480), .ZN(n10462) );
  NAND2_X1 U12913 ( .A1(n14759), .A2(n10462), .ZN(n14848) );
  XNOR2_X1 U12914 ( .A(n15046), .B(n14710), .ZN(n14913) );
  XNOR2_X1 U12915 ( .A(n15057), .B(n14489), .ZN(n14745) );
  INV_X1 U12916 ( .A(n10463), .ZN(n14950) );
  NAND2_X1 U12917 ( .A1(n14741), .A2(n10464), .ZN(n12692) );
  INV_X1 U12918 ( .A(n14551), .ZN(n15305) );
  XNOR2_X1 U12919 ( .A(n15342), .B(n15305), .ZN(n12620) );
  XNOR2_X1 U12920 ( .A(n12687), .B(n14552), .ZN(n12615) );
  INV_X1 U12921 ( .A(n14554), .ZN(n12601) );
  OR2_X1 U12922 ( .A1(n15543), .A2(n12601), .ZN(n12529) );
  NAND2_X1 U12923 ( .A1(n15543), .A2(n12601), .ZN(n10465) );
  XNOR2_X1 U12924 ( .A(n12248), .B(n12247), .ZN(n12242) );
  INV_X1 U12925 ( .A(n14556), .ZN(n12551) );
  XNOR2_X1 U12926 ( .A(n12302), .B(n12551), .ZN(n12297) );
  INV_X1 U12927 ( .A(n11506), .ZN(n12115) );
  INV_X1 U12928 ( .A(n11912), .ZN(n10466) );
  OAI21_X1 U12929 ( .B1(n11616), .B2(n12115), .A(n10466), .ZN(n11445) );
  NOR4_X1 U12930 ( .A1(n11445), .A2(n12130), .A3(n11919), .A4(n15500), .ZN(
        n10468) );
  NAND2_X1 U12931 ( .A1(n12083), .A2(n14559), .ZN(n10467) );
  NAND2_X1 U12932 ( .A1(n11696), .A2(n12006), .ZN(n12000) );
  XNOR2_X1 U12933 ( .A(n12055), .B(n14558), .ZN(n12049) );
  XNOR2_X2 U12934 ( .A(n14560), .B(n14508), .ZN(n12163) );
  NAND4_X1 U12935 ( .A1(n10468), .A2(n12003), .A3(n12049), .A4(n12163), .ZN(
        n10469) );
  NOR4_X1 U12936 ( .A1(n12526), .A2(n12242), .A3(n12297), .A4(n10469), .ZN(
        n10470) );
  XNOR2_X1 U12937 ( .A(n15403), .B(n14553), .ZN(n12531) );
  XNOR2_X1 U12938 ( .A(n12554), .B(n14555), .ZN(n12301) );
  NAND4_X1 U12939 ( .A1(n12615), .A2(n10470), .A3(n12531), .A4(n12301), .ZN(
        n10471) );
  NOR4_X1 U12940 ( .A1(n12692), .A2(n7014), .A3(n12620), .A4(n10471), .ZN(
        n10472) );
  XNOR2_X1 U12941 ( .A(n15371), .B(n14703), .ZN(n14961) );
  NAND3_X1 U12942 ( .A1(n14950), .A2(n10472), .A3(n14961), .ZN(n10473) );
  NOR4_X1 U12943 ( .A1(n14913), .A2(n14928), .A3(n14745), .A4(n10473), .ZN(
        n10474) );
  XNOR2_X1 U12944 ( .A(n15024), .B(n14717), .ZN(n14864) );
  XNOR2_X1 U12945 ( .A(n14884), .B(n14714), .ZN(n14877) );
  NAND4_X1 U12946 ( .A1(n10474), .A2(n14864), .A3(n14877), .A4(n14891), .ZN(
        n10475) );
  NOR4_X1 U12947 ( .A1(n14807), .A2(n14838), .A3(n14848), .A4(n10475), .ZN(
        n10477) );
  NAND2_X1 U12948 ( .A1(n14779), .A2(n14789), .ZN(n14724) );
  OR2_X1 U12949 ( .A1(n14779), .A2(n14789), .ZN(n10476) );
  NAND2_X1 U12950 ( .A1(n14724), .A2(n10476), .ZN(n14770) );
  NAND4_X1 U12951 ( .A1(n14765), .A2(n10477), .A3(n14770), .A4(n14794), .ZN(
        n10478) );
  XOR2_X1 U12952 ( .A(n14814), .B(n10481), .Z(n10483) );
  INV_X1 U12953 ( .A(n10482), .ZN(n10579) );
  NAND2_X1 U12954 ( .A1(n10483), .A2(n10579), .ZN(n10484) );
  INV_X1 U12955 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n10488) );
  INV_X1 U12956 ( .A(n10782), .ZN(n10490) );
  NAND2_X1 U12957 ( .A1(n10490), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12630) );
  INV_X1 U12958 ( .A(n10578), .ZN(n10783) );
  NAND2_X1 U12959 ( .A1(n12393), .A2(n14973), .ZN(n10564) );
  NAND2_X1 U12960 ( .A1(n10783), .A2(n10564), .ZN(n11435) );
  INV_X1 U12961 ( .A(n10492), .ZN(n10493) );
  NAND2_X1 U12962 ( .A1(n10493), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10494) );
  XNOR2_X1 U12963 ( .A(n10494), .B(P1_IR_REG_25__SCAN_IN), .ZN(n10561) );
  NAND2_X1 U12964 ( .A1(n10495), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10496) );
  XNOR2_X1 U12965 ( .A(n10496), .B(P1_IR_REG_24__SCAN_IN), .ZN(n10559) );
  NAND2_X1 U12966 ( .A1(n10497), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10498) );
  AND2_X1 U12967 ( .A1(n10782), .A2(n10543), .ZN(n10500) );
  NAND2_X1 U12968 ( .A1(n11435), .A2(n10500), .ZN(n10574) );
  INV_X1 U12969 ( .A(n6678), .ZN(n15443) );
  NAND2_X1 U12970 ( .A1(n15443), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10502) );
  NOR3_X1 U12971 ( .A1(n10574), .A2(n14966), .A3(n10502), .ZN(n10504) );
  OAI21_X1 U12972 ( .B1(n12630), .B2(n10412), .A(P1_B_REG_SCAN_IN), .ZN(n10503) );
  OR2_X1 U12973 ( .A1(n10504), .A2(n10503), .ZN(n10505) );
  NAND2_X1 U12974 ( .A1(n10506), .A2(n10505), .ZN(P1_U3242) );
  INV_X1 U12975 ( .A(n10543), .ZN(n10508) );
  AND2_X2 U12976 ( .A1(n10790), .A2(n10508), .ZN(P1_U4016) );
  INV_X2 U12977 ( .A(n12787), .ZN(n10525) );
  NAND2_X1 U12978 ( .A1(n10509), .A2(n10543), .ZN(n10512) );
  OR2_X1 U12979 ( .A1(n15518), .A2(n12785), .ZN(n10510) );
  NAND2_X1 U12980 ( .A1(n11439), .A2(n10509), .ZN(n10528) );
  INV_X2 U12981 ( .A(n12819), .ZN(n12672) );
  INV_X4 U12982 ( .A(n12788), .ZN(n12848) );
  NAND2_X1 U12983 ( .A1(n14561), .A2(n12848), .ZN(n10514) );
  OR2_X1 U12984 ( .A1(n15518), .A2(n12787), .ZN(n10513) );
  NAND2_X1 U12985 ( .A1(n10514), .A2(n10513), .ZN(n11667) );
  XNOR2_X1 U12986 ( .A(n11668), .B(n11667), .ZN(n10569) );
  OAI22_X1 U12987 ( .A1(n11508), .A2(n12788), .B1(n11920), .B2(n12787), .ZN(
        n10515) );
  INV_X1 U12988 ( .A(n10515), .ZN(n10532) );
  NAND2_X1 U12989 ( .A1(n11443), .A2(n10525), .ZN(n10517) );
  OAI22_X1 U12990 ( .A1(n11506), .A2(n12785), .B1(n10543), .B2(n10523), .ZN(
        n10524) );
  INV_X1 U12991 ( .A(n11373), .ZN(n10530) );
  NAND2_X1 U12992 ( .A1(n11372), .A2(n10531), .ZN(n11612) );
  INV_X1 U12993 ( .A(n10533), .ZN(n10534) );
  NAND2_X1 U12994 ( .A1(n10536), .A2(n10525), .ZN(n10538) );
  OR2_X1 U12995 ( .A1(n15513), .A2(n12785), .ZN(n10537) );
  NAND2_X1 U12996 ( .A1(n10538), .A2(n10537), .ZN(n10539) );
  XNOR2_X1 U12997 ( .A(n10539), .B(n12672), .ZN(n10540) );
  AOI22_X1 U12998 ( .A1(n10536), .A2(n12848), .B1(n11936), .B2(n10525), .ZN(
        n10541) );
  XNOR2_X1 U12999 ( .A(n10540), .B(n10541), .ZN(n11379) );
  INV_X1 U13000 ( .A(n10540), .ZN(n10542) );
  NAND2_X1 U13001 ( .A1(n10542), .A2(n10541), .ZN(n11675) );
  NAND2_X1 U13002 ( .A1(n11683), .A2(n11675), .ZN(n10568) );
  AND2_X1 U13003 ( .A1(n10790), .A2(n10543), .ZN(n10780) );
  INV_X1 U13004 ( .A(P1_B_REG_SCAN_IN), .ZN(n14688) );
  NOR2_X1 U13005 ( .A1(n10561), .A2(n14688), .ZN(n10544) );
  MUX2_X1 U13006 ( .A(n10544), .B(n14688), .S(n10559), .Z(n10545) );
  INV_X1 U13007 ( .A(n10545), .ZN(n10546) );
  NOR2_X1 U13008 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n10550) );
  NOR4_X1 U13009 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n10549) );
  NOR4_X1 U13010 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n10548) );
  NOR4_X1 U13011 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n10547) );
  NAND4_X1 U13012 ( .A1(n10550), .A2(n10549), .A3(n10548), .A4(n10547), .ZN(
        n10556) );
  NOR4_X1 U13013 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n10554) );
  NOR4_X1 U13014 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n10553) );
  NOR4_X1 U13015 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n10552) );
  NOR4_X1 U13016 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n10551) );
  NAND4_X1 U13017 ( .A1(n10554), .A2(n10553), .A3(n10552), .A4(n10551), .ZN(
        n10555) );
  NOR2_X1 U13018 ( .A1(n10556), .A2(n10555), .ZN(n10572) );
  NAND2_X1 U13019 ( .A1(n10780), .A2(n10572), .ZN(n10557) );
  OR2_X1 U13020 ( .A1(n10571), .A2(P1_D_REG_0__SCAN_IN), .ZN(n10560) );
  INV_X1 U13021 ( .A(n10558), .ZN(n15097) );
  INV_X1 U13022 ( .A(n10559), .ZN(n15105) );
  NAND2_X1 U13023 ( .A1(n15097), .A2(n15105), .ZN(n10785) );
  OR2_X1 U13024 ( .A1(n10571), .A2(P1_D_REG_1__SCAN_IN), .ZN(n10562) );
  INV_X1 U13025 ( .A(n10561), .ZN(n15100) );
  NAND2_X1 U13026 ( .A1(n15097), .A2(n15100), .ZN(n10788) );
  AND2_X1 U13027 ( .A1(n10562), .A2(n10788), .ZN(n11433) );
  AND2_X1 U13028 ( .A1(n14732), .A2(n11433), .ZN(n10570) );
  INV_X1 U13029 ( .A(n10570), .ZN(n10580) );
  AND2_X1 U13030 ( .A1(n12513), .A2(n10564), .ZN(n10565) );
  NAND2_X1 U13031 ( .A1(n15545), .A2(n10578), .ZN(n10566) );
  NOR2_X1 U13032 ( .A1(n10580), .A2(n10566), .ZN(n10567) );
  AOI211_X1 U13033 ( .C1(n10569), .C2(n10568), .A(n15337), .B(n11688), .ZN(
        n10587) );
  OAI21_X1 U13034 ( .B1(n10572), .B2(n10571), .A(n10570), .ZN(n10573) );
  NAND2_X1 U13035 ( .A1(n10573), .A2(n11436), .ZN(n10576) );
  INV_X1 U13036 ( .A(n10574), .ZN(n10575) );
  NAND2_X1 U13037 ( .A1(n10576), .A2(n10575), .ZN(n11374) );
  INV_X1 U13038 ( .A(n15369), .ZN(n14532) );
  MUX2_X1 U13039 ( .A(n14532), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n10586) );
  AND2_X1 U13040 ( .A1(n11435), .A2(n11433), .ZN(n10577) );
  NAND2_X1 U13041 ( .A1(n15348), .A2(n14825), .ZN(n15361) );
  INV_X1 U13042 ( .A(n10536), .ZN(n11615) );
  NOR2_X1 U13043 ( .A1(n15361), .A2(n11615), .ZN(n10585) );
  NAND2_X1 U13044 ( .A1(n15348), .A2(n14827), .ZN(n15360) );
  INV_X1 U13045 ( .A(n14560), .ZN(n11929) );
  NAND2_X1 U13046 ( .A1(n10563), .A2(n10579), .ZN(n11826) );
  NOR2_X1 U13047 ( .A1(n10580), .A2(n11826), .ZN(n10581) );
  NAND2_X1 U13048 ( .A1(n11438), .A2(n10581), .ZN(n10583) );
  INV_X1 U13049 ( .A(n15351), .ZN(n15358) );
  OAI22_X1 U13050 ( .A1(n15360), .A2(n11929), .B1(n15518), .B2(n15358), .ZN(
        n10584) );
  OR4_X1 U13051 ( .A1(n10587), .A2(n10586), .A3(n10585), .A4(n10584), .ZN(
        P1_U3218) );
  INV_X1 U13052 ( .A(n13685), .ZN(n11266) );
  NAND2_X1 U13053 ( .A1(n10712), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10598) );
  OAI21_X1 U13054 ( .B1(n10712), .B2(P3_REG1_REG_6__SCAN_IN), .A(n10598), .ZN(
        n11290) );
  NAND2_X1 U13055 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n7369), .ZN(n11245) );
  NAND2_X1 U13056 ( .A1(n11023), .A2(n11245), .ZN(n10591) );
  INV_X1 U13057 ( .A(n11245), .ZN(n10589) );
  NAND2_X1 U13058 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10589), .ZN(n10590) );
  NAND2_X1 U13059 ( .A1(n10591), .A2(n10590), .ZN(n11007) );
  NAND2_X1 U13060 ( .A1(n11007), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n11006) );
  OR2_X1 U13061 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n11245), .ZN(n10592) );
  NAND2_X1 U13062 ( .A1(n11006), .A2(n10592), .ZN(n11056) );
  OR2_X1 U13063 ( .A1(n11069), .A2(n10640), .ZN(n10593) );
  NAND2_X1 U13064 ( .A1(n11055), .A2(n10593), .ZN(n10594) );
  NAND2_X1 U13065 ( .A1(n10594), .A2(n11030), .ZN(n11146) );
  OR2_X1 U13066 ( .A1(n10594), .A2(n11030), .ZN(n10595) );
  XNOR2_X1 U13067 ( .A(n11162), .B(n11552), .ZN(n11147) );
  NOR2_X1 U13068 ( .A1(n10597), .A2(n11202), .ZN(n11291) );
  INV_X1 U13069 ( .A(n10598), .ZN(n10599) );
  NOR2_X1 U13070 ( .A1(n11315), .A2(n10600), .ZN(n10601) );
  NAND2_X1 U13071 ( .A1(n10737), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n10602) );
  OAI21_X1 U13072 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n10737), .A(n10602), .ZN(
        n11405) );
  NOR2_X1 U13073 ( .A1(n10677), .A2(n10603), .ZN(n10604) );
  OR2_X1 U13074 ( .A1(n10681), .A2(n15852), .ZN(n12410) );
  NAND2_X1 U13075 ( .A1(n10681), .A2(n15852), .ZN(n10605) );
  NAND2_X1 U13076 ( .A1(n12410), .A2(n10605), .ZN(n10606) );
  NAND2_X1 U13077 ( .A1(n10607), .A2(n10606), .ZN(n10613) );
  NAND2_X1 U13078 ( .A1(n10608), .A2(n13245), .ZN(n10692) );
  OR2_X1 U13079 ( .A1(n13228), .A2(n10609), .ZN(n10610) );
  AND2_X1 U13080 ( .A1(n10611), .A2(n10610), .ZN(n10690) );
  NAND2_X1 U13081 ( .A1(n10692), .A2(n10690), .ZN(n10688) );
  AOI21_X1 U13082 ( .B1(n12411), .B2(n10613), .A(n15744), .ZN(n10697) );
  INV_X1 U13083 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11701) );
  NAND2_X1 U13084 ( .A1(n10712), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10620) );
  OAI21_X1 U13085 ( .B1(n10712), .B2(P3_REG2_REG_6__SCAN_IN), .A(n10620), .ZN(
        n11286) );
  XNOR2_X1 U13086 ( .A(n11069), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n11053) );
  INV_X1 U13087 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11470) );
  NOR2_X1 U13088 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n11470), .ZN(n11240) );
  NAND2_X1 U13089 ( .A1(n10614), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10615) );
  OAI21_X1 U13090 ( .B1(n11023), .B2(n11240), .A(n10615), .ZN(n11016) );
  INV_X1 U13091 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n11015) );
  OR2_X1 U13092 ( .A1(n11016), .A2(n11015), .ZN(n11018) );
  NAND2_X1 U13093 ( .A1(n11018), .A2(n10615), .ZN(n11052) );
  NAND2_X1 U13094 ( .A1(n11053), .A2(n11052), .ZN(n11051) );
  INV_X1 U13095 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10641) );
  OR2_X1 U13096 ( .A1(n11069), .A2(n10641), .ZN(n10616) );
  INV_X1 U13097 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10652) );
  XNOR2_X1 U13098 ( .A(n11162), .B(n10652), .ZN(n11141) );
  AOI21_X1 U13099 ( .B1(n11142), .B2(n11140), .A(n11141), .ZN(n11144) );
  AOI21_X1 U13100 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n10706), .A(n11144), .ZN(
        n10617) );
  NOR2_X1 U13101 ( .A1(n10617), .A2(n11209), .ZN(n10619) );
  INV_X1 U13102 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11200) );
  INV_X1 U13103 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11307) );
  NAND2_X1 U13104 ( .A1(n10737), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n10622) );
  OAI21_X1 U13105 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n10737), .A(n10622), .ZN(
        n11408) );
  NOR2_X1 U13106 ( .A1(n11701), .A2(n11700), .ZN(n11699) );
  NOR2_X1 U13107 ( .A1(n10677), .A2(n10625), .ZN(n10626) );
  INV_X1 U13108 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n12327) );
  OR2_X1 U13109 ( .A1(n10681), .A2(n12327), .ZN(n12423) );
  NAND2_X1 U13110 ( .A1(n10681), .A2(n12327), .ZN(n10627) );
  NAND2_X1 U13111 ( .A1(n12423), .A2(n10627), .ZN(n10630) );
  INV_X1 U13112 ( .A(n10630), .ZN(n10628) );
  NAND2_X1 U13113 ( .A1(n10631), .A2(n10630), .ZN(n10633) );
  AOI21_X1 U13114 ( .B1(n12424), .B2(n10633), .A(n15752), .ZN(n10696) );
  MUX2_X1 U13115 ( .A(n11015), .B(n10634), .S(n6671), .Z(n10636) );
  INV_X1 U13116 ( .A(n11023), .ZN(n10635) );
  NAND2_X1 U13117 ( .A1(n10636), .A2(n10635), .ZN(n11060) );
  INV_X1 U13118 ( .A(n10636), .ZN(n10637) );
  NAND2_X1 U13119 ( .A1(n10637), .A2(n11023), .ZN(n10638) );
  NAND2_X1 U13120 ( .A1(n11060), .A2(n10638), .ZN(n11009) );
  MUX2_X1 U13121 ( .A(n11470), .B(n10639), .S(n6671), .Z(n11246) );
  NAND2_X1 U13122 ( .A1(n11246), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11239) );
  MUX2_X1 U13123 ( .A(n10641), .B(n10640), .S(n6671), .Z(n10642) );
  NAND2_X1 U13124 ( .A1(n10642), .A2(n11069), .ZN(n10645) );
  INV_X1 U13125 ( .A(n10642), .ZN(n10643) );
  INV_X1 U13126 ( .A(n11069), .ZN(n10727) );
  NAND2_X1 U13127 ( .A1(n10643), .A2(n10727), .ZN(n10644) );
  NAND2_X1 U13128 ( .A1(n10645), .A2(n10644), .ZN(n11059) );
  AOI21_X1 U13129 ( .B1(n11061), .B2(n11060), .A(n11059), .ZN(n11063) );
  INV_X1 U13130 ( .A(n10645), .ZN(n11035) );
  INV_X1 U13131 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10647) );
  MUX2_X1 U13132 ( .A(n10647), .B(n10646), .S(n6670), .Z(n10649) );
  NAND2_X1 U13133 ( .A1(n10649), .A2(n10648), .ZN(n11156) );
  INV_X1 U13134 ( .A(n10649), .ZN(n10650) );
  NAND2_X1 U13135 ( .A1(n10650), .A2(n11030), .ZN(n10651) );
  AND2_X1 U13136 ( .A1(n11156), .A2(n10651), .ZN(n11034) );
  OAI21_X1 U13137 ( .B1(n11063), .B2(n11035), .A(n11034), .ZN(n11157) );
  MUX2_X1 U13138 ( .A(n10652), .B(n11552), .S(n8267), .Z(n10653) );
  NAND2_X1 U13139 ( .A1(n10653), .A2(n11162), .ZN(n10656) );
  INV_X1 U13140 ( .A(n10653), .ZN(n10654) );
  NAND2_X1 U13141 ( .A1(n10654), .A2(n10706), .ZN(n10655) );
  NAND2_X1 U13142 ( .A1(n10656), .A2(n10655), .ZN(n11155) );
  INV_X1 U13143 ( .A(n10656), .ZN(n11211) );
  MUX2_X1 U13144 ( .A(n11200), .B(n10657), .S(n8267), .Z(n10658) );
  NAND2_X1 U13145 ( .A1(n10658), .A2(n11209), .ZN(n11297) );
  INV_X1 U13146 ( .A(n10658), .ZN(n10659) );
  NAND2_X1 U13147 ( .A1(n10659), .A2(n10703), .ZN(n10660) );
  AND2_X1 U13148 ( .A1(n11297), .A2(n10660), .ZN(n11210) );
  OAI21_X1 U13149 ( .B1(n11212), .B2(n11211), .A(n11210), .ZN(n11298) );
  INV_X1 U13150 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11772) );
  MUX2_X1 U13151 ( .A(n11772), .B(n10661), .S(n10612), .Z(n10662) );
  INV_X1 U13152 ( .A(n10712), .ZN(n11303) );
  NAND2_X1 U13153 ( .A1(n10662), .A2(n11303), .ZN(n10665) );
  INV_X1 U13154 ( .A(n10662), .ZN(n10663) );
  NAND2_X1 U13155 ( .A1(n10663), .A2(n10712), .ZN(n10664) );
  NAND2_X1 U13156 ( .A1(n10665), .A2(n10664), .ZN(n11296) );
  AOI21_X1 U13157 ( .B1(n11298), .B2(n11297), .A(n11296), .ZN(n11310) );
  INV_X1 U13158 ( .A(n10665), .ZN(n11309) );
  MUX2_X1 U13159 ( .A(n11307), .B(n10666), .S(n10612), .Z(n10667) );
  NAND2_X1 U13160 ( .A1(n10667), .A2(n11315), .ZN(n11416) );
  INV_X1 U13161 ( .A(n10667), .ZN(n10668) );
  NAND2_X1 U13162 ( .A1(n10668), .A2(n10733), .ZN(n10669) );
  AND2_X1 U13163 ( .A1(n11416), .A2(n10669), .ZN(n11308) );
  OAI21_X1 U13164 ( .B1(n11310), .B2(n11309), .A(n11308), .ZN(n11417) );
  INV_X1 U13165 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n15758) );
  MUX2_X1 U13166 ( .A(n15758), .B(n10670), .S(n10612), .Z(n10671) );
  INV_X1 U13167 ( .A(n10737), .ZN(n11414) );
  NAND2_X1 U13168 ( .A1(n10671), .A2(n11414), .ZN(n10674) );
  INV_X1 U13169 ( .A(n10671), .ZN(n10672) );
  NAND2_X1 U13170 ( .A1(n10672), .A2(n10737), .ZN(n10673) );
  NAND2_X1 U13171 ( .A1(n10674), .A2(n10673), .ZN(n11415) );
  INV_X1 U13172 ( .A(n10674), .ZN(n11706) );
  MUX2_X1 U13173 ( .A(n11701), .B(n10675), .S(n10612), .Z(n10676) );
  NAND2_X1 U13174 ( .A1(n10676), .A2(n10677), .ZN(n10685) );
  INV_X1 U13175 ( .A(n10676), .ZN(n10678) );
  NAND2_X1 U13176 ( .A1(n10678), .A2(n10623), .ZN(n10679) );
  AND2_X1 U13177 ( .A1(n10685), .A2(n10679), .ZN(n11705) );
  OAI21_X1 U13178 ( .B1(n11707), .B2(n11706), .A(n11705), .ZN(n11704) );
  MUX2_X1 U13179 ( .A(n12327), .B(n15852), .S(n10612), .Z(n10680) );
  NAND2_X1 U13180 ( .A1(n10680), .A2(n10681), .ZN(n12417) );
  INV_X1 U13181 ( .A(n10680), .ZN(n10682) );
  INV_X1 U13182 ( .A(n10681), .ZN(n10721) );
  NAND2_X1 U13183 ( .A1(n10682), .A2(n10721), .ZN(n10683) );
  NAND2_X1 U13184 ( .A1(n12417), .A2(n10683), .ZN(n10684) );
  AOI21_X1 U13185 ( .B1(n11704), .B2(n10685), .A(n10684), .ZN(n12419) );
  INV_X1 U13186 ( .A(n12419), .ZN(n10687) );
  NAND3_X1 U13187 ( .A1(n11704), .A2(n10685), .A3(n10684), .ZN(n10686) );
  INV_X1 U13188 ( .A(n8266), .ZN(n13240) );
  NOR2_X2 U13189 ( .A1(n10689), .A2(n13240), .ZN(n13395) );
  INV_X1 U13190 ( .A(n13395), .ZN(n15746) );
  AOI21_X1 U13191 ( .B1(n10687), .B2(n10686), .A(n15746), .ZN(n10695) );
  MUX2_X1 U13192 ( .A(n10689), .B(n10688), .S(n8266), .Z(n15738) );
  NAND2_X1 U13193 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n12519)
         );
  INV_X1 U13194 ( .A(n10690), .ZN(n10691) );
  NAND2_X1 U13195 ( .A1(n15732), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n10693) );
  OAI211_X1 U13196 ( .C1(n15738), .C2(n10721), .A(n12519), .B(n10693), .ZN(
        n10694) );
  OR4_X1 U13197 ( .A1(n10697), .A2(n10696), .A3(n10695), .A4(n10694), .ZN(
        P3_U3192) );
  AND2_X1 U13198 ( .A1(n10717), .A2(P2_U3088), .ZN(n14414) );
  INV_X2 U13199 ( .A(n14414), .ZN(n14428) );
  NOR2_X1 U13200 ( .A1(n10717), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14421) );
  INV_X1 U13201 ( .A(n14421), .ZN(n14434) );
  OAI222_X1 U13202 ( .A1(n14428), .A2(n10722), .B1(n15562), .B2(P2_U3088), 
        .C1(n10698), .C2(n14434), .ZN(P2_U3326) );
  NOR2_X1 U13203 ( .A1(n10717), .A2(P3_STATE_REG_SCAN_IN), .ZN(n15121) );
  INV_X2 U13204 ( .A(n15121), .ZN(n13712) );
  INV_X1 U13205 ( .A(SI_3_), .ZN(n10699) );
  NAND2_X1 U13206 ( .A1(n10717), .A2(P3_U3151), .ZN(n13715) );
  OAI222_X1 U13207 ( .A1(n11030), .A2(P3_U3151), .B1(n13712), .B2(n10700), 
        .C1(n10699), .C2(n13715), .ZN(P3_U3292) );
  OAI222_X1 U13208 ( .A1(n10703), .A2(P3_U3151), .B1(n13712), .B2(n10702), 
        .C1(n10701), .C2(n13715), .ZN(P3_U3290) );
  OAI222_X1 U13209 ( .A1(n10706), .A2(P3_U3151), .B1(n13712), .B2(n10705), 
        .C1(n10704), .C2(n13715), .ZN(P3_U3291) );
  INV_X1 U13210 ( .A(n10707), .ZN(n10708) );
  OAI222_X1 U13211 ( .A1(P3_U3151), .A2(n7369), .B1(n13712), .B2(n10708), .C1(
        n9388), .C2(n13715), .ZN(P3_U3295) );
  INV_X1 U13212 ( .A(n10709), .ZN(n10711) );
  OAI222_X1 U13213 ( .A1(P3_U3151), .A2(n10712), .B1(n13712), .B2(n10711), 
        .C1(n10710), .C2(n13715), .ZN(P3_U3289) );
  AOI22_X1 U13214 ( .A1(n14421), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n10812), .ZN(n10714) );
  OAI21_X1 U13215 ( .B1(n9964), .B2(n14428), .A(n10714), .ZN(P2_U3325) );
  AOI22_X1 U13216 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n14421), .B1(n13950), 
        .B2(P2_STATE_REG_SCAN_IN), .ZN(n10716) );
  OAI21_X1 U13217 ( .B1(n9976), .B2(n14428), .A(n10716), .ZN(P2_U3324) );
  NAND2_X1 U13218 ( .A1(n10717), .A2(P1_U3086), .ZN(n15086) );
  INV_X1 U13219 ( .A(n15086), .ZN(n10850) );
  INV_X1 U13220 ( .A(n10850), .ZN(n15101) );
  NOR2_X1 U13221 ( .A1(n10717), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15090) );
  OAI222_X1 U13222 ( .A1(n15101), .A2(n10718), .B1(n15104), .B2(n9964), .C1(
        P1_U3086), .C2(n14584), .ZN(P1_U3353) );
  OAI222_X1 U13223 ( .A1(P3_U3151), .A2(n10721), .B1(n13715), .B2(n10720), 
        .C1(n13712), .C2(n10719), .ZN(P3_U3285) );
  OAI222_X1 U13224 ( .A1(P1_U3086), .A2(n14598), .B1(n15104), .B2(n9976), .C1(
        n6986), .C2(n15086), .ZN(P1_U3352) );
  OAI222_X1 U13225 ( .A1(n15086), .A2(n8403), .B1(n15104), .B2(n10722), .C1(
        P1_U3086), .C2(n10920), .ZN(P1_U3354) );
  AOI22_X1 U13226 ( .A1(n13964), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n14421), .ZN(n10723) );
  OAI21_X1 U13227 ( .B1(n9996), .B2(n14428), .A(n10723), .ZN(P2_U3323) );
  INV_X1 U13228 ( .A(n13715), .ZN(n15120) );
  INV_X1 U13229 ( .A(n15120), .ZN(n13709) );
  OAI222_X1 U13230 ( .A1(n12426), .A2(P3_U3151), .B1(n13712), .B2(n10725), 
        .C1(n13709), .C2(n10724), .ZN(P3_U3284) );
  OAI222_X1 U13231 ( .A1(n10727), .A2(P3_U3151), .B1(n13712), .B2(n10726), 
        .C1(n7663), .C2(n13709), .ZN(P3_U3293) );
  OAI222_X1 U13232 ( .A1(n13712), .A2(n7761), .B1(n13709), .B2(n10728), .C1(
        P3_U3151), .C2(n11023), .ZN(P3_U3294) );
  INV_X1 U13233 ( .A(n15459), .ZN(n10730) );
  INV_X1 U13234 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10729) );
  OAI222_X1 U13235 ( .A1(P1_U3086), .A2(n10730), .B1(n15104), .B2(n9996), .C1(
        n10729), .C2(n15086), .ZN(P1_U3351) );
  OAI222_X1 U13236 ( .A1(P3_U3151), .A2(n10733), .B1(n13715), .B2(n10732), 
        .C1(n13712), .C2(n10731), .ZN(P3_U3288) );
  INV_X1 U13237 ( .A(n10734), .ZN(n10735) );
  OAI222_X1 U13238 ( .A1(P3_U3151), .A2(n10737), .B1(n13709), .B2(n10736), 
        .C1(n13712), .C2(n10735), .ZN(P3_U3287) );
  INV_X1 U13239 ( .A(SI_9_), .ZN(n10739) );
  OAI222_X1 U13240 ( .A1(P3_U3151), .A2(n10623), .B1(n13715), .B2(n10739), 
        .C1(n13712), .C2(n10738), .ZN(P3_U3286) );
  INV_X1 U13241 ( .A(n10740), .ZN(n10741) );
  OAI222_X1 U13242 ( .A1(n13715), .A2(n10742), .B1(n13712), .B2(n10741), .C1(
        P3_U3151), .C2(n13255), .ZN(P3_U3283) );
  INV_X1 U13243 ( .A(n10743), .ZN(n10745) );
  AOI22_X1 U13244 ( .A1(n13980), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n14421), .ZN(n10744) );
  OAI21_X1 U13245 ( .B1(n10745), .B2(n14428), .A(n10744), .ZN(P2_U3322) );
  INV_X1 U13246 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10746) );
  INV_X1 U13247 ( .A(n14610), .ZN(n10908) );
  OAI222_X1 U13248 ( .A1(n15101), .A2(n10746), .B1(n15104), .B2(n10745), .C1(
        P1_U3086), .C2(n10908), .ZN(P1_U3350) );
  INV_X1 U13249 ( .A(n10923), .ZN(n11081) );
  OAI222_X1 U13250 ( .A1(P1_U3086), .A2(n11081), .B1(n15104), .B2(n10748), 
        .C1(n10747), .C2(n15086), .ZN(P1_U3349) );
  INV_X1 U13251 ( .A(n13995), .ZN(n10749) );
  OAI222_X1 U13252 ( .A1(n14434), .A2(n10750), .B1(n10749), .B2(P2_U3088), 
        .C1(n14428), .C2(n10748), .ZN(P2_U3321) );
  INV_X1 U13253 ( .A(n14627), .ZN(n14623) );
  OAI222_X1 U13254 ( .A1(P1_U3086), .A2(n14623), .B1(n15104), .B2(n10752), 
        .C1(n10751), .C2(n15086), .ZN(P1_U3348) );
  INV_X1 U13255 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10753) );
  INV_X1 U13256 ( .A(n14011), .ZN(n14003) );
  OAI222_X1 U13257 ( .A1(n14434), .A2(n10753), .B1(n14003), .B2(P2_U3088), 
        .C1(n14428), .C2(n10752), .ZN(P2_U3320) );
  INV_X1 U13258 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10754) );
  OR2_X1 U13259 ( .A1(n15562), .A2(n10754), .ZN(n10758) );
  NAND2_X1 U13260 ( .A1(n15562), .A2(n10754), .ZN(n10755) );
  NAND2_X1 U13261 ( .A1(n10758), .A2(n10755), .ZN(n15566) );
  INV_X1 U13262 ( .A(n15566), .ZN(n10757) );
  AND2_X1 U13263 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n15565), .ZN(n10756) );
  NAND2_X1 U13264 ( .A1(n10757), .A2(n10756), .ZN(n15569) );
  NAND2_X1 U13265 ( .A1(n15569), .A2(n10758), .ZN(n10811) );
  INV_X1 U13266 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10759) );
  XNOR2_X1 U13267 ( .A(n10812), .B(n10759), .ZN(n10810) );
  XNOR2_X1 U13268 ( .A(n10811), .B(n10810), .ZN(n10779) );
  OAI21_X1 U13269 ( .B1(n10762), .B2(n10761), .A(n10760), .ZN(n10763) );
  INV_X1 U13270 ( .A(n10769), .ZN(n10768) );
  NAND2_X1 U13271 ( .A1(n10765), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14416) );
  INV_X1 U13272 ( .A(n14416), .ZN(n10766) );
  AND2_X1 U13273 ( .A1(n10768), .A2(n10766), .ZN(n10774) );
  NAND2_X1 U13274 ( .A1(n10774), .A2(n10767), .ZN(n12583) );
  AND2_X1 U13275 ( .A1(n9203), .A2(n10768), .ZN(n15561) );
  NAND2_X1 U13276 ( .A1(n15561), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14004) );
  INV_X1 U13277 ( .A(n14004), .ZN(n15641) );
  AND2_X1 U13278 ( .A1(n10769), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15635) );
  INV_X1 U13279 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11638) );
  OAI22_X1 U13280 ( .A1(n15592), .A2(n7312), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11638), .ZN(n10770) );
  AOI21_X1 U13281 ( .B1(n10812), .B2(n15641), .A(n10770), .ZN(n10778) );
  INV_X1 U13282 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10771) );
  MUX2_X1 U13283 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10771), .S(n10812), .Z(
        n10776) );
  XNOR2_X1 U13284 ( .A(n15562), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n15572) );
  AND2_X1 U13285 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n15565), .ZN(n15571) );
  NAND2_X1 U13286 ( .A1(n15572), .A2(n15571), .ZN(n15570) );
  NAND2_X1 U13287 ( .A1(n7592), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10772) );
  NAND2_X1 U13288 ( .A1(n15570), .A2(n10772), .ZN(n10775) );
  AND2_X1 U13289 ( .A1(n10774), .A2(n10773), .ZN(n15644) );
  NAND2_X1 U13290 ( .A1(n10775), .A2(n10776), .ZN(n13953) );
  OAI211_X1 U13291 ( .C1(n10776), .C2(n10775), .A(n15644), .B(n13953), .ZN(
        n10777) );
  OAI211_X1 U13292 ( .C1(n10779), .C2(n12583), .A(n10778), .B(n10777), .ZN(
        P2_U3216) );
  OR2_X1 U13293 ( .A1(n10780), .A2(n10491), .ZN(n10914) );
  AOI21_X1 U13294 ( .B1(n10783), .B2(n10782), .A(n10781), .ZN(n10913) );
  INV_X1 U13295 ( .A(n10913), .ZN(n10784) );
  AND2_X1 U13296 ( .A1(n10914), .A2(n10784), .ZN(n15450) );
  NOR2_X1 U13297 ( .A1(n15450), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U13298 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10787) );
  INV_X1 U13299 ( .A(n10785), .ZN(n10786) );
  AOI22_X1 U13300 ( .A1(n15510), .A2(n10787), .B1(n10786), .B2(n10790), .ZN(
        P1_U3445) );
  INV_X1 U13301 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10791) );
  INV_X1 U13302 ( .A(n10788), .ZN(n10789) );
  AOI22_X1 U13303 ( .A1(n15510), .A2(n10791), .B1(n10790), .B2(n10789), .ZN(
        P1_U3446) );
  AOI22_X1 U13304 ( .A1(n10942), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10850), .ZN(n10792) );
  OAI21_X1 U13305 ( .B1(n10793), .B2(n15104), .A(n10792), .ZN(P1_U3347) );
  INV_X1 U13306 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10795) );
  INV_X1 U13307 ( .A(n14026), .ZN(n10794) );
  OAI222_X1 U13308 ( .A1(n14434), .A2(n10795), .B1(n10794), .B2(P2_U3088), 
        .C1(n14428), .C2(n10793), .ZN(P2_U3319) );
  INV_X1 U13309 ( .A(n15644), .ZN(n12371) );
  INV_X1 U13310 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10796) );
  NOR2_X1 U13311 ( .A1(n12371), .A2(n10796), .ZN(n10834) );
  NAND2_X1 U13312 ( .A1(n10812), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n13951) );
  NAND2_X1 U13313 ( .A1(n13953), .A2(n13951), .ZN(n10798) );
  INV_X1 U13314 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11572) );
  MUX2_X1 U13315 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11572), .S(n13950), .Z(
        n10797) );
  NAND2_X1 U13316 ( .A1(n10798), .A2(n10797), .ZN(n13968) );
  NAND2_X1 U13317 ( .A1(n13950), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n13967) );
  NAND2_X1 U13318 ( .A1(n13968), .A2(n13967), .ZN(n10800) );
  INV_X1 U13319 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n13965) );
  MUX2_X1 U13320 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n13965), .S(n13964), .Z(
        n10799) );
  NAND2_X1 U13321 ( .A1(n10800), .A2(n10799), .ZN(n13978) );
  NAND2_X1 U13322 ( .A1(n13964), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n13977) );
  NAND2_X1 U13323 ( .A1(n13978), .A2(n13977), .ZN(n10802) );
  INV_X1 U13324 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11589) );
  MUX2_X1 U13325 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11589), .S(n13980), .Z(
        n10801) );
  NAND2_X1 U13326 ( .A1(n10802), .A2(n10801), .ZN(n13993) );
  NAND2_X1 U13327 ( .A1(n13980), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n13992) );
  NAND2_X1 U13328 ( .A1(n13993), .A2(n13992), .ZN(n10804) );
  INV_X1 U13329 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11578) );
  MUX2_X1 U13330 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11578), .S(n13995), .Z(
        n10803) );
  NAND2_X1 U13331 ( .A1(n10804), .A2(n10803), .ZN(n14009) );
  NAND2_X1 U13332 ( .A1(n13995), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n14008) );
  NAND2_X1 U13333 ( .A1(n14009), .A2(n14008), .ZN(n10806) );
  INV_X1 U13334 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11601) );
  MUX2_X1 U13335 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11601), .S(n14011), .Z(
        n10805) );
  NAND2_X1 U13336 ( .A1(n10806), .A2(n10805), .ZN(n14023) );
  NAND2_X1 U13337 ( .A1(n14011), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n14022) );
  NAND2_X1 U13338 ( .A1(n14023), .A2(n14022), .ZN(n10808) );
  INV_X1 U13339 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11867) );
  MUX2_X1 U13340 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11867), .S(n14026), .Z(
        n10807) );
  NAND2_X1 U13341 ( .A1(n10808), .A2(n10807), .ZN(n14025) );
  NAND2_X1 U13342 ( .A1(n14026), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10809) );
  NAND2_X1 U13343 ( .A1(n14025), .A2(n10809), .ZN(n10841) );
  INV_X1 U13344 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10832) );
  NAND2_X1 U13345 ( .A1(n10811), .A2(n10810), .ZN(n10814) );
  NAND2_X1 U13346 ( .A1(n10812), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10813) );
  NAND2_X1 U13347 ( .A1(n10814), .A2(n10813), .ZN(n13948) );
  INV_X1 U13348 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10815) );
  MUX2_X1 U13349 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10815), .S(n13950), .Z(
        n13949) );
  NAND2_X1 U13350 ( .A1(n13948), .A2(n13949), .ZN(n13961) );
  NAND2_X1 U13351 ( .A1(n13950), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n13960) );
  NAND2_X1 U13352 ( .A1(n13961), .A2(n13960), .ZN(n10818) );
  INV_X1 U13353 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10816) );
  MUX2_X1 U13354 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10816), .S(n13964), .Z(
        n10817) );
  NAND2_X1 U13355 ( .A1(n10818), .A2(n10817), .ZN(n13984) );
  NAND2_X1 U13356 ( .A1(n13964), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n13983) );
  NAND2_X1 U13357 ( .A1(n13984), .A2(n13983), .ZN(n10820) );
  INV_X1 U13358 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n13981) );
  MUX2_X1 U13359 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n13981), .S(n13980), .Z(
        n10819) );
  NAND2_X1 U13360 ( .A1(n10820), .A2(n10819), .ZN(n13998) );
  NAND2_X1 U13361 ( .A1(n13980), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n13997) );
  NAND2_X1 U13362 ( .A1(n13998), .A2(n13997), .ZN(n10823) );
  INV_X1 U13363 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10821) );
  MUX2_X1 U13364 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10821), .S(n13995), .Z(
        n10822) );
  NAND2_X1 U13365 ( .A1(n10823), .A2(n10822), .ZN(n14014) );
  NAND2_X1 U13366 ( .A1(n13995), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n14013) );
  NAND2_X1 U13367 ( .A1(n14014), .A2(n14013), .ZN(n10826) );
  INV_X1 U13368 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10824) );
  MUX2_X1 U13369 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10824), .S(n14011), .Z(
        n10825) );
  NAND2_X1 U13370 ( .A1(n10826), .A2(n10825), .ZN(n14029) );
  NAND2_X1 U13371 ( .A1(n14011), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n14028) );
  NAND2_X1 U13372 ( .A1(n14029), .A2(n14028), .ZN(n10829) );
  INV_X1 U13373 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10827) );
  MUX2_X1 U13374 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10827), .S(n14026), .Z(
        n10828) );
  NAND2_X1 U13375 ( .A1(n10829), .A2(n10828), .ZN(n14031) );
  NAND2_X1 U13376 ( .A1(n14026), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10830) );
  NAND2_X1 U13377 ( .A1(n14031), .A2(n10830), .ZN(n10836) );
  INV_X1 U13378 ( .A(n10836), .ZN(n10831) );
  NOR3_X1 U13379 ( .A1(n12583), .A2(n10832), .A3(n10831), .ZN(n10833) );
  AOI211_X1 U13380 ( .C1(n10834), .C2(n10841), .A(n15641), .B(n10833), .ZN(
        n10847) );
  INV_X1 U13381 ( .A(n10871), .ZN(n10854) );
  NAND2_X1 U13382 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n11762) );
  INV_X1 U13383 ( .A(n11762), .ZN(n10839) );
  MUX2_X1 U13384 ( .A(n10832), .B(P2_REG1_REG_9__SCAN_IN), .S(n10871), .Z(
        n10835) );
  NAND3_X1 U13385 ( .A1(n10836), .A2(n10832), .A3(n10854), .ZN(n10837) );
  AOI21_X1 U13386 ( .B1(n10873), .B2(n10837), .A(n12583), .ZN(n10838) );
  AOI211_X1 U13387 ( .C1(n15635), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n10839), .B(
        n10838), .ZN(n10846) );
  MUX2_X1 U13388 ( .A(n10796), .B(P2_REG2_REG_9__SCAN_IN), .S(n10871), .Z(
        n10840) );
  INV_X1 U13389 ( .A(n10866), .ZN(n10844) );
  INV_X1 U13390 ( .A(n10841), .ZN(n10842) );
  NOR3_X1 U13391 ( .A1(n10842), .A2(P2_REG2_REG_9__SCAN_IN), .A3(n10871), .ZN(
        n10843) );
  OAI21_X1 U13392 ( .B1(n10844), .B2(n10843), .A(n15644), .ZN(n10845) );
  OAI211_X1 U13393 ( .C1(n10847), .C2(n10854), .A(n10846), .B(n10845), .ZN(
        P2_U3223) );
  AND2_X1 U13394 ( .A1(n10984), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U13395 ( .A1(n10984), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U13396 ( .A1(n10984), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U13397 ( .A1(n10984), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U13398 ( .A1(n10984), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U13399 ( .A1(n10984), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U13400 ( .A1(n10984), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U13401 ( .A1(n10984), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U13402 ( .A1(n10984), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U13403 ( .A1(n10984), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U13404 ( .A1(n10984), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  INV_X1 U13405 ( .A(n13270), .ZN(n13293) );
  OAI222_X1 U13406 ( .A1(P3_U3151), .A2(n13293), .B1(n13715), .B2(n10849), 
        .C1(n13712), .C2(n10848), .ZN(P3_U3281) );
  AOI22_X1 U13407 ( .A1(n10993), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n10850), .ZN(n10851) );
  OAI21_X1 U13408 ( .B1(n10853), .B2(n15104), .A(n10851), .ZN(P1_U3346) );
  INV_X1 U13409 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13041) );
  NAND2_X1 U13410 ( .A1(n14690), .A2(P1_U4016), .ZN(n10852) );
  OAI21_X1 U13411 ( .B1(P1_U4016), .B2(n13041), .A(n10852), .ZN(P1_U3591) );
  INV_X1 U13412 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10855) );
  OAI222_X1 U13413 ( .A1(n14434), .A2(n10855), .B1(n10854), .B2(P2_U3088), 
        .C1(n14428), .C2(n10853), .ZN(P2_U3318) );
  INV_X1 U13414 ( .A(n12583), .ZN(n15639) );
  AOI22_X1 U13415 ( .A1(n15639), .A2(P2_REG1_REG_0__SCAN_IN), .B1(n15644), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n10860) );
  INV_X1 U13416 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10856) );
  NAND2_X1 U13417 ( .A1(n15644), .A2(n10856), .ZN(n10857) );
  OAI211_X1 U13418 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n12583), .A(n10857), .B(
        n14004), .ZN(n10858) );
  INV_X1 U13419 ( .A(n10858), .ZN(n10859) );
  MUX2_X1 U13420 ( .A(n10860), .B(n10859), .S(n15565), .Z(n10862) );
  AOI22_X1 U13421 ( .A1(n15635), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n10861) );
  NAND2_X1 U13422 ( .A1(n10862), .A2(n10861), .ZN(P2_U3214) );
  OAI222_X1 U13423 ( .A1(P3_U3151), .A2(n15146), .B1(n13715), .B2(n10864), 
        .C1(n13712), .C2(n10863), .ZN(P3_U3280) );
  OR2_X1 U13424 ( .A1(n10871), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10865) );
  NAND2_X1 U13425 ( .A1(n10866), .A2(n10865), .ZN(n10870) );
  INV_X1 U13426 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10867) );
  MUX2_X1 U13427 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n10867), .S(n10885), .Z(
        n10869) );
  INV_X1 U13428 ( .A(n12352), .ZN(n10868) );
  AOI211_X1 U13429 ( .C1(n10870), .C2(n10869), .A(n10868), .B(n12371), .ZN(
        n10881) );
  OR2_X1 U13430 ( .A1(n10871), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n10872) );
  NAND2_X1 U13431 ( .A1(n10873), .A2(n10872), .ZN(n10877) );
  INV_X1 U13432 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10874) );
  MUX2_X1 U13433 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n10874), .S(n10885), .Z(
        n10876) );
  INV_X1 U13434 ( .A(n14043), .ZN(n10875) );
  AOI211_X1 U13435 ( .C1(n10877), .C2(n10876), .A(n10875), .B(n12583), .ZN(
        n10880) );
  AND2_X1 U13436 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n11906) );
  AOI21_X1 U13437 ( .B1(n15635), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n11906), 
        .ZN(n10878) );
  OAI21_X1 U13438 ( .B1(n10885), .B2(n14004), .A(n10878), .ZN(n10879) );
  OR3_X1 U13439 ( .A1(n10881), .A2(n10880), .A3(n10879), .ZN(P2_U3224) );
  MUX2_X1 U13440 ( .A(n12317), .B(n14489), .S(P1_U4016), .Z(n10882) );
  INV_X1 U13441 ( .A(n10882), .ZN(P1_U3578) );
  INV_X1 U13442 ( .A(n10994), .ZN(n11047) );
  OAI222_X1 U13443 ( .A1(n15086), .A2(n10883), .B1(n15104), .B2(n10884), .C1(
        P1_U3086), .C2(n11047), .ZN(P1_U3345) );
  INV_X1 U13444 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10886) );
  OAI222_X1 U13445 ( .A1(n14434), .A2(n10886), .B1(n10885), .B2(P2_U3088), 
        .C1(n14428), .C2(n10884), .ZN(P2_U3317) );
  XNOR2_X1 U13446 ( .A(n10888), .B(n10887), .ZN(n11645) );
  AOI21_X1 U13447 ( .B1(n15711), .B2(n15710), .A(n11645), .ZN(n10893) );
  XNOR2_X1 U13448 ( .A(n10889), .B(n10890), .ZN(n10891) );
  AOI22_X1 U13449 ( .A1(n13906), .A2(n9686), .B1(n13945), .B2(n13907), .ZN(
        n11166) );
  OAI21_X1 U13450 ( .B1(n10891), .B2(n15668), .A(n11166), .ZN(n11642) );
  INV_X1 U13451 ( .A(n15281), .ZN(n15718) );
  OAI211_X1 U13452 ( .C1(n6915), .C2(n11836), .A(n14293), .B(n11562), .ZN(
        n11639) );
  OAI21_X1 U13453 ( .B1(n6915), .B2(n15718), .A(n11639), .ZN(n10892) );
  NOR3_X1 U13454 ( .A1(n10893), .A2(n11642), .A3(n10892), .ZN(n15705) );
  NOR2_X1 U13455 ( .A1(n15685), .A2(P2_U3088), .ZN(n10894) );
  AND2_X1 U13456 ( .A1(n10960), .A2(n10894), .ZN(n10895) );
  NAND2_X1 U13457 ( .A1(n15729), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10897) );
  OAI21_X1 U13458 ( .B1(n15705), .B2(n15729), .A(n10897), .ZN(P2_U3501) );
  MUX2_X1 U13459 ( .A(n7674), .B(P1_REG2_REG_2__SCAN_IN), .S(n14584), .Z(
        n10900) );
  MUX2_X1 U13460 ( .A(n11827), .B(P1_REG2_REG_1__SCAN_IN), .S(n10920), .Z(
        n14564) );
  AND2_X1 U13461 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10898) );
  NAND2_X1 U13462 ( .A1(n14564), .A2(n10898), .ZN(n14586) );
  OR2_X1 U13463 ( .A1(n10920), .A2(n11827), .ZN(n14585) );
  NAND2_X1 U13464 ( .A1(n14586), .A2(n14585), .ZN(n10899) );
  NAND2_X1 U13465 ( .A1(n10900), .A2(n10899), .ZN(n14593) );
  INV_X1 U13466 ( .A(n14584), .ZN(n14578) );
  NAND2_X1 U13467 ( .A1(n14578), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14592) );
  NAND2_X1 U13468 ( .A1(n14593), .A2(n14592), .ZN(n10903) );
  MUX2_X1 U13469 ( .A(n10901), .B(P1_REG2_REG_3__SCAN_IN), .S(n14598), .Z(
        n10902) );
  NAND2_X1 U13470 ( .A1(n10903), .A2(n10902), .ZN(n15456) );
  OR2_X1 U13471 ( .A1(n14598), .A2(n10901), .ZN(n15455) );
  NAND2_X1 U13472 ( .A1(n15456), .A2(n15455), .ZN(n10906) );
  INV_X1 U13473 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10904) );
  MUX2_X1 U13474 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10904), .S(n15459), .Z(
        n10905) );
  NAND2_X1 U13475 ( .A1(n10906), .A2(n10905), .ZN(n15458) );
  NAND2_X1 U13476 ( .A1(n15459), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n14616) );
  MUX2_X1 U13477 ( .A(n10907), .B(P1_REG2_REG_5__SCAN_IN), .S(n14610), .Z(
        n14617) );
  AOI21_X1 U13478 ( .B1(n15458), .B2(n14616), .A(n14617), .ZN(n14615) );
  NOR2_X1 U13479 ( .A1(n10908), .A2(n10907), .ZN(n11074) );
  INV_X1 U13480 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n12013) );
  MUX2_X1 U13481 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n12013), .S(n10923), .Z(
        n11073) );
  OAI21_X1 U13482 ( .B1(n14615), .B2(n11074), .A(n11073), .ZN(n14636) );
  NAND2_X1 U13483 ( .A1(n10923), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n14635) );
  INV_X1 U13484 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10909) );
  MUX2_X1 U13485 ( .A(n10909), .B(P1_REG2_REG_7__SCAN_IN), .S(n14627), .Z(
        n14634) );
  AOI21_X1 U13486 ( .B1(n14636), .B2(n14635), .A(n14634), .ZN(n14633) );
  NOR2_X1 U13487 ( .A1(n14623), .A2(n10909), .ZN(n10943) );
  MUX2_X1 U13488 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10910), .S(n10942), .Z(
        n10911) );
  OAI21_X1 U13489 ( .B1(n14633), .B2(n10943), .A(n10911), .ZN(n10946) );
  NAND2_X1 U13490 ( .A1(n10942), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10918) );
  INV_X1 U13491 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10912) );
  MUX2_X1 U13492 ( .A(n10912), .B(P1_REG2_REG_9__SCAN_IN), .S(n10993), .Z(
        n10917) );
  AOI21_X1 U13493 ( .B1(n10946), .B2(n10918), .A(n10917), .ZN(n10988) );
  NAND2_X1 U13494 ( .A1(n10914), .A2(n10913), .ZN(n15453) );
  INV_X1 U13495 ( .A(n15453), .ZN(n10916) );
  NOR2_X1 U13496 ( .A1(n10501), .A2(n6678), .ZN(n10915) );
  NAND2_X1 U13497 ( .A1(n10916), .A2(n10915), .ZN(n15481) );
  NAND3_X1 U13498 ( .A1(n10946), .A2(n10918), .A3(n10917), .ZN(n10919) );
  NAND2_X1 U13499 ( .A1(n15462), .A2(n10919), .ZN(n10936) );
  MUX2_X1 U13500 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9941), .S(n10920), .Z(
        n14566) );
  NAND2_X1 U13501 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14565) );
  OR2_X1 U13502 ( .A1(n14566), .A2(n14565), .ZN(n14581) );
  NAND2_X1 U13503 ( .A1(n7504), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n14580) );
  MUX2_X1 U13504 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10921), .S(n14584), .Z(
        n14582) );
  AOI21_X1 U13505 ( .B1(n14581), .B2(n14580), .A(n14582), .ZN(n14579) );
  NOR2_X1 U13506 ( .A1(n14584), .A2(n10921), .ZN(n14597) );
  MUX2_X1 U13507 ( .A(n15553), .B(P1_REG1_REG_3__SCAN_IN), .S(n14598), .Z(
        n10922) );
  OAI21_X1 U13508 ( .B1(n14579), .B2(n14597), .A(n10922), .ZN(n15466) );
  INV_X1 U13509 ( .A(n14598), .ZN(n14596) );
  NAND2_X1 U13510 ( .A1(n14596), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n15465) );
  MUX2_X1 U13511 ( .A(n10000), .B(P1_REG1_REG_4__SCAN_IN), .S(n15459), .Z(
        n15464) );
  AOI21_X1 U13512 ( .B1(n15466), .B2(n15465), .A(n15464), .ZN(n15463) );
  AOI21_X1 U13513 ( .B1(n15459), .B2(P1_REG1_REG_4__SCAN_IN), .A(n15463), .ZN(
        n14612) );
  MUX2_X1 U13514 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10018), .S(n14610), .Z(
        n14613) );
  NAND2_X1 U13515 ( .A1(n14612), .A2(n14613), .ZN(n14611) );
  OAI21_X1 U13516 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n14610), .A(n14611), .ZN(
        n11072) );
  MUX2_X1 U13517 ( .A(n10037), .B(P1_REG1_REG_6__SCAN_IN), .S(n10923), .Z(
        n11071) );
  NOR2_X1 U13518 ( .A1(n11072), .A2(n11071), .ZN(n14632) );
  NOR2_X1 U13519 ( .A1(n11081), .A2(n10037), .ZN(n14626) );
  MUX2_X1 U13520 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10924), .S(n14627), .Z(
        n10925) );
  OAI21_X1 U13521 ( .B1(n14632), .B2(n14626), .A(n10925), .ZN(n14630) );
  OAI21_X1 U13522 ( .B1(n10924), .B2(n14623), .A(n14630), .ZN(n10938) );
  MUX2_X1 U13523 ( .A(n10926), .B(P1_REG1_REG_8__SCAN_IN), .S(n10942), .Z(
        n10939) );
  NOR2_X1 U13524 ( .A1(n10938), .A2(n10939), .ZN(n10937) );
  NOR2_X1 U13525 ( .A1(n10942), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10927) );
  MUX2_X1 U13526 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10084), .S(n10993), .Z(
        n10928) );
  OAI21_X1 U13527 ( .B1(n10937), .B2(n10927), .A(n10928), .ZN(n10992) );
  INV_X1 U13528 ( .A(n10992), .ZN(n10930) );
  NOR3_X1 U13529 ( .A1(n10937), .A2(n10928), .A3(n10927), .ZN(n10929) );
  NOR2_X2 U13530 ( .A1(n15453), .A2(n15443), .ZN(n15469) );
  OAI21_X1 U13531 ( .B1(n10930), .B2(n10929), .A(n15469), .ZN(n10935) );
  NOR2_X1 U13532 ( .A1(n15453), .A2(n10931), .ZN(n15460) );
  INV_X1 U13533 ( .A(n15450), .ZN(n15489) );
  INV_X1 U13534 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10932) );
  NAND2_X1 U13535 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n12549) );
  OAI21_X1 U13536 ( .B1(n15489), .B2(n10932), .A(n12549), .ZN(n10933) );
  AOI21_X1 U13537 ( .B1(n10993), .B2(n15460), .A(n10933), .ZN(n10934) );
  OAI211_X1 U13538 ( .C1(n10988), .C2(n10936), .A(n10935), .B(n10934), .ZN(
        P1_U3252) );
  AOI21_X1 U13539 ( .B1(n10939), .B2(n10938), .A(n10937), .ZN(n10950) );
  INV_X1 U13540 ( .A(n15469), .ZN(n15483) );
  INV_X1 U13541 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10940) );
  NAND2_X1 U13542 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n12237) );
  OAI21_X1 U13543 ( .B1(n15489), .B2(n10940), .A(n12237), .ZN(n10941) );
  AOI21_X1 U13544 ( .B1(n10942), .B2(n15460), .A(n10941), .ZN(n10949) );
  MUX2_X1 U13545 ( .A(n10910), .B(P1_REG2_REG_8__SCAN_IN), .S(n10942), .Z(
        n10945) );
  INV_X1 U13546 ( .A(n10943), .ZN(n10944) );
  NAND2_X1 U13547 ( .A1(n10945), .A2(n10944), .ZN(n10947) );
  OAI211_X1 U13548 ( .C1(n14633), .C2(n10947), .A(n15462), .B(n10946), .ZN(
        n10948) );
  OAI211_X1 U13549 ( .C1(n10950), .C2(n15483), .A(n10949), .B(n10948), .ZN(
        P1_U3251) );
  INV_X1 U13550 ( .A(n15688), .ZN(n10951) );
  NAND2_X1 U13551 ( .A1(n10952), .A2(n10951), .ZN(n11554) );
  INV_X1 U13552 ( .A(n15685), .ZN(n10953) );
  NAND2_X1 U13553 ( .A1(n15689), .A2(n10953), .ZN(n10954) );
  NOR2_X1 U13554 ( .A1(n15281), .A2(n10955), .ZN(n10956) );
  NAND2_X2 U13555 ( .A1(n10968), .A2(n10956), .ZN(n13916) );
  INV_X1 U13556 ( .A(n13916), .ZN(n13880) );
  NAND2_X1 U13557 ( .A1(n7043), .A2(n8434), .ZN(n10958) );
  OR2_X1 U13558 ( .A1(n11841), .A2(n14078), .ZN(n11135) );
  AND2_X1 U13559 ( .A1(n10958), .A2(n11135), .ZN(n10959) );
  XNOR2_X1 U13560 ( .A(n11110), .B(n9178), .ZN(n11106) );
  NAND2_X1 U13561 ( .A1(n9686), .A2(n13804), .ZN(n11107) );
  OAI21_X1 U13562 ( .B1(n11554), .B2(n15685), .A(n10964), .ZN(n10961) );
  NAND2_X1 U13563 ( .A1(n10961), .A2(n10960), .ZN(n11123) );
  OR2_X1 U13564 ( .A1(n11123), .A2(P2_U3088), .ZN(n11168) );
  AOI22_X1 U13565 ( .A1(n13880), .A2(n10962), .B1(n11168), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n10972) );
  AND2_X1 U13566 ( .A1(n15690), .A2(n10963), .ZN(n11560) );
  NAND2_X1 U13567 ( .A1(n10968), .A2(n11560), .ZN(n10966) );
  INV_X1 U13568 ( .A(n10964), .ZN(n10965) );
  NAND2_X2 U13569 ( .A1(n15689), .A2(n10965), .ZN(n15676) );
  NAND2_X1 U13570 ( .A1(n13946), .A2(n13907), .ZN(n10970) );
  NAND2_X1 U13571 ( .A1(n13947), .A2(n13906), .ZN(n10969) );
  NAND2_X1 U13572 ( .A1(n10970), .A2(n10969), .ZN(n11834) );
  AOI22_X1 U13573 ( .A1(n9178), .A2(n13914), .B1(n13910), .B2(n11834), .ZN(
        n10971) );
  NAND2_X1 U13574 ( .A1(n10972), .A2(n10971), .ZN(P2_U3194) );
  INV_X1 U13575 ( .A(n10973), .ZN(n10974) );
  OAI222_X1 U13576 ( .A1(P3_U3151), .A2(n13333), .B1(n13709), .B2(n10975), 
        .C1(n13712), .C2(n10974), .ZN(P3_U3279) );
  OAI222_X1 U13577 ( .A1(P3_U3151), .A2(n13361), .B1(n13715), .B2(n10977), 
        .C1(n13712), .C2(n10976), .ZN(P3_U3278) );
  INV_X1 U13578 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10979) );
  INV_X1 U13579 ( .A(n10978), .ZN(n10980) );
  INV_X1 U13580 ( .A(n14648), .ZN(n10995) );
  OAI222_X1 U13581 ( .A1(n15086), .A2(n10979), .B1(n15104), .B2(n10980), .C1(
        P1_U3086), .C2(n10995), .ZN(P1_U3344) );
  INV_X1 U13582 ( .A(n14040), .ZN(n12353) );
  OAI222_X1 U13583 ( .A1(n14434), .A2(n10981), .B1(n14428), .B2(n10980), .C1(
        P2_U3088), .C2(n12353), .ZN(P2_U3316) );
  NAND2_X1 U13584 ( .A1(n13518), .A2(P3_U3897), .ZN(n10982) );
  OAI21_X1 U13585 ( .B1(P3_U3897), .B2(n10983), .A(n10982), .ZN(P3_U3510) );
  INV_X1 U13586 ( .A(n10985), .ZN(n10986) );
  AOI22_X1 U13587 ( .A1(n10984), .A2(n10987), .B1(n13685), .B2(n10986), .ZN(
        P3_U3377) );
  MUX2_X1 U13588 ( .A(n12538), .B(P1_REG2_REG_12__SCAN_IN), .S(n11000), .Z(
        n10991) );
  AOI21_X1 U13589 ( .B1(n10993), .B2(P1_REG2_REG_9__SCAN_IN), .A(n10988), .ZN(
        n11044) );
  MUX2_X1 U13590 ( .A(n12479), .B(P1_REG2_REG_10__SCAN_IN), .S(n10994), .Z(
        n11043) );
  NOR2_X1 U13591 ( .A1(n11044), .A2(n11043), .ZN(n14651) );
  NOR2_X1 U13592 ( .A1(n11047), .A2(n12479), .ZN(n14650) );
  MUX2_X1 U13593 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n10989), .S(n14648), .Z(
        n14649) );
  OAI21_X1 U13594 ( .B1(n14651), .B2(n14650), .A(n14649), .ZN(n14653) );
  OAI21_X1 U13595 ( .B1(n10995), .B2(n10989), .A(n14653), .ZN(n10990) );
  NOR2_X1 U13596 ( .A1(n10990), .A2(n10991), .ZN(n11083) );
  AOI21_X1 U13597 ( .B1(n10991), .B2(n10990), .A(n11083), .ZN(n11005) );
  OAI21_X1 U13598 ( .B1(n10993), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10992), .ZN(
        n11042) );
  MUX2_X1 U13599 ( .A(n10105), .B(P1_REG1_REG_10__SCAN_IN), .S(n10994), .Z(
        n11041) );
  NOR2_X1 U13600 ( .A1(n11042), .A2(n11041), .ZN(n11040) );
  AOI21_X1 U13601 ( .B1(n10994), .B2(P1_REG1_REG_10__SCAN_IN), .A(n11040), 
        .ZN(n14643) );
  MUX2_X1 U13602 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10118), .S(n14648), .Z(
        n14644) );
  NAND2_X1 U13603 ( .A1(n14643), .A2(n14644), .ZN(n14642) );
  NAND2_X1 U13604 ( .A1(n10995), .A2(n10118), .ZN(n10997) );
  MUX2_X1 U13605 ( .A(n10996), .B(P1_REG1_REG_12__SCAN_IN), .S(n11000), .Z(
        n10998) );
  AOI21_X1 U13606 ( .B1(n14642), .B2(n10997), .A(n10998), .ZN(n11082) );
  AND3_X1 U13607 ( .A1(n14642), .A2(n10998), .A3(n10997), .ZN(n10999) );
  OAI21_X1 U13608 ( .B1(n11082), .B2(n10999), .A(n15469), .ZN(n11004) );
  NOR2_X1 U13609 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n12683), .ZN(n11002) );
  INV_X1 U13610 ( .A(n11000), .ZN(n11180) );
  NOR2_X1 U13611 ( .A1(n15485), .A2(n11180), .ZN(n11001) );
  AOI211_X1 U13612 ( .C1(n15450), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n11002), 
        .B(n11001), .ZN(n11003) );
  OAI211_X1 U13613 ( .C1(n11005), .C2(n15481), .A(n11004), .B(n11003), .ZN(
        P1_U3255) );
  INV_X1 U13614 ( .A(n15744), .ZN(n11149) );
  OAI21_X1 U13615 ( .B1(n11007), .B2(P3_REG1_REG_1__SCAN_IN), .A(n11006), .ZN(
        n11021) );
  NAND2_X1 U13616 ( .A1(n15732), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n11013) );
  NAND2_X1 U13617 ( .A1(n11009), .A2(n11239), .ZN(n11010) );
  NAND2_X1 U13618 ( .A1(n11061), .A2(n11010), .ZN(n11011) );
  NAND2_X1 U13619 ( .A1(n13395), .A2(n11011), .ZN(n11012) );
  OAI211_X1 U13620 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n11014), .A(n11013), .B(
        n11012), .ZN(n11020) );
  NAND2_X1 U13621 ( .A1(n11016), .A2(n11015), .ZN(n11017) );
  AOI21_X1 U13622 ( .B1(n11018), .B2(n11017), .A(n15752), .ZN(n11019) );
  AOI211_X1 U13623 ( .C1(n11149), .C2(n11021), .A(n11020), .B(n11019), .ZN(
        n11022) );
  OAI21_X1 U13624 ( .B1(n11023), .B2(n15738), .A(n11022), .ZN(P3_U3183) );
  AND2_X1 U13625 ( .A1(n10984), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U13626 ( .A1(n10984), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U13627 ( .A1(n10984), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U13628 ( .A1(n10984), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U13629 ( .A1(n10984), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U13630 ( .A1(n10984), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U13631 ( .A1(n10984), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U13632 ( .A1(n10984), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U13633 ( .A1(n10984), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U13634 ( .A1(n10984), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U13635 ( .A1(n10984), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U13636 ( .A1(n10984), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U13637 ( .A1(n10984), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U13638 ( .A1(n10984), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U13639 ( .A1(n10984), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U13640 ( .A1(n10984), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U13641 ( .A1(n10984), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U13642 ( .A1(n10984), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U13643 ( .A1(n10984), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  INV_X1 U13644 ( .A(n15752), .ZN(n12430) );
  OAI21_X1 U13645 ( .B1(n11024), .B2(P3_REG2_REG_3__SCAN_IN), .A(n11142), .ZN(
        n11033) );
  NAND2_X1 U13646 ( .A1(n11025), .A2(n10646), .ZN(n11026) );
  AND2_X1 U13647 ( .A1(n11148), .A2(n11026), .ZN(n11029) );
  NOR2_X1 U13648 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11740), .ZN(n11732) );
  INV_X1 U13649 ( .A(n11732), .ZN(n11028) );
  NAND2_X1 U13650 ( .A1(n15732), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n11027) );
  OAI211_X1 U13651 ( .C1(n15744), .C2(n11029), .A(n11028), .B(n11027), .ZN(
        n11032) );
  NOR2_X1 U13652 ( .A1(n15738), .A2(n11030), .ZN(n11031) );
  AOI211_X1 U13653 ( .C1(n12430), .C2(n11033), .A(n11032), .B(n11031), .ZN(
        n11039) );
  INV_X1 U13654 ( .A(n11157), .ZN(n11037) );
  NOR3_X1 U13655 ( .A1(n11063), .A2(n11035), .A3(n11034), .ZN(n11036) );
  OAI21_X1 U13656 ( .B1(n11037), .B2(n11036), .A(n13395), .ZN(n11038) );
  NAND2_X1 U13657 ( .A1(n11039), .A2(n11038), .ZN(P3_U3185) );
  AOI211_X1 U13658 ( .C1(n11042), .C2(n11041), .A(n15483), .B(n11040), .ZN(
        n11050) );
  NAND2_X1 U13659 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n15319)
         );
  AOI211_X1 U13660 ( .C1(n11044), .C2(n11043), .A(n15481), .B(n14651), .ZN(
        n11045) );
  INV_X1 U13661 ( .A(n11045), .ZN(n11046) );
  NAND2_X1 U13662 ( .A1(n15319), .A2(n11046), .ZN(n11049) );
  OAI22_X1 U13663 ( .A1(n15485), .A2(n11047), .B1(n15489), .B2(n9229), .ZN(
        n11048) );
  OR3_X1 U13664 ( .A1(n11050), .A2(n11049), .A3(n11048), .ZN(P1_U3253) );
  OAI21_X1 U13665 ( .B1(n11053), .B2(n11052), .A(n11051), .ZN(n11054) );
  NAND2_X1 U13666 ( .A1(n12430), .A2(n11054), .ZN(n11067) );
  OAI21_X1 U13667 ( .B1(n11057), .B2(n11056), .A(n11055), .ZN(n11058) );
  NAND2_X1 U13668 ( .A1(n11149), .A2(n11058), .ZN(n11066) );
  AOI22_X1 U13669 ( .A1(n15732), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n11065) );
  AND3_X1 U13670 ( .A1(n11061), .A2(n11060), .A3(n11059), .ZN(n11062) );
  OAI21_X1 U13671 ( .B1(n11063), .B2(n11062), .A(n13395), .ZN(n11064) );
  NAND4_X1 U13672 ( .A1(n11067), .A2(n11066), .A3(n11065), .A4(n11064), .ZN(
        n11068) );
  AOI21_X1 U13673 ( .B1(n11069), .B2(n13349), .A(n11068), .ZN(n11070) );
  INV_X1 U13674 ( .A(n11070), .ZN(P3_U3184) );
  AOI211_X1 U13675 ( .C1(n11072), .C2(n11071), .A(n14632), .B(n15483), .ZN(
        n11078) );
  INV_X1 U13676 ( .A(n14636), .ZN(n11076) );
  NOR3_X1 U13677 ( .A1(n14615), .A2(n11074), .A3(n11073), .ZN(n11075) );
  NOR3_X1 U13678 ( .A1(n15481), .A2(n11076), .A3(n11075), .ZN(n11077) );
  NOR2_X1 U13679 ( .A1(n11078), .A2(n11077), .ZN(n11080) );
  AND2_X1 U13680 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n11950) );
  AOI21_X1 U13681 ( .B1(n15450), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n11950), .ZN(
        n11079) );
  OAI211_X1 U13682 ( .C1(n11081), .C2(n15485), .A(n11080), .B(n11079), .ZN(
        P1_U3249) );
  MUX2_X1 U13683 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10152), .S(n11257), .Z(
        n11184) );
  AOI21_X1 U13684 ( .B1(n10996), .B2(n11180), .A(n11082), .ZN(n11186) );
  XOR2_X1 U13685 ( .A(n11184), .B(n11186), .Z(n11091) );
  NOR2_X1 U13686 ( .A1(n15485), .A2(n11257), .ZN(n11089) );
  NAND2_X1 U13687 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n15343)
         );
  AOI21_X1 U13688 ( .B1(n12538), .B2(n11180), .A(n11083), .ZN(n11086) );
  MUX2_X1 U13689 ( .A(n11084), .B(P1_REG2_REG_13__SCAN_IN), .S(n11257), .Z(
        n11085) );
  NAND2_X1 U13690 ( .A1(n11086), .A2(n11085), .ZN(n11190) );
  OAI211_X1 U13691 ( .C1(n11086), .C2(n11085), .A(n11190), .B(n15462), .ZN(
        n11087) );
  NAND2_X1 U13692 ( .A1(n15343), .A2(n11087), .ZN(n11088) );
  AOI211_X1 U13693 ( .C1(n15450), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n11089), 
        .B(n11088), .ZN(n11090) );
  OAI21_X1 U13694 ( .B1(n11091), .B2(n15483), .A(n11090), .ZN(P1_U3256) );
  XNOR2_X1 U13695 ( .A(n11092), .B(n11093), .ZN(n15658) );
  XNOR2_X1 U13696 ( .A(n11094), .B(n11093), .ZN(n11097) );
  NAND2_X1 U13697 ( .A1(n13943), .A2(n13907), .ZN(n11096) );
  NAND2_X1 U13698 ( .A1(n13945), .A2(n13906), .ZN(n11095) );
  NAND2_X1 U13699 ( .A1(n11096), .A2(n11095), .ZN(n11124) );
  AOI21_X1 U13700 ( .B1(n11097), .B2(n15256), .A(n11124), .ZN(n15657) );
  OAI211_X1 U13701 ( .C1(n15662), .C2(n11563), .A(n14293), .B(n11326), .ZN(
        n15653) );
  OAI211_X1 U13702 ( .C1(n15285), .C2(n15658), .A(n15657), .B(n15653), .ZN(
        n11102) );
  NAND2_X1 U13703 ( .A1(n15731), .A2(n15281), .ZN(n14351) );
  OAI22_X1 U13704 ( .A1(n14351), .A2(n15662), .B1(n15731), .B2(n10816), .ZN(
        n11098) );
  AOI21_X1 U13705 ( .B1(n11102), .B2(n15731), .A(n11098), .ZN(n11099) );
  INV_X1 U13706 ( .A(n11099), .ZN(P2_U3503) );
  INV_X1 U13707 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n11100) );
  OAI22_X1 U13708 ( .A1(n14401), .A2(n15662), .B1(n15724), .B2(n11100), .ZN(
        n11101) );
  AOI21_X1 U13709 ( .B1(n11102), .B2(n15724), .A(n11101), .ZN(n11103) );
  INV_X1 U13710 ( .A(n11103), .ZN(P2_U3442) );
  INV_X1 U13711 ( .A(n11104), .ZN(n11179) );
  AOI22_X1 U13712 ( .A1(n15586), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n14421), .ZN(n11105) );
  OAI21_X1 U13713 ( .B1(n11179), .B2(n14428), .A(n11105), .ZN(P2_U3315) );
  XNOR2_X1 U13714 ( .A(n11125), .B(n13806), .ZN(n11227) );
  NAND2_X1 U13715 ( .A1(n13944), .A2(n13804), .ZN(n11217) );
  XNOR2_X1 U13716 ( .A(n11227), .B(n11217), .ZN(n11128) );
  INV_X1 U13717 ( .A(n11106), .ZN(n11169) );
  NAND2_X1 U13718 ( .A1(n11169), .A2(n11107), .ZN(n11108) );
  NAND2_X1 U13719 ( .A1(n11172), .A2(n11108), .ZN(n11111) );
  XNOR2_X1 U13720 ( .A(n11110), .B(n11109), .ZN(n11112) );
  NAND2_X1 U13721 ( .A1(n13946), .A2(n13804), .ZN(n11113) );
  XNOR2_X1 U13722 ( .A(n11112), .B(n11113), .ZN(n11171) );
  INV_X1 U13723 ( .A(n11112), .ZN(n11114) );
  NAND2_X1 U13724 ( .A1(n11114), .A2(n11113), .ZN(n11115) );
  XNOR2_X1 U13725 ( .A(n13783), .B(n13806), .ZN(n11116) );
  AND2_X1 U13726 ( .A1(n13945), .A2(n13804), .ZN(n11117) );
  NAND2_X1 U13727 ( .A1(n11116), .A2(n11117), .ZN(n11121) );
  INV_X1 U13728 ( .A(n11116), .ZN(n11129) );
  INV_X1 U13729 ( .A(n11117), .ZN(n11118) );
  NAND2_X1 U13730 ( .A1(n11129), .A2(n11118), .ZN(n11119) );
  NAND2_X1 U13731 ( .A1(n11121), .A2(n11119), .ZN(n13778) );
  AND2_X1 U13732 ( .A1(n11128), .A2(n11121), .ZN(n11122) );
  NAND2_X1 U13733 ( .A1(n13780), .A2(n11122), .ZN(n11220) );
  OAI21_X1 U13734 ( .B1(n11128), .B2(n13780), .A(n11220), .ZN(n11133) );
  AND2_X1 U13735 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n13963) );
  AOI21_X1 U13736 ( .B1(n13910), .B2(n11124), .A(n13963), .ZN(n11127) );
  NAND2_X1 U13737 ( .A1(n13914), .A2(n11125), .ZN(n11126) );
  OAI211_X1 U13738 ( .C1(n13912), .C2(n15661), .A(n11127), .B(n11126), .ZN(
        n11132) );
  OR2_X1 U13739 ( .A1(n13916), .A2(n14078), .ZN(n13844) );
  NOR4_X1 U13740 ( .A1(n13844), .A2(n11130), .A3(n11129), .A4(n11128), .ZN(
        n11131) );
  AOI211_X1 U13741 ( .C1(n13880), .C2(n11133), .A(n11132), .B(n11131), .ZN(
        n11134) );
  INV_X1 U13742 ( .A(n11134), .ZN(P2_U3202) );
  INV_X1 U13743 ( .A(n11135), .ZN(n11139) );
  INV_X1 U13744 ( .A(n13844), .ZN(n13877) );
  AOI22_X1 U13745 ( .A1(n13877), .A2(n13947), .B1(n13880), .B2(n15691), .ZN(
        n11138) );
  NAND2_X1 U13746 ( .A1(n9686), .A2(n13907), .ZN(n15669) );
  OAI22_X1 U13747 ( .A1(n13901), .A2(n8434), .B1(n13884), .B2(n15669), .ZN(
        n11136) );
  AOI21_X1 U13748 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n11168), .A(n11136), .ZN(
        n11137) );
  OAI21_X1 U13749 ( .B1(n11139), .B2(n11138), .A(n11137), .ZN(P2_U3204) );
  AND3_X1 U13750 ( .A1(n11142), .A2(n11141), .A3(n11140), .ZN(n11143) );
  OAI21_X1 U13751 ( .B1(n11144), .B2(n11143), .A(n12430), .ZN(n11154) );
  INV_X1 U13752 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n11145) );
  NOR2_X1 U13753 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11145), .ZN(n11797) );
  AOI21_X1 U13754 ( .B1(n15732), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n11797), .ZN(
        n11153) );
  AND3_X1 U13755 ( .A1(n11148), .A2(n11147), .A3(n11146), .ZN(n11150) );
  OAI21_X1 U13756 ( .B1(n11151), .B2(n11150), .A(n11149), .ZN(n11152) );
  NAND3_X1 U13757 ( .A1(n11154), .A2(n11153), .A3(n11152), .ZN(n11161) );
  INV_X1 U13758 ( .A(n11212), .ZN(n11159) );
  NAND3_X1 U13759 ( .A1(n11157), .A2(n11156), .A3(n11155), .ZN(n11158) );
  AOI21_X1 U13760 ( .B1(n11159), .B2(n11158), .A(n15746), .ZN(n11160) );
  AOI211_X1 U13761 ( .C1(n13349), .C2(n11162), .A(n11161), .B(n11160), .ZN(
        n11163) );
  INV_X1 U13762 ( .A(n11163), .ZN(P3_U3186) );
  NAND2_X1 U13763 ( .A1(n13466), .A2(P3_U3897), .ZN(n11164) );
  OAI21_X1 U13764 ( .B1(P3_U3897), .B2(n11165), .A(n11164), .ZN(P3_U3514) );
  OAI22_X1 U13765 ( .A1(n6915), .A2(n13901), .B1(n13884), .B2(n11166), .ZN(
        n11167) );
  AOI21_X1 U13766 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n11168), .A(n11167), .ZN(
        n11176) );
  INV_X1 U13767 ( .A(n9686), .ZN(n11170) );
  OAI22_X1 U13768 ( .A1(n13844), .A2(n11170), .B1(n11169), .B2(n13916), .ZN(
        n11174) );
  INV_X1 U13769 ( .A(n11171), .ZN(n11173) );
  NAND3_X1 U13770 ( .A1(n11174), .A2(n11173), .A3(n11172), .ZN(n11175) );
  OAI211_X1 U13771 ( .C1(n13916), .C2(n11177), .A(n11176), .B(n11175), .ZN(
        P2_U3209) );
  OAI222_X1 U13772 ( .A1(P1_U3086), .A2(n11180), .B1(n15104), .B2(n11179), 
        .C1(n11178), .C2(n15086), .ZN(P1_U3343) );
  INV_X1 U13773 ( .A(n11181), .ZN(n11182) );
  OAI222_X1 U13774 ( .A1(P3_U3151), .A2(n13380), .B1(n13709), .B2(n11183), 
        .C1(n13712), .C2(n11182), .ZN(P3_U3277) );
  INV_X1 U13775 ( .A(n11195), .ZN(n12217) );
  AOI22_X1 U13776 ( .A1(n11195), .A2(n10176), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n12217), .ZN(n11189) );
  INV_X1 U13777 ( .A(n11184), .ZN(n11185) );
  NAND2_X1 U13778 ( .A1(n11186), .A2(n11185), .ZN(n11187) );
  OAI21_X1 U13779 ( .B1(n11257), .B2(n10152), .A(n11187), .ZN(n11188) );
  NOR2_X1 U13780 ( .A1(n11189), .A2(n11188), .ZN(n12216) );
  AOI21_X1 U13781 ( .B1(n11189), .B2(n11188), .A(n12216), .ZN(n11198) );
  OAI21_X1 U13782 ( .B1(n11257), .B2(n11084), .A(n11190), .ZN(n11192) );
  MUX2_X1 U13783 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n12613), .S(n11195), .Z(
        n11191) );
  NAND2_X1 U13784 ( .A1(n11191), .A2(n11192), .ZN(n12209) );
  OAI211_X1 U13785 ( .C1(n11192), .C2(n11191), .A(n15462), .B(n12209), .ZN(
        n11197) );
  NAND2_X1 U13786 ( .A1(n15450), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n11193) );
  NAND2_X1 U13787 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n15309)
         );
  NAND2_X1 U13788 ( .A1(n11193), .A2(n15309), .ZN(n11194) );
  AOI21_X1 U13789 ( .B1(n11195), .B2(n15460), .A(n11194), .ZN(n11196) );
  OAI211_X1 U13790 ( .C1(n11198), .C2(n15483), .A(n11197), .B(n11196), .ZN(
        P1_U3257) );
  AOI21_X1 U13791 ( .B1(n11201), .B2(n11200), .A(n11199), .ZN(n11207) );
  NOR2_X1 U13792 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7924), .ZN(n11977) );
  AOI21_X1 U13793 ( .B1(n11203), .B2(n10657), .A(n11202), .ZN(n11204) );
  NOR2_X1 U13794 ( .A1(n11204), .A2(n15744), .ZN(n11205) );
  AOI211_X1 U13795 ( .C1(n15732), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n11977), .B(
        n11205), .ZN(n11206) );
  OAI21_X1 U13796 ( .B1(n11207), .B2(n15752), .A(n11206), .ZN(n11208) );
  AOI21_X1 U13797 ( .B1(n11209), .B2(n13349), .A(n11208), .ZN(n11216) );
  INV_X1 U13798 ( .A(n11298), .ZN(n11214) );
  NOR3_X1 U13799 ( .A1(n11212), .A2(n11211), .A3(n11210), .ZN(n11213) );
  OAI21_X1 U13800 ( .B1(n11214), .B2(n11213), .A(n13395), .ZN(n11215) );
  NAND2_X1 U13801 ( .A1(n11216), .A2(n11215), .ZN(P3_U3187) );
  INV_X1 U13802 ( .A(n11227), .ZN(n11218) );
  NAND2_X1 U13803 ( .A1(n11218), .A2(n11217), .ZN(n11219) );
  NAND2_X1 U13804 ( .A1(n11220), .A2(n11219), .ZN(n11221) );
  XNOR2_X1 U13805 ( .A(n11590), .B(n13806), .ZN(n11336) );
  NAND2_X1 U13806 ( .A1(n13943), .A2(n13804), .ZN(n11337) );
  XNOR2_X1 U13807 ( .A(n11336), .B(n11337), .ZN(n11228) );
  INV_X1 U13808 ( .A(n13912), .ZN(n13886) );
  INV_X1 U13809 ( .A(n11591), .ZN(n11233) );
  NAND2_X1 U13810 ( .A1(n13914), .A2(n11590), .ZN(n11226) );
  NAND2_X1 U13811 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n13974) );
  NAND2_X1 U13812 ( .A1(n13942), .A2(n13907), .ZN(n11223) );
  NAND2_X1 U13813 ( .A1(n13944), .A2(n13906), .ZN(n11222) );
  AND2_X1 U13814 ( .A1(n11223), .A2(n11222), .ZN(n11329) );
  INV_X1 U13815 ( .A(n11329), .ZN(n11224) );
  NAND2_X1 U13816 ( .A1(n13910), .A2(n11224), .ZN(n11225) );
  NAND3_X1 U13817 ( .A1(n11226), .A2(n13974), .A3(n11225), .ZN(n11232) );
  AOI22_X1 U13818 ( .A1(n13877), .A2(n13944), .B1(n13880), .B2(n11227), .ZN(
        n11230) );
  INV_X1 U13819 ( .A(n11220), .ZN(n11229) );
  NOR3_X1 U13820 ( .A1(n11230), .A2(n11229), .A3(n11228), .ZN(n11231) );
  AOI211_X1 U13821 ( .C1(n13886), .C2(n11233), .A(n11232), .B(n11231), .ZN(
        n11234) );
  OAI21_X1 U13822 ( .B1(n11340), .B2(n13916), .A(n11234), .ZN(P2_U3199) );
  NAND2_X1 U13823 ( .A1(n15807), .A2(n11475), .ZN(n13099) );
  AND2_X1 U13824 ( .A1(n15803), .A2(n13099), .ZN(n13061) );
  NAND2_X1 U13825 ( .A1(n11235), .A2(n15815), .ZN(n11236) );
  OAI22_X1 U13826 ( .A1(n13061), .A2(n11236), .B1(n15790), .B2(n15787), .ZN(
        n11473) );
  NOR2_X1 U13827 ( .A1(n15854), .A2(n10639), .ZN(n11237) );
  AOI21_X1 U13828 ( .B1(n15854), .B2(n11473), .A(n11237), .ZN(n11238) );
  OAI21_X1 U13829 ( .B1(n11475), .B2(n13626), .A(n11238), .ZN(P3_U3459) );
  INV_X1 U13830 ( .A(n11239), .ZN(n11251) );
  NAND3_X1 U13831 ( .A1(n15746), .A2(n15752), .A3(n15744), .ZN(n11250) );
  NAND2_X1 U13832 ( .A1(n12430), .A2(n11240), .ZN(n11244) );
  NOR2_X1 U13833 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11241), .ZN(n11242) );
  AOI21_X1 U13834 ( .B1(n15732), .B2(P3_ADDR_REG_0__SCAN_IN), .A(n11242), .ZN(
        n11243) );
  OAI211_X1 U13835 ( .C1(n11245), .C2(n15744), .A(n11244), .B(n11243), .ZN(
        n11249) );
  NOR2_X1 U13836 ( .A1(n15746), .A2(n11246), .ZN(n11247) );
  MUX2_X1 U13837 ( .A(n11247), .B(n13349), .S(P3_IR_REG_0__SCAN_IN), .Z(n11248) );
  AOI211_X1 U13838 ( .C1(n11251), .C2(n11250), .A(n11249), .B(n11248), .ZN(
        n11252) );
  INV_X1 U13839 ( .A(n11252), .ZN(P3_U3182) );
  INV_X1 U13840 ( .A(n11253), .ZN(n11255) );
  OAI222_X1 U13841 ( .A1(n13712), .A2(n11255), .B1(n13709), .B2(n11254), .C1(
        P3_U3151), .C2(n13393), .ZN(P3_U3276) );
  INV_X1 U13842 ( .A(n11256), .ZN(n11271) );
  OAI222_X1 U13843 ( .A1(n15086), .A2(n11258), .B1(P1_U3086), .B2(n11257), 
        .C1(n11271), .C2(n15104), .ZN(P1_U3342) );
  INV_X1 U13844 ( .A(n15805), .ZN(n11264) );
  INV_X1 U13845 ( .A(n11259), .ZN(n15804) );
  NOR3_X1 U13846 ( .A1(n15804), .A2(n12862), .A3(n11260), .ZN(n11262) );
  AOI211_X1 U13847 ( .C1(n11264), .C2(n11263), .A(n11262), .B(n11261), .ZN(
        n11270) );
  INV_X1 U13848 ( .A(n13028), .ZN(n13014) );
  OAI22_X1 U13849 ( .A1(n13016), .A2(n7377), .B1(n13035), .B2(n15816), .ZN(
        n11265) );
  AOI21_X1 U13850 ( .B1(n13014), .B2(n15807), .A(n11265), .ZN(n11269) );
  OR2_X1 U13851 ( .A1(n11267), .A2(n11266), .ZN(n11500) );
  NAND2_X1 U13852 ( .A1(n11500), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n11268) );
  OAI211_X1 U13853 ( .C1(n11270), .C2(n13008), .A(n11269), .B(n11268), .ZN(
        P3_U3162) );
  INV_X1 U13854 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n11272) );
  INV_X1 U13855 ( .A(n15594), .ZN(n12356) );
  OAI222_X1 U13856 ( .A1(n14434), .A2(n11272), .B1(n12356), .B2(P2_U3088), 
        .C1(n14428), .C2(n11271), .ZN(P2_U3314) );
  NAND2_X1 U13857 ( .A1(n11500), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n11274) );
  AOI22_X1 U13858 ( .A1(n13026), .A2(n11400), .B1(n13006), .B2(n11467), .ZN(
        n11273) );
  OAI211_X1 U13859 ( .C1(n13061), .C2(n13008), .A(n11274), .B(n11273), .ZN(
        P3_U3172) );
  NAND2_X1 U13860 ( .A1(n13560), .A2(P3_U3897), .ZN(n11275) );
  OAI21_X1 U13861 ( .B1(P3_U3897), .B2(n11276), .A(n11275), .ZN(P3_U3509) );
  NAND2_X1 U13862 ( .A1(n13532), .A2(P3_U3897), .ZN(n11277) );
  OAI21_X1 U13863 ( .B1(P3_U3897), .B2(n11278), .A(n11277), .ZN(P3_U3511) );
  NAND2_X1 U13864 ( .A1(n11427), .A2(P3_U3897), .ZN(n11279) );
  OAI21_X1 U13865 ( .B1(P3_U3897), .B2(n11280), .A(n11279), .ZN(P3_U3495) );
  NAND2_X1 U13866 ( .A1(n15808), .A2(P3_U3897), .ZN(n11281) );
  OAI21_X1 U13867 ( .B1(P3_U3897), .B2(n11282), .A(n11281), .ZN(P3_U3493) );
  INV_X1 U13868 ( .A(P3_DATAO_REG_22__SCAN_IN), .ZN(n11284) );
  NAND2_X1 U13869 ( .A1(n13482), .A2(P3_U3897), .ZN(n11283) );
  OAI21_X1 U13870 ( .B1(P3_U3897), .B2(n11284), .A(n11283), .ZN(P3_U3513) );
  AOI21_X1 U13871 ( .B1(n11287), .B2(n11286), .A(n11285), .ZN(n11295) );
  NOR2_X1 U13872 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11288), .ZN(n12028) );
  AOI21_X1 U13873 ( .B1(n11291), .B2(n11290), .A(n11289), .ZN(n11292) );
  NOR2_X1 U13874 ( .A1(n15744), .A2(n11292), .ZN(n11293) );
  AOI211_X1 U13875 ( .C1(n15732), .C2(P3_ADDR_REG_6__SCAN_IN), .A(n12028), .B(
        n11293), .ZN(n11294) );
  OAI21_X1 U13876 ( .B1(n11295), .B2(n15752), .A(n11294), .ZN(n11302) );
  INV_X1 U13877 ( .A(n11310), .ZN(n11300) );
  NAND3_X1 U13878 ( .A1(n11298), .A2(n11297), .A3(n11296), .ZN(n11299) );
  AOI21_X1 U13879 ( .B1(n11300), .B2(n11299), .A(n15746), .ZN(n11301) );
  AOI211_X1 U13880 ( .C1(n13349), .C2(n11303), .A(n11302), .B(n11301), .ZN(
        n11304) );
  INV_X1 U13881 ( .A(n11304), .ZN(P3_U3188) );
  AOI21_X1 U13882 ( .B1(n11307), .B2(n11306), .A(n11305), .ZN(n11322) );
  INV_X1 U13883 ( .A(n11417), .ZN(n11312) );
  NOR3_X1 U13884 ( .A1(n11310), .A2(n11309), .A3(n11308), .ZN(n11311) );
  OAI21_X1 U13885 ( .B1(n11312), .B2(n11311), .A(n13395), .ZN(n11321) );
  AOI21_X1 U13886 ( .B1(n10666), .B2(n11314), .A(n11313), .ZN(n11318) );
  AND2_X1 U13887 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n12155) );
  AOI21_X1 U13888 ( .B1(n15732), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n12155), .ZN(
        n11317) );
  NAND2_X1 U13889 ( .A1(n13349), .A2(n11315), .ZN(n11316) );
  OAI211_X1 U13890 ( .C1(n11318), .C2(n15744), .A(n11317), .B(n11316), .ZN(
        n11319) );
  INV_X1 U13891 ( .A(n11319), .ZN(n11320) );
  OAI211_X1 U13892 ( .C1(n11322), .C2(n15752), .A(n11321), .B(n11320), .ZN(
        P3_U3189) );
  NAND2_X1 U13893 ( .A1(n13483), .A2(P3_U3897), .ZN(n11323) );
  OAI21_X1 U13894 ( .B1(P3_U3897), .B2(n11324), .A(n11323), .ZN(P3_U3515) );
  XOR2_X1 U13895 ( .A(n11325), .B(n11328), .Z(n11586) );
  AOI211_X1 U13896 ( .C1(n11590), .C2(n11326), .A(n15263), .B(n11386), .ZN(
        n11594) );
  XOR2_X1 U13897 ( .A(n11328), .B(n11327), .Z(n11330) );
  OAI21_X1 U13898 ( .B1(n11330), .B2(n15668), .A(n11329), .ZN(n11587) );
  AOI211_X1 U13899 ( .C1(n11586), .C2(n15722), .A(n11594), .B(n11587), .ZN(
        n11335) );
  AOI22_X1 U13900 ( .A1(n14333), .A2(n11590), .B1(n15729), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n11331) );
  OAI21_X1 U13901 ( .B1(n11335), .B2(n15729), .A(n11331), .ZN(P2_U3504) );
  INV_X1 U13902 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11332) );
  NOR2_X1 U13903 ( .A1(n15724), .A2(n11332), .ZN(n11333) );
  AOI21_X1 U13904 ( .B1(n9774), .B2(n11590), .A(n11333), .ZN(n11334) );
  OAI21_X1 U13905 ( .B1(n11335), .B2(n9771), .A(n11334), .ZN(P2_U3445) );
  INV_X1 U13906 ( .A(n11336), .ZN(n11338) );
  NAND2_X1 U13907 ( .A1(n11338), .A2(n11337), .ZN(n11339) );
  XNOR2_X1 U13908 ( .A(n11395), .B(n13806), .ZN(n11341) );
  AND2_X1 U13909 ( .A1(n13942), .A2(n13804), .ZN(n11342) );
  NAND2_X1 U13910 ( .A1(n11341), .A2(n11342), .ZN(n11482) );
  INV_X1 U13911 ( .A(n11341), .ZN(n11481) );
  INV_X1 U13912 ( .A(n11342), .ZN(n11343) );
  NAND2_X1 U13913 ( .A1(n11481), .A2(n11343), .ZN(n11344) );
  NAND2_X1 U13914 ( .A1(n11482), .A2(n11344), .ZN(n11346) );
  AOI21_X1 U13915 ( .B1(n11345), .B2(n11346), .A(n13916), .ZN(n11348) );
  NAND2_X1 U13916 ( .A1(n11348), .A2(n11483), .ZN(n11351) );
  AOI22_X1 U13917 ( .A1(n13906), .A2(n13943), .B1(n13941), .B2(n13907), .ZN(
        n11390) );
  NAND2_X1 U13918 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n13989) );
  OAI21_X1 U13919 ( .B1(n13884), .B2(n11390), .A(n13989), .ZN(n11349) );
  AOI21_X1 U13920 ( .B1(n11395), .B2(n13914), .A(n11349), .ZN(n11350) );
  OAI211_X1 U13921 ( .C1(n13912), .C2(n11579), .A(n11351), .B(n11350), .ZN(
        P2_U3211) );
  NAND2_X1 U13922 ( .A1(n15807), .A2(P3_U3897), .ZN(n11352) );
  OAI21_X1 U13923 ( .B1(P3_U3897), .B2(n11353), .A(n11352), .ZN(P3_U3491) );
  NAND2_X1 U13924 ( .A1(n13148), .A2(P3_U3897), .ZN(n11354) );
  OAI21_X1 U13925 ( .B1(P3_U3897), .B2(n11355), .A(n11354), .ZN(P3_U3500) );
  NAND2_X1 U13926 ( .A1(n13559), .A2(P3_U3897), .ZN(n11356) );
  OAI21_X1 U13927 ( .B1(P3_U3897), .B2(n11357), .A(n11356), .ZN(P3_U3507) );
  NAND2_X1 U13928 ( .A1(n13574), .A2(P3_U3897), .ZN(n11358) );
  OAI21_X1 U13929 ( .B1(P3_U3897), .B2(n11359), .A(n11358), .ZN(P3_U3508) );
  NAND2_X1 U13930 ( .A1(n11628), .A2(P3_U3897), .ZN(n11360) );
  OAI21_X1 U13931 ( .B1(P3_U3897), .B2(n11361), .A(n11360), .ZN(P3_U3496) );
  NAND2_X1 U13932 ( .A1(n11963), .A2(P3_U3897), .ZN(n11362) );
  OAI21_X1 U13933 ( .B1(P3_U3897), .B2(n11363), .A(n11362), .ZN(P3_U3497) );
  NAND2_X1 U13934 ( .A1(n15173), .A2(P3_U3897), .ZN(n11364) );
  OAI21_X1 U13935 ( .B1(P3_U3897), .B2(n11365), .A(n11364), .ZN(P3_U3506) );
  NAND2_X1 U13936 ( .A1(n15187), .A2(P3_U3897), .ZN(n11366) );
  OAI21_X1 U13937 ( .B1(P3_U3897), .B2(n11367), .A(n11366), .ZN(P3_U3505) );
  INV_X1 U13938 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n11369) );
  NAND2_X1 U13939 ( .A1(n15199), .A2(P3_U3897), .ZN(n11368) );
  OAI21_X1 U13940 ( .B1(P3_U3897), .B2(n11369), .A(n11368), .ZN(P3_U3504) );
  NAND2_X1 U13941 ( .A1(n12286), .A2(P3_U3897), .ZN(n11370) );
  OAI21_X1 U13942 ( .B1(P3_U3897), .B2(n11371), .A(n11370), .ZN(P3_U3498) );
  OAI21_X1 U13943 ( .B1(n7767), .B2(n11373), .A(n11372), .ZN(n14572) );
  NAND2_X1 U13944 ( .A1(n14572), .A2(n15365), .ZN(n11377) );
  NOR2_X1 U13945 ( .A1(n11374), .A2(P1_U3086), .ZN(n11614) );
  INV_X1 U13946 ( .A(n11614), .ZN(n11375) );
  AOI22_X1 U13947 ( .A1(n11375), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n12115), 
        .B2(n15351), .ZN(n11376) );
  OAI211_X1 U13948 ( .C1(n11508), .C2(n15360), .A(n11377), .B(n11376), .ZN(
        P1_U3232) );
  XNOR2_X1 U13949 ( .A(n11378), .B(n11379), .ZN(n11380) );
  NAND2_X1 U13950 ( .A1(n11380), .A2(n15365), .ZN(n11383) );
  INV_X1 U13951 ( .A(n14561), .ZN(n11381) );
  OAI22_X1 U13952 ( .A1(n11381), .A2(n14967), .B1(n11508), .B2(n14966), .ZN(
        n15492) );
  AOI22_X1 U13953 ( .A1(n15492), .A2(n15348), .B1(n11936), .B2(n15351), .ZN(
        n11382) );
  OAI211_X1 U13954 ( .C1(n11614), .C2(n14576), .A(n11383), .B(n11382), .ZN(
        P1_U3237) );
  XNOR2_X1 U13955 ( .A(n11385), .B(n11384), .ZN(n11575) );
  OAI211_X1 U13956 ( .C1(n11580), .C2(n11386), .A(n14293), .B(n11524), .ZN(
        n11387) );
  INV_X1 U13957 ( .A(n11387), .ZN(n11582) );
  XNOR2_X1 U13958 ( .A(n11389), .B(n11388), .ZN(n11391) );
  OAI21_X1 U13959 ( .B1(n11391), .B2(n15668), .A(n11390), .ZN(n11576) );
  AOI211_X1 U13960 ( .C1(n15722), .C2(n11575), .A(n11582), .B(n11576), .ZN(
        n11397) );
  INV_X1 U13961 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n11392) );
  OAI22_X1 U13962 ( .A1(n14401), .A2(n11580), .B1(n15724), .B2(n11392), .ZN(
        n11393) );
  INV_X1 U13963 ( .A(n11393), .ZN(n11394) );
  OAI21_X1 U13964 ( .B1(n11397), .B2(n9771), .A(n11394), .ZN(P2_U3448) );
  AOI22_X1 U13965 ( .A1(n14333), .A2(n11395), .B1(n15729), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n11396) );
  OAI21_X1 U13966 ( .B1(n11397), .B2(n15729), .A(n11396), .ZN(P2_U3505) );
  NAND2_X1 U13967 ( .A1(n11796), .A2(P3_U3897), .ZN(n11398) );
  OAI21_X1 U13968 ( .B1(P3_U3897), .B2(n11399), .A(n11398), .ZN(P3_U3494) );
  NAND2_X1 U13969 ( .A1(n11400), .A2(P3_U3897), .ZN(n11401) );
  OAI21_X1 U13970 ( .B1(P3_U3897), .B2(n11402), .A(n11401), .ZN(P3_U3492) );
  INV_X1 U13971 ( .A(n11403), .ZN(n11404) );
  AOI21_X1 U13972 ( .B1(n11406), .B2(n11405), .A(n11404), .ZN(n11421) );
  INV_X1 U13973 ( .A(n15732), .ZN(n15737) );
  OR2_X1 U13974 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11407), .ZN(n12269) );
  OAI21_X1 U13975 ( .B1(n15737), .B2(n9565), .A(n12269), .ZN(n11413) );
  NAND2_X1 U13976 ( .A1(n11409), .A2(n11408), .ZN(n11410) );
  AOI21_X1 U13977 ( .B1(n11411), .B2(n11410), .A(n15752), .ZN(n11412) );
  AOI211_X1 U13978 ( .C1(n13349), .C2(n11414), .A(n11413), .B(n11412), .ZN(
        n11420) );
  AND3_X1 U13979 ( .A1(n11417), .A2(n11416), .A3(n11415), .ZN(n11418) );
  OAI21_X1 U13980 ( .B1(n11707), .B2(n11418), .A(n13395), .ZN(n11419) );
  OAI211_X1 U13981 ( .C1(n11421), .C2(n15744), .A(n11420), .B(n11419), .ZN(
        P3_U3190) );
  OAI21_X1 U13982 ( .B1(n11423), .B2(n13063), .A(n11422), .ZN(n15773) );
  NAND2_X1 U13983 ( .A1(n11425), .A2(n11424), .ZN(n11426) );
  AOI21_X1 U13984 ( .B1(n11426), .B2(n13063), .A(n15811), .ZN(n11430) );
  INV_X1 U13985 ( .A(n11427), .ZN(n11976) );
  OAI22_X1 U13986 ( .A1(n7377), .A2(n15789), .B1(n11976), .B2(n15787), .ZN(
        n11428) );
  AOI21_X1 U13987 ( .B1(n11430), .B2(n11429), .A(n11428), .ZN(n15774) );
  INV_X1 U13988 ( .A(n15774), .ZN(n11431) );
  AOI21_X1 U13989 ( .B1(n15241), .B2(n15773), .A(n11431), .ZN(n11550) );
  INV_X1 U13990 ( .A(n13626), .ZN(n13635) );
  AOI22_X1 U13991 ( .A1(n13635), .A2(n15779), .B1(n15851), .B2(
        P3_REG1_REG_3__SCAN_IN), .ZN(n11432) );
  OAI21_X1 U13992 ( .B1(n11550), .B2(n15851), .A(n11432), .ZN(P3_U3462) );
  INV_X1 U13993 ( .A(n11433), .ZN(n11434) );
  INV_X2 U13994 ( .A(n15550), .ZN(n15541) );
  INV_X1 U13995 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n11448) );
  OR2_X1 U13996 ( .A1(n11439), .A2(n10509), .ZN(n11440) );
  NAND2_X1 U13997 ( .A1(n10412), .A2(n14814), .ZN(n11442) );
  OR2_X1 U13998 ( .A1(n12513), .A2(n12393), .ZN(n11441) );
  NAND2_X1 U13999 ( .A1(n15529), .A2(n15393), .ZN(n11444) );
  AOI22_X1 U14000 ( .A1(n11445), .A2(n11444), .B1(n14827), .B2(n14562), .ZN(
        n12118) );
  NAND3_X1 U14001 ( .A1(n12115), .A2(n10563), .A3(n12513), .ZN(n11446) );
  NAND2_X1 U14002 ( .A1(n12118), .A2(n11446), .ZN(n15069) );
  NAND2_X1 U14003 ( .A1(n15069), .A2(n15541), .ZN(n11447) );
  OAI21_X1 U14004 ( .B1(n15541), .B2(n11448), .A(n11447), .ZN(P1_U3459) );
  NAND2_X1 U14005 ( .A1(n15209), .A2(P3_U3897), .ZN(n11449) );
  OAI21_X1 U14006 ( .B1(P3_U3897), .B2(n11450), .A(n11449), .ZN(P3_U3503) );
  INV_X1 U14007 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n11452) );
  NAND2_X1 U14008 ( .A1(n15198), .A2(P3_U3897), .ZN(n11451) );
  OAI21_X1 U14009 ( .B1(P3_U3897), .B2(n11452), .A(n11451), .ZN(P3_U3502) );
  NAND2_X1 U14010 ( .A1(n15208), .A2(P3_U3897), .ZN(n11453) );
  OAI21_X1 U14011 ( .B1(P3_U3897), .B2(n11454), .A(n11453), .ZN(P3_U3501) );
  NAND2_X1 U14012 ( .A1(n13143), .A2(P3_U3897), .ZN(n11455) );
  OAI21_X1 U14013 ( .B1(P3_U3897), .B2(n11456), .A(n11455), .ZN(P3_U3499) );
  INV_X1 U14014 ( .A(n11457), .ZN(n11460) );
  NAND2_X1 U14015 ( .A1(n11461), .A2(n11458), .ZN(n11459) );
  OAI21_X1 U14016 ( .B1(n11461), .B2(n11460), .A(n11459), .ZN(n11462) );
  INV_X1 U14017 ( .A(n11462), .ZN(n11463) );
  INV_X1 U14018 ( .A(n15817), .ZN(n15798) );
  INV_X1 U14019 ( .A(n15760), .ZN(n15780) );
  NAND2_X1 U14020 ( .A1(n15780), .A2(n11467), .ZN(n11469) );
  INV_X2 U14021 ( .A(n15782), .ZN(n15818) );
  AOI22_X1 U14022 ( .A1(n15801), .A2(n11473), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(n15818), .ZN(n11468) );
  OAI211_X1 U14023 ( .C1(n11470), .C2(n15801), .A(n11469), .B(n11468), .ZN(
        P3_U3233) );
  INV_X1 U14024 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11471) );
  NOR2_X1 U14025 ( .A1(n15846), .A2(n11471), .ZN(n11472) );
  AOI21_X1 U14026 ( .B1(n15846), .B2(n11473), .A(n11472), .ZN(n11474) );
  OAI21_X1 U14027 ( .B1(n11475), .B2(n13676), .A(n11474), .ZN(P3_U3390) );
  XNOR2_X1 U14028 ( .A(n11534), .B(n13806), .ZN(n11476) );
  AND2_X1 U14029 ( .A1(n13941), .A2(n13804), .ZN(n11477) );
  NAND2_X1 U14030 ( .A1(n11476), .A2(n11477), .ZN(n11742) );
  INV_X1 U14031 ( .A(n11476), .ZN(n11747) );
  INV_X1 U14032 ( .A(n11477), .ZN(n11478) );
  NAND2_X1 U14033 ( .A1(n11747), .A2(n11478), .ZN(n11479) );
  AND2_X1 U14034 ( .A1(n11742), .A2(n11479), .ZN(n11484) );
  INV_X1 U14035 ( .A(n11484), .ZN(n11480) );
  AOI21_X1 U14036 ( .B1(n11483), .B2(n11480), .A(n13916), .ZN(n11487) );
  NOR3_X1 U14037 ( .A1(n13844), .A2(n11488), .A3(n11481), .ZN(n11486) );
  NAND2_X1 U14038 ( .A1(n11483), .A2(n11482), .ZN(n11485) );
  OAI21_X1 U14039 ( .B1(n11487), .B2(n11486), .A(n11745), .ZN(n11492) );
  INV_X1 U14040 ( .A(n13906), .ZN(n13857) );
  OAI22_X1 U14041 ( .A1(n11488), .A2(n13857), .B1(n11759), .B2(n13855), .ZN(
        n11528) );
  NOR2_X1 U14042 ( .A1(n11489), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14006) );
  NOR2_X1 U14043 ( .A1(n13912), .A2(n11602), .ZN(n11490) );
  AOI211_X1 U14044 ( .C1(n13910), .C2(n11528), .A(n14006), .B(n11490), .ZN(
        n11491) );
  OAI211_X1 U14045 ( .C1(n7469), .C2(n13901), .A(n11492), .B(n11491), .ZN(
        P2_U3185) );
  INV_X1 U14046 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n11495) );
  NAND2_X1 U14047 ( .A1(n13467), .A2(P3_U3897), .ZN(n11494) );
  OAI21_X1 U14048 ( .B1(P3_U3897), .B2(n11495), .A(n11494), .ZN(P3_U3516) );
  XOR2_X1 U14049 ( .A(n11497), .B(n11496), .Z(n11502) );
  AOI22_X1 U14050 ( .A1(n13026), .A2(n11796), .B1(n13006), .B2(n15797), .ZN(
        n11498) );
  OAI21_X1 U14051 ( .B1(n15790), .B2(n13028), .A(n11498), .ZN(n11499) );
  AOI21_X1 U14052 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n11500), .A(n11499), .ZN(
        n11501) );
  OAI21_X1 U14053 ( .B1(n11502), .B2(n13008), .A(n11501), .ZN(P3_U3177) );
  NAND2_X1 U14054 ( .A1(n14563), .A2(n12115), .ZN(n11918) );
  AND3_X1 U14055 ( .A1(n11919), .A2(n15549), .A3(n11918), .ZN(n11513) );
  NAND2_X1 U14056 ( .A1(n15549), .A2(n12115), .ZN(n11504) );
  MUX2_X1 U14057 ( .A(n11504), .B(n15393), .S(n11919), .Z(n11505) );
  NAND2_X1 U14058 ( .A1(n11505), .A2(n14966), .ZN(n11511) );
  NAND2_X1 U14059 ( .A1(n11920), .A2(n11506), .ZN(n15501) );
  OR2_X1 U14060 ( .A1(n11920), .A2(n11506), .ZN(n11507) );
  NAND2_X1 U14061 ( .A1(n15501), .A2(n11507), .ZN(n11514) );
  XNOR2_X1 U14062 ( .A(n11508), .B(n11514), .ZN(n11509) );
  NOR2_X1 U14063 ( .A1(n11509), .A2(n15393), .ZN(n11510) );
  MUX2_X1 U14064 ( .A(n11511), .B(n11510), .S(n11616), .Z(n11512) );
  AOI211_X1 U14065 ( .C1(n14827), .C2(n10536), .A(n11513), .B(n11512), .ZN(
        n11828) );
  INV_X1 U14066 ( .A(n11514), .ZN(n11830) );
  NAND2_X1 U14067 ( .A1(n11830), .A2(n15503), .ZN(n11515) );
  OAI211_X1 U14068 ( .C1(n11920), .C2(n15545), .A(n11828), .B(n11515), .ZN(
        n11517) );
  NAND2_X1 U14069 ( .A1(n11517), .A2(n15559), .ZN(n11516) );
  OAI21_X1 U14070 ( .B1(n15559), .B2(n9941), .A(n11516), .ZN(P1_U3529) );
  INV_X1 U14071 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n11519) );
  NAND2_X1 U14072 ( .A1(n11517), .A2(n15541), .ZN(n11518) );
  OAI21_X1 U14073 ( .B1(n15541), .B2(n11519), .A(n11518), .ZN(P1_U3462) );
  NAND2_X1 U14074 ( .A1(n11520), .A2(P3_U3897), .ZN(n11521) );
  OAI21_X1 U14075 ( .B1(P3_U3897), .B2(n11522), .A(n11521), .ZN(P3_U3517) );
  XNOR2_X1 U14076 ( .A(n11523), .B(n6939), .ZN(n11598) );
  AOI21_X1 U14077 ( .B1(n11534), .B2(n11524), .A(n15263), .ZN(n11525) );
  AND2_X1 U14078 ( .A1(n11654), .A2(n11525), .ZN(n11604) );
  XNOR2_X1 U14079 ( .A(n11527), .B(n11526), .ZN(n11530) );
  INV_X1 U14080 ( .A(n11528), .ZN(n11529) );
  OAI21_X1 U14081 ( .B1(n11530), .B2(n15668), .A(n11529), .ZN(n11599) );
  AOI211_X1 U14082 ( .C1(n15722), .C2(n11598), .A(n11604), .B(n11599), .ZN(
        n11536) );
  INV_X1 U14083 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n11531) );
  OAI22_X1 U14084 ( .A1(n14401), .A2(n7469), .B1(n15724), .B2(n11531), .ZN(
        n11532) );
  INV_X1 U14085 ( .A(n11532), .ZN(n11533) );
  OAI21_X1 U14086 ( .B1(n11536), .B2(n9771), .A(n11533), .ZN(P2_U3451) );
  AOI22_X1 U14087 ( .A1(n14333), .A2(n11534), .B1(n15729), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n11535) );
  OAI21_X1 U14088 ( .B1(n11536), .B2(n15729), .A(n11535), .ZN(P2_U3506) );
  OAI21_X1 U14089 ( .B1(n11538), .B2(n13059), .A(n11537), .ZN(n12113) );
  OAI211_X1 U14090 ( .C1(n13116), .C2(n11539), .A(n11540), .B(n15211), .ZN(
        n11542) );
  AOI22_X1 U14091 ( .A1(n15809), .A2(n11628), .B1(n11796), .B2(n15806), .ZN(
        n11541) );
  NAND2_X1 U14092 ( .A1(n11542), .A2(n11541), .ZN(n12110) );
  AOI21_X1 U14093 ( .B1(n15241), .B2(n12113), .A(n12110), .ZN(n11551) );
  INV_X1 U14094 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n11543) );
  OAI22_X1 U14095 ( .A1(n13676), .A2(n12109), .B1(n15846), .B2(n11543), .ZN(
        n11544) );
  INV_X1 U14096 ( .A(n11544), .ZN(n11545) );
  OAI21_X1 U14097 ( .B1(n11551), .B2(n15844), .A(n11545), .ZN(P3_U3402) );
  INV_X1 U14098 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n11546) );
  OAI22_X1 U14099 ( .A1(n13676), .A2(n11547), .B1(n15846), .B2(n11546), .ZN(
        n11548) );
  INV_X1 U14100 ( .A(n11548), .ZN(n11549) );
  OAI21_X1 U14101 ( .B1(n11550), .B2(n15844), .A(n11549), .ZN(P3_U3399) );
  MUX2_X1 U14102 ( .A(n11552), .B(n11551), .S(n15854), .Z(n11553) );
  OAI21_X1 U14103 ( .B1(n13626), .B2(n12109), .A(n11553), .ZN(P3_U3463) );
  INV_X1 U14104 ( .A(n11554), .ZN(n11555) );
  NAND2_X1 U14105 ( .A1(n11556), .A2(n11555), .ZN(n11561) );
  NAND2_X1 U14106 ( .A1(n11557), .A2(n14272), .ZN(n15651) );
  AND2_X1 U14107 ( .A1(n15711), .A2(n15651), .ZN(n11558) );
  XNOR2_X1 U14108 ( .A(n11559), .B(n11568), .ZN(n15709) );
  INV_X1 U14109 ( .A(n11560), .ZN(n15672) );
  INV_X1 U14110 ( .A(n11562), .ZN(n11565) );
  INV_X1 U14111 ( .A(n11563), .ZN(n11564) );
  OAI211_X1 U14112 ( .C1(n15708), .C2(n11565), .A(n11564), .B(n14293), .ZN(
        n15706) );
  OAI22_X1 U14113 ( .A1(n15654), .A2(n15706), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n15676), .ZN(n11566) );
  AOI21_X1 U14114 ( .B1(n15261), .B2(n13783), .A(n11566), .ZN(n11574) );
  XNOR2_X1 U14115 ( .A(n11567), .B(n11568), .ZN(n11571) );
  NAND2_X1 U14116 ( .A1(n13944), .A2(n13907), .ZN(n11570) );
  NAND2_X1 U14117 ( .A1(n13946), .A2(n13906), .ZN(n11569) );
  NAND2_X1 U14118 ( .A1(n11570), .A2(n11569), .ZN(n13782) );
  AOI21_X1 U14119 ( .B1(n11571), .B2(n15256), .A(n13782), .ZN(n15707) );
  MUX2_X1 U14120 ( .A(n15707), .B(n11572), .S(n15678), .Z(n11573) );
  OAI211_X1 U14121 ( .C1(n14261), .C2(n15709), .A(n11574), .B(n11573), .ZN(
        P2_U3262) );
  INV_X1 U14122 ( .A(n11575), .ZN(n11585) );
  INV_X1 U14123 ( .A(n11576), .ZN(n11577) );
  MUX2_X1 U14124 ( .A(n11578), .B(n11577), .S(n15659), .Z(n11584) );
  OAI22_X1 U14125 ( .A1(n15663), .A2(n11580), .B1(n15676), .B2(n11579), .ZN(
        n11581) );
  AOI21_X1 U14126 ( .B1(n11582), .B2(n15270), .A(n11581), .ZN(n11583) );
  OAI211_X1 U14127 ( .C1(n11585), .C2(n14261), .A(n11584), .B(n11583), .ZN(
        P2_U3259) );
  INV_X1 U14128 ( .A(n11586), .ZN(n11597) );
  INV_X1 U14129 ( .A(n11587), .ZN(n11588) );
  MUX2_X1 U14130 ( .A(n11589), .B(n11588), .S(n15659), .Z(n11596) );
  INV_X1 U14131 ( .A(n11590), .ZN(n11592) );
  OAI22_X1 U14132 ( .A1(n15663), .A2(n11592), .B1(n11591), .B2(n15676), .ZN(
        n11593) );
  AOI21_X1 U14133 ( .B1(n11594), .B2(n15270), .A(n11593), .ZN(n11595) );
  OAI211_X1 U14134 ( .C1(n14261), .C2(n11597), .A(n11596), .B(n11595), .ZN(
        P2_U3260) );
  INV_X1 U14135 ( .A(n11598), .ZN(n11607) );
  INV_X1 U14136 ( .A(n11599), .ZN(n11600) );
  MUX2_X1 U14137 ( .A(n11601), .B(n11600), .S(n15659), .Z(n11606) );
  OAI22_X1 U14138 ( .A1(n7469), .A2(n15663), .B1(n11602), .B2(n15676), .ZN(
        n11603) );
  AOI21_X1 U14139 ( .B1(n11604), .B2(n15270), .A(n11603), .ZN(n11605) );
  OAI211_X1 U14140 ( .C1(n11607), .C2(n14261), .A(n11606), .B(n11605), .ZN(
        P2_U3258) );
  INV_X1 U14141 ( .A(n11608), .ZN(n11623) );
  OAI222_X1 U14142 ( .A1(P1_U3086), .A2(n12217), .B1(n15104), .B2(n11623), 
        .C1(n11609), .C2(n15086), .ZN(P1_U3341) );
  OAI21_X1 U14143 ( .B1(n11610), .B2(n11612), .A(n11611), .ZN(n11619) );
  OAI22_X1 U14144 ( .A1(n15358), .A2(n11920), .B1(n11614), .B2(n11613), .ZN(
        n11618) );
  OAI22_X1 U14145 ( .A1(n11616), .A2(n15361), .B1(n15360), .B2(n11615), .ZN(
        n11617) );
  AOI211_X1 U14146 ( .C1(n11619), .C2(n15365), .A(n11618), .B(n11617), .ZN(
        n11620) );
  INV_X1 U14147 ( .A(n11620), .ZN(P1_U3222) );
  NAND2_X1 U14148 ( .A1(n12868), .A2(P3_U3897), .ZN(n11621) );
  OAI21_X1 U14149 ( .B1(P3_U3897), .B2(n11622), .A(n11621), .ZN(P3_U3518) );
  INV_X1 U14150 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11624) );
  INV_X1 U14151 ( .A(n15605), .ZN(n12358) );
  OAI222_X1 U14152 ( .A1(n14434), .A2(n11624), .B1(n12358), .B2(P2_U3088), 
        .C1(n14428), .C2(n11623), .ZN(P2_U3313) );
  NAND2_X1 U14153 ( .A1(n11625), .A2(n13062), .ZN(n11626) );
  NAND3_X1 U14154 ( .A1(n11627), .A2(n15211), .A3(n11626), .ZN(n11630) );
  AOI22_X1 U14155 ( .A1(n15806), .A2(n11628), .B1(n12286), .B2(n15809), .ZN(
        n11629) );
  AND2_X1 U14156 ( .A1(n11630), .A2(n11629), .ZN(n11773) );
  OR2_X1 U14157 ( .A1(n11631), .A2(n13062), .ZN(n11632) );
  NAND2_X1 U14158 ( .A1(n11633), .A2(n11632), .ZN(n11771) );
  NAND2_X1 U14159 ( .A1(n11771), .A2(n15241), .ZN(n11634) );
  NAND2_X1 U14160 ( .A1(n11773), .A2(n11634), .ZN(n11845) );
  INV_X1 U14161 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n11635) );
  OAI22_X1 U14162 ( .A1(n13676), .A2(n12030), .B1(n15846), .B2(n11635), .ZN(
        n11636) );
  AOI21_X1 U14163 ( .B1(n11845), .B2(n15846), .A(n11636), .ZN(n11637) );
  INV_X1 U14164 ( .A(n11637), .ZN(P3_U3408) );
  OAI22_X1 U14165 ( .A1(n15654), .A2(n11639), .B1(n11638), .B2(n15676), .ZN(
        n11641) );
  NOR2_X1 U14166 ( .A1(n15663), .A2(n6915), .ZN(n11640) );
  AOI211_X1 U14167 ( .C1(n15652), .C2(P2_REG2_REG_2__SCAN_IN), .A(n11641), .B(
        n11640), .ZN(n11644) );
  NAND2_X1 U14168 ( .A1(n11642), .A2(n15659), .ZN(n11643) );
  OAI211_X1 U14169 ( .C1(n14261), .C2(n11645), .A(n11644), .B(n11643), .ZN(
        P2_U3263) );
  XNOR2_X1 U14170 ( .A(n11646), .B(n7517), .ZN(n11871) );
  XNOR2_X1 U14171 ( .A(n11648), .B(n11647), .ZN(n11652) );
  NAND2_X1 U14172 ( .A1(n13941), .A2(n13906), .ZN(n11650) );
  NAND2_X1 U14173 ( .A1(n13939), .A2(n13907), .ZN(n11649) );
  NAND2_X1 U14174 ( .A1(n11650), .A2(n11649), .ZN(n11743) );
  INV_X1 U14175 ( .A(n11743), .ZN(n11651) );
  OAI21_X1 U14176 ( .B1(n11652), .B2(n15668), .A(n11651), .ZN(n11864) );
  INV_X1 U14177 ( .A(n11808), .ZN(n11653) );
  AOI211_X1 U14178 ( .C1(n11754), .C2(n11654), .A(n15263), .B(n11653), .ZN(
        n11870) );
  AOI211_X1 U14179 ( .C1(n15722), .C2(n11871), .A(n11864), .B(n11870), .ZN(
        n11659) );
  INV_X1 U14180 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n11655) );
  OAI22_X1 U14181 ( .A1(n11865), .A2(n14401), .B1(n15724), .B2(n11655), .ZN(
        n11656) );
  INV_X1 U14182 ( .A(n11656), .ZN(n11657) );
  OAI21_X1 U14183 ( .B1(n11659), .B2(n9771), .A(n11657), .ZN(P2_U3454) );
  AOI22_X1 U14184 ( .A1(n14333), .A2(n11754), .B1(n15729), .B2(
        P2_REG1_REG_8__SCAN_IN), .ZN(n11658) );
  OAI21_X1 U14185 ( .B1(n11659), .B2(n15729), .A(n11658), .ZN(P2_U3507) );
  INV_X1 U14186 ( .A(n11660), .ZN(n11662) );
  OAI222_X1 U14187 ( .A1(P3_U3151), .A2(n11663), .B1(n13712), .B2(n11662), 
        .C1(n11661), .C2(n13715), .ZN(P3_U3275) );
  OAI22_X1 U14188 ( .A1(n12083), .A2(n12785), .B1(n12006), .B2(n12787), .ZN(
        n11664) );
  XNOR2_X1 U14189 ( .A(n11664), .B(n12672), .ZN(n11938) );
  OAI22_X1 U14190 ( .A1(n12083), .A2(n12787), .B1(n12006), .B2(n12788), .ZN(
        n11939) );
  XNOR2_X1 U14191 ( .A(n11938), .B(n11939), .ZN(n11691) );
  NAND2_X1 U14192 ( .A1(n14560), .A2(n12848), .ZN(n11666) );
  NAND2_X1 U14193 ( .A1(n14508), .A2(n12849), .ZN(n11665) );
  NAND2_X1 U14194 ( .A1(n11666), .A2(n11665), .ZN(n11686) );
  AND2_X1 U14195 ( .A1(n11685), .A2(n11686), .ZN(n11672) );
  INV_X1 U14196 ( .A(n11672), .ZN(n11682) );
  INV_X1 U14197 ( .A(n11675), .ZN(n11671) );
  INV_X1 U14198 ( .A(n11686), .ZN(n11676) );
  INV_X1 U14199 ( .A(n11668), .ZN(n11674) );
  OAI21_X1 U14200 ( .B1(n11676), .B2(n11667), .A(n11674), .ZN(n11670) );
  INV_X1 U14201 ( .A(n11667), .ZN(n11673) );
  OAI21_X1 U14202 ( .B1(n11673), .B2(n11686), .A(n11668), .ZN(n11669) );
  NAND2_X1 U14203 ( .A1(n11674), .A2(n11673), .ZN(n11678) );
  AND2_X1 U14204 ( .A1(n11678), .A2(n11677), .ZN(n11679) );
  NAND2_X1 U14205 ( .A1(n11683), .A2(n11679), .ZN(n11680) );
  AOI22_X1 U14206 ( .A1(n14560), .A2(n12849), .B1(n12846), .B2(n14508), .ZN(
        n11684) );
  XOR2_X1 U14207 ( .A(n12672), .B(n11684), .Z(n14506) );
  NAND2_X1 U14208 ( .A1(n14507), .A2(n14506), .ZN(n14505) );
  AOI21_X1 U14209 ( .B1(n11691), .B2(n11690), .A(n11942), .ZN(n11698) );
  INV_X1 U14210 ( .A(n11692), .ZN(n12081) );
  INV_X1 U14211 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n11693) );
  OAI22_X1 U14212 ( .A1(n15369), .A2(n12081), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11693), .ZN(n11695) );
  INV_X1 U14213 ( .A(n14558), .ZN(n12076) );
  OAI22_X1 U14214 ( .A1(n11929), .A2(n15361), .B1(n15360), .B2(n12076), .ZN(
        n11694) );
  AOI211_X1 U14215 ( .C1(n11696), .C2(n15351), .A(n11695), .B(n11694), .ZN(
        n11697) );
  OAI21_X1 U14216 ( .B1(n11698), .B2(n15337), .A(n11697), .ZN(P1_U3227) );
  AOI21_X1 U14217 ( .B1(n11701), .B2(n11700), .A(n11699), .ZN(n11716) );
  AOI21_X1 U14218 ( .B1(n10675), .B2(n11703), .A(n11702), .ZN(n11713) );
  INV_X1 U14219 ( .A(n11704), .ZN(n11709) );
  NOR3_X1 U14220 ( .A1(n11707), .A2(n11706), .A3(n11705), .ZN(n11708) );
  OAI21_X1 U14221 ( .B1(n11709), .B2(n11708), .A(n13395), .ZN(n11712) );
  NOR2_X1 U14222 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7986), .ZN(n12457) );
  NOR2_X1 U14223 ( .A1(n15738), .A2(n10623), .ZN(n11710) );
  AOI211_X1 U14224 ( .C1(n15732), .C2(P3_ADDR_REG_9__SCAN_IN), .A(n12457), .B(
        n11710), .ZN(n11711) );
  OAI211_X1 U14225 ( .C1(n11713), .C2(n15744), .A(n11712), .B(n11711), .ZN(
        n11714) );
  INV_X1 U14226 ( .A(n11714), .ZN(n11715) );
  OAI21_X1 U14227 ( .B1(n11716), .B2(n15752), .A(n11715), .ZN(P3_U3191) );
  INV_X1 U14228 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n11720) );
  NAND2_X1 U14229 ( .A1(n7898), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n11719) );
  NAND2_X1 U14230 ( .A1(n11717), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n11718) );
  OAI211_X1 U14231 ( .C1(n11720), .C2(n7909), .A(n11719), .B(n11718), .ZN(
        n11721) );
  INV_X1 U14232 ( .A(n11721), .ZN(n11722) );
  INV_X1 U14233 ( .A(n15161), .ZN(n11724) );
  NAND2_X1 U14234 ( .A1(n11724), .A2(P3_U3897), .ZN(n11725) );
  OAI21_X1 U14235 ( .B1(P3_U3897), .B2(n11726), .A(n11725), .ZN(P3_U3522) );
  INV_X1 U14236 ( .A(n13051), .ZN(n13052) );
  NAND2_X1 U14237 ( .A1(n13052), .A2(P3_U3897), .ZN(n11727) );
  OAI21_X1 U14238 ( .B1(P3_U3897), .B2(n11728), .A(n11727), .ZN(P3_U3521) );
  INV_X1 U14239 ( .A(n13411), .ZN(n11729) );
  NAND2_X1 U14240 ( .A1(n11729), .A2(P3_U3897), .ZN(n11730) );
  OAI21_X1 U14241 ( .B1(P3_U3897), .B2(n11731), .A(n11730), .ZN(P3_U3520) );
  AOI21_X1 U14242 ( .B1(n13006), .B2(n15779), .A(n11732), .ZN(n11734) );
  NAND2_X1 U14243 ( .A1(n13014), .A2(n15808), .ZN(n11733) );
  OAI211_X1 U14244 ( .C1(n11976), .C2(n13016), .A(n11734), .B(n11733), .ZN(
        n11739) );
  AOI211_X1 U14245 ( .C1(n11737), .C2(n11735), .A(n13008), .B(n11736), .ZN(
        n11738) );
  AOI211_X1 U14246 ( .C1(n11740), .C2(n13031), .A(n11739), .B(n11738), .ZN(
        n11741) );
  INV_X1 U14247 ( .A(n11741), .ZN(P3_U3158) );
  XNOR2_X1 U14248 ( .A(n11754), .B(n13806), .ZN(n11764) );
  NAND2_X1 U14249 ( .A1(n13940), .A2(n13804), .ZN(n11756) );
  XNOR2_X1 U14250 ( .A(n11764), .B(n11756), .ZN(n11750) );
  NAND2_X1 U14251 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n14019) );
  NAND2_X1 U14252 ( .A1(n13910), .A2(n11743), .ZN(n11744) );
  OAI211_X1 U14253 ( .C1(n13912), .C2(n11866), .A(n14019), .B(n11744), .ZN(
        n11753) );
  INV_X1 U14254 ( .A(n11745), .ZN(n11749) );
  NOR3_X1 U14255 ( .A1(n11747), .A2(n13844), .A3(n11746), .ZN(n11748) );
  AOI21_X1 U14256 ( .B1(n11749), .B2(n13880), .A(n11748), .ZN(n11751) );
  NOR2_X1 U14257 ( .A1(n11751), .A2(n11750), .ZN(n11752) );
  AOI211_X1 U14258 ( .C1(n11754), .C2(n13914), .A(n11753), .B(n11752), .ZN(
        n11755) );
  OAI21_X1 U14259 ( .B1(n11763), .B2(n13916), .A(n11755), .ZN(P2_U3193) );
  INV_X1 U14260 ( .A(n11764), .ZN(n11757) );
  NAND2_X1 U14261 ( .A1(n11757), .A2(n11756), .ZN(n11758) );
  XNOR2_X1 U14262 ( .A(n11879), .B(n13806), .ZN(n11896) );
  NAND2_X1 U14263 ( .A1(n13939), .A2(n13804), .ZN(n11897) );
  XNOR2_X1 U14264 ( .A(n11896), .B(n11897), .ZN(n11765) );
  OAI22_X1 U14265 ( .A1(n11760), .A2(n13855), .B1(n11759), .B2(n13857), .ZN(
        n11811) );
  NAND2_X1 U14266 ( .A1(n13910), .A2(n11811), .ZN(n11761) );
  OAI211_X1 U14267 ( .C1(n13912), .C2(n11877), .A(n11762), .B(n11761), .ZN(
        n11769) );
  INV_X1 U14268 ( .A(n11763), .ZN(n11767) );
  AOI22_X1 U14269 ( .A1(n13880), .A2(n11764), .B1(n13877), .B2(n13940), .ZN(
        n11766) );
  NOR3_X1 U14270 ( .A1(n11767), .A2(n11766), .A3(n11765), .ZN(n11768) );
  AOI211_X1 U14271 ( .C1(n11879), .C2(n13914), .A(n11769), .B(n11768), .ZN(
        n11770) );
  OAI21_X1 U14272 ( .B1(n11900), .B2(n13916), .A(n11770), .ZN(P2_U3203) );
  NOR2_X1 U14273 ( .A1(n15817), .A2(n11788), .ZN(n15795) );
  OR2_X1 U14274 ( .A1(n15814), .A2(n15795), .ZN(n15754) );
  INV_X1 U14275 ( .A(n15218), .ZN(n13420) );
  INV_X1 U14276 ( .A(n11771), .ZN(n11776) );
  MUX2_X1 U14277 ( .A(n11773), .B(n11772), .S(n15822), .Z(n11775) );
  AOI22_X1 U14278 ( .A1(n15780), .A2(n11847), .B1(n15818), .B2(n12023), .ZN(
        n11774) );
  OAI211_X1 U14279 ( .C1(n13420), .C2(n11776), .A(n11775), .B(n11774), .ZN(
        P3_U3227) );
  XNOR2_X1 U14280 ( .A(n11777), .B(n11779), .ZN(n15834) );
  INV_X1 U14281 ( .A(n15819), .ZN(n11786) );
  OAI21_X1 U14282 ( .B1(n11780), .B2(n11779), .A(n11778), .ZN(n11783) );
  OAI22_X1 U14283 ( .A1(n11976), .A2(n15789), .B1(n12154), .B2(n15787), .ZN(
        n11782) );
  INV_X1 U14284 ( .A(n15814), .ZN(n13486) );
  NOR2_X1 U14285 ( .A1(n15834), .A2(n13486), .ZN(n11781) );
  AOI211_X1 U14286 ( .C1(n15211), .C2(n11783), .A(n11782), .B(n11781), .ZN(
        n15835) );
  MUX2_X1 U14287 ( .A(n11200), .B(n15835), .S(n15801), .Z(n11785) );
  NOR2_X1 U14288 ( .A1(n11979), .A2(n15815), .ZN(n15837) );
  AOI22_X1 U14289 ( .A1(n15217), .A2(n15837), .B1(n15818), .B2(n11982), .ZN(
        n11784) );
  OAI211_X1 U14290 ( .C1(n15834), .C2(n11786), .A(n11785), .B(n11784), .ZN(
        P3_U3228) );
  INV_X1 U14291 ( .A(n11787), .ZN(n11790) );
  OAI222_X1 U14292 ( .A1(n13712), .A2(n11790), .B1(n13709), .B2(n11789), .C1(
        P3_U3151), .C2(n11788), .ZN(P3_U3274) );
  INV_X1 U14293 ( .A(n11791), .ZN(n12108) );
  OAI21_X1 U14294 ( .B1(n11794), .B2(n11793), .A(n11792), .ZN(n11795) );
  NAND2_X1 U14295 ( .A1(n11795), .A2(n13023), .ZN(n11802) );
  INV_X1 U14296 ( .A(n11796), .ZN(n15788) );
  OAI22_X1 U14297 ( .A1(n12027), .A2(n13016), .B1(n13028), .B2(n15788), .ZN(
        n11800) );
  INV_X1 U14298 ( .A(n11797), .ZN(n11798) );
  OAI21_X1 U14299 ( .B1(n13035), .B2(n12109), .A(n11798), .ZN(n11799) );
  NOR2_X1 U14300 ( .A1(n11800), .A2(n11799), .ZN(n11801) );
  OAI211_X1 U14301 ( .C1(n12108), .C2(n12958), .A(n11802), .B(n11801), .ZN(
        P3_U3170) );
  INV_X1 U14302 ( .A(n12218), .ZN(n15484) );
  INV_X1 U14303 ( .A(n11803), .ZN(n11819) );
  OAI222_X1 U14304 ( .A1(P1_U3086), .A2(n15484), .B1(n15104), .B2(n11819), 
        .C1(n11804), .C2(n15101), .ZN(P1_U3340) );
  XNOR2_X1 U14305 ( .A(n11805), .B(n11806), .ZN(n11880) );
  AOI211_X1 U14306 ( .C1(n11879), .C2(n11808), .A(n15263), .B(n11807), .ZN(
        n11876) );
  XNOR2_X1 U14307 ( .A(n11810), .B(n11809), .ZN(n11813) );
  INV_X1 U14308 ( .A(n11811), .ZN(n11812) );
  OAI21_X1 U14309 ( .B1(n11813), .B2(n15668), .A(n11812), .ZN(n11875) );
  AOI211_X1 U14310 ( .C1(n15722), .C2(n11880), .A(n11876), .B(n11875), .ZN(
        n11818) );
  AOI22_X1 U14311 ( .A1(n11879), .A2(n14333), .B1(n15729), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11814) );
  OAI21_X1 U14312 ( .B1(n11818), .B2(n15729), .A(n11814), .ZN(P2_U3508) );
  INV_X1 U14313 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11815) );
  NOR2_X1 U14314 ( .A1(n15724), .A2(n11815), .ZN(n11816) );
  AOI21_X1 U14315 ( .B1(n11879), .B2(n9774), .A(n11816), .ZN(n11817) );
  OAI21_X1 U14316 ( .B1(n11818), .B2(n9771), .A(n11817), .ZN(P2_U3457) );
  INV_X1 U14317 ( .A(n15615), .ZN(n12362) );
  OAI222_X1 U14318 ( .A1(n14434), .A2(n11820), .B1(n12362), .B2(P2_U3088), 
        .C1(n14428), .C2(n11819), .ZN(P2_U3312) );
  NAND2_X1 U14319 ( .A1(n11821), .A2(P3_U3897), .ZN(n11822) );
  OAI21_X1 U14320 ( .B1(P3_U3897), .B2(n11823), .A(n11822), .ZN(P3_U3519) );
  NAND2_X1 U14321 ( .A1(n14735), .A2(n11824), .ZN(n11825) );
  MUX2_X1 U14322 ( .A(n11828), .B(n11827), .S(n15509), .Z(n11832) );
  NOR2_X1 U14323 ( .A1(n14732), .A2(n14814), .ZN(n11829) );
  AND2_X1 U14324 ( .A1(n15505), .A2(n15503), .ZN(n14946) );
  INV_X1 U14325 ( .A(n14975), .ZN(n15494) );
  AOI22_X1 U14326 ( .A1(n14946), .A2(n11830), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n15494), .ZN(n11831) );
  OAI211_X1 U14327 ( .C1(n11920), .C2(n15497), .A(n11832), .B(n11831), .ZN(
        P1_U3292) );
  XNOR2_X1 U14328 ( .A(n11842), .B(n11833), .ZN(n11835) );
  AOI21_X1 U14329 ( .B1(n11835), .B2(n15256), .A(n11834), .ZN(n15699) );
  OAI21_X1 U14330 ( .B1(n15698), .B2(n8434), .A(n14293), .ZN(n11837) );
  OR2_X1 U14331 ( .A1(n11837), .A2(n11836), .ZN(n15697) );
  INV_X1 U14332 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11838) );
  OAI22_X1 U14333 ( .A1(n15654), .A2(n15697), .B1(n11838), .B2(n15676), .ZN(
        n11840) );
  NOR2_X1 U14334 ( .A1(n15663), .A2(n15698), .ZN(n11839) );
  AOI211_X1 U14335 ( .C1(n15652), .C2(P2_REG2_REG_1__SCAN_IN), .A(n11840), .B(
        n11839), .ZN(n11844) );
  XNOR2_X1 U14336 ( .A(n11842), .B(n11841), .ZN(n15702) );
  NAND2_X1 U14337 ( .A1(n15269), .A2(n15702), .ZN(n11843) );
  OAI211_X1 U14338 ( .C1(n15678), .C2(n15699), .A(n11844), .B(n11843), .ZN(
        P2_U3264) );
  MUX2_X1 U14339 ( .A(n11845), .B(P3_REG1_REG_6__SCAN_IN), .S(n15851), .Z(
        n11846) );
  AOI21_X1 U14340 ( .B1(n13635), .B2(n11847), .A(n11846), .ZN(n11848) );
  INV_X1 U14341 ( .A(n11848), .ZN(P3_U3465) );
  XNOR2_X1 U14342 ( .A(n11850), .B(n11849), .ZN(n11854) );
  OAI22_X1 U14343 ( .A1(n11852), .A2(n13855), .B1(n11851), .B2(n13857), .ZN(
        n11907) );
  INV_X1 U14344 ( .A(n11907), .ZN(n11853) );
  OAI21_X1 U14345 ( .B1(n11854), .B2(n15668), .A(n11853), .ZN(n11989) );
  INV_X1 U14346 ( .A(n11989), .ZN(n11863) );
  INV_X1 U14347 ( .A(n11888), .ZN(n11855) );
  AOI211_X1 U14348 ( .C1(n11991), .C2(n11856), .A(n15263), .B(n11855), .ZN(
        n11988) );
  NOR2_X1 U14349 ( .A1(n11994), .A2(n15663), .ZN(n11858) );
  OAI22_X1 U14350 ( .A1(n15659), .A2(n10867), .B1(n11904), .B2(n15676), .ZN(
        n11857) );
  AOI211_X1 U14351 ( .C1(n11988), .C2(n15270), .A(n11858), .B(n11857), .ZN(
        n11862) );
  XNOR2_X1 U14352 ( .A(n11860), .B(n11859), .ZN(n11990) );
  NAND2_X1 U14353 ( .A1(n11990), .A2(n15269), .ZN(n11861) );
  OAI211_X1 U14354 ( .C1(n15678), .C2(n11863), .A(n11862), .B(n11861), .ZN(
        P2_U3255) );
  INV_X1 U14355 ( .A(n11864), .ZN(n11874) );
  NOR2_X1 U14356 ( .A1(n11865), .A2(n15663), .ZN(n11869) );
  OAI22_X1 U14357 ( .A1(n15659), .A2(n11867), .B1(n11866), .B2(n15676), .ZN(
        n11868) );
  AOI211_X1 U14358 ( .C1(n11870), .C2(n15270), .A(n11869), .B(n11868), .ZN(
        n11873) );
  NAND2_X1 U14359 ( .A1(n11871), .A2(n15269), .ZN(n11872) );
  OAI211_X1 U14360 ( .C1(n15678), .C2(n11874), .A(n11873), .B(n11872), .ZN(
        P2_U3257) );
  AOI21_X1 U14361 ( .B1(n11876), .B2(n9162), .A(n11875), .ZN(n11883) );
  OAI22_X1 U14362 ( .A1(n15659), .A2(n10796), .B1(n11877), .B2(n15676), .ZN(
        n11878) );
  AOI21_X1 U14363 ( .B1(n11879), .B2(n15261), .A(n11878), .ZN(n11882) );
  NAND2_X1 U14364 ( .A1(n11880), .A2(n15269), .ZN(n11881) );
  OAI211_X1 U14365 ( .C1(n11883), .C2(n15678), .A(n11882), .B(n11881), .ZN(
        P2_U3256) );
  XNOR2_X1 U14366 ( .A(n11884), .B(n11892), .ZN(n11887) );
  NAND2_X1 U14367 ( .A1(n13936), .A2(n13907), .ZN(n11886) );
  NAND2_X1 U14368 ( .A1(n13938), .A2(n13906), .ZN(n11885) );
  NAND2_X1 U14369 ( .A1(n11886), .A2(n11885), .ZN(n12101) );
  AOI21_X1 U14370 ( .B1(n11887), .B2(n15256), .A(n12101), .ZN(n15715) );
  AOI211_X1 U14371 ( .C1(n12105), .C2(n11888), .A(n15263), .B(n6825), .ZN(
        n15716) );
  NOR2_X1 U14372 ( .A1(n7476), .A2(n15663), .ZN(n11891) );
  INV_X1 U14373 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11889) );
  OAI22_X1 U14374 ( .A1(n15659), .A2(n11889), .B1(n12103), .B2(n15676), .ZN(
        n11890) );
  AOI211_X1 U14375 ( .C1(n15716), .C2(n15270), .A(n11891), .B(n11890), .ZN(
        n11895) );
  XNOR2_X1 U14376 ( .A(n11893), .B(n11892), .ZN(n15721) );
  NAND2_X1 U14377 ( .A1(n15721), .A2(n15269), .ZN(n11894) );
  OAI211_X1 U14378 ( .C1(n15678), .C2(n15715), .A(n11895), .B(n11894), .ZN(
        P2_U3254) );
  INV_X1 U14379 ( .A(n11896), .ZN(n11898) );
  NAND2_X1 U14380 ( .A1(n11898), .A2(n11897), .ZN(n11899) );
  XNOR2_X1 U14381 ( .A(n11991), .B(n7043), .ZN(n12094) );
  NAND2_X1 U14382 ( .A1(n13938), .A2(n13804), .ZN(n12095) );
  XNOR2_X1 U14383 ( .A(n12094), .B(n12095), .ZN(n11902) );
  AOI21_X1 U14384 ( .B1(n11901), .B2(n11902), .A(n13916), .ZN(n11903) );
  NAND2_X1 U14385 ( .A1(n11903), .A2(n12099), .ZN(n11909) );
  NOR2_X1 U14386 ( .A1(n13912), .A2(n11904), .ZN(n11905) );
  AOI211_X1 U14387 ( .C1(n13910), .C2(n11907), .A(n11906), .B(n11905), .ZN(
        n11908) );
  OAI211_X1 U14388 ( .C1(n11994), .C2(n13901), .A(n11909), .B(n11908), .ZN(
        P2_U3189) );
  OAI21_X1 U14389 ( .B1(n11912), .B2(n11911), .A(n11910), .ZN(n15491) );
  NAND2_X1 U14390 ( .A1(n12138), .A2(n12137), .ZN(n12136) );
  OR2_X1 U14391 ( .A1(n14561), .A2(n15518), .ZN(n11914) );
  NAND2_X1 U14392 ( .A1(n12136), .A2(n11914), .ZN(n12164) );
  NAND2_X1 U14393 ( .A1(n12164), .A2(n12163), .ZN(n11916) );
  NAND2_X1 U14394 ( .A1(n11929), .A2(n14508), .ZN(n11915) );
  NAND2_X1 U14395 ( .A1(n11916), .A2(n11915), .ZN(n11917) );
  NAND2_X1 U14396 ( .A1(n11917), .A2(n12003), .ZN(n12001) );
  OAI21_X1 U14397 ( .B1(n12003), .B2(n11917), .A(n12001), .ZN(n11935) );
  OAI22_X1 U14398 ( .A1(n12076), .A2(n14967), .B1(n11929), .B2(n14966), .ZN(
        n11934) );
  NAND2_X1 U14399 ( .A1(n11919), .A2(n11918), .ZN(n11923) );
  INV_X1 U14400 ( .A(n11920), .ZN(n11921) );
  OR2_X1 U14401 ( .A1(n14562), .A2(n11921), .ZN(n11922) );
  NAND2_X1 U14402 ( .A1(n11923), .A2(n11922), .ZN(n15499) );
  OR2_X1 U14403 ( .A1(n10536), .A2(n11936), .ZN(n11924) );
  NAND2_X1 U14404 ( .A1(n11925), .A2(n11924), .ZN(n12129) );
  NAND2_X1 U14405 ( .A1(n12129), .A2(n12130), .ZN(n11927) );
  OR2_X1 U14406 ( .A1(n14561), .A2(n12131), .ZN(n11926) );
  NAND2_X1 U14407 ( .A1(n11927), .A2(n11926), .ZN(n12162) );
  INV_X1 U14408 ( .A(n12163), .ZN(n11928) );
  NAND2_X1 U14409 ( .A1(n12162), .A2(n11928), .ZN(n11931) );
  INV_X1 U14410 ( .A(n14508), .ZN(n15528) );
  NAND2_X1 U14411 ( .A1(n11929), .A2(n15528), .ZN(n11930) );
  XNOR2_X1 U14412 ( .A(n12005), .B(n12003), .ZN(n11932) );
  NOR2_X1 U14413 ( .A1(n11932), .A2(n15529), .ZN(n11933) );
  AOI211_X1 U14414 ( .C1(n15534), .C2(n11935), .A(n11934), .B(n11933), .ZN(
        n12089) );
  OAI211_X1 U14415 ( .C1(n12170), .C2(n12083), .A(n15503), .B(n11998), .ZN(
        n12086) );
  OAI211_X1 U14416 ( .C1(n12083), .C2(n15545), .A(n12089), .B(n12086), .ZN(
        n11954) );
  NAND2_X1 U14417 ( .A1(n11954), .A2(n15559), .ZN(n11937) );
  OAI21_X1 U14418 ( .B1(n15559), .B2(n10018), .A(n11937), .ZN(P1_U3533) );
  INV_X1 U14419 ( .A(n12055), .ZN(n12052) );
  INV_X1 U14420 ( .A(n11938), .ZN(n11941) );
  INV_X1 U14421 ( .A(n11939), .ZN(n11940) );
  NAND2_X1 U14422 ( .A1(n12055), .A2(n12846), .ZN(n11944) );
  NAND2_X1 U14423 ( .A1(n14558), .A2(n12849), .ZN(n11943) );
  NAND2_X1 U14424 ( .A1(n11944), .A2(n11943), .ZN(n11945) );
  XNOR2_X1 U14425 ( .A(n11945), .B(n12672), .ZN(n12067) );
  AND2_X1 U14426 ( .A1(n14558), .A2(n12848), .ZN(n11946) );
  AOI21_X1 U14427 ( .B1(n12055), .B2(n12849), .A(n11946), .ZN(n12068) );
  XNOR2_X1 U14428 ( .A(n12067), .B(n12068), .ZN(n11947) );
  OAI211_X1 U14429 ( .C1(n11948), .C2(n11947), .A(n12071), .B(n15365), .ZN(
        n11953) );
  INV_X1 U14430 ( .A(n12014), .ZN(n11951) );
  OAI22_X1 U14431 ( .A1(n12006), .A2(n15361), .B1(n15360), .B2(n12247), .ZN(
        n11949) );
  AOI211_X1 U14432 ( .C1(n14532), .C2(n11951), .A(n11950), .B(n11949), .ZN(
        n11952) );
  OAI211_X1 U14433 ( .C1(n12052), .C2(n15358), .A(n11953), .B(n11952), .ZN(
        P1_U3239) );
  NAND2_X1 U14434 ( .A1(n11954), .A2(n15541), .ZN(n11955) );
  OAI21_X1 U14435 ( .B1(n15541), .B2(n10019), .A(n11955), .ZN(P1_U3474) );
  INV_X1 U14436 ( .A(n11956), .ZN(n11958) );
  OAI22_X1 U14437 ( .A1(n13243), .A2(P3_U3151), .B1(SI_22_), .B2(n13709), .ZN(
        n11957) );
  AOI21_X1 U14438 ( .B1(n11958), .B2(n15121), .A(n11957), .ZN(P3_U3273) );
  OAI21_X1 U14439 ( .B1(n11960), .B2(n13060), .A(n11959), .ZN(n15765) );
  OAI211_X1 U14440 ( .C1(n11962), .C2(n13134), .A(n11961), .B(n15211), .ZN(
        n11965) );
  AOI22_X1 U14441 ( .A1(n15806), .A2(n11963), .B1(n13143), .B2(n15809), .ZN(
        n11964) );
  AND2_X1 U14442 ( .A1(n11965), .A2(n11964), .ZN(n15766) );
  INV_X1 U14443 ( .A(n15766), .ZN(n11966) );
  AOI21_X1 U14444 ( .B1(n15241), .B2(n15765), .A(n11966), .ZN(n11971) );
  INV_X1 U14445 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n11967) );
  OAI22_X1 U14446 ( .A1(n13676), .A2(n12157), .B1(n15846), .B2(n11967), .ZN(
        n11968) );
  INV_X1 U14447 ( .A(n11968), .ZN(n11969) );
  OAI21_X1 U14448 ( .B1(n11971), .B2(n15844), .A(n11969), .ZN(P3_U3411) );
  AOI22_X1 U14449 ( .A1(n13635), .A2(n15770), .B1(n15851), .B2(
        P3_REG1_REG_7__SCAN_IN), .ZN(n11970) );
  OAI21_X1 U14450 ( .B1(n11971), .B2(n15851), .A(n11970), .ZN(P3_U3466) );
  INV_X1 U14451 ( .A(n14661), .ZN(n12221) );
  INV_X1 U14452 ( .A(n11972), .ZN(n11986) );
  OAI222_X1 U14453 ( .A1(P1_U3086), .A2(n12221), .B1(n15104), .B2(n11986), 
        .C1(n11973), .C2(n15101), .ZN(P1_U3339) );
  XOR2_X1 U14454 ( .A(n11975), .B(n11974), .Z(n11985) );
  OAI22_X1 U14455 ( .A1(n11976), .A2(n13028), .B1(n13016), .B2(n12154), .ZN(
        n11981) );
  INV_X1 U14456 ( .A(n11977), .ZN(n11978) );
  OAI21_X1 U14457 ( .B1(n13035), .B2(n11979), .A(n11978), .ZN(n11980) );
  NOR2_X1 U14458 ( .A1(n11981), .A2(n11980), .ZN(n11984) );
  NAND2_X1 U14459 ( .A1(n13031), .A2(n11982), .ZN(n11983) );
  OAI211_X1 U14460 ( .C1(n11985), .C2(n13008), .A(n11984), .B(n11983), .ZN(
        P3_U3167) );
  INV_X1 U14461 ( .A(n15627), .ZN(n12365) );
  OAI222_X1 U14462 ( .A1(n14434), .A2(n11987), .B1(n12365), .B2(P2_U3088), 
        .C1(n14428), .C2(n11986), .ZN(P2_U3311) );
  AOI211_X1 U14463 ( .C1(n15722), .C2(n11990), .A(n11989), .B(n11988), .ZN(
        n11997) );
  AOI22_X1 U14464 ( .A1(n11991), .A2(n14333), .B1(n15729), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n11992) );
  OAI21_X1 U14465 ( .B1(n11997), .B2(n15729), .A(n11992), .ZN(P2_U3509) );
  INV_X1 U14466 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11993) );
  OAI22_X1 U14467 ( .A1(n11994), .A2(n14401), .B1(n15724), .B2(n11993), .ZN(
        n11995) );
  INV_X1 U14468 ( .A(n11995), .ZN(n11996) );
  OAI21_X1 U14469 ( .B1(n11997), .B2(n9771), .A(n11996), .ZN(P2_U3460) );
  INV_X1 U14470 ( .A(n11998), .ZN(n11999) );
  OAI211_X1 U14471 ( .C1(n11999), .C2(n12052), .A(n15503), .B(n12048), .ZN(
        n12018) );
  NAND2_X1 U14472 ( .A1(n12001), .A2(n12000), .ZN(n12002) );
  OAI21_X1 U14473 ( .B1(n12002), .B2(n12049), .A(n12057), .ZN(n12012) );
  OAI22_X1 U14474 ( .A1(n12247), .A2(n14967), .B1(n12006), .B2(n14966), .ZN(
        n12011) );
  INV_X1 U14475 ( .A(n12003), .ZN(n12004) );
  NAND2_X1 U14476 ( .A1(n12005), .A2(n12004), .ZN(n12008) );
  NAND2_X1 U14477 ( .A1(n12083), .A2(n12006), .ZN(n12007) );
  NAND2_X1 U14478 ( .A1(n12008), .A2(n12007), .ZN(n12051) );
  XNOR2_X1 U14479 ( .A(n12051), .B(n12049), .ZN(n12009) );
  NOR2_X1 U14480 ( .A1(n12009), .A2(n15529), .ZN(n12010) );
  AOI211_X1 U14481 ( .C1(n15534), .C2(n12012), .A(n12011), .B(n12010), .ZN(
        n12019) );
  INV_X2 U14482 ( .A(n15495), .ZN(n14922) );
  MUX2_X1 U14483 ( .A(n12013), .B(n12019), .S(n14922), .Z(n12017) );
  OAI22_X1 U14484 ( .A1(n15497), .A2(n12052), .B1(n14975), .B2(n12014), .ZN(
        n12015) );
  INV_X1 U14485 ( .A(n12015), .ZN(n12016) );
  OAI211_X1 U14486 ( .C1(n14873), .C2(n12018), .A(n12017), .B(n12016), .ZN(
        P1_U3287) );
  OAI211_X1 U14487 ( .C1(n12052), .C2(n15545), .A(n12019), .B(n12018), .ZN(
        n12021) );
  NAND2_X1 U14488 ( .A1(n12021), .A2(n15559), .ZN(n12020) );
  OAI21_X1 U14489 ( .B1(n15559), .B2(n10037), .A(n12020), .ZN(P1_U3534) );
  NAND2_X1 U14490 ( .A1(n12021), .A2(n15541), .ZN(n12022) );
  OAI21_X1 U14491 ( .B1(n15541), .B2(n10043), .A(n12022), .ZN(P1_U3477) );
  INV_X1 U14492 ( .A(n12023), .ZN(n12035) );
  OAI211_X1 U14493 ( .C1(n12026), .C2(n12025), .A(n12024), .B(n13023), .ZN(
        n12034) );
  INV_X1 U14494 ( .A(n12286), .ZN(n12268) );
  OAI22_X1 U14495 ( .A1(n12027), .A2(n13028), .B1(n13016), .B2(n12268), .ZN(
        n12032) );
  INV_X1 U14496 ( .A(n12028), .ZN(n12029) );
  OAI21_X1 U14497 ( .B1(n13035), .B2(n12030), .A(n12029), .ZN(n12031) );
  NOR2_X1 U14498 ( .A1(n12032), .A2(n12031), .ZN(n12033) );
  OAI211_X1 U14499 ( .C1(n12035), .C2(n12958), .A(n12034), .B(n12033), .ZN(
        P3_U3179) );
  INV_X1 U14500 ( .A(n12036), .ZN(n12065) );
  OAI222_X1 U14501 ( .A1(P1_U3086), .A2(n12503), .B1(n15104), .B2(n12065), 
        .C1(n12037), .C2(n15086), .ZN(P1_U3338) );
  XOR2_X1 U14502 ( .A(n12042), .B(n12038), .Z(n12041) );
  NAND2_X1 U14503 ( .A1(n13935), .A2(n13907), .ZN(n12040) );
  NAND2_X1 U14504 ( .A1(n13937), .A2(n13906), .ZN(n12039) );
  NAND2_X1 U14505 ( .A1(n12040), .A2(n12039), .ZN(n12187) );
  AOI21_X1 U14506 ( .B1(n12041), .B2(n15256), .A(n12187), .ZN(n15290) );
  XOR2_X1 U14507 ( .A(n12043), .B(n12042), .Z(n15291) );
  INV_X1 U14508 ( .A(n15291), .ZN(n15294) );
  OAI211_X1 U14509 ( .C1(n15289), .C2(n6825), .A(n14293), .B(n12197), .ZN(
        n15288) );
  INV_X1 U14510 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n12354) );
  OAI22_X1 U14511 ( .A1(n15659), .A2(n12354), .B1(n12189), .B2(n15676), .ZN(
        n12044) );
  AOI21_X1 U14512 ( .B1(n12191), .B2(n15261), .A(n12044), .ZN(n12045) );
  OAI21_X1 U14513 ( .B1(n15288), .B2(n15654), .A(n12045), .ZN(n12046) );
  AOI21_X1 U14514 ( .B1(n15294), .B2(n15269), .A(n12046), .ZN(n12047) );
  OAI21_X1 U14515 ( .B1(n15678), .B2(n15290), .A(n12047), .ZN(P2_U3253) );
  AOI211_X1 U14516 ( .C1(n12248), .C2(n12048), .A(n15061), .B(n12258), .ZN(
        n12149) );
  INV_X1 U14517 ( .A(n12049), .ZN(n12050) );
  NAND2_X1 U14518 ( .A1(n12051), .A2(n12050), .ZN(n12054) );
  NAND2_X1 U14519 ( .A1(n12052), .A2(n12076), .ZN(n12053) );
  XNOR2_X1 U14520 ( .A(n12243), .B(n7349), .ZN(n12061) );
  NAND2_X1 U14521 ( .A1(n12055), .A2(n12076), .ZN(n12056) );
  XNOR2_X1 U14522 ( .A(n12246), .B(n7349), .ZN(n12058) );
  NAND2_X1 U14523 ( .A1(n12058), .A2(n15534), .ZN(n12060) );
  AOI22_X1 U14524 ( .A1(n14825), .A2(n14558), .B1(n14556), .B2(n14827), .ZN(
        n12059) );
  OAI211_X1 U14525 ( .C1(n12061), .C2(n15529), .A(n12060), .B(n12059), .ZN(
        n12146) );
  AOI211_X1 U14526 ( .C1(n15387), .C2(n12248), .A(n12149), .B(n12146), .ZN(
        n12063) );
  OR2_X1 U14527 ( .A1(n12063), .A2(n15557), .ZN(n12062) );
  OAI21_X1 U14528 ( .B1(n15559), .B2(n10924), .A(n12062), .ZN(P1_U3535) );
  OR2_X1 U14529 ( .A1(n12063), .A2(n15550), .ZN(n12064) );
  OAI21_X1 U14530 ( .B1(n15541), .B2(n10056), .A(n12064), .ZN(P1_U3480) );
  INV_X1 U14531 ( .A(n15640), .ZN(n12368) );
  OAI222_X1 U14532 ( .A1(n14434), .A2(n12066), .B1(n12368), .B2(P2_U3088), 
        .C1(n14428), .C2(n12065), .ZN(P2_U3310) );
  INV_X1 U14533 ( .A(n12248), .ZN(n12245) );
  NAND2_X1 U14534 ( .A1(n12067), .A2(n12069), .ZN(n12070) );
  AND2_X1 U14535 ( .A1(n14557), .A2(n12848), .ZN(n12072) );
  AOI21_X1 U14536 ( .B1(n12248), .B2(n12849), .A(n12072), .ZN(n12231) );
  AOI22_X1 U14537 ( .A1(n12248), .A2(n12846), .B1(n12849), .B2(n14557), .ZN(
        n12073) );
  XNOR2_X1 U14538 ( .A(n12073), .B(n12672), .ZN(n12232) );
  XOR2_X1 U14539 ( .A(n12231), .B(n12232), .Z(n12074) );
  NAND2_X1 U14540 ( .A1(n12075), .A2(n12074), .ZN(n12234) );
  OAI211_X1 U14541 ( .C1(n12075), .C2(n12074), .A(n12234), .B(n15365), .ZN(
        n12080) );
  INV_X1 U14542 ( .A(n12145), .ZN(n12078) );
  AND2_X1 U14543 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n14625) );
  OAI22_X1 U14544 ( .A1(n12076), .A2(n15361), .B1(n15360), .B2(n12551), .ZN(
        n12077) );
  AOI211_X1 U14545 ( .C1(n14532), .C2(n12078), .A(n14625), .B(n12077), .ZN(
        n12079) );
  OAI211_X1 U14546 ( .C1(n12245), .C2(n15358), .A(n12080), .B(n12079), .ZN(
        P1_U3213) );
  NOR2_X1 U14547 ( .A1(n14975), .A2(n12081), .ZN(n12082) );
  AOI21_X1 U14548 ( .B1(n15495), .B2(P1_REG2_REG_5__SCAN_IN), .A(n12082), .ZN(
        n12085) );
  OR2_X1 U14549 ( .A1(n15497), .A2(n12083), .ZN(n12084) );
  OAI211_X1 U14550 ( .C1(n12086), .C2(n14873), .A(n12085), .B(n12084), .ZN(
        n12087) );
  INV_X1 U14551 ( .A(n12087), .ZN(n12088) );
  OAI21_X1 U14552 ( .B1(n12089), .B2(n15509), .A(n12088), .ZN(P1_U3288) );
  XNOR2_X1 U14553 ( .A(n12105), .B(n7043), .ZN(n12090) );
  NAND2_X1 U14554 ( .A1(n13937), .A2(n13804), .ZN(n12091) );
  NAND2_X1 U14555 ( .A1(n12090), .A2(n12091), .ZN(n12182) );
  INV_X1 U14556 ( .A(n12090), .ZN(n12093) );
  INV_X1 U14557 ( .A(n12091), .ZN(n12092) );
  NAND2_X1 U14558 ( .A1(n12093), .A2(n12092), .ZN(n12184) );
  NAND2_X1 U14559 ( .A1(n12182), .A2(n12184), .ZN(n12100) );
  INV_X1 U14560 ( .A(n12094), .ZN(n12097) );
  INV_X1 U14561 ( .A(n12095), .ZN(n12096) );
  NAND2_X1 U14562 ( .A1(n12097), .A2(n12096), .ZN(n12098) );
  XOR2_X1 U14563 ( .A(n12100), .B(n12183), .Z(n12107) );
  NAND2_X1 U14564 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n14035)
         );
  NAND2_X1 U14565 ( .A1(n13910), .A2(n12101), .ZN(n12102) );
  OAI211_X1 U14566 ( .C1(n13912), .C2(n12103), .A(n14035), .B(n12102), .ZN(
        n12104) );
  AOI21_X1 U14567 ( .B1(n12105), .B2(n13914), .A(n12104), .ZN(n12106) );
  OAI21_X1 U14568 ( .B1(n12107), .B2(n13916), .A(n12106), .ZN(P2_U3208) );
  OAI22_X1 U14569 ( .A1(n15760), .A2(n12109), .B1(n12108), .B2(n15782), .ZN(
        n12112) );
  MUX2_X1 U14570 ( .A(n12110), .B(P3_REG2_REG_4__SCAN_IN), .S(n15822), .Z(
        n12111) );
  AOI211_X1 U14571 ( .C1(n15218), .C2(n12113), .A(n12112), .B(n12111), .ZN(
        n12114) );
  INV_X1 U14572 ( .A(n12114), .ZN(P3_U3229) );
  OAI21_X1 U14573 ( .B1(n14963), .B2(n14946), .A(n12115), .ZN(n12117) );
  AOI22_X1 U14574 ( .A1(n15509), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n15494), .ZN(n12116) );
  OAI211_X1 U14575 ( .C1(n15509), .C2(n12118), .A(n12117), .B(n12116), .ZN(
        P1_U3293) );
  NAND2_X1 U14576 ( .A1(n12119), .A2(n13066), .ZN(n12120) );
  NAND3_X1 U14577 ( .A1(n12121), .A2(n15211), .A3(n12120), .ZN(n12123) );
  AOI22_X1 U14578 ( .A1(n15806), .A2(n13143), .B1(n15208), .B2(n15809), .ZN(
        n12122) );
  NAND2_X1 U14579 ( .A1(n12123), .A2(n12122), .ZN(n12276) );
  INV_X1 U14580 ( .A(n12276), .ZN(n12128) );
  XNOR2_X1 U14581 ( .A(n12124), .B(n13066), .ZN(n12274) );
  AOI22_X1 U14582 ( .A1(n15822), .A2(P3_REG2_REG_9__SCAN_IN), .B1(n15818), 
        .B2(n12459), .ZN(n12125) );
  OAI21_X1 U14583 ( .B1(n15760), .B2(n13147), .A(n12125), .ZN(n12126) );
  AOI21_X1 U14584 ( .B1(n12274), .B2(n15218), .A(n12126), .ZN(n12127) );
  OAI21_X1 U14585 ( .B1(n12128), .B2(n15822), .A(n12127), .ZN(P3_U3224) );
  XNOR2_X1 U14586 ( .A(n12129), .B(n12130), .ZN(n15521) );
  NAND2_X1 U14587 ( .A1(n15502), .A2(n12131), .ZN(n12132) );
  NAND2_X1 U14588 ( .A1(n12132), .A2(n15503), .ZN(n12133) );
  NOR2_X1 U14589 ( .A1(n12169), .A2(n12133), .ZN(n15520) );
  INV_X1 U14590 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U14591 ( .A1(n15520), .A2(n15505), .B1(n15494), .B2(n12134), .ZN(
        n12135) );
  OAI21_X1 U14592 ( .B1(n15518), .B2(n15497), .A(n12135), .ZN(n12143) );
  OAI21_X1 U14593 ( .B1(n12138), .B2(n12137), .A(n12136), .ZN(n12139) );
  NAND2_X1 U14594 ( .A1(n12139), .A2(n15534), .ZN(n12141) );
  AOI22_X1 U14595 ( .A1(n14825), .A2(n10536), .B1(n14560), .B2(n14827), .ZN(
        n12140) );
  NAND2_X1 U14596 ( .A1(n12141), .A2(n12140), .ZN(n15517) );
  MUX2_X1 U14597 ( .A(n15517), .B(P1_REG2_REG_3__SCAN_IN), .S(n15509), .Z(
        n12142) );
  AOI211_X1 U14598 ( .C1(n15506), .C2(n15521), .A(n12143), .B(n12142), .ZN(
        n12144) );
  INV_X1 U14599 ( .A(n12144), .ZN(P1_U3290) );
  OAI22_X1 U14600 ( .A1(n15497), .A2(n12245), .B1(n12145), .B2(n14975), .ZN(
        n12148) );
  MUX2_X1 U14601 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n12146), .S(n14922), .Z(
        n12147) );
  AOI211_X1 U14602 ( .C1(n15505), .C2(n12149), .A(n12148), .B(n12147), .ZN(
        n12150) );
  INV_X1 U14603 ( .A(n12150), .ZN(P1_U3286) );
  OAI211_X1 U14604 ( .C1(n12153), .C2(n12152), .A(n12151), .B(n13023), .ZN(
        n12161) );
  INV_X1 U14605 ( .A(n13143), .ZN(n12455) );
  OAI22_X1 U14606 ( .A1(n12154), .A2(n13028), .B1(n13016), .B2(n12455), .ZN(
        n12159) );
  INV_X1 U14607 ( .A(n12155), .ZN(n12156) );
  OAI21_X1 U14608 ( .B1(n13035), .B2(n12157), .A(n12156), .ZN(n12158) );
  NOR2_X1 U14609 ( .A1(n12159), .A2(n12158), .ZN(n12160) );
  OAI211_X1 U14610 ( .C1(n15772), .C2(n12958), .A(n12161), .B(n12160), .ZN(
        P3_U3153) );
  XNOR2_X1 U14611 ( .A(n12162), .B(n12163), .ZN(n15530) );
  XNOR2_X1 U14612 ( .A(n12164), .B(n12163), .ZN(n15533) );
  NAND2_X1 U14613 ( .A1(n14561), .A2(n14825), .ZN(n12166) );
  NAND2_X1 U14614 ( .A1(n14559), .A2(n14827), .ZN(n12165) );
  NAND2_X1 U14615 ( .A1(n12166), .A2(n12165), .ZN(n15525) );
  INV_X1 U14616 ( .A(n14509), .ZN(n12167) );
  AOI22_X1 U14617 ( .A1(n14922), .A2(n15525), .B1(n12167), .B2(n15494), .ZN(
        n12168) );
  OAI21_X1 U14618 ( .B1(n10904), .B2(n14922), .A(n12168), .ZN(n12173) );
  OAI21_X1 U14619 ( .B1(n12169), .B2(n15528), .A(n15503), .ZN(n12171) );
  OR2_X1 U14620 ( .A1(n12171), .A2(n12170), .ZN(n15527) );
  OAI22_X1 U14621 ( .A1(n15497), .A2(n15528), .B1(n15527), .B2(n14873), .ZN(
        n12172) );
  AOI211_X1 U14622 ( .C1(n15533), .C2(n14958), .A(n12173), .B(n12172), .ZN(
        n12174) );
  OAI21_X1 U14623 ( .B1(n14960), .B2(n15530), .A(n12174), .ZN(P1_U3289) );
  NAND2_X1 U14624 ( .A1(n12175), .A2(n15121), .ZN(n12176) );
  OAI211_X1 U14625 ( .C1(n12177), .C2(n13709), .A(n12176), .B(n13245), .ZN(
        P3_U3272) );
  XNOR2_X1 U14626 ( .A(n12191), .B(n7043), .ZN(n12181) );
  INV_X1 U14627 ( .A(n12181), .ZN(n12179) );
  NAND2_X1 U14628 ( .A1(n13936), .A2(n13804), .ZN(n12180) );
  INV_X1 U14629 ( .A(n12180), .ZN(n12178) );
  NAND2_X1 U14630 ( .A1(n12179), .A2(n12178), .ZN(n12401) );
  NAND2_X1 U14631 ( .A1(n12181), .A2(n12180), .ZN(n12399) );
  NAND2_X1 U14632 ( .A1(n12401), .A2(n12399), .ZN(n12186) );
  XOR2_X1 U14633 ( .A(n12186), .B(n12400), .Z(n12193) );
  NAND2_X1 U14634 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n15590)
         );
  NAND2_X1 U14635 ( .A1(n13910), .A2(n12187), .ZN(n12188) );
  OAI211_X1 U14636 ( .C1(n13912), .C2(n12189), .A(n15590), .B(n12188), .ZN(
        n12190) );
  AOI21_X1 U14637 ( .B1(n12191), .B2(n13914), .A(n12190), .ZN(n12192) );
  OAI21_X1 U14638 ( .B1(n12193), .B2(n13916), .A(n12192), .ZN(P2_U3196) );
  XOR2_X1 U14639 ( .A(n12196), .B(n12194), .Z(n12195) );
  AOI22_X1 U14640 ( .A1(n13906), .A2(n13936), .B1(n13934), .B2(n13907), .ZN(
        n12405) );
  OAI21_X1 U14641 ( .B1(n12195), .B2(n15668), .A(n12405), .ZN(n12379) );
  INV_X1 U14642 ( .A(n12379), .ZN(n12204) );
  XNOR2_X1 U14643 ( .A(n6818), .B(n12196), .ZN(n12381) );
  AOI21_X1 U14644 ( .B1(n12197), .B2(n12394), .A(n15263), .ZN(n12198) );
  AND2_X1 U14645 ( .A1(n12198), .A2(n15264), .ZN(n12380) );
  NAND2_X1 U14646 ( .A1(n12380), .A2(n15270), .ZN(n12201) );
  INV_X1 U14647 ( .A(n12199), .ZN(n12407) );
  INV_X1 U14648 ( .A(n15676), .ZN(n15260) );
  AOI22_X1 U14649 ( .A1(n15652), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n12407), 
        .B2(n15260), .ZN(n12200) );
  OAI211_X1 U14650 ( .C1(n7473), .C2(n15663), .A(n12201), .B(n12200), .ZN(
        n12202) );
  AOI21_X1 U14651 ( .B1(n12381), .B2(n15269), .A(n12202), .ZN(n12203) );
  OAI21_X1 U14652 ( .B1(n12204), .B2(n15678), .A(n12203), .ZN(P2_U3252) );
  NOR2_X1 U14653 ( .A1(n12503), .A2(n12205), .ZN(n12206) );
  AOI21_X1 U14654 ( .B1(n12205), .B2(n12503), .A(n12206), .ZN(n12213) );
  OR2_X1 U14655 ( .A1(n14661), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n12208) );
  NAND2_X1 U14656 ( .A1(n14661), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n12207) );
  AND2_X1 U14657 ( .A1(n12208), .A2(n12207), .ZN(n14663) );
  OAI21_X1 U14658 ( .B1(n12613), .B2(n12217), .A(n12209), .ZN(n12210) );
  NOR2_X1 U14659 ( .A1(n12218), .A2(n12210), .ZN(n12211) );
  XNOR2_X1 U14660 ( .A(n12210), .B(n12218), .ZN(n15479) );
  NOR2_X1 U14661 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n15479), .ZN(n15478) );
  NOR2_X1 U14662 ( .A1(n12211), .A2(n15478), .ZN(n14664) );
  NAND2_X1 U14663 ( .A1(n14663), .A2(n14664), .ZN(n14662) );
  OAI21_X1 U14664 ( .B1(n12221), .B2(n10223), .A(n14662), .ZN(n12212) );
  NAND2_X1 U14665 ( .A1(n12213), .A2(n12212), .ZN(n12500) );
  OAI211_X1 U14666 ( .C1(n12213), .C2(n12212), .A(n15462), .B(n12500), .ZN(
        n12227) );
  NAND2_X1 U14667 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14490)
         );
  XNOR2_X1 U14668 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n12503), .ZN(n12223) );
  NOR2_X1 U14669 ( .A1(n12221), .A2(n12214), .ZN(n12215) );
  AOI21_X1 U14670 ( .B1(n12214), .B2(n12221), .A(n12215), .ZN(n14658) );
  AOI21_X1 U14671 ( .B1(n12217), .B2(n10176), .A(n12216), .ZN(n12219) );
  NOR2_X1 U14672 ( .A1(n12218), .A2(n12219), .ZN(n12220) );
  XOR2_X1 U14673 ( .A(n12219), .B(n15484), .Z(n15477) );
  NOR2_X1 U14674 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n15477), .ZN(n15476) );
  NOR2_X1 U14675 ( .A1(n12220), .A2(n15476), .ZN(n14659) );
  NAND2_X1 U14676 ( .A1(n14658), .A2(n14659), .ZN(n14657) );
  OAI21_X1 U14677 ( .B1(n12214), .B2(n12221), .A(n14657), .ZN(n12222) );
  NAND2_X1 U14678 ( .A1(n12223), .A2(n12222), .ZN(n12502) );
  OAI211_X1 U14679 ( .C1(n12223), .C2(n12222), .A(n12502), .B(n15469), .ZN(
        n12224) );
  NAND2_X1 U14680 ( .A1(n14490), .A2(n12224), .ZN(n12225) );
  AOI21_X1 U14681 ( .B1(n15450), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n12225), 
        .ZN(n12226) );
  OAI211_X1 U14682 ( .C1(n15485), .C2(n12503), .A(n12227), .B(n12226), .ZN(
        P1_U3260) );
  AOI22_X1 U14683 ( .A1(n12302), .A2(n12849), .B1(n12848), .B2(n14556), .ZN(
        n12543) );
  NAND2_X1 U14684 ( .A1(n12302), .A2(n12846), .ZN(n12229) );
  NAND2_X1 U14685 ( .A1(n14556), .A2(n12849), .ZN(n12228) );
  NAND2_X1 U14686 ( .A1(n12229), .A2(n12228), .ZN(n12230) );
  XNOR2_X1 U14687 ( .A(n12230), .B(n12672), .ZN(n12542) );
  XOR2_X1 U14688 ( .A(n12543), .B(n12542), .Z(n12236) );
  AOI21_X1 U14689 ( .B1(n12236), .B2(n12235), .A(n12545), .ZN(n12241) );
  OAI21_X1 U14690 ( .B1(n15369), .B2(n12259), .A(n12237), .ZN(n12239) );
  INV_X1 U14691 ( .A(n14555), .ZN(n15313) );
  OAI22_X1 U14692 ( .A1(n12247), .A2(n15361), .B1(n15360), .B2(n15313), .ZN(
        n12238) );
  AOI211_X1 U14693 ( .C1(n12302), .C2(n15351), .A(n12239), .B(n12238), .ZN(
        n12240) );
  OAI21_X1 U14694 ( .B1(n12241), .B2(n15337), .A(n12240), .ZN(P1_U3221) );
  NAND2_X1 U14695 ( .A1(n12245), .A2(n12247), .ZN(n12244) );
  XNOR2_X1 U14696 ( .A(n12298), .B(n12297), .ZN(n12256) );
  OAI22_X1 U14697 ( .A1(n15313), .A2(n14967), .B1(n12247), .B2(n14966), .ZN(
        n12255) );
  NAND2_X1 U14698 ( .A1(n12248), .A2(n12247), .ZN(n12249) );
  INV_X1 U14699 ( .A(n12253), .ZN(n12251) );
  INV_X1 U14700 ( .A(n12304), .ZN(n12252) );
  AOI211_X1 U14701 ( .C1(n12297), .C2(n12253), .A(n15393), .B(n12252), .ZN(
        n12254) );
  AOI211_X1 U14702 ( .C1(n12256), .C2(n15549), .A(n12255), .B(n12254), .ZN(
        n12332) );
  INV_X1 U14703 ( .A(n12332), .ZN(n12261) );
  INV_X1 U14704 ( .A(n12302), .ZN(n12333) );
  AND2_X1 U14705 ( .A1(n12258), .A2(n12333), .ZN(n12310) );
  INV_X1 U14706 ( .A(n12310), .ZN(n12257) );
  OAI211_X1 U14707 ( .C1(n12333), .C2(n12258), .A(n12257), .B(n15503), .ZN(
        n12331) );
  OAI22_X1 U14708 ( .A1(n12331), .A2(n14814), .B1(n14975), .B2(n12259), .ZN(
        n12260) );
  OAI21_X1 U14709 ( .B1(n12261), .B2(n12260), .A(n14922), .ZN(n12263) );
  NAND2_X1 U14710 ( .A1(n14963), .A2(n12302), .ZN(n12262) );
  OAI211_X1 U14711 ( .C1(n10910), .C2(n14922), .A(n12263), .B(n12262), .ZN(
        P1_U3285) );
  INV_X1 U14712 ( .A(n12264), .ZN(n15764) );
  OAI211_X1 U14713 ( .C1(n12267), .C2(n12266), .A(n12265), .B(n13023), .ZN(
        n12273) );
  OAI22_X1 U14714 ( .A1(n12268), .A2(n13028), .B1(n13016), .B2(n9803), .ZN(
        n12271) );
  OAI21_X1 U14715 ( .B1(n13035), .B2(n15759), .A(n12269), .ZN(n12270) );
  NOR2_X1 U14716 ( .A1(n12271), .A2(n12270), .ZN(n12272) );
  OAI211_X1 U14717 ( .C1(n15764), .C2(n12958), .A(n12273), .B(n12272), .ZN(
        P3_U3161) );
  AND2_X1 U14718 ( .A1(n12274), .A2(n15241), .ZN(n12275) );
  NOR2_X1 U14719 ( .A1(n12276), .A2(n12275), .ZN(n12279) );
  INV_X1 U14720 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n12277) );
  MUX2_X1 U14721 ( .A(n12279), .B(n12277), .S(n15844), .Z(n12278) );
  OAI21_X1 U14722 ( .B1(n13676), .B2(n13147), .A(n12278), .ZN(P3_U3417) );
  MUX2_X1 U14723 ( .A(n10675), .B(n12279), .S(n15854), .Z(n12280) );
  OAI21_X1 U14724 ( .B1(n13626), .B2(n13147), .A(n12280), .ZN(P3_U3468) );
  OAI21_X1 U14725 ( .B1(n12282), .B2(n6953), .A(n12281), .ZN(n15755) );
  OAI21_X1 U14726 ( .B1(n13144), .B2(n12284), .A(n12283), .ZN(n12287) );
  NAND2_X1 U14727 ( .A1(n13148), .A2(n13221), .ZN(n13149) );
  INV_X1 U14728 ( .A(n13149), .ZN(n12322) );
  AOI222_X1 U14729 ( .A1(n15211), .A2(n12287), .B1(n12286), .B2(n15806), .C1(
        n12285), .C2(n12322), .ZN(n15756) );
  INV_X1 U14730 ( .A(n15756), .ZN(n12288) );
  AOI21_X1 U14731 ( .B1(n15241), .B2(n15755), .A(n12288), .ZN(n12294) );
  AOI22_X1 U14732 ( .A1(n13635), .A2(n12289), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n15851), .ZN(n12290) );
  OAI21_X1 U14733 ( .B1(n12294), .B2(n15851), .A(n12290), .ZN(P3_U3467) );
  INV_X1 U14734 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n12291) );
  OAI22_X1 U14735 ( .A1(n13676), .A2(n15759), .B1(n15846), .B2(n12291), .ZN(
        n12292) );
  INV_X1 U14736 ( .A(n12292), .ZN(n12293) );
  OAI21_X1 U14737 ( .B1(n12294), .B2(n15844), .A(n12293), .ZN(P3_U3414) );
  INV_X1 U14738 ( .A(n12295), .ZN(n12316) );
  INV_X1 U14739 ( .A(n14674), .ZN(n12510) );
  OAI222_X1 U14740 ( .A1(n15086), .A2(n12296), .B1(n15104), .B2(n12316), .C1(
        P1_U3086), .C2(n12510), .ZN(P1_U3337) );
  OR2_X1 U14741 ( .A1(n12302), .A2(n14556), .ZN(n12299) );
  NAND2_X1 U14742 ( .A1(n12300), .A2(n12299), .ZN(n12467) );
  XNOR2_X1 U14743 ( .A(n12467), .B(n12466), .ZN(n15535) );
  INV_X1 U14744 ( .A(n15535), .ZN(n12315) );
  OR2_X1 U14745 ( .A1(n12302), .A2(n12551), .ZN(n12303) );
  NAND2_X1 U14746 ( .A1(n12305), .A2(n12466), .ZN(n12306) );
  NAND2_X1 U14747 ( .A1(n12470), .A2(n12306), .ZN(n12307) );
  NAND2_X1 U14748 ( .A1(n12307), .A2(n15534), .ZN(n12309) );
  AOI22_X1 U14749 ( .A1(n14825), .A2(n14556), .B1(n14554), .B2(n14827), .ZN(
        n12308) );
  NAND2_X1 U14750 ( .A1(n12309), .A2(n12308), .ZN(n15540) );
  INV_X1 U14751 ( .A(n12554), .ZN(n15537) );
  OAI211_X1 U14752 ( .C1(n12310), .C2(n15537), .A(n15503), .B(n12475), .ZN(
        n15536) );
  OAI22_X1 U14753 ( .A1(n14922), .A2(n10912), .B1(n12550), .B2(n14975), .ZN(
        n12311) );
  AOI21_X1 U14754 ( .B1(n12554), .B2(n14963), .A(n12311), .ZN(n12312) );
  OAI21_X1 U14755 ( .B1(n15536), .B2(n14873), .A(n12312), .ZN(n12313) );
  AOI21_X1 U14756 ( .B1(n15540), .B2(n14922), .A(n12313), .ZN(n12314) );
  OAI21_X1 U14757 ( .B1(n14960), .B2(n12315), .A(n12314), .ZN(P1_U3284) );
  INV_X1 U14758 ( .A(n12579), .ZN(n12374) );
  OAI222_X1 U14759 ( .A1(n14434), .A2(n12317), .B1(n12374), .B2(P2_U3088), 
        .C1(n14428), .C2(n12316), .ZN(P2_U3309) );
  XNOR2_X1 U14760 ( .A(n12318), .B(n13151), .ZN(n12325) );
  OAI211_X1 U14761 ( .C1(n12320), .C2(n13151), .A(n12319), .B(n15211), .ZN(
        n12324) );
  AOI22_X1 U14762 ( .A1(n12322), .A2(n12321), .B1(n15809), .B2(n15198), .ZN(
        n12323) );
  OAI211_X1 U14763 ( .C1(n13486), .C2(n12325), .A(n12324), .B(n12323), .ZN(
        n15840) );
  INV_X1 U14764 ( .A(n15840), .ZN(n12330) );
  INV_X1 U14765 ( .A(n12325), .ZN(n15843) );
  NOR2_X1 U14766 ( .A1(n12520), .A2(n15815), .ZN(n15841) );
  AOI22_X1 U14767 ( .A1(n15217), .A2(n15841), .B1(n15818), .B2(n12514), .ZN(
        n12326) );
  OAI21_X1 U14768 ( .B1(n12327), .B2(n15801), .A(n12326), .ZN(n12328) );
  AOI21_X1 U14769 ( .B1(n15843), .B2(n15819), .A(n12328), .ZN(n12329) );
  OAI21_X1 U14770 ( .B1(n12330), .B2(n15822), .A(n12329), .ZN(P3_U3223) );
  OAI211_X1 U14771 ( .C1(n12333), .C2(n15545), .A(n12332), .B(n12331), .ZN(
        n12335) );
  NAND2_X1 U14772 ( .A1(n12335), .A2(n15559), .ZN(n12334) );
  OAI21_X1 U14773 ( .B1(n15559), .B2(n10926), .A(n12334), .ZN(P1_U3536) );
  INV_X1 U14774 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n12337) );
  NAND2_X1 U14775 ( .A1(n12335), .A2(n15541), .ZN(n12336) );
  OAI21_X1 U14776 ( .B1(n15541), .B2(n12337), .A(n12336), .ZN(P1_U3483) );
  XNOR2_X1 U14777 ( .A(n12365), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n15629) );
  INV_X1 U14778 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n15287) );
  INV_X1 U14779 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n12342) );
  INV_X1 U14780 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n15295) );
  INV_X1 U14781 ( .A(n15586), .ZN(n12355) );
  NAND2_X1 U14782 ( .A1(n12350), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n14042) );
  NAND2_X1 U14783 ( .A1(n14043), .A2(n14042), .ZN(n12340) );
  INV_X1 U14784 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n12338) );
  MUX2_X1 U14785 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n12338), .S(n14040), .Z(
        n12339) );
  NAND2_X1 U14786 ( .A1(n12340), .A2(n12339), .ZN(n14045) );
  NAND2_X1 U14787 ( .A1(n14040), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n12341) );
  MUX2_X1 U14788 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n15295), .S(n15586), .Z(
        n15577) );
  AOI21_X1 U14789 ( .B1(n15295), .B2(n12355), .A(n15580), .ZN(n15597) );
  MUX2_X1 U14790 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n12342), .S(n15594), .Z(
        n15596) );
  NAND2_X1 U14791 ( .A1(n15597), .A2(n15596), .ZN(n15595) );
  OAI21_X1 U14792 ( .B1(n12342), .B2(n12356), .A(n15595), .ZN(n15610) );
  OR2_X1 U14793 ( .A1(n15605), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n12344) );
  NAND2_X1 U14794 ( .A1(n15605), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n12343) );
  AND2_X1 U14795 ( .A1(n12344), .A2(n12343), .ZN(n15609) );
  NAND2_X1 U14796 ( .A1(n15610), .A2(n15609), .ZN(n15608) );
  OAI21_X1 U14797 ( .B1(n15287), .B2(n12358), .A(n15608), .ZN(n12345) );
  NAND2_X1 U14798 ( .A1(n15615), .A2(n12345), .ZN(n12346) );
  XNOR2_X1 U14799 ( .A(n12345), .B(n12362), .ZN(n15619) );
  NAND2_X1 U14800 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n15619), .ZN(n15618) );
  NAND2_X1 U14801 ( .A1(n12346), .A2(n15618), .ZN(n15630) );
  NAND2_X1 U14802 ( .A1(n15629), .A2(n15630), .ZN(n15628) );
  INV_X1 U14803 ( .A(n15628), .ZN(n12347) );
  AOI21_X1 U14804 ( .B1(n15627), .B2(P2_REG1_REG_16__SCAN_IN), .A(n12347), 
        .ZN(n15636) );
  XNOR2_X1 U14805 ( .A(n15640), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15637) );
  INV_X1 U14806 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n12348) );
  OAI22_X1 U14807 ( .A1(n15636), .A2(n15637), .B1(n12348), .B2(n12368), .ZN(
        n12578) );
  XOR2_X1 U14808 ( .A(n12579), .B(n12578), .Z(n12349) );
  NAND2_X1 U14809 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n12349), .ZN(n12581) );
  OAI21_X1 U14810 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n12349), .A(n12581), 
        .ZN(n12378) );
  INV_X1 U14811 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n12369) );
  INV_X1 U14812 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n12364) );
  XOR2_X1 U14813 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n15627), .Z(n15625) );
  INV_X1 U14814 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n12357) );
  NAND2_X1 U14815 ( .A1(n12350), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n12351) );
  MUX2_X1 U14816 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n11889), .S(n14040), .Z(
        n14037) );
  NAND2_X1 U14817 ( .A1(n14038), .A2(n14037), .ZN(n15583) );
  NAND2_X1 U14818 ( .A1(n12353), .A2(n11889), .ZN(n15581) );
  MUX2_X1 U14819 ( .A(n12354), .B(P2_REG2_REG_12__SCAN_IN), .S(n15586), .Z(
        n15582) );
  AOI21_X1 U14820 ( .B1(n15583), .B2(n15581), .A(n15582), .ZN(n15585) );
  AOI21_X1 U14821 ( .B1(n12354), .B2(n12355), .A(n15585), .ZN(n15600) );
  MUX2_X1 U14822 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n12357), .S(n15594), .Z(
        n15599) );
  NAND2_X1 U14823 ( .A1(n15600), .A2(n15599), .ZN(n15598) );
  OAI21_X1 U14824 ( .B1(n12357), .B2(n12356), .A(n15598), .ZN(n12359) );
  NAND2_X1 U14825 ( .A1(n15605), .A2(n12359), .ZN(n12360) );
  XNOR2_X1 U14826 ( .A(n12359), .B(n12358), .ZN(n15607) );
  NAND2_X1 U14827 ( .A1(n15607), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n15606) );
  NAND2_X1 U14828 ( .A1(n12360), .A2(n15606), .ZN(n12361) );
  NAND2_X1 U14829 ( .A1(n15615), .A2(n12361), .ZN(n12363) );
  XNOR2_X1 U14830 ( .A(n12362), .B(n12361), .ZN(n15617) );
  NAND2_X1 U14831 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n15617), .ZN(n15616) );
  NAND2_X1 U14832 ( .A1(n12363), .A2(n15616), .ZN(n15626) );
  NAND2_X1 U14833 ( .A1(n15625), .A2(n15626), .ZN(n15624) );
  OAI21_X1 U14834 ( .B1(n12365), .B2(n12364), .A(n15624), .ZN(n15645) );
  INV_X1 U14835 ( .A(n15645), .ZN(n12367) );
  NAND2_X1 U14836 ( .A1(n15640), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n12366) );
  OAI21_X1 U14837 ( .B1(n15640), .B2(P2_REG2_REG_17__SCAN_IN), .A(n12366), 
        .ZN(n15642) );
  OAI21_X1 U14838 ( .B1(n12369), .B2(n12368), .A(n15643), .ZN(n12574) );
  XNOR2_X1 U14839 ( .A(n12579), .B(n12574), .ZN(n12370) );
  NOR2_X1 U14840 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n12370), .ZN(n12576) );
  AOI21_X1 U14841 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n12370), .A(n12576), 
        .ZN(n12372) );
  OR2_X1 U14842 ( .A1(n12372), .A2(n12371), .ZN(n12377) );
  NOR2_X1 U14843 ( .A1(n12373), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13898) );
  NOR2_X1 U14844 ( .A1(n14004), .A2(n12374), .ZN(n12375) );
  AOI211_X1 U14845 ( .C1(n15635), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n13898), 
        .B(n12375), .ZN(n12376) );
  OAI211_X1 U14846 ( .C1(n12378), .C2(n12583), .A(n12377), .B(n12376), .ZN(
        P2_U3232) );
  AOI211_X1 U14847 ( .C1(n12381), .C2(n15722), .A(n12380), .B(n12379), .ZN(
        n12386) );
  AOI22_X1 U14848 ( .A1(n12394), .A2(n14333), .B1(n15729), .B2(
        P2_REG1_REG_13__SCAN_IN), .ZN(n12382) );
  OAI21_X1 U14849 ( .B1(n12386), .B2(n15729), .A(n12382), .ZN(P2_U3512) );
  INV_X1 U14850 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n12383) );
  OAI22_X1 U14851 ( .A1(n7473), .A2(n14401), .B1(n15724), .B2(n12383), .ZN(
        n12384) );
  INV_X1 U14852 ( .A(n12384), .ZN(n12385) );
  OAI21_X1 U14853 ( .B1(n12386), .B2(n9771), .A(n12385), .ZN(P2_U3469) );
  INV_X1 U14854 ( .A(n12387), .ZN(n12389) );
  OAI222_X1 U14855 ( .A1(P1_U3086), .A2(n14973), .B1(n15104), .B2(n12389), 
        .C1(n12388), .C2(n15101), .ZN(P1_U3336) );
  OAI222_X1 U14856 ( .A1(n14434), .A2(n12390), .B1(n14428), .B2(n12389), .C1(
        P2_U3088), .C2(n9162), .ZN(P2_U3308) );
  INV_X1 U14857 ( .A(n12391), .ZN(n12708) );
  OAI222_X1 U14858 ( .A1(n12393), .A2(P1_U3086), .B1(n15104), .B2(n12708), 
        .C1(n12392), .C2(n15101), .ZN(P1_U3335) );
  XNOR2_X1 U14859 ( .A(n12394), .B(n13806), .ZN(n12440) );
  AND2_X1 U14860 ( .A1(n13935), .A2(n13804), .ZN(n12395) );
  NAND2_X1 U14861 ( .A1(n12440), .A2(n12395), .ZN(n12439) );
  INV_X1 U14862 ( .A(n12440), .ZN(n12397) );
  INV_X1 U14863 ( .A(n12395), .ZN(n12396) );
  NAND2_X1 U14864 ( .A1(n12397), .A2(n12396), .ZN(n12398) );
  AND2_X1 U14865 ( .A1(n12439), .A2(n12398), .ZN(n12403) );
  OAI211_X1 U14866 ( .C1(n12403), .C2(n12402), .A(n6812), .B(n13880), .ZN(
        n12409) );
  OAI22_X1 U14867 ( .A1(n13884), .A2(n12405), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12404), .ZN(n12406) );
  AOI21_X1 U14868 ( .B1(n12407), .B2(n13886), .A(n12406), .ZN(n12408) );
  OAI211_X1 U14869 ( .C1(n7473), .C2(n13901), .A(n12409), .B(n12408), .ZN(
        P2_U3206) );
  MUX2_X1 U14870 ( .A(n12413), .B(P3_REG1_REG_12__SCAN_IN), .S(n13255), .Z(
        n12415) );
  INV_X1 U14871 ( .A(n13247), .ZN(n12414) );
  AOI21_X1 U14872 ( .B1(n12416), .B2(n12415), .A(n12414), .ZN(n12438) );
  INV_X1 U14873 ( .A(n12417), .ZN(n12418) );
  NOR2_X1 U14874 ( .A1(n12419), .A2(n12418), .ZN(n15741) );
  MUX2_X1 U14875 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n10612), .Z(n12420) );
  XOR2_X1 U14876 ( .A(n12425), .B(n12420), .Z(n15740) );
  NOR2_X1 U14877 ( .A1(n12420), .A2(n12426), .ZN(n12422) );
  MUX2_X1 U14878 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n10612), .Z(n13250) );
  XNOR2_X1 U14879 ( .A(n13250), .B(n13255), .ZN(n12421) );
  NOR3_X1 U14880 ( .A1(n15739), .A2(n12422), .A3(n12421), .ZN(n13249) );
  NOR2_X1 U14881 ( .A1(n13249), .A2(n15746), .ZN(n12436) );
  OAI21_X1 U14882 ( .B1(n15739), .B2(n12422), .A(n12421), .ZN(n12435) );
  NOR2_X1 U14883 ( .A1(n12425), .A2(n6748), .ZN(n12427) );
  INV_X1 U14884 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n15735) );
  INV_X1 U14885 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12428) );
  MUX2_X1 U14886 ( .A(n12428), .B(P3_REG2_REG_12__SCAN_IN), .S(n13255), .Z(
        n13257) );
  XNOR2_X1 U14887 ( .A(n13258), .B(n13257), .ZN(n12429) );
  NAND2_X1 U14888 ( .A1(n12430), .A2(n12429), .ZN(n12433) );
  NOR2_X1 U14889 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12431), .ZN(n12915) );
  AOI21_X1 U14890 ( .B1(n15732), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n12915), 
        .ZN(n12432) );
  OAI211_X1 U14891 ( .C1(n15738), .C2(n13255), .A(n12433), .B(n12432), .ZN(
        n12434) );
  AOI21_X1 U14892 ( .B1(n12436), .B2(n12435), .A(n12434), .ZN(n12437) );
  OAI21_X1 U14893 ( .B1(n12438), .B2(n15744), .A(n12437), .ZN(P3_U3194) );
  XNOR2_X1 U14894 ( .A(n15280), .B(n7043), .ZN(n12561) );
  NAND2_X1 U14895 ( .A1(n13934), .A2(n13804), .ZN(n12560) );
  XNOR2_X1 U14896 ( .A(n12561), .B(n12560), .ZN(n12447) );
  NAND3_X1 U14897 ( .A1(n12440), .A2(n13877), .A3(n13935), .ZN(n12441) );
  OAI21_X1 U14898 ( .B1(n6812), .B2(n13916), .A(n12441), .ZN(n12448) );
  NAND2_X1 U14899 ( .A1(n15280), .A2(n13914), .ZN(n12445) );
  NAND2_X1 U14900 ( .A1(n13933), .A2(n13907), .ZN(n12443) );
  NAND2_X1 U14901 ( .A1(n13935), .A2(n13906), .ZN(n12442) );
  NAND2_X1 U14902 ( .A1(n12443), .A2(n12442), .ZN(n15255) );
  AOI22_X1 U14903 ( .A1(n13910), .A2(n15255), .B1(P2_REG3_REG_14__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12444) );
  OAI211_X1 U14904 ( .C1(n13912), .C2(n15258), .A(n12445), .B(n12444), .ZN(
        n12446) );
  AOI21_X1 U14905 ( .B1(n12448), .B2(n12447), .A(n12446), .ZN(n12449) );
  OAI21_X1 U14906 ( .B1(n12562), .B2(n13916), .A(n12449), .ZN(P2_U3187) );
  INV_X1 U14907 ( .A(n12450), .ZN(n12451) );
  AOI21_X1 U14908 ( .B1(n12453), .B2(n12452), .A(n12451), .ZN(n12462) );
  INV_X1 U14909 ( .A(n15208), .ZN(n12454) );
  OAI22_X1 U14910 ( .A1(n12455), .A2(n13028), .B1(n13016), .B2(n12454), .ZN(
        n12456) );
  AOI211_X1 U14911 ( .C1(n13006), .C2(n12458), .A(n12457), .B(n12456), .ZN(
        n12461) );
  NAND2_X1 U14912 ( .A1(n13031), .A2(n12459), .ZN(n12460) );
  OAI211_X1 U14913 ( .C1(n12462), .C2(n13008), .A(n12461), .B(n12460), .ZN(
        P3_U3171) );
  INV_X1 U14914 ( .A(n12463), .ZN(n12512) );
  OAI222_X1 U14915 ( .A1(n14434), .A2(n12465), .B1(n14428), .B2(n12512), .C1(
        P2_U3088), .C2(n12464), .ZN(P2_U3306) );
  OR2_X1 U14916 ( .A1(n12554), .A2(n14555), .ZN(n12468) );
  XOR2_X1 U14917 ( .A(n12527), .B(n12526), .Z(n15542) );
  NAND2_X1 U14918 ( .A1(n12554), .A2(n15313), .ZN(n12469) );
  NAND2_X1 U14919 ( .A1(n12470), .A2(n12469), .ZN(n12474) );
  INV_X1 U14920 ( .A(n12474), .ZN(n12472) );
  NAND2_X1 U14921 ( .A1(n12472), .A2(n12471), .ZN(n12530) );
  INV_X1 U14922 ( .A(n12530), .ZN(n12473) );
  AOI211_X1 U14923 ( .C1(n12526), .C2(n12474), .A(n15393), .B(n12473), .ZN(
        n15546) );
  AOI21_X1 U14924 ( .B1(n12475), .B2(n15543), .A(n15061), .ZN(n12477) );
  INV_X1 U14925 ( .A(n14553), .ZN(n15312) );
  OAI22_X1 U14926 ( .A1(n15312), .A2(n14967), .B1(n15313), .B2(n14966), .ZN(
        n12476) );
  AOI21_X1 U14927 ( .B1(n12477), .B2(n12592), .A(n12476), .ZN(n15544) );
  NOR2_X1 U14928 ( .A1(n15544), .A2(n14814), .ZN(n12478) );
  OAI21_X1 U14929 ( .B1(n15546), .B2(n12478), .A(n14922), .ZN(n12482) );
  OAI22_X1 U14930 ( .A1(n14922), .A2(n12479), .B1(n15321), .B2(n14975), .ZN(
        n12480) );
  AOI21_X1 U14931 ( .B1(n15543), .B2(n14963), .A(n12480), .ZN(n12481) );
  OAI211_X1 U14932 ( .C1(n15542), .C2(n14960), .A(n12482), .B(n12481), .ZN(
        P1_U3283) );
  OAI21_X1 U14933 ( .B1(n12484), .B2(n9666), .A(n12483), .ZN(n15277) );
  INV_X1 U14934 ( .A(n15277), .ZN(n12494) );
  OAI21_X1 U14935 ( .B1(n12487), .B2(n12486), .A(n12485), .ZN(n12488) );
  NAND2_X1 U14936 ( .A1(n12488), .A2(n15256), .ZN(n12489) );
  AOI22_X1 U14937 ( .A1(n13932), .A2(n13907), .B1(n13906), .B2(n13934), .ZN(
        n12567) );
  NAND2_X1 U14938 ( .A1(n12489), .A2(n12567), .ZN(n15275) );
  INV_X1 U14939 ( .A(n12570), .ZN(n15274) );
  INV_X1 U14940 ( .A(n12490), .ZN(n15262) );
  OAI211_X1 U14941 ( .C1(n15274), .C2(n15262), .A(n14293), .B(n14269), .ZN(
        n15273) );
  OAI22_X1 U14942 ( .A1(n15273), .A2(n14272), .B1(n15676), .B2(n12565), .ZN(
        n12491) );
  OAI21_X1 U14943 ( .B1(n15275), .B2(n12491), .A(n15659), .ZN(n12493) );
  AOI22_X1 U14944 ( .A1(n12570), .A2(n15261), .B1(P2_REG2_REG_15__SCAN_IN), 
        .B2(n15678), .ZN(n12492) );
  OAI211_X1 U14945 ( .C1(n12494), .C2(n14261), .A(n12493), .B(n12492), .ZN(
        P2_U3250) );
  INV_X1 U14946 ( .A(n12495), .ZN(n12499) );
  INV_X1 U14947 ( .A(n12496), .ZN(n12497) );
  OAI222_X1 U14948 ( .A1(n13712), .A2(n12499), .B1(n13709), .B2(n12498), .C1(
        P3_U3151), .C2(n12497), .ZN(P3_U3271) );
  OAI21_X1 U14949 ( .B1(n12205), .B2(n12503), .A(n12500), .ZN(n14673) );
  XNOR2_X1 U14950 ( .A(n12510), .B(n14673), .ZN(n12501) );
  NAND2_X1 U14951 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n12501), .ZN(n14676) );
  OAI211_X1 U14952 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n12501), .A(n15462), 
        .B(n14676), .ZN(n12509) );
  NAND2_X1 U14953 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14534)
         );
  OAI21_X1 U14954 ( .B1(n12504), .B2(n12503), .A(n12502), .ZN(n14668) );
  XNOR2_X1 U14955 ( .A(n14668), .B(n12510), .ZN(n12505) );
  NAND2_X1 U14956 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n12505), .ZN(n14670) );
  OAI211_X1 U14957 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n12505), .A(n15469), 
        .B(n14670), .ZN(n12506) );
  NAND2_X1 U14958 ( .A1(n14534), .A2(n12506), .ZN(n12507) );
  AOI21_X1 U14959 ( .B1(n15450), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n12507), 
        .ZN(n12508) );
  OAI211_X1 U14960 ( .C1(n15485), .C2(n12510), .A(n12509), .B(n12508), .ZN(
        P1_U3261) );
  OAI222_X1 U14961 ( .A1(P1_U3086), .A2(n12513), .B1(n15104), .B2(n12512), 
        .C1(n12511), .C2(n15101), .ZN(P1_U3334) );
  INV_X1 U14962 ( .A(n12514), .ZN(n12525) );
  AOI21_X1 U14963 ( .B1(n12516), .B2(n12515), .A(n13008), .ZN(n12518) );
  NAND2_X1 U14964 ( .A1(n12518), .A2(n12517), .ZN(n12524) );
  OAI22_X1 U14965 ( .A1(n9803), .A2(n13028), .B1(n13016), .B2(n12991), .ZN(
        n12522) );
  OAI21_X1 U14966 ( .B1(n13035), .B2(n12520), .A(n12519), .ZN(n12521) );
  NOR2_X1 U14967 ( .A1(n12522), .A2(n12521), .ZN(n12523) );
  OAI211_X1 U14968 ( .C1(n12525), .C2(n12958), .A(n12524), .B(n12523), .ZN(
        P3_U3157) );
  INV_X1 U14969 ( .A(n12531), .ZN(n12599) );
  OR2_X1 U14970 ( .A1(n15403), .A2(n14553), .ZN(n12528) );
  XNOR2_X1 U14971 ( .A(n12617), .B(n12615), .ZN(n12536) );
  NAND2_X1 U14972 ( .A1(n12530), .A2(n12529), .ZN(n12598) );
  OR2_X1 U14973 ( .A1(n15403), .A2(n15312), .ZN(n12532) );
  OAI211_X1 U14974 ( .C1(n12533), .C2(n12615), .A(n12607), .B(n15534), .ZN(
        n12535) );
  AOI22_X1 U14975 ( .A1(n14825), .A2(n14553), .B1(n14551), .B2(n14827), .ZN(
        n12534) );
  OAI211_X1 U14976 ( .C1(n12536), .C2(n15529), .A(n12535), .B(n12534), .ZN(
        n12537) );
  INV_X1 U14977 ( .A(n12537), .ZN(n12652) );
  OAI22_X1 U14978 ( .A1(n14922), .A2(n12538), .B1(n12684), .B2(n14975), .ZN(
        n12540) );
  INV_X1 U14979 ( .A(n12687), .ZN(n12653) );
  OAI211_X1 U14980 ( .C1(n12653), .C2(n6826), .A(n15503), .B(n12644), .ZN(
        n12651) );
  NOR2_X1 U14981 ( .A1(n12651), .A2(n14873), .ZN(n12539) );
  AOI211_X1 U14982 ( .C1(n14963), .C2(n12687), .A(n12540), .B(n12539), .ZN(
        n12541) );
  OAI21_X1 U14983 ( .B1(n12652), .B2(n15509), .A(n12541), .ZN(P1_U3281) );
  INV_X1 U14984 ( .A(n12542), .ZN(n12544) );
  AND2_X1 U14985 ( .A1(n14555), .A2(n12848), .ZN(n12546) );
  AOI21_X1 U14986 ( .B1(n12554), .B2(n12849), .A(n12546), .ZN(n12659) );
  AOI22_X1 U14987 ( .A1(n12554), .A2(n12846), .B1(n12849), .B2(n14555), .ZN(
        n12548) );
  XNOR2_X1 U14988 ( .A(n12548), .B(n12672), .ZN(n12662) );
  XOR2_X1 U14989 ( .A(n12663), .B(n12662), .Z(n12556) );
  OAI21_X1 U14990 ( .B1(n15369), .B2(n12550), .A(n12549), .ZN(n12553) );
  OAI22_X1 U14991 ( .A1(n12551), .A2(n15361), .B1(n15360), .B2(n12601), .ZN(
        n12552) );
  AOI211_X1 U14992 ( .C1(n12554), .C2(n15351), .A(n12553), .B(n12552), .ZN(
        n12555) );
  OAI21_X1 U14993 ( .B1(n12556), .B2(n15337), .A(n12555), .ZN(P1_U3231) );
  INV_X1 U14994 ( .A(n12557), .ZN(n12558) );
  OAI222_X1 U14995 ( .A1(n14434), .A2(n12559), .B1(n14428), .B2(n12558), .C1(
        P2_U3088), .C2(n7046), .ZN(P2_U3305) );
  XNOR2_X1 U14996 ( .A(n12570), .B(n13806), .ZN(n13720) );
  XNOR2_X1 U14997 ( .A(n13719), .B(n13720), .ZN(n12564) );
  AOI22_X1 U14998 ( .A1(n12564), .A2(n13880), .B1(n13877), .B2(n13933), .ZN(
        n12573) );
  AND2_X1 U14999 ( .A1(n13933), .A2(n13804), .ZN(n12563) );
  NAND2_X1 U15000 ( .A1(n12564), .A2(n12563), .ZN(n13723) );
  INV_X1 U15001 ( .A(n13723), .ZN(n12572) );
  NOR2_X1 U15002 ( .A1(n13912), .A2(n12565), .ZN(n12569) );
  OAI22_X1 U15003 ( .A1(n13884), .A2(n12567), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12566), .ZN(n12568) );
  AOI211_X1 U15004 ( .C1(n12570), .C2(n13914), .A(n12569), .B(n12568), .ZN(
        n12571) );
  OAI21_X1 U15005 ( .B1(n12573), .B2(n12572), .A(n12571), .ZN(P2_U3213) );
  NOR2_X1 U15006 ( .A1(n12579), .A2(n12574), .ZN(n12575) );
  NOR2_X1 U15007 ( .A1(n12576), .A2(n12575), .ZN(n12577) );
  XOR2_X1 U15008 ( .A(n12577), .B(P2_REG2_REG_19__SCAN_IN), .Z(n12587) );
  INV_X1 U15009 ( .A(n12587), .ZN(n12585) );
  NAND2_X1 U15010 ( .A1(n12579), .A2(n12578), .ZN(n12580) );
  NAND2_X1 U15011 ( .A1(n12581), .A2(n12580), .ZN(n12582) );
  XNOR2_X1 U15012 ( .A(n12582), .B(n14349), .ZN(n12586) );
  OAI21_X1 U15013 ( .B1(n12586), .B2(n12583), .A(n14004), .ZN(n12584) );
  AOI21_X1 U15014 ( .B1(n12585), .B2(n15644), .A(n12584), .ZN(n12589) );
  AOI22_X1 U15015 ( .A1(n12587), .A2(n15644), .B1(n15639), .B2(n12586), .ZN(
        n12588) );
  MUX2_X1 U15016 ( .A(n12589), .B(n12588), .S(n9162), .Z(n12590) );
  NAND2_X1 U15017 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13793)
         );
  OAI211_X1 U15018 ( .C1(n7836), .C2(n15592), .A(n12590), .B(n13793), .ZN(
        P2_U3233) );
  XNOR2_X1 U15019 ( .A(n12591), .B(n12599), .ZN(n15407) );
  NAND2_X1 U15020 ( .A1(n15403), .A2(n12592), .ZN(n12593) );
  NAND2_X1 U15021 ( .A1(n12593), .A2(n15503), .ZN(n12594) );
  OR2_X1 U15022 ( .A1(n6826), .A2(n12594), .ZN(n15404) );
  NAND2_X1 U15023 ( .A1(n15495), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n12595) );
  OAI21_X1 U15024 ( .B1(n14975), .B2(n15354), .A(n12595), .ZN(n12596) );
  AOI21_X1 U15025 ( .B1(n15403), .B2(n14963), .A(n12596), .ZN(n12597) );
  OAI21_X1 U15026 ( .B1(n15404), .B2(n14873), .A(n12597), .ZN(n12605) );
  INV_X1 U15027 ( .A(n12598), .ZN(n12600) );
  AOI21_X1 U15028 ( .B1(n12600), .B2(n12599), .A(n15393), .ZN(n12603) );
  INV_X1 U15029 ( .A(n14552), .ZN(n15333) );
  OAI22_X1 U15030 ( .A1(n15333), .A2(n14967), .B1(n12601), .B2(n14966), .ZN(
        n15349) );
  AOI21_X1 U15031 ( .B1(n12603), .B2(n12602), .A(n15349), .ZN(n15405) );
  NOR2_X1 U15032 ( .A1(n15405), .A2(n15509), .ZN(n12604) );
  AOI211_X1 U15033 ( .C1(n15407), .C2(n15506), .A(n12605), .B(n12604), .ZN(
        n12606) );
  INV_X1 U15034 ( .A(n12606), .ZN(P1_U3282) );
  INV_X1 U15035 ( .A(n12620), .ZN(n12642) );
  NAND2_X1 U15036 ( .A1(n12643), .A2(n12642), .ZN(n12641) );
  OR2_X1 U15037 ( .A1(n15342), .A2(n15305), .ZN(n12608) );
  NAND2_X1 U15038 ( .A1(n12641), .A2(n12608), .ZN(n12609) );
  NAND2_X1 U15039 ( .A1(n12609), .A2(n12623), .ZN(n12694) );
  OAI21_X1 U15040 ( .B1(n12609), .B2(n12623), .A(n12694), .ZN(n15392) );
  AOI211_X1 U15041 ( .C1(n15386), .C2(n12645), .A(n15061), .B(n7289), .ZN(
        n15384) );
  NAND2_X1 U15042 ( .A1(n15386), .A2(n14963), .ZN(n12612) );
  NOR2_X1 U15043 ( .A1(n14975), .A2(n15311), .ZN(n12610) );
  OAI22_X1 U15044 ( .A1(n15305), .A2(n14966), .B1(n15326), .B2(n14967), .ZN(
        n15385) );
  OAI21_X1 U15045 ( .B1(n12610), .B2(n15385), .A(n14922), .ZN(n12611) );
  OAI211_X1 U15046 ( .C1(n14922), .C2(n12613), .A(n12612), .B(n12611), .ZN(
        n12614) );
  AOI21_X1 U15047 ( .B1(n15384), .B2(n15505), .A(n12614), .ZN(n12626) );
  INV_X1 U15048 ( .A(n12615), .ZN(n12616) );
  OR2_X1 U15049 ( .A1(n12687), .A2(n14552), .ZN(n12618) );
  NAND2_X1 U15050 ( .A1(n12619), .A2(n12618), .ZN(n12640) );
  NAND2_X1 U15051 ( .A1(n12640), .A2(n12620), .ZN(n12622) );
  OR2_X1 U15052 ( .A1(n15342), .A2(n14551), .ZN(n12621) );
  NAND2_X1 U15053 ( .A1(n12624), .A2(n12623), .ZN(n15388) );
  NAND3_X1 U15054 ( .A1(n15389), .A2(n15388), .A3(n15506), .ZN(n12625) );
  OAI211_X1 U15055 ( .C1(n15392), .C2(n14979), .A(n12626), .B(n12625), .ZN(
        P1_U3279) );
  NAND2_X1 U15056 ( .A1(n12629), .A2(n14414), .ZN(n12627) );
  OAI211_X1 U15057 ( .C1(n12628), .C2(n14434), .A(n12627), .B(n9166), .ZN(
        P2_U3304) );
  NAND2_X1 U15058 ( .A1(n12629), .A2(n15090), .ZN(n12631) );
  OAI211_X1 U15059 ( .C1(n12632), .C2(n15101), .A(n12631), .B(n12630), .ZN(
        P1_U3332) );
  XNOR2_X1 U15060 ( .A(n12633), .B(n12636), .ZN(n12634) );
  AOI222_X1 U15061 ( .A1(n15211), .A2(n12634), .B1(n15187), .B2(n15806), .C1(
        n13559), .C2(n15809), .ZN(n13640) );
  XNOR2_X1 U15062 ( .A(n12635), .B(n12636), .ZN(n13638) );
  AOI22_X1 U15063 ( .A1(n15822), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15818), 
        .B2(n13032), .ZN(n12637) );
  OAI21_X1 U15064 ( .B1(n13179), .B2(n15760), .A(n12637), .ZN(n12638) );
  AOI21_X1 U15065 ( .B1(n13638), .B2(n15218), .A(n12638), .ZN(n12639) );
  OAI21_X1 U15066 ( .B1(n13640), .B2(n15822), .A(n12639), .ZN(P3_U3218) );
  XNOR2_X1 U15067 ( .A(n12640), .B(n12642), .ZN(n15395) );
  OAI211_X1 U15068 ( .C1(n12643), .C2(n12642), .A(n15534), .B(n12641), .ZN(
        n15399) );
  INV_X1 U15069 ( .A(n15362), .ZN(n14550) );
  AOI22_X1 U15070 ( .A1(n14550), .A2(n14827), .B1(n14825), .B2(n14552), .ZN(
        n15396) );
  OAI211_X1 U15071 ( .C1(n14975), .C2(n15345), .A(n15399), .B(n15396), .ZN(
        n12649) );
  INV_X1 U15072 ( .A(n12644), .ZN(n12646) );
  INV_X1 U15073 ( .A(n15342), .ZN(n15398) );
  OAI211_X1 U15074 ( .C1(n12646), .C2(n15398), .A(n15503), .B(n12645), .ZN(
        n15397) );
  AOI22_X1 U15075 ( .A1(n15342), .A2(n14963), .B1(P1_REG2_REG_13__SCAN_IN), 
        .B2(n15495), .ZN(n12647) );
  OAI21_X1 U15076 ( .B1(n15397), .B2(n14873), .A(n12647), .ZN(n12648) );
  AOI21_X1 U15077 ( .B1(n12649), .B2(n14922), .A(n12648), .ZN(n12650) );
  OAI21_X1 U15078 ( .B1(n14960), .B2(n15395), .A(n12650), .ZN(P1_U3280) );
  OAI211_X1 U15079 ( .C1(n12653), .C2(n15545), .A(n12652), .B(n12651), .ZN(
        n12655) );
  NAND2_X1 U15080 ( .A1(n12655), .A2(n15559), .ZN(n12654) );
  OAI21_X1 U15081 ( .B1(n15559), .B2(n10996), .A(n12654), .ZN(P1_U3540) );
  INV_X1 U15082 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n12657) );
  NAND2_X1 U15083 ( .A1(n12655), .A2(n15541), .ZN(n12656) );
  OAI21_X1 U15084 ( .B1(n15541), .B2(n12657), .A(n12656), .ZN(P1_U3495) );
  AOI21_X2 U15085 ( .B1(n12663), .B2(n12662), .A(n12661), .ZN(n15315) );
  AOI22_X1 U15086 ( .A1(n15543), .A2(n12849), .B1(n12848), .B2(n14554), .ZN(
        n12667) );
  NAND2_X1 U15087 ( .A1(n15543), .A2(n12846), .ZN(n12665) );
  NAND2_X1 U15088 ( .A1(n14554), .A2(n12849), .ZN(n12664) );
  NAND2_X1 U15089 ( .A1(n12665), .A2(n12664), .ZN(n12666) );
  XNOR2_X1 U15090 ( .A(n12666), .B(n12672), .ZN(n12669) );
  XOR2_X1 U15091 ( .A(n12667), .B(n12669), .Z(n15314) );
  INV_X1 U15092 ( .A(n12667), .ZN(n12668) );
  NAND2_X1 U15093 ( .A1(n15403), .A2(n12846), .ZN(n12671) );
  NAND2_X1 U15094 ( .A1(n14553), .A2(n12849), .ZN(n12670) );
  NAND2_X1 U15095 ( .A1(n12671), .A2(n12670), .ZN(n12673) );
  XNOR2_X1 U15096 ( .A(n12673), .B(n12672), .ZN(n12674) );
  AOI22_X1 U15097 ( .A1(n15403), .A2(n12849), .B1(n12848), .B2(n14553), .ZN(
        n12675) );
  XNOR2_X1 U15098 ( .A(n12674), .B(n12675), .ZN(n15347) );
  INV_X1 U15099 ( .A(n12674), .ZN(n12676) );
  NAND2_X1 U15100 ( .A1(n12687), .A2(n12846), .ZN(n12678) );
  NAND2_X1 U15101 ( .A1(n14552), .A2(n12849), .ZN(n12677) );
  NAND2_X1 U15102 ( .A1(n12678), .A2(n12677), .ZN(n12679) );
  XNOR2_X1 U15103 ( .A(n12679), .B(n10529), .ZN(n12725) );
  AND2_X1 U15104 ( .A1(n14552), .A2(n12848), .ZN(n12680) );
  AOI21_X1 U15105 ( .B1(n12687), .B2(n12849), .A(n12680), .ZN(n12723) );
  XNOR2_X1 U15106 ( .A(n12725), .B(n12723), .ZN(n12681) );
  OAI211_X1 U15107 ( .C1(n12682), .C2(n12681), .A(n12727), .B(n15365), .ZN(
        n12689) );
  OAI22_X1 U15108 ( .A1(n15369), .A2(n12684), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12683), .ZN(n12686) );
  OAI22_X1 U15109 ( .A1(n15312), .A2(n15361), .B1(n15360), .B2(n15305), .ZN(
        n12685) );
  AOI211_X1 U15110 ( .C1(n12687), .C2(n15351), .A(n12686), .B(n12685), .ZN(
        n12688) );
  NAND2_X1 U15111 ( .A1(n12689), .A2(n12688), .ZN(P1_U3224) );
  NAND2_X1 U15112 ( .A1(n15386), .A2(n14550), .ZN(n12690) );
  INV_X1 U15113 ( .A(n12692), .ZN(n12695) );
  OAI21_X1 U15114 ( .B1(n7364), .B2(n12692), .A(n14702), .ZN(n15383) );
  INV_X1 U15115 ( .A(n15383), .ZN(n12704) );
  NAND2_X1 U15116 ( .A1(n12694), .A2(n12693), .ZN(n12696) );
  NOR2_X1 U15117 ( .A1(n12696), .A2(n12695), .ZN(n15380) );
  INV_X1 U15118 ( .A(n14742), .ZN(n15379) );
  OR3_X1 U15119 ( .A1(n15380), .A2(n15379), .A3(n14979), .ZN(n12703) );
  INV_X1 U15120 ( .A(n14700), .ZN(n15378) );
  OAI211_X1 U15121 ( .C1(n15378), .C2(n7289), .A(n15503), .B(n14972), .ZN(
        n15377) );
  AOI22_X1 U15122 ( .A1(n14550), .A2(n14825), .B1(n14827), .B2(n14703), .ZN(
        n15376) );
  INV_X1 U15123 ( .A(n15368), .ZN(n12698) );
  NAND2_X1 U15124 ( .A1(n15494), .A2(n12698), .ZN(n12699) );
  OAI211_X1 U15125 ( .C1(n15377), .C2(n14814), .A(n15376), .B(n12699), .ZN(
        n12701) );
  OAI22_X1 U15126 ( .A1(n15378), .A2(n15497), .B1(n10195), .B2(n14922), .ZN(
        n12700) );
  AOI21_X1 U15127 ( .B1(n12701), .B2(n14922), .A(n12700), .ZN(n12702) );
  OAI211_X1 U15128 ( .C1(n12704), .C2(n14960), .A(n12703), .B(n12702), .ZN(
        P1_U3278) );
  INV_X1 U15129 ( .A(n12705), .ZN(n12718) );
  OAI222_X1 U15130 ( .A1(P1_U3086), .A2(n12706), .B1(n15104), .B2(n12718), 
        .C1(n13040), .C2(n15086), .ZN(P1_U3325) );
  OAI222_X1 U15131 ( .A1(n14428), .A2(n12708), .B1(n12707), .B2(P2_U3088), 
        .C1(n7818), .C2(n14434), .ZN(P2_U3307) );
  AOI21_X1 U15132 ( .B1(n13466), .B2(n12709), .A(n7769), .ZN(n12715) );
  AOI22_X1 U15133 ( .A1(n13483), .A2(n13026), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12711) );
  NAND2_X1 U15134 ( .A1(n13031), .A2(n13488), .ZN(n12710) );
  OAI211_X1 U15135 ( .C1(n13507), .C2(n13028), .A(n12711), .B(n12710), .ZN(
        n12712) );
  AOI21_X1 U15136 ( .B1(n12713), .B2(n13006), .A(n12712), .ZN(n12714) );
  OAI21_X1 U15137 ( .B1(n12715), .B2(n13008), .A(n12714), .ZN(P3_U3156) );
  INV_X1 U15138 ( .A(n14415), .ZN(n12717) );
  OAI222_X1 U15139 ( .A1(P1_U3086), .A2(n10501), .B1(n15104), .B2(n12717), 
        .C1(n12716), .C2(n15101), .ZN(P1_U3327) );
  OAI222_X1 U15140 ( .A1(n14428), .A2(n12718), .B1(n8415), .B2(P2_U3088), .C1(
        n13038), .C2(n14434), .ZN(P2_U3297) );
  NAND2_X1 U15141 ( .A1(n15342), .A2(n12846), .ZN(n12720) );
  NAND2_X1 U15142 ( .A1(n14551), .A2(n12849), .ZN(n12719) );
  NAND2_X1 U15143 ( .A1(n12720), .A2(n12719), .ZN(n12721) );
  XNOR2_X1 U15144 ( .A(n12721), .B(n10529), .ZN(n12730) );
  AND2_X1 U15145 ( .A1(n14551), .A2(n12848), .ZN(n12722) );
  AOI21_X1 U15146 ( .B1(n15342), .B2(n12849), .A(n12722), .ZN(n12728) );
  XNOR2_X1 U15147 ( .A(n12730), .B(n12728), .ZN(n15334) );
  INV_X1 U15148 ( .A(n12723), .ZN(n12724) );
  NAND2_X1 U15149 ( .A1(n12725), .A2(n12724), .ZN(n15335) );
  AND2_X1 U15150 ( .A1(n15334), .A2(n15335), .ZN(n12726) );
  INV_X1 U15151 ( .A(n12728), .ZN(n12729) );
  INV_X1 U15152 ( .A(n15386), .ZN(n15304) );
  OAI22_X1 U15153 ( .A1(n15304), .A2(n12787), .B1(n15362), .B2(n12788), .ZN(
        n12735) );
  NAND2_X1 U15154 ( .A1(n15386), .A2(n12846), .ZN(n12733) );
  OR2_X1 U15155 ( .A1(n15362), .A2(n12787), .ZN(n12732) );
  NAND2_X1 U15156 ( .A1(n12733), .A2(n12732), .ZN(n12734) );
  XNOR2_X1 U15157 ( .A(n12734), .B(n10529), .ZN(n12736) );
  XOR2_X1 U15158 ( .A(n12735), .B(n12736), .Z(n15303) );
  NAND2_X1 U15159 ( .A1(n14700), .A2(n12846), .ZN(n12738) );
  OR2_X1 U15160 ( .A1(n15326), .A2(n12787), .ZN(n12737) );
  NAND2_X1 U15161 ( .A1(n12738), .A2(n12737), .ZN(n12739) );
  XNOR2_X1 U15162 ( .A(n12739), .B(n10529), .ZN(n12740) );
  XNOR2_X1 U15163 ( .A(n12742), .B(n12740), .ZN(n15356) );
  INV_X1 U15164 ( .A(n15326), .ZN(n14699) );
  AOI22_X1 U15165 ( .A1(n14700), .A2(n12849), .B1(n12848), .B2(n14699), .ZN(
        n15357) );
  NAND2_X1 U15166 ( .A1(n15356), .A2(n15357), .ZN(n15355) );
  INV_X1 U15167 ( .A(n12740), .ZN(n12741) );
  NAND2_X1 U15168 ( .A1(n12742), .A2(n12741), .ZN(n12743) );
  NAND2_X1 U15169 ( .A1(n15355), .A2(n12743), .ZN(n15322) );
  OAI22_X1 U15170 ( .A1(n15324), .A2(n12787), .B1(n15359), .B2(n12788), .ZN(
        n12748) );
  NAND2_X1 U15171 ( .A1(n15371), .A2(n12846), .ZN(n12745) );
  NAND2_X1 U15172 ( .A1(n14703), .A2(n12849), .ZN(n12744) );
  NAND2_X1 U15173 ( .A1(n12745), .A2(n12744), .ZN(n12746) );
  XNOR2_X1 U15174 ( .A(n12746), .B(n10529), .ZN(n12747) );
  XOR2_X1 U15175 ( .A(n12748), .B(n12747), .Z(n15323) );
  NAND2_X1 U15176 ( .A1(n15322), .A2(n15323), .ZN(n12752) );
  INV_X1 U15177 ( .A(n12747), .ZN(n12750) );
  INV_X1 U15178 ( .A(n12748), .ZN(n12749) );
  NAND2_X1 U15179 ( .A1(n12750), .A2(n12749), .ZN(n12751) );
  NAND2_X1 U15180 ( .A1(n12752), .A2(n12751), .ZN(n14485) );
  NAND2_X1 U15181 ( .A1(n15064), .A2(n12846), .ZN(n12754) );
  NAND2_X1 U15182 ( .A1(n14705), .A2(n12849), .ZN(n12753) );
  NAND2_X1 U15183 ( .A1(n12754), .A2(n12753), .ZN(n12755) );
  XNOR2_X1 U15184 ( .A(n12755), .B(n10529), .ZN(n14487) );
  NAND2_X1 U15185 ( .A1(n15064), .A2(n12849), .ZN(n12757) );
  NAND2_X1 U15186 ( .A1(n14705), .A2(n12848), .ZN(n12756) );
  NAND2_X1 U15187 ( .A1(n12757), .A2(n12756), .ZN(n14486) );
  NOR2_X1 U15188 ( .A1(n14487), .A2(n14486), .ZN(n12759) );
  NAND2_X1 U15189 ( .A1(n14487), .A2(n14486), .ZN(n12758) );
  OAI22_X1 U15190 ( .A1(n14944), .A2(n12785), .B1(n14489), .B2(n12787), .ZN(
        n12760) );
  XNOR2_X1 U15191 ( .A(n12760), .B(n10529), .ZN(n12767) );
  OR2_X1 U15192 ( .A1(n14944), .A2(n12787), .ZN(n12762) );
  OR2_X1 U15193 ( .A1(n14489), .A2(n12788), .ZN(n12761) );
  NAND2_X1 U15194 ( .A1(n12762), .A2(n12761), .ZN(n12766) );
  XNOR2_X1 U15195 ( .A(n12767), .B(n12766), .ZN(n14531) );
  AOI22_X1 U15196 ( .A1(n15052), .A2(n12846), .B1(n12849), .B2(n14709), .ZN(
        n12764) );
  XNOR2_X1 U15197 ( .A(n12764), .B(n10529), .ZN(n12769) );
  AND2_X1 U15198 ( .A1(n14709), .A2(n12848), .ZN(n12765) );
  AOI21_X1 U15199 ( .B1(n15052), .B2(n12849), .A(n12765), .ZN(n12770) );
  XNOR2_X1 U15200 ( .A(n12769), .B(n12770), .ZN(n14455) );
  NOR2_X1 U15201 ( .A1(n12767), .A2(n12766), .ZN(n14456) );
  NOR2_X1 U15202 ( .A1(n14455), .A2(n14456), .ZN(n12768) );
  INV_X1 U15203 ( .A(n12770), .ZN(n12771) );
  NAND2_X1 U15204 ( .A1(n12772), .A2(n12771), .ZN(n12773) );
  OAI22_X1 U15205 ( .A1(n14911), .A2(n12787), .B1(n14710), .B2(n12788), .ZN(
        n12775) );
  OAI22_X1 U15206 ( .A1(n14911), .A2(n12785), .B1(n14710), .B2(n12787), .ZN(
        n12774) );
  XNOR2_X1 U15207 ( .A(n12774), .B(n10529), .ZN(n12776) );
  XOR2_X1 U15208 ( .A(n12775), .B(n12776), .Z(n14514) );
  NAND2_X1 U15209 ( .A1(n12776), .A2(n12775), .ZN(n12777) );
  NAND2_X1 U15210 ( .A1(n15041), .A2(n12846), .ZN(n12780) );
  NAND2_X1 U15211 ( .A1(n14712), .A2(n12849), .ZN(n12779) );
  NAND2_X1 U15212 ( .A1(n12780), .A2(n12779), .ZN(n12781) );
  XNOR2_X1 U15213 ( .A(n12781), .B(n7239), .ZN(n12784) );
  AND2_X1 U15214 ( .A1(n14712), .A2(n12848), .ZN(n12782) );
  AOI21_X1 U15215 ( .B1(n15041), .B2(n12849), .A(n12782), .ZN(n12783) );
  NAND2_X1 U15216 ( .A1(n12784), .A2(n12783), .ZN(n14525) );
  OAI21_X1 U15217 ( .B1(n12784), .B2(n12783), .A(n14525), .ZN(n14465) );
  OAI22_X1 U15218 ( .A1(n14884), .A2(n12785), .B1(n14714), .B2(n12787), .ZN(
        n12786) );
  XNOR2_X1 U15219 ( .A(n12786), .B(n12819), .ZN(n12791) );
  OR2_X1 U15220 ( .A1(n14884), .A2(n12787), .ZN(n12790) );
  OR2_X1 U15221 ( .A1(n14714), .A2(n12788), .ZN(n12789) );
  AND2_X1 U15222 ( .A1(n12790), .A2(n12789), .ZN(n12792) );
  NAND2_X1 U15223 ( .A1(n12791), .A2(n12792), .ZN(n14450) );
  INV_X1 U15224 ( .A(n12791), .ZN(n12794) );
  INV_X1 U15225 ( .A(n12792), .ZN(n12793) );
  NAND2_X1 U15226 ( .A1(n12794), .A2(n12793), .ZN(n12795) );
  AND2_X1 U15227 ( .A1(n14450), .A2(n12795), .ZN(n14523) );
  NAND2_X1 U15228 ( .A1(n12796), .A2(n14523), .ZN(n14447) );
  NAND2_X1 U15229 ( .A1(n14447), .A2(n14450), .ZN(n12806) );
  NAND2_X1 U15230 ( .A1(n15024), .A2(n12846), .ZN(n12798) );
  NAND2_X1 U15231 ( .A1(n14717), .A2(n12849), .ZN(n12797) );
  NAND2_X1 U15232 ( .A1(n12798), .A2(n12797), .ZN(n12799) );
  XNOR2_X1 U15233 ( .A(n12799), .B(n12819), .ZN(n12801) );
  AND2_X1 U15234 ( .A1(n14717), .A2(n12848), .ZN(n12800) );
  AOI21_X1 U15235 ( .B1(n15024), .B2(n12849), .A(n12800), .ZN(n12802) );
  NAND2_X1 U15236 ( .A1(n12801), .A2(n12802), .ZN(n14495) );
  INV_X1 U15237 ( .A(n12801), .ZN(n12804) );
  INV_X1 U15238 ( .A(n12802), .ZN(n12803) );
  NAND2_X1 U15239 ( .A1(n12804), .A2(n12803), .ZN(n12805) );
  NAND2_X1 U15240 ( .A1(n12806), .A2(n14448), .ZN(n14446) );
  NAND2_X1 U15241 ( .A1(n14446), .A2(n14495), .ZN(n12816) );
  NAND2_X1 U15242 ( .A1(n14859), .A2(n12846), .ZN(n12808) );
  NAND2_X1 U15243 ( .A1(n14826), .A2(n12849), .ZN(n12807) );
  NAND2_X1 U15244 ( .A1(n12808), .A2(n12807), .ZN(n12809) );
  XNOR2_X1 U15245 ( .A(n12809), .B(n12819), .ZN(n12811) );
  AND2_X1 U15246 ( .A1(n14826), .A2(n12848), .ZN(n12810) );
  AOI21_X1 U15247 ( .B1(n14859), .B2(n12849), .A(n12810), .ZN(n12812) );
  NAND2_X1 U15248 ( .A1(n12811), .A2(n12812), .ZN(n14472) );
  INV_X1 U15249 ( .A(n12811), .ZN(n12814) );
  INV_X1 U15250 ( .A(n12812), .ZN(n12813) );
  NAND2_X1 U15251 ( .A1(n12814), .A2(n12813), .ZN(n12815) );
  NAND2_X1 U15252 ( .A1(n12816), .A2(n14497), .ZN(n14475) );
  NAND2_X1 U15253 ( .A1(n14475), .A2(n14472), .ZN(n12827) );
  NAND2_X1 U15254 ( .A1(n15014), .A2(n12846), .ZN(n12818) );
  NAND2_X1 U15255 ( .A1(n14720), .A2(n12849), .ZN(n12817) );
  NAND2_X1 U15256 ( .A1(n12818), .A2(n12817), .ZN(n12820) );
  XNOR2_X1 U15257 ( .A(n12820), .B(n12819), .ZN(n12822) );
  AND2_X1 U15258 ( .A1(n14720), .A2(n12848), .ZN(n12821) );
  AOI21_X1 U15259 ( .B1(n15014), .B2(n12849), .A(n12821), .ZN(n12823) );
  NAND2_X1 U15260 ( .A1(n12822), .A2(n12823), .ZN(n12828) );
  INV_X1 U15261 ( .A(n12822), .ZN(n12825) );
  INV_X1 U15262 ( .A(n12823), .ZN(n12824) );
  NAND2_X1 U15263 ( .A1(n12825), .A2(n12824), .ZN(n12826) );
  NAND2_X1 U15264 ( .A1(n12827), .A2(n14474), .ZN(n14476) );
  NAND2_X1 U15265 ( .A1(n14476), .A2(n12828), .ZN(n14540) );
  NAND2_X1 U15266 ( .A1(n14762), .A2(n12846), .ZN(n12830) );
  NAND2_X1 U15267 ( .A1(n14828), .A2(n12849), .ZN(n12829) );
  NAND2_X1 U15268 ( .A1(n12830), .A2(n12829), .ZN(n12831) );
  XNOR2_X1 U15269 ( .A(n12831), .B(n10529), .ZN(n12835) );
  NAND2_X1 U15270 ( .A1(n14762), .A2(n12849), .ZN(n12833) );
  NAND2_X1 U15271 ( .A1(n14828), .A2(n12848), .ZN(n12832) );
  NAND2_X1 U15272 ( .A1(n12833), .A2(n12832), .ZN(n12834) );
  NOR2_X1 U15273 ( .A1(n12835), .A2(n12834), .ZN(n12836) );
  AOI21_X1 U15274 ( .B1(n12835), .B2(n12834), .A(n12836), .ZN(n14541) );
  INV_X1 U15275 ( .A(n12836), .ZN(n12837) );
  NAND2_X1 U15276 ( .A1(n14802), .A2(n12846), .ZN(n12839) );
  NAND2_X1 U15277 ( .A1(n14764), .A2(n12849), .ZN(n12838) );
  NAND2_X1 U15278 ( .A1(n12839), .A2(n12838), .ZN(n12840) );
  XNOR2_X1 U15279 ( .A(n12840), .B(n10529), .ZN(n12844) );
  NAND2_X1 U15280 ( .A1(n14802), .A2(n12849), .ZN(n12842) );
  NAND2_X1 U15281 ( .A1(n14764), .A2(n12848), .ZN(n12841) );
  NAND2_X1 U15282 ( .A1(n12842), .A2(n12841), .ZN(n12843) );
  NOR2_X1 U15283 ( .A1(n12844), .A2(n12843), .ZN(n12845) );
  AOI21_X1 U15284 ( .B1(n12844), .B2(n12843), .A(n12845), .ZN(n14436) );
  AOI22_X1 U15285 ( .A1(n14779), .A2(n12846), .B1(n12849), .B2(n14789), .ZN(
        n12847) );
  XNOR2_X1 U15286 ( .A(n12847), .B(n10529), .ZN(n12851) );
  AOI22_X1 U15287 ( .A1(n14779), .A2(n12849), .B1(n12848), .B2(n14789), .ZN(
        n12850) );
  XNOR2_X1 U15288 ( .A(n12851), .B(n12850), .ZN(n12852) );
  OR2_X1 U15289 ( .A1(n12853), .A2(n14967), .ZN(n12855) );
  NAND2_X1 U15290 ( .A1(n14764), .A2(n14825), .ZN(n12854) );
  NAND2_X1 U15291 ( .A1(n12855), .A2(n12854), .ZN(n14774) );
  AOI22_X1 U15292 ( .A1(n15348), .A2(n14774), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12856) );
  OAI21_X1 U15293 ( .B1(n14775), .B2(n15369), .A(n12856), .ZN(n12857) );
  AOI21_X1 U15294 ( .B1(n14779), .B2(n15351), .A(n12857), .ZN(n12858) );
  OAI21_X1 U15295 ( .B1(n12859), .B2(n15337), .A(n12858), .ZN(P1_U3220) );
  INV_X1 U15296 ( .A(n12860), .ZN(n14413) );
  OAI222_X1 U15297 ( .A1(P1_U3086), .A2(n9904), .B1(n15104), .B2(n14413), .C1(
        n12861), .C2(n15101), .ZN(P1_U3326) );
  XNOR2_X1 U15298 ( .A(n13407), .B(n12862), .ZN(n12870) );
  INV_X1 U15299 ( .A(n12870), .ZN(n12863) );
  NAND2_X1 U15300 ( .A1(n12863), .A2(n13023), .ZN(n12875) );
  INV_X1 U15301 ( .A(n12864), .ZN(n12865) );
  AOI22_X1 U15302 ( .A1(n12868), .A2(n13014), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12867) );
  NAND2_X1 U15303 ( .A1(n13416), .A2(n13031), .ZN(n12866) );
  OAI211_X1 U15304 ( .C1(n13411), .C2(n13016), .A(n12867), .B(n12866), .ZN(
        n12872) );
  NOR4_X1 U15305 ( .A1(n12870), .A2(n12869), .A3(n12868), .A4(n13008), .ZN(
        n12871) );
  AOI211_X1 U15306 ( .C1(n13006), .C2(n13415), .A(n12872), .B(n12871), .ZN(
        n12873) );
  OR2_X1 U15307 ( .A1(n12876), .A2(n12877), .ZN(n12880) );
  NAND2_X1 U15308 ( .A1(n12880), .A2(n12878), .ZN(n12881) );
  AND2_X1 U15309 ( .A1(n12880), .A2(n12879), .ZN(n13021) );
  AOI21_X1 U15310 ( .B1(n12882), .B2(n12881), .A(n13021), .ZN(n12889) );
  NOR2_X1 U15311 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12883), .ZN(n13290) );
  AOI21_X1 U15312 ( .B1(n13026), .B2(n15173), .A(n13290), .ZN(n12884) );
  OAI21_X1 U15313 ( .B1(n12885), .B2(n13028), .A(n12884), .ZN(n12887) );
  NOR2_X1 U15314 ( .A1(n15178), .A2(n13035), .ZN(n12886) );
  AOI211_X1 U15315 ( .C1(n15175), .C2(n13031), .A(n12887), .B(n12886), .ZN(
        n12888) );
  OAI21_X1 U15316 ( .B1(n12889), .B2(n13008), .A(n12888), .ZN(P3_U3155) );
  INV_X1 U15317 ( .A(n12890), .ZN(n12891) );
  AOI21_X1 U15318 ( .B1(n12893), .B2(n12892), .A(n12891), .ZN(n12900) );
  NAND2_X1 U15319 ( .A1(n13031), .A2(n13537), .ZN(n12896) );
  NOR2_X1 U15320 ( .A1(n12894), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13391) );
  AOI21_X1 U15321 ( .B1(n13026), .B2(n13532), .A(n13391), .ZN(n12895) );
  OAI211_X1 U15322 ( .C1(n12897), .C2(n13028), .A(n12896), .B(n12895), .ZN(
        n12898) );
  AOI21_X1 U15323 ( .B1(n13671), .B2(n13006), .A(n12898), .ZN(n12899) );
  OAI21_X1 U15324 ( .B1(n12900), .B2(n13008), .A(n12899), .ZN(P3_U3159) );
  INV_X1 U15325 ( .A(n12901), .ZN(n12902) );
  AOI21_X1 U15326 ( .B1(n12904), .B2(n12903), .A(n12902), .ZN(n12909) );
  NAND2_X1 U15327 ( .A1(n13031), .A2(n13511), .ZN(n12906) );
  AOI22_X1 U15328 ( .A1(n13026), .A2(n13482), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12905) );
  OAI211_X1 U15329 ( .C1(n13508), .C2(n13028), .A(n12906), .B(n12905), .ZN(
        n12907) );
  AOI21_X1 U15330 ( .B1(n13086), .B2(n13006), .A(n12907), .ZN(n12908) );
  OAI21_X1 U15331 ( .B1(n12909), .B2(n13008), .A(n12908), .ZN(P3_U3163) );
  INV_X1 U15332 ( .A(n12911), .ZN(n12912) );
  AOI21_X1 U15333 ( .B1(n12913), .B2(n12910), .A(n12912), .ZN(n12919) );
  NOR2_X1 U15334 ( .A1(n13028), .A2(n12991), .ZN(n12914) );
  AOI211_X1 U15335 ( .C1(n13026), .C2(n15199), .A(n12915), .B(n12914), .ZN(
        n12916) );
  OAI21_X1 U15336 ( .B1(n15204), .B2(n13035), .A(n12916), .ZN(n12917) );
  AOI21_X1 U15337 ( .B1(n15201), .B2(n13031), .A(n12917), .ZN(n12918) );
  OAI21_X1 U15338 ( .B1(n12919), .B2(n13008), .A(n12918), .ZN(P3_U3164) );
  NAND2_X1 U15339 ( .A1(n12922), .A2(n12921), .ZN(n12955) );
  INV_X1 U15340 ( .A(n12923), .ZN(n12925) );
  NOR3_X1 U15341 ( .A1(n12955), .A2(n12925), .A3(n12924), .ZN(n12928) );
  INV_X1 U15342 ( .A(n12926), .ZN(n12927) );
  OAI21_X1 U15343 ( .B1(n12928), .B2(n12927), .A(n13023), .ZN(n12933) );
  INV_X1 U15344 ( .A(n13453), .ZN(n12929) );
  NOR2_X1 U15345 ( .A1(n12929), .A2(n12958), .ZN(n12931) );
  OAI22_X1 U15346 ( .A1(n13448), .A2(n13016), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9525), .ZN(n12930) );
  AOI211_X1 U15347 ( .C1(n13014), .C2(n13483), .A(n12931), .B(n12930), .ZN(
        n12932) );
  OAI211_X1 U15348 ( .C1(n13651), .C2(n13035), .A(n12933), .B(n12932), .ZN(
        P3_U3165) );
  XNOR2_X1 U15349 ( .A(n12934), .B(n12935), .ZN(n12941) );
  NAND2_X1 U15350 ( .A1(n13031), .A2(n13581), .ZN(n12938) );
  NOR2_X1 U15351 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12936), .ZN(n13316) );
  AOI21_X1 U15352 ( .B1(n13026), .B2(n13574), .A(n13316), .ZN(n12937) );
  OAI211_X1 U15353 ( .C1(n13180), .C2(n13028), .A(n12938), .B(n12937), .ZN(
        n12939) );
  AOI21_X1 U15354 ( .B1(n13681), .B2(n13006), .A(n12939), .ZN(n12940) );
  OAI21_X1 U15355 ( .B1(n12941), .B2(n13008), .A(n12940), .ZN(P3_U3166) );
  XNOR2_X1 U15356 ( .A(n12942), .B(n12943), .ZN(n12950) );
  INV_X1 U15357 ( .A(n13568), .ZN(n13627) );
  NAND2_X1 U15358 ( .A1(n13031), .A2(n13566), .ZN(n12946) );
  NOR2_X1 U15359 ( .A1(n12944), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13338) );
  AOI21_X1 U15360 ( .B1(n13026), .B2(n13560), .A(n13338), .ZN(n12945) );
  OAI211_X1 U15361 ( .C1(n12947), .C2(n13028), .A(n12946), .B(n12945), .ZN(
        n12948) );
  AOI21_X1 U15362 ( .B1(n13627), .B2(n13006), .A(n12948), .ZN(n12949) );
  OAI21_X1 U15363 ( .B1(n12950), .B2(n13008), .A(n12949), .ZN(P3_U3168) );
  INV_X1 U15364 ( .A(n12952), .ZN(n12954) );
  NOR3_X1 U15365 ( .A1(n7769), .A2(n12954), .A3(n12953), .ZN(n12956) );
  OAI21_X1 U15366 ( .B1(n12956), .B2(n12955), .A(n13023), .ZN(n12963) );
  INV_X1 U15367 ( .A(n13471), .ZN(n12957) );
  NOR2_X1 U15368 ( .A1(n12958), .A2(n12957), .ZN(n12961) );
  OAI22_X1 U15369 ( .A1(n13433), .A2(n13016), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12959), .ZN(n12960) );
  AOI211_X1 U15370 ( .C1(n13014), .C2(n13466), .A(n12961), .B(n12960), .ZN(
        n12962) );
  OAI211_X1 U15371 ( .C1(n13655), .C2(n13035), .A(n12963), .B(n12962), .ZN(
        P3_U3169) );
  NAND2_X1 U15372 ( .A1(n12890), .A2(n12964), .ZN(n12966) );
  AOI21_X1 U15373 ( .B1(n12966), .B2(n12965), .A(n13008), .ZN(n12968) );
  NAND2_X1 U15374 ( .A1(n12968), .A2(n12967), .ZN(n12972) );
  AOI22_X1 U15375 ( .A1(n13026), .A2(n13519), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12969) );
  OAI21_X1 U15376 ( .B1(n13547), .B2(n13028), .A(n12969), .ZN(n12970) );
  AOI21_X1 U15377 ( .B1(n13526), .B2(n13031), .A(n12970), .ZN(n12971) );
  OAI211_X1 U15378 ( .C1(n13528), .C2(n13035), .A(n12972), .B(n12971), .ZN(
        P3_U3173) );
  XNOR2_X1 U15379 ( .A(n12973), .B(n15199), .ZN(n12974) );
  XNOR2_X1 U15380 ( .A(n12876), .B(n12974), .ZN(n12981) );
  NOR2_X1 U15381 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12975), .ZN(n13253) );
  AOI21_X1 U15382 ( .B1(n13026), .B2(n15187), .A(n13253), .ZN(n12976) );
  OAI21_X1 U15383 ( .B1(n12994), .B2(n13028), .A(n12976), .ZN(n12978) );
  NOR2_X1 U15384 ( .A1(n15194), .A2(n13035), .ZN(n12977) );
  AOI211_X1 U15385 ( .C1(n12979), .C2(n13031), .A(n12978), .B(n12977), .ZN(
        n12980) );
  OAI21_X1 U15386 ( .B1(n12981), .B2(n13008), .A(n12980), .ZN(P3_U3174) );
  AOI21_X1 U15387 ( .B1(n13482), .B2(n12982), .A(n6728), .ZN(n12987) );
  NAND2_X1 U15388 ( .A1(n13031), .A2(n13500), .ZN(n12984) );
  AOI22_X1 U15389 ( .A1(n13026), .A2(n13466), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12983) );
  OAI211_X1 U15390 ( .C1(n13496), .C2(n13028), .A(n12984), .B(n12983), .ZN(
        n12985) );
  AOI21_X1 U15391 ( .B1(n13499), .B2(n13006), .A(n12985), .ZN(n12986) );
  OAI21_X1 U15392 ( .B1(n12987), .B2(n13008), .A(n12986), .ZN(P3_U3175) );
  INV_X1 U15393 ( .A(n12988), .ZN(n12990) );
  NAND2_X1 U15394 ( .A1(n12990), .A2(n12989), .ZN(n12992) );
  XNOR2_X1 U15395 ( .A(n12992), .B(n12991), .ZN(n12999) );
  NOR2_X1 U15396 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12993), .ZN(n15750) );
  NOR2_X1 U15397 ( .A1(n13016), .A2(n12994), .ZN(n12995) );
  AOI211_X1 U15398 ( .C1(n13014), .C2(n15208), .A(n15750), .B(n12995), .ZN(
        n12996) );
  OAI21_X1 U15399 ( .B1(n15216), .B2(n13035), .A(n12996), .ZN(n12997) );
  AOI21_X1 U15400 ( .B1(n15212), .B2(n13031), .A(n12997), .ZN(n12998) );
  OAI21_X1 U15401 ( .B1(n12999), .B2(n13008), .A(n12998), .ZN(P3_U3176) );
  XNOR2_X1 U15402 ( .A(n13000), .B(n13001), .ZN(n13009) );
  NAND2_X1 U15403 ( .A1(n13031), .A2(n13551), .ZN(n13004) );
  NOR2_X1 U15404 ( .A1(n13002), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13368) );
  AOI21_X1 U15405 ( .B1(n13026), .B2(n13518), .A(n13368), .ZN(n13003) );
  OAI211_X1 U15406 ( .C1(n13546), .C2(n13028), .A(n13004), .B(n13003), .ZN(
        n13005) );
  AOI21_X1 U15407 ( .B1(n13550), .B2(n13006), .A(n13005), .ZN(n13007) );
  OAI21_X1 U15408 ( .B1(n13009), .B2(n13008), .A(n13007), .ZN(P3_U3178) );
  AOI22_X1 U15409 ( .A1(n13467), .A2(n13014), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13015) );
  OAI21_X1 U15410 ( .B1(n13434), .B2(n13016), .A(n13015), .ZN(n13017) );
  AOI21_X1 U15411 ( .B1(n13438), .B2(n13031), .A(n13017), .ZN(n13018) );
  OAI21_X1 U15412 ( .B1(n13021), .B2(n13020), .A(n13019), .ZN(n13024) );
  NAND3_X1 U15413 ( .A1(n13024), .A2(n13023), .A3(n13022), .ZN(n13034) );
  NOR2_X1 U15414 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13025), .ZN(n15157) );
  AOI21_X1 U15415 ( .B1(n13026), .B2(n13559), .A(n15157), .ZN(n13027) );
  OAI21_X1 U15416 ( .B1(n13029), .B2(n13028), .A(n13027), .ZN(n13030) );
  AOI21_X1 U15417 ( .B1(n13032), .B2(n13031), .A(n13030), .ZN(n13033) );
  OAI211_X1 U15418 ( .C1(n13035), .C2(n13179), .A(n13034), .B(n13033), .ZN(
        P3_U3181) );
  OAI22_X1 U15419 ( .A1(n13040), .A2(n13038), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13047) );
  OAI21_X1 U15420 ( .B1(n13040), .B2(P1_DATAO_REG_30__SCAN_IN), .A(n13039), 
        .ZN(n13043) );
  AOI22_X1 U15421 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(
        P1_DATAO_REG_31__SCAN_IN), .B1(n13041), .B2(n15087), .ZN(n13042) );
  XOR2_X1 U15422 ( .A(n13043), .B(n13042), .Z(n13687) );
  NAND2_X1 U15423 ( .A1(n13687), .A2(n6677), .ZN(n13046) );
  INV_X1 U15424 ( .A(SI_31_), .ZN(n13692) );
  OR2_X1 U15425 ( .A1(n13044), .A2(n13692), .ZN(n13045) );
  INV_X1 U15426 ( .A(n13057), .ZN(n13058) );
  XOR2_X1 U15427 ( .A(n13048), .B(n13047), .Z(n13694) );
  OR2_X1 U15428 ( .A1(n13044), .A2(n13693), .ZN(n13049) );
  OAI21_X1 U15429 ( .B1(n13694), .B2(n13050), .A(n13049), .ZN(n15167) );
  NOR2_X1 U15430 ( .A1(n13053), .A2(n13411), .ZN(n13232) );
  INV_X1 U15431 ( .A(n15167), .ZN(n15223) );
  OAI22_X1 U15432 ( .A1(n15223), .A2(n13052), .B1(n13057), .B2(n15161), .ZN(
        n13234) );
  INV_X1 U15433 ( .A(n13234), .ZN(n13055) );
  AND2_X1 U15434 ( .A1(n13053), .A2(n13411), .ZN(n13231) );
  AOI21_X1 U15435 ( .B1(n15167), .B2(n15161), .A(n13231), .ZN(n13054) );
  NAND2_X1 U15436 ( .A1(n13057), .A2(n15161), .ZN(n13233) );
  XNOR2_X1 U15437 ( .A(n13086), .B(n13496), .ZN(n13510) );
  NAND2_X1 U15438 ( .A1(n13205), .A2(n13202), .ZN(n13497) );
  INV_X1 U15439 ( .A(n13535), .ZN(n13073) );
  NAND4_X1 U15440 ( .A1(n13060), .A2(n13059), .A3(n15785), .A4(n13124), .ZN(
        n13065) );
  NAND4_X1 U15441 ( .A1(n15804), .A2(n13063), .A3(n13062), .A4(n13061), .ZN(
        n13064) );
  NOR3_X1 U15442 ( .A1(n13065), .A2(n13064), .A3(n13144), .ZN(n13069) );
  INV_X1 U15443 ( .A(n13151), .ZN(n13067) );
  NAND2_X1 U15444 ( .A1(n13067), .A2(n13066), .ZN(n13160) );
  INV_X1 U15445 ( .A(n13160), .ZN(n13068) );
  NAND4_X1 U15446 ( .A1(n13069), .A2(n15214), .A3(n15202), .A4(n13068), .ZN(
        n13070) );
  OR3_X1 U15447 ( .A1(n15176), .A2(n15193), .A3(n13070), .ZN(n13071) );
  NOR4_X1 U15448 ( .A1(n13094), .A2(n13176), .A3(n8240), .A4(n13071), .ZN(
        n13072) );
  NAND4_X1 U15449 ( .A1(n13196), .A2(n13564), .A3(n13073), .A4(n13072), .ZN(
        n13074) );
  NOR4_X1 U15450 ( .A1(n13510), .A2(n13497), .A3(n13481), .A4(n13074), .ZN(
        n13075) );
  NAND4_X1 U15451 ( .A1(n13214), .A2(n13432), .A3(n13075), .A4(n13459), .ZN(
        n13076) );
  NOR2_X1 U15452 ( .A1(n13077), .A2(n13076), .ZN(n13078) );
  NAND4_X1 U15453 ( .A1(n6725), .A2(n13407), .A3(n13078), .A4(n13233), .ZN(
        n13080) );
  XNOR2_X1 U15454 ( .A(n13082), .B(n13081), .ZN(n13237) );
  XNOR2_X1 U15455 ( .A(n13083), .B(n13228), .ZN(n13212) );
  OR2_X1 U15456 ( .A1(n13496), .A2(n13221), .ZN(n13085) );
  NAND3_X1 U15457 ( .A1(n13086), .A2(n13496), .A3(n13221), .ZN(n13084) );
  OAI21_X1 U15458 ( .B1(n13086), .B2(n13085), .A(n13084), .ZN(n13087) );
  NOR2_X1 U15459 ( .A1(n13497), .A2(n13087), .ZN(n13201) );
  INV_X1 U15460 ( .A(n13510), .ZN(n13200) );
  OAI21_X1 U15461 ( .B1(n13546), .B2(n13627), .A(n13088), .ZN(n13089) );
  NAND2_X1 U15462 ( .A1(n13089), .A2(n13092), .ZN(n13090) );
  NAND2_X1 U15463 ( .A1(n13091), .A2(n13090), .ZN(n13096) );
  OAI211_X1 U15464 ( .C1(n13094), .C2(n13093), .A(n13191), .B(n13092), .ZN(
        n13095) );
  MUX2_X1 U15465 ( .A(n13096), .B(n13095), .S(n13228), .Z(n13097) );
  INV_X1 U15466 ( .A(n13097), .ZN(n13195) );
  MUX2_X1 U15467 ( .A(n13100), .B(n13098), .S(n13228), .Z(n13107) );
  NAND2_X1 U15468 ( .A1(n13099), .A2(n13243), .ZN(n13103) );
  NAND2_X1 U15469 ( .A1(n13099), .A2(n13105), .ZN(n13101) );
  NAND3_X1 U15470 ( .A1(n13101), .A2(n13228), .A3(n13100), .ZN(n13102) );
  OAI21_X1 U15471 ( .B1(n11259), .B2(n13103), .A(n13102), .ZN(n13104) );
  OAI21_X1 U15472 ( .B1(n13105), .B2(n15803), .A(n13104), .ZN(n13106) );
  NAND2_X1 U15473 ( .A1(n13115), .A2(n13108), .ZN(n13109) );
  NAND2_X1 U15474 ( .A1(n13109), .A2(n13228), .ZN(n13110) );
  NAND2_X1 U15475 ( .A1(n13112), .A2(n13111), .ZN(n13113) );
  NAND2_X1 U15476 ( .A1(n13113), .A2(n13221), .ZN(n13114) );
  NOR2_X1 U15477 ( .A1(n13115), .A2(n13228), .ZN(n13117) );
  NOR2_X1 U15478 ( .A1(n13117), .A2(n13116), .ZN(n13118) );
  NAND2_X1 U15479 ( .A1(n13119), .A2(n13118), .ZN(n13125) );
  NAND3_X1 U15480 ( .A1(n13125), .A2(n13124), .A3(n13120), .ZN(n13122) );
  NAND3_X1 U15481 ( .A1(n13122), .A2(n13127), .A3(n13121), .ZN(n13132) );
  NAND3_X1 U15482 ( .A1(n13125), .A2(n13124), .A3(n13123), .ZN(n13130) );
  AND2_X1 U15483 ( .A1(n13133), .A2(n13126), .ZN(n13129) );
  INV_X1 U15484 ( .A(n13127), .ZN(n13128) );
  AOI21_X1 U15485 ( .B1(n13130), .B2(n13129), .A(n13128), .ZN(n13131) );
  NOR2_X1 U15486 ( .A1(n13133), .A2(n13228), .ZN(n13135) );
  NOR2_X1 U15487 ( .A1(n13135), .A2(n13134), .ZN(n13141) );
  INV_X1 U15488 ( .A(n13136), .ZN(n13139) );
  INV_X1 U15489 ( .A(n13137), .ZN(n13138) );
  MUX2_X1 U15490 ( .A(n13139), .B(n13138), .S(n13221), .Z(n13140) );
  AOI21_X1 U15491 ( .B1(n13142), .B2(n13141), .A(n13140), .ZN(n13146) );
  XNOR2_X1 U15492 ( .A(n13143), .B(n13221), .ZN(n13145) );
  MUX2_X1 U15493 ( .A(n13146), .B(n13145), .S(n13144), .Z(n13161) );
  MUX2_X1 U15494 ( .A(n13221), .B(n13148), .S(n13147), .Z(n13150) );
  NAND2_X1 U15495 ( .A1(n13150), .A2(n13149), .ZN(n13152) );
  OAI21_X1 U15496 ( .B1(n13152), .B2(n13151), .A(n15214), .ZN(n13158) );
  INV_X1 U15497 ( .A(n13153), .ZN(n13156) );
  INV_X1 U15498 ( .A(n13154), .ZN(n13155) );
  MUX2_X1 U15499 ( .A(n13156), .B(n13155), .S(n13221), .Z(n13157) );
  NOR2_X1 U15500 ( .A1(n13158), .A2(n13157), .ZN(n13159) );
  NAND2_X1 U15501 ( .A1(n13166), .A2(n13162), .ZN(n13163) );
  NAND2_X1 U15502 ( .A1(n13163), .A2(n13228), .ZN(n13164) );
  AOI21_X1 U15503 ( .B1(n6792), .B2(n13165), .A(n13228), .ZN(n13169) );
  NOR2_X1 U15504 ( .A1(n13166), .A2(n13228), .ZN(n13167) );
  NOR2_X1 U15505 ( .A1(n15193), .A2(n13167), .ZN(n13168) );
  MUX2_X1 U15506 ( .A(n13171), .B(n13170), .S(n13221), .Z(n13172) );
  INV_X1 U15507 ( .A(n13173), .ZN(n13174) );
  MUX2_X1 U15508 ( .A(n13175), .B(n13174), .S(n13228), .Z(n13177) );
  OR3_X1 U15509 ( .A1(n13178), .A2(n13177), .A3(n13176), .ZN(n13184) );
  INV_X1 U15510 ( .A(n13179), .ZN(n13637) );
  OAI21_X1 U15511 ( .B1(n13180), .B2(n13637), .A(n13187), .ZN(n13181) );
  NAND2_X1 U15512 ( .A1(n13181), .A2(n13228), .ZN(n13183) );
  AOI21_X1 U15513 ( .B1(n13184), .B2(n13183), .A(n13182), .ZN(n13189) );
  AOI21_X1 U15514 ( .B1(n13186), .B2(n13185), .A(n13228), .ZN(n13188) );
  OAI22_X1 U15515 ( .A1(n13189), .A2(n13188), .B1(n13228), .B2(n13187), .ZN(
        n13190) );
  INV_X1 U15516 ( .A(n13191), .ZN(n13193) );
  MUX2_X1 U15517 ( .A(n13193), .B(n13192), .S(n13228), .Z(n13194) );
  MUX2_X1 U15518 ( .A(n13198), .B(n13197), .S(n13221), .Z(n13199) );
  INV_X1 U15519 ( .A(n13202), .ZN(n13203) );
  NOR2_X1 U15520 ( .A1(n13481), .A2(n13203), .ZN(n13204) );
  AND2_X1 U15521 ( .A1(n13206), .A2(n13204), .ZN(n13210) );
  NAND3_X1 U15522 ( .A1(n13206), .A2(n13476), .A3(n13205), .ZN(n13208) );
  NAND2_X1 U15523 ( .A1(n13208), .A2(n13207), .ZN(n13209) );
  MUX2_X1 U15524 ( .A(n13210), .B(n13209), .S(n13221), .Z(n13211) );
  NAND3_X1 U15525 ( .A1(n13432), .A2(n13218), .A3(n13217), .ZN(n13220) );
  NAND2_X1 U15526 ( .A1(n13220), .A2(n13219), .ZN(n13222) );
  OAI21_X1 U15527 ( .B1(n13226), .B2(n13228), .A(n13225), .ZN(n13227) );
  INV_X1 U15528 ( .A(n13407), .ZN(n13229) );
  NAND3_X1 U15529 ( .A1(n13241), .A2(n13240), .A3(n10612), .ZN(n13242) );
  OAI211_X1 U15530 ( .C1(n13243), .C2(n13245), .A(n13242), .B(P3_B_REG_SCAN_IN), .ZN(n13244) );
  MUX2_X1 U15531 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n13519), .S(P3_U3897), .Z(
        P3_U3512) );
  NAND2_X1 U15532 ( .A1(n13255), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n13246) );
  AOI21_X1 U15533 ( .B1(n8048), .B2(n13248), .A(n13268), .ZN(n13266) );
  AOI21_X1 U15534 ( .B1(n13250), .B2(n13255), .A(n13249), .ZN(n13252) );
  MUX2_X1 U15535 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n10612), .Z(n13280) );
  XNOR2_X1 U15536 ( .A(n13280), .B(n13281), .ZN(n13251) );
  NAND2_X1 U15537 ( .A1(n13252), .A2(n13251), .ZN(n13287) );
  OAI21_X1 U15538 ( .B1(n13252), .B2(n13251), .A(n13287), .ZN(n13264) );
  AOI21_X1 U15539 ( .B1(n15732), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n13253), 
        .ZN(n13254) );
  OAI21_X1 U15540 ( .B1(n15738), .B2(n15124), .A(n13254), .ZN(n13263) );
  INV_X1 U15541 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n15190) );
  NAND2_X1 U15542 ( .A1(n13255), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n13256) );
  AOI21_X1 U15543 ( .B1(n15190), .B2(n13260), .A(n13277), .ZN(n13261) );
  NOR2_X1 U15544 ( .A1(n13261), .A2(n15752), .ZN(n13262) );
  AOI211_X1 U15545 ( .C1(n13395), .C2(n13264), .A(n13263), .B(n13262), .ZN(
        n13265) );
  OAI21_X1 U15546 ( .B1(n13266), .B2(n15744), .A(n13265), .ZN(P3_U3195) );
  OR2_X1 U15547 ( .A1(n13270), .A2(n13269), .ZN(n13319) );
  NAND2_X1 U15548 ( .A1(n13270), .A2(n13269), .ZN(n13271) );
  AND2_X1 U15549 ( .A1(n13319), .A2(n13271), .ZN(n13284) );
  INV_X1 U15550 ( .A(n13284), .ZN(n13273) );
  INV_X1 U15551 ( .A(n13318), .ZN(n13272) );
  AOI21_X1 U15552 ( .B1(n13274), .B2(n13273), .A(n13272), .ZN(n13297) );
  NOR2_X1 U15553 ( .A1(n13281), .A2(n13275), .ZN(n13276) );
  NAND2_X1 U15554 ( .A1(n13293), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n13304) );
  OAI21_X1 U15555 ( .B1(n13293), .B2(P3_REG2_REG_14__SCAN_IN), .A(n13304), 
        .ZN(n13283) );
  AOI21_X1 U15556 ( .B1(n13278), .B2(n13283), .A(n13298), .ZN(n13279) );
  NOR2_X1 U15557 ( .A1(n13279), .A2(n15752), .ZN(n13295) );
  INV_X1 U15558 ( .A(n13280), .ZN(n13282) );
  NAND2_X1 U15559 ( .A1(n13282), .A2(n13281), .ZN(n13286) );
  AND2_X1 U15560 ( .A1(n13287), .A2(n13286), .ZN(n13289) );
  INV_X1 U15561 ( .A(n13283), .ZN(n13285) );
  MUX2_X1 U15562 ( .A(n13285), .B(n13284), .S(n10612), .Z(n13288) );
  NAND3_X1 U15563 ( .A1(n13287), .A2(n13286), .A3(n13288), .ZN(n13306) );
  OAI211_X1 U15564 ( .C1(n13289), .C2(n13288), .A(n13395), .B(n13306), .ZN(
        n13292) );
  AOI21_X1 U15565 ( .B1(n15732), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n13290), 
        .ZN(n13291) );
  OAI211_X1 U15566 ( .C1(n15738), .C2(n13293), .A(n13292), .B(n13291), .ZN(
        n13294) );
  NOR2_X1 U15567 ( .A1(n13295), .A2(n13294), .ZN(n13296) );
  OAI21_X1 U15568 ( .B1(n13297), .B2(n15744), .A(n13296), .ZN(P3_U3196) );
  XNOR2_X1 U15569 ( .A(n13333), .B(P3_REG2_REG_16__SCAN_IN), .ZN(n13303) );
  AND2_X1 U15570 ( .A1(n15146), .A2(n13299), .ZN(n13300) );
  INV_X1 U15571 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n15144) );
  NOR2_X1 U15572 ( .A1(n13300), .A2(n15142), .ZN(n13302) );
  INV_X1 U15573 ( .A(n13335), .ZN(n13301) );
  AOI21_X1 U15574 ( .B1(n13303), .B2(n13302), .A(n13301), .ZN(n13328) );
  MUX2_X1 U15575 ( .A(n13304), .B(n13319), .S(n10612), .Z(n13305) );
  NAND2_X1 U15576 ( .A1(n13306), .A2(n13305), .ZN(n13307) );
  INV_X1 U15577 ( .A(n13307), .ZN(n13309) );
  XNOR2_X1 U15578 ( .A(n13307), .B(n15146), .ZN(n15151) );
  MUX2_X1 U15579 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n10612), .Z(n15152) );
  AOI21_X1 U15580 ( .B1(n13309), .B2(n13308), .A(n15150), .ZN(n13343) );
  INV_X1 U15581 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13311) );
  MUX2_X1 U15582 ( .A(n13311), .B(n13310), .S(n10612), .Z(n13313) );
  INV_X1 U15583 ( .A(n13333), .ZN(n13312) );
  NOR2_X1 U15584 ( .A1(n13313), .A2(n13312), .ZN(n13342) );
  INV_X1 U15585 ( .A(n13342), .ZN(n13314) );
  NAND2_X1 U15586 ( .A1(n13313), .A2(n13312), .ZN(n13341) );
  NAND2_X1 U15587 ( .A1(n13314), .A2(n13341), .ZN(n13315) );
  XNOR2_X1 U15588 ( .A(n13343), .B(n13315), .ZN(n13326) );
  AOI21_X1 U15589 ( .B1(n15732), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n13316), 
        .ZN(n13317) );
  OAI21_X1 U15590 ( .B1(n15738), .B2(n13333), .A(n13317), .ZN(n13325) );
  XNOR2_X1 U15591 ( .A(n13333), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n13321) );
  NAND2_X1 U15592 ( .A1(n13322), .A2(n13321), .ZN(n13323) );
  AOI21_X1 U15593 ( .B1(n13330), .B2(n13323), .A(n15744), .ZN(n13324) );
  AOI211_X1 U15594 ( .C1(n13395), .C2(n13326), .A(n13325), .B(n13324), .ZN(
        n13327) );
  OAI21_X1 U15595 ( .B1(n13328), .B2(n15752), .A(n13327), .ZN(P3_U3198) );
  NAND2_X1 U15596 ( .A1(n13333), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n13329) );
  AOI21_X1 U15597 ( .B1(n13332), .B2(n13331), .A(n13352), .ZN(n13351) );
  NAND2_X1 U15598 ( .A1(n13333), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n13334) );
  INV_X1 U15599 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13336) );
  AOI21_X1 U15600 ( .B1(n13337), .B2(n13336), .A(n13360), .ZN(n13340) );
  AOI21_X1 U15601 ( .B1(n15732), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n13338), 
        .ZN(n13339) );
  OAI21_X1 U15602 ( .B1(n13340), .B2(n15752), .A(n13339), .ZN(n13347) );
  MUX2_X1 U15603 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n10612), .Z(n13356) );
  XNOR2_X1 U15604 ( .A(n13356), .B(n13361), .ZN(n13345) );
  OAI21_X1 U15605 ( .B1(n13343), .B2(n13342), .A(n13341), .ZN(n13344) );
  NOR2_X1 U15606 ( .A1(n13344), .A2(n13345), .ZN(n13355) );
  AOI211_X1 U15607 ( .C1(n13345), .C2(n13344), .A(n15746), .B(n13355), .ZN(
        n13346) );
  AOI211_X1 U15608 ( .C1(n13349), .C2(n13348), .A(n13347), .B(n13346), .ZN(
        n13350) );
  OAI21_X1 U15609 ( .B1(n13351), .B2(n15744), .A(n13350), .ZN(P3_U3199) );
  NAND2_X1 U15610 ( .A1(n13380), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n13375) );
  OAI21_X1 U15611 ( .B1(n13380), .B2(P3_REG1_REG_18__SCAN_IN), .A(n13375), 
        .ZN(n13354) );
  AOI21_X1 U15612 ( .B1(n6795), .B2(n13354), .A(n13377), .ZN(n13374) );
  MUX2_X1 U15613 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n10612), .Z(n13358) );
  XOR2_X1 U15614 ( .A(n13380), .B(n13383), .Z(n13357) );
  NOR2_X1 U15615 ( .A1(n13357), .A2(n13358), .ZN(n13381) );
  AOI21_X1 U15616 ( .B1(n13358), .B2(n13357), .A(n13381), .ZN(n13359) );
  INV_X1 U15617 ( .A(n13359), .ZN(n13372) );
  NAND2_X1 U15618 ( .A1(n13380), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n13387) );
  OAI21_X1 U15619 ( .B1(n13380), .B2(P3_REG2_REG_18__SCAN_IN), .A(n13387), 
        .ZN(n13365) );
  NAND2_X1 U15620 ( .A1(n13366), .A2(n13365), .ZN(n13367) );
  AOI21_X1 U15621 ( .B1(n13388), .B2(n13367), .A(n15752), .ZN(n13371) );
  AOI21_X1 U15622 ( .B1(n15732), .B2(P3_ADDR_REG_18__SCAN_IN), .A(n13368), 
        .ZN(n13369) );
  OAI21_X1 U15623 ( .B1(n15738), .B2(n13380), .A(n13369), .ZN(n13370) );
  AOI211_X1 U15624 ( .C1(n13372), .C2(n13395), .A(n13371), .B(n13370), .ZN(
        n13373) );
  OAI21_X1 U15625 ( .B1(n13374), .B2(n15744), .A(n13373), .ZN(P3_U3200) );
  INV_X1 U15626 ( .A(n13375), .ZN(n13376) );
  XNOR2_X1 U15627 ( .A(n13393), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13384) );
  INV_X1 U15628 ( .A(n13384), .ZN(n13378) );
  XNOR2_X1 U15629 ( .A(n13379), .B(n13378), .ZN(n13397) );
  INV_X1 U15630 ( .A(n13380), .ZN(n13382) );
  AOI21_X1 U15631 ( .B1(n13383), .B2(n13382), .A(n13381), .ZN(n13386) );
  XNOR2_X1 U15632 ( .A(n13393), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n13389) );
  MUX2_X1 U15633 ( .A(n13389), .B(n13384), .S(n10612), .Z(n13385) );
  XNOR2_X1 U15634 ( .A(n13386), .B(n13385), .ZN(n13396) );
  NAND2_X1 U15635 ( .A1(n13388), .A2(n13387), .ZN(n13390) );
  AOI21_X1 U15636 ( .B1(n15732), .B2(P3_ADDR_REG_19__SCAN_IN), .A(n13391), 
        .ZN(n13392) );
  OAI21_X1 U15637 ( .B1(n15738), .B2(n13393), .A(n13392), .ZN(n13394) );
  INV_X1 U15638 ( .A(n13398), .ZN(n13404) );
  AOI22_X1 U15639 ( .A1(n15162), .A2(n15818), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n15822), .ZN(n13399) );
  OAI21_X1 U15640 ( .B1(n13400), .B2(n15760), .A(n13399), .ZN(n13401) );
  AOI21_X1 U15641 ( .B1(n13402), .B2(n15218), .A(n13401), .ZN(n13403) );
  OAI21_X1 U15642 ( .B1(n13404), .B2(n15822), .A(n13403), .ZN(P3_U3204) );
  XNOR2_X1 U15643 ( .A(n13407), .B(n13406), .ZN(n13586) );
  INV_X1 U15644 ( .A(n13586), .ZN(n13421) );
  NAND2_X1 U15645 ( .A1(n13408), .A2(n15211), .ZN(n13409) );
  OAI22_X1 U15646 ( .A1(n13411), .A2(n15787), .B1(n13434), .B2(n15789), .ZN(
        n13412) );
  INV_X1 U15647 ( .A(n13412), .ZN(n13413) );
  NAND2_X1 U15648 ( .A1(n13414), .A2(n13413), .ZN(n13587) );
  INV_X1 U15649 ( .A(n13415), .ZN(n13643) );
  AOI22_X1 U15650 ( .A1(n13416), .A2(n15818), .B1(n15822), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n13417) );
  OAI21_X1 U15651 ( .B1(n13643), .B2(n15760), .A(n13417), .ZN(n13418) );
  AOI21_X1 U15652 ( .B1(n13587), .B2(n15801), .A(n13418), .ZN(n13419) );
  OAI21_X1 U15653 ( .B1(n13421), .B2(n13420), .A(n13419), .ZN(P3_U3205) );
  INV_X1 U15654 ( .A(n13422), .ZN(n13429) );
  AOI22_X1 U15655 ( .A1(n13423), .A2(n15818), .B1(n15822), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13424) );
  OAI21_X1 U15656 ( .B1(n13425), .B2(n15760), .A(n13424), .ZN(n13426) );
  AOI21_X1 U15657 ( .B1(n13427), .B2(n15819), .A(n13426), .ZN(n13428) );
  OAI21_X1 U15658 ( .B1(n13429), .B2(n15822), .A(n13428), .ZN(P3_U3206) );
  XOR2_X1 U15659 ( .A(n13430), .B(n13432), .Z(n13437) );
  XNOR2_X1 U15660 ( .A(n13432), .B(n13431), .ZN(n13590) );
  OAI22_X1 U15661 ( .A1(n13434), .A2(n15787), .B1(n13433), .B2(n15789), .ZN(
        n13435) );
  AOI21_X1 U15662 ( .B1(n13590), .B2(n15814), .A(n13435), .ZN(n13436) );
  OAI21_X1 U15663 ( .B1(n13437), .B2(n15811), .A(n13436), .ZN(n13589) );
  INV_X1 U15664 ( .A(n13589), .ZN(n13442) );
  AOI22_X1 U15665 ( .A1(n15822), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n13438), 
        .B2(n15818), .ZN(n13439) );
  OAI21_X1 U15666 ( .B1(n13647), .B2(n15760), .A(n13439), .ZN(n13440) );
  AOI21_X1 U15667 ( .B1(n13590), .B2(n15819), .A(n13440), .ZN(n13441) );
  OAI21_X1 U15668 ( .B1(n13442), .B2(n15822), .A(n13441), .ZN(P3_U3207) );
  XNOR2_X1 U15669 ( .A(n13445), .B(n13443), .ZN(n13452) );
  OAI211_X1 U15670 ( .C1(n13446), .C2(n13445), .A(n13444), .B(n15211), .ZN(
        n13451) );
  OAI22_X1 U15671 ( .A1(n13448), .A2(n15787), .B1(n13447), .B2(n15789), .ZN(
        n13449) );
  INV_X1 U15672 ( .A(n13449), .ZN(n13450) );
  OAI211_X1 U15673 ( .C1(n13486), .C2(n13452), .A(n13451), .B(n13450), .ZN(
        n13593) );
  INV_X1 U15674 ( .A(n13593), .ZN(n13457) );
  INV_X1 U15675 ( .A(n13452), .ZN(n13594) );
  AOI22_X1 U15676 ( .A1(n15822), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n13453), 
        .B2(n15818), .ZN(n13454) );
  OAI21_X1 U15677 ( .B1(n13651), .B2(n15760), .A(n13454), .ZN(n13455) );
  AOI21_X1 U15678 ( .B1(n13594), .B2(n15819), .A(n13455), .ZN(n13456) );
  OAI21_X1 U15679 ( .B1(n13457), .B2(n15822), .A(n13456), .ZN(P3_U3208) );
  INV_X1 U15680 ( .A(n13458), .ZN(n13462) );
  AOI21_X1 U15681 ( .B1(n13479), .B2(n13460), .A(n13459), .ZN(n13461) );
  NOR2_X1 U15682 ( .A1(n13462), .A2(n13461), .ZN(n13470) );
  OAI211_X1 U15683 ( .C1(n13465), .C2(n13464), .A(n13463), .B(n15211), .ZN(
        n13469) );
  AOI22_X1 U15684 ( .A1(n13467), .A2(n15809), .B1(n15806), .B2(n13466), .ZN(
        n13468) );
  OAI211_X1 U15685 ( .C1(n13486), .C2(n13470), .A(n13469), .B(n13468), .ZN(
        n13597) );
  INV_X1 U15686 ( .A(n13597), .ZN(n13475) );
  INV_X1 U15687 ( .A(n13470), .ZN(n13598) );
  AOI22_X1 U15688 ( .A1(n15822), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n15818), 
        .B2(n13471), .ZN(n13472) );
  OAI21_X1 U15689 ( .B1(n13655), .B2(n15760), .A(n13472), .ZN(n13473) );
  AOI21_X1 U15690 ( .B1(n13598), .B2(n15819), .A(n13473), .ZN(n13474) );
  OAI21_X1 U15691 ( .B1(n13475), .B2(n15822), .A(n13474), .ZN(P3_U3209) );
  OR2_X1 U15692 ( .A1(n13477), .A2(n13476), .ZN(n13478) );
  NAND2_X1 U15693 ( .A1(n13479), .A2(n13478), .ZN(n13487) );
  OAI211_X1 U15694 ( .C1(n6806), .C2(n13481), .A(n13480), .B(n15211), .ZN(
        n13485) );
  AOI22_X1 U15695 ( .A1(n13483), .A2(n15809), .B1(n13482), .B2(n15806), .ZN(
        n13484) );
  OAI211_X1 U15696 ( .C1(n13486), .C2(n13487), .A(n13485), .B(n13484), .ZN(
        n13601) );
  INV_X1 U15697 ( .A(n13601), .ZN(n13492) );
  INV_X1 U15698 ( .A(n13487), .ZN(n13602) );
  AOI22_X1 U15699 ( .A1(n15822), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n15818), 
        .B2(n13488), .ZN(n13489) );
  OAI21_X1 U15700 ( .B1(n13659), .B2(n15760), .A(n13489), .ZN(n13490) );
  AOI21_X1 U15701 ( .B1(n13602), .B2(n15819), .A(n13490), .ZN(n13491) );
  OAI21_X1 U15702 ( .B1(n13492), .B2(n15822), .A(n13491), .ZN(P3_U3210) );
  XNOR2_X1 U15703 ( .A(n13493), .B(n13497), .ZN(n13494) );
  OAI222_X1 U15704 ( .A1(n15789), .A2(n13496), .B1(n15787), .B2(n13495), .C1(
        n13494), .C2(n15811), .ZN(n13605) );
  INV_X1 U15705 ( .A(n13605), .ZN(n13504) );
  XNOR2_X1 U15706 ( .A(n13498), .B(n13497), .ZN(n13606) );
  INV_X1 U15707 ( .A(n13499), .ZN(n13663) );
  AOI22_X1 U15708 ( .A1(n15822), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15818), 
        .B2(n13500), .ZN(n13501) );
  OAI21_X1 U15709 ( .B1(n13663), .B2(n15760), .A(n13501), .ZN(n13502) );
  AOI21_X1 U15710 ( .B1(n13606), .B2(n15218), .A(n13502), .ZN(n13503) );
  OAI21_X1 U15711 ( .B1(n13504), .B2(n15822), .A(n13503), .ZN(P3_U3211) );
  XNOR2_X1 U15712 ( .A(n13505), .B(n13510), .ZN(n13506) );
  OAI222_X1 U15713 ( .A1(n15789), .A2(n13508), .B1(n15787), .B2(n13507), .C1(
        n15811), .C2(n13506), .ZN(n13609) );
  INV_X1 U15714 ( .A(n13609), .ZN(n13515) );
  XNOR2_X1 U15715 ( .A(n13509), .B(n13510), .ZN(n13610) );
  AOI22_X1 U15716 ( .A1(n15822), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15818), 
        .B2(n13511), .ZN(n13512) );
  OAI21_X1 U15717 ( .B1(n13667), .B2(n15760), .A(n13512), .ZN(n13513) );
  AOI21_X1 U15718 ( .B1(n13610), .B2(n15218), .A(n13513), .ZN(n13514) );
  OAI21_X1 U15719 ( .B1(n13515), .B2(n15822), .A(n13514), .ZN(P3_U3212) );
  OAI211_X1 U15720 ( .C1(n13525), .C2(n13517), .A(n13516), .B(n15211), .ZN(
        n13521) );
  AOI22_X1 U15721 ( .A1(n13519), .A2(n15809), .B1(n15806), .B2(n13518), .ZN(
        n13520) );
  INV_X1 U15722 ( .A(n13523), .ZN(n13524) );
  AOI21_X1 U15723 ( .B1(n13525), .B2(n13522), .A(n13524), .ZN(n13614) );
  AOI22_X1 U15724 ( .A1(n15822), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15818), 
        .B2(n13526), .ZN(n13527) );
  OAI21_X1 U15725 ( .B1(n13528), .B2(n15760), .A(n13527), .ZN(n13529) );
  AOI21_X1 U15726 ( .B1(n13614), .B2(n15218), .A(n13529), .ZN(n13530) );
  OAI21_X1 U15727 ( .B1(n13616), .B2(n15822), .A(n13530), .ZN(P3_U3213) );
  OAI211_X1 U15728 ( .C1(n6821), .C2(n13535), .A(n13531), .B(n15211), .ZN(
        n13534) );
  AOI22_X1 U15729 ( .A1(n13532), .A2(n15809), .B1(n15806), .B2(n13560), .ZN(
        n13533) );
  AND2_X1 U15730 ( .A1(n13534), .A2(n13533), .ZN(n13619) );
  XNOR2_X1 U15731 ( .A(n13536), .B(n13535), .ZN(n13617) );
  INV_X1 U15732 ( .A(n13671), .ZN(n13539) );
  AOI22_X1 U15733 ( .A1(n15822), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15818), 
        .B2(n13537), .ZN(n13538) );
  OAI21_X1 U15734 ( .B1(n13539), .B2(n15760), .A(n13538), .ZN(n13540) );
  AOI21_X1 U15735 ( .B1(n13617), .B2(n15218), .A(n13540), .ZN(n13541) );
  OAI21_X1 U15736 ( .B1(n13619), .B2(n15822), .A(n13541), .ZN(P3_U3214) );
  INV_X1 U15737 ( .A(n13542), .ZN(n13543) );
  AOI21_X1 U15738 ( .B1(n13548), .B2(n13544), .A(n13543), .ZN(n13545) );
  OAI222_X1 U15739 ( .A1(n15787), .A2(n13547), .B1(n15789), .B2(n13546), .C1(
        n15811), .C2(n13545), .ZN(n13622) );
  INV_X1 U15740 ( .A(n13622), .ZN(n13555) );
  XNOR2_X1 U15741 ( .A(n13549), .B(n13548), .ZN(n13623) );
  INV_X1 U15742 ( .A(n13550), .ZN(n13677) );
  AOI22_X1 U15743 ( .A1(n15822), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15818), 
        .B2(n13551), .ZN(n13552) );
  OAI21_X1 U15744 ( .B1(n13677), .B2(n15760), .A(n13552), .ZN(n13553) );
  AOI21_X1 U15745 ( .B1(n13623), .B2(n15218), .A(n13553), .ZN(n13554) );
  OAI21_X1 U15746 ( .B1(n13555), .B2(n15822), .A(n13554), .ZN(P3_U3215) );
  OAI211_X1 U15747 ( .C1(n13558), .C2(n13557), .A(n13556), .B(n15211), .ZN(
        n13562) );
  AOI22_X1 U15748 ( .A1(n15809), .A2(n13560), .B1(n13559), .B2(n15806), .ZN(
        n13561) );
  AND2_X1 U15749 ( .A1(n13562), .A2(n13561), .ZN(n13630) );
  OAI21_X1 U15750 ( .B1(n13565), .B2(n13564), .A(n13563), .ZN(n13628) );
  AOI22_X1 U15751 ( .A1(n15822), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15818), 
        .B2(n13566), .ZN(n13567) );
  OAI21_X1 U15752 ( .B1(n13568), .B2(n15760), .A(n13567), .ZN(n13569) );
  AOI21_X1 U15753 ( .B1(n13628), .B2(n15218), .A(n13569), .ZN(n13570) );
  OAI21_X1 U15754 ( .B1(n13630), .B2(n15822), .A(n13570), .ZN(P3_U3216) );
  NAND2_X1 U15755 ( .A1(n13571), .A2(n13577), .ZN(n13572) );
  NAND3_X1 U15756 ( .A1(n13573), .A2(n15211), .A3(n13572), .ZN(n13576) );
  AOI22_X1 U15757 ( .A1(n15809), .A2(n13574), .B1(n15173), .B2(n15806), .ZN(
        n13575) );
  AND2_X1 U15758 ( .A1(n13576), .A2(n13575), .ZN(n13633) );
  OR2_X1 U15759 ( .A1(n13578), .A2(n13577), .ZN(n13579) );
  NAND2_X1 U15760 ( .A1(n13580), .A2(n13579), .ZN(n13631) );
  INV_X1 U15761 ( .A(n13681), .ZN(n13583) );
  AOI22_X1 U15762 ( .A1(n15822), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15818), 
        .B2(n13581), .ZN(n13582) );
  OAI21_X1 U15763 ( .B1(n13583), .B2(n15760), .A(n13582), .ZN(n13584) );
  AOI21_X1 U15764 ( .B1(n13631), .B2(n15218), .A(n13584), .ZN(n13585) );
  OAI21_X1 U15765 ( .B1(n13633), .B2(n15822), .A(n13585), .ZN(P3_U3217) );
  AOI21_X1 U15766 ( .B1(n15842), .B2(n13590), .A(n13589), .ZN(n13644) );
  MUX2_X1 U15767 ( .A(n13591), .B(n13644), .S(n15854), .Z(n13592) );
  OAI21_X1 U15768 ( .B1(n13647), .B2(n13626), .A(n13592), .ZN(P3_U3485) );
  AOI21_X1 U15769 ( .B1(n15842), .B2(n13594), .A(n13593), .ZN(n13648) );
  MUX2_X1 U15770 ( .A(n13595), .B(n13648), .S(n15854), .Z(n13596) );
  OAI21_X1 U15771 ( .B1(n13651), .B2(n13626), .A(n13596), .ZN(P3_U3484) );
  AOI21_X1 U15772 ( .B1(n15842), .B2(n13598), .A(n13597), .ZN(n13652) );
  MUX2_X1 U15773 ( .A(n13599), .B(n13652), .S(n15854), .Z(n13600) );
  OAI21_X1 U15774 ( .B1(n13655), .B2(n13626), .A(n13600), .ZN(P3_U3483) );
  AOI21_X1 U15775 ( .B1(n15842), .B2(n13602), .A(n13601), .ZN(n13656) );
  MUX2_X1 U15776 ( .A(n13603), .B(n13656), .S(n15854), .Z(n13604) );
  OAI21_X1 U15777 ( .B1(n13659), .B2(n13626), .A(n13604), .ZN(P3_U3482) );
  AOI21_X1 U15778 ( .B1(n15241), .B2(n13606), .A(n13605), .ZN(n13660) );
  MUX2_X1 U15779 ( .A(n13607), .B(n13660), .S(n15854), .Z(n13608) );
  OAI21_X1 U15780 ( .B1(n13663), .B2(n13626), .A(n13608), .ZN(P3_U3481) );
  INV_X1 U15781 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13611) );
  AOI21_X1 U15782 ( .B1(n13610), .B2(n15241), .A(n13609), .ZN(n13664) );
  MUX2_X1 U15783 ( .A(n13611), .B(n13664), .S(n15854), .Z(n13612) );
  OAI21_X1 U15784 ( .B1(n13667), .B2(n13626), .A(n13612), .ZN(P3_U3480) );
  AOI22_X1 U15785 ( .A1(n13614), .A2(n15241), .B1(n15796), .B2(n13613), .ZN(
        n13615) );
  NAND2_X1 U15786 ( .A1(n13616), .A2(n13615), .ZN(n13668) );
  MUX2_X1 U15787 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n13668), .S(n15854), .Z(
        P3_U3479) );
  NAND2_X1 U15788 ( .A1(n13617), .A2(n15241), .ZN(n13618) );
  NAND2_X1 U15789 ( .A1(n13619), .A2(n13618), .ZN(n13669) );
  MUX2_X1 U15790 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n13669), .S(n15854), .Z(
        n13620) );
  AOI21_X1 U15791 ( .B1(n13635), .B2(n13671), .A(n13620), .ZN(n13621) );
  INV_X1 U15792 ( .A(n13621), .ZN(P3_U3478) );
  AOI21_X1 U15793 ( .B1(n13623), .B2(n15241), .A(n13622), .ZN(n13673) );
  MUX2_X1 U15794 ( .A(n13624), .B(n13673), .S(n15854), .Z(n13625) );
  OAI21_X1 U15795 ( .B1(n13677), .B2(n13626), .A(n13625), .ZN(P3_U3477) );
  AOI22_X1 U15796 ( .A1(n13628), .A2(n15241), .B1(n13627), .B2(n15796), .ZN(
        n13629) );
  NAND2_X1 U15797 ( .A1(n13630), .A2(n13629), .ZN(n13678) );
  MUX2_X1 U15798 ( .A(n13678), .B(P3_REG1_REG_17__SCAN_IN), .S(n15851), .Z(
        P3_U3476) );
  NAND2_X1 U15799 ( .A1(n13631), .A2(n15241), .ZN(n13632) );
  NAND2_X1 U15800 ( .A1(n13633), .A2(n13632), .ZN(n13679) );
  MUX2_X1 U15801 ( .A(n13679), .B(P3_REG1_REG_16__SCAN_IN), .S(n15851), .Z(
        n13634) );
  AOI21_X1 U15802 ( .B1(n13635), .B2(n13681), .A(n13634), .ZN(n13636) );
  INV_X1 U15803 ( .A(n13636), .ZN(P3_U3475) );
  AOI22_X1 U15804 ( .A1(n13638), .A2(n15241), .B1(n13637), .B2(n15796), .ZN(
        n13639) );
  NAND2_X1 U15805 ( .A1(n13640), .A2(n13639), .ZN(n13684) );
  MUX2_X1 U15806 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n13684), .S(n15854), .Z(
        P3_U3474) );
  INV_X1 U15807 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13642) );
  INV_X1 U15808 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13645) );
  MUX2_X1 U15809 ( .A(n13645), .B(n13644), .S(n15846), .Z(n13646) );
  OAI21_X1 U15810 ( .B1(n13647), .B2(n13676), .A(n13646), .ZN(P3_U3453) );
  INV_X1 U15811 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13649) );
  MUX2_X1 U15812 ( .A(n13649), .B(n13648), .S(n15846), .Z(n13650) );
  OAI21_X1 U15813 ( .B1(n13651), .B2(n13676), .A(n13650), .ZN(P3_U3452) );
  INV_X1 U15814 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13653) );
  MUX2_X1 U15815 ( .A(n13653), .B(n13652), .S(n15846), .Z(n13654) );
  OAI21_X1 U15816 ( .B1(n13655), .B2(n13676), .A(n13654), .ZN(P3_U3451) );
  INV_X1 U15817 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13657) );
  MUX2_X1 U15818 ( .A(n13657), .B(n13656), .S(n15846), .Z(n13658) );
  OAI21_X1 U15819 ( .B1(n13659), .B2(n13676), .A(n13658), .ZN(P3_U3450) );
  INV_X1 U15820 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13661) );
  MUX2_X1 U15821 ( .A(n13661), .B(n13660), .S(n15846), .Z(n13662) );
  OAI21_X1 U15822 ( .B1(n13663), .B2(n13676), .A(n13662), .ZN(P3_U3449) );
  INV_X1 U15823 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13665) );
  MUX2_X1 U15824 ( .A(n13665), .B(n13664), .S(n15846), .Z(n13666) );
  OAI21_X1 U15825 ( .B1(n13667), .B2(n13676), .A(n13666), .ZN(P3_U3448) );
  MUX2_X1 U15826 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n13668), .S(n15846), .Z(
        P3_U3447) );
  INV_X1 U15827 ( .A(n13676), .ZN(n13682) );
  MUX2_X1 U15828 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n13669), .S(n15846), .Z(
        n13670) );
  AOI21_X1 U15829 ( .B1(n13682), .B2(n13671), .A(n13670), .ZN(n13672) );
  INV_X1 U15830 ( .A(n13672), .ZN(P3_U3446) );
  INV_X1 U15831 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13674) );
  MUX2_X1 U15832 ( .A(n13674), .B(n13673), .S(n15846), .Z(n13675) );
  OAI21_X1 U15833 ( .B1(n13677), .B2(n13676), .A(n13675), .ZN(P3_U3444) );
  MUX2_X1 U15834 ( .A(n13678), .B(P3_REG0_REG_17__SCAN_IN), .S(n15844), .Z(
        P3_U3441) );
  MUX2_X1 U15835 ( .A(n13679), .B(P3_REG0_REG_16__SCAN_IN), .S(n15844), .Z(
        n13680) );
  AOI21_X1 U15836 ( .B1(n13682), .B2(n13681), .A(n13680), .ZN(n13683) );
  INV_X1 U15837 ( .A(n13683), .ZN(P3_U3438) );
  MUX2_X1 U15838 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n13684), .S(n15846), .Z(
        P3_U3435) );
  MUX2_X1 U15839 ( .A(P3_D_REG_0__SCAN_IN), .B(n13686), .S(n13685), .Z(
        P3_U3376) );
  NAND2_X1 U15840 ( .A1(n13687), .A2(n15121), .ZN(n13691) );
  NAND2_X1 U15841 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_STATE_REG_SCAN_IN), 
        .ZN(n13688) );
  OR3_X1 U15842 ( .A1(n13689), .A2(P3_IR_REG_30__SCAN_IN), .A3(n13688), .ZN(
        n13690) );
  OAI211_X1 U15843 ( .C1(n13692), .C2(n13709), .A(n13691), .B(n13690), .ZN(
        P3_U3264) );
  OAI222_X1 U15844 ( .A1(P3_U3151), .A2(n13695), .B1(n13712), .B2(n13694), 
        .C1(n13693), .C2(n13709), .ZN(P3_U3265) );
  INV_X1 U15845 ( .A(n13696), .ZN(n13698) );
  OAI222_X1 U15846 ( .A1(n13715), .A2(n13699), .B1(n13712), .B2(n13698), .C1(
        n13697), .C2(P3_U3151), .ZN(P3_U3266) );
  INV_X1 U15847 ( .A(n13700), .ZN(n13703) );
  OAI222_X1 U15848 ( .A1(n13712), .A2(n13703), .B1(P3_U3151), .B2(n8266), .C1(
        n13701), .C2(n13709), .ZN(P3_U3267) );
  INV_X1 U15849 ( .A(n13704), .ZN(n13706) );
  OAI222_X1 U15850 ( .A1(P3_U3151), .A2(n10612), .B1(n13712), .B2(n13706), 
        .C1(n13705), .C2(n13709), .ZN(P3_U3268) );
  INV_X1 U15851 ( .A(n13707), .ZN(n13713) );
  INV_X1 U15852 ( .A(n13708), .ZN(n13711) );
  OAI222_X1 U15853 ( .A1(n13713), .A2(P3_U3151), .B1(n13712), .B2(n13711), 
        .C1(n13710), .C2(n13709), .ZN(P3_U3269) );
  INV_X1 U15854 ( .A(n13714), .ZN(n13717) );
  OAI222_X1 U15855 ( .A1(P3_U3151), .A2(n13718), .B1(n13712), .B2(n13717), 
        .C1(n13716), .C2(n13715), .ZN(P3_U3270) );
  XNOR2_X1 U15856 ( .A(n14394), .B(n7043), .ZN(n13749) );
  NAND2_X1 U15857 ( .A1(n13926), .A2(n13804), .ZN(n13879) );
  INV_X1 U15858 ( .A(n13719), .ZN(n13721) );
  NAND2_X1 U15859 ( .A1(n13721), .A2(n13720), .ZN(n13722) );
  XNOR2_X1 U15860 ( .A(n14364), .B(n7043), .ZN(n13846) );
  NAND2_X1 U15861 ( .A1(n13932), .A2(n13804), .ZN(n13725) );
  XNOR2_X1 U15862 ( .A(n13846), .B(n13725), .ZN(n13833) );
  NAND2_X1 U15863 ( .A1(n13846), .A2(n13725), .ZN(n13726) );
  XNOR2_X1 U15864 ( .A(n14359), .B(n13806), .ZN(n13728) );
  NAND2_X1 U15865 ( .A1(n13931), .A2(n13804), .ZN(n13729) );
  XNOR2_X1 U15866 ( .A(n13728), .B(n13729), .ZN(n13843) );
  NAND2_X1 U15867 ( .A1(n13727), .A2(n13843), .ZN(n13851) );
  INV_X1 U15868 ( .A(n13728), .ZN(n13730) );
  NAND2_X1 U15869 ( .A1(n13730), .A2(n13729), .ZN(n13731) );
  XNOR2_X1 U15870 ( .A(n14353), .B(n13806), .ZN(n13787) );
  AND2_X1 U15871 ( .A1(n13930), .A2(n13804), .ZN(n13732) );
  NAND2_X1 U15872 ( .A1(n13787), .A2(n13732), .ZN(n13737) );
  INV_X1 U15873 ( .A(n13787), .ZN(n13734) );
  INV_X1 U15874 ( .A(n13732), .ZN(n13733) );
  NAND2_X1 U15875 ( .A1(n13734), .A2(n13733), .ZN(n13735) );
  NAND2_X1 U15876 ( .A1(n13737), .A2(n13735), .ZN(n13891) );
  XNOR2_X1 U15877 ( .A(n14345), .B(n13806), .ZN(n13738) );
  NAND2_X1 U15878 ( .A1(n13929), .A2(n13804), .ZN(n13739) );
  XNOR2_X1 U15879 ( .A(n13738), .B(n13739), .ZN(n13789) );
  INV_X1 U15880 ( .A(n13738), .ZN(n13740) );
  NAND2_X1 U15881 ( .A1(n13740), .A2(n13739), .ZN(n13741) );
  XNOR2_X1 U15882 ( .A(n14341), .B(n7043), .ZN(n13742) );
  NAND2_X1 U15883 ( .A1(n13928), .A2(n13804), .ZN(n13743) );
  NAND2_X1 U15884 ( .A1(n13742), .A2(n13743), .ZN(n13864) );
  INV_X1 U15885 ( .A(n13742), .ZN(n13745) );
  INV_X1 U15886 ( .A(n13743), .ZN(n13744) );
  NAND2_X1 U15887 ( .A1(n13745), .A2(n13744), .ZN(n13863) );
  XNOR2_X1 U15888 ( .A(n14337), .B(n13806), .ZN(n13748) );
  NAND2_X1 U15889 ( .A1(n13927), .A2(n13804), .ZN(n13746) );
  XNOR2_X1 U15890 ( .A(n13748), .B(n13746), .ZN(n13816) );
  NAND2_X1 U15891 ( .A1(n13815), .A2(n13816), .ZN(n13874) );
  INV_X1 U15892 ( .A(n13746), .ZN(n13747) );
  NAND2_X1 U15893 ( .A1(n13748), .A2(n13747), .ZN(n13873) );
  OAI211_X1 U15894 ( .C1(n13749), .C2(n13879), .A(n13874), .B(n13873), .ZN(
        n13751) );
  INV_X1 U15895 ( .A(n13749), .ZN(n13875) );
  INV_X1 U15896 ( .A(n13879), .ZN(n13750) );
  NAND2_X1 U15897 ( .A1(n13925), .A2(n13804), .ZN(n13769) );
  XNOR2_X1 U15898 ( .A(n14316), .B(n7043), .ZN(n13754) );
  NAND2_X1 U15899 ( .A1(n13924), .A2(n13804), .ZN(n13753) );
  NAND2_X1 U15900 ( .A1(n13754), .A2(n13753), .ZN(n13755) );
  OAI21_X1 U15901 ( .B1(n13754), .B2(n13753), .A(n13755), .ZN(n13854) );
  INV_X1 U15902 ( .A(n13755), .ZN(n13756) );
  XNOR2_X1 U15903 ( .A(n14310), .B(n13806), .ZN(n13759) );
  NAND2_X1 U15904 ( .A1(n13923), .A2(n13804), .ZN(n13757) );
  XNOR2_X1 U15905 ( .A(n13759), .B(n13757), .ZN(n13822) );
  INV_X1 U15906 ( .A(n13757), .ZN(n13758) );
  AND2_X1 U15907 ( .A1(n13922), .A2(n13804), .ZN(n13761) );
  XNOR2_X1 U15908 ( .A(n14108), .B(n13806), .ZN(n13760) );
  NOR2_X1 U15909 ( .A1(n13760), .A2(n13761), .ZN(n13762) );
  AOI21_X1 U15910 ( .B1(n13761), .B2(n13760), .A(n13762), .ZN(n13903) );
  NAND2_X1 U15911 ( .A1(n13921), .A2(n13804), .ZN(n13800) );
  XNOR2_X1 U15912 ( .A(n14091), .B(n13806), .ZN(n13799) );
  XOR2_X1 U15913 ( .A(n13800), .B(n13799), .Z(n13802) );
  XNOR2_X1 U15914 ( .A(n13803), .B(n13802), .ZN(n13768) );
  OAI22_X1 U15915 ( .A1(n13764), .A2(n13857), .B1(n13763), .B2(n13855), .ZN(
        n14086) );
  AOI22_X1 U15916 ( .A1(n13910), .A2(n14086), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13765) );
  OAI21_X1 U15917 ( .B1(n14092), .B2(n13912), .A(n13765), .ZN(n13766) );
  AOI21_X1 U15918 ( .B1(n14091), .B2(n13914), .A(n13766), .ZN(n13767) );
  OAI21_X1 U15919 ( .B1(n13768), .B2(n13916), .A(n13767), .ZN(P2_U3186) );
  NAND2_X1 U15920 ( .A1(n13769), .A2(n13880), .ZN(n13772) );
  NAND2_X1 U15921 ( .A1(n13877), .A2(n13925), .ZN(n13771) );
  MUX2_X1 U15922 ( .A(n13772), .B(n13771), .S(n13770), .Z(n13777) );
  AND2_X1 U15923 ( .A1(n13924), .A2(n13907), .ZN(n13773) );
  AOI21_X1 U15924 ( .B1(n13926), .B2(n13906), .A(n13773), .ZN(n14152) );
  OAI22_X1 U15925 ( .A1(n13884), .A2(n14152), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13774), .ZN(n13775) );
  AOI21_X1 U15926 ( .B1(n14155), .B2(n13886), .A(n13775), .ZN(n13776) );
  OAI211_X1 U15927 ( .C1(n14391), .C2(n13901), .A(n13777), .B(n13776), .ZN(
        P2_U3188) );
  AOI21_X1 U15928 ( .B1(n13779), .B2(n13778), .A(n13916), .ZN(n13781) );
  NAND2_X1 U15929 ( .A1(n13781), .A2(n13780), .ZN(n13786) );
  AOI22_X1 U15930 ( .A1(n13783), .A2(n13914), .B1(n13910), .B2(n13782), .ZN(
        n13785) );
  MUX2_X1 U15931 ( .A(n13912), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n13784) );
  NAND3_X1 U15932 ( .A1(n13786), .A2(n13785), .A3(n13784), .ZN(P2_U3190) );
  NAND3_X1 U15933 ( .A1(n13787), .A2(n13877), .A3(n13930), .ZN(n13788) );
  OAI21_X1 U15934 ( .B1(n13893), .B2(n13916), .A(n13788), .ZN(n13791) );
  INV_X1 U15935 ( .A(n13789), .ZN(n13790) );
  NAND2_X1 U15936 ( .A1(n13791), .A2(n13790), .ZN(n13797) );
  NOR2_X1 U15937 ( .A1(n13912), .A2(n14219), .ZN(n13795) );
  AND2_X1 U15938 ( .A1(n13930), .A2(n13906), .ZN(n13792) );
  AOI21_X1 U15939 ( .B1(n13928), .B2(n13907), .A(n13792), .ZN(n14216) );
  OAI21_X1 U15940 ( .B1(n13884), .B2(n14216), .A(n13793), .ZN(n13794) );
  AOI211_X1 U15941 ( .C1(n14345), .C2(n13914), .A(n13795), .B(n13794), .ZN(
        n13796) );
  OAI211_X1 U15942 ( .C1(n13798), .C2(n13916), .A(n13797), .B(n13796), .ZN(
        P2_U3191) );
  INV_X1 U15943 ( .A(n13799), .ZN(n13801) );
  NAND2_X1 U15944 ( .A1(n13920), .A2(n13804), .ZN(n13805) );
  XNOR2_X1 U15945 ( .A(n13806), .B(n13805), .ZN(n13807) );
  XNOR2_X1 U15946 ( .A(n14292), .B(n13807), .ZN(n13808) );
  OAI22_X1 U15947 ( .A1(n13810), .A2(n13857), .B1(n13809), .B2(n13855), .ZN(
        n14075) );
  AOI22_X1 U15948 ( .A1(n13910), .A2(n14075), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13811) );
  OAI21_X1 U15949 ( .B1(n14080), .B2(n13912), .A(n13811), .ZN(n13812) );
  AOI21_X1 U15950 ( .B1(n14292), .B2(n13914), .A(n13812), .ZN(n13813) );
  OAI21_X1 U15951 ( .B1(n13814), .B2(n13916), .A(n13813), .ZN(P2_U3192) );
  XNOR2_X1 U15952 ( .A(n13815), .B(n13816), .ZN(n13821) );
  AOI22_X1 U15953 ( .A1(n13926), .A2(n13907), .B1(n13906), .B2(n13928), .ZN(
        n14183) );
  INV_X1 U15954 ( .A(n14183), .ZN(n13817) );
  AOI22_X1 U15955 ( .A1(n13817), .A2(n13910), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13818) );
  OAI21_X1 U15956 ( .B1(n14187), .B2(n13912), .A(n13818), .ZN(n13819) );
  AOI21_X1 U15957 ( .B1(n14337), .B2(n13914), .A(n13819), .ZN(n13820) );
  OAI21_X1 U15958 ( .B1(n13821), .B2(n13916), .A(n13820), .ZN(P2_U3195) );
  XNOR2_X1 U15959 ( .A(n13823), .B(n13822), .ZN(n13829) );
  NAND2_X1 U15960 ( .A1(n13922), .A2(n13907), .ZN(n13825) );
  NAND2_X1 U15961 ( .A1(n13924), .A2(n13906), .ZN(n13824) );
  NAND2_X1 U15962 ( .A1(n13825), .A2(n13824), .ZN(n14114) );
  AOI22_X1 U15963 ( .A1(n13910), .A2(n14114), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13826) );
  OAI21_X1 U15964 ( .B1(n14121), .B2(n13912), .A(n13826), .ZN(n13827) );
  AOI21_X1 U15965 ( .B1(n14310), .B2(n13914), .A(n13827), .ZN(n13828) );
  OAI21_X1 U15966 ( .B1(n13829), .B2(n13916), .A(n13828), .ZN(P2_U3197) );
  INV_X1 U15967 ( .A(n13830), .ZN(n13831) );
  AOI21_X1 U15968 ( .B1(n13833), .B2(n13832), .A(n13831), .ZN(n13839) );
  NAND2_X1 U15969 ( .A1(n13931), .A2(n13907), .ZN(n13835) );
  NAND2_X1 U15970 ( .A1(n13933), .A2(n13906), .ZN(n13834) );
  NAND2_X1 U15971 ( .A1(n13835), .A2(n13834), .ZN(n14266) );
  AOI22_X1 U15972 ( .A1(n13910), .A2(n14266), .B1(P2_REG3_REG_16__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13836) );
  OAI21_X1 U15973 ( .B1(n14271), .B2(n13912), .A(n13836), .ZN(n13837) );
  AOI21_X1 U15974 ( .B1(n14364), .B2(n13914), .A(n13837), .ZN(n13838) );
  OAI21_X1 U15975 ( .B1(n13839), .B2(n13916), .A(n13838), .ZN(P2_U3198) );
  OAI22_X1 U15976 ( .A1(n13840), .A2(n13855), .B1(n13845), .B2(n13857), .ZN(
        n14246) );
  AOI22_X1 U15977 ( .A1(n13910), .A2(n14246), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13841) );
  OAI21_X1 U15978 ( .B1(n14253), .B2(n13912), .A(n13841), .ZN(n13842) );
  AOI21_X1 U15979 ( .B1(n14359), .B2(n13914), .A(n13842), .ZN(n13850) );
  INV_X1 U15980 ( .A(n13843), .ZN(n13848) );
  OAI22_X1 U15981 ( .A1(n13846), .A2(n13916), .B1(n13845), .B2(n13844), .ZN(
        n13847) );
  NAND3_X1 U15982 ( .A1(n13830), .A2(n13848), .A3(n13847), .ZN(n13849) );
  OAI211_X1 U15983 ( .C1(n13851), .C2(n13916), .A(n13850), .B(n13849), .ZN(
        P2_U3200) );
  AOI21_X1 U15984 ( .B1(n13854), .B2(n13853), .A(n13852), .ZN(n13862) );
  OAI22_X1 U15985 ( .A1(n13858), .A2(n13857), .B1(n13856), .B2(n13855), .ZN(
        n14131) );
  AOI22_X1 U15986 ( .A1(n14131), .A2(n13910), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13859) );
  OAI21_X1 U15987 ( .B1(n14136), .B2(n13912), .A(n13859), .ZN(n13860) );
  AOI21_X1 U15988 ( .B1(n14316), .B2(n13914), .A(n13860), .ZN(n13861) );
  OAI21_X1 U15989 ( .B1(n13862), .B2(n13916), .A(n13861), .ZN(P2_U3201) );
  NAND2_X1 U15990 ( .A1(n13864), .A2(n13863), .ZN(n13866) );
  XOR2_X1 U15991 ( .A(n13866), .B(n13865), .Z(n13872) );
  AND2_X1 U15992 ( .A1(n13929), .A2(n13906), .ZN(n13867) );
  AOI21_X1 U15993 ( .B1(n13927), .B2(n13907), .A(n13867), .ZN(n14199) );
  OAI22_X1 U15994 ( .A1(n13884), .A2(n14199), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13868), .ZN(n13869) );
  AOI21_X1 U15995 ( .B1(n14205), .B2(n13886), .A(n13869), .ZN(n13871) );
  NAND2_X1 U15996 ( .A1(n14341), .A2(n13914), .ZN(n13870) );
  OAI211_X1 U15997 ( .C1(n13872), .C2(n13916), .A(n13871), .B(n13870), .ZN(
        P2_U3205) );
  NAND2_X1 U15998 ( .A1(n13874), .A2(n13873), .ZN(n13876) );
  XNOR2_X1 U15999 ( .A(n13876), .B(n13875), .ZN(n13878) );
  NAND3_X1 U16000 ( .A1(n13878), .A2(n13877), .A3(n13926), .ZN(n13890) );
  INV_X1 U16001 ( .A(n13878), .ZN(n13881) );
  NAND3_X1 U16002 ( .A1(n13881), .A2(n13880), .A3(n13879), .ZN(n13889) );
  AND2_X1 U16003 ( .A1(n13927), .A2(n13906), .ZN(n13882) );
  AOI21_X1 U16004 ( .B1(n13925), .B2(n13907), .A(n13882), .ZN(n14170) );
  OAI22_X1 U16005 ( .A1(n14170), .A2(n13884), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13883), .ZN(n13885) );
  AOI21_X1 U16006 ( .B1(n14173), .B2(n13886), .A(n13885), .ZN(n13888) );
  NAND2_X1 U16007 ( .A1(n14394), .A2(n13914), .ZN(n13887) );
  NAND4_X1 U16008 ( .A1(n13890), .A2(n13889), .A3(n13888), .A4(n13887), .ZN(
        P2_U3207) );
  INV_X1 U16009 ( .A(n14353), .ZN(n14236) );
  AOI21_X1 U16010 ( .B1(n13892), .B2(n13891), .A(n13916), .ZN(n13894) );
  NAND2_X1 U16011 ( .A1(n13894), .A2(n13893), .ZN(n13900) );
  NAND2_X1 U16012 ( .A1(n13929), .A2(n13907), .ZN(n13896) );
  NAND2_X1 U16013 ( .A1(n13931), .A2(n13906), .ZN(n13895) );
  NAND2_X1 U16014 ( .A1(n13896), .A2(n13895), .ZN(n14230) );
  NOR2_X1 U16015 ( .A1(n13912), .A2(n14233), .ZN(n13897) );
  AOI211_X1 U16016 ( .C1(n13910), .C2(n14230), .A(n13898), .B(n13897), .ZN(
        n13899) );
  OAI211_X1 U16017 ( .C1(n14236), .C2(n13901), .A(n13900), .B(n13899), .ZN(
        P2_U3210) );
  OAI21_X1 U16018 ( .B1(n13904), .B2(n13903), .A(n13902), .ZN(n13905) );
  INV_X1 U16019 ( .A(n13905), .ZN(n13917) );
  NAND2_X1 U16020 ( .A1(n13923), .A2(n13906), .ZN(n13909) );
  NAND2_X1 U16021 ( .A1(n13921), .A2(n13907), .ZN(n13908) );
  NAND2_X1 U16022 ( .A1(n13909), .A2(n13908), .ZN(n14100) );
  AOI22_X1 U16023 ( .A1(n13910), .A2(n14100), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13911) );
  OAI21_X1 U16024 ( .B1(n14106), .B2(n13912), .A(n13911), .ZN(n13913) );
  AOI21_X1 U16025 ( .B1(n14108), .B2(n13914), .A(n13913), .ZN(n13915) );
  OAI21_X1 U16026 ( .B1(n13917), .B2(n13916), .A(n13915), .ZN(P2_U3212) );
  MUX2_X1 U16027 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n14052), .S(n15560), .Z(
        P2_U3562) );
  MUX2_X1 U16028 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13918), .S(n15560), .Z(
        P2_U3561) );
  MUX2_X1 U16029 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13919), .S(n15560), .Z(
        P2_U3560) );
  MUX2_X1 U16030 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13920), .S(n15560), .Z(
        P2_U3559) );
  MUX2_X1 U16031 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13921), .S(n15560), .Z(
        P2_U3558) );
  MUX2_X1 U16032 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13922), .S(n15560), .Z(
        P2_U3557) );
  MUX2_X1 U16033 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13923), .S(n15560), .Z(
        P2_U3556) );
  MUX2_X1 U16034 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13924), .S(n15560), .Z(
        P2_U3555) );
  MUX2_X1 U16035 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13925), .S(n15560), .Z(
        P2_U3554) );
  MUX2_X1 U16036 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13926), .S(n15560), .Z(
        P2_U3553) );
  MUX2_X1 U16037 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13927), .S(n15560), .Z(
        P2_U3552) );
  MUX2_X1 U16038 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13928), .S(n15560), .Z(
        P2_U3551) );
  MUX2_X1 U16039 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13929), .S(n15560), .Z(
        P2_U3550) );
  MUX2_X1 U16040 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13930), .S(n15560), .Z(
        P2_U3549) );
  MUX2_X1 U16041 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13931), .S(n15560), .Z(
        P2_U3548) );
  MUX2_X1 U16042 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13932), .S(n15560), .Z(
        P2_U3547) );
  MUX2_X1 U16043 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13933), .S(n15560), .Z(
        P2_U3546) );
  MUX2_X1 U16044 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13934), .S(n15560), .Z(
        P2_U3545) );
  MUX2_X1 U16045 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13935), .S(n15560), .Z(
        P2_U3544) );
  MUX2_X1 U16046 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13936), .S(n15560), .Z(
        P2_U3543) );
  MUX2_X1 U16047 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13937), .S(n15560), .Z(
        P2_U3542) );
  MUX2_X1 U16048 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13938), .S(n15560), .Z(
        P2_U3541) );
  MUX2_X1 U16049 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13939), .S(P2_U3947), .Z(
        P2_U3540) );
  MUX2_X1 U16050 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13940), .S(P2_U3947), .Z(
        P2_U3539) );
  MUX2_X1 U16051 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13941), .S(P2_U3947), .Z(
        P2_U3538) );
  MUX2_X1 U16052 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13942), .S(n15560), .Z(
        P2_U3537) );
  MUX2_X1 U16053 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13943), .S(P2_U3947), .Z(
        P2_U3536) );
  MUX2_X1 U16054 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13944), .S(P2_U3947), .Z(
        P2_U3535) );
  MUX2_X1 U16055 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13945), .S(P2_U3947), .Z(
        P2_U3534) );
  MUX2_X1 U16056 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13946), .S(P2_U3947), .Z(
        P2_U3533) );
  MUX2_X1 U16057 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n9686), .S(P2_U3947), .Z(
        P2_U3532) );
  MUX2_X1 U16058 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n13947), .S(P2_U3947), .Z(
        P2_U3531) );
  OAI211_X1 U16059 ( .C1(n13949), .C2(n13948), .A(n15639), .B(n13961), .ZN(
        n13958) );
  AOI22_X1 U16060 ( .A1(n15635), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(P2_U3088), .ZN(n13957) );
  NAND2_X1 U16061 ( .A1(n15641), .A2(n13950), .ZN(n13956) );
  MUX2_X1 U16062 ( .A(n11572), .B(P2_REG2_REG_3__SCAN_IN), .S(n13950), .Z(
        n13952) );
  NAND3_X1 U16063 ( .A1(n13953), .A2(n13952), .A3(n13951), .ZN(n13954) );
  NAND3_X1 U16064 ( .A1(n15644), .A2(n13968), .A3(n13954), .ZN(n13955) );
  NAND4_X1 U16065 ( .A1(n13958), .A2(n13957), .A3(n13956), .A4(n13955), .ZN(
        P2_U3217) );
  MUX2_X1 U16066 ( .A(n10816), .B(P2_REG1_REG_4__SCAN_IN), .S(n13964), .Z(
        n13959) );
  NAND3_X1 U16067 ( .A1(n13961), .A2(n13960), .A3(n13959), .ZN(n13962) );
  NAND3_X1 U16068 ( .A1(n15639), .A2(n13984), .A3(n13962), .ZN(n13973) );
  NAND2_X1 U16069 ( .A1(n15641), .A2(n13964), .ZN(n13972) );
  AOI21_X1 U16070 ( .B1(n15635), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n13963), .ZN(
        n13971) );
  MUX2_X1 U16071 ( .A(n13965), .B(P2_REG2_REG_4__SCAN_IN), .S(n13964), .Z(
        n13966) );
  NAND3_X1 U16072 ( .A1(n13968), .A2(n13967), .A3(n13966), .ZN(n13969) );
  NAND3_X1 U16073 ( .A1(n15644), .A2(n13978), .A3(n13969), .ZN(n13970) );
  NAND4_X1 U16074 ( .A1(n13973), .A2(n13972), .A3(n13971), .A4(n13970), .ZN(
        P2_U3218) );
  OAI21_X1 U16075 ( .B1(n15592), .B2(n15859), .A(n13974), .ZN(n13975) );
  AOI21_X1 U16076 ( .B1(n13980), .B2(n15641), .A(n13975), .ZN(n13988) );
  MUX2_X1 U16077 ( .A(n11589), .B(P2_REG2_REG_5__SCAN_IN), .S(n13980), .Z(
        n13976) );
  NAND3_X1 U16078 ( .A1(n13978), .A2(n13977), .A3(n13976), .ZN(n13979) );
  NAND3_X1 U16079 ( .A1(n15644), .A2(n13993), .A3(n13979), .ZN(n13987) );
  MUX2_X1 U16080 ( .A(n13981), .B(P2_REG1_REG_5__SCAN_IN), .S(n13980), .Z(
        n13982) );
  NAND3_X1 U16081 ( .A1(n13984), .A2(n13983), .A3(n13982), .ZN(n13985) );
  NAND3_X1 U16082 ( .A1(n15639), .A2(n13998), .A3(n13985), .ZN(n13986) );
  NAND3_X1 U16083 ( .A1(n13988), .A2(n13987), .A3(n13986), .ZN(P2_U3219) );
  OAI21_X1 U16084 ( .B1(n15592), .B2(n9280), .A(n13989), .ZN(n13990) );
  AOI21_X1 U16085 ( .B1(n13995), .B2(n15641), .A(n13990), .ZN(n14002) );
  MUX2_X1 U16086 ( .A(n11578), .B(P2_REG2_REG_6__SCAN_IN), .S(n13995), .Z(
        n13991) );
  NAND3_X1 U16087 ( .A1(n13993), .A2(n13992), .A3(n13991), .ZN(n13994) );
  NAND3_X1 U16088 ( .A1(n15644), .A2(n14009), .A3(n13994), .ZN(n14001) );
  MUX2_X1 U16089 ( .A(n10821), .B(P2_REG1_REG_6__SCAN_IN), .S(n13995), .Z(
        n13996) );
  NAND3_X1 U16090 ( .A1(n13998), .A2(n13997), .A3(n13996), .ZN(n13999) );
  NAND3_X1 U16091 ( .A1(n15639), .A2(n14014), .A3(n13999), .ZN(n14000) );
  NAND3_X1 U16092 ( .A1(n14002), .A2(n14001), .A3(n14000), .ZN(P2_U3220) );
  NOR2_X1 U16093 ( .A1(n14004), .A2(n14003), .ZN(n14005) );
  AOI211_X1 U16094 ( .C1(n15635), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n14006), .B(
        n14005), .ZN(n14018) );
  MUX2_X1 U16095 ( .A(n11601), .B(P2_REG2_REG_7__SCAN_IN), .S(n14011), .Z(
        n14007) );
  NAND3_X1 U16096 ( .A1(n14009), .A2(n14008), .A3(n14007), .ZN(n14010) );
  NAND3_X1 U16097 ( .A1(n15644), .A2(n14023), .A3(n14010), .ZN(n14017) );
  MUX2_X1 U16098 ( .A(n10824), .B(P2_REG1_REG_7__SCAN_IN), .S(n14011), .Z(
        n14012) );
  NAND3_X1 U16099 ( .A1(n14014), .A2(n14013), .A3(n14012), .ZN(n14015) );
  NAND3_X1 U16100 ( .A1(n15639), .A2(n14029), .A3(n14015), .ZN(n14016) );
  NAND3_X1 U16101 ( .A1(n14018), .A2(n14017), .A3(n14016), .ZN(P2_U3221) );
  OAI21_X1 U16102 ( .B1(n15592), .B2(n15129), .A(n14019), .ZN(n14020) );
  AOI21_X1 U16103 ( .B1(n14026), .B2(n15641), .A(n14020), .ZN(n14034) );
  MUX2_X1 U16104 ( .A(n11867), .B(P2_REG2_REG_8__SCAN_IN), .S(n14026), .Z(
        n14021) );
  NAND3_X1 U16105 ( .A1(n14023), .A2(n14022), .A3(n14021), .ZN(n14024) );
  NAND3_X1 U16106 ( .A1(n15644), .A2(n14025), .A3(n14024), .ZN(n14033) );
  MUX2_X1 U16107 ( .A(n10827), .B(P2_REG1_REG_8__SCAN_IN), .S(n14026), .Z(
        n14027) );
  NAND3_X1 U16108 ( .A1(n14029), .A2(n14028), .A3(n14027), .ZN(n14030) );
  NAND3_X1 U16109 ( .A1(n15639), .A2(n14031), .A3(n14030), .ZN(n14032) );
  NAND3_X1 U16110 ( .A1(n14034), .A2(n14033), .A3(n14032), .ZN(P2_U3222) );
  OAI21_X1 U16111 ( .B1(n15592), .B2(n15422), .A(n14035), .ZN(n14036) );
  AOI21_X1 U16112 ( .B1(n14040), .B2(n15641), .A(n14036), .ZN(n14048) );
  OAI21_X1 U16113 ( .B1(n14038), .B2(n14037), .A(n15583), .ZN(n14039) );
  NAND2_X1 U16114 ( .A1(n14039), .A2(n15644), .ZN(n14047) );
  MUX2_X1 U16115 ( .A(n12338), .B(P2_REG1_REG_11__SCAN_IN), .S(n14040), .Z(
        n14041) );
  NAND3_X1 U16116 ( .A1(n14043), .A2(n14042), .A3(n14041), .ZN(n14044) );
  NAND3_X1 U16117 ( .A1(n15639), .A2(n14045), .A3(n14044), .ZN(n14046) );
  NAND3_X1 U16118 ( .A1(n14048), .A2(n14047), .A3(n14046), .ZN(P2_U3225) );
  NAND2_X1 U16119 ( .A1(n14280), .A2(n15270), .ZN(n14055) );
  AND2_X1 U16120 ( .A1(n14053), .A2(n14052), .ZN(n14279) );
  INV_X1 U16121 ( .A(n14279), .ZN(n14283) );
  NOR2_X1 U16122 ( .A1(n15678), .A2(n14283), .ZN(n14059) );
  AOI21_X1 U16123 ( .B1(n15652), .B2(P2_REG2_REG_31__SCAN_IN), .A(n14059), 
        .ZN(n14054) );
  OAI211_X1 U16124 ( .C1(n14373), .C2(n15663), .A(n14055), .B(n14054), .ZN(
        P2_U3234) );
  OAI211_X1 U16125 ( .C1(n14377), .C2(n14057), .A(n14293), .B(n14056), .ZN(
        n14284) );
  NOR2_X1 U16126 ( .A1(n14377), .A2(n15663), .ZN(n14058) );
  AOI211_X1 U16127 ( .C1(n15652), .C2(P2_REG2_REG_30__SCAN_IN), .A(n14059), 
        .B(n14058), .ZN(n14060) );
  OAI21_X1 U16128 ( .B1(n15654), .B2(n14284), .A(n14060), .ZN(P2_U3235) );
  NOR2_X1 U16129 ( .A1(n14061), .A2(n15654), .ZN(n14066) );
  NOR2_X1 U16130 ( .A1(n15676), .A2(n14062), .ZN(n14063) );
  AOI21_X1 U16131 ( .B1(n15652), .B2(P2_REG2_REG_29__SCAN_IN), .A(n14063), 
        .ZN(n14064) );
  OAI21_X1 U16132 ( .B1(n14291), .B2(n15663), .A(n14064), .ZN(n14065) );
  OAI21_X1 U16133 ( .B1(n14069), .B2(n15678), .A(n14068), .ZN(P2_U3236) );
  XNOR2_X1 U16134 ( .A(n14071), .B(n14070), .ZN(n14297) );
  AOI21_X1 U16135 ( .B1(n14084), .B2(n14073), .A(n14072), .ZN(n14074) );
  NOR3_X1 U16136 ( .A1(n14074), .A2(n6745), .A3(n15668), .ZN(n14076) );
  NOR2_X1 U16137 ( .A1(n14076), .A2(n14075), .ZN(n14296) );
  AOI21_X1 U16138 ( .B1(n14292), .B2(n14090), .A(n14077), .ZN(n14294) );
  NAND2_X1 U16139 ( .A1(n14294), .A2(n14078), .ZN(n14079) );
  OAI211_X1 U16140 ( .C1(n15676), .C2(n14080), .A(n14296), .B(n14079), .ZN(
        n14081) );
  NAND2_X1 U16141 ( .A1(n14081), .A2(n15659), .ZN(n14083) );
  AOI22_X1 U16142 ( .A1(n14292), .A2(n15261), .B1(n15652), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n14082) );
  OAI211_X1 U16143 ( .C1(n14261), .C2(n14297), .A(n14083), .B(n14082), .ZN(
        P2_U3237) );
  OAI21_X1 U16144 ( .B1(n14085), .B2(n14088), .A(n14084), .ZN(n14087) );
  NAND2_X1 U16145 ( .A1(n14300), .A2(n15269), .ZN(n14097) );
  AOI211_X1 U16146 ( .C1(n14091), .C2(n14104), .A(n15263), .B(n9746), .ZN(
        n14299) );
  INV_X1 U16147 ( .A(n14091), .ZN(n14381) );
  INV_X1 U16148 ( .A(n14092), .ZN(n14093) );
  AOI22_X1 U16149 ( .A1(n15652), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n14093), 
        .B2(n15260), .ZN(n14094) );
  OAI21_X1 U16150 ( .B1(n14381), .B2(n15663), .A(n14094), .ZN(n14095) );
  AOI21_X1 U16151 ( .B1(n14299), .B2(n15270), .A(n14095), .ZN(n14096) );
  OAI211_X1 U16152 ( .C1(n15678), .C2(n14298), .A(n14097), .B(n14096), .ZN(
        P2_U3238) );
  INV_X1 U16153 ( .A(n14102), .ZN(n14098) );
  XNOR2_X1 U16154 ( .A(n14099), .B(n14098), .ZN(n14101) );
  AOI21_X1 U16155 ( .B1(n14101), .B2(n15256), .A(n14100), .ZN(n14304) );
  XNOR2_X1 U16156 ( .A(n14103), .B(n14102), .ZN(n14302) );
  OAI211_X1 U16157 ( .C1(n14385), .C2(n14125), .A(n14293), .B(n14104), .ZN(
        n14303) );
  NAND2_X1 U16158 ( .A1(n15652), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n14105) );
  OAI21_X1 U16159 ( .B1(n15676), .B2(n14106), .A(n14105), .ZN(n14107) );
  AOI21_X1 U16160 ( .B1(n14108), .B2(n15261), .A(n14107), .ZN(n14109) );
  OAI21_X1 U16161 ( .B1(n14303), .B2(n15654), .A(n14109), .ZN(n14110) );
  AOI21_X1 U16162 ( .B1(n14302), .B2(n15269), .A(n14110), .ZN(n14111) );
  OAI21_X1 U16163 ( .B1(n15652), .B2(n14304), .A(n14111), .ZN(P2_U3239) );
  XNOR2_X1 U16164 ( .A(n14113), .B(n14112), .ZN(n14115) );
  AOI21_X1 U16165 ( .B1(n14115), .B2(n15256), .A(n14114), .ZN(n14312) );
  OAI21_X1 U16166 ( .B1(n14118), .B2(n14117), .A(n14116), .ZN(n14119) );
  INV_X1 U16167 ( .A(n14119), .ZN(n14313) );
  NAND2_X1 U16168 ( .A1(n15652), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n14120) );
  OAI21_X1 U16169 ( .B1(n15676), .B2(n14121), .A(n14120), .ZN(n14122) );
  AOI21_X1 U16170 ( .B1(n14310), .B2(n15261), .A(n14122), .ZN(n14127) );
  NAND2_X1 U16171 ( .A1(n14310), .A2(n14134), .ZN(n14123) );
  NAND2_X1 U16172 ( .A1(n14123), .A2(n14293), .ZN(n14124) );
  NOR2_X1 U16173 ( .A1(n14125), .A2(n14124), .ZN(n14309) );
  NAND2_X1 U16174 ( .A1(n14309), .A2(n15270), .ZN(n14126) );
  OAI211_X1 U16175 ( .C1(n14313), .C2(n14261), .A(n14127), .B(n14126), .ZN(
        n14128) );
  INV_X1 U16176 ( .A(n14128), .ZN(n14129) );
  OAI21_X1 U16177 ( .B1(n15652), .B2(n14312), .A(n14129), .ZN(P2_U3240) );
  XNOR2_X1 U16178 ( .A(n14130), .B(n14139), .ZN(n14132) );
  AOI21_X1 U16179 ( .B1(n14132), .B2(n15256), .A(n14131), .ZN(n14319) );
  INV_X1 U16180 ( .A(n14319), .ZN(n14138) );
  AOI21_X1 U16181 ( .B1(n14316), .B2(n14133), .A(n15263), .ZN(n14135) );
  NAND2_X1 U16182 ( .A1(n14135), .A2(n14134), .ZN(n14317) );
  OAI22_X1 U16183 ( .A1(n14317), .A2(n14272), .B1(n15676), .B2(n14136), .ZN(
        n14137) );
  OAI21_X1 U16184 ( .B1(n14138), .B2(n14137), .A(n15659), .ZN(n14143) );
  AOI22_X1 U16185 ( .A1(n14316), .A2(n15261), .B1(n15652), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n14142) );
  NAND2_X1 U16186 ( .A1(n14140), .A2(n14139), .ZN(n14314) );
  NAND3_X1 U16187 ( .A1(n14315), .A2(n15269), .A3(n14314), .ZN(n14141) );
  NAND3_X1 U16188 ( .A1(n14143), .A2(n14142), .A3(n14141), .ZN(P2_U3241) );
  NAND2_X1 U16189 ( .A1(n14145), .A2(n14144), .ZN(n14146) );
  NAND2_X1 U16190 ( .A1(n14147), .A2(n14146), .ZN(n14321) );
  INV_X1 U16191 ( .A(n14321), .ZN(n14162) );
  NAND2_X1 U16192 ( .A1(n14148), .A2(n7008), .ZN(n14149) );
  NAND2_X1 U16193 ( .A1(n14150), .A2(n14149), .ZN(n14151) );
  NAND2_X1 U16194 ( .A1(n14151), .A2(n15256), .ZN(n14323) );
  INV_X1 U16195 ( .A(n14323), .ZN(n14158) );
  XNOR2_X1 U16196 ( .A(n6706), .B(n14391), .ZN(n14154) );
  INV_X1 U16197 ( .A(n14152), .ZN(n14153) );
  AOI21_X1 U16198 ( .B1(n14154), .B2(n14293), .A(n14153), .ZN(n14322) );
  INV_X1 U16199 ( .A(n14155), .ZN(n14156) );
  OAI22_X1 U16200 ( .A1(n14322), .A2(n14272), .B1(n15676), .B2(n14156), .ZN(
        n14157) );
  OAI21_X1 U16201 ( .B1(n14158), .B2(n14157), .A(n15659), .ZN(n14161) );
  AOI22_X1 U16202 ( .A1(n14159), .A2(n15261), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n15678), .ZN(n14160) );
  OAI211_X1 U16203 ( .C1(n14162), .C2(n14261), .A(n14161), .B(n14160), .ZN(
        P2_U3242) );
  OR2_X1 U16204 ( .A1(n14163), .A2(n14166), .ZN(n14164) );
  NAND2_X1 U16205 ( .A1(n14165), .A2(n14164), .ZN(n14331) );
  NAND2_X1 U16206 ( .A1(n14167), .A2(n14166), .ZN(n14168) );
  NAND3_X1 U16207 ( .A1(n14169), .A2(n15256), .A3(n14168), .ZN(n14171) );
  NAND2_X1 U16208 ( .A1(n14171), .A2(n14170), .ZN(n14329) );
  INV_X1 U16209 ( .A(n14394), .ZN(n14176) );
  AOI21_X1 U16210 ( .B1(n14186), .B2(n14394), .A(n15263), .ZN(n14172) );
  AND2_X1 U16211 ( .A1(n14172), .A2(n6706), .ZN(n14328) );
  NAND2_X1 U16212 ( .A1(n14328), .A2(n15270), .ZN(n14175) );
  AOI22_X1 U16213 ( .A1(n14173), .A2(n15260), .B1(n15652), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n14174) );
  OAI211_X1 U16214 ( .C1(n14176), .C2(n15663), .A(n14175), .B(n14174), .ZN(
        n14177) );
  AOI21_X1 U16215 ( .B1(n14329), .B2(n15659), .A(n14177), .ZN(n14178) );
  OAI21_X1 U16216 ( .B1(n14261), .B2(n14331), .A(n14178), .ZN(P2_U3243) );
  XNOR2_X1 U16217 ( .A(n14180), .B(n14179), .ZN(n14339) );
  XNOR2_X1 U16218 ( .A(n14182), .B(n14181), .ZN(n14184) );
  OAI21_X1 U16219 ( .B1(n14184), .B2(n15668), .A(n14183), .ZN(n14335) );
  OR2_X1 U16220 ( .A1(n14204), .A2(n14191), .ZN(n14185) );
  NAND2_X1 U16221 ( .A1(n14336), .A2(n15270), .ZN(n14190) );
  INV_X1 U16222 ( .A(n14187), .ZN(n14188) );
  AOI22_X1 U16223 ( .A1(P2_REG2_REG_21__SCAN_IN), .A2(n15678), .B1(n14188), 
        .B2(n15260), .ZN(n14189) );
  OAI211_X1 U16224 ( .C1(n14191), .C2(n15663), .A(n14190), .B(n14189), .ZN(
        n14192) );
  AOI21_X1 U16225 ( .B1(n14335), .B2(n15659), .A(n14192), .ZN(n14193) );
  OAI21_X1 U16226 ( .B1(n14261), .B2(n14339), .A(n14193), .ZN(P2_U3244) );
  XNOR2_X1 U16227 ( .A(n14195), .B(n14194), .ZN(n14344) );
  OAI21_X1 U16228 ( .B1(n14198), .B2(n14197), .A(n14196), .ZN(n14201) );
  INV_X1 U16229 ( .A(n14199), .ZN(n14200) );
  AOI21_X1 U16230 ( .B1(n14201), .B2(n15256), .A(n14200), .ZN(n14343) );
  INV_X1 U16231 ( .A(n14343), .ZN(n14210) );
  INV_X1 U16232 ( .A(n14341), .ZN(n14208) );
  NAND2_X1 U16233 ( .A1(n14223), .A2(n14341), .ZN(n14202) );
  NAND2_X1 U16234 ( .A1(n14202), .A2(n14293), .ZN(n14203) );
  NOR2_X1 U16235 ( .A1(n14204), .A2(n14203), .ZN(n14340) );
  NAND2_X1 U16236 ( .A1(n14340), .A2(n15270), .ZN(n14207) );
  AOI22_X1 U16237 ( .A1(n15652), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14205), 
        .B2(n15260), .ZN(n14206) );
  OAI211_X1 U16238 ( .C1(n14208), .C2(n15663), .A(n14207), .B(n14206), .ZN(
        n14209) );
  AOI21_X1 U16239 ( .B1(n14210), .B2(n15659), .A(n14209), .ZN(n14211) );
  OAI21_X1 U16240 ( .B1(n14344), .B2(n14261), .A(n14211), .ZN(P2_U3245) );
  INV_X1 U16241 ( .A(n14212), .ZN(n14214) );
  AOI22_X1 U16242 ( .A1(n14222), .A2(n14215), .B1(n14214), .B2(n14213), .ZN(
        n14217) );
  OAI21_X1 U16243 ( .B1(n14217), .B2(n15668), .A(n14216), .ZN(n14346) );
  NAND2_X1 U16244 ( .A1(n14346), .A2(n15659), .ZN(n14228) );
  NAND2_X1 U16245 ( .A1(n15652), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n14218) );
  OAI21_X1 U16246 ( .B1(n15676), .B2(n14219), .A(n14218), .ZN(n14220) );
  AOI21_X1 U16247 ( .B1(n14345), .B2(n15261), .A(n14220), .ZN(n14227) );
  XNOR2_X1 U16248 ( .A(n14222), .B(n14221), .ZN(n14348) );
  NAND2_X1 U16249 ( .A1(n14348), .A2(n15269), .ZN(n14226) );
  AOI21_X1 U16250 ( .B1(n14345), .B2(n14232), .A(n15263), .ZN(n14224) );
  AND2_X1 U16251 ( .A1(n14224), .A2(n14223), .ZN(n14347) );
  NAND2_X1 U16252 ( .A1(n14347), .A2(n15270), .ZN(n14225) );
  NAND4_X1 U16253 ( .A1(n14228), .A2(n14227), .A3(n14226), .A4(n14225), .ZN(
        P2_U3246) );
  XNOR2_X1 U16254 ( .A(n14229), .B(n14238), .ZN(n14231) );
  AOI21_X1 U16255 ( .B1(n14231), .B2(n15256), .A(n14230), .ZN(n14354) );
  AOI211_X1 U16256 ( .C1(n14353), .C2(n14258), .A(n15263), .B(n7467), .ZN(
        n14352) );
  INV_X1 U16257 ( .A(n14233), .ZN(n14234) );
  AOI22_X1 U16258 ( .A1(n15652), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14234), 
        .B2(n15260), .ZN(n14235) );
  OAI21_X1 U16259 ( .B1(n14236), .B2(n15663), .A(n14235), .ZN(n14241) );
  OAI21_X1 U16260 ( .B1(n14238), .B2(n6824), .A(n14237), .ZN(n14239) );
  INV_X1 U16261 ( .A(n14239), .ZN(n14356) );
  NOR2_X1 U16262 ( .A1(n14356), .A2(n14261), .ZN(n14240) );
  AOI211_X1 U16263 ( .C1(n14352), .C2(n15270), .A(n14241), .B(n14240), .ZN(
        n14242) );
  OAI21_X1 U16264 ( .B1(n15678), .B2(n14354), .A(n14242), .ZN(P2_U3247) );
  OAI211_X1 U16265 ( .C1(n14245), .C2(n14244), .A(n14243), .B(n15256), .ZN(
        n14248) );
  INV_X1 U16266 ( .A(n14246), .ZN(n14247) );
  NAND2_X1 U16267 ( .A1(n14248), .A2(n14247), .ZN(n14357) );
  OR2_X1 U16268 ( .A1(n14249), .A2(n7136), .ZN(n14251) );
  NAND2_X1 U16269 ( .A1(n14251), .A2(n14250), .ZN(n14361) );
  NAND2_X1 U16270 ( .A1(n15678), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n14252) );
  OAI21_X1 U16271 ( .B1(n15676), .B2(n14253), .A(n14252), .ZN(n14254) );
  AOI21_X1 U16272 ( .B1(n14359), .B2(n15261), .A(n14254), .ZN(n14260) );
  OR2_X1 U16273 ( .A1(n14256), .A2(n14255), .ZN(n14257) );
  AND3_X1 U16274 ( .A1(n14258), .A2(n14257), .A3(n14293), .ZN(n14358) );
  NAND2_X1 U16275 ( .A1(n14358), .A2(n15270), .ZN(n14259) );
  OAI211_X1 U16276 ( .C1(n14361), .C2(n14261), .A(n14260), .B(n14259), .ZN(
        n14262) );
  AOI21_X1 U16277 ( .B1(n15659), .B2(n14357), .A(n14262), .ZN(n14263) );
  INV_X1 U16278 ( .A(n14263), .ZN(P2_U3248) );
  XNOR2_X1 U16279 ( .A(n14264), .B(n14274), .ZN(n14265) );
  NAND2_X1 U16280 ( .A1(n14265), .A2(n15256), .ZN(n14268) );
  INV_X1 U16281 ( .A(n14266), .ZN(n14267) );
  NAND2_X1 U16282 ( .A1(n14268), .A2(n14267), .ZN(n14368) );
  XNOR2_X1 U16283 ( .A(n14364), .B(n14269), .ZN(n14270) );
  OR2_X1 U16284 ( .A1(n14270), .A2(n15263), .ZN(n14365) );
  OAI22_X1 U16285 ( .A1(n14365), .A2(n14272), .B1(n15676), .B2(n14271), .ZN(
        n14273) );
  OAI21_X1 U16286 ( .B1(n14368), .B2(n14273), .A(n15659), .ZN(n14278) );
  AOI22_X1 U16287 ( .A1(n14364), .A2(n15261), .B1(n15652), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n14277) );
  NAND2_X1 U16288 ( .A1(n14275), .A2(n14274), .ZN(n14362) );
  NAND3_X1 U16289 ( .A1(n14363), .A2(n14362), .A3(n15269), .ZN(n14276) );
  NAND3_X1 U16290 ( .A1(n14278), .A2(n14277), .A3(n14276), .ZN(P2_U3249) );
  NOR2_X1 U16291 ( .A1(n14280), .A2(n14279), .ZN(n14370) );
  MUX2_X1 U16292 ( .A(n14281), .B(n14370), .S(n15731), .Z(n14282) );
  OAI21_X1 U16293 ( .B1(n14373), .B2(n14351), .A(n14282), .ZN(P2_U3530) );
  AND2_X1 U16294 ( .A1(n14284), .A2(n14283), .ZN(n14374) );
  MUX2_X1 U16295 ( .A(n14285), .B(n14374), .S(n15731), .Z(n14286) );
  OAI21_X1 U16296 ( .B1(n14377), .B2(n14351), .A(n14286), .ZN(P2_U3529) );
  NAND2_X1 U16297 ( .A1(n15729), .A2(n14288), .ZN(n14289) );
  OAI21_X1 U16298 ( .B1(n14291), .B2(n14351), .A(n14290), .ZN(P2_U3528) );
  AOI22_X1 U16299 ( .A1(n14294), .A2(n14293), .B1(n15281), .B2(n14292), .ZN(
        n14295) );
  OAI211_X1 U16300 ( .C1(n15285), .C2(n14297), .A(n14296), .B(n14295), .ZN(
        n14378) );
  MUX2_X1 U16301 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n14378), .S(n15731), .Z(
        P2_U3527) );
  INV_X1 U16302 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n14301) );
  NAND2_X1 U16303 ( .A1(n14302), .A2(n15722), .ZN(n14306) );
  AND2_X1 U16304 ( .A1(n14304), .A2(n14303), .ZN(n14305) );
  NAND2_X1 U16305 ( .A1(n14306), .A2(n14305), .ZN(n14382) );
  MUX2_X1 U16306 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14382), .S(n15731), .Z(
        n14307) );
  INV_X1 U16307 ( .A(n14307), .ZN(n14308) );
  OAI21_X1 U16308 ( .B1(n14385), .B2(n14351), .A(n14308), .ZN(P2_U3525) );
  AOI21_X1 U16309 ( .B1(n15281), .B2(n14310), .A(n14309), .ZN(n14311) );
  OAI211_X1 U16310 ( .C1(n14313), .C2(n15285), .A(n14312), .B(n14311), .ZN(
        n14386) );
  MUX2_X1 U16311 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14386), .S(n15731), .Z(
        P2_U3524) );
  NAND3_X1 U16312 ( .A1(n14315), .A2(n15722), .A3(n14314), .ZN(n14320) );
  NAND2_X1 U16313 ( .A1(n14316), .A2(n15281), .ZN(n14318) );
  NAND4_X1 U16314 ( .A1(n14320), .A2(n14319), .A3(n14318), .A4(n14317), .ZN(
        n14387) );
  MUX2_X1 U16315 ( .A(n14387), .B(P2_REG1_REG_24__SCAN_IN), .S(n15729), .Z(
        P2_U3523) );
  NAND2_X1 U16316 ( .A1(n14321), .A2(n15722), .ZN(n14325) );
  AND2_X1 U16317 ( .A1(n14323), .A2(n14322), .ZN(n14324) );
  NAND2_X1 U16318 ( .A1(n14325), .A2(n14324), .ZN(n14388) );
  MUX2_X1 U16319 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14388), .S(n15731), .Z(
        n14326) );
  INV_X1 U16320 ( .A(n14326), .ZN(n14327) );
  OAI21_X1 U16321 ( .B1(n14391), .B2(n14351), .A(n14327), .ZN(P2_U3522) );
  NOR2_X1 U16322 ( .A1(n14329), .A2(n14328), .ZN(n14330) );
  OAI21_X1 U16323 ( .B1(n14331), .B2(n15285), .A(n14330), .ZN(n14392) );
  MUX2_X1 U16324 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14392), .S(n15731), .Z(
        n14332) );
  AOI21_X1 U16325 ( .B1(n14333), .B2(n14394), .A(n14332), .ZN(n14334) );
  INV_X1 U16326 ( .A(n14334), .ZN(P2_U3521) );
  AOI211_X1 U16327 ( .C1(n15281), .C2(n14337), .A(n14336), .B(n14335), .ZN(
        n14338) );
  OAI21_X1 U16328 ( .B1(n15285), .B2(n14339), .A(n14338), .ZN(n14396) );
  MUX2_X1 U16329 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14396), .S(n15731), .Z(
        P2_U3520) );
  AOI21_X1 U16330 ( .B1(n15281), .B2(n14341), .A(n14340), .ZN(n14342) );
  OAI211_X1 U16331 ( .C1(n14344), .C2(n15285), .A(n14343), .B(n14342), .ZN(
        n14397) );
  MUX2_X1 U16332 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14397), .S(n15731), .Z(
        P2_U3519) );
  AOI211_X1 U16333 ( .C1(n14348), .C2(n15722), .A(n14347), .B(n14346), .ZN(
        n14398) );
  MUX2_X1 U16334 ( .A(n14349), .B(n14398), .S(n15731), .Z(n14350) );
  OAI21_X1 U16335 ( .B1(n7466), .B2(n14351), .A(n14350), .ZN(P2_U3518) );
  AOI21_X1 U16336 ( .B1(n15281), .B2(n14353), .A(n14352), .ZN(n14355) );
  OAI211_X1 U16337 ( .C1(n15285), .C2(n14356), .A(n14355), .B(n14354), .ZN(
        n14402) );
  MUX2_X1 U16338 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14402), .S(n15731), .Z(
        P2_U3517) );
  AOI211_X1 U16339 ( .C1(n15281), .C2(n14359), .A(n14358), .B(n14357), .ZN(
        n14360) );
  OAI21_X1 U16340 ( .B1(n15285), .B2(n14361), .A(n14360), .ZN(n14403) );
  MUX2_X1 U16341 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14403), .S(n15731), .Z(
        P2_U3516) );
  NAND3_X1 U16342 ( .A1(n14363), .A2(n14362), .A3(n15722), .ZN(n14367) );
  NAND2_X1 U16343 ( .A1(n14364), .A2(n15281), .ZN(n14366) );
  NAND3_X1 U16344 ( .A1(n14367), .A2(n14366), .A3(n14365), .ZN(n14369) );
  MUX2_X1 U16345 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14404), .S(n15731), .Z(
        P2_U3515) );
  INV_X1 U16346 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n14371) );
  MUX2_X1 U16347 ( .A(n14371), .B(n14370), .S(n15724), .Z(n14372) );
  INV_X1 U16348 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n14375) );
  MUX2_X1 U16349 ( .A(n14375), .B(n14374), .S(n15724), .Z(n14376) );
  OAI21_X1 U16350 ( .B1(n14377), .B2(n14401), .A(n14376), .ZN(P2_U3497) );
  MUX2_X1 U16351 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n14378), .S(n15724), .Z(
        P2_U3495) );
  INV_X1 U16352 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n14380) );
  MUX2_X1 U16353 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14382), .S(n15724), .Z(
        n14383) );
  INV_X1 U16354 ( .A(n14383), .ZN(n14384) );
  OAI21_X1 U16355 ( .B1(n14385), .B2(n14401), .A(n14384), .ZN(P2_U3493) );
  MUX2_X1 U16356 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14386), .S(n15724), .Z(
        P2_U3492) );
  MUX2_X1 U16357 ( .A(n14387), .B(P2_REG0_REG_24__SCAN_IN), .S(n9771), .Z(
        P2_U3491) );
  MUX2_X1 U16358 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14388), .S(n15724), .Z(
        n14389) );
  INV_X1 U16359 ( .A(n14389), .ZN(n14390) );
  OAI21_X1 U16360 ( .B1(n14391), .B2(n14401), .A(n14390), .ZN(P2_U3490) );
  MUX2_X1 U16361 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14392), .S(n15724), .Z(
        n14393) );
  AOI21_X1 U16362 ( .B1(n9774), .B2(n14394), .A(n14393), .ZN(n14395) );
  INV_X1 U16363 ( .A(n14395), .ZN(P2_U3489) );
  MUX2_X1 U16364 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14396), .S(n15724), .Z(
        P2_U3488) );
  MUX2_X1 U16365 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14397), .S(n15724), .Z(
        P2_U3487) );
  INV_X1 U16366 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14399) );
  MUX2_X1 U16367 ( .A(n14399), .B(n14398), .S(n15724), .Z(n14400) );
  OAI21_X1 U16368 ( .B1(n7466), .B2(n14401), .A(n14400), .ZN(P2_U3486) );
  MUX2_X1 U16369 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14402), .S(n15724), .Z(
        P2_U3484) );
  MUX2_X1 U16370 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14403), .S(n15724), .Z(
        P2_U3481) );
  MUX2_X1 U16371 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14404), .S(n15724), .Z(
        P2_U3478) );
  INV_X1 U16372 ( .A(n10409), .ZN(n14410) );
  INV_X1 U16373 ( .A(n14405), .ZN(n14407) );
  NOR4_X1 U16374 ( .A1(n14407), .A2(P2_IR_REG_30__SCAN_IN), .A3(n14406), .A4(
        P2_U3088), .ZN(n14408) );
  AOI21_X1 U16375 ( .B1(n14421), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14408), 
        .ZN(n14409) );
  OAI21_X1 U16376 ( .B1(n14410), .B2(n14428), .A(n14409), .ZN(P2_U3296) );
  OAI222_X1 U16377 ( .A1(n14428), .A2(n14413), .B1(n14412), .B2(P2_U3088), 
        .C1(n14411), .C2(n14434), .ZN(P2_U3298) );
  NAND2_X1 U16378 ( .A1(n14415), .A2(n14414), .ZN(n14417) );
  OAI211_X1 U16379 ( .C1(n14434), .C2(n14418), .A(n14417), .B(n14416), .ZN(
        P2_U3299) );
  INV_X1 U16380 ( .A(n14419), .ZN(n15093) );
  AOI21_X1 U16381 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n14421), .A(n14420), 
        .ZN(n14422) );
  OAI21_X1 U16382 ( .B1(n15093), .B2(n14428), .A(n14422), .ZN(P2_U3300) );
  INV_X1 U16383 ( .A(n14423), .ZN(n15096) );
  OAI222_X1 U16384 ( .A1(n14434), .A2(n14425), .B1(n14424), .B2(P2_U3088), 
        .C1(n14428), .C2(n15096), .ZN(P2_U3301) );
  INV_X1 U16385 ( .A(n14426), .ZN(n15099) );
  OAI222_X1 U16386 ( .A1(n14434), .A2(n14429), .B1(n14428), .B2(n15099), .C1(
        P2_U3088), .C2(n14427), .ZN(P2_U3302) );
  INV_X1 U16387 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n14433) );
  INV_X1 U16388 ( .A(n14430), .ZN(n15103) );
  OAI222_X1 U16389 ( .A1(n14434), .A2(n14433), .B1(n14428), .B2(n15103), .C1(
        P2_U3088), .C2(n14431), .ZN(P2_U3303) );
  MUX2_X1 U16390 ( .A(n14435), .B(n15565), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3327) );
  NAND2_X1 U16391 ( .A1(n14437), .A2(n15365), .ZN(n14442) );
  NOR2_X1 U16392 ( .A1(n15369), .A2(n14799), .ZN(n14440) );
  INV_X1 U16393 ( .A(n14789), .ZN(n14438) );
  OAI22_X1 U16394 ( .A1(n14761), .A2(n15361), .B1(n15360), .B2(n14438), .ZN(
        n14439) );
  AOI211_X1 U16395 ( .C1(P1_REG3_REG_27__SCAN_IN), .C2(P1_U3086), .A(n14440), 
        .B(n14439), .ZN(n14441) );
  OAI211_X1 U16396 ( .C1(n15001), .C2(n15358), .A(n14442), .B(n14441), .ZN(
        P1_U3214) );
  OR2_X1 U16397 ( .A1(n14714), .A2(n14966), .ZN(n14444) );
  NAND2_X1 U16398 ( .A1(n14826), .A2(n14827), .ZN(n14443) );
  NAND2_X1 U16399 ( .A1(n14444), .A2(n14443), .ZN(n15023) );
  AOI22_X1 U16400 ( .A1(n15348), .A2(n15023), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14445) );
  OAI21_X1 U16401 ( .B1(n14866), .B2(n15369), .A(n14445), .ZN(n14453) );
  INV_X1 U16402 ( .A(n14448), .ZN(n14449) );
  NAND3_X1 U16403 ( .A1(n14447), .A2(n14450), .A3(n14449), .ZN(n14451) );
  AOI21_X1 U16404 ( .B1(n14446), .B2(n14451), .A(n15337), .ZN(n14452) );
  AOI211_X1 U16405 ( .C1(n15024), .C2(n15351), .A(n14453), .B(n14452), .ZN(
        n14454) );
  INV_X1 U16406 ( .A(n14454), .ZN(P1_U3216) );
  INV_X1 U16407 ( .A(n15052), .ZN(n14926) );
  OAI21_X1 U16408 ( .B1(n6707), .B2(n14456), .A(n14455), .ZN(n14458) );
  NAND3_X1 U16409 ( .A1(n14458), .A2(n15365), .A3(n14457), .ZN(n14462) );
  OAI22_X1 U16410 ( .A1(n14710), .A2(n14967), .B1(n14489), .B2(n14966), .ZN(
        n15051) );
  NOR2_X1 U16411 ( .A1(n14459), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14684) );
  NOR2_X1 U16412 ( .A1(n15369), .A2(n14921), .ZN(n14460) );
  AOI211_X1 U16413 ( .C1(n15051), .C2(n15348), .A(n14684), .B(n14460), .ZN(
        n14461) );
  OAI211_X1 U16414 ( .C1(n14926), .C2(n15358), .A(n14462), .B(n14461), .ZN(
        P1_U3219) );
  INV_X1 U16415 ( .A(n14463), .ZN(n14464) );
  AOI21_X1 U16416 ( .B1(n14466), .B2(n14465), .A(n14464), .ZN(n14471) );
  INV_X1 U16417 ( .A(n14895), .ZN(n14468) );
  OAI22_X1 U16418 ( .A1(n14710), .A2(n14966), .B1(n14714), .B2(n14967), .ZN(
        n15040) );
  AOI22_X1 U16419 ( .A1(n15040), .A2(n15348), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14467) );
  OAI21_X1 U16420 ( .B1(n14468), .B2(n15369), .A(n14467), .ZN(n14469) );
  AOI21_X1 U16421 ( .B1(n15041), .B2(n15351), .A(n14469), .ZN(n14470) );
  OAI21_X1 U16422 ( .B1(n14471), .B2(n15337), .A(n14470), .ZN(P1_U3223) );
  INV_X1 U16423 ( .A(n14472), .ZN(n14473) );
  NOR2_X1 U16424 ( .A1(n14474), .A2(n14473), .ZN(n14478) );
  INV_X1 U16425 ( .A(n14476), .ZN(n14477) );
  AOI21_X1 U16426 ( .B1(n14478), .B2(n14475), .A(n14477), .ZN(n14484) );
  INV_X1 U16427 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14479) );
  OAI22_X1 U16428 ( .A1(n15369), .A2(n14833), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14479), .ZN(n14482) );
  OAI22_X1 U16429 ( .A1(n14480), .A2(n15361), .B1(n15360), .B2(n14761), .ZN(
        n14481) );
  AOI211_X1 U16430 ( .C1(n15014), .C2(n15351), .A(n14482), .B(n14481), .ZN(
        n14483) );
  OAI21_X1 U16431 ( .B1(n14484), .B2(n15337), .A(n14483), .ZN(P1_U3225) );
  XNOR2_X1 U16432 ( .A(n14487), .B(n14486), .ZN(n14488) );
  XNOR2_X1 U16433 ( .A(n14485), .B(n14488), .ZN(n14494) );
  OAI22_X1 U16434 ( .A1(n14489), .A2(n14967), .B1(n15359), .B2(n14966), .ZN(
        n15063) );
  NAND2_X1 U16435 ( .A1(n15063), .A2(n15348), .ZN(n14491) );
  OAI211_X1 U16436 ( .C1(n15369), .C2(n14953), .A(n14491), .B(n14490), .ZN(
        n14492) );
  AOI21_X1 U16437 ( .B1(n15064), .B2(n15351), .A(n14492), .ZN(n14493) );
  OAI21_X1 U16438 ( .B1(n14494), .B2(n15337), .A(n14493), .ZN(P1_U3228) );
  INV_X1 U16439 ( .A(n14495), .ZN(n14496) );
  NOR2_X1 U16440 ( .A1(n14497), .A2(n14496), .ZN(n14499) );
  INV_X1 U16441 ( .A(n14475), .ZN(n14498) );
  AOI21_X1 U16442 ( .B1(n14499), .B2(n14446), .A(n14498), .ZN(n14504) );
  INV_X1 U16443 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14500) );
  OAI22_X1 U16444 ( .A1(n15369), .A2(n14854), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14500), .ZN(n14502) );
  INV_X1 U16445 ( .A(n14717), .ZN(n14845) );
  OAI22_X1 U16446 ( .A1(n14845), .A2(n15361), .B1(n15360), .B2(n14846), .ZN(
        n14501) );
  AOI211_X1 U16447 ( .C1(n14859), .C2(n15351), .A(n14502), .B(n14501), .ZN(
        n14503) );
  OAI21_X1 U16448 ( .B1(n14504), .B2(n15337), .A(n14503), .ZN(P1_U3229) );
  OAI211_X1 U16449 ( .C1(n14507), .C2(n14506), .A(n14505), .B(n15365), .ZN(
        n14513) );
  AOI22_X1 U16450 ( .A1(n15351), .A2(n14508), .B1(P1_REG3_REG_4__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14512) );
  OR2_X1 U16451 ( .A1(n15369), .A2(n14509), .ZN(n14511) );
  NAND2_X1 U16452 ( .A1(n15348), .A2(n15525), .ZN(n14510) );
  NAND4_X1 U16453 ( .A1(n14513), .A2(n14512), .A3(n14511), .A4(n14510), .ZN(
        P1_U3230) );
  XNOR2_X1 U16454 ( .A(n14515), .B(n14514), .ZN(n14521) );
  NAND2_X1 U16455 ( .A1(n14712), .A2(n14827), .ZN(n14517) );
  NAND2_X1 U16456 ( .A1(n14709), .A2(n14825), .ZN(n14516) );
  NAND2_X1 U16457 ( .A1(n14517), .A2(n14516), .ZN(n14902) );
  AOI22_X1 U16458 ( .A1(n14902), .A2(n15348), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14518) );
  OAI21_X1 U16459 ( .B1(n14908), .B2(n15369), .A(n14518), .ZN(n14519) );
  AOI21_X1 U16460 ( .B1(n15046), .B2(n15351), .A(n14519), .ZN(n14520) );
  OAI21_X1 U16461 ( .B1(n14521), .B2(n15337), .A(n14520), .ZN(P1_U3233) );
  INV_X1 U16462 ( .A(n14712), .ZN(n14752) );
  OAI22_X1 U16463 ( .A1(n14752), .A2(n14966), .B1(n14845), .B2(n14967), .ZN(
        n15032) );
  AOI22_X1 U16464 ( .A1(n15032), .A2(n15348), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14522) );
  OAI21_X1 U16465 ( .B1(n14880), .B2(n15369), .A(n14522), .ZN(n14528) );
  INV_X1 U16466 ( .A(n14523), .ZN(n14524) );
  NAND3_X1 U16467 ( .A1(n14463), .A2(n14525), .A3(n14524), .ZN(n14526) );
  AOI21_X1 U16468 ( .B1(n14447), .B2(n14526), .A(n15337), .ZN(n14527) );
  AOI211_X1 U16469 ( .C1(n15033), .C2(n15351), .A(n14528), .B(n14527), .ZN(
        n14529) );
  INV_X1 U16470 ( .A(n14529), .ZN(P1_U3235) );
  AOI21_X1 U16471 ( .B1(n14531), .B2(n14530), .A(n6707), .ZN(n14538) );
  AOI22_X1 U16472 ( .A1(n14825), .A2(n14705), .B1(n14709), .B2(n14827), .ZN(
        n14939) );
  INV_X1 U16473 ( .A(n15348), .ZN(n14535) );
  NAND2_X1 U16474 ( .A1(n14532), .A2(n14942), .ZN(n14533) );
  OAI211_X1 U16475 ( .C1(n14939), .C2(n14535), .A(n14534), .B(n14533), .ZN(
        n14536) );
  AOI21_X1 U16476 ( .B1(n15057), .B2(n15351), .A(n14536), .ZN(n14537) );
  OAI21_X1 U16477 ( .B1(n14538), .B2(n15337), .A(n14537), .ZN(P1_U3238) );
  OAI21_X1 U16478 ( .B1(n14541), .B2(n14540), .A(n14539), .ZN(n14547) );
  NAND2_X1 U16479 ( .A1(n14762), .A2(n15351), .ZN(n14545) );
  NAND2_X1 U16480 ( .A1(n14764), .A2(n14827), .ZN(n14543) );
  NAND2_X1 U16481 ( .A1(n14720), .A2(n14825), .ZN(n14542) );
  NAND2_X1 U16482 ( .A1(n14543), .A2(n14542), .ZN(n14813) );
  AOI22_X1 U16483 ( .A1(n15348), .A2(n14813), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14544) );
  OAI211_X1 U16484 ( .C1(n15369), .C2(n14815), .A(n14545), .B(n14544), .ZN(
        n14546) );
  AOI21_X1 U16485 ( .B1(n14547), .B2(n15365), .A(n14546), .ZN(n14548) );
  INV_X1 U16486 ( .A(n14548), .ZN(P1_U3240) );
  MUX2_X1 U16487 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14731), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16488 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14549), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16489 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14789), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16490 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14764), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16491 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14828), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16492 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14720), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16493 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14826), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16494 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14717), .S(P1_U4016), .Z(
        P1_U3583) );
  INV_X1 U16495 ( .A(n14714), .ZN(n14755) );
  MUX2_X1 U16496 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14755), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16497 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14712), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16498 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14750), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16499 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14709), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16500 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14705), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16501 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14703), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16502 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14699), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16503 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14550), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16504 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14551), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16505 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14552), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16506 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14553), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16507 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14554), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16508 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14555), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16509 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14556), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16510 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14557), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16511 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14558), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16512 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14559), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16513 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14560), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16514 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14561), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16515 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n10536), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16516 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14562), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16517 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14563), .S(P1_U4016), .Z(
        P1_U3560) );
  NAND2_X1 U16518 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14573) );
  OAI211_X1 U16519 ( .C1(n10898), .C2(n14564), .A(n15462), .B(n14586), .ZN(
        n14571) );
  AOI22_X1 U16520 ( .A1(n15450), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14570) );
  NAND2_X1 U16521 ( .A1(n15460), .A2(n7504), .ZN(n14569) );
  NAND2_X1 U16522 ( .A1(n14566), .A2(n14565), .ZN(n14567) );
  NAND3_X1 U16523 ( .A1(n15469), .A2(n14581), .A3(n14567), .ZN(n14568) );
  NAND4_X1 U16524 ( .A1(n14571), .A2(n14570), .A3(n14569), .A4(n14568), .ZN(
        P1_U3244) );
  MUX2_X1 U16525 ( .A(n14573), .B(n14572), .S(n6678), .Z(n14575) );
  NOR2_X1 U16526 ( .A1(n6678), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n14574) );
  OR2_X1 U16527 ( .A1(n14574), .A2(n10501), .ZN(n15444) );
  NAND2_X1 U16528 ( .A1(n15444), .A2(n7693), .ZN(n15448) );
  OAI211_X1 U16529 ( .C1(n14575), .C2(n10501), .A(P1_U4016), .B(n15448), .ZN(
        n15472) );
  OAI22_X1 U16530 ( .A1(n15489), .A2(n9208), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14576), .ZN(n14577) );
  AOI21_X1 U16531 ( .B1(n14578), .B2(n15460), .A(n14577), .ZN(n14591) );
  INV_X1 U16532 ( .A(n14579), .ZN(n14601) );
  NAND3_X1 U16533 ( .A1(n14582), .A2(n14581), .A3(n14580), .ZN(n14583) );
  NAND3_X1 U16534 ( .A1(n15469), .A2(n14601), .A3(n14583), .ZN(n14590) );
  MUX2_X1 U16535 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n7674), .S(n14584), .Z(
        n14587) );
  NAND3_X1 U16536 ( .A1(n14587), .A2(n14586), .A3(n14585), .ZN(n14588) );
  NAND3_X1 U16537 ( .A1(n15462), .A2(n14593), .A3(n14588), .ZN(n14589) );
  NAND4_X1 U16538 ( .A1(n15472), .A2(n14591), .A3(n14590), .A4(n14589), .ZN(
        P1_U3245) );
  MUX2_X1 U16539 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10901), .S(n14598), .Z(
        n14594) );
  NAND3_X1 U16540 ( .A1(n14594), .A2(n14593), .A3(n14592), .ZN(n14595) );
  NAND3_X1 U16541 ( .A1(n15462), .A2(n15456), .A3(n14595), .ZN(n14606) );
  AOI22_X1 U16542 ( .A1(n15450), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(P1_U3086), .ZN(n14605) );
  NAND2_X1 U16543 ( .A1(n15460), .A2(n14596), .ZN(n14604) );
  INV_X1 U16544 ( .A(n14597), .ZN(n14600) );
  INV_X1 U16545 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n15553) );
  MUX2_X1 U16546 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n15553), .S(n14598), .Z(
        n14599) );
  NAND3_X1 U16547 ( .A1(n14601), .A2(n14600), .A3(n14599), .ZN(n14602) );
  NAND3_X1 U16548 ( .A1(n15469), .A2(n15466), .A3(n14602), .ZN(n14603) );
  NAND4_X1 U16549 ( .A1(n14606), .A2(n14605), .A3(n14604), .A4(n14603), .ZN(
        P1_U3246) );
  NAND2_X1 U16550 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n14607) );
  OAI21_X1 U16551 ( .B1(n15489), .B2(n14608), .A(n14607), .ZN(n14609) );
  AOI21_X1 U16552 ( .B1(n14610), .B2(n15460), .A(n14609), .ZN(n14622) );
  OAI21_X1 U16553 ( .B1(n14613), .B2(n14612), .A(n14611), .ZN(n14614) );
  NAND2_X1 U16554 ( .A1(n15469), .A2(n14614), .ZN(n14621) );
  INV_X1 U16555 ( .A(n14615), .ZN(n14619) );
  NAND3_X1 U16556 ( .A1(n15458), .A2(n14617), .A3(n14616), .ZN(n14618) );
  NAND3_X1 U16557 ( .A1(n15462), .A2(n14619), .A3(n14618), .ZN(n14620) );
  NAND3_X1 U16558 ( .A1(n14622), .A2(n14621), .A3(n14620), .ZN(P1_U3248) );
  NOR2_X1 U16559 ( .A1(n15485), .A2(n14623), .ZN(n14624) );
  AOI211_X1 U16560 ( .C1(n15450), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n14625), .B(
        n14624), .ZN(n14641) );
  INV_X1 U16561 ( .A(n14626), .ZN(n14629) );
  MUX2_X1 U16562 ( .A(n10924), .B(P1_REG1_REG_7__SCAN_IN), .S(n14627), .Z(
        n14628) );
  NAND2_X1 U16563 ( .A1(n14629), .A2(n14628), .ZN(n14631) );
  OAI211_X1 U16564 ( .C1(n14632), .C2(n14631), .A(n15469), .B(n14630), .ZN(
        n14640) );
  INV_X1 U16565 ( .A(n14633), .ZN(n14638) );
  NAND3_X1 U16566 ( .A1(n14636), .A2(n14635), .A3(n14634), .ZN(n14637) );
  NAND3_X1 U16567 ( .A1(n15462), .A2(n14638), .A3(n14637), .ZN(n14639) );
  NAND3_X1 U16568 ( .A1(n14641), .A2(n14640), .A3(n14639), .ZN(P1_U3250) );
  OAI21_X1 U16569 ( .B1(n14644), .B2(n14643), .A(n14642), .ZN(n14645) );
  NAND2_X1 U16570 ( .A1(n14645), .A2(n15469), .ZN(n14656) );
  INV_X1 U16571 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14646) );
  NAND2_X1 U16572 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n15352)
         );
  OAI21_X1 U16573 ( .B1(n15489), .B2(n14646), .A(n15352), .ZN(n14647) );
  AOI21_X1 U16574 ( .B1(n15460), .B2(n14648), .A(n14647), .ZN(n14655) );
  OR3_X1 U16575 ( .A1(n14651), .A2(n14650), .A3(n14649), .ZN(n14652) );
  NAND3_X1 U16576 ( .A1(n14653), .A2(n15462), .A3(n14652), .ZN(n14654) );
  NAND3_X1 U16577 ( .A1(n14656), .A2(n14655), .A3(n14654), .ZN(P1_U3254) );
  NAND2_X1 U16578 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n15330)
         );
  OAI211_X1 U16579 ( .C1(n14659), .C2(n14658), .A(n15469), .B(n14657), .ZN(
        n14660) );
  AND2_X1 U16580 ( .A1(n15330), .A2(n14660), .ZN(n14667) );
  AOI22_X1 U16581 ( .A1(n15460), .A2(n14661), .B1(n15450), .B2(
        P1_ADDR_REG_16__SCAN_IN), .ZN(n14666) );
  OAI211_X1 U16582 ( .C1(n14664), .C2(n14663), .A(n15462), .B(n14662), .ZN(
        n14665) );
  NAND3_X1 U16583 ( .A1(n14667), .A2(n14666), .A3(n14665), .ZN(P1_U3259) );
  NAND2_X1 U16584 ( .A1(n14674), .A2(n14668), .ZN(n14669) );
  NAND2_X1 U16585 ( .A1(n14670), .A2(n14669), .ZN(n14672) );
  INV_X1 U16586 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14671) );
  XNOR2_X1 U16587 ( .A(n14672), .B(n14671), .ZN(n14681) );
  INV_X1 U16588 ( .A(n14681), .ZN(n14679) );
  NAND2_X1 U16589 ( .A1(n14674), .A2(n14673), .ZN(n14675) );
  NAND2_X1 U16590 ( .A1(n14676), .A2(n14675), .ZN(n14677) );
  XOR2_X1 U16591 ( .A(n14677), .B(P1_REG2_REG_19__SCAN_IN), .Z(n14680) );
  NOR2_X1 U16592 ( .A1(n14680), .A2(n15481), .ZN(n14678) );
  AOI211_X1 U16593 ( .C1(n15469), .C2(n14679), .A(n15460), .B(n14678), .ZN(
        n14683) );
  AOI22_X1 U16594 ( .A1(n14681), .A2(n15469), .B1(n15462), .B2(n14680), .ZN(
        n14682) );
  MUX2_X1 U16595 ( .A(n14683), .B(n14682), .S(n14973), .Z(n14686) );
  INV_X1 U16596 ( .A(n14684), .ZN(n14685) );
  OAI211_X1 U16597 ( .C1(n7835), .C2(n15489), .A(n14686), .B(n14685), .ZN(
        P1_U3262) );
  INV_X1 U16598 ( .A(n14762), .ZN(n15008) );
  NAND2_X1 U16599 ( .A1(n14944), .A2(n14952), .ZN(n14941) );
  INV_X1 U16600 ( .A(n15024), .ZN(n14868) );
  NOR2_X2 U16601 ( .A1(n7758), .A2(n15014), .ZN(n14832) );
  NAND2_X1 U16602 ( .A1(n14985), .A2(n14727), .ZN(n14693) );
  XNOR2_X1 U16603 ( .A(n14982), .B(n14693), .ZN(n14980) );
  NAND2_X1 U16604 ( .A1(n14980), .A2(n14946), .ZN(n14692) );
  NOR2_X1 U16605 ( .A1(n6678), .A2(n14688), .ZN(n14689) );
  NOR2_X1 U16606 ( .A1(n14967), .A2(n14689), .ZN(n14730) );
  NAND2_X1 U16607 ( .A1(n14690), .A2(n14730), .ZN(n14983) );
  NOR2_X1 U16608 ( .A1(n15509), .A2(n14983), .ZN(n14694) );
  AOI21_X1 U16609 ( .B1(n15495), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14694), 
        .ZN(n14691) );
  OAI211_X1 U16610 ( .C1(n14982), .C2(n15497), .A(n14692), .B(n14691), .ZN(
        P1_U3263) );
  OAI211_X1 U16611 ( .C1(n14985), .C2(n14727), .A(n15503), .B(n14693), .ZN(
        n14984) );
  NAND2_X1 U16612 ( .A1(n15495), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n14696) );
  INV_X1 U16613 ( .A(n14694), .ZN(n14695) );
  OAI211_X1 U16614 ( .C1(n14985), .C2(n15497), .A(n14696), .B(n14695), .ZN(
        n14697) );
  INV_X1 U16615 ( .A(n14697), .ZN(n14698) );
  OAI21_X1 U16616 ( .B1(n14984), .B2(n14873), .A(n14698), .ZN(P1_U3264) );
  OR2_X1 U16617 ( .A1(n14700), .A2(n14699), .ZN(n14701) );
  INV_X1 U16618 ( .A(n14961), .ZN(n14965) );
  OR2_X1 U16619 ( .A1(n15371), .A2(n14703), .ZN(n14704) );
  NAND2_X1 U16620 ( .A1(n15064), .A2(n14705), .ZN(n14706) );
  NAND2_X2 U16621 ( .A1(n14914), .A2(n14913), .ZN(n14912) );
  OR2_X1 U16622 ( .A1(n14911), .A2(n14710), .ZN(n14711) );
  OR2_X1 U16623 ( .A1(n15041), .A2(n14712), .ZN(n14713) );
  INV_X1 U16624 ( .A(n14877), .ZN(n14878) );
  NAND2_X1 U16625 ( .A1(n14884), .A2(n14714), .ZN(n14715) );
  NAND2_X2 U16626 ( .A1(n14716), .A2(n7705), .ZN(n15026) );
  NAND2_X1 U16627 ( .A1(n15024), .A2(n14717), .ZN(n14718) );
  OR2_X1 U16628 ( .A1(n14859), .A2(n14826), .ZN(n14719) );
  NAND2_X1 U16629 ( .A1(n15014), .A2(n14720), .ZN(n14721) );
  NAND2_X1 U16630 ( .A1(n14762), .A2(n14828), .ZN(n14722) );
  INV_X1 U16631 ( .A(n14764), .ZN(n14723) );
  NAND2_X1 U16632 ( .A1(n14781), .A2(n14724), .ZN(n14726) );
  INV_X1 U16633 ( .A(n14773), .ZN(n14728) );
  AOI211_X1 U16634 ( .C1(n14729), .C2(n14728), .A(n15061), .B(n14727), .ZN(
        n14986) );
  NAND2_X1 U16635 ( .A1(n14789), .A2(n14825), .ZN(n14988) );
  NAND2_X1 U16636 ( .A1(n14731), .A2(n14730), .ZN(n14987) );
  NOR2_X1 U16637 ( .A1(n14987), .A2(n14732), .ZN(n14736) );
  INV_X1 U16638 ( .A(n14733), .ZN(n14734) );
  AOI22_X1 U16639 ( .A1(n14736), .A2(n14735), .B1(n14734), .B2(n15494), .ZN(
        n14737) );
  OAI21_X1 U16640 ( .B1(n15495), .B2(n14988), .A(n14737), .ZN(n14738) );
  AOI21_X1 U16641 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n15495), .A(n14738), 
        .ZN(n14739) );
  OAI21_X1 U16642 ( .B1(n14989), .B2(n15497), .A(n14739), .ZN(n14740) );
  AOI21_X1 U16643 ( .B1(n14986), .B2(n15505), .A(n14740), .ZN(n14768) );
  INV_X1 U16644 ( .A(n14745), .ZN(n14936) );
  NAND2_X1 U16645 ( .A1(n14932), .A2(n14936), .ZN(n14748) );
  NAND2_X1 U16646 ( .A1(n14944), .A2(n14746), .ZN(n14747) );
  NAND2_X1 U16647 ( .A1(n14911), .A2(n14750), .ZN(n14751) );
  NAND2_X1 U16648 ( .A1(n14903), .A2(n14751), .ZN(n14892) );
  NAND2_X1 U16649 ( .A1(n14892), .A2(n14891), .ZN(n14754) );
  OR2_X1 U16650 ( .A1(n15041), .A2(n14752), .ZN(n14753) );
  OR2_X1 U16651 ( .A1(n14884), .A2(n14755), .ZN(n14756) );
  NAND2_X1 U16652 ( .A1(n15024), .A2(n14845), .ZN(n14847) );
  INV_X1 U16653 ( .A(n14848), .ZN(n14757) );
  NAND2_X1 U16654 ( .A1(n14758), .A2(n14757), .ZN(n14850) );
  NAND2_X1 U16655 ( .A1(n14850), .A2(n14759), .ZN(n14824) );
  INV_X1 U16656 ( .A(n14838), .ZN(n14823) );
  NAND2_X1 U16657 ( .A1(n14824), .A2(n14823), .ZN(n14822) );
  NAND2_X1 U16658 ( .A1(n15014), .A2(n14846), .ZN(n14760) );
  NAND2_X1 U16659 ( .A1(n14822), .A2(n14760), .ZN(n14811) );
  INV_X1 U16660 ( .A(n14807), .ZN(n14810) );
  NAND2_X1 U16661 ( .A1(n14811), .A2(n14810), .ZN(n14809) );
  NAND2_X1 U16662 ( .A1(n14762), .A2(n14761), .ZN(n14763) );
  NAND2_X1 U16663 ( .A1(n14809), .A2(n14763), .ZN(n14786) );
  INV_X1 U16664 ( .A(n14779), .ZN(n14995) );
  XNOR2_X1 U16665 ( .A(n14766), .B(n14765), .ZN(n14991) );
  NAND2_X1 U16666 ( .A1(n14991), .A2(n14958), .ZN(n14767) );
  OAI211_X1 U16667 ( .C1(n14992), .C2(n14960), .A(n14768), .B(n14767), .ZN(
        P1_U3356) );
  OAI21_X1 U16668 ( .B1(n14771), .B2(n14770), .A(n14769), .ZN(n14997) );
  AND2_X1 U16669 ( .A1(n14779), .A2(n14797), .ZN(n14772) );
  OR3_X1 U16670 ( .A1(n14773), .A2(n14772), .A3(n15061), .ZN(n14994) );
  INV_X1 U16671 ( .A(n14774), .ZN(n14993) );
  NAND2_X1 U16672 ( .A1(n15495), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n14777) );
  OR2_X1 U16673 ( .A1(n14975), .A2(n14775), .ZN(n14776) );
  OAI211_X1 U16674 ( .C1(n15509), .C2(n14993), .A(n14777), .B(n14776), .ZN(
        n14778) );
  AOI21_X1 U16675 ( .B1(n14779), .B2(n14963), .A(n14778), .ZN(n14780) );
  OAI21_X1 U16676 ( .B1(n14994), .B2(n14873), .A(n14780), .ZN(n14784) );
  OAI21_X1 U16677 ( .B1(n14782), .B2(n7714), .A(n14781), .ZN(n14999) );
  NOR2_X1 U16678 ( .A1(n14999), .A2(n14960), .ZN(n14783) );
  INV_X1 U16679 ( .A(n14785), .ZN(P1_U3265) );
  OR2_X1 U16680 ( .A1(n14786), .A2(n14794), .ZN(n14787) );
  NAND2_X1 U16681 ( .A1(n14788), .A2(n14787), .ZN(n14793) );
  NAND2_X1 U16682 ( .A1(n14828), .A2(n14825), .ZN(n14791) );
  NAND2_X1 U16683 ( .A1(n14789), .A2(n14827), .ZN(n14790) );
  NAND2_X1 U16684 ( .A1(n14791), .A2(n14790), .ZN(n14792) );
  AOI21_X1 U16685 ( .B1(n14793), .B2(n15534), .A(n14792), .ZN(n15005) );
  OR2_X1 U16686 ( .A1(n14796), .A2(n14795), .ZN(n15003) );
  AOI21_X1 U16687 ( .B1(n14802), .B2(n14812), .A(n15061), .ZN(n14798) );
  NAND2_X1 U16688 ( .A1(n14798), .A2(n14797), .ZN(n15000) );
  OAI22_X1 U16689 ( .A1(n14922), .A2(n14800), .B1(n14799), .B2(n14975), .ZN(
        n14801) );
  AOI21_X1 U16690 ( .B1(n14802), .B2(n14963), .A(n14801), .ZN(n14803) );
  OAI21_X1 U16691 ( .B1(n15000), .B2(n14873), .A(n14803), .ZN(n14804) );
  AOI21_X1 U16692 ( .B1(n15003), .B2(n15506), .A(n14804), .ZN(n14805) );
  OAI21_X1 U16693 ( .B1(n15005), .B2(n15509), .A(n14805), .ZN(P1_U3266) );
  OAI21_X1 U16694 ( .B1(n14808), .B2(n14807), .A(n14806), .ZN(n15012) );
  OAI21_X1 U16695 ( .B1(n14811), .B2(n14810), .A(n14809), .ZN(n15010) );
  NAND2_X1 U16696 ( .A1(n15010), .A2(n14958), .ZN(n14821) );
  OAI211_X1 U16697 ( .C1(n15008), .C2(n14832), .A(n15503), .B(n14812), .ZN(
        n15007) );
  INV_X1 U16698 ( .A(n14813), .ZN(n15006) );
  OAI21_X1 U16699 ( .B1(n15007), .B2(n14814), .A(n15006), .ZN(n14819) );
  NOR2_X1 U16700 ( .A1(n15008), .A2(n15497), .ZN(n14818) );
  OAI22_X1 U16701 ( .A1(n14922), .A2(n14816), .B1(n14815), .B2(n14975), .ZN(
        n14817) );
  AOI211_X1 U16702 ( .C1(n14819), .C2(n14922), .A(n14818), .B(n14817), .ZN(
        n14820) );
  OAI211_X1 U16703 ( .C1(n15012), .C2(n14960), .A(n14821), .B(n14820), .ZN(
        P1_U3267) );
  OAI21_X1 U16704 ( .B1(n14824), .B2(n14823), .A(n14822), .ZN(n14829) );
  AOI222_X1 U16705 ( .A1(n15534), .A2(n14829), .B1(n14828), .B2(n14827), .C1(
        n14826), .C2(n14825), .ZN(n15018) );
  NAND2_X1 U16706 ( .A1(n15014), .A2(n7758), .ZN(n14830) );
  NAND2_X1 U16707 ( .A1(n14830), .A2(n15503), .ZN(n14831) );
  NOR2_X1 U16708 ( .A1(n14832), .A2(n14831), .ZN(n15013) );
  OAI22_X1 U16709 ( .A1(n14922), .A2(n14834), .B1(n14833), .B2(n14975), .ZN(
        n14837) );
  INV_X1 U16710 ( .A(n15014), .ZN(n14835) );
  NOR2_X1 U16711 ( .A1(n14835), .A2(n15497), .ZN(n14836) );
  AOI211_X1 U16712 ( .C1(n15013), .C2(n15505), .A(n14837), .B(n14836), .ZN(
        n14842) );
  OR2_X1 U16713 ( .A1(n14839), .A2(n14838), .ZN(n15015) );
  NAND3_X1 U16714 ( .A1(n15015), .A2(n15506), .A3(n14840), .ZN(n14841) );
  OAI211_X1 U16715 ( .C1(n15018), .C2(n15495), .A(n14842), .B(n14841), .ZN(
        P1_U3268) );
  OAI21_X1 U16716 ( .B1(n14844), .B2(n14848), .A(n14843), .ZN(n14853) );
  OAI22_X1 U16717 ( .A1(n14846), .A2(n14967), .B1(n14845), .B2(n14966), .ZN(
        n14852) );
  NAND3_X1 U16718 ( .A1(n14861), .A2(n14848), .A3(n14847), .ZN(n14849) );
  AOI21_X1 U16719 ( .B1(n14850), .B2(n14849), .A(n15393), .ZN(n14851) );
  AOI211_X1 U16720 ( .C1(n15549), .C2(n14853), .A(n14852), .B(n14851), .ZN(
        n15020) );
  OAI22_X1 U16721 ( .A1(n14922), .A2(n14855), .B1(n14854), .B2(n14975), .ZN(
        n14858) );
  INV_X1 U16722 ( .A(n14859), .ZN(n15021) );
  INV_X1 U16723 ( .A(n14863), .ZN(n14856) );
  OAI211_X1 U16724 ( .C1(n15021), .C2(n14856), .A(n7758), .B(n15503), .ZN(
        n15019) );
  NOR2_X1 U16725 ( .A1(n15019), .A2(n14873), .ZN(n14857) );
  AOI211_X1 U16726 ( .C1(n14963), .C2(n14859), .A(n14858), .B(n14857), .ZN(
        n14860) );
  OAI21_X1 U16727 ( .B1(n15020), .B2(n15509), .A(n14860), .ZN(P1_U3269) );
  OAI21_X1 U16728 ( .B1(n14862), .B2(n14864), .A(n14861), .ZN(n15022) );
  OAI211_X1 U16729 ( .C1(n6708), .C2(n14868), .A(n15503), .B(n14863), .ZN(
        n15027) );
  NAND2_X1 U16730 ( .A1(n14865), .A2(n14864), .ZN(n15025) );
  NAND3_X1 U16731 ( .A1(n15026), .A2(n15025), .A3(n15506), .ZN(n14872) );
  INV_X1 U16732 ( .A(n15023), .ZN(n14867) );
  OAI22_X1 U16733 ( .A1(n15495), .A2(n14867), .B1(n14866), .B2(n14975), .ZN(
        n14870) );
  NOR2_X1 U16734 ( .A1(n14868), .A2(n15497), .ZN(n14869) );
  AOI211_X1 U16735 ( .C1(n15495), .C2(P1_REG2_REG_23__SCAN_IN), .A(n14870), 
        .B(n14869), .ZN(n14871) );
  OAI211_X1 U16736 ( .C1(n15027), .C2(n14873), .A(n14872), .B(n14871), .ZN(
        n14874) );
  AOI21_X1 U16737 ( .B1(n15022), .B2(n14958), .A(n14874), .ZN(n14875) );
  INV_X1 U16738 ( .A(n14875), .ZN(P1_U3270) );
  XNOR2_X1 U16739 ( .A(n14876), .B(n14877), .ZN(n15037) );
  XNOR2_X1 U16740 ( .A(n14879), .B(n14878), .ZN(n15034) );
  NAND2_X1 U16741 ( .A1(n15034), .A2(n14958), .ZN(n14887) );
  AOI211_X1 U16742 ( .C1(n15033), .C2(n14893), .A(n15061), .B(n6708), .ZN(
        n15031) );
  INV_X1 U16743 ( .A(n15032), .ZN(n14881) );
  OAI22_X1 U16744 ( .A1(n14881), .A2(n15495), .B1(n14880), .B2(n14975), .ZN(
        n14882) );
  AOI21_X1 U16745 ( .B1(P1_REG2_REG_22__SCAN_IN), .B2(n15495), .A(n14882), 
        .ZN(n14883) );
  OAI21_X1 U16746 ( .B1(n14884), .B2(n15497), .A(n14883), .ZN(n14885) );
  AOI21_X1 U16747 ( .B1(n15031), .B2(n15505), .A(n14885), .ZN(n14886) );
  OAI211_X1 U16748 ( .C1(n15037), .C2(n14960), .A(n14887), .B(n14886), .ZN(
        P1_U3271) );
  INV_X1 U16749 ( .A(n14888), .ZN(n14889) );
  AOI21_X1 U16750 ( .B1(n14891), .B2(n14890), .A(n14889), .ZN(n15044) );
  XOR2_X1 U16751 ( .A(n14892), .B(n14891), .Z(n15038) );
  NAND2_X1 U16752 ( .A1(n15038), .A2(n14958), .ZN(n14901) );
  INV_X1 U16753 ( .A(n14893), .ZN(n14894) );
  AOI211_X1 U16754 ( .C1(n15041), .C2(n14906), .A(n15061), .B(n14894), .ZN(
        n15039) );
  INV_X1 U16755 ( .A(n15041), .ZN(n14898) );
  AOI22_X1 U16756 ( .A1(n15040), .A2(n14922), .B1(n14895), .B2(n15494), .ZN(
        n14897) );
  NAND2_X1 U16757 ( .A1(n15495), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n14896) );
  OAI211_X1 U16758 ( .C1(n14898), .C2(n15497), .A(n14897), .B(n14896), .ZN(
        n14899) );
  AOI21_X1 U16759 ( .B1(n15039), .B2(n15505), .A(n14899), .ZN(n14900) );
  OAI211_X1 U16760 ( .C1(n15044), .C2(n14960), .A(n14901), .B(n14900), .ZN(
        P1_U3272) );
  AOI21_X1 U16761 ( .B1(n6816), .B2(n14913), .A(n15393), .ZN(n14904) );
  AOI21_X1 U16762 ( .B1(n14904), .B2(n14903), .A(n14902), .ZN(n15048) );
  INV_X1 U16763 ( .A(n14905), .ZN(n14920) );
  INV_X1 U16764 ( .A(n14906), .ZN(n14907) );
  AOI211_X1 U16765 ( .C1(n15046), .C2(n14920), .A(n15061), .B(n14907), .ZN(
        n15045) );
  INV_X1 U16766 ( .A(n14908), .ZN(n14909) );
  AOI22_X1 U16767 ( .A1(n15495), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14909), 
        .B2(n15494), .ZN(n14910) );
  OAI21_X1 U16768 ( .B1(n14911), .B2(n15497), .A(n14910), .ZN(n14916) );
  OAI21_X1 U16769 ( .B1(n14914), .B2(n14913), .A(n14912), .ZN(n15049) );
  NOR2_X1 U16770 ( .A1(n15049), .A2(n14960), .ZN(n14915) );
  AOI211_X1 U16771 ( .C1(n15045), .C2(n15505), .A(n14916), .B(n14915), .ZN(
        n14917) );
  OAI21_X1 U16772 ( .B1(n15509), .B2(n15048), .A(n14917), .ZN(P1_U3273) );
  XNOR2_X1 U16773 ( .A(n14919), .B(n14918), .ZN(n15056) );
  AOI211_X1 U16774 ( .C1(n15052), .C2(n14941), .A(n15061), .B(n14905), .ZN(
        n15050) );
  NAND2_X1 U16775 ( .A1(n15495), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n14925) );
  NOR2_X1 U16776 ( .A1(n14975), .A2(n14921), .ZN(n14923) );
  OAI21_X1 U16777 ( .B1(n15051), .B2(n14923), .A(n14922), .ZN(n14924) );
  OAI211_X1 U16778 ( .C1(n14926), .C2(n15497), .A(n14925), .B(n14924), .ZN(
        n14927) );
  AOI21_X1 U16779 ( .B1(n15050), .B2(n15505), .A(n14927), .ZN(n14931) );
  XNOR2_X1 U16780 ( .A(n14929), .B(n14928), .ZN(n15053) );
  NAND2_X1 U16781 ( .A1(n15053), .A2(n14958), .ZN(n14930) );
  OAI211_X1 U16782 ( .C1(n15056), .C2(n14960), .A(n14931), .B(n14930), .ZN(
        P1_U3274) );
  INV_X1 U16783 ( .A(n14933), .ZN(n14934) );
  AOI22_X1 U16784 ( .A1(n14932), .A2(n15534), .B1(n14934), .B2(n15549), .ZN(
        n14938) );
  INV_X1 U16785 ( .A(n14932), .ZN(n14935) );
  AOI22_X1 U16786 ( .A1(n14935), .A2(n15534), .B1(n15549), .B2(n14933), .ZN(
        n14937) );
  MUX2_X1 U16787 ( .A(n14938), .B(n14937), .S(n14936), .Z(n14940) );
  OAI21_X1 U16788 ( .B1(n14944), .B2(n14952), .A(n14941), .ZN(n15060) );
  INV_X1 U16789 ( .A(n15060), .ZN(n14947) );
  AOI22_X1 U16790 ( .A1(n15495), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14942), 
        .B2(n15494), .ZN(n14943) );
  OAI21_X1 U16791 ( .B1(n14944), .B2(n15497), .A(n14943), .ZN(n14945) );
  AOI21_X1 U16792 ( .B1(n14947), .B2(n14946), .A(n14945), .ZN(n14948) );
  OAI21_X1 U16793 ( .B1(n15059), .B2(n15495), .A(n14948), .ZN(P1_U3275) );
  XNOR2_X1 U16794 ( .A(n14949), .B(n14950), .ZN(n15068) );
  XNOR2_X1 U16795 ( .A(n14951), .B(n14950), .ZN(n15065) );
  AOI211_X1 U16796 ( .C1(n15064), .C2(n14970), .A(n15061), .B(n14952), .ZN(
        n15062) );
  NOR2_X1 U16797 ( .A1(n14975), .A2(n14953), .ZN(n14954) );
  AOI211_X1 U16798 ( .C1(n15062), .C2(n14973), .A(n14954), .B(n15063), .ZN(
        n14956) );
  AOI22_X1 U16799 ( .A1(n15064), .A2(n14963), .B1(P1_REG2_REG_17__SCAN_IN), 
        .B2(n15495), .ZN(n14955) );
  OAI21_X1 U16800 ( .B1(n14956), .B2(n15495), .A(n14955), .ZN(n14957) );
  AOI21_X1 U16801 ( .B1(n14958), .B2(n15065), .A(n14957), .ZN(n14959) );
  OAI21_X1 U16802 ( .B1(n14960), .B2(n15068), .A(n14959), .ZN(P1_U3276) );
  XNOR2_X1 U16803 ( .A(n14962), .B(n14961), .ZN(n15374) );
  AOI22_X1 U16804 ( .A1(n15371), .A2(n14963), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n15495), .ZN(n14978) );
  XNOR2_X1 U16805 ( .A(n14964), .B(n14965), .ZN(n14969) );
  OAI22_X1 U16806 ( .A1(n15325), .A2(n14967), .B1(n15326), .B2(n14966), .ZN(
        n14968) );
  AOI21_X1 U16807 ( .B1(n14969), .B2(n15549), .A(n14968), .ZN(n15373) );
  INV_X1 U16808 ( .A(n14970), .ZN(n14971) );
  AOI211_X1 U16809 ( .C1(n15371), .C2(n14972), .A(n15061), .B(n14971), .ZN(
        n15370) );
  NAND2_X1 U16810 ( .A1(n15370), .A2(n14973), .ZN(n14974) );
  OAI211_X1 U16811 ( .C1(n14975), .C2(n15332), .A(n15373), .B(n14974), .ZN(
        n14976) );
  NAND2_X1 U16812 ( .A1(n14976), .A2(n14922), .ZN(n14977) );
  OAI211_X1 U16813 ( .C1(n15374), .C2(n14979), .A(n14978), .B(n14977), .ZN(
        P1_U3277) );
  NAND2_X1 U16814 ( .A1(n14980), .A2(n15503), .ZN(n14981) );
  OAI211_X1 U16815 ( .C1(n14982), .C2(n15545), .A(n14981), .B(n14983), .ZN(
        n15070) );
  MUX2_X1 U16816 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15070), .S(n15559), .Z(
        P1_U3559) );
  OAI211_X1 U16817 ( .C1(n14985), .C2(n15545), .A(n14984), .B(n14983), .ZN(
        n15071) );
  MUX2_X1 U16818 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15071), .S(n15559), .Z(
        P1_U3558) );
  OAI211_X1 U16819 ( .C1(n14989), .C2(n15545), .A(n14988), .B(n14987), .ZN(
        n14990) );
  MUX2_X1 U16820 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n15072), .S(n15559), .Z(
        P1_U3557) );
  OAI211_X1 U16821 ( .C1(n14995), .C2(n15545), .A(n14994), .B(n14993), .ZN(
        n14996) );
  AOI21_X1 U16822 ( .B1(n14997), .B2(n15534), .A(n14996), .ZN(n14998) );
  OAI21_X1 U16823 ( .B1(n14999), .B2(n15529), .A(n14998), .ZN(n15073) );
  MUX2_X1 U16824 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15073), .S(n15559), .Z(
        P1_U3556) );
  OAI21_X1 U16825 ( .B1(n15001), .B2(n15545), .A(n15000), .ZN(n15002) );
  NAND2_X1 U16826 ( .A1(n15005), .A2(n15004), .ZN(n15074) );
  MUX2_X1 U16827 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15074), .S(n15559), .Z(
        P1_U3555) );
  OAI211_X1 U16828 ( .C1(n15008), .C2(n15545), .A(n15007), .B(n15006), .ZN(
        n15009) );
  AOI21_X1 U16829 ( .B1(n15010), .B2(n15534), .A(n15009), .ZN(n15011) );
  OAI21_X1 U16830 ( .B1(n15529), .B2(n15012), .A(n15011), .ZN(n15075) );
  MUX2_X1 U16831 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15075), .S(n15559), .Z(
        P1_U3554) );
  AOI21_X1 U16832 ( .B1(n15387), .B2(n15014), .A(n15013), .ZN(n15017) );
  NAND3_X1 U16833 ( .A1(n15015), .A2(n15549), .A3(n14840), .ZN(n15016) );
  NAND3_X1 U16834 ( .A1(n15018), .A2(n15017), .A3(n15016), .ZN(n15076) );
  MUX2_X1 U16835 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15076), .S(n15559), .Z(
        P1_U3553) );
  OAI211_X1 U16836 ( .C1(n15021), .C2(n15545), .A(n15020), .B(n15019), .ZN(
        n15077) );
  MUX2_X1 U16837 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15077), .S(n15559), .Z(
        P1_U3552) );
  NAND2_X1 U16838 ( .A1(n15022), .A2(n15534), .ZN(n15030) );
  AOI21_X1 U16839 ( .B1(n15024), .B2(n15387), .A(n15023), .ZN(n15029) );
  NAND3_X1 U16840 ( .A1(n15026), .A2(n15549), .A3(n15025), .ZN(n15028) );
  NAND4_X1 U16841 ( .A1(n15030), .A2(n15029), .A3(n15028), .A4(n15027), .ZN(
        n15078) );
  MUX2_X1 U16842 ( .A(n15078), .B(P1_REG1_REG_23__SCAN_IN), .S(n15557), .Z(
        P1_U3551) );
  AOI211_X1 U16843 ( .C1(n15387), .C2(n15033), .A(n15032), .B(n15031), .ZN(
        n15036) );
  NAND2_X1 U16844 ( .A1(n15034), .A2(n15534), .ZN(n15035) );
  OAI211_X1 U16845 ( .C1(n15037), .C2(n15529), .A(n15036), .B(n15035), .ZN(
        n15079) );
  MUX2_X1 U16846 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15079), .S(n15559), .Z(
        P1_U3550) );
  NAND2_X1 U16847 ( .A1(n15038), .A2(n15534), .ZN(n15043) );
  AOI211_X1 U16848 ( .C1(n15387), .C2(n15041), .A(n15040), .B(n15039), .ZN(
        n15042) );
  OAI211_X1 U16849 ( .C1(n15044), .C2(n15529), .A(n15043), .B(n15042), .ZN(
        n15080) );
  MUX2_X1 U16850 ( .A(n15080), .B(P1_REG1_REG_21__SCAN_IN), .S(n15557), .Z(
        P1_U3549) );
  AOI21_X1 U16851 ( .B1(n15387), .B2(n15046), .A(n15045), .ZN(n15047) );
  OAI211_X1 U16852 ( .C1(n15529), .C2(n15049), .A(n15048), .B(n15047), .ZN(
        n15081) );
  MUX2_X1 U16853 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15081), .S(n15559), .Z(
        P1_U3548) );
  AOI211_X1 U16854 ( .C1(n15387), .C2(n15052), .A(n15051), .B(n15050), .ZN(
        n15055) );
  NAND2_X1 U16855 ( .A1(n15053), .A2(n15534), .ZN(n15054) );
  OAI211_X1 U16856 ( .C1(n15056), .C2(n15529), .A(n15055), .B(n15054), .ZN(
        n15082) );
  MUX2_X1 U16857 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15082), .S(n15559), .Z(
        P1_U3547) );
  NAND2_X1 U16858 ( .A1(n15057), .A2(n15387), .ZN(n15058) );
  OAI211_X1 U16859 ( .C1(n15061), .C2(n15060), .A(n15059), .B(n15058), .ZN(
        n15083) );
  MUX2_X1 U16860 ( .A(n15083), .B(P1_REG1_REG_18__SCAN_IN), .S(n15557), .Z(
        P1_U3546) );
  AOI211_X1 U16861 ( .C1(n15387), .C2(n15064), .A(n15063), .B(n15062), .ZN(
        n15067) );
  NAND2_X1 U16862 ( .A1(n15065), .A2(n15534), .ZN(n15066) );
  OAI211_X1 U16863 ( .C1(n15529), .C2(n15068), .A(n15067), .B(n15066), .ZN(
        n15084) );
  MUX2_X1 U16864 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15084), .S(n15559), .Z(
        P1_U3545) );
  MUX2_X1 U16865 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n15069), .S(n15559), .Z(
        P1_U3528) );
  MUX2_X1 U16866 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15070), .S(n15541), .Z(
        P1_U3527) );
  MUX2_X1 U16867 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15071), .S(n15541), .Z(
        P1_U3526) );
  MUX2_X1 U16868 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n15072), .S(n15541), .Z(
        P1_U3525) );
  MUX2_X1 U16869 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15073), .S(n15541), .Z(
        P1_U3524) );
  MUX2_X1 U16870 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15074), .S(n15541), .Z(
        P1_U3523) );
  MUX2_X1 U16871 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15075), .S(n15541), .Z(
        P1_U3522) );
  MUX2_X1 U16872 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15076), .S(n15541), .Z(
        P1_U3521) );
  MUX2_X1 U16873 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15077), .S(n15541), .Z(
        P1_U3520) );
  MUX2_X1 U16874 ( .A(n15078), .B(P1_REG0_REG_23__SCAN_IN), .S(n15550), .Z(
        P1_U3519) );
  MUX2_X1 U16875 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15079), .S(n15541), .Z(
        P1_U3518) );
  MUX2_X1 U16876 ( .A(n15080), .B(P1_REG0_REG_21__SCAN_IN), .S(n15550), .Z(
        P1_U3517) );
  MUX2_X1 U16877 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15081), .S(n15541), .Z(
        P1_U3516) );
  MUX2_X1 U16878 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15082), .S(n15541), .Z(
        P1_U3515) );
  MUX2_X1 U16879 ( .A(n15083), .B(P1_REG0_REG_18__SCAN_IN), .S(n15550), .Z(
        P1_U3513) );
  MUX2_X1 U16880 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15084), .S(n15541), .Z(
        P1_U3510) );
  NAND3_X1 U16881 ( .A1(n9899), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n15088) );
  OAI22_X1 U16882 ( .A1(n15085), .A2(n15088), .B1(n15087), .B2(n15086), .ZN(
        n15089) );
  AOI21_X1 U16883 ( .B1(n10409), .B2(n15090), .A(n15089), .ZN(n15091) );
  INV_X1 U16884 ( .A(n15091), .ZN(P1_U3324) );
  OAI222_X1 U16885 ( .A1(P1_U3086), .A2(n6678), .B1(n15104), .B2(n15093), .C1(
        n15092), .C2(n15101), .ZN(P1_U3328) );
  OAI222_X1 U16886 ( .A1(n15097), .A2(P1_U3086), .B1(n15104), .B2(n15096), 
        .C1(n15095), .C2(n15101), .ZN(P1_U3329) );
  OAI222_X1 U16887 ( .A1(P1_U3086), .A2(n15100), .B1(n15104), .B2(n15099), 
        .C1(n15098), .C2(n15101), .ZN(P1_U3330) );
  OAI222_X1 U16888 ( .A1(P1_U3086), .A2(n15105), .B1(n15104), .B2(n15103), 
        .C1(n15102), .C2(n15101), .ZN(P1_U3331) );
  MUX2_X1 U16889 ( .A(n15106), .B(n10412), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16890 ( .A(n15107), .ZN(n15108) );
  MUX2_X1 U16891 ( .A(n15108), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U16892 ( .A(n15112), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16893 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15113) );
  OAI21_X1 U16894 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n15113), 
        .ZN(U28) );
  AOI21_X1 U16895 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n15114) );
  OAI21_X1 U16896 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n15114), 
        .ZN(U29) );
  OAI21_X1 U16897 ( .B1(n15117), .B2(n15116), .A(n15115), .ZN(n15118) );
  XNOR2_X1 U16898 ( .A(n15118), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  INV_X1 U16899 ( .A(n15119), .ZN(n15122) );
  AOI22_X1 U16900 ( .A1(n15122), .A2(n15121), .B1(SI_13_), .B2(n15120), .ZN(
        n15123) );
  OAI21_X1 U16901 ( .B1(P3_U3151), .B2(n15124), .A(n15123), .ZN(P3_U3282) );
  AOI21_X1 U16902 ( .B1(n15127), .B2(n15126), .A(n15125), .ZN(SUB_1596_U57) );
  AOI21_X1 U16903 ( .B1(n15130), .B2(n15129), .A(n15128), .ZN(SUB_1596_U55) );
  OAI21_X1 U16904 ( .B1(n15133), .B2(n15132), .A(n15131), .ZN(SUB_1596_U54) );
  OAI222_X1 U16905 ( .A1(n15137), .A2(n15136), .B1(n15137), .B2(n15135), .C1(
        n6730), .C2(n15134), .ZN(SUB_1596_U70) );
  AOI21_X1 U16906 ( .B1(n15140), .B2(n15139), .A(n15138), .ZN(n15141) );
  XOR2_X1 U16907 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n15141), .Z(SUB_1596_U63)
         );
  AOI21_X1 U16908 ( .B1(n15144), .B2(n15143), .A(n15142), .ZN(n15159) );
  OAI22_X1 U16909 ( .A1(n15738), .A2(n15146), .B1(n15737), .B2(n15145), .ZN(
        n15156) );
  AOI21_X1 U16910 ( .B1(n15149), .B2(n15148), .A(n15147), .ZN(n15154) );
  AOI21_X1 U16911 ( .B1(n15152), .B2(n15151), .A(n15150), .ZN(n15153) );
  OAI22_X1 U16912 ( .A1(n15154), .A2(n15744), .B1(n15153), .B2(n15746), .ZN(
        n15155) );
  NOR3_X1 U16913 ( .A1(n15157), .A2(n15156), .A3(n15155), .ZN(n15158) );
  OAI21_X1 U16914 ( .B1(n15159), .B2(n15752), .A(n15158), .ZN(P3_U3197) );
  INV_X1 U16915 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n15165) );
  NAND2_X1 U16916 ( .A1(n15162), .A2(n15818), .ZN(n15163) );
  AOI21_X1 U16917 ( .B1(n15222), .B2(n15163), .A(n15822), .ZN(n15166) );
  AOI21_X1 U16918 ( .B1(n13057), .B2(n15780), .A(n15166), .ZN(n15164) );
  OAI21_X1 U16919 ( .B1(n15165), .B2(n15801), .A(n15164), .ZN(P3_U3202) );
  INV_X1 U16920 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n15169) );
  AOI21_X1 U16921 ( .B1(n15167), .B2(n15780), .A(n15166), .ZN(n15168) );
  OAI21_X1 U16922 ( .B1(n15169), .B2(n15801), .A(n15168), .ZN(P3_U3203) );
  AND2_X1 U16923 ( .A1(n15171), .A2(n15170), .ZN(n15172) );
  XOR2_X1 U16924 ( .A(n15176), .B(n15172), .Z(n15174) );
  AOI222_X1 U16925 ( .A1(n15211), .A2(n15174), .B1(n15199), .B2(n15806), .C1(
        n15173), .C2(n15809), .ZN(n15225) );
  AOI22_X1 U16926 ( .A1(n15822), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15818), 
        .B2(n15175), .ZN(n15180) );
  XNOR2_X1 U16927 ( .A(n15177), .B(n15176), .ZN(n15228) );
  NOR2_X1 U16928 ( .A1(n15178), .A2(n15815), .ZN(n15227) );
  AOI22_X1 U16929 ( .A1(n15228), .A2(n15218), .B1(n15217), .B2(n15227), .ZN(
        n15179) );
  OAI211_X1 U16930 ( .C1(n15822), .C2(n15225), .A(n15180), .B(n15179), .ZN(
        P3_U3219) );
  NAND2_X1 U16931 ( .A1(n15182), .A2(n15181), .ZN(n15197) );
  NAND2_X1 U16932 ( .A1(n15197), .A2(n15183), .ZN(n15185) );
  NAND2_X1 U16933 ( .A1(n15185), .A2(n15184), .ZN(n15186) );
  XOR2_X1 U16934 ( .A(n15193), .B(n15186), .Z(n15188) );
  AOI222_X1 U16935 ( .A1(n15211), .A2(n15188), .B1(n15187), .B2(n15809), .C1(
        n15209), .C2(n15806), .ZN(n15229) );
  OAI22_X1 U16936 ( .A1(n15190), .A2(n15801), .B1(n15782), .B2(n15189), .ZN(
        n15191) );
  INV_X1 U16937 ( .A(n15191), .ZN(n15196) );
  XOR2_X1 U16938 ( .A(n15192), .B(n15193), .Z(n15232) );
  NOR2_X1 U16939 ( .A1(n15194), .A2(n15815), .ZN(n15231) );
  AOI22_X1 U16940 ( .A1(n15232), .A2(n15218), .B1(n15217), .B2(n15231), .ZN(
        n15195) );
  OAI211_X1 U16941 ( .C1(n15822), .C2(n15229), .A(n15196), .B(n15195), .ZN(
        P3_U3220) );
  XNOR2_X1 U16942 ( .A(n15197), .B(n15202), .ZN(n15200) );
  AOI222_X1 U16943 ( .A1(n15211), .A2(n15200), .B1(n15199), .B2(n15809), .C1(
        n15198), .C2(n15806), .ZN(n15233) );
  AOI22_X1 U16944 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n15822), .B1(n15818), 
        .B2(n15201), .ZN(n15206) );
  XNOR2_X1 U16945 ( .A(n15203), .B(n15202), .ZN(n15236) );
  NOR2_X1 U16946 ( .A1(n15204), .A2(n15815), .ZN(n15235) );
  AOI22_X1 U16947 ( .A1(n15236), .A2(n15218), .B1(n15217), .B2(n15235), .ZN(
        n15205) );
  OAI211_X1 U16948 ( .C1(n15822), .C2(n15233), .A(n15206), .B(n15205), .ZN(
        P3_U3221) );
  XNOR2_X1 U16949 ( .A(n15207), .B(n15214), .ZN(n15210) );
  AOI222_X1 U16950 ( .A1(n15211), .A2(n15210), .B1(n15209), .B2(n15809), .C1(
        n15208), .C2(n15806), .ZN(n15237) );
  AOI22_X1 U16951 ( .A1(n15822), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n15818), 
        .B2(n15212), .ZN(n15220) );
  OAI21_X1 U16952 ( .B1(n15215), .B2(n15214), .A(n15213), .ZN(n15240) );
  NOR2_X1 U16953 ( .A1(n15216), .A2(n15815), .ZN(n15239) );
  AOI22_X1 U16954 ( .A1(n15240), .A2(n15218), .B1(n15217), .B2(n15239), .ZN(
        n15219) );
  OAI211_X1 U16955 ( .C1(n15822), .C2(n15237), .A(n15220), .B(n15219), .ZN(
        P3_U3222) );
  INV_X1 U16956 ( .A(n15222), .ZN(n15221) );
  AOI21_X1 U16957 ( .B1(n13057), .B2(n15796), .A(n15221), .ZN(n15243) );
  AOI22_X1 U16958 ( .A1(n15854), .A2(n15243), .B1(n11720), .B2(n15851), .ZN(
        P3_U3490) );
  OAI21_X1 U16959 ( .B1(n15223), .B2(n15815), .A(n15222), .ZN(n15244) );
  OAI22_X1 U16960 ( .A1(n15851), .A2(n15244), .B1(P3_REG1_REG_30__SCAN_IN), 
        .B2(n15854), .ZN(n15224) );
  INV_X1 U16961 ( .A(n15224), .ZN(P3_U3489) );
  INV_X1 U16962 ( .A(n15225), .ZN(n15226) );
  AOI211_X1 U16963 ( .C1(n15241), .C2(n15228), .A(n15227), .B(n15226), .ZN(
        n15247) );
  AOI22_X1 U16964 ( .A1(n15854), .A2(n15247), .B1(n13269), .B2(n15851), .ZN(
        P3_U3473) );
  INV_X1 U16965 ( .A(n15229), .ZN(n15230) );
  AOI211_X1 U16966 ( .C1(n15232), .C2(n15241), .A(n15231), .B(n15230), .ZN(
        n15249) );
  AOI22_X1 U16967 ( .A1(n15854), .A2(n15249), .B1(n8048), .B2(n15851), .ZN(
        P3_U3472) );
  INV_X1 U16968 ( .A(n15233), .ZN(n15234) );
  AOI211_X1 U16969 ( .C1(n15236), .C2(n15241), .A(n15235), .B(n15234), .ZN(
        n15251) );
  AOI22_X1 U16970 ( .A1(n15854), .A2(n15251), .B1(n12413), .B2(n15851), .ZN(
        P3_U3471) );
  INV_X1 U16971 ( .A(n15237), .ZN(n15238) );
  AOI211_X1 U16972 ( .C1(n15241), .C2(n15240), .A(n15239), .B(n15238), .ZN(
        n15253) );
  AOI22_X1 U16973 ( .A1(n15854), .A2(n15253), .B1(n8015), .B2(n15851), .ZN(
        P3_U3470) );
  INV_X1 U16974 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n15242) );
  AOI22_X1 U16975 ( .A1(n15846), .A2(n15243), .B1(n15242), .B2(n15844), .ZN(
        P3_U3458) );
  OAI22_X1 U16976 ( .A1(n15844), .A2(n15244), .B1(P3_REG0_REG_30__SCAN_IN), 
        .B2(n15846), .ZN(n15245) );
  INV_X1 U16977 ( .A(n15245), .ZN(P3_U3457) );
  INV_X1 U16978 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n15246) );
  AOI22_X1 U16979 ( .A1(n15846), .A2(n15247), .B1(n15246), .B2(n15844), .ZN(
        P3_U3432) );
  INV_X1 U16980 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n15248) );
  AOI22_X1 U16981 ( .A1(n15846), .A2(n15249), .B1(n15248), .B2(n15844), .ZN(
        P3_U3429) );
  INV_X1 U16982 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n15250) );
  AOI22_X1 U16983 ( .A1(n15846), .A2(n15251), .B1(n15250), .B2(n15844), .ZN(
        P3_U3426) );
  INV_X1 U16984 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n15252) );
  AOI22_X1 U16985 ( .A1(n15846), .A2(n15253), .B1(n15252), .B2(n15844), .ZN(
        P3_U3423) );
  XNOR2_X1 U16986 ( .A(n15267), .B(n15254), .ZN(n15257) );
  AOI21_X1 U16987 ( .B1(n15257), .B2(n15256), .A(n15255), .ZN(n15282) );
  INV_X1 U16988 ( .A(n15258), .ZN(n15259) );
  AOI222_X1 U16989 ( .A1(n15280), .A2(n15261), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n15678), .C1(n15260), .C2(n15259), .ZN(n15272) );
  AOI211_X1 U16990 ( .C1(n15280), .C2(n15264), .A(n15263), .B(n15262), .ZN(
        n15279) );
  OAI21_X1 U16991 ( .B1(n15267), .B2(n15266), .A(n15265), .ZN(n15284) );
  INV_X1 U16992 ( .A(n15284), .ZN(n15268) );
  AOI22_X1 U16993 ( .A1(n15279), .A2(n15270), .B1(n15269), .B2(n15268), .ZN(
        n15271) );
  OAI211_X1 U16994 ( .C1(n15678), .C2(n15282), .A(n15272), .B(n15271), .ZN(
        P2_U3251) );
  OAI21_X1 U16995 ( .B1(n15274), .B2(n15718), .A(n15273), .ZN(n15276) );
  AOI211_X1 U16996 ( .C1(n15722), .C2(n15277), .A(n15276), .B(n15275), .ZN(
        n15297) );
  INV_X1 U16997 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n15278) );
  AOI22_X1 U16998 ( .A1(n15731), .A2(n15297), .B1(n15278), .B2(n15729), .ZN(
        P2_U3514) );
  AOI21_X1 U16999 ( .B1(n15281), .B2(n15280), .A(n15279), .ZN(n15283) );
  OAI211_X1 U17000 ( .C1(n15285), .C2(n15284), .A(n15283), .B(n15282), .ZN(
        n15286) );
  INV_X1 U17001 ( .A(n15286), .ZN(n15299) );
  AOI22_X1 U17002 ( .A1(n15731), .A2(n15299), .B1(n15287), .B2(n15729), .ZN(
        P2_U3513) );
  INV_X1 U17003 ( .A(n15710), .ZN(n15692) );
  OAI21_X1 U17004 ( .B1(n15289), .B2(n15718), .A(n15288), .ZN(n15293) );
  OAI21_X1 U17005 ( .B1(n15291), .B2(n15711), .A(n15290), .ZN(n15292) );
  AOI211_X1 U17006 ( .C1(n15692), .C2(n15294), .A(n15293), .B(n15292), .ZN(
        n15301) );
  AOI22_X1 U17007 ( .A1(n15731), .A2(n15301), .B1(n15295), .B2(n15729), .ZN(
        P2_U3511) );
  INV_X1 U17008 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n15296) );
  AOI22_X1 U17009 ( .A1(n15724), .A2(n15297), .B1(n15296), .B2(n9771), .ZN(
        P2_U3475) );
  INV_X1 U17010 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n15298) );
  AOI22_X1 U17011 ( .A1(n15724), .A2(n15299), .B1(n15298), .B2(n9771), .ZN(
        P2_U3472) );
  INV_X1 U17012 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n15300) );
  AOI22_X1 U17013 ( .A1(n15724), .A2(n15301), .B1(n15300), .B2(n9771), .ZN(
        P2_U3466) );
  XNOR2_X1 U17014 ( .A(n15302), .B(n15303), .ZN(n15308) );
  NOR2_X1 U17015 ( .A1(n15304), .A2(n15358), .ZN(n15307) );
  OAI22_X1 U17016 ( .A1(n15305), .A2(n15361), .B1(n15360), .B2(n15326), .ZN(
        n15306) );
  AOI211_X1 U17017 ( .C1(n15308), .C2(n15365), .A(n15307), .B(n15306), .ZN(
        n15310) );
  OAI211_X1 U17018 ( .C1(n15369), .C2(n15311), .A(n15310), .B(n15309), .ZN(
        P1_U3215) );
  OAI22_X1 U17019 ( .A1(n15313), .A2(n15361), .B1(n15360), .B2(n15312), .ZN(
        n15318) );
  XOR2_X1 U17020 ( .A(n15315), .B(n15314), .Z(n15316) );
  NOR2_X1 U17021 ( .A1(n15316), .A2(n15337), .ZN(n15317) );
  AOI211_X1 U17022 ( .C1(n15543), .C2(n15351), .A(n15318), .B(n15317), .ZN(
        n15320) );
  OAI211_X1 U17023 ( .C1(n15369), .C2(n15321), .A(n15320), .B(n15319), .ZN(
        P1_U3217) );
  XNOR2_X1 U17024 ( .A(n15322), .B(n15323), .ZN(n15329) );
  NOR2_X1 U17025 ( .A1(n15324), .A2(n15358), .ZN(n15328) );
  OAI22_X1 U17026 ( .A1(n15326), .A2(n15361), .B1(n15360), .B2(n15325), .ZN(
        n15327) );
  AOI211_X1 U17027 ( .C1(n15329), .C2(n15365), .A(n15328), .B(n15327), .ZN(
        n15331) );
  OAI211_X1 U17028 ( .C1(n15369), .C2(n15332), .A(n15331), .B(n15330), .ZN(
        P1_U3226) );
  OAI22_X1 U17029 ( .A1(n15333), .A2(n15361), .B1(n15360), .B2(n15362), .ZN(
        n15341) );
  AOI21_X1 U17030 ( .B1(n12727), .B2(n15335), .A(n15334), .ZN(n15336) );
  INV_X1 U17031 ( .A(n15336), .ZN(n15339) );
  AOI21_X1 U17032 ( .B1(n15339), .B2(n15338), .A(n15337), .ZN(n15340) );
  AOI211_X1 U17033 ( .C1(n15342), .C2(n15351), .A(n15341), .B(n15340), .ZN(
        n15344) );
  OAI211_X1 U17034 ( .C1(n15369), .C2(n15345), .A(n15344), .B(n15343), .ZN(
        P1_U3234) );
  XNOR2_X1 U17035 ( .A(n15346), .B(n15347), .ZN(n15350) );
  AOI222_X1 U17036 ( .A1(n15351), .A2(n15403), .B1(n15365), .B2(n15350), .C1(
        n15349), .C2(n15348), .ZN(n15353) );
  OAI211_X1 U17037 ( .C1(n15369), .C2(n15354), .A(n15353), .B(n15352), .ZN(
        P1_U3236) );
  OAI21_X1 U17038 ( .B1(n15357), .B2(n15356), .A(n15355), .ZN(n15366) );
  NOR2_X1 U17039 ( .A1(n15378), .A2(n15358), .ZN(n15364) );
  OAI22_X1 U17040 ( .A1(n15362), .A2(n15361), .B1(n15360), .B2(n15359), .ZN(
        n15363) );
  AOI211_X1 U17041 ( .C1(n15366), .C2(n15365), .A(n15364), .B(n15363), .ZN(
        n15367) );
  NAND2_X1 U17042 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n15487)
         );
  OAI211_X1 U17043 ( .C1(n15369), .C2(n15368), .A(n15367), .B(n15487), .ZN(
        P1_U3241) );
  AOI21_X1 U17044 ( .B1(n15387), .B2(n15371), .A(n15370), .ZN(n15372) );
  OAI211_X1 U17045 ( .C1(n15374), .C2(n15393), .A(n15373), .B(n15372), .ZN(
        n15375) );
  INV_X1 U17046 ( .A(n15375), .ZN(n15409) );
  AOI22_X1 U17047 ( .A1(n15559), .A2(n15409), .B1(n12214), .B2(n15557), .ZN(
        P1_U3544) );
  OAI211_X1 U17048 ( .C1(n15378), .C2(n15545), .A(n15377), .B(n15376), .ZN(
        n15382) );
  NOR3_X1 U17049 ( .A1(n15380), .A2(n15379), .A3(n15393), .ZN(n15381) );
  AOI211_X1 U17050 ( .C1(n15549), .C2(n15383), .A(n15382), .B(n15381), .ZN(
        n15411) );
  AOI22_X1 U17051 ( .A1(n15559), .A2(n15411), .B1(n10191), .B2(n15557), .ZN(
        P1_U3543) );
  AOI211_X1 U17052 ( .C1(n15387), .C2(n15386), .A(n15385), .B(n15384), .ZN(
        n15391) );
  NAND3_X1 U17053 ( .A1(n15389), .A2(n15388), .A3(n15549), .ZN(n15390) );
  OAI211_X1 U17054 ( .C1(n15393), .C2(n15392), .A(n15391), .B(n15390), .ZN(
        n15394) );
  INV_X1 U17055 ( .A(n15394), .ZN(n15413) );
  AOI22_X1 U17056 ( .A1(n15559), .A2(n15413), .B1(n10176), .B2(n15557), .ZN(
        P1_U3542) );
  INV_X1 U17057 ( .A(n15395), .ZN(n15402) );
  OAI211_X1 U17058 ( .C1(n15398), .C2(n15545), .A(n15397), .B(n15396), .ZN(
        n15401) );
  INV_X1 U17059 ( .A(n15399), .ZN(n15400) );
  AOI211_X1 U17060 ( .C1(n15402), .C2(n15549), .A(n15401), .B(n15400), .ZN(
        n15415) );
  AOI22_X1 U17061 ( .A1(n15559), .A2(n15415), .B1(n10152), .B2(n15557), .ZN(
        P1_U3541) );
  OAI211_X1 U17062 ( .C1(n7295), .C2(n15545), .A(n15405), .B(n15404), .ZN(
        n15406) );
  AOI21_X1 U17063 ( .B1(n15549), .B2(n15407), .A(n15406), .ZN(n15417) );
  AOI22_X1 U17064 ( .A1(n15559), .A2(n15417), .B1(n10118), .B2(n15557), .ZN(
        P1_U3539) );
  INV_X1 U17065 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n15408) );
  AOI22_X1 U17066 ( .A1(n15541), .A2(n15409), .B1(n15408), .B2(n15550), .ZN(
        P1_U3507) );
  INV_X1 U17067 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n15410) );
  AOI22_X1 U17068 ( .A1(n15541), .A2(n15411), .B1(n15410), .B2(n15550), .ZN(
        P1_U3504) );
  INV_X1 U17069 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n15412) );
  AOI22_X1 U17070 ( .A1(n15541), .A2(n15413), .B1(n15412), .B2(n15550), .ZN(
        P1_U3501) );
  INV_X1 U17071 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n15414) );
  AOI22_X1 U17072 ( .A1(n15541), .A2(n15415), .B1(n15414), .B2(n15550), .ZN(
        P1_U3498) );
  INV_X1 U17073 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n15416) );
  AOI22_X1 U17074 ( .A1(n15541), .A2(n15417), .B1(n15416), .B2(n15550), .ZN(
        P1_U3492) );
  OAI222_X1 U17075 ( .A1(n15422), .A2(n15421), .B1(n15422), .B2(n15420), .C1(
        n15419), .C2(n15418), .ZN(SUB_1596_U69) );
  AOI21_X1 U17076 ( .B1(n15425), .B2(n15424), .A(n15423), .ZN(n15426) );
  XOR2_X1 U17077 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n15426), .Z(SUB_1596_U68)
         );
  OAI21_X1 U17078 ( .B1(n15429), .B2(n15428), .A(n15427), .ZN(n15430) );
  XNOR2_X1 U17079 ( .A(n15430), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  OAI21_X1 U17080 ( .B1(n15433), .B2(n15432), .A(n15431), .ZN(n15434) );
  XNOR2_X1 U17081 ( .A(n15434), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI21_X1 U17082 ( .B1(n15437), .B2(n15436), .A(n15435), .ZN(n15438) );
  XNOR2_X1 U17083 ( .A(n15438), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(SUB_1596_U65)
         );
  OAI21_X1 U17084 ( .B1(n15441), .B2(n15440), .A(n15439), .ZN(n15442) );
  XNOR2_X1 U17085 ( .A(n15442), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  NOR2_X1 U17086 ( .A1(n15443), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n15445) );
  OR2_X1 U17087 ( .A1(n15444), .A2(n15445), .ZN(n15447) );
  INV_X1 U17088 ( .A(n15445), .ZN(n15446) );
  MUX2_X1 U17089 ( .A(n15447), .B(n15446), .S(n7693), .Z(n15449) );
  NAND2_X1 U17090 ( .A1(n15449), .A2(n15448), .ZN(n15452) );
  AOI22_X1 U17091 ( .A1(n15450), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15451) );
  OAI21_X1 U17092 ( .B1(n15453), .B2(n15452), .A(n15451), .ZN(P1_U3243) );
  MUX2_X1 U17093 ( .A(n10904), .B(P1_REG2_REG_4__SCAN_IN), .S(n15459), .Z(
        n15454) );
  NAND3_X1 U17094 ( .A1(n15456), .A2(n15455), .A3(n15454), .ZN(n15457) );
  AND2_X1 U17095 ( .A1(n15458), .A2(n15457), .ZN(n15461) );
  AOI22_X1 U17096 ( .A1(n15462), .A2(n15461), .B1(n15460), .B2(n15459), .ZN(
        n15471) );
  INV_X1 U17097 ( .A(n15463), .ZN(n15468) );
  NAND3_X1 U17098 ( .A1(n15466), .A2(n15465), .A3(n15464), .ZN(n15467) );
  NAND3_X1 U17099 ( .A1(n15469), .A2(n15468), .A3(n15467), .ZN(n15470) );
  AND3_X1 U17100 ( .A1(n15472), .A2(n15471), .A3(n15470), .ZN(n15474) );
  NAND2_X1 U17101 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n15473) );
  OAI211_X1 U17102 ( .C1(n15489), .C2(n15475), .A(n15474), .B(n15473), .ZN(
        P1_U3247) );
  AOI21_X1 U17103 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n15477), .A(n15476), 
        .ZN(n15482) );
  AOI21_X1 U17104 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n15479), .A(n15478), 
        .ZN(n15480) );
  OAI222_X1 U17105 ( .A1(n15485), .A2(n15484), .B1(n15483), .B2(n15482), .C1(
        n15481), .C2(n15480), .ZN(n15486) );
  INV_X1 U17106 ( .A(n15486), .ZN(n15488) );
  OAI211_X1 U17107 ( .C1(n15490), .C2(n15489), .A(n15488), .B(n15487), .ZN(
        P1_U3258) );
  XNOR2_X1 U17108 ( .A(n15491), .B(n15500), .ZN(n15493) );
  AOI21_X1 U17109 ( .B1(n15493), .B2(n15534), .A(n15492), .ZN(n15512) );
  AOI22_X1 U17110 ( .A1(n15495), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n15494), .ZN(n15496) );
  OAI21_X1 U17111 ( .B1(n15497), .B2(n15513), .A(n15496), .ZN(n15498) );
  INV_X1 U17112 ( .A(n15498), .ZN(n15508) );
  XNOR2_X1 U17113 ( .A(n15499), .B(n15500), .ZN(n15515) );
  OAI211_X1 U17114 ( .C1(n7292), .C2(n15513), .A(n15503), .B(n15502), .ZN(
        n15511) );
  INV_X1 U17115 ( .A(n15511), .ZN(n15504) );
  AOI22_X1 U17116 ( .A1(n15506), .A2(n15515), .B1(n15505), .B2(n15504), .ZN(
        n15507) );
  OAI211_X1 U17117 ( .C1(n15509), .C2(n15512), .A(n15508), .B(n15507), .ZN(
        P1_U3291) );
  AND2_X1 U17118 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15510), .ZN(P1_U3294) );
  AND2_X1 U17119 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15510), .ZN(P1_U3295) );
  AND2_X1 U17120 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15510), .ZN(P1_U3296) );
  AND2_X1 U17121 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15510), .ZN(P1_U3297) );
  AND2_X1 U17122 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15510), .ZN(P1_U3298) );
  AND2_X1 U17123 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15510), .ZN(P1_U3299) );
  AND2_X1 U17124 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15510), .ZN(P1_U3300) );
  AND2_X1 U17125 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15510), .ZN(P1_U3301) );
  AND2_X1 U17126 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15510), .ZN(P1_U3302) );
  AND2_X1 U17127 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15510), .ZN(P1_U3303) );
  AND2_X1 U17128 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15510), .ZN(P1_U3304) );
  AND2_X1 U17129 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15510), .ZN(P1_U3305) );
  AND2_X1 U17130 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15510), .ZN(P1_U3306) );
  AND2_X1 U17131 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15510), .ZN(P1_U3307) );
  AND2_X1 U17132 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15510), .ZN(P1_U3308) );
  AND2_X1 U17133 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15510), .ZN(P1_U3309) );
  AND2_X1 U17134 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15510), .ZN(P1_U3310) );
  AND2_X1 U17135 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15510), .ZN(P1_U3311) );
  AND2_X1 U17136 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15510), .ZN(P1_U3312) );
  AND2_X1 U17137 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15510), .ZN(P1_U3313) );
  AND2_X1 U17138 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15510), .ZN(P1_U3314) );
  AND2_X1 U17139 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15510), .ZN(P1_U3315) );
  AND2_X1 U17140 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15510), .ZN(P1_U3316) );
  AND2_X1 U17141 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15510), .ZN(P1_U3317) );
  AND2_X1 U17142 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15510), .ZN(P1_U3318) );
  AND2_X1 U17143 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15510), .ZN(P1_U3319) );
  AND2_X1 U17144 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15510), .ZN(P1_U3320) );
  AND2_X1 U17145 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15510), .ZN(P1_U3321) );
  AND2_X1 U17146 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15510), .ZN(P1_U3322) );
  AND2_X1 U17147 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15510), .ZN(P1_U3323) );
  OAI211_X1 U17148 ( .C1(n15513), .C2(n15545), .A(n15512), .B(n15511), .ZN(
        n15514) );
  AOI21_X1 U17149 ( .B1(n15549), .B2(n15515), .A(n15514), .ZN(n15552) );
  INV_X1 U17150 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n15516) );
  AOI22_X1 U17151 ( .A1(n15541), .A2(n15552), .B1(n15516), .B2(n15550), .ZN(
        P1_U3465) );
  INV_X1 U17152 ( .A(n15517), .ZN(n15524) );
  NOR2_X1 U17153 ( .A1(n15518), .A2(n15545), .ZN(n15519) );
  NOR2_X1 U17154 ( .A1(n15520), .A2(n15519), .ZN(n15523) );
  NAND2_X1 U17155 ( .A1(n15521), .A2(n15549), .ZN(n15522) );
  AND3_X1 U17156 ( .A1(n15524), .A2(n15523), .A3(n15522), .ZN(n15554) );
  AOI22_X1 U17157 ( .A1(n15541), .A2(n15554), .B1(n9969), .B2(n15550), .ZN(
        P1_U3468) );
  INV_X1 U17158 ( .A(n15525), .ZN(n15526) );
  OAI211_X1 U17159 ( .C1(n15528), .C2(n15545), .A(n15527), .B(n15526), .ZN(
        n15532) );
  NOR2_X1 U17160 ( .A1(n15530), .A2(n15529), .ZN(n15531) );
  AOI211_X1 U17161 ( .C1(n15534), .C2(n15533), .A(n15532), .B(n15531), .ZN(
        n15555) );
  AOI22_X1 U17162 ( .A1(n15541), .A2(n15555), .B1(n10001), .B2(n15550), .ZN(
        P1_U3471) );
  AND2_X1 U17163 ( .A1(n15535), .A2(n15549), .ZN(n15539) );
  OAI21_X1 U17164 ( .B1(n15537), .B2(n15545), .A(n15536), .ZN(n15538) );
  NOR3_X1 U17165 ( .A1(n15540), .A2(n15539), .A3(n15538), .ZN(n15556) );
  AOI22_X1 U17166 ( .A1(n15541), .A2(n15556), .B1(n10087), .B2(n15550), .ZN(
        P1_U3486) );
  INV_X1 U17167 ( .A(n15542), .ZN(n15548) );
  OAI21_X1 U17168 ( .B1(n7296), .B2(n15545), .A(n15544), .ZN(n15547) );
  AOI211_X1 U17169 ( .C1(n15549), .C2(n15548), .A(n15547), .B(n15546), .ZN(
        n15558) );
  INV_X1 U17170 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n15551) );
  AOI22_X1 U17171 ( .A1(n15541), .A2(n15558), .B1(n15551), .B2(n15550), .ZN(
        P1_U3489) );
  AOI22_X1 U17172 ( .A1(n15559), .A2(n15552), .B1(n10921), .B2(n15557), .ZN(
        P1_U3530) );
  AOI22_X1 U17173 ( .A1(n15559), .A2(n15554), .B1(n15553), .B2(n15557), .ZN(
        P1_U3531) );
  AOI22_X1 U17174 ( .A1(n15559), .A2(n15555), .B1(n10000), .B2(n15557), .ZN(
        P1_U3532) );
  AOI22_X1 U17175 ( .A1(n15559), .A2(n15556), .B1(n10084), .B2(n15557), .ZN(
        P1_U3537) );
  AOI22_X1 U17176 ( .A1(n15559), .A2(n15558), .B1(n10105), .B2(n15557), .ZN(
        P1_U3538) );
  NOR2_X1 U17177 ( .A1(n15635), .A2(n15560), .ZN(P2_U3087) );
  INV_X1 U17178 ( .A(n15561), .ZN(n15563) );
  OAI21_X1 U17179 ( .B1(n15563), .B2(n15562), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15564) );
  OAI21_X1 U17180 ( .B1(P2_STATE_REG_SCAN_IN), .B2(P2_REG3_REG_1__SCAN_IN), 
        .A(n15564), .ZN(n15576) );
  INV_X1 U17181 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n15725) );
  INV_X1 U17182 ( .A(n15565), .ZN(n15567) );
  OAI21_X1 U17183 ( .B1(n15725), .B2(n15567), .A(n15566), .ZN(n15568) );
  NAND3_X1 U17184 ( .A1(n15639), .A2(n15569), .A3(n15568), .ZN(n15575) );
  OAI211_X1 U17185 ( .C1(n15572), .C2(n15571), .A(n15644), .B(n15570), .ZN(
        n15574) );
  NAND2_X1 U17186 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n15635), .ZN(n15573) );
  NAND4_X1 U17187 ( .A1(n15576), .A2(n15575), .A3(n15574), .A4(n15573), .ZN(
        P2_U3215) );
  INV_X1 U17188 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15593) );
  NOR2_X1 U17189 ( .A1(n15578), .A2(n15577), .ZN(n15579) );
  OAI21_X1 U17190 ( .B1(n15580), .B2(n15579), .A(n15639), .ZN(n15589) );
  AND3_X1 U17191 ( .A1(n15583), .A2(n15582), .A3(n15581), .ZN(n15584) );
  OAI21_X1 U17192 ( .B1(n15585), .B2(n15584), .A(n15644), .ZN(n15588) );
  NAND2_X1 U17193 ( .A1(n15641), .A2(n15586), .ZN(n15587) );
  AND3_X1 U17194 ( .A1(n15589), .A2(n15588), .A3(n15587), .ZN(n15591) );
  OAI211_X1 U17195 ( .C1(n15593), .C2(n15592), .A(n15591), .B(n15590), .ZN(
        P2_U3226) );
  AOI22_X1 U17196 ( .A1(n15635), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3088), .ZN(n15604) );
  NAND2_X1 U17197 ( .A1(n15641), .A2(n15594), .ZN(n15603) );
  OAI211_X1 U17198 ( .C1(n15597), .C2(n15596), .A(n15595), .B(n15639), .ZN(
        n15602) );
  OAI211_X1 U17199 ( .C1(n15600), .C2(n15599), .A(n15598), .B(n15644), .ZN(
        n15601) );
  NAND4_X1 U17200 ( .A1(n15604), .A2(n15603), .A3(n15602), .A4(n15601), .ZN(
        P2_U3227) );
  AOI22_X1 U17201 ( .A1(n15635), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(P2_U3088), .ZN(n15614) );
  NAND2_X1 U17202 ( .A1(n15641), .A2(n15605), .ZN(n15613) );
  OAI211_X1 U17203 ( .C1(n15607), .C2(P2_REG2_REG_14__SCAN_IN), .A(n15606), 
        .B(n15644), .ZN(n15612) );
  OAI211_X1 U17204 ( .C1(n15610), .C2(n15609), .A(n15608), .B(n15639), .ZN(
        n15611) );
  NAND4_X1 U17205 ( .A1(n15614), .A2(n15613), .A3(n15612), .A4(n15611), .ZN(
        P2_U3228) );
  AOI22_X1 U17206 ( .A1(n15635), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n15623) );
  NAND2_X1 U17207 ( .A1(n15641), .A2(n15615), .ZN(n15622) );
  OAI211_X1 U17208 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n15617), .A(n15644), 
        .B(n15616), .ZN(n15621) );
  OAI211_X1 U17209 ( .C1(n15619), .C2(P2_REG1_REG_15__SCAN_IN), .A(n15639), 
        .B(n15618), .ZN(n15620) );
  NAND4_X1 U17210 ( .A1(n15623), .A2(n15622), .A3(n15621), .A4(n15620), .ZN(
        P2_U3229) );
  AOI22_X1 U17211 ( .A1(n15635), .A2(P2_ADDR_REG_16__SCAN_IN), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(P2_U3088), .ZN(n15634) );
  OAI211_X1 U17212 ( .C1(n15626), .C2(n15625), .A(n15644), .B(n15624), .ZN(
        n15633) );
  NAND2_X1 U17213 ( .A1(n15641), .A2(n15627), .ZN(n15632) );
  OAI211_X1 U17214 ( .C1(n15630), .C2(n15629), .A(n15639), .B(n15628), .ZN(
        n15631) );
  NAND4_X1 U17215 ( .A1(n15634), .A2(n15633), .A3(n15632), .A4(n15631), .ZN(
        P2_U3230) );
  AOI22_X1 U17216 ( .A1(n15635), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(P2_U3088), .ZN(n15650) );
  XOR2_X1 U17217 ( .A(n15637), .B(n15636), .Z(n15638) );
  NAND2_X1 U17218 ( .A1(n15639), .A2(n15638), .ZN(n15649) );
  NAND2_X1 U17219 ( .A1(n15641), .A2(n15640), .ZN(n15648) );
  INV_X1 U17220 ( .A(n15642), .ZN(n15646) );
  OAI211_X1 U17221 ( .C1(n15646), .C2(n15645), .A(n15644), .B(n15643), .ZN(
        n15647) );
  NAND4_X1 U17222 ( .A1(n15650), .A2(n15649), .A3(n15648), .A4(n15647), .ZN(
        P2_U3231) );
  NOR2_X1 U17223 ( .A1(n15652), .A2(n15651), .ZN(n15679) );
  INV_X1 U17224 ( .A(n15679), .ZN(n15655) );
  OAI22_X1 U17225 ( .A1(n15658), .A2(n15655), .B1(n15654), .B2(n15653), .ZN(
        n15656) );
  INV_X1 U17226 ( .A(n15656), .ZN(n15667) );
  OAI21_X1 U17227 ( .B1(n15711), .B2(n15658), .A(n15657), .ZN(n15660) );
  MUX2_X1 U17228 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n15660), .S(n15659), .Z(
        n15665) );
  OAI22_X1 U17229 ( .A1(n15663), .A2(n15662), .B1(n15676), .B2(n15661), .ZN(
        n15664) );
  NOR2_X1 U17230 ( .A1(n15665), .A2(n15664), .ZN(n15666) );
  NAND2_X1 U17231 ( .A1(n15667), .A2(n15666), .ZN(P2_U3261) );
  INV_X1 U17232 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n15675) );
  NAND2_X1 U17233 ( .A1(n15711), .A2(n15668), .ZN(n15671) );
  INV_X1 U17234 ( .A(n15669), .ZN(n15670) );
  AOI21_X1 U17235 ( .B1(n15693), .B2(n15671), .A(n15670), .ZN(n15695) );
  NAND2_X1 U17236 ( .A1(n15672), .A2(n13804), .ZN(n15673) );
  NAND2_X1 U17237 ( .A1(n15673), .A2(n15691), .ZN(n15674) );
  OAI211_X1 U17238 ( .C1(n15676), .C2(n15675), .A(n15695), .B(n15674), .ZN(
        n15677) );
  INV_X1 U17239 ( .A(n15677), .ZN(n15681) );
  AOI22_X1 U17240 ( .A1(n15679), .A2(n15693), .B1(P2_REG2_REG_0__SCAN_IN), 
        .B2(n15678), .ZN(n15680) );
  OAI21_X1 U17241 ( .B1(n15678), .B2(n15681), .A(n15680), .ZN(P2_U3265) );
  AND2_X1 U17242 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15683), .ZN(P2_U3266) );
  AND2_X1 U17243 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15683), .ZN(P2_U3267) );
  AND2_X1 U17244 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15683), .ZN(P2_U3268) );
  AND2_X1 U17245 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15683), .ZN(P2_U3269) );
  AND2_X1 U17246 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15683), .ZN(P2_U3270) );
  AND2_X1 U17247 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15683), .ZN(P2_U3271) );
  AND2_X1 U17248 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15683), .ZN(P2_U3272) );
  AND2_X1 U17249 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15683), .ZN(P2_U3273) );
  AND2_X1 U17250 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15683), .ZN(P2_U3274) );
  AND2_X1 U17251 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15683), .ZN(P2_U3275) );
  AND2_X1 U17252 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15683), .ZN(P2_U3276) );
  AND2_X1 U17253 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15683), .ZN(P2_U3277) );
  AND2_X1 U17254 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15683), .ZN(P2_U3278) );
  AND2_X1 U17255 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15683), .ZN(P2_U3279) );
  AND2_X1 U17256 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15683), .ZN(P2_U3280) );
  AND2_X1 U17257 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15683), .ZN(P2_U3281) );
  AND2_X1 U17258 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15683), .ZN(P2_U3282) );
  AND2_X1 U17259 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15683), .ZN(P2_U3283) );
  AND2_X1 U17260 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15683), .ZN(P2_U3284) );
  AND2_X1 U17261 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15683), .ZN(P2_U3285) );
  AND2_X1 U17262 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15683), .ZN(P2_U3286) );
  AND2_X1 U17263 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15683), .ZN(P2_U3287) );
  AND2_X1 U17264 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15683), .ZN(P2_U3288) );
  AND2_X1 U17265 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15683), .ZN(P2_U3289) );
  AND2_X1 U17266 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15683), .ZN(P2_U3290) );
  AND2_X1 U17267 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15683), .ZN(P2_U3291) );
  AND2_X1 U17268 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15683), .ZN(P2_U3292) );
  AND2_X1 U17269 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15683), .ZN(P2_U3293) );
  AND2_X1 U17270 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15683), .ZN(P2_U3294) );
  AND2_X1 U17271 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15683), .ZN(P2_U3295) );
  AOI22_X1 U17272 ( .A1(n15689), .A2(n15685), .B1(n15684), .B2(n15686), .ZN(
        P2_U3416) );
  AOI22_X1 U17273 ( .A1(n15689), .A2(n15688), .B1(n15687), .B2(n15686), .ZN(
        P2_U3417) );
  AOI22_X1 U17274 ( .A1(n15693), .A2(n15692), .B1(n15691), .B2(n15690), .ZN(
        n15694) );
  AND2_X1 U17275 ( .A1(n15695), .A2(n15694), .ZN(n15726) );
  INV_X1 U17276 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15696) );
  AOI22_X1 U17277 ( .A1(n15724), .A2(n15726), .B1(n15696), .B2(n9771), .ZN(
        P2_U3430) );
  OAI21_X1 U17278 ( .B1(n15698), .B2(n15718), .A(n15697), .ZN(n15701) );
  INV_X1 U17279 ( .A(n15699), .ZN(n15700) );
  AOI211_X1 U17280 ( .C1(n15702), .C2(n15722), .A(n15701), .B(n15700), .ZN(
        n15727) );
  INV_X1 U17281 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n15703) );
  AOI22_X1 U17282 ( .A1(n15724), .A2(n15727), .B1(n15703), .B2(n9771), .ZN(
        P2_U3433) );
  INV_X1 U17283 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15704) );
  AOI22_X1 U17284 ( .A1(n15724), .A2(n15705), .B1(n15704), .B2(n9771), .ZN(
        P2_U3436) );
  OAI211_X1 U17285 ( .C1(n15708), .C2(n15718), .A(n15707), .B(n15706), .ZN(
        n15713) );
  AOI21_X1 U17286 ( .B1(n15711), .B2(n15710), .A(n15709), .ZN(n15712) );
  NOR2_X1 U17287 ( .A1(n15713), .A2(n15712), .ZN(n15728) );
  INV_X1 U17288 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15714) );
  AOI22_X1 U17289 ( .A1(n15724), .A2(n15728), .B1(n15714), .B2(n9771), .ZN(
        P2_U3439) );
  INV_X1 U17290 ( .A(n15715), .ZN(n15720) );
  INV_X1 U17291 ( .A(n15716), .ZN(n15717) );
  OAI21_X1 U17292 ( .B1(n7476), .B2(n15718), .A(n15717), .ZN(n15719) );
  AOI211_X1 U17293 ( .C1(n15722), .C2(n15721), .A(n15720), .B(n15719), .ZN(
        n15730) );
  INV_X1 U17294 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n15723) );
  AOI22_X1 U17295 ( .A1(n15724), .A2(n15730), .B1(n15723), .B2(n9771), .ZN(
        P2_U3463) );
  AOI22_X1 U17296 ( .A1(n15731), .A2(n15726), .B1(n15725), .B2(n15729), .ZN(
        P2_U3499) );
  AOI22_X1 U17297 ( .A1(n15731), .A2(n15727), .B1(n10754), .B2(n15729), .ZN(
        P2_U3500) );
  AOI22_X1 U17298 ( .A1(n15731), .A2(n15728), .B1(n10815), .B2(n15729), .ZN(
        P2_U3502) );
  AOI22_X1 U17299 ( .A1(n15731), .A2(n15730), .B1(n12338), .B2(n15729), .ZN(
        P2_U3510) );
  NOR2_X1 U17300 ( .A1(P3_U3897), .A2(n15732), .ZN(P3_U3150) );
  AOI21_X1 U17301 ( .B1(n15735), .B2(n15734), .A(n15733), .ZN(n15753) );
  OAI22_X1 U17302 ( .A1(n15738), .A2(n12426), .B1(n15737), .B2(n15736), .ZN(
        n15749) );
  AOI21_X1 U17303 ( .B1(n15741), .B2(n15740), .A(n15739), .ZN(n15747) );
  AOI21_X1 U17304 ( .B1(n8015), .B2(n15743), .A(n15742), .ZN(n15745) );
  OAI22_X1 U17305 ( .A1(n15747), .A2(n15746), .B1(n15745), .B2(n15744), .ZN(
        n15748) );
  NOR3_X1 U17306 ( .A1(n15750), .A2(n15749), .A3(n15748), .ZN(n15751) );
  OAI21_X1 U17307 ( .B1(n15753), .B2(n15752), .A(n15751), .ZN(P3_U3193) );
  INV_X1 U17308 ( .A(n15754), .ZN(n15775) );
  INV_X1 U17309 ( .A(n15755), .ZN(n15757) );
  OAI21_X1 U17310 ( .B1(n15775), .B2(n15757), .A(n15756), .ZN(n15762) );
  OAI22_X1 U17311 ( .A1(n15760), .A2(n15759), .B1(n15758), .B2(n15801), .ZN(
        n15761) );
  AOI21_X1 U17312 ( .B1(n15762), .B2(n15801), .A(n15761), .ZN(n15763) );
  OAI21_X1 U17313 ( .B1(n15764), .B2(n15782), .A(n15763), .ZN(P3_U3225) );
  INV_X1 U17314 ( .A(n15765), .ZN(n15767) );
  OAI21_X1 U17315 ( .B1(n15775), .B2(n15767), .A(n15766), .ZN(n15768) );
  MUX2_X1 U17316 ( .A(n15768), .B(P3_REG2_REG_7__SCAN_IN), .S(n15822), .Z(
        n15769) );
  AOI21_X1 U17317 ( .B1(n15780), .B2(n15770), .A(n15769), .ZN(n15771) );
  OAI21_X1 U17318 ( .B1(n15772), .B2(n15782), .A(n15771), .ZN(P3_U3226) );
  INV_X1 U17319 ( .A(n15773), .ZN(n15776) );
  OAI21_X1 U17320 ( .B1(n15776), .B2(n15775), .A(n15774), .ZN(n15777) );
  MUX2_X1 U17321 ( .A(P3_REG2_REG_3__SCAN_IN), .B(n15777), .S(n15801), .Z(
        n15778) );
  AOI21_X1 U17322 ( .B1(n15780), .B2(n15779), .A(n15778), .ZN(n15781) );
  OAI21_X1 U17323 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(n15782), .A(n15781), .ZN(
        P3_U3230) );
  XNOR2_X1 U17324 ( .A(n15783), .B(n15785), .ZN(n15793) );
  OAI21_X1 U17325 ( .B1(n15786), .B2(n15785), .A(n15784), .ZN(n15794) );
  OAI22_X1 U17326 ( .A1(n15790), .A2(n15789), .B1(n15788), .B2(n15787), .ZN(
        n15791) );
  AOI21_X1 U17327 ( .B1(n15794), .B2(n15814), .A(n15791), .ZN(n15792) );
  OAI21_X1 U17328 ( .B1(n15811), .B2(n15793), .A(n15792), .ZN(n15828) );
  INV_X1 U17329 ( .A(n15794), .ZN(n15832) );
  INV_X1 U17330 ( .A(n15795), .ZN(n15799) );
  NAND2_X1 U17331 ( .A1(n15797), .A2(n15796), .ZN(n15829) );
  OAI22_X1 U17332 ( .A1(n15832), .A2(n15799), .B1(n15798), .B2(n15829), .ZN(
        n15800) );
  AOI211_X1 U17333 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15818), .A(n15828), .B(
        n15800), .ZN(n15802) );
  AOI22_X1 U17334 ( .A1(n15822), .A2(n10641), .B1(n15802), .B2(n15801), .ZN(
        P3_U3231) );
  XNOR2_X1 U17335 ( .A(n11259), .B(n15803), .ZN(n15826) );
  XNOR2_X1 U17336 ( .A(n15805), .B(n15804), .ZN(n15812) );
  AOI22_X1 U17337 ( .A1(n15809), .A2(n15808), .B1(n15807), .B2(n15806), .ZN(
        n15810) );
  OAI21_X1 U17338 ( .B1(n15812), .B2(n15811), .A(n15810), .ZN(n15813) );
  AOI21_X1 U17339 ( .B1(n15814), .B2(n15826), .A(n15813), .ZN(n15823) );
  NOR2_X1 U17340 ( .A1(n15816), .A2(n15815), .ZN(n15825) );
  AOI22_X1 U17341 ( .A1(n15818), .A2(P3_REG3_REG_1__SCAN_IN), .B1(n15825), 
        .B2(n15817), .ZN(n15821) );
  AOI22_X1 U17342 ( .A1(n15819), .A2(n15826), .B1(n15822), .B2(
        P3_REG2_REG_1__SCAN_IN), .ZN(n15820) );
  OAI221_X1 U17343 ( .B1(n15822), .B2(n15823), .C1(n15822), .C2(n15821), .A(
        n15820), .ZN(P3_U3232) );
  INV_X1 U17344 ( .A(n15823), .ZN(n15824) );
  AOI211_X1 U17345 ( .C1(n15842), .C2(n15826), .A(n15825), .B(n15824), .ZN(
        n15847) );
  INV_X1 U17346 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15827) );
  AOI22_X1 U17347 ( .A1(n15846), .A2(n15847), .B1(n15827), .B2(n15844), .ZN(
        P3_U3393) );
  INV_X1 U17348 ( .A(n15828), .ZN(n15830) );
  OAI211_X1 U17349 ( .C1(n15832), .C2(n15831), .A(n15830), .B(n15829), .ZN(
        n15848) );
  OAI22_X1 U17350 ( .A1(n15844), .A2(n15848), .B1(P3_REG0_REG_2__SCAN_IN), 
        .B2(n15846), .ZN(n15833) );
  INV_X1 U17351 ( .A(n15833), .ZN(P3_U3396) );
  INV_X1 U17352 ( .A(n15834), .ZN(n15838) );
  INV_X1 U17353 ( .A(n15835), .ZN(n15836) );
  AOI211_X1 U17354 ( .C1(n15838), .C2(n15842), .A(n15837), .B(n15836), .ZN(
        n15850) );
  INV_X1 U17355 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15839) );
  AOI22_X1 U17356 ( .A1(n15846), .A2(n15850), .B1(n15839), .B2(n15844), .ZN(
        P3_U3405) );
  AOI211_X1 U17357 ( .C1(n15843), .C2(n15842), .A(n15841), .B(n15840), .ZN(
        n15853) );
  INV_X1 U17358 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15845) );
  AOI22_X1 U17359 ( .A1(n15846), .A2(n15853), .B1(n15845), .B2(n15844), .ZN(
        P3_U3420) );
  AOI22_X1 U17360 ( .A1(n15854), .A2(n15847), .B1(n10634), .B2(n15851), .ZN(
        P3_U3460) );
  OAI22_X1 U17361 ( .A1(n15851), .A2(n15848), .B1(P3_REG1_REG_2__SCAN_IN), 
        .B2(n15854), .ZN(n15849) );
  INV_X1 U17362 ( .A(n15849), .ZN(P3_U3461) );
  AOI22_X1 U17363 ( .A1(n15854), .A2(n15850), .B1(n10657), .B2(n15851), .ZN(
        P3_U3464) );
  AOI22_X1 U17364 ( .A1(n15854), .A2(n15853), .B1(n15852), .B2(n15851), .ZN(
        P3_U3469) );
  AOI21_X1 U17365 ( .B1(n15857), .B2(n15856), .A(n15855), .ZN(SUB_1596_U59) );
  OAI21_X1 U17366 ( .B1(n15860), .B2(n15859), .A(n15858), .ZN(SUB_1596_U58) );
  XNOR2_X1 U17367 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15861), .ZN(SUB_1596_U53)
         );
  OAI21_X1 U17368 ( .B1(n15864), .B2(n15863), .A(n15862), .ZN(SUB_1596_U56) );
  AOI21_X1 U17369 ( .B1(n15867), .B2(n15866), .A(n15865), .ZN(n15868) );
  XOR2_X1 U17370 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15868), .Z(SUB_1596_U60) );
  AOI21_X1 U17371 ( .B1(n15871), .B2(n15870), .A(n15869), .ZN(SUB_1596_U5) );
  CLKBUF_X1 U7417 ( .A(n8267), .Z(n10612) );
  CLKBUF_X1 U7434 ( .A(n10512), .Z(n12785) );
  CLKBUF_X1 U7435 ( .A(n8062), .Z(n8328) );
  NOR2_X2 U7438 ( .A1(n14134), .A2(n14310), .ZN(n14125) );
  CLKBUF_X1 U7478 ( .A(n7909), .Z(n8331) );
  CLKBUF_X1 U7805 ( .A(n10069), .Z(n10418) );
  XNOR2_X1 U9387 ( .A(n7234), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9931) );
endmodule

