

module b17_C_gen_AntiSAT_k_128_10 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput_f0, keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, 
        keyinput_f5, keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, 
        keyinput_f10, keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, 
        keyinput_f15, keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, 
        keyinput_f20, keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, 
        keyinput_f25, keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, 
        keyinput_f30, keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, 
        keyinput_f35, keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, 
        keyinput_f40, keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, 
        keyinput_f45, keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, 
        keyinput_f50, keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, 
        keyinput_f55, keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, 
        keyinput_f60, keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, 
        keyinput_g1, keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, 
        keyinput_g6, keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, 
        keyinput_g11, keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, 
        keyinput_g16, keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, 
        keyinput_g21, keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, 
        keyinput_g26, keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, 
        keyinput_g31, keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, 
        keyinput_g36, keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, 
        keyinput_g41, keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, 
        keyinput_g46, keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, 
        keyinput_g51, keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, 
        keyinput_g56, keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, 
        keyinput_g61, keyinput_g62, keyinput_g63, U355, U356, U357, U358, U359, 
        U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, 
        U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, 
        U376, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, 
        U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, 
        U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, 
        U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, 
        U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, 
        U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, 
        P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, 
        P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, 
        P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, 
        P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, 
        P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, 
        P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, 
        P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, 
        P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, 
        P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, 
        P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, 
        P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, 
        P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, 
        P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, 
        P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, 
        P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, 
        P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, 
        P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, 
        P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, 
        P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, 
        P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, 
        P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, 
        P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, 
        P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, 
        P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, 
        P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, 
        P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, 
        P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, 
        P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, 
        P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, 
        P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, 
        P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, 
        P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, 
        P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, 
        P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, 
        P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, 
        P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, 
        P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, 
        P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, 
        P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, 
        P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, 
        P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, 
        P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, 
        P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, 
        P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, 
        P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, 
        P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, 
        P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, 
        P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, 
        P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, 
        P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, 
        P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, 
        P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, 
        P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, 
        P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, 
        P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, 
        P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, 
        P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, 
        P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, 
        P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, 
        P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, 
        P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, 
        P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, 
        P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, 
        P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, 
        P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, 
        P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, 
        P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, 
        P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, 
        P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, 
        P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, 
        P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, 
        P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, 
        P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, 
        P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, 
        P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, 
        P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, 
        P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, 
        P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, 
        P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, 
        P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, 
        P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, 
        P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, 
        P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, 
        P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, 
        P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, 
        P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, 
        P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, 
        P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, 
        P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, 
        P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, 
        P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, 
        P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, 
        P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, 
        P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, 
        P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, 
        P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, 
        P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, 
        P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, 
        P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, 
        P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, 
        P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, 
        P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, 
        P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, 
        P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, 
        P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, 
        P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, 
        P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, 
        P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, 
        P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, 
        P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, 
        P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, 
        P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, 
        P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, 
        P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, 
        P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, 
        P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, 
        P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, 
        P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, 
        P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, 
        P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, 
        P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, 
        P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, 
        P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, 
        P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, 
        P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, 
        P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, 
        P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, 
        P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, 
        P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, 
        P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, 
        P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, 
        P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, 
        P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, 
        P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, 
        P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, 
        P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, 
        P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, 
        P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, 
        P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, 
        P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, 
        P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, 
        P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, 
        P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, 
        P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, 
        P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, 
        P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, 
        P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, 
        P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, 
        P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, 
        P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, 
        P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, 
        P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, 
        P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, 
        P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, 
        P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, 
        P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, 
        P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, 
        P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, 
        P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, 
        P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, 
        P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, 
        P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, 
        P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, 
        P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, 
        P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, 
        P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, 
        P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, 
        P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, 
        P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, 
        P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, 
        P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, 
        P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, 
        P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, 
        P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, 
        P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, 
        P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, 
        P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, 
        P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, 
        P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, 
        P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, 
        P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9649, n9650,
         n9651, n9652, n9653, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
         n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
         n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
         n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
         n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
         n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938,
         n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
         n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954,
         n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
         n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970,
         n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978,
         n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986,
         n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
         n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002,
         n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010,
         n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
         n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026,
         n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
         n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
         n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050,
         n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058,
         n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
         n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074,
         n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082,
         n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
         n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098,
         n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
         n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114,
         n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122,
         n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130,
         n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
         n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146,
         n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154,
         n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
         n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
         n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
         n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186,
         n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194,
         n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
         n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
         n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218,
         n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226,
         n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
         n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
         n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258,
         n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266,
         n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274,
         n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
         n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
         n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
         n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
         n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314,
         n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322,
         n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330,
         n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338,
         n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346,
         n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
         n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362,
         n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
         n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
         n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386,
         n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
         n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402,
         n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
         n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418,
         n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
         n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434,
         n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442,
         n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
         n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458,
         n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
         n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474,
         n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
         n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
         n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
         n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506,
         n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
         n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
         n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530,
         n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538,
         n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546,
         n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
         n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562,
         n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
         n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578,
         n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
         n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
         n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
         n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
         n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618,
         n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
         n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
         n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
         n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650,
         n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658,
         n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
         n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674,
         n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682,
         n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690,
         n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
         n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
         n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
         n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
         n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
         n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
         n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762,
         n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770,
         n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
         n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
         n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794,
         n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
         n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
         n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
         n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
         n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
         n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
         n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
         n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
         n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
         n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
         n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
         n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
         n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
         n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
         n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
         n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
         n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
         n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
         n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026,
         n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
         n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
         n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
         n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058,
         n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066,
         n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074,
         n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
         n21083;

  CLKBUF_X1 U11074 ( .A(n17900), .Z(n9676) );
  NOR2_X2 U11075 ( .A1(n12576), .A2(n14718), .ZN(n12577) );
  OR2_X1 U11076 ( .A1(n16070), .A2(n10188), .ZN(n10186) );
  OR2_X1 U11077 ( .A1(n15259), .A2(n16198), .ZN(n10295) );
  NOR2_X1 U11078 ( .A1(n18723), .A2(n18114), .ZN(n18202) );
  NOR2_X1 U11079 ( .A1(n20051), .A2(n12464), .ZN(n20016) );
  INV_X1 U11080 ( .A(n18906), .ZN(n16530) );
  NAND2_X2 U11081 ( .A1(n10178), .A2(n10177), .ZN(n14079) );
  NAND4_X1 U11082 ( .A1(n11686), .A2(n9816), .A3(n9815), .A4(n9814), .ZN(
        n11794) );
  AND2_X1 U11083 ( .A1(n10667), .A2(n12910), .ZN(n19752) );
  AND2_X1 U11084 ( .A1(n10671), .A2(n12910), .ZN(n19525) );
  AND2_X1 U11085 ( .A1(n10669), .A2(n12910), .ZN(n19584) );
  INV_X1 U11086 ( .A(n13380), .ZN(n19956) );
  AOI211_X1 U11087 ( .C1(n11207), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n11234), .B(n11233), .ZN(n17387) );
  CLKBUF_X2 U11089 ( .A(n12668), .Z(n10770) );
  INV_X1 U11090 ( .A(n13803), .ZN(n11643) );
  AND2_X1 U11091 ( .A1(n9656), .A2(n10510), .ZN(n10721) );
  AND2_X1 U11092 ( .A1(n9656), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10382) );
  AND2_X1 U11093 ( .A1(n13187), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10381) );
  AND2_X1 U11094 ( .A1(n10543), .A2(n10510), .ZN(n13039) );
  BUF_X1 U11095 ( .A(n10546), .Z(n13116) );
  NAND2_X2 U11096 ( .A1(n12442), .A2(n9662), .ZN(n12446) );
  INV_X2 U11097 ( .A(n11148), .ZN(n17133) );
  BUF_X1 U11098 ( .A(n11189), .Z(n9644) );
  INV_X4 U11099 ( .A(n9746), .ZN(n17212) );
  INV_X2 U11100 ( .A(n17223), .ZN(n17167) );
  NAND2_X1 U11101 ( .A1(n10568), .A2(n16342), .ZN(n13347) );
  AND2_X1 U11102 ( .A1(n10569), .A2(n19237), .ZN(n10603) );
  BUF_X1 U11103 ( .A(n12089), .Z(n9666) );
  INV_X2 U11104 ( .A(n19237), .ZN(n13586) );
  CLKBUF_X2 U11105 ( .A(n12261), .Z(n9669) );
  CLKBUF_X2 U11106 ( .A(n11571), .Z(n9673) );
  CLKBUF_X2 U11107 ( .A(n11531), .Z(n9661) );
  INV_X1 U11108 ( .A(n12186), .ZN(n12259) );
  INV_X1 U11109 ( .A(n12190), .ZN(n12232) );
  INV_X1 U11110 ( .A(n12190), .ZN(n12261) );
  BUF_X1 U11112 ( .A(n10542), .Z(n9651) );
  BUF_X1 U11113 ( .A(n10542), .Z(n9653) );
  NOR2_X2 U11114 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14180) );
  INV_X1 U11115 ( .A(n18759), .ZN(n9630) );
  INV_X1 U11116 ( .A(n9630), .ZN(n9631) );
  INV_X1 U11117 ( .A(n9630), .ZN(n9632) );
  INV_X1 U11118 ( .A(n19823), .ZN(n9633) );
  INV_X1 U11119 ( .A(n9633), .ZN(n9634) );
  INV_X1 U11120 ( .A(n9633), .ZN(n9635) );
  AND2_X1 U11121 ( .A1(n13806), .A2(n11513), .ZN(n11571) );
  CLKBUF_X2 U11122 ( .A(n11570), .Z(n12237) );
  INV_X1 U11123 ( .A(n10423), .ZN(n13036) );
  AOI21_X1 U11124 ( .B1(n11112), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n10597), .ZN(n10600) );
  AND2_X1 U11125 ( .A1(n13810), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13672) );
  AND2_X1 U11126 ( .A1(n9645), .A2(n10517), .ZN(n10421) );
  AND2_X1 U11127 ( .A1(n9652), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12716) );
  AND2_X1 U11128 ( .A1(n10673), .A2(n12910), .ZN(n19654) );
  AND2_X1 U11129 ( .A1(n12910), .A2(n19193), .ZN(n10675) );
  NOR2_X1 U11130 ( .A1(n10509), .A2(n10508), .ZN(n10581) );
  NAND2_X1 U11132 ( .A1(n20220), .A2(n13654), .ZN(n13770) );
  NAND2_X1 U11133 ( .A1(n10000), .A2(n11655), .ZN(n11800) );
  INV_X2 U11134 ( .A(n17116), .ZN(n17214) );
  BUF_X1 U11135 ( .A(n18114), .Z(n9640) );
  NAND2_X1 U11136 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18690) );
  INV_X1 U11137 ( .A(n20027), .ZN(n20053) );
  INV_X1 U11138 ( .A(n13717), .ZN(n12361) );
  OAI21_X1 U11139 ( .B1(n15162), .B2(n10928), .A(n9731), .ZN(n9893) );
  INV_X1 U11140 ( .A(n12794), .ZN(n12877) );
  INV_X1 U11141 ( .A(n11287), .ZN(n17213) );
  AND2_X1 U11142 ( .A1(n14217), .A2(n12484), .ZN(n20027) );
  BUF_X1 U11143 ( .A(n12589), .Z(n9641) );
  NAND2_X2 U11144 ( .A1(n10064), .A2(n11586), .ZN(n13654) );
  AND2_X1 U11145 ( .A1(n15534), .A2(n10104), .ZN(n15175) );
  INV_X2 U11146 ( .A(n16846), .ZN(n16858) );
  INV_X1 U11147 ( .A(n17673), .ZN(n17890) );
  NAND2_X1 U11148 ( .A1(n18202), .A2(n18703), .ZN(n18125) );
  NOR2_X1 U11149 ( .A1(n17644), .A2(n17614), .ZN(n17673) );
  AND2_X1 U11150 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n9636) );
  BUF_X1 U11151 ( .A(n11028), .Z(n11105) );
  XNOR2_X1 U11152 ( .A(n10657), .B(n9865), .ZN(n10664) );
  CLKBUF_X3 U11153 ( .A(n11543), .Z(n9675) );
  CLKBUF_X3 U11154 ( .A(n11543), .Z(n12116) );
  NOR2_X1 U11155 ( .A1(n18880), .A2(n18872), .ZN(n18691) );
  NOR2_X2 U11156 ( .A1(n14361), .A2(n10265), .ZN(n14310) );
  NOR2_X4 U11157 ( .A1(n15025), .A2(n12941), .ZN(n15004) );
  NAND2_X2 U11159 ( .A1(n10244), .A2(n9769), .ZN(n11719) );
  OR3_X2 U11160 ( .A1(n11215), .A2(n11214), .A3(n11213), .ZN(n17409) );
  NOR3_X2 U11161 ( .A1(n14275), .A2(n20948), .A3(n20835), .ZN(n14250) );
  AND2_X2 U11162 ( .A1(n14181), .A2(n10639), .ZN(n9637) );
  NAND2_X1 U11163 ( .A1(n11604), .A2(n13654), .ZN(n12442) );
  NOR2_X2 U11164 ( .A1(n15181), .A2(n15374), .ZN(n10915) );
  AND2_X2 U11165 ( .A1(n15582), .A2(n10325), .ZN(n9656) );
  AND2_X2 U11166 ( .A1(n15582), .A2(n10325), .ZN(n9657) );
  AND2_X1 U11167 ( .A1(n13672), .A2(n13807), .ZN(n9639) );
  NOR2_X2 U11168 ( .A1(n15174), .A2(n14858), .ZN(n14857) );
  AND2_X2 U11169 ( .A1(n10192), .A2(n10190), .ZN(n14858) );
  AND2_X2 U11170 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14181) );
  NOR2_X1 U11171 ( .A1(n15218), .A2(n13255), .ZN(n13254) );
  AND2_X4 U11172 ( .A1(n14180), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10478) );
  OAI21_X1 U11173 ( .B1(n18682), .B2(n18694), .A(n18681), .ZN(n18114) );
  AND2_X2 U11174 ( .A1(n10675), .A2(n10674), .ZN(n19552) );
  NOR2_X2 U11175 ( .A1(n18993), .A2(n16056), .ZN(n12661) );
  INV_X1 U11176 ( .A(n11105), .ZN(n9642) );
  INV_X2 U11177 ( .A(n9642), .ZN(n9643) );
  NOR3_X1 U11178 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n18690), .ZN(n11189) );
  XNOR2_X2 U11179 ( .A(n11800), .B(n11801), .ZN(n12509) );
  AND2_X4 U11180 ( .A1(n10328), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13066) );
  NAND2_X1 U11181 ( .A1(n14557), .A2(n10254), .ZN(n14387) );
  NAND2_X1 U11182 ( .A1(n10237), .A2(n10236), .ZN(n13860) );
  INV_X4 U11183 ( .A(n10313), .ZN(n15883) );
  OAI22_X1 U11184 ( .A1(n17762), .A2(n17901), .B1(n17809), .B2(n17760), .ZN(
        n17773) );
  NOR2_X1 U11185 ( .A1(n18733), .A2(n18747), .ZN(n11490) );
  NAND2_X1 U11186 ( .A1(n20075), .A2(n13725), .ZN(n14480) );
  NOR2_X2 U11187 ( .A1(n16530), .A2(n18125), .ZN(n18722) );
  NAND2_X1 U11188 ( .A1(n11681), .A2(n20315), .ZN(n11704) );
  NAND2_X1 U11189 ( .A1(n17381), .A2(n11463), .ZN(n17737) );
  NOR2_X1 U11190 ( .A1(n17478), .A2(n11435), .ZN(n16510) );
  CLKBUF_X1 U11191 ( .A(n11112), .Z(n11118) );
  AOI211_X1 U11192 ( .C1(n18245), .C2(n11408), .A(n11407), .B(n11406), .ZN(
        n11436) );
  NOR2_X1 U11193 ( .A1(n9916), .A2(n11616), .ZN(n11617) );
  OR2_X1 U11194 ( .A1(n11613), .A2(n13542), .ZN(n9916) );
  BUF_X1 U11195 ( .A(n18250), .Z(n9677) );
  INV_X1 U11196 ( .A(n13770), .ZN(n20873) );
  NAND2_X2 U11197 ( .A1(n11724), .A2(n12496), .ZN(n12335) );
  NAND2_X4 U11198 ( .A1(n9689), .A2(n9727), .ZN(n9926) );
  INV_X1 U11199 ( .A(n10587), .ZN(n12670) );
  NAND2_X2 U11200 ( .A1(n10006), .A2(n10009), .ZN(n10559) );
  AOI211_X1 U11201 ( .C1(n17049), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n11295), .B(n11294), .ZN(n11296) );
  AND2_X1 U11202 ( .A1(n10373), .A2(n10010), .ZN(n10554) );
  INV_X1 U11203 ( .A(n19220), .ZN(n16342) );
  NAND2_X2 U11204 ( .A1(n9960), .A2(n9959), .ZN(n11576) );
  NAND2_X1 U11205 ( .A1(n10489), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10009) );
  CLKBUF_X3 U11207 ( .A(n17206), .Z(n9649) );
  INV_X4 U11208 ( .A(n17191), .ZN(n11202) );
  BUF_X2 U11209 ( .A(n13046), .Z(n9650) );
  BUF_X2 U11210 ( .A(n11993), .Z(n12208) );
  CLKBUF_X2 U11211 ( .A(n11846), .Z(n12250) );
  CLKBUF_X2 U11212 ( .A(n11571), .Z(n9674) );
  CLKBUF_X2 U11213 ( .A(n13047), .Z(n10330) );
  BUF_X2 U11214 ( .A(n11531), .Z(n9660) );
  CLKBUF_X2 U11215 ( .A(n11664), .Z(n12094) );
  CLKBUF_X2 U11216 ( .A(n11879), .Z(n12165) );
  CLKBUF_X2 U11217 ( .A(n10542), .Z(n9652) );
  BUF_X2 U11218 ( .A(n11531), .Z(n9659) );
  BUF_X4 U11220 ( .A(n10542), .Z(n9645) );
  INV_X2 U11221 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13807) );
  NOR2_X4 U11222 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11513) );
  OR2_X1 U11223 ( .A1(n15136), .A2(n10279), .ZN(n10275) );
  AOI21_X1 U11224 ( .B1(n15155), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n9891), .ZN(n15147) );
  OAI21_X1 U11225 ( .B1(n15333), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15150), .ZN(n15319) );
  AND2_X1 U11226 ( .A1(n9893), .A2(n15144), .ZN(n9891) );
  XNOR2_X1 U11227 ( .A(n9893), .B(n9892), .ZN(n15155) );
  AND2_X1 U11228 ( .A1(n16181), .A2(n16180), .ZN(n16273) );
  NOR2_X1 U11229 ( .A1(n15161), .A2(n15311), .ZN(n15333) );
  AND2_X1 U11230 ( .A1(n14257), .A2(n12590), .ZN(n12591) );
  NOR2_X1 U11231 ( .A1(n15161), .A2(n9883), .ZN(n15138) );
  XNOR2_X1 U11232 ( .A(n12280), .B(n12279), .ZN(n13218) );
  AND2_X1 U11233 ( .A1(n15474), .A2(n15511), .ZN(n15499) );
  CLKBUF_X1 U11234 ( .A(n14297), .Z(n14298) );
  NAND2_X1 U11235 ( .A1(n9981), .A2(n9694), .ZN(n15492) );
  NAND2_X1 U11236 ( .A1(n9983), .A2(n11009), .ZN(n15534) );
  NAND2_X1 U11237 ( .A1(n9897), .A2(n15200), .ZN(n15512) );
  NOR2_X1 U11238 ( .A1(n14625), .A2(n14577), .ZN(n14599) );
  OAI21_X1 U11239 ( .B1(n15772), .B2(n11474), .A(n9929), .ZN(n11501) );
  NAND2_X1 U11240 ( .A1(n10091), .A2(n11005), .ZN(n16194) );
  NAND2_X1 U11241 ( .A1(n14637), .A2(n12575), .ZN(n14625) );
  NAND2_X1 U11242 ( .A1(n12575), .A2(n15883), .ZN(n14608) );
  NAND2_X1 U11243 ( .A1(n14636), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12575) );
  NAND2_X1 U11244 ( .A1(n9911), .A2(n15883), .ZN(n14636) );
  AND2_X1 U11245 ( .A1(n10125), .A2(n18134), .ZN(n11464) );
  NOR2_X1 U11246 ( .A1(n14938), .A2(n12664), .ZN(n12663) );
  AOI21_X1 U11247 ( .B1(n9991), .B2(n10313), .A(n10299), .ZN(n9990) );
  AND2_X1 U11248 ( .A1(n10816), .A2(n10823), .ZN(n9890) );
  OAI21_X1 U11249 ( .B1(n9999), .B2(n9998), .A(n9921), .ZN(n9991) );
  AOI21_X1 U11250 ( .B1(n15567), .B2(n9680), .A(n9688), .ZN(n9880) );
  XNOR2_X1 U11251 ( .A(n10789), .B(n10994), .ZN(n15558) );
  AND2_X1 U11252 ( .A1(n14355), .A2(n9837), .ZN(n14301) );
  OR2_X1 U11253 ( .A1(n13282), .A2(n10194), .ZN(n10192) );
  AOI21_X1 U11254 ( .B1(n10131), .B2(n12571), .A(n9787), .ZN(n9921) );
  NAND2_X1 U11255 ( .A1(n10764), .A2(n19043), .ZN(n10789) );
  NAND2_X1 U11256 ( .A1(n10993), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10998) );
  OR2_X1 U11257 ( .A1(n12573), .A2(n14668), .ZN(n10299) );
  AND2_X1 U11258 ( .A1(n10989), .A2(n10769), .ZN(n16218) );
  NOR2_X2 U11259 ( .A1(n14681), .A2(n12503), .ZN(n14788) );
  NAND2_X1 U11260 ( .A1(n13884), .A2(n13885), .ZN(n13963) );
  NOR2_X1 U11261 ( .A1(n18993), .A2(n13254), .ZN(n13269) );
  OAI211_X1 U11262 ( .C1(n12546), .C2(n11955), .A(n11845), .B(n11844), .ZN(
        n13980) );
  NAND2_X1 U11263 ( .A1(n11823), .A2(n11822), .ZN(n13885) );
  AND2_X1 U11264 ( .A1(n10761), .A2(n10760), .ZN(n10792) );
  AOI21_X1 U11265 ( .B1(n12548), .B2(n11971), .A(n11785), .ZN(n14125) );
  NAND2_X2 U11266 ( .A1(n13704), .A2(n10235), .ZN(n10237) );
  NAND2_X1 U11267 ( .A1(n11838), .A2(n11781), .ZN(n12548) );
  OR2_X1 U11268 ( .A1(n13272), .A2(n10899), .ZN(n10906) );
  OAI21_X1 U11269 ( .B1(n14089), .B2(n9924), .A(n12508), .ZN(n12531) );
  AOI21_X1 U11270 ( .B1(n12533), .B2(n11971), .A(n11834), .ZN(n13964) );
  NAND2_X1 U11271 ( .A1(n11824), .A2(n10004), .ZN(n14089) );
  AND4_X1 U11272 ( .A1(n10796), .A2(n10795), .A3(n10794), .A4(n10793), .ZN(
        n10809) );
  AND2_X1 U11273 ( .A1(n13749), .A2(n12917), .ZN(n13706) );
  XNOR2_X1 U11274 ( .A(n12549), .B(n11772), .ZN(n12559) );
  INV_X1 U11275 ( .A(n17822), .ZN(n17891) );
  AOI21_X1 U11276 ( .B1(n17614), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n18257), .ZN(n17729) );
  OAI21_X1 U11277 ( .B1(n11786), .B2(n10005), .A(n13868), .ZN(n10004) );
  NAND2_X1 U11278 ( .A1(n11813), .A2(n9845), .ZN(n12549) );
  INV_X1 U11279 ( .A(n17761), .ZN(n17809) );
  AND2_X1 U11280 ( .A1(n10689), .A2(n10688), .ZN(n10742) );
  XNOR2_X1 U11281 ( .A(n20162), .B(n12518), .ZN(n13330) );
  AND2_X1 U11282 ( .A1(n10690), .A2(n13648), .ZN(n10737) );
  AND3_X1 U11283 ( .A1(n11812), .A2(n9767), .A3(n13866), .ZN(n9845) );
  NOR2_X1 U11284 ( .A1(n18971), .A2(n14904), .ZN(n14891) );
  AND2_X1 U11285 ( .A1(n10690), .A2(n10688), .ZN(n19446) );
  AND2_X1 U11286 ( .A1(n10663), .A2(n10676), .ZN(n19613) );
  NAND2_X1 U11287 ( .A1(n10225), .A2(n10229), .ZN(n12916) );
  INV_X1 U11288 ( .A(n17897), .ZN(n17857) );
  AND2_X1 U11289 ( .A1(n12934), .A2(n9965), .ZN(n13647) );
  NAND2_X1 U11290 ( .A1(n9989), .A2(n11735), .ZN(n13866) );
  NOR2_X2 U11291 ( .A1(n15720), .A2(n9676), .ZN(n17806) );
  NAND2_X1 U11292 ( .A1(n20163), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n20162) );
  NAND2_X2 U11293 ( .A1(n11794), .A2(n11793), .ZN(n20283) );
  OAI21_X1 U11294 ( .B1(n12509), .B2(n9924), .A(n12511), .ZN(n20163) );
  NAND2_X1 U11295 ( .A1(n17804), .A2(n17805), .ZN(n17803) );
  NAND2_X1 U11296 ( .A1(n9896), .A2(n9895), .ZN(n9894) );
  INV_X1 U11297 ( .A(n11490), .ZN(n16511) );
  OR2_X1 U11298 ( .A1(n11264), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17697) );
  OR2_X1 U11299 ( .A1(n11807), .A2(n12056), .ZN(n11808) );
  NAND2_X1 U11300 ( .A1(n18906), .A2(n11490), .ZN(n17901) );
  NOR2_X1 U11301 ( .A1(n20353), .A2(n20214), .ZN(n20712) );
  OR2_X1 U11302 ( .A1(n20147), .A2(n9926), .ZN(n20148) );
  NOR2_X1 U11303 ( .A1(n20353), .A2(n20246), .ZN(n20756) );
  NOR2_X1 U11304 ( .A1(n20353), .A2(n20120), .ZN(n20732) );
  NAND2_X1 U11305 ( .A1(n11704), .A2(n11702), .ZN(n11698) );
  NOR2_X2 U11306 ( .A1(n10884), .A2(n10882), .ZN(n10881) );
  CLKBUF_X2 U11307 ( .A(n11803), .Z(n9664) );
  NAND2_X1 U11308 ( .A1(n10840), .A2(n9759), .ZN(n10884) );
  OR2_X1 U11309 ( .A1(n11699), .A2(n11700), .ZN(n11697) );
  OR2_X1 U11310 ( .A1(n10473), .A2(n10154), .ZN(n10840) );
  XNOR2_X1 U11311 ( .A(n11680), .B(n11630), .ZN(n11803) );
  NOR2_X2 U11312 ( .A1(n13352), .A2(n19956), .ZN(n11014) );
  OR2_X1 U11313 ( .A1(n16013), .A2(n14210), .ZN(n14476) );
  NAND2_X1 U11314 ( .A1(n9840), .A2(n12340), .ZN(n13715) );
  NOR2_X2 U11315 ( .A1(n19233), .A2(n19618), .ZN(n19234) );
  NOR2_X2 U11316 ( .A1(n19225), .A2(n19618), .ZN(n19226) );
  NOR2_X2 U11317 ( .A1(n19238), .A2(n19618), .ZN(n19239) );
  NAND2_X1 U11318 ( .A1(n10127), .A2(n11621), .ZN(n11680) );
  INV_X2 U11319 ( .A(n15036), .ZN(n14987) );
  OAI21_X1 U11320 ( .B1(n12339), .B2(n12337), .A(n12336), .ZN(n9840) );
  NAND2_X1 U11321 ( .A1(n10172), .A2(n10647), .ZN(n10650) );
  OR2_X1 U11322 ( .A1(n13889), .A2(n10085), .ZN(n16026) );
  NAND2_X1 U11323 ( .A1(n10601), .A2(n10600), .ZN(n10630) );
  OR2_X1 U11324 ( .A1(n12331), .A2(n12330), .ZN(n12339) );
  INV_X2 U11325 ( .A(n19031), .ZN(n9646) );
  NOR2_X2 U11326 ( .A1(n16510), .A2(n18914), .ZN(n17416) );
  AND2_X1 U11327 ( .A1(n10164), .A2(n10163), .ZN(n10161) );
  AND2_X1 U11328 ( .A1(n13578), .A2(n11141), .ZN(n16340) );
  AND2_X1 U11329 ( .A1(n16530), .A2(n17478), .ZN(n16526) );
  OR2_X1 U11330 ( .A1(n17390), .A2(n11255), .ZN(n11236) );
  NAND2_X1 U11331 ( .A1(n18241), .A2(n11402), .ZN(n11400) );
  NAND2_X1 U11332 ( .A1(n9995), .A2(n11602), .ZN(n9994) );
  NOR2_X1 U11333 ( .A1(n14178), .A2(n10591), .ZN(n15585) );
  BUF_X4 U11334 ( .A(n10631), .Z(n11113) );
  AND2_X1 U11335 ( .A1(n13594), .A2(n10621), .ZN(n10624) );
  XNOR2_X1 U11336 ( .A(n11255), .B(n11361), .ZN(n17835) );
  NOR2_X1 U11337 ( .A1(n15611), .A2(n11391), .ZN(n11402) );
  AND2_X2 U11338 ( .A1(n13207), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10631) );
  AND2_X1 U11339 ( .A1(n10592), .A2(n11126), .ZN(n13207) );
  INV_X1 U11340 ( .A(n11599), .ZN(n9996) );
  OR2_X1 U11341 ( .A1(n11623), .A2(n11615), .ZN(n13307) );
  AND2_X1 U11342 ( .A1(n13804), .A2(n11606), .ZN(n10309) );
  CLKBUF_X1 U11343 ( .A(n10965), .Z(n16343) );
  NOR2_X1 U11344 ( .A1(n17397), .A2(n9797), .ZN(n11252) );
  INV_X1 U11345 ( .A(n17418), .ZN(n18234) );
  AND2_X1 U11346 ( .A1(n11126), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10604) );
  NOR2_X1 U11347 ( .A1(n18266), .A2(n18245), .ZN(n11399) );
  NOR2_X1 U11348 ( .A1(n13448), .A2(n10591), .ZN(n10592) );
  AND2_X1 U11349 ( .A1(n13298), .A2(n11597), .ZN(n11599) );
  INV_X1 U11350 ( .A(n11454), .ZN(n18241) );
  AND2_X1 U11351 ( .A1(n13717), .A2(n12360), .ZN(n12439) );
  NOR2_X1 U11352 ( .A1(n12671), .A2(n10559), .ZN(n9889) );
  AND2_X1 U11353 ( .A1(n11554), .A2(n13725), .ZN(n11614) );
  OAI211_X1 U11354 ( .C1(n17015), .C2(n17179), .A(n11297), .B(n11296), .ZN(
        n11454) );
  INV_X1 U11355 ( .A(n10603), .ZN(n10591) );
  INV_X1 U11356 ( .A(n13617), .ZN(n11126) );
  INV_X1 U11357 ( .A(n11610), .ZN(n13319) );
  NAND2_X1 U11358 ( .A1(n11604), .A2(n14820), .ZN(n11605) );
  NAND2_X2 U11359 ( .A1(n10471), .A2(n10470), .ZN(n10947) );
  AOI211_X2 U11360 ( .C1(n17212), .C2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n11359), .B(n11358), .ZN(n18245) );
  INV_X1 U11361 ( .A(n13412), .ZN(n12360) );
  OAI211_X1 U11362 ( .C1(n17223), .C2(n15655), .A(n11317), .B(n11316), .ZN(
        n17418) );
  OAI211_X1 U11363 ( .C1(n17116), .C2(n17031), .A(n11185), .B(n11184), .ZN(
        n11364) );
  INV_X1 U11364 ( .A(n11612), .ZN(n13336) );
  NAND2_X1 U11365 ( .A1(n14820), .A2(n20227), .ZN(n12592) );
  NAND2_X2 U11366 ( .A1(n12670), .A2(n19220), .ZN(n13617) );
  AND2_X1 U11368 ( .A1(n16342), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9874) );
  OR2_X1 U11369 ( .A1(n11553), .A2(n11552), .ZN(n13725) );
  INV_X1 U11370 ( .A(n10554), .ZN(n10558) );
  OR2_X1 U11371 ( .A1(n11653), .A2(n11652), .ZN(n12569) );
  AND4_X1 U11372 ( .A1(n11563), .A2(n11562), .A3(n11561), .A4(n11560), .ZN(
        n11565) );
  AND4_X1 U11373 ( .A1(n11535), .A2(n11534), .A3(n11533), .A4(n11532), .ZN(
        n11542) );
  INV_X2 U11374 ( .A(U212), .ZN(n16446) );
  OR2_X2 U11375 ( .A1(n16459), .A2(n16408), .ZN(n16461) );
  AND4_X1 U11376 ( .A1(n11582), .A2(n11583), .A3(n11585), .A4(n11584), .ZN(
        n11586) );
  AND2_X1 U11377 ( .A1(n10065), .A2(n10315), .ZN(n10064) );
  OR2_X2 U11378 ( .A1(n11530), .A2(n11529), .ZN(n11600) );
  OAI21_X1 U11379 ( .B1(n10529), .B2(n10528), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10536) );
  NAND3_X1 U11380 ( .A1(n10549), .A2(n10548), .A3(n10547), .ZN(n10550) );
  AND3_X1 U11381 ( .A1(n11519), .A2(n11518), .A3(n11506), .ZN(n9959) );
  AND4_X1 U11382 ( .A1(n9961), .A2(n11520), .A3(n11509), .A4(n11517), .ZN(
        n9960) );
  AND3_X1 U11383 ( .A1(n11579), .A2(n11580), .A3(n11581), .ZN(n10065) );
  AND4_X1 U11384 ( .A1(n11539), .A2(n11538), .A3(n11537), .A4(n11536), .ZN(
        n11541) );
  BUF_X2 U11385 ( .A(n12261), .Z(n9670) );
  INV_X2 U11386 ( .A(n17199), .ZN(n17149) );
  BUF_X2 U11387 ( .A(n12089), .Z(n9667) );
  AND2_X1 U11388 ( .A1(n9811), .A2(n9810), .ZN(n11521) );
  AND2_X1 U11389 ( .A1(n10364), .A2(n10365), .ZN(n10011) );
  AND2_X1 U11390 ( .A1(n10371), .A2(n10370), .ZN(n10372) );
  AND4_X1 U11391 ( .A1(n10344), .A2(n10343), .A3(n10342), .A4(n10341), .ZN(
        n10345) );
  AND3_X1 U11392 ( .A1(n10545), .A2(n10517), .A3(n10544), .ZN(n10549) );
  AND4_X1 U11393 ( .A1(n10349), .A2(n10348), .A3(n10347), .A4(n10346), .ZN(
        n10350) );
  INV_X2 U11394 ( .A(n20815), .ZN(n20838) );
  INV_X1 U11395 ( .A(n18851), .ZN(n18759) );
  CLKBUF_X3 U11396 ( .A(n11571), .Z(n9672) );
  INV_X2 U11397 ( .A(n18217), .ZN(n9647) );
  INV_X2 U11398 ( .A(n16495), .ZN(U215) );
  NOR2_X1 U11399 ( .A1(n18865), .A2(n17896), .ZN(n18903) );
  NAND2_X1 U11400 ( .A1(n9803), .A2(n11153), .ZN(n17223) );
  NAND2_X2 U11401 ( .A1(n19974), .A2(n19839), .ZN(n19886) );
  INV_X1 U11402 ( .A(n17210), .ZN(n17199) );
  INV_X1 U11403 ( .A(n19897), .ZN(n19823) );
  CLKBUF_X1 U11404 ( .A(n13525), .Z(n19217) );
  AND2_X2 U11405 ( .A1(n10546), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10380) );
  INV_X2 U11406 ( .A(n16499), .ZN(n16501) );
  INV_X2 U11407 ( .A(n18896), .ZN(n18830) );
  OR2_X1 U11408 ( .A1(n11155), .A2(n11154), .ZN(n9746) );
  OR2_X1 U11409 ( .A1(n11154), .A2(n18690), .ZN(n17188) );
  INV_X1 U11410 ( .A(n9644), .ZN(n17135) );
  OAI21_X1 U11411 ( .B1(n13240), .B2(n13239), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13525) );
  NAND2_X1 U11412 ( .A1(n10247), .A2(n13805), .ZN(n12186) );
  INV_X2 U11413 ( .A(n12139), .ZN(n11760) );
  AND2_X2 U11414 ( .A1(n11504), .A2(n13674), .ZN(n11846) );
  INV_X1 U11415 ( .A(n12139), .ZN(n9671) );
  NAND4_X1 U11416 ( .A1(n13807), .A2(n13576), .A3(n9913), .A4(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12139) );
  AND2_X1 U11417 ( .A1(n13807), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11504) );
  AND3_X1 U11418 ( .A1(n11687), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11503) );
  NAND2_X1 U11419 ( .A1(n13805), .A2(n11516), .ZN(n12184) );
  AND2_X1 U11420 ( .A1(n9913), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13806) );
  AND2_X1 U11421 ( .A1(n10317), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10328) );
  AND2_X2 U11422 ( .A1(n10321), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10542) );
  NOR2_X1 U11423 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10321) );
  INV_X1 U11424 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10639) );
  NOR2_X1 U11425 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11516) );
  AND2_X1 U11426 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11512) );
  NOR2_X1 U11427 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11511) );
  AND2_X2 U11428 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13810) );
  AND2_X1 U11429 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15582) );
  AOI21_X1 U11430 ( .B1(n15883), .B2(n14569), .A(n14568), .ZN(n14570) );
  AND2_X1 U11431 ( .A1(n11507), .A2(n11508), .ZN(n9961) );
  NOR2_X2 U11432 ( .A1(n14297), .A2(n14299), .ZN(n14282) );
  NAND2_X2 U11433 ( .A1(n11698), .A2(n11697), .ZN(n9915) );
  AOI21_X1 U11434 ( .B1(n14705), .B2(n20156), .A(n13225), .ZN(n13226) );
  XNOR2_X1 U11435 ( .A(n13222), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14705) );
  NOR2_X4 U11436 ( .A1(n16896), .A2(n11154), .ZN(n11217) );
  OAI22_X2 U11437 ( .A1(n10915), .A2(n15179), .B1(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n10914), .ZN(n15162) );
  NAND2_X1 U11438 ( .A1(n10178), .A2(n10177), .ZN(n9655) );
  OAI21_X2 U11439 ( .B1(n15452), .B2(n15453), .A(n15211), .ZN(n16115) );
  OAI21_X2 U11440 ( .B1(n15209), .B2(n15208), .A(n15207), .ZN(n15452) );
  OAI22_X2 U11441 ( .A1(n14003), .A2(n14002), .B1(n14056), .B2(n14014), .ZN(
        n15557) );
  OR2_X2 U11442 ( .A1(n12622), .A2(n10196), .ZN(n12621) );
  NOR2_X2 U11443 ( .A1(n15153), .A2(n14843), .ZN(n14842) );
  NAND2_X2 U11444 ( .A1(n9992), .A2(n9728), .ZN(n12594) );
  INV_X1 U11445 ( .A(n13803), .ZN(n9658) );
  AND2_X1 U11446 ( .A1(n13672), .A2(n13807), .ZN(n11588) );
  AND2_X1 U11447 ( .A1(n11513), .A2(n11512), .ZN(n11531) );
  INV_X1 U11448 ( .A(n13412), .ZN(n9662) );
  CLKBUF_X1 U11449 ( .A(n17158), .Z(n9663) );
  INV_X1 U11450 ( .A(n11186), .ZN(n17158) );
  INV_X1 U11451 ( .A(n10947), .ZN(n9665) );
  INV_X1 U11452 ( .A(n12141), .ZN(n12089) );
  AND2_X1 U11453 ( .A1(n11511), .A2(n13810), .ZN(n11879) );
  INV_X4 U11455 ( .A(n12186), .ZN(n12160) );
  INV_X2 U11456 ( .A(n11600), .ZN(n11606) );
  INV_X1 U11457 ( .A(n12139), .ZN(n12260) );
  NOR2_X2 U11458 ( .A1(n12640), .A2(n12642), .ZN(n12639) );
  NAND2_X1 U11459 ( .A1(n13806), .A2(n11515), .ZN(n12188) );
  AND2_X4 U11460 ( .A1(n11503), .A2(n13807), .ZN(n11543) );
  NOR2_X2 U11461 ( .A1(n12637), .A2(n15240), .ZN(n12636) );
  NOR2_X2 U11462 ( .A1(n14124), .A2(n14147), .ZN(n14148) );
  NOR2_X2 U11463 ( .A1(n14589), .A2(n9919), .ZN(n14568) );
  NOR2_X4 U11464 ( .A1(n9717), .A2(n16150), .ZN(n12646) );
  OR2_X2 U11465 ( .A1(n12648), .A2(n10179), .ZN(n9717) );
  NOR2_X2 U11466 ( .A1(n12643), .A2(n18960), .ZN(n12645) );
  XNOR2_X2 U11467 ( .A(n11786), .B(n11812), .ZN(n12521) );
  NAND2_X2 U11468 ( .A1(n11794), .A2(n11686), .ZN(n11786) );
  NOR2_X2 U11469 ( .A1(n12634), .A2(n15215), .ZN(n12633) );
  NOR2_X2 U11470 ( .A1(n12631), .A2(n15188), .ZN(n12629) );
  NOR2_X2 U11471 ( .A1(n12650), .A2(n15264), .ZN(n12652) );
  NOR2_X2 U11472 ( .A1(n12627), .A2(n14863), .ZN(n12625) );
  INV_X4 U11473 ( .A(n14079), .ZN(n18993) );
  NOR2_X1 U11474 ( .A1(n20147), .A2(n9926), .ZN(n9678) );
  NOR2_X1 U11475 ( .A1(n11236), .A2(n17387), .ZN(n11463) );
  NOR2_X1 U11476 ( .A1(n11786), .A2(n9844), .ZN(n11759) );
  INV_X1 U11477 ( .A(n11897), .ZN(n10251) );
  NAND2_X1 U11478 ( .A1(n10641), .A2(n10640), .ZN(n10658) );
  CLKBUF_X1 U11479 ( .A(n9713), .Z(n17015) );
  NAND2_X1 U11480 ( .A1(n9800), .A2(n9799), .ZN(n11275) );
  INV_X1 U11481 ( .A(n11274), .ZN(n9800) );
  AND2_X1 U11482 ( .A1(n17805), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10126) );
  AOI21_X1 U11483 ( .B1(n11452), .B2(n11451), .A(n11450), .ZN(n18727) );
  NOR2_X1 U11484 ( .A1(n13586), .A2(n19220), .ZN(n9873) );
  NAND2_X1 U11485 ( .A1(n19584), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n9861) );
  NAND2_X1 U11486 ( .A1(n19525), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n9862) );
  NAND2_X1 U11487 ( .A1(n19752), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n9863) );
  NAND2_X1 U11488 ( .A1(n19654), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n9864) );
  NAND2_X1 U11489 ( .A1(n13571), .A2(n20227), .ZN(n9995) );
  NOR2_X1 U11490 ( .A1(n12670), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12672) );
  NAND2_X1 U11491 ( .A1(n10264), .A2(n14283), .ZN(n10263) );
  INV_X1 U11492 ( .A(n14273), .ZN(n10264) );
  AND2_X1 U11493 ( .A1(n10252), .A2(n10251), .ZN(n10250) );
  INV_X1 U11494 ( .A(n13963), .ZN(n9826) );
  XNOR2_X1 U11495 ( .A(n11824), .B(n11825), .ZN(n12533) );
  NOR2_X1 U11496 ( .A1(n11576), .A2(n11773), .ZN(n11971) );
  NAND2_X1 U11497 ( .A1(n9985), .A2(n12570), .ZN(n10131) );
  NAND2_X1 U11498 ( .A1(n9988), .A2(n9986), .ZN(n9985) );
  OR2_X1 U11499 ( .A1(n15883), .A2(n16019), .ZN(n12570) );
  NAND2_X1 U11500 ( .A1(n9917), .A2(n14198), .ZN(n9988) );
  NAND2_X1 U11501 ( .A1(n13307), .A2(n13571), .ZN(n11629) );
  NAND2_X1 U11502 ( .A1(n13800), .A2(n16055), .ZN(n9989) );
  INV_X1 U11503 ( .A(n15159), .ZN(n10189) );
  AND2_X1 U11504 ( .A1(n10157), .A2(n10873), .ZN(n10156) );
  INV_X1 U11505 ( .A(n10854), .ZN(n10153) );
  AND2_X1 U11506 ( .A1(n10472), .A2(n10165), .ZN(n10164) );
  INV_X1 U11507 ( .A(n10762), .ZN(n10165) );
  AND2_X1 U11508 ( .A1(n9756), .A2(n16161), .ZN(n10291) );
  AND2_X1 U11509 ( .A1(n10294), .A2(n10830), .ZN(n10293) );
  INV_X1 U11510 ( .A(n15530), .ZN(n10294) );
  OR3_X1 U11511 ( .A1(n11008), .A2(n10899), .A3(n11007), .ZN(n11009) );
  OR2_X1 U11512 ( .A1(n11008), .A2(n10899), .ZN(n11006) );
  OAI21_X1 U11513 ( .B1(n10991), .B2(n10016), .A(n11002), .ZN(n10015) );
  INV_X1 U11514 ( .A(n10792), .ZN(n10016) );
  NAND2_X1 U11515 ( .A1(n10657), .A2(n10659), .ZN(n10017) );
  INV_X1 U11516 ( .A(n10657), .ZN(n10018) );
  AND2_X1 U11517 ( .A1(n11019), .A2(n10652), .ZN(n10231) );
  NAND2_X1 U11518 ( .A1(n12672), .A2(n12668), .ZN(n12842) );
  CLKBUF_X2 U11519 ( .A(n12712), .Z(n12871) );
  NOR2_X1 U11520 ( .A1(n12697), .A2(n12696), .ZN(n12702) );
  NAND2_X1 U11521 ( .A1(n9962), .A2(n12923), .ZN(n12934) );
  XNOR2_X1 U11522 ( .A(n11236), .B(n9928), .ZN(n11256) );
  INV_X1 U11523 ( .A(n17387), .ZN(n9928) );
  NAND2_X1 U11524 ( .A1(n14217), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13928) );
  INV_X1 U11525 ( .A(n10316), .ZN(n11987) );
  AND2_X1 U11526 ( .A1(n11773), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12277) );
  AND2_X1 U11527 ( .A1(n14625), .A2(n10061), .ZN(n14578) );
  NAND2_X1 U11528 ( .A1(n15883), .A2(n14718), .ZN(n10061) );
  AND2_X1 U11529 ( .A1(n13312), .A2(n19975), .ZN(n13338) );
  NAND2_X1 U11530 ( .A1(n13715), .A2(n9757), .ZN(n13310) );
  NOR2_X1 U11531 ( .A1(n9818), .A2(n9817), .ZN(n9816) );
  INV_X1 U11532 ( .A(n11685), .ZN(n9817) );
  INV_X1 U11533 ( .A(n9819), .ZN(n9818) );
  OR2_X1 U11534 ( .A1(n15070), .A2(n15071), .ZN(n15068) );
  NAND2_X1 U11535 ( .A1(n12905), .A2(n19931), .ZN(n12928) );
  AND2_X1 U11536 ( .A1(n19904), .A2(n19933), .ZN(n19415) );
  NAND2_X1 U11537 ( .A1(n11450), .A2(n11442), .ZN(n18725) );
  NOR3_X1 U11538 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n11155), .ZN(n17206) );
  INV_X1 U11539 ( .A(n17737), .ZN(n17805) );
  NAND2_X1 U11540 ( .A1(n10121), .A2(n17837), .ZN(n10120) );
  INV_X1 U11541 ( .A(n17835), .ZN(n10121) );
  NAND2_X1 U11542 ( .A1(n17835), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10119) );
  XNOR2_X1 U11543 ( .A(n11256), .B(n18150), .ZN(n17824) );
  NOR2_X1 U11544 ( .A1(n18752), .A2(n18749), .ZN(n18901) );
  AOI21_X1 U11545 ( .B1(n14747), .B2(n20047), .A(n9832), .ZN(n9831) );
  OAI21_X1 U11546 ( .B1(n20053), .B2(n14573), .A(n9833), .ZN(n9832) );
  NAND2_X1 U11547 ( .A1(n15848), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n9833) );
  AND2_X1 U11548 ( .A1(n12666), .A2(n12665), .ZN(n15301) );
  OAI211_X1 U11549 ( .C1(n17015), .C2(n18580), .A(n11165), .B(n11164), .ZN(
        n17381) );
  AOI21_X1 U11550 ( .B1(n11464), .B2(n11463), .A(n11462), .ZN(n11465) );
  NAND2_X1 U11551 ( .A1(n10559), .A2(n10558), .ZN(n10560) );
  NAND2_X1 U11552 ( .A1(n12911), .A2(n13379), .ZN(n10561) );
  INV_X1 U11553 ( .A(n12454), .ZN(n9922) );
  NAND2_X1 U11554 ( .A1(n10406), .A2(n10405), .ZN(n10419) );
  NAND2_X1 U11555 ( .A1(n10026), .A2(n10025), .ZN(n10024) );
  NAND2_X1 U11556 ( .A1(n10674), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10026) );
  NAND2_X1 U11557 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10025) );
  NAND2_X1 U11558 ( .A1(n10675), .A2(n10020), .ZN(n10019) );
  NAND2_X1 U11559 ( .A1(n10022), .A2(n10021), .ZN(n10020) );
  NAND2_X1 U11560 ( .A1(n10674), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10022) );
  NAND2_X1 U11561 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10021) );
  AOI22_X1 U11562 ( .A1(n13066), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10365) );
  AND2_X1 U11563 ( .A1(n10363), .A2(n10517), .ZN(n10367) );
  AOI21_X1 U11564 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n18714), .A(
        n11419), .ZN(n11420) );
  NOR2_X1 U11565 ( .A1(n11427), .A2(n11426), .ZN(n11419) );
  OR2_X1 U11566 ( .A1(n12291), .A2(n12290), .ZN(n12298) );
  NAND2_X1 U11567 ( .A1(n13806), .A2(n13810), .ZN(n12190) );
  AND2_X1 U11568 ( .A1(n13576), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10247) );
  AND2_X1 U11569 ( .A1(n11612), .A2(n11600), .ZN(n11610) );
  NOR2_X1 U11570 ( .A1(n11687), .A2(n16055), .ZN(n9908) );
  NAND2_X1 U11571 ( .A1(n11618), .A2(n9908), .ZN(n9906) );
  NAND2_X1 U11572 ( .A1(n11510), .A2(n13806), .ZN(n12141) );
  NOR2_X1 U11573 ( .A1(n11514), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11510) );
  INV_X1 U11574 ( .A(n12710), .ZN(n10810) );
  OAI22_X1 U11575 ( .A1(n10419), .A2(n10418), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n10517), .ZN(n10954) );
  AND3_X1 U11577 ( .A1(n10573), .A2(n12911), .A3(n9873), .ZN(n9872) );
  INV_X1 U11578 ( .A(n10173), .ZN(n10172) );
  OAI21_X1 U11579 ( .B1(n10635), .B2(n10175), .A(n10174), .ZN(n10173) );
  AND2_X1 U11580 ( .A1(n10646), .A2(n10645), .ZN(n10648) );
  NAND3_X1 U11581 ( .A1(n12668), .A2(n10552), .A3(n9887), .ZN(n10965) );
  NAND2_X1 U11582 ( .A1(n9888), .A2(n9885), .ZN(n13206) );
  INV_X1 U11583 ( .A(n10593), .ZN(n9888) );
  NAND2_X1 U11584 ( .A1(n10965), .A2(n9886), .ZN(n9885) );
  AND2_X1 U11585 ( .A1(n12670), .A2(n19237), .ZN(n9886) );
  NAND2_X1 U11586 ( .A1(n10231), .A2(n9704), .ZN(n10227) );
  NAND2_X1 U11587 ( .A1(n12912), .A2(n12911), .ZN(n12927) );
  NOR2_X1 U11588 ( .A1(n13380), .A2(n9877), .ZN(n12912) );
  NAND2_X1 U11589 ( .A1(n10688), .A2(n13613), .ZN(n10677) );
  NAND2_X1 U11590 ( .A1(n11238), .A2(n17409), .ZN(n9797) );
  NAND2_X1 U11591 ( .A1(n10083), .A2(n14335), .ZN(n10082) );
  INV_X1 U11592 ( .A(n14440), .ZN(n10083) );
  NAND2_X1 U11593 ( .A1(n12130), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12174) );
  NAND2_X1 U11594 ( .A1(n10270), .A2(n14338), .ZN(n10269) );
  INV_X1 U11595 ( .A(n10271), .ZN(n10270) );
  NOR2_X1 U11596 ( .A1(n10256), .A2(n10255), .ZN(n10254) );
  INV_X1 U11597 ( .A(n14459), .ZN(n10255) );
  OR2_X1 U11598 ( .A1(n13725), .A2(n11773), .ZN(n10316) );
  AND2_X1 U11599 ( .A1(n11815), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11829) );
  OR2_X1 U11600 ( .A1(n12512), .A2(n20220), .ZN(n9912) );
  AND2_X1 U11601 ( .A1(n14667), .A2(n14689), .ZN(n14805) );
  NAND2_X1 U11602 ( .A1(n10076), .A2(n14464), .ZN(n10075) );
  INV_X1 U11603 ( .A(n14475), .ZN(n10076) );
  NAND2_X1 U11604 ( .A1(n15893), .A2(n10132), .ZN(n9999) );
  NOR2_X1 U11605 ( .A1(n10133), .A2(n10134), .ZN(n10132) );
  NOR2_X1 U11606 ( .A1(n10313), .A2(n9754), .ZN(n9917) );
  NAND2_X1 U11607 ( .A1(n13412), .A2(n13717), .ZN(n12443) );
  NAND2_X1 U11608 ( .A1(n9923), .A2(n13553), .ZN(n13296) );
  AND2_X1 U11609 ( .A1(n11812), .A2(n13866), .ZN(n10248) );
  INV_X1 U11610 ( .A(n11605), .ZN(n13804) );
  INV_X1 U11611 ( .A(n12509), .ZN(n14090) );
  NAND2_X1 U11612 ( .A1(n10840), .A2(n10847), .ZN(n10855) );
  NOR2_X1 U11613 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n10838), .ZN(n10473) );
  NOR2_X1 U11614 ( .A1(n10831), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10834) );
  INV_X1 U11615 ( .A(n10763), .ZN(n10162) );
  NAND2_X1 U11616 ( .A1(n10637), .A2(n10636), .ZN(n9866) );
  NOR2_X1 U11617 ( .A1(n12937), .A2(n10238), .ZN(n10235) );
  INV_X1 U11618 ( .A(n12935), .ZN(n10238) );
  AND3_X1 U11619 ( .A1(n10218), .A2(n9778), .A3(n10221), .ZN(n9691) );
  INV_X1 U11620 ( .A(n14968), .ZN(n10222) );
  AND2_X1 U11621 ( .A1(n10232), .A2(n14986), .ZN(n9970) );
  AND2_X1 U11622 ( .A1(n10234), .A2(n10233), .ZN(n10232) );
  INV_X1 U11623 ( .A(n14991), .ZN(n10233) );
  NOR2_X1 U11624 ( .A1(n10438), .A2(n10437), .ZN(n12676) );
  INV_X1 U11625 ( .A(n13258), .ZN(n10197) );
  AND2_X1 U11626 ( .A1(n14893), .A2(n10199), .ZN(n10198) );
  INV_X1 U11627 ( .A(n14879), .ZN(n10199) );
  NAND2_X1 U11628 ( .A1(n10288), .A2(n10302), .ZN(n10287) );
  OR2_X1 U11629 ( .A1(n15144), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10302) );
  INV_X1 U11630 ( .A(n10928), .ZN(n10288) );
  INV_X1 U11631 ( .A(n15081), .ZN(n10045) );
  INV_X1 U11632 ( .A(n10051), .ZN(n10050) );
  NAND2_X1 U11633 ( .A1(n9735), .A2(n11002), .ZN(n11008) );
  OR2_X1 U11634 ( .A1(n10661), .A2(n10660), .ZN(n10665) );
  NAND2_X1 U11635 ( .A1(n10660), .A2(n10661), .ZN(n10662) );
  CLKBUF_X1 U11636 ( .A(n13207), .Z(n15584) );
  INV_X1 U11637 ( .A(n10677), .ZN(n10676) );
  AOI22_X1 U11638 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13047), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10544) );
  AND3_X1 U11639 ( .A1(n10553), .A2(n19237), .A3(n19242), .ZN(n10552) );
  INV_X1 U11640 ( .A(n11151), .ZN(n9803) );
  NAND2_X1 U11641 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18887), .ZN(
        n11155) );
  NAND2_X1 U11642 ( .A1(n18860), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11154) );
  INV_X1 U11643 ( .A(n11222), .ZN(n9936) );
  AOI21_X1 U11644 ( .B1(n11202), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n9938), .ZN(n9937) );
  INV_X1 U11645 ( .A(n11267), .ZN(n9796) );
  NOR2_X1 U11646 ( .A1(n17697), .A2(n9941), .ZN(n11262) );
  NAND2_X1 U11647 ( .A1(n17878), .A2(n11248), .ZN(n11249) );
  XNOR2_X1 U11648 ( .A(n17409), .B(n11238), .ZN(n11239) );
  OAI21_X1 U11649 ( .B1(n18245), .B2(n11409), .A(n11436), .ZN(n11411) );
  AND2_X1 U11650 ( .A1(n9859), .A2(n15707), .ZN(n16525) );
  INV_X1 U11651 ( .A(n18694), .ZN(n9859) );
  INV_X1 U11652 ( .A(n18904), .ZN(n17415) );
  NAND2_X1 U11653 ( .A1(n9996), .A2(n9723), .ZN(n9993) );
  NOR2_X1 U11654 ( .A1(n14304), .A2(n21010), .ZN(n9837) );
  AND3_X1 U11655 ( .A1(n14104), .A2(n11612), .A3(n11576), .ZN(n13716) );
  NAND2_X1 U11656 ( .A1(n9761), .A2(n9828), .ZN(n9827) );
  INV_X1 U11657 ( .A(n14299), .ZN(n9828) );
  NAND2_X1 U11658 ( .A1(n12224), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12274) );
  INV_X1 U11659 ( .A(n15921), .ZN(n10146) );
  OR2_X1 U11660 ( .A1(n10251), .A2(n10252), .ZN(n10249) );
  NAND2_X1 U11661 ( .A1(n11814), .A2(n11971), .ZN(n11823) );
  OR2_X1 U11662 ( .A1(n13715), .A2(n15762), .ZN(n13650) );
  AND2_X1 U11663 ( .A1(n9692), .A2(n14737), .ZN(n9848) );
  AND2_X1 U11664 ( .A1(n14287), .A2(n14269), .ZN(n14271) );
  INV_X1 U11665 ( .A(n12565), .ZN(n10134) );
  INV_X1 U11666 ( .A(n9988), .ZN(n10133) );
  INV_X1 U11667 ( .A(n9917), .ZN(n14194) );
  INV_X1 U11668 ( .A(n10089), .ZN(n10086) );
  XNOR2_X1 U11669 ( .A(n12540), .B(n13915), .ZN(n13907) );
  NAND2_X1 U11670 ( .A1(n13907), .A2(n13908), .ZN(n13906) );
  NAND2_X1 U11671 ( .A1(n11691), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10127) );
  OAI211_X1 U11672 ( .C1(n11629), .C2(n20220), .A(n11628), .B(n11627), .ZN(
        n11679) );
  NOR2_X1 U11673 ( .A1(n11625), .A2(n9916), .ZN(n11628) );
  OAI211_X1 U11674 ( .C1(n12315), .C2(n20218), .A(n11658), .B(n11657), .ZN(
        n11801) );
  NOR2_X1 U11675 ( .A1(n11674), .A2(n9747), .ZN(n9820) );
  NAND2_X1 U11676 ( .A1(n20256), .A2(n11704), .ZN(n20455) );
  NAND2_X1 U11677 ( .A1(n12521), .A2(n13868), .ZN(n20426) );
  INV_X1 U11678 ( .A(n20554), .ZN(n20509) );
  OR2_X1 U11679 ( .A1(n20283), .A2(n12509), .ZN(n20641) );
  NOR2_X1 U11680 ( .A1(n20514), .A2(n20353), .ZN(n20678) );
  NAND2_X1 U11681 ( .A1(n16055), .A2(n14103), .ZN(n20353) );
  AND2_X1 U11682 ( .A1(n11136), .A2(n10960), .ZN(n16333) );
  NOR2_X1 U11683 ( .A1(n10185), .A2(n18993), .ZN(n10184) );
  INV_X1 U11684 ( .A(n10187), .ZN(n10185) );
  NOR2_X1 U11685 ( .A1(n10191), .A2(n18993), .ZN(n10190) );
  INV_X1 U11686 ( .A(n10193), .ZN(n10191) );
  OR2_X1 U11687 ( .A1(n10825), .A2(n19251), .ZN(n10924) );
  NAND2_X1 U11688 ( .A1(n10881), .A2(n9760), .ZN(n10871) );
  INV_X1 U11689 ( .A(n10869), .ZN(n10155) );
  NAND2_X1 U11690 ( .A1(n10834), .A2(n14142), .ZN(n10838) );
  AND2_X1 U11691 ( .A1(n19251), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10824) );
  AOI21_X1 U11692 ( .B1(n10034), .B2(n10037), .A(n9762), .ZN(n13989) );
  NOR2_X1 U11693 ( .A1(n10035), .A2(n10040), .ZN(n10034) );
  NAND2_X1 U11694 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10177) );
  AND2_X1 U11695 ( .A1(n16333), .A2(n19819), .ZN(n13348) );
  NOR2_X1 U11696 ( .A1(n13860), .A2(n9966), .ZN(n14164) );
  NAND2_X1 U11697 ( .A1(n9967), .A2(n14167), .ZN(n9966) );
  INV_X1 U11698 ( .A(n9968), .ZN(n9967) );
  NAND2_X1 U11699 ( .A1(n13878), .A2(n13900), .ZN(n10224) );
  NAND2_X1 U11700 ( .A1(n10243), .A2(n10242), .ZN(n10241) );
  INV_X1 U11701 ( .A(n14950), .ZN(n10242) );
  NAND2_X1 U11702 ( .A1(n10032), .A2(n10031), .ZN(n10035) );
  INV_X1 U11703 ( .A(n12703), .ZN(n10032) );
  AND2_X1 U11704 ( .A1(n13943), .A2(n10036), .ZN(n10031) );
  INV_X1 U11705 ( .A(n13946), .ZN(n10036) );
  NAND4_X1 U11706 ( .A1(n13465), .A2(n10553), .A3(n10573), .A4(n12904), .ZN(
        n13448) );
  INV_X1 U11707 ( .A(n14170), .ZN(n10206) );
  XNOR2_X1 U11708 ( .A(n9711), .B(n14835), .ZN(n15282) );
  NAND2_X1 U11709 ( .A1(n9884), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9883) );
  NAND2_X1 U11710 ( .A1(n9882), .A2(n9884), .ZN(n15150) );
  INV_X1 U11711 ( .A(n15144), .ZN(n9892) );
  AND2_X1 U11712 ( .A1(n9710), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10104) );
  NAND2_X1 U11713 ( .A1(n15534), .A2(n9710), .ZN(n15178) );
  AND2_X1 U11714 ( .A1(n15534), .A2(n10105), .ZN(n15193) );
  NAND2_X1 U11715 ( .A1(n9901), .A2(n9898), .ZN(n15186) );
  INV_X1 U11716 ( .A(n9899), .ZN(n9898) );
  NAND2_X1 U11717 ( .A1(n16153), .A2(n9902), .ZN(n9901) );
  OAI21_X1 U11718 ( .B1(n9687), .B2(n9900), .A(n10282), .ZN(n9899) );
  NAND2_X1 U11719 ( .A1(n15534), .A2(n11013), .ZN(n15398) );
  INV_X1 U11720 ( .A(n15512), .ZN(n10858) );
  AND2_X1 U11721 ( .A1(n15492), .A2(n15426), .ZN(n16121) );
  NAND2_X1 U11722 ( .A1(n14171), .A2(n15037), .ZN(n15038) );
  AND2_X1 U11723 ( .A1(n11057), .A2(n11056), .ZN(n15029) );
  NOR2_X1 U11724 ( .A1(n15038), .A2(n15029), .ZN(n15030) );
  INV_X1 U11725 ( .A(n16176), .ZN(n10292) );
  NAND2_X1 U11726 ( .A1(n15570), .A2(n10998), .ZN(n10999) );
  INV_X1 U11727 ( .A(n10231), .ZN(n9895) );
  NAND2_X1 U11728 ( .A1(n10644), .A2(n10643), .ZN(n9896) );
  INV_X1 U11729 ( .A(n15579), .ZN(n13409) );
  AND2_X1 U11730 ( .A1(n10665), .A2(n10662), .ZN(n19063) );
  AOI21_X1 U11731 ( .B1(n19193), .B2(n12931), .A(n12930), .ZN(n13468) );
  NAND2_X1 U11732 ( .A1(n13469), .A2(n13468), .ZN(n13470) );
  NAND2_X1 U11733 ( .A1(n19519), .A2(n19479), .ZN(n19652) );
  AND2_X1 U11734 ( .A1(n11143), .A2(n9877), .ZN(n19761) );
  OR2_X1 U11735 ( .A1(n16362), .A2(n11142), .ZN(n11143) );
  INV_X1 U11736 ( .A(n19761), .ZN(n19618) );
  NOR2_X2 U11737 ( .A1(n19219), .A2(n19218), .ZN(n19258) );
  NOR2_X2 U11738 ( .A1(n19217), .A2(n19218), .ZN(n19259) );
  AOI21_X1 U11739 ( .B1(n11202), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n10110), .ZN(n10109) );
  INV_X1 U11740 ( .A(n11244), .ZN(n10111) );
  OR3_X1 U11741 ( .A1(n17345), .A2(n15611), .A3(n15610), .ZN(n15612) );
  OAI21_X1 U11742 ( .B1(n16525), .B2(n16526), .A(n9858), .ZN(n15799) );
  AND2_X1 U11743 ( .A1(n18725), .A2(n18907), .ZN(n9858) );
  NAND2_X1 U11744 ( .A1(n17672), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17651) );
  INV_X1 U11745 ( .A(n17730), .ZN(n9947) );
  NOR2_X1 U11746 ( .A1(n17821), .A2(n17827), .ZN(n17794) );
  OR2_X1 U11747 ( .A1(n17843), .A2(n17842), .ZN(n17821) );
  NOR2_X1 U11748 ( .A1(n17574), .A2(n11271), .ZN(n11272) );
  NAND2_X1 U11749 ( .A1(n10114), .A2(n9792), .ZN(n17823) );
  AND2_X1 U11750 ( .A1(n10113), .A2(n17824), .ZN(n9792) );
  NAND2_X1 U11751 ( .A1(n10118), .A2(n10119), .ZN(n10113) );
  OR2_X1 U11752 ( .A1(n17840), .A2(n17841), .ZN(n9806) );
  NAND2_X1 U11753 ( .A1(n17849), .A2(n11254), .ZN(n17836) );
  INV_X1 U11754 ( .A(n15800), .ZN(n17895) );
  INV_X1 U11755 ( .A(n15762), .ZN(n19975) );
  OR2_X1 U11756 ( .A1(n14259), .A2(n20963), .ZN(n9834) );
  AND2_X1 U11757 ( .A1(n14217), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20048) );
  AND2_X1 U11758 ( .A1(n14217), .A2(n12356), .ZN(n20041) );
  INV_X1 U11759 ( .A(n20049), .ZN(n20040) );
  AND2_X1 U11760 ( .A1(n12462), .A2(n12452), .ZN(n20047) );
  XOR2_X1 U11761 ( .A(n12450), .B(n12449), .Z(n14706) );
  NAND3_X1 U11762 ( .A1(n10068), .A2(n10067), .A3(n10069), .ZN(n12449) );
  NAND2_X1 U11763 ( .A1(n10071), .A2(n13412), .ZN(n10069) );
  XNOR2_X1 U11764 ( .A(n9641), .B(n12479), .ZN(n14241) );
  XNOR2_X1 U11765 ( .A(n14583), .B(n14582), .ZN(n14755) );
  NAND2_X1 U11766 ( .A1(n14581), .A2(n14580), .ZN(n14583) );
  NAND2_X1 U11767 ( .A1(n14579), .A2(n15883), .ZN(n14580) );
  XNOR2_X1 U11768 ( .A(n14591), .B(n14764), .ZN(n14762) );
  OR2_X1 U11769 ( .A1(n12580), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20170) );
  AND2_X1 U11770 ( .A1(n13338), .A2(n13333), .ZN(n20188) );
  INV_X1 U11771 ( .A(n16001), .ZN(n14787) );
  INV_X1 U11772 ( .A(n20455), .ZN(n20674) );
  AND2_X1 U11773 ( .A1(n16335), .A2(n13348), .ZN(n19965) );
  INV_X1 U11774 ( .A(n19035), .ZN(n19054) );
  INV_X1 U11775 ( .A(n19933), .ZN(n19479) );
  INV_X1 U11776 ( .A(n19218), .ZN(n19194) );
  AND2_X1 U11777 ( .A1(n19194), .A2(n10093), .ZN(n10097) );
  AND2_X1 U11778 ( .A1(n16227), .A2(n13485), .ZN(n19195) );
  NAND2_X1 U11779 ( .A1(n16308), .A2(n19188), .ZN(n10098) );
  NAND3_X1 U11780 ( .A1(n19902), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19761), 
        .ZN(n19218) );
  OR2_X1 U11781 ( .A1(n10148), .A2(n10280), .ZN(n10279) );
  NAND2_X1 U11782 ( .A1(n10277), .A2(n10278), .ZN(n10274) );
  NAND2_X1 U11783 ( .A1(n10148), .A2(n10298), .ZN(n10278) );
  NAND2_X1 U11784 ( .A1(n9736), .A2(n10147), .ZN(n10277) );
  INV_X1 U11785 ( .A(n10148), .ZN(n10147) );
  XNOR2_X1 U11786 ( .A(n10103), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15296) );
  NAND2_X1 U11787 ( .A1(n15138), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10103) );
  OAI21_X1 U11788 ( .B1(n15294), .B2(n19206), .A(n10101), .ZN(n10100) );
  NOR2_X1 U11789 ( .A1(n15295), .A2(n15293), .ZN(n10101) );
  OAI211_X1 U11790 ( .C1(n10056), .C2(n19206), .A(n15299), .B(n10055), .ZN(
        n10054) );
  INV_X1 U11791 ( .A(n15301), .ZN(n10056) );
  OR2_X1 U11792 ( .A1(n15302), .A2(n15303), .ZN(n10055) );
  NAND2_X1 U11793 ( .A1(n9711), .A2(n12881), .ZN(n15300) );
  OAI21_X1 U11794 ( .B1(n15328), .B2(n15314), .A(n10210), .ZN(n10209) );
  NOR2_X1 U11795 ( .A1(n15309), .A2(n10211), .ZN(n10210) );
  INV_X1 U11796 ( .A(n15313), .ZN(n10211) );
  NAND2_X1 U11797 ( .A1(n14937), .A2(n14938), .ZN(n15308) );
  OR2_X1 U11798 ( .A1(n16131), .A2(n19209), .ZN(n9978) );
  NOR2_X1 U11799 ( .A1(n15462), .A2(n9976), .ZN(n9975) );
  NOR2_X1 U11800 ( .A1(n9977), .A2(n19206), .ZN(n9976) );
  INV_X1 U11801 ( .A(n18950), .ZN(n9977) );
  AOI21_X1 U11802 ( .B1(n16127), .B2(n15459), .A(n15458), .ZN(n15464) );
  INV_X1 U11803 ( .A(n19204), .ZN(n16301) );
  INV_X1 U11804 ( .A(n19202), .ZN(n16306) );
  AND2_X1 U11805 ( .A1(n13618), .A2(n19944), .ZN(n19204) );
  INV_X1 U11806 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19939) );
  NOR2_X1 U11807 ( .A1(n13628), .A2(n12703), .ZN(n13944) );
  NAND2_X1 U11808 ( .A1(n13704), .A2(n13707), .ZN(n19904) );
  NOR2_X1 U11809 ( .A1(n17426), .A2(n9712), .ZN(n17285) );
  NAND2_X1 U11810 ( .A1(n17262), .A2(n17384), .ZN(n17377) );
  AND2_X1 U11811 ( .A1(n17345), .A2(n17262), .ZN(n17376) );
  XNOR2_X1 U11812 ( .A(n9807), .B(n18863), .ZN(n11499) );
  NAND2_X1 U11813 ( .A1(n16400), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9807) );
  OAI21_X1 U11814 ( .B1(n9931), .B2(n11471), .A(n9930), .ZN(n9929) );
  INV_X1 U11815 ( .A(n11473), .ZN(n9930) );
  NAND2_X1 U11816 ( .A1(n10125), .A2(n10124), .ZN(n10123) );
  INV_X1 U11817 ( .A(n11458), .ZN(n10122) );
  OAI221_X2 U11818 ( .B1(n11456), .B2(n18727), .C1(n11456), .C2(n11455), .A(
        n18901), .ZN(n18218) );
  NAND2_X1 U11819 ( .A1(n12288), .A2(n12287), .ZN(n12294) );
  NAND2_X1 U11820 ( .A1(n11113), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10174) );
  OR2_X1 U11821 ( .A1(n10631), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10606) );
  NOR2_X1 U11822 ( .A1(n10677), .A2(n12910), .ZN(n10681) );
  AND2_X1 U11823 ( .A1(n11514), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11515) );
  AOI22_X1 U11824 ( .A1(n11588), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11587), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11577) );
  NAND2_X1 U11825 ( .A1(n11759), .A2(n11758), .ZN(n11838) );
  OR2_X1 U11826 ( .A1(n11670), .A2(n11669), .ZN(n12514) );
  OR2_X1 U11827 ( .A1(n11715), .A2(n11714), .ZN(n11716) );
  INV_X1 U11828 ( .A(n11716), .ZN(n12522) );
  OR2_X1 U11829 ( .A1(n12294), .A2(n20220), .ZN(n12329) );
  NOR2_X1 U11830 ( .A1(n13315), .A2(n12592), .ZN(n12579) );
  NAND2_X1 U11831 ( .A1(n9813), .A2(n9812), .ZN(n11602) );
  NAND2_X1 U11832 ( .A1(n11601), .A2(n14820), .ZN(n9813) );
  NAND2_X1 U11833 ( .A1(n11600), .A2(n11576), .ZN(n11601) );
  OR2_X1 U11834 ( .A1(n11734), .A2(n11733), .ZN(n12534) );
  AND3_X1 U11835 ( .A1(n13654), .A2(n13336), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12326) );
  OR2_X1 U11836 ( .A1(n11127), .A2(n10957), .ZN(n10958) );
  NAND2_X1 U11837 ( .A1(n13617), .A2(n10949), .ZN(n10152) );
  INV_X1 U11838 ( .A(n10952), .ZN(n11131) );
  AOI21_X1 U11839 ( .B1(n10624), .B2(n16342), .A(n9877), .ZN(n10566) );
  NAND2_X1 U11840 ( .A1(n10568), .A2(n9874), .ZN(n9876) );
  NOR2_X1 U11841 ( .A1(n10027), .A2(n9860), .ZN(n10694) );
  NAND2_X1 U11842 ( .A1(n10023), .A2(n10019), .ZN(n10027) );
  NAND2_X1 U11843 ( .A1(n10663), .A2(n10024), .ZN(n10023) );
  OR2_X1 U11844 ( .A1(n10336), .A2(n10335), .ZN(n10734) );
  INV_X1 U11845 ( .A(n9866), .ZN(n10659) );
  OR2_X1 U11846 ( .A1(n10401), .A2(n10400), .ZN(n10696) );
  NAND2_X1 U11847 ( .A1(n10311), .A2(n10372), .ZN(n10373) );
  NAND2_X1 U11848 ( .A1(n13387), .A2(n10553), .ZN(n13392) );
  NAND2_X1 U11849 ( .A1(n10484), .A2(n10517), .ZN(n10008) );
  NAND2_X1 U11850 ( .A1(n10483), .A2(n10510), .ZN(n10007) );
  INV_X1 U11851 ( .A(n10479), .ZN(n10484) );
  OAI211_X1 U11852 ( .C1(n16983), .C2(n17134), .A(n9939), .B(n9726), .ZN(n9938) );
  NAND2_X1 U11853 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n9939) );
  AND2_X1 U11854 ( .A1(n9802), .A2(n9801), .ZN(n11191) );
  NAND2_X1 U11855 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n9802) );
  INV_X1 U11856 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n9942) );
  AOI21_X1 U11857 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18709), .A(
        n11418), .ZN(n11427) );
  AOI21_X1 U11858 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18718), .A(
        n11422), .ZN(n11431) );
  OAI21_X1 U11859 ( .B1(n11454), .B2(n17418), .A(n18702), .ZN(n11401) );
  NAND2_X1 U11860 ( .A1(n14348), .A2(n10272), .ZN(n10271) );
  INV_X1 U11861 ( .A(n14444), .ZN(n10272) );
  NAND2_X1 U11862 ( .A1(n11587), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n9811) );
  NAND2_X1 U11863 ( .A1(n9639), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n9810) );
  NOR2_X1 U11864 ( .A1(n10263), .A2(n10262), .ZN(n10261) );
  INV_X1 U11865 ( .A(n14258), .ZN(n10262) );
  INV_X1 U11866 ( .A(n12590), .ZN(n9829) );
  NAND2_X1 U11867 ( .A1(n10259), .A2(n10257), .ZN(n10256) );
  INV_X1 U11868 ( .A(n14463), .ZN(n10257) );
  AND2_X1 U11869 ( .A1(n14401), .A2(n14558), .ZN(n10259) );
  AND2_X1 U11870 ( .A1(n14209), .A2(n14193), .ZN(n10252) );
  AND2_X1 U11871 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11774), .ZN(
        n11815) );
  AND2_X1 U11872 ( .A1(n12571), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9843) );
  NAND2_X1 U11873 ( .A1(n11612), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12496) );
  INV_X1 U11874 ( .A(n12541), .ZN(n10142) );
  NAND2_X1 U11875 ( .A1(n10088), .A2(n13909), .ZN(n10089) );
  NOR2_X1 U11876 ( .A1(n13888), .A2(n16039), .ZN(n10088) );
  NAND2_X1 U11877 ( .A1(n13331), .A2(n12520), .ZN(n12529) );
  NAND2_X1 U11878 ( .A1(n11610), .A2(n13412), .ZN(n13326) );
  AND3_X1 U11879 ( .A1(n11642), .A2(n11641), .A3(n11640), .ZN(n11656) );
  AND4_X1 U11880 ( .A1(n11639), .A2(n11638), .A3(n11637), .A4(n11636), .ZN(
        n11641) );
  INV_X1 U11881 ( .A(n11655), .ZN(n10003) );
  AND2_X1 U11882 ( .A1(n11801), .A2(n10002), .ZN(n10001) );
  NAND2_X1 U11883 ( .A1(n11655), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10002) );
  NAND2_X1 U11884 ( .A1(n11693), .A2(n11692), .ZN(n11699) );
  XNOR2_X1 U11885 ( .A(n11678), .B(n11677), .ZN(n20315) );
  INV_X1 U11886 ( .A(n12592), .ZN(n10143) );
  NAND2_X1 U11887 ( .A1(n10956), .A2(n10955), .ZN(n11136) );
  NAND2_X1 U11888 ( .A1(n10951), .A2(n10950), .ZN(n11135) );
  NOR2_X1 U11889 ( .A1(n10907), .A2(n10168), .ZN(n10167) );
  INV_X1 U11890 ( .A(n15561), .ZN(n10040) );
  OR2_X1 U11891 ( .A1(n10450), .A2(n10449), .ZN(n12710) );
  NAND2_X1 U11892 ( .A1(n10150), .A2(n10149), .ZN(n10780) );
  NAND2_X1 U11893 ( .A1(n19251), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10149) );
  NAND2_X1 U11894 ( .A1(n10151), .A2(n10770), .ZN(n10150) );
  OAI21_X1 U11895 ( .B1(n10696), .B2(n13617), .A(n10152), .ZN(n10151) );
  OR2_X1 U11896 ( .A1(n10954), .A2(n10955), .ZN(n10951) );
  OR2_X1 U11897 ( .A1(n10417), .A2(n10416), .ZN(n10988) );
  OR2_X1 U11898 ( .A1(n10389), .A2(n10388), .ZN(n10981) );
  AND2_X1 U11899 ( .A1(n12991), .A2(n13004), .ZN(n10234) );
  AND2_X1 U11900 ( .A1(n13920), .A2(n13902), .ZN(n10207) );
  NAND2_X1 U11901 ( .A1(n10180), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10179) );
  INV_X1 U11902 ( .A(n10181), .ZN(n10180) );
  OR2_X1 U11903 ( .A1(n10182), .A2(n16171), .ZN(n10181) );
  NAND2_X1 U11904 ( .A1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10182) );
  INV_X1 U11905 ( .A(n14848), .ZN(n10058) );
  INV_X1 U11906 ( .A(n13248), .ZN(n10059) );
  NOR2_X1 U11907 ( .A1(n15311), .A2(n15327), .ZN(n9884) );
  NAND2_X1 U11908 ( .A1(n10927), .A2(n10926), .ZN(n10928) );
  AND2_X1 U11909 ( .A1(n14865), .A2(n10217), .ZN(n10216) );
  INV_X1 U11910 ( .A(n14954), .ZN(n10217) );
  AND2_X1 U11911 ( .A1(n10216), .A2(n10215), .ZN(n10214) );
  INV_X1 U11912 ( .A(n13246), .ZN(n10215) );
  AND2_X1 U11913 ( .A1(n12861), .A2(n13261), .ZN(n10046) );
  AND2_X1 U11914 ( .A1(n11013), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10105) );
  OAI21_X1 U11915 ( .B1(n10310), .B2(n10284), .A(n15395), .ZN(n10283) );
  NAND2_X1 U11916 ( .A1(n16151), .A2(n15200), .ZN(n9900) );
  NOR2_X1 U11917 ( .A1(n9687), .A2(n9903), .ZN(n9902) );
  AND2_X1 U11918 ( .A1(n13260), .A2(n13261), .ZN(n13275) );
  AND2_X1 U11919 ( .A1(n12851), .A2(n12850), .ZN(n14895) );
  INV_X1 U11920 ( .A(n15114), .ZN(n10043) );
  NAND2_X1 U11921 ( .A1(n10295), .A2(n10291), .ZN(n15201) );
  NOR2_X1 U11922 ( .A1(n14114), .A2(n10052), .ZN(n10051) );
  INV_X1 U11923 ( .A(n15539), .ZN(n10052) );
  NOR2_X1 U11924 ( .A1(n10203), .A2(n11031), .ZN(n10202) );
  INV_X1 U11925 ( .A(n10204), .ZN(n10203) );
  NOR2_X1 U11926 ( .A1(n13758), .A2(n10205), .ZN(n10204) );
  INV_X1 U11927 ( .A(n13784), .ZN(n10205) );
  OR2_X1 U11928 ( .A1(n10987), .A2(n14014), .ZN(n9871) );
  INV_X1 U11929 ( .A(n10650), .ZN(n10649) );
  NAND2_X1 U11930 ( .A1(n10766), .A2(n10765), .ZN(n10989) );
  NAND2_X1 U11931 ( .A1(n12686), .A2(n12685), .ZN(n13457) );
  OR2_X1 U11932 ( .A1(n12877), .A2(n10595), .ZN(n12689) );
  INV_X1 U11933 ( .A(n10696), .ZN(n12707) );
  AND3_X1 U11934 ( .A1(n10573), .A2(n12911), .A3(n16342), .ZN(n10608) );
  AND2_X1 U11935 ( .A1(n9887), .A2(n10573), .ZN(n9878) );
  NAND2_X1 U11936 ( .A1(n9704), .A2(n10230), .ZN(n10229) );
  NAND2_X1 U11937 ( .A1(n10226), .A2(n11020), .ZN(n10225) );
  OR2_X1 U11938 ( .A1(n12927), .A2(n12913), .ZN(n12915) );
  NAND2_X1 U11939 ( .A1(n10352), .A2(n10351), .ZN(n10587) );
  AOI22_X1 U11940 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9637), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10525) );
  NOR2_X1 U11941 ( .A1(n10499), .A2(n10498), .ZN(n10578) );
  INV_X1 U11942 ( .A(n19904), .ZN(n19519) );
  OR2_X1 U11943 ( .A1(n10952), .A2(n11135), .ZN(n10961) );
  INV_X1 U11944 ( .A(n11136), .ZN(n11140) );
  NAND2_X1 U11945 ( .A1(n18872), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11151) );
  NOR2_X1 U11946 ( .A1(n17040), .A2(n17209), .ZN(n10110) );
  NAND4_X1 U11947 ( .A1(n18872), .A2(n18880), .A3(n18860), .A4(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17155) );
  INV_X1 U11948 ( .A(n11399), .ZN(n11392) );
  OR2_X1 U11949 ( .A1(n16395), .A2(n16574), .ZN(n11491) );
  NAND2_X1 U11950 ( .A1(n17823), .A2(n11257), .ZN(n11260) );
  INV_X1 U11951 ( .A(n10120), .ZN(n10118) );
  NOR2_X1 U11952 ( .A1(n10116), .A2(n9798), .ZN(n10115) );
  INV_X1 U11953 ( .A(n11254), .ZN(n10116) );
  INV_X1 U11954 ( .A(n10119), .ZN(n9798) );
  AND2_X1 U11955 ( .A1(n9806), .A2(n9766), .ZN(n11378) );
  XNOR2_X1 U11956 ( .A(n9797), .B(n11364), .ZN(n11250) );
  NOR3_X1 U11957 ( .A1(n11392), .A2(n11443), .A3(n18683), .ZN(n15609) );
  AND2_X1 U11958 ( .A1(n12348), .A2(n12347), .ZN(n13422) );
  NAND2_X1 U11959 ( .A1(n14301), .A2(n12469), .ZN(n14275) );
  INV_X1 U11960 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15841) );
  OR3_X1 U11961 ( .A1(n20802), .A2(n12464), .A3(n20022), .ZN(n19998) );
  NAND2_X1 U11962 ( .A1(n14407), .A2(n12463), .ZN(n20051) );
  OR2_X1 U11963 ( .A1(n20869), .A2(n12352), .ZN(n14217) );
  NOR2_X1 U11964 ( .A1(n13928), .A2(n20212), .ZN(n12462) );
  INV_X1 U11965 ( .A(n14248), .ZN(n10072) );
  NAND2_X1 U11966 ( .A1(n10081), .A2(n10080), .ZN(n10079) );
  INV_X1 U11967 ( .A(n10082), .ZN(n10081) );
  NOR2_X1 U11968 ( .A1(n10084), .A2(n14324), .ZN(n10080) );
  AND2_X1 U11969 ( .A1(n12411), .A2(n12410), .ZN(n14390) );
  NOR2_X1 U11970 ( .A1(n14460), .A2(n14390), .ZN(n14392) );
  INV_X1 U11971 ( .A(n12025), .ZN(n14446) );
  AND3_X1 U11972 ( .A1(n11860), .A2(n11859), .A3(n11858), .ZN(n14147) );
  NAND2_X1 U11973 ( .A1(n13651), .A2(n9752), .ZN(n13653) );
  OR2_X1 U11974 ( .A1(n13650), .A2(n9925), .ZN(n13651) );
  NAND2_X1 U11975 ( .A1(n14282), .A2(n10261), .ZN(n14257) );
  AND2_X1 U11976 ( .A1(n12223), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12224) );
  INV_X1 U11977 ( .A(n10263), .ZN(n10260) );
  AND2_X1 U11978 ( .A1(n12175), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12176) );
  NAND2_X1 U11979 ( .A1(n12176), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12222) );
  NAND2_X1 U11980 ( .A1(n10267), .A2(n10266), .ZN(n10265) );
  INV_X1 U11981 ( .A(n10269), .ZN(n10267) );
  INV_X1 U11982 ( .A(n14323), .ZN(n10266) );
  NAND2_X1 U11983 ( .A1(n12084), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12129) );
  AND2_X1 U11984 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12083), .ZN(
        n12084) );
  INV_X1 U11985 ( .A(n12069), .ZN(n12083) );
  NOR2_X1 U11986 ( .A1(n12040), .A2(n14369), .ZN(n12041) );
  NAND2_X1 U11987 ( .A1(n12041), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12069) );
  NOR2_X1 U11988 ( .A1(n12009), .A2(n14383), .ZN(n12010) );
  NAND2_X1 U11989 ( .A1(n12505), .A2(n14793), .ZN(n14669) );
  CLKBUF_X1 U11990 ( .A(n14375), .Z(n14376) );
  NAND2_X1 U11991 ( .A1(n11959), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11974) );
  NAND2_X1 U11992 ( .A1(n10313), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14806) );
  AND2_X1 U11993 ( .A1(n9850), .A2(n9849), .ZN(n14809) );
  INV_X1 U11994 ( .A(n14688), .ZN(n9850) );
  NOR2_X1 U11995 ( .A1(n15873), .A2(n14690), .ZN(n9849) );
  NOR2_X1 U11996 ( .A1(n11942), .A2(n14405), .ZN(n11959) );
  INV_X1 U11997 ( .A(n14558), .ZN(n10258) );
  AND2_X1 U11998 ( .A1(n11891), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11892) );
  NAND2_X1 U11999 ( .A1(n11892), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11937) );
  INV_X1 U12000 ( .A(n14472), .ZN(n11909) );
  NOR2_X1 U12001 ( .A1(n11887), .A2(n11886), .ZN(n11891) );
  INV_X1 U12002 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11775) );
  AOI21_X1 U12003 ( .B1(n12559), .B2(n11971), .A(n11780), .ZN(n14126) );
  NAND2_X1 U12004 ( .A1(n11839), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11782) );
  XNOR2_X1 U12005 ( .A(n12529), .B(n20191), .ZN(n13894) );
  AOI21_X1 U12006 ( .B1(n11791), .B2(n11955), .A(n9823), .ZN(n9822) );
  INV_X1 U12007 ( .A(n11811), .ZN(n9823) );
  NAND2_X1 U12008 ( .A1(n13330), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13331) );
  NAND2_X1 U12009 ( .A1(n14568), .A2(n14566), .ZN(n9918) );
  NAND2_X1 U12010 ( .A1(n14764), .A2(n14582), .ZN(n9919) );
  AND2_X1 U12011 ( .A1(n12577), .A2(n9920), .ZN(n14567) );
  NAND2_X1 U12012 ( .A1(n14764), .A2(n12435), .ZN(n10060) );
  AND2_X1 U12013 ( .A1(n14295), .A2(n14289), .ZN(n14287) );
  NAND2_X1 U12014 ( .A1(n14599), .A2(n12576), .ZN(n14589) );
  OR2_X1 U12015 ( .A1(n9714), .A2(n14314), .ZN(n14312) );
  NOR2_X1 U12016 ( .A1(n14312), .A2(n14294), .ZN(n14295) );
  NAND2_X1 U12017 ( .A1(n14662), .A2(n10145), .ZN(n9911) );
  AND2_X1 U12018 ( .A1(n9724), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10145) );
  OR2_X1 U12019 ( .A1(n14662), .A2(n9789), .ZN(n9927) );
  NOR2_X1 U12020 ( .A1(n14441), .A2(n14440), .ZN(n14442) );
  NOR3_X1 U12021 ( .A1(n14441), .A2(n10084), .A3(n14440), .ZN(n14351) );
  OR2_X1 U12022 ( .A1(n14448), .A2(n14364), .ZN(n14441) );
  NAND2_X1 U12023 ( .A1(n14662), .A2(n14661), .ZN(n14651) );
  AND2_X1 U12024 ( .A1(n14392), .A2(n14380), .ZN(n14450) );
  NAND2_X1 U12025 ( .A1(n14450), .A2(n14449), .ZN(n14448) );
  NAND2_X1 U12026 ( .A1(n12402), .A2(n10077), .ZN(n10074) );
  INV_X1 U12027 ( .A(n14461), .ZN(n10077) );
  NOR3_X1 U12028 ( .A1(n14476), .A2(n10078), .A3(n14475), .ZN(n14465) );
  OAI21_X1 U12029 ( .B1(n10313), .B2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n14806), .ZN(n14690) );
  NOR2_X1 U12030 ( .A1(n14476), .A2(n14475), .ZN(n15840) );
  AND2_X1 U12031 ( .A1(n12394), .A2(n12393), .ZN(n14210) );
  INV_X1 U12032 ( .A(n10131), .ZN(n10130) );
  NOR2_X1 U12033 ( .A1(n16026), .A2(n14150), .ZN(n16011) );
  AND2_X1 U12034 ( .A1(n12384), .A2(n12383), .ZN(n16022) );
  OR2_X1 U12035 ( .A1(n13889), .A2(n10089), .ZN(n16042) );
  OR2_X1 U12036 ( .A1(n13889), .A2(n10090), .ZN(n16040) );
  NAND2_X1 U12037 ( .A1(n10087), .A2(n13909), .ZN(n10090) );
  INV_X1 U12038 ( .A(n13888), .ZN(n10087) );
  NOR2_X1 U12039 ( .A1(n13889), .A2(n13888), .ZN(n13910) );
  AND2_X1 U12040 ( .A1(n12368), .A2(n12367), .ZN(n13852) );
  NAND2_X1 U12041 ( .A1(n12370), .A2(n12369), .ZN(n13889) );
  INV_X1 U12042 ( .A(n13852), .ZN(n12369) );
  INV_X1 U12043 ( .A(n10066), .ZN(n12370) );
  OR2_X1 U12044 ( .A1(n13334), .A2(n15785), .ZN(n16001) );
  CLKBUF_X1 U12045 ( .A(n12341), .Z(n13420) );
  NAND2_X1 U12046 ( .A1(n9814), .A2(n11685), .ZN(n12512) );
  NAND2_X1 U12047 ( .A1(n11674), .A2(n9747), .ZN(n9819) );
  AND2_X1 U12048 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20721), .ZN(n13869) );
  INV_X1 U12049 ( .A(n11812), .ZN(n10005) );
  INV_X1 U12050 ( .A(n12599), .ZN(n10128) );
  AND2_X1 U12051 ( .A1(n14089), .A2(n14816), .ZN(n20314) );
  INV_X1 U12052 ( .A(n20508), .ZN(n20670) );
  NAND2_X1 U12053 ( .A1(n20283), .A2(n14090), .ZN(n20553) );
  NAND2_X1 U12054 ( .A1(n20154), .A2(n14481), .ZN(n20247) );
  INV_X1 U12055 ( .A(n20719), .ZN(n20721) );
  INV_X1 U12056 ( .A(n20321), .ZN(n20717) );
  NAND2_X1 U12057 ( .A1(n10924), .A2(n9716), .ZN(n10918) );
  NAND2_X1 U12058 ( .A1(n10942), .A2(n10941), .ZN(n10945) );
  NOR2_X1 U12059 ( .A1(n10932), .A2(n10933), .ZN(n10942) );
  NAND2_X1 U12060 ( .A1(n10918), .A2(n10929), .ZN(n10932) );
  NAND2_X1 U12061 ( .A1(n18993), .A2(n10189), .ZN(n10187) );
  NAND2_X1 U12062 ( .A1(n10189), .A2(n12626), .ZN(n10188) );
  NAND2_X1 U12063 ( .A1(n12630), .A2(n10195), .ZN(n10194) );
  INV_X1 U12064 ( .A(n15192), .ZN(n10195) );
  NAND2_X1 U12065 ( .A1(n18993), .A2(n12630), .ZN(n10193) );
  NAND2_X1 U12066 ( .A1(n10861), .A2(n10167), .ZN(n10911) );
  NOR2_X1 U12067 ( .A1(n13282), .A2(n15192), .ZN(n13281) );
  NOR2_X2 U12068 ( .A1(n10868), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10864) );
  NOR2_X1 U12069 ( .A1(n10475), .A2(n10158), .ZN(n10157) );
  NAND2_X1 U12070 ( .A1(n10881), .A2(n10156), .ZN(n10875) );
  CLKBUF_X1 U12071 ( .A(n12640), .Z(n12641) );
  NAND2_X1 U12072 ( .A1(n10881), .A2(n10880), .ZN(n10878) );
  INV_X1 U12073 ( .A(n10473), .ZN(n10848) );
  INV_X1 U12074 ( .A(n10924), .ZN(n10154) );
  NAND2_X1 U12075 ( .A1(n10162), .A2(n10164), .ZN(n10825) );
  INV_X1 U12076 ( .A(n10824), .ZN(n10163) );
  NOR2_X1 U12077 ( .A1(n10763), .A2(n10762), .ZN(n10819) );
  XNOR2_X1 U12078 ( .A(n9866), .B(n10658), .ZN(n9865) );
  INV_X1 U12079 ( .A(n11113), .ZN(n11121) );
  AND2_X1 U12080 ( .A1(n11081), .A2(n11080), .ZN(n13258) );
  AND2_X1 U12081 ( .A1(n11070), .A2(n11069), .ZN(n14908) );
  NAND2_X1 U12082 ( .A1(n9764), .A2(n13862), .ZN(n9968) );
  INV_X1 U12083 ( .A(n10224), .ZN(n10223) );
  AND2_X1 U12084 ( .A1(n13901), .A2(n13902), .ZN(n13921) );
  AND2_X1 U12085 ( .A1(n9705), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10236) );
  AND2_X1 U12086 ( .A1(n9708), .A2(n14860), .ZN(n10044) );
  NAND2_X1 U12087 ( .A1(n10222), .A2(n10220), .ZN(n10219) );
  INV_X1 U12088 ( .A(n14979), .ZN(n10220) );
  AND2_X1 U12089 ( .A1(n15004), .A2(n9770), .ZN(n13065) );
  INV_X1 U12090 ( .A(n13087), .ZN(n9969) );
  NOR2_X1 U12091 ( .A1(n15485), .A2(n14922), .ZN(n15113) );
  NAND2_X1 U12092 ( .A1(n15484), .A2(n15486), .ZN(n15485) );
  AND2_X1 U12093 ( .A1(n13147), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13750) );
  AND2_X1 U12094 ( .A1(n13475), .A2(n19955), .ZN(n19140) );
  AND2_X1 U12095 ( .A1(n12887), .A2(n13348), .ZN(n13355) );
  INV_X1 U12096 ( .A(n13525), .ZN(n19219) );
  CLKBUF_X1 U12097 ( .A(n12622), .Z(n12623) );
  CLKBUF_X1 U12098 ( .A(n12627), .Z(n12628) );
  NAND2_X1 U12099 ( .A1(n14973), .A2(n14865), .ZN(n14864) );
  OR2_X1 U12100 ( .A1(n13285), .A2(n13286), .ZN(n14972) );
  NOR2_X1 U12101 ( .A1(n14972), .A2(n14971), .ZN(n14973) );
  CLKBUF_X1 U12102 ( .A(n12631), .Z(n12632) );
  CLKBUF_X1 U12103 ( .A(n12634), .Z(n12635) );
  AND2_X1 U12104 ( .A1(n11077), .A2(n11076), .ZN(n14879) );
  NAND2_X1 U12105 ( .A1(n14909), .A2(n10198), .ZN(n14877) );
  CLKBUF_X1 U12106 ( .A(n12637), .Z(n12638) );
  AND2_X1 U12107 ( .A1(n11066), .A2(n11065), .ZN(n15016) );
  NAND2_X1 U12108 ( .A1(n10171), .A2(n10170), .ZN(n15013) );
  INV_X1 U12109 ( .A(n15016), .ZN(n10170) );
  INV_X1 U12110 ( .A(n15015), .ZN(n10171) );
  CLKBUF_X1 U12111 ( .A(n12643), .Z(n12644) );
  AND2_X1 U12112 ( .A1(n11050), .A2(n11049), .ZN(n14170) );
  NAND2_X1 U12113 ( .A1(n13901), .A2(n9749), .ZN(n14169) );
  AND2_X1 U12114 ( .A1(n13901), .A2(n10207), .ZN(n14021) );
  CLKBUF_X1 U12115 ( .A(n9717), .Z(n12660) );
  CLKBUF_X1 U12116 ( .A(n12648), .Z(n12659) );
  NOR2_X1 U12117 ( .A1(n13757), .A2(n10201), .ZN(n13857) );
  INV_X1 U12118 ( .A(n10202), .ZN(n10201) );
  CLKBUF_X1 U12119 ( .A(n12650), .Z(n12651) );
  CLKBUF_X1 U12120 ( .A(n12654), .Z(n12655) );
  INV_X1 U12121 ( .A(n10298), .ZN(n10280) );
  INV_X1 U12122 ( .A(n15134), .ZN(n10281) );
  XNOR2_X1 U12123 ( .A(n10477), .B(n15289), .ZN(n10148) );
  NOR2_X1 U12124 ( .A1(n14841), .A2(n10899), .ZN(n10477) );
  OR3_X1 U12125 ( .A1(n12896), .A2(n10899), .A3(n15280), .ZN(n15123) );
  AND2_X1 U12126 ( .A1(n14973), .A2(n10212), .ZN(n14936) );
  AND2_X1 U12127 ( .A1(n10214), .A2(n10213), .ZN(n10212) );
  INV_X1 U12128 ( .A(n14845), .ZN(n10213) );
  NOR2_X1 U12129 ( .A1(n14856), .A2(n10899), .ZN(n15145) );
  NOR2_X1 U12130 ( .A1(n13244), .A2(n10899), .ZN(n15144) );
  NAND2_X1 U12131 ( .A1(n14973), .A2(n10216), .ZN(n14956) );
  NAND2_X1 U12132 ( .A1(n14973), .A2(n10214), .ZN(n14846) );
  NAND2_X1 U12133 ( .A1(n13260), .A2(n10046), .ZN(n15082) );
  INV_X1 U12134 ( .A(n13275), .ZN(n13288) );
  NOR2_X1 U12135 ( .A1(n14911), .A2(n14895), .ZN(n14882) );
  NAND2_X1 U12136 ( .A1(n14909), .A2(n14893), .ZN(n14876) );
  NAND2_X1 U12137 ( .A1(n10042), .A2(n10041), .ZN(n14911) );
  NOR2_X1 U12138 ( .A1(n9701), .A2(n9786), .ZN(n10041) );
  INV_X1 U12139 ( .A(n15485), .ZN(n10042) );
  NAND2_X1 U12140 ( .A1(n15030), .A2(n14925), .ZN(n15015) );
  NAND2_X1 U12141 ( .A1(n16240), .A2(n15519), .ZN(n15518) );
  AND2_X1 U12142 ( .A1(n9721), .A2(n15423), .ZN(n9982) );
  AOI21_X1 U12143 ( .B1(n16198), .B2(n10291), .A(n10030), .ZN(n10029) );
  INV_X1 U12144 ( .A(n15202), .ZN(n10030) );
  NOR2_X1 U12145 ( .A1(n9748), .A2(n10049), .ZN(n10048) );
  INV_X1 U12146 ( .A(n16255), .ZN(n10049) );
  NOR2_X1 U12147 ( .A1(n16254), .A2(n16241), .ZN(n16240) );
  NAND2_X1 U12148 ( .A1(n9979), .A2(n9686), .ZN(n16165) );
  NAND2_X1 U12149 ( .A1(n16194), .A2(n9721), .ZN(n9979) );
  NAND2_X1 U12150 ( .A1(n10290), .A2(n10293), .ZN(n16173) );
  AND2_X1 U12151 ( .A1(n10845), .A2(n16269), .ZN(n16176) );
  AND3_X1 U12152 ( .A1(n12763), .A2(n12762), .A3(n12761), .ZN(n14134) );
  NAND2_X1 U12153 ( .A1(n10047), .A2(n10051), .ZN(n15538) );
  NOR2_X1 U12154 ( .A1(n16289), .A2(n9748), .ZN(n16256) );
  NAND2_X1 U12155 ( .A1(n16194), .A2(n16192), .ZN(n9983) );
  OAI22_X1 U12156 ( .A1(n13989), .A2(n12715), .B1(n10899), .B2(n12842), .ZN(
        n16291) );
  XNOR2_X1 U12157 ( .A(n11008), .B(n10899), .ZN(n15256) );
  OR2_X1 U12158 ( .A1(n14007), .A2(n19201), .ZN(n16257) );
  NAND2_X1 U12159 ( .A1(n10200), .A2(n10204), .ZN(n13782) );
  NOR2_X1 U12160 ( .A1(n13757), .A2(n13758), .ZN(n13783) );
  NAND2_X1 U12161 ( .A1(n15566), .A2(n9680), .ZN(n9881) );
  NAND2_X1 U12162 ( .A1(n9974), .A2(n9973), .ZN(n15570) );
  AND2_X1 U12163 ( .A1(n11020), .A2(n11019), .ZN(n13755) );
  NAND2_X1 U12164 ( .A1(n12794), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12688) );
  AND2_X1 U12165 ( .A1(n13457), .A2(n13458), .ZN(n13456) );
  INV_X1 U12166 ( .A(n14079), .ZN(n18971) );
  NAND2_X1 U12167 ( .A1(n10653), .A2(n10656), .ZN(n19193) );
  INV_X1 U12168 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14182) );
  NOR2_X1 U12169 ( .A1(n12923), .A2(n9964), .ZN(n9963) );
  AND2_X1 U12170 ( .A1(n13470), .A2(n12933), .ZN(n13646) );
  NAND2_X1 U12171 ( .A1(n13645), .A2(n12934), .ZN(n13705) );
  AND2_X1 U12172 ( .A1(n19913), .A2(n19903), .ZN(n19276) );
  AND2_X1 U12173 ( .A1(n19904), .A2(n19479), .ZN(n19454) );
  INV_X1 U12174 ( .A(n19276), .ZN(n19520) );
  AND2_X1 U12175 ( .A1(n19913), .A2(n19923), .ZN(n19899) );
  OR2_X1 U12176 ( .A1(n19913), .A2(n19923), .ZN(n19651) );
  NAND2_X2 U12177 ( .A1(n10551), .A2(n10550), .ZN(n19237) );
  NAND2_X1 U12178 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19761), .ZN(n19250) );
  NOR2_X1 U12179 ( .A1(n19904), .A2(n19479), .ZN(n19712) );
  INV_X1 U12180 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16351) );
  NOR2_X1 U12181 ( .A1(n17889), .A2(n11491), .ZN(n16391) );
  AND2_X1 U12182 ( .A1(n16846), .A2(n9944), .ZN(n16659) );
  NAND2_X1 U12183 ( .A1(n16548), .A2(n16890), .ZN(n9944) );
  NOR2_X1 U12184 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16715), .ZN(n16704) );
  NAND2_X1 U12185 ( .A1(n16391), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16374) );
  NOR2_X1 U12186 ( .A1(n17422), .A2(n17424), .ZN(n9851) );
  NAND2_X1 U12187 ( .A1(n9856), .A2(n9854), .ZN(n17266) );
  NOR2_X1 U12188 ( .A1(n11338), .A2(n9855), .ZN(n9854) );
  INV_X1 U12189 ( .A(n11337), .ZN(n9856) );
  AND2_X1 U12190 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n9855) );
  NAND3_X1 U12191 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18691), .A3(
        n18887), .ZN(n17191) );
  INV_X1 U12192 ( .A(n11224), .ZN(n9940) );
  NOR2_X1 U12193 ( .A1(n11201), .A2(n11200), .ZN(n11237) );
  NAND2_X1 U12194 ( .A1(n11199), .A2(n11198), .ZN(n11200) );
  NAND2_X1 U12195 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11198) );
  NAND2_X1 U12196 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11211) );
  NAND2_X1 U12197 ( .A1(n18259), .A2(n17266), .ZN(n18702) );
  NOR2_X1 U12198 ( .A1(n17479), .A2(n17417), .ZN(n17446) );
  OR2_X1 U12199 ( .A1(n17538), .A2(n17539), .ZN(n16395) );
  AND2_X1 U12200 ( .A1(n17641), .A2(n9948), .ZN(n17563) );
  AND2_X1 U12201 ( .A1(n9700), .A2(n9949), .ZN(n9948) );
  INV_X1 U12202 ( .A(n17581), .ZN(n9949) );
  NOR2_X1 U12203 ( .A1(n17616), .A2(n9951), .ZN(n9950) );
  NAND2_X1 U12204 ( .A1(n17641), .A2(n9700), .ZN(n17580) );
  NAND2_X1 U12205 ( .A1(n17641), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17615) );
  NAND2_X1 U12206 ( .A1(n17794), .A2(n9682), .ZN(n17728) );
  NAND2_X1 U12207 ( .A1(n11264), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17760) );
  NOR2_X1 U12208 ( .A1(n11469), .A2(n17737), .ZN(n11471) );
  NAND2_X1 U12209 ( .A1(n9933), .A2(n9932), .ZN(n9931) );
  INV_X1 U12210 ( .A(n11485), .ZN(n9932) );
  NAND2_X1 U12211 ( .A1(n11472), .A2(n11478), .ZN(n9933) );
  NOR2_X1 U12212 ( .A1(n11445), .A2(n11434), .ZN(n11489) );
  NAND2_X1 U12213 ( .A1(n17577), .A2(n17908), .ZN(n17911) );
  NOR2_X1 U12214 ( .A1(n17591), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17590) );
  NOR2_X1 U12215 ( .A1(n17609), .A2(n17627), .ZN(n17667) );
  NOR2_X1 U12216 ( .A1(n11268), .A2(n9794), .ZN(n9793) );
  NAND2_X1 U12217 ( .A1(n9796), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9795) );
  AND2_X1 U12218 ( .A1(n17805), .A2(n18040), .ZN(n9794) );
  AND2_X1 U12219 ( .A1(n9804), .A2(n17685), .ZN(n17968) );
  AOI21_X1 U12220 ( .B1(n11410), .B2(n16530), .A(n11411), .ZN(n18681) );
  NOR2_X1 U12221 ( .A1(n11385), .A2(n9805), .ZN(n17802) );
  AND2_X1 U12222 ( .A1(n11386), .A2(n11387), .ZN(n9805) );
  NOR2_X1 U12223 ( .A1(n17802), .A2(n18130), .ZN(n17801) );
  XNOR2_X1 U12224 ( .A(n11260), .B(n11259), .ZN(n17811) );
  NAND2_X1 U12225 ( .A1(n17811), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17810) );
  XNOR2_X1 U12226 ( .A(n11378), .B(n11379), .ZN(n17830) );
  NOR2_X1 U12227 ( .A1(n17830), .A2(n18150), .ZN(n17829) );
  XNOR2_X1 U12228 ( .A(n11249), .B(n10106), .ZN(n17866) );
  INV_X1 U12229 ( .A(n11250), .ZN(n10106) );
  NAND2_X1 U12230 ( .A1(n17885), .A2(n11247), .ZN(n17879) );
  NAND2_X1 U12231 ( .A1(n17879), .A2(n17880), .ZN(n17878) );
  NOR2_X1 U12232 ( .A1(n11411), .A2(n11412), .ZN(n15707) );
  NAND2_X1 U12233 ( .A1(n11398), .A2(n11397), .ZN(n18694) );
  INV_X1 U12234 ( .A(n18188), .ZN(n18723) );
  NAND2_X1 U12235 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18691), .ZN(
        n18686) );
  AOI211_X1 U12236 ( .C1(n17184), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n11328), .B(n11327), .ZN(n18250) );
  INV_X1 U12237 ( .A(n17266), .ZN(n18254) );
  INV_X1 U12238 ( .A(n11391), .ZN(n18259) );
  INV_X1 U12239 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18749) );
  NAND2_X1 U12240 ( .A1(n9839), .A2(n9838), .ZN(n13773) );
  NOR2_X1 U12241 ( .A1(n13420), .A2(n15762), .ZN(n9838) );
  INV_X1 U12242 ( .A(n13715), .ZN(n9839) );
  OR2_X1 U12243 ( .A1(n13415), .A2(n15762), .ZN(n13375) );
  INV_X1 U12244 ( .A(n13417), .ZN(n11607) );
  NAND2_X1 U12245 ( .A1(n13773), .A2(n13375), .ZN(n20869) );
  INV_X1 U12246 ( .A(n14241), .ZN(n12480) );
  AND2_X1 U12247 ( .A1(n12467), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n14355) );
  NOR2_X1 U12248 ( .A1(n15828), .A2(n12466), .ZN(n15815) );
  NAND2_X1 U12249 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n9722), .ZN(n15828) );
  NOR2_X1 U12250 ( .A1(n20008), .A2(n9836), .ZN(n15837) );
  NAND2_X1 U12251 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .ZN(n9836) );
  INV_X1 U12252 ( .A(n14407), .ZN(n14416) );
  CLKBUF_X1 U12253 ( .A(n13800), .Z(n20454) );
  AND2_X1 U12254 ( .A1(n12462), .A2(n12460), .ZN(n14407) );
  INV_X1 U12255 ( .A(n20048), .ZN(n20000) );
  INV_X1 U12256 ( .A(n20054), .ZN(n15848) );
  INV_X1 U12257 ( .A(n14467), .ZN(n20070) );
  AND2_X2 U12258 ( .A1(n13720), .A2(n19975), .ZN(n20075) );
  NAND2_X1 U12259 ( .A1(n20075), .A2(n14104), .ZN(n14467) );
  OR2_X1 U12260 ( .A1(n12615), .A2(n14481), .ZN(n14532) );
  INV_X1 U12261 ( .A(n14530), .ZN(n14540) );
  INV_X1 U12262 ( .A(n14524), .ZN(n14543) );
  NAND2_X1 U12263 ( .A1(n14550), .A2(n13743), .ZN(n14562) );
  BUF_X1 U12264 ( .A(n20102), .Z(n20872) );
  CLKBUF_X1 U12265 ( .A(n15781), .Z(n20101) );
  XNOR2_X1 U12266 ( .A(n12355), .B(n12354), .ZN(n13224) );
  OR2_X1 U12267 ( .A1(n12353), .A2(n12485), .ZN(n12355) );
  NAND2_X1 U12268 ( .A1(n9641), .A2(n12479), .ZN(n12280) );
  AND2_X1 U12269 ( .A1(n14662), .A2(n9724), .ZN(n14644) );
  NOR2_X1 U12270 ( .A1(n13963), .A2(n13964), .ZN(n13981) );
  INV_X1 U12271 ( .A(n12495), .ZN(n20154) );
  OAI21_X1 U12272 ( .B1(n15893), .B2(n9986), .A(n10129), .ZN(n14228) );
  AOI21_X1 U12273 ( .B1(n10135), .B2(n10134), .A(n10133), .ZN(n10129) );
  NAND2_X1 U12274 ( .A1(n10136), .A2(n12566), .ZN(n14196) );
  NAND2_X1 U12275 ( .A1(n15893), .A2(n12565), .ZN(n10136) );
  NAND2_X1 U12276 ( .A1(n13906), .A2(n12541), .ZN(n15904) );
  INV_X1 U12277 ( .A(n16014), .ZN(n20203) );
  INV_X1 U12278 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20634) );
  NAND2_X1 U12279 ( .A1(n11803), .A2(n16055), .ZN(n10000) );
  INV_X1 U12280 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20582) );
  NAND2_X1 U12281 ( .A1(n11773), .A2(n20590), .ZN(n20719) );
  OR2_X1 U12282 ( .A1(n13715), .A2(n20590), .ZN(n13837) );
  OR2_X1 U12283 ( .A1(n9915), .A2(n20579), .ZN(n13642) );
  OAI21_X1 U12284 ( .B1(n20289), .B2(n20288), .A(n20287), .ZN(n20309) );
  OAI21_X1 U12285 ( .B1(n20370), .B2(n20354), .A(n20678), .ZN(n20372) );
  OAI211_X1 U12286 ( .C1(n20420), .C2(n20590), .A(n20678), .B(n20405), .ZN(
        n20422) );
  OAI211_X1 U12287 ( .C1(n20479), .C2(n20590), .A(n20516), .B(n20463), .ZN(
        n20481) );
  INV_X1 U12288 ( .A(n20520), .ZN(n20542) );
  NAND2_X1 U12289 ( .A1(n20243), .A2(n11576), .ZN(n20620) );
  OAI211_X1 U12290 ( .C1(n20591), .C2(n20590), .A(n20678), .B(n20589), .ZN(
        n20629) );
  OAI211_X1 U12291 ( .C1(n20703), .C2(n20679), .A(n20678), .B(n20677), .ZN(
        n20705) );
  INV_X1 U12292 ( .A(n20605), .ZN(n20739) );
  INV_X1 U12293 ( .A(n20620), .ZN(n20757) );
  INV_X1 U12294 ( .A(n20762), .ZN(n20769) );
  OR2_X1 U12295 ( .A1(n20716), .A2(n20553), .ZN(n20773) );
  OR2_X1 U12296 ( .A1(n20775), .A2(n16055), .ZN(n15762) );
  INV_X1 U12297 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16053) );
  INV_X1 U12298 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20590) );
  OAI21_X1 U12299 ( .B1(n10160), .B2(n10770), .A(n10159), .ZN(n14841) );
  NAND2_X1 U12300 ( .A1(n10918), .A2(n10770), .ZN(n10159) );
  NOR2_X1 U12301 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n10945), .ZN(n10160) );
  NOR2_X1 U12302 ( .A1(n16070), .A2(n16071), .ZN(n16069) );
  INV_X1 U12303 ( .A(n18944), .ZN(n10176) );
  AND2_X1 U12304 ( .A1(n19965), .A2(n16361), .ZN(n19056) );
  INV_X1 U12305 ( .A(n19822), .ZN(n19049) );
  OR2_X1 U12306 ( .A1(n19965), .A2(n12885), .ZN(n19035) );
  CLKBUF_X1 U12307 ( .A(n18996), .Z(n19068) );
  CLKBUF_X1 U12308 ( .A(n15025), .Z(n15026) );
  CLKBUF_X1 U12309 ( .A(n14164), .Z(n14165) );
  OR2_X1 U12310 ( .A1(n12759), .A2(n12758), .ZN(n13900) );
  INV_X1 U12311 ( .A(n15019), .ZN(n15041) );
  INV_X1 U12312 ( .A(n19193), .ZN(n19207) );
  INV_X1 U12313 ( .A(n19923), .ZN(n19903) );
  XNOR2_X1 U12314 ( .A(n9972), .B(n9971), .ZN(n15058) );
  INV_X1 U12315 ( .A(n14945), .ZN(n9971) );
  NAND2_X1 U12316 ( .A1(n10240), .A2(n14944), .ZN(n9972) );
  NOR2_X1 U12317 ( .A1(n13166), .A2(n10241), .ZN(n14949) );
  INV_X1 U12318 ( .A(n19077), .ZN(n15116) );
  INV_X1 U12319 ( .A(n10035), .ZN(n10033) );
  NOR2_X1 U12320 ( .A1(n19085), .A2(n19131), .ZN(n19119) );
  NOR2_X1 U12321 ( .A1(n12703), .A2(n10039), .ZN(n10038) );
  OR2_X1 U12322 ( .A1(n13452), .A2(n13451), .ZN(n13453) );
  INV_X1 U12323 ( .A(n19135), .ZN(n19085) );
  INV_X1 U12324 ( .A(n19122), .ZN(n19131) );
  NOR2_X1 U12325 ( .A1(n19140), .A2(n19968), .ZN(n19154) );
  CLKBUF_X1 U12327 ( .A(n13701), .Z(n19968) );
  INV_X1 U12328 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16171) );
  INV_X1 U12329 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15264) );
  INV_X1 U12330 ( .A(n19195), .ZN(n19182) );
  INV_X1 U12331 ( .A(n16227), .ZN(n19187) );
  INV_X1 U12332 ( .A(n16209), .ZN(n19188) );
  NAND2_X1 U12333 ( .A1(n10286), .A2(n10310), .ZN(n15393) );
  NAND2_X1 U12334 ( .A1(n10858), .A2(n10285), .ZN(n10286) );
  AND2_X1 U12335 ( .A1(n15032), .A2(n15031), .ZN(n18957) );
  AND2_X1 U12336 ( .A1(n10290), .A2(n9756), .ZN(n16159) );
  NAND2_X1 U12337 ( .A1(n10290), .A2(n10830), .ZN(n15533) );
  NAND2_X1 U12338 ( .A1(n16216), .A2(n10987), .ZN(n14000) );
  AND2_X1 U12339 ( .A1(n19192), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10095) );
  INV_X1 U12340 ( .A(n10688), .ZN(n13648) );
  NAND2_X1 U12341 ( .A1(n13409), .A2(n13408), .ZN(n19933) );
  INV_X1 U12342 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19929) );
  OR2_X1 U12343 ( .A1(n19913), .A2(n19903), .ZN(n19905) );
  NAND2_X1 U12344 ( .A1(n12925), .A2(n12924), .ZN(n15579) );
  NAND2_X1 U12345 ( .A1(n19063), .A2(n12931), .ZN(n12925) );
  NAND2_X1 U12346 ( .A1(n13471), .A2(n13470), .ZN(n19923) );
  OR2_X1 U12347 ( .A1(n13469), .A2(n13468), .ZN(n13471) );
  AOI21_X1 U12348 ( .B1(n10093), .B2(n15605), .A(n15604), .ZN(n16323) );
  OR2_X1 U12349 ( .A1(n19306), .A2(n19618), .ZN(n19324) );
  OAI21_X1 U12350 ( .B1(n19367), .B2(n19366), .A(n19365), .ZN(n19385) );
  OR3_X1 U12351 ( .A1(n19422), .A2(n19421), .A3(n19618), .ZN(n19441) );
  OAI21_X1 U12352 ( .B1(n19623), .B2(n19931), .A(n19622), .ZN(n19648) );
  INV_X1 U12353 ( .A(n19802), .ZN(n19699) );
  INV_X1 U12354 ( .A(n19690), .ZN(n19708) );
  INV_X1 U12355 ( .A(n19782), .ZN(n19733) );
  OAI21_X1 U12356 ( .B1(n19723), .B2(n19722), .A(n19721), .ZN(n19748) );
  INV_X1 U12357 ( .A(n19674), .ZN(n19768) );
  INV_X1 U12358 ( .A(n19740), .ZN(n19785) );
  INV_X1 U12359 ( .A(n19249), .ZN(n19791) );
  NAND2_X1 U12360 ( .A1(n19712), .A2(n19756), .ZN(n19801) );
  INV_X1 U12361 ( .A(n19812), .ZN(n19798) );
  AND3_X1 U12362 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n19713), .ZN(n19804) );
  INV_X1 U12363 ( .A(n19801), .ZN(n19808) );
  OR2_X1 U12364 ( .A1(n19652), .A2(n19905), .ZN(n19812) );
  INV_X1 U12365 ( .A(n19260), .ZN(n19807) );
  NOR2_X1 U12366 ( .A1(n16340), .A2(n19931), .ZN(n16362) );
  NAND2_X1 U12367 ( .A1(n18921), .A2(n17418), .ZN(n18919) );
  INV_X1 U12368 ( .A(n18921), .ZN(n18916) );
  NAND2_X1 U12369 ( .A1(n18901), .A2(n18725), .ZN(n17479) );
  NOR2_X1 U12370 ( .A1(n18919), .A2(n18741), .ZN(n16874) );
  INV_X1 U12371 ( .A(n16874), .ZN(n16895) );
  NAND2_X1 U12372 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n16909), .ZN(n16878) );
  NAND4_X1 U12373 ( .A1(n18217), .A2(n18916), .A3(n18755), .A4(n18745), .ZN(
        n16909) );
  NOR2_X1 U12374 ( .A1(n16916), .A2(n16971), .ZN(n16976) );
  INV_X1 U12375 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17252) );
  NOR2_X2 U12376 ( .A1(n18266), .A2(n17079), .ZN(n17257) );
  INV_X1 U12377 ( .A(n17272), .ZN(n17268) );
  NAND2_X1 U12378 ( .A1(n17285), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n17280) );
  NAND2_X1 U12379 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(P3_EAX_REG_25__SCAN_IN), 
        .ZN(n9852) );
  NOR3_X1 U12380 ( .A1(n17299), .A2(n17345), .A3(n9853), .ZN(n17290) );
  NOR3_X1 U12381 ( .A1(n17432), .A2(n17304), .A3(n17311), .ZN(n17300) );
  NOR2_X1 U12382 ( .A1(n17345), .A2(n17304), .ZN(n17338) );
  NOR2_X2 U12383 ( .A1(n18259), .A2(n17407), .ZN(n17337) );
  NOR2_X1 U12384 ( .A1(n17350), .A2(n17531), .ZN(n17340) );
  INV_X1 U12385 ( .A(n18266), .ZN(n17345) );
  NAND2_X1 U12386 ( .A1(n17375), .A2(n9857), .ZN(n17350) );
  AND2_X1 U12387 ( .A1(n17349), .A2(P3_EAX_REG_14__SCAN_IN), .ZN(n9857) );
  NOR2_X1 U12388 ( .A1(n17377), .A2(n17459), .ZN(n17375) );
  INV_X1 U12389 ( .A(n11361), .ZN(n17390) );
  INV_X1 U12390 ( .A(n17410), .ZN(n17402) );
  INV_X2 U12391 ( .A(n17376), .ZN(n17407) );
  NOR2_X1 U12392 ( .A1(n10111), .A2(n10108), .ZN(n10107) );
  NOR2_X1 U12393 ( .A1(n11245), .A2(n9725), .ZN(n10112) );
  OAI21_X1 U12394 ( .B1(n15799), .B2(n18747), .A(n15798), .ZN(n17262) );
  INV_X1 U12395 ( .A(n17405), .ZN(n17411) );
  NOR2_X1 U12396 ( .A1(n18903), .A2(n17446), .ZN(n17442) );
  CLKBUF_X1 U12397 ( .A(n17442), .Z(n17472) );
  NOR2_X1 U12398 ( .A1(n17479), .A2(n18740), .ZN(n17515) );
  CLKBUF_X1 U12399 ( .A(n17518), .Z(n17527) );
  NOR2_X1 U12400 ( .A1(n17527), .A2(n18906), .ZN(n17528) );
  NOR2_X1 U12401 ( .A1(n17911), .A2(n11482), .ZN(n16400) );
  INV_X1 U12402 ( .A(n10125), .ZN(n17535) );
  NOR2_X1 U12403 ( .A1(n17651), .A2(n17652), .ZN(n17641) );
  AND3_X1 U12404 ( .A1(n17794), .A2(n9682), .A3(n9744), .ZN(n17672) );
  NOR2_X1 U12405 ( .A1(n17689), .A2(n9946), .ZN(n9945) );
  INV_X1 U12406 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n9946) );
  AND3_X1 U12407 ( .A1(n17794), .A2(n9682), .A3(n9947), .ZN(n17711) );
  INV_X1 U12408 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17827) );
  NAND2_X1 U12409 ( .A1(n18525), .A2(n18585), .ZN(n18263) );
  INV_X1 U12410 ( .A(n17901), .ZN(n17888) );
  AND2_X1 U12411 ( .A1(n11272), .A2(n9934), .ZN(n17567) );
  OAI21_X1 U12412 ( .B1(n18045), .B2(n18020), .A(n18196), .ZN(n18120) );
  INV_X1 U12413 ( .A(n17804), .ZN(n18138) );
  NAND2_X1 U12414 ( .A1(n10117), .A2(n10119), .ZN(n17825) );
  NAND2_X1 U12415 ( .A1(n17836), .A2(n10120), .ZN(n10117) );
  INV_X1 U12416 ( .A(n9806), .ZN(n17839) );
  NAND2_X1 U12417 ( .A1(n17836), .A2(n17835), .ZN(n17834) );
  NOR2_X1 U12418 ( .A1(n15707), .A2(n18694), .ZN(n18703) );
  INV_X1 U12419 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18707) );
  INV_X1 U12420 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18714) );
  AOI211_X1 U12421 ( .C1(n18901), .C2(n18734), .A(n18233), .B(n15711), .ZN(
        n18888) );
  INV_X1 U12422 ( .A(n16893), .ZN(n18755) );
  NOR2_X1 U12425 ( .A1(n9835), .A2(n9830), .ZN(n14252) );
  INV_X1 U12426 ( .A(n14251), .ZN(n9835) );
  NAND2_X1 U12427 ( .A1(n9834), .A2(n9831), .ZN(n9830) );
  NOR2_X1 U12428 ( .A1(n20008), .A2(n20804), .ZN(n14222) );
  INV_X1 U12429 ( .A(n12586), .ZN(n12587) );
  OAI21_X1 U12430 ( .B1(n14743), .B2(n20172), .A(n12585), .ZN(n12586) );
  INV_X1 U12431 ( .A(n14705), .ZN(n14734) );
  OAI21_X1 U12432 ( .B1(n14755), .B2(n20208), .A(n10062), .ZN(P1_U3003) );
  NOR2_X1 U12433 ( .A1(n10063), .A2(n14756), .ZN(n10062) );
  AND2_X1 U12434 ( .A1(n14765), .A2(n14757), .ZN(n10063) );
  OAI21_X1 U12435 ( .B1(n14762), .B2(n20208), .A(n9733), .ZN(P1_U3004) );
  AND2_X1 U12436 ( .A1(n14765), .A2(n14764), .ZN(n9914) );
  OR2_X1 U12437 ( .A1(n14086), .A2(n9779), .ZN(n10094) );
  AND2_X1 U12438 ( .A1(n13210), .A2(n13209), .ZN(n13211) );
  INV_X1 U12439 ( .A(n10093), .ZN(n13709) );
  AND2_X1 U12440 ( .A1(n10098), .A2(n10096), .ZN(n16225) );
  AOI21_X1 U12441 ( .B1(n16302), .B2(n11014), .A(n10097), .ZN(n10096) );
  AOI21_X1 U12442 ( .B1(n19073), .B2(n19202), .A(n10100), .ZN(n10099) );
  NAND2_X1 U12443 ( .A1(n15296), .A2(n19204), .ZN(n10102) );
  OAI21_X1 U12444 ( .B1(n15300), .B2(n16306), .A(n10053), .ZN(n15304) );
  INV_X1 U12445 ( .A(n10054), .ZN(n10053) );
  OAI21_X1 U12446 ( .B1(n15308), .B2(n19206), .A(n10208), .ZN(n15315) );
  AOI21_X1 U12447 ( .B1(n15310), .B2(n19202), .A(n10209), .ZN(n10208) );
  OAI21_X1 U12448 ( .B1(n15460), .B2(n9693), .A(n9734), .ZN(P2_U3029) );
  AOI21_X1 U12449 ( .B1(n16303), .B2(n10093), .A(n10095), .ZN(n16304) );
  AND2_X1 U12450 ( .A1(n11497), .A2(n11496), .ZN(n11498) );
  OR2_X1 U12451 ( .A1(n11481), .A2(n18218), .ZN(n9808) );
  NAND2_X1 U12452 ( .A1(n11501), .A2(n18134), .ZN(n9809) );
  AOI21_X1 U12453 ( .B1(n10123), .B2(n10122), .A(n9647), .ZN(n11459) );
  INV_X2 U12454 ( .A(n17040), .ZN(n11207) );
  INV_X1 U12455 ( .A(n11587), .ZN(n12258) );
  AND2_X1 U12456 ( .A1(n11513), .A2(n11511), .ZN(n11664) );
  OR2_X1 U12457 ( .A1(n14361), .A2(n10269), .ZN(n14322) );
  AND2_X1 U12458 ( .A1(n9825), .A2(n13980), .ZN(n9679) );
  AND2_X1 U12459 ( .A1(n10996), .A2(n10998), .ZN(n9680) );
  AND4_X1 U12460 ( .A1(n11575), .A2(n11574), .A3(n11573), .A4(n11572), .ZN(
        n9681) );
  NAND2_X1 U12461 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10320), .ZN(
        n10423) );
  INV_X2 U12462 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n9877) );
  AND2_X1 U12463 ( .A1(n17755), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9682) );
  NOR2_X1 U12464 ( .A1(n10253), .A2(n10258), .ZN(n14399) );
  OR2_X1 U12465 ( .A1(n12648), .A2(n10182), .ZN(n9683) );
  NOR2_X1 U12466 ( .A1(n10253), .A2(n10256), .ZN(n14458) );
  NOR2_X1 U12467 ( .A1(n14361), .A2(n14444), .ZN(n9684) );
  AND3_X1 U12468 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12658) );
  NOR2_X1 U12469 ( .A1(n14387), .A2(n14388), .ZN(n9685) );
  OR2_X1 U12470 ( .A1(n11009), .A2(n9984), .ZN(n9686) );
  NAND2_X1 U12471 ( .A1(n10285), .A2(n15394), .ZN(n9687) );
  AND2_X1 U12472 ( .A1(n15569), .A2(n10013), .ZN(n9688) );
  NAND2_X1 U12473 ( .A1(n14697), .A2(n12571), .ZN(n14667) );
  AND4_X1 U12474 ( .A1(n11596), .A2(n11595), .A3(n11594), .A4(n11593), .ZN(
        n9689) );
  AND4_X1 U12475 ( .A1(n11569), .A2(n11568), .A3(n11567), .A4(n11566), .ZN(
        n9690) );
  INV_X1 U12476 ( .A(n11588), .ZN(n13803) );
  INV_X1 U12477 ( .A(n10268), .ZN(n14337) );
  AND2_X1 U12478 ( .A1(n14565), .A2(n9920), .ZN(n9692) );
  INV_X1 U12479 ( .A(n12571), .ZN(n9998) );
  AND2_X1 U12480 ( .A1(n15464), .A2(n15461), .ZN(n9693) );
  INV_X1 U12481 ( .A(n17409), .ZN(n11369) );
  OR2_X1 U12482 ( .A1(n9686), .A2(n9980), .ZN(n9694) );
  NOR2_X1 U12483 ( .A1(n14662), .A2(n9785), .ZN(n9695) );
  AND2_X1 U12484 ( .A1(n10202), .A2(n13858), .ZN(n9696) );
  AND2_X1 U12485 ( .A1(n10792), .A2(n10013), .ZN(n9697) );
  NOR2_X1 U12486 ( .A1(n14126), .A2(n14125), .ZN(n9698) );
  NAND2_X1 U12487 ( .A1(n10987), .A2(n14014), .ZN(n9699) );
  NAND2_X1 U12488 ( .A1(n10237), .A2(n13750), .ZN(n13752) );
  OR2_X1 U12489 ( .A1(n13861), .A2(n10224), .ZN(n13899) );
  NAND2_X1 U12490 ( .A1(n15004), .A2(n10234), .ZN(n14990) );
  NOR3_X1 U12491 ( .A1(n12622), .A2(n13243), .A3(n15149), .ZN(n12620) );
  AND2_X1 U12492 ( .A1(n13901), .A2(n9768), .ZN(n14171) );
  AND2_X1 U12493 ( .A1(n9950), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9700) );
  OR2_X1 U12494 ( .A1(n14922), .A2(n10043), .ZN(n9701) );
  AND2_X1 U12495 ( .A1(n10198), .A2(n10197), .ZN(n9702) );
  OR3_X1 U12496 ( .A1(n14476), .A2(n10075), .A3(n10078), .ZN(n9703) );
  AND2_X1 U12497 ( .A1(n12909), .A2(n12908), .ZN(n9704) );
  NAND2_X1 U12498 ( .A1(n13725), .A2(n11576), .ZN(n13298) );
  INV_X1 U12499 ( .A(n13298), .ZN(n9956) );
  AND2_X1 U12500 ( .A1(n13750), .A2(n9780), .ZN(n9705) );
  AND2_X1 U12501 ( .A1(n9702), .A2(n13273), .ZN(n9706) );
  AND2_X1 U12502 ( .A1(n10167), .A2(n10166), .ZN(n9707) );
  AND2_X1 U12503 ( .A1(n10046), .A2(n10045), .ZN(n9708) );
  AND2_X1 U12504 ( .A1(n9707), .A2(n11096), .ZN(n9709) );
  AND2_X1 U12505 ( .A1(n10105), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9710) );
  NAND2_X2 U12506 ( .A1(n19974), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n19884) );
  AND2_X2 U12507 ( .A1(n10328), .A2(n10318), .ZN(n10319) );
  INV_X1 U12508 ( .A(n11112), .ZN(n10635) );
  OR3_X1 U12509 ( .A1(n15068), .A2(n10057), .A3(n12880), .ZN(n9711) );
  OR3_X1 U12510 ( .A1(n17299), .A2(n17345), .A3(n9852), .ZN(n9712) );
  AND2_X1 U12511 ( .A1(n13187), .A2(n10510), .ZN(n10720) );
  OR3_X1 U12512 ( .A1(n16896), .A2(n18872), .A3(n18860), .ZN(n9713) );
  OR2_X1 U12513 ( .A1(n14441), .A2(n10079), .ZN(n9714) );
  AND2_X1 U12514 ( .A1(n12547), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9715) );
  OR2_X1 U12515 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n10916), .ZN(n9716) );
  NAND2_X1 U12516 ( .A1(n10654), .A2(n10662), .ZN(n10653) );
  NAND2_X1 U12517 ( .A1(n10183), .A2(n9636), .ZN(n12653) );
  NAND2_X1 U12518 ( .A1(n10858), .A2(n10857), .ZN(n15474) );
  NOR2_X1 U12519 ( .A1(n12648), .A2(n16191), .ZN(n12649) );
  NOR2_X1 U12520 ( .A1(n12648), .A2(n10181), .ZN(n12647) );
  AND2_X1 U12521 ( .A1(n14287), .A2(n10070), .ZN(n9718) );
  NAND2_X1 U12522 ( .A1(n10575), .A2(n13617), .ZN(n10609) );
  INV_X1 U12523 ( .A(n9935), .ZN(n17394) );
  AND2_X1 U12524 ( .A1(n17285), .A2(n9851), .ZN(n9719) );
  NOR2_X1 U12525 ( .A1(n15125), .A2(n10281), .ZN(n9720) );
  AND2_X1 U12526 ( .A1(n10602), .A2(n10630), .ZN(n10654) );
  AND2_X1 U12527 ( .A1(n13147), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12923) );
  AND2_X1 U12528 ( .A1(n16192), .A2(n15411), .ZN(n9721) );
  NOR2_X1 U12529 ( .A1(n14375), .A2(n14446), .ZN(n14360) );
  INV_X1 U12530 ( .A(n10573), .ZN(n12668) );
  AND2_X1 U12531 ( .A1(n15837), .A2(n12465), .ZN(n9722) );
  NOR2_X1 U12532 ( .A1(n13319), .A2(n13654), .ZN(n9723) );
  BUF_X1 U12533 ( .A(n10559), .Z(n12904) );
  NAND2_X1 U12534 ( .A1(n9957), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11677) );
  AND2_X1 U12535 ( .A1(n14661), .A2(n10146), .ZN(n9724) );
  AND2_X1 U12536 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n9725) );
  INV_X1 U12537 ( .A(n14557), .ZN(n10253) );
  INV_X1 U12538 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12656) );
  OR2_X1 U12539 ( .A1(n17053), .A2(n11221), .ZN(n9726) );
  INV_X1 U12540 ( .A(n20227), .ZN(n11604) );
  INV_X1 U12541 ( .A(n13654), .ZN(n20212) );
  AND4_X1 U12542 ( .A1(n11592), .A2(n11591), .A3(n11590), .A4(n11589), .ZN(
        n9727) );
  AND2_X1 U12543 ( .A1(n10689), .A2(n13648), .ZN(n10741) );
  INV_X1 U12544 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10517) );
  AND3_X1 U12545 ( .A1(n9996), .A2(n9723), .A3(n20220), .ZN(n9728) );
  AND2_X1 U12546 ( .A1(n14282), .A2(n10260), .ZN(n14256) );
  OR2_X1 U12547 ( .A1(n15068), .A2(n13248), .ZN(n9729) );
  OR2_X1 U12548 ( .A1(n14361), .A2(n10271), .ZN(n10268) );
  OR2_X1 U12549 ( .A1(n15068), .A2(n10057), .ZN(n9730) );
  NAND2_X1 U12550 ( .A1(n10130), .A2(n9999), .ZN(n14697) );
  AND2_X1 U12551 ( .A1(n15170), .A2(n10939), .ZN(n9731) );
  AND2_X1 U12552 ( .A1(n10092), .A2(n10594), .ZN(n9732) );
  INV_X1 U12553 ( .A(n14820), .ZN(n13561) );
  AND3_X2 U12554 ( .A1(n10314), .A2(n11565), .A3(n11564), .ZN(n14820) );
  INV_X1 U12555 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11687) );
  NOR2_X1 U12556 ( .A1(n14763), .A2(n9914), .ZN(n9733) );
  NOR2_X1 U12557 ( .A1(n12670), .A2(n19220), .ZN(n10574) );
  INV_X1 U12558 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9913) );
  NAND2_X1 U12559 ( .A1(n10861), .A2(n9707), .ZN(n10169) );
  AND2_X1 U12560 ( .A1(n9978), .A2(n9975), .ZN(n9734) );
  INV_X1 U12561 ( .A(n15567), .ZN(n9973) );
  AND2_X1 U12562 ( .A1(n10995), .A2(n10994), .ZN(n15567) );
  NAND2_X1 U12563 ( .A1(n15175), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15161) );
  INV_X1 U12564 ( .A(n15161), .ZN(n9882) );
  INV_X1 U12565 ( .A(n11237), .ZN(n11238) );
  AND2_X1 U12566 ( .A1(n10014), .A2(n10792), .ZN(n9735) );
  INV_X1 U12567 ( .A(n11786), .ZN(n11813) );
  INV_X1 U12568 ( .A(n15566), .ZN(n9974) );
  NAND2_X1 U12569 ( .A1(n9868), .A2(n9867), .ZN(n15566) );
  OR2_X1 U12570 ( .A1(n9720), .A2(n10280), .ZN(n9736) );
  AND3_X1 U12571 ( .A1(n11223), .A2(n9937), .A3(n9936), .ZN(n9737) );
  INV_X1 U12572 ( .A(n11153), .ZN(n16896) );
  NOR2_X1 U12573 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11153) );
  AND2_X1 U12574 ( .A1(n10148), .A2(n9720), .ZN(n9738) );
  AND2_X1 U12575 ( .A1(n10881), .A2(n10157), .ZN(n9739) );
  NOR2_X1 U12576 ( .A1(n14662), .A2(n12574), .ZN(n9740) );
  AND2_X1 U12577 ( .A1(n16021), .A2(n16022), .ZN(n9741) );
  NOR2_X1 U12578 ( .A1(n16069), .A2(n18993), .ZN(n9742) );
  AND2_X1 U12579 ( .A1(n10812), .A2(n10811), .ZN(n11002) );
  INV_X1 U12580 ( .A(n11002), .ZN(n10013) );
  INV_X1 U12581 ( .A(n15394), .ZN(n10284) );
  NAND2_X1 U12582 ( .A1(n20220), .A2(n9922), .ZN(n9743) );
  AND2_X1 U12583 ( .A1(n9947), .A2(n9945), .ZN(n9744) );
  AND2_X1 U12584 ( .A1(n9918), .A2(n9846), .ZN(n9745) );
  INV_X1 U12585 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13576) );
  INV_X1 U12586 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16214) );
  INV_X1 U12587 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18860) );
  INV_X1 U12588 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18880) );
  INV_X2 U12589 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18872) );
  AND2_X1 U12590 ( .A1(n13454), .A2(n12672), .ZN(n12794) );
  INV_X1 U12591 ( .A(n9924), .ZN(n13305) );
  NOR2_X1 U12592 ( .A1(n9994), .A2(n9993), .ZN(n12342) );
  OR2_X1 U12593 ( .A1(n12729), .A2(n12728), .ZN(n13862) );
  NAND2_X1 U12594 ( .A1(n9826), .A2(n9679), .ZN(n13979) );
  NAND2_X1 U12595 ( .A1(n12579), .A2(n11599), .ZN(n13297) );
  AND2_X1 U12596 ( .A1(n14148), .A2(n14193), .ZN(n14191) );
  NAND2_X1 U12597 ( .A1(n15004), .A2(n12991), .ZN(n14994) );
  NAND2_X1 U12598 ( .A1(n9915), .A2(n11705), .ZN(n10245) );
  AND2_X1 U12599 ( .A1(n15004), .A2(n10232), .ZN(n14984) );
  NOR2_X1 U12600 ( .A1(n15518), .A2(n15500), .ZN(n15484) );
  INV_X1 U12601 ( .A(n9804), .ZN(n17762) );
  OR2_X1 U12602 ( .A1(n17801), .A2(n11388), .ZN(n9804) );
  AND2_X1 U12603 ( .A1(n11684), .A2(n12569), .ZN(n9747) );
  OR2_X1 U12604 ( .A1(n10050), .A2(n14134), .ZN(n9748) );
  AND2_X1 U12605 ( .A1(n10207), .A2(n14020), .ZN(n9749) );
  NAND2_X1 U12606 ( .A1(n11747), .A2(n11746), .ZN(n11825) );
  AND2_X1 U12607 ( .A1(n14909), .A2(n9702), .ZN(n9750) );
  INV_X1 U12608 ( .A(n15200), .ZN(n9903) );
  AND2_X1 U12609 ( .A1(n13260), .A2(n9708), .ZN(n9751) );
  INV_X1 U12610 ( .A(n10880), .ZN(n10158) );
  NOR2_X1 U12611 ( .A1(n14977), .A2(n14979), .ZN(n14978) );
  OR2_X1 U12612 ( .A1(n13773), .A2(n9926), .ZN(n9752) );
  OR3_X1 U12613 ( .A1(n14441), .A2(n10082), .A3(n10084), .ZN(n9753) );
  AND3_X1 U12614 ( .A1(n20873), .A2(n12569), .A3(n12568), .ZN(n9754) );
  NAND2_X1 U12615 ( .A1(n10817), .A2(n10816), .ZN(n15260) );
  NOR2_X1 U12616 ( .A1(n13065), .A2(n14978), .ZN(n9755) );
  AND2_X1 U12617 ( .A1(n10292), .A2(n10293), .ZN(n9756) );
  AND2_X1 U12618 ( .A1(n13547), .A2(n9926), .ZN(n9757) );
  OR2_X1 U12619 ( .A1(n15485), .A2(n9701), .ZN(n9758) );
  AND2_X1 U12620 ( .A1(n10847), .A2(n10153), .ZN(n9759) );
  AND2_X1 U12621 ( .A1(n14882), .A2(n14881), .ZN(n13260) );
  AND2_X1 U12622 ( .A1(n10156), .A2(n10155), .ZN(n9760) );
  INV_X1 U12623 ( .A(n14167), .ZN(n12940) );
  OR2_X1 U12624 ( .A1(n12806), .A2(n12805), .ZN(n14167) );
  AND2_X1 U12625 ( .A1(n10261), .A2(n9829), .ZN(n9761) );
  INV_X1 U12626 ( .A(n9986), .ZN(n10135) );
  NAND2_X1 U12627 ( .A1(n9987), .A2(n12566), .ZN(n9986) );
  AND2_X1 U12628 ( .A1(n12711), .A2(n12710), .ZN(n9762) );
  INV_X1 U12629 ( .A(n12402), .ZN(n10078) );
  NOR2_X1 U12630 ( .A1(n14024), .A2(n14023), .ZN(n9763) );
  AND2_X1 U12631 ( .A1(n9763), .A2(n10223), .ZN(n9764) );
  INV_X1 U12632 ( .A(n13878), .ZN(n12939) );
  OR2_X1 U12633 ( .A1(n12743), .A2(n12742), .ZN(n13878) );
  NAND2_X1 U12634 ( .A1(n13647), .A2(n13646), .ZN(n13645) );
  NOR2_X1 U12635 ( .A1(n13281), .A2(n18993), .ZN(n9765) );
  NAND2_X1 U12636 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n11363), .ZN(
        n9766) );
  AND2_X1 U12637 ( .A1(n10246), .A2(n11825), .ZN(n9767) );
  AND2_X1 U12638 ( .A1(n9749), .A2(n10206), .ZN(n9768) );
  OR2_X1 U12639 ( .A1(n12522), .A2(n12496), .ZN(n9769) );
  AND2_X1 U12640 ( .A1(n9970), .A2(n9969), .ZN(n9770) );
  AND2_X1 U12641 ( .A1(n12008), .A2(n11992), .ZN(n9771) );
  AND2_X1 U12642 ( .A1(n9871), .A2(n14014), .ZN(n9772) );
  INV_X1 U12643 ( .A(n13943), .ZN(n10039) );
  OR2_X1 U12644 ( .A1(n12709), .A2(n12708), .ZN(n13943) );
  NOR2_X1 U12645 ( .A1(n13861), .A2(n12939), .ZN(n9773) );
  INV_X1 U12646 ( .A(n12188), .ZN(n11570) );
  INV_X1 U12647 ( .A(n12275), .ZN(n12056) );
  INV_X1 U12648 ( .A(n12056), .ZN(n12350) );
  INV_X1 U12649 ( .A(n11971), .ZN(n11955) );
  AND2_X1 U12650 ( .A1(n17641), .A2(n9950), .ZN(n9774) );
  INV_X1 U12651 ( .A(n13628), .ZN(n10037) );
  INV_X1 U12652 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n9951) );
  AND2_X1 U12653 ( .A1(n13618), .A2(n19943), .ZN(n16309) );
  AND2_X1 U12654 ( .A1(n10237), .A2(n9705), .ZN(n13762) );
  OR2_X1 U12655 ( .A1(n13860), .A2(n12938), .ZN(n13861) );
  OR2_X1 U12656 ( .A1(n13860), .A2(n9968), .ZN(n14022) );
  NOR2_X1 U12657 ( .A1(n16289), .A2(n14114), .ZN(n14113) );
  AND2_X1 U12658 ( .A1(n14253), .A2(n14269), .ZN(n9775) );
  AND2_X1 U12659 ( .A1(n10037), .A2(n10038), .ZN(n9776) );
  AND2_X1 U12660 ( .A1(n10037), .A2(n10033), .ZN(n9777) );
  NAND2_X1 U12661 ( .A1(n16291), .A2(n16290), .ZN(n16289) );
  NAND2_X1 U12662 ( .A1(n13755), .A2(n13754), .ZN(n13757) );
  NAND2_X1 U12663 ( .A1(n13851), .A2(n11811), .ZN(n13884) );
  NAND2_X1 U12664 ( .A1(n13704), .A2(n12935), .ZN(n13748) );
  OR3_X1 U12665 ( .A1(n13087), .A2(n13086), .A3(n14970), .ZN(n9778) );
  AND2_X1 U12666 ( .A1(n10093), .A2(n19062), .ZN(n9779) );
  INV_X1 U12667 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11787) );
  INV_X1 U12668 ( .A(n10903), .ZN(n10168) );
  INV_X1 U12669 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n16055) );
  INV_X1 U12670 ( .A(n9925), .ZN(n15727) );
  NOR3_X1 U12671 ( .A1(n14476), .A2(n10075), .A3(n10074), .ZN(n10073) );
  OR2_X1 U12672 ( .A1(n12838), .A2(n12837), .ZN(n15028) );
  INV_X1 U12673 ( .A(n15028), .ZN(n12941) );
  OAI21_X1 U12674 ( .B1(n12521), .B2(n11790), .A(n9822), .ZN(n13849) );
  AND2_X1 U12675 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9780) );
  NAND2_X1 U12676 ( .A1(n11607), .A2(n10309), .ZN(n13543) );
  INV_X1 U12677 ( .A(n13543), .ZN(n9953) );
  OR2_X1 U12678 ( .A1(n12622), .A2(n13243), .ZN(n9781) );
  INV_X1 U12679 ( .A(n10071), .ZN(n10070) );
  NAND2_X1 U12680 ( .A1(n10072), .A2(n9775), .ZN(n10071) );
  OR2_X1 U12681 ( .A1(n11468), .A2(n10126), .ZN(n9782) );
  NOR2_X1 U12682 ( .A1(n14085), .A2(n10094), .ZN(n9783) );
  AND2_X1 U12683 ( .A1(n10070), .A2(n12482), .ZN(n9784) );
  INV_X1 U12684 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10175) );
  INV_X1 U12685 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n9952) );
  OR2_X1 U12686 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n12574), .ZN(
        n9785) );
  AND2_X1 U12687 ( .A1(n12849), .A2(n12848), .ZN(n9786) );
  NAND2_X1 U12688 ( .A1(n10559), .A2(n10556), .ZN(n13455) );
  INV_X1 U12689 ( .A(n13455), .ZN(n9887) );
  INV_X1 U12690 ( .A(n9958), .ZN(n13335) );
  NAND2_X1 U12691 ( .A1(n9953), .A2(n9956), .ZN(n9958) );
  OR2_X1 U12692 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n9787) );
  AND2_X1 U12693 ( .A1(n9955), .A2(n12594), .ZN(n9788) );
  OR2_X1 U12694 ( .A1(n9785), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9789) );
  INV_X1 U12695 ( .A(n15411), .ZN(n9984) );
  INV_X1 U12696 ( .A(n15423), .ZN(n9980) );
  AND2_X1 U12697 ( .A1(n9877), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12931) );
  INV_X1 U12698 ( .A(n12931), .ZN(n10230) );
  INV_X1 U12699 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10166) );
  INV_X1 U12700 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n9943) );
  INV_X1 U12701 ( .A(n14724), .ZN(n9920) );
  INV_X1 U12702 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n9853) );
  AND2_X1 U12703 ( .A1(n9851), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n9790) );
  OR2_X1 U12704 ( .A1(n14577), .A2(n10060), .ZN(n9791) );
  NAND2_X2 U12705 ( .A1(n18918), .A2(n16528), .ZN(n18217) );
  OAI22_X2 U12706 ( .A1(n14237), .A2(n20248), .B1(n21027), .B2(n20247), .ZN(
        n20698) );
  OAI22_X2 U12707 ( .A1(n16426), .A2(n20248), .B1(n20959), .B2(n20247), .ZN(
        n20734) );
  OAI22_X2 U12708 ( .A1(n21033), .A2(n20247), .B1(n20219), .B2(n20248), .ZN(
        n20728) );
  NAND2_X1 U12709 ( .A1(n20154), .A2(n14547), .ZN(n20248) );
  OAI22_X2 U12710 ( .A1(n20933), .A2(n20247), .B1(n20211), .B2(n20248), .ZN(
        n20722) );
  OAI22_X2 U12711 ( .A1(n20239), .A2(n20247), .B1(n20238), .B2(n20248), .ZN(
        n20752) );
  OAI22_X2 U12712 ( .A1(n20226), .A2(n20248), .B1(n20922), .B2(n20247), .ZN(
        n20688) );
  OAI22_X2 U12713 ( .A1(n20234), .A2(n20248), .B1(n20233), .B2(n20247), .ZN(
        n20694) );
  OAI22_X2 U12714 ( .A1(n14494), .A2(n20248), .B1(n21014), .B2(n20247), .ZN(
        n20684) );
  NAND2_X1 U12715 ( .A1(n10137), .A2(n9997), .ZN(n15896) );
  NAND2_X2 U12716 ( .A1(n10128), .A2(n11598), .ZN(n13571) );
  NAND2_X2 U12717 ( .A1(n10698), .A2(n10697), .ZN(n10765) );
  NAND2_X1 U12718 ( .A1(n11001), .A2(n11000), .ZN(n15258) );
  NAND2_X2 U12719 ( .A1(n17675), .A2(n17737), .ZN(n17636) );
  NAND2_X2 U12720 ( .A1(n17676), .A2(n18016), .ZN(n17675) );
  AND2_X2 U12721 ( .A1(n9795), .A2(n9793), .ZN(n17676) );
  XNOR2_X2 U12722 ( .A(n11264), .B(n18130), .ZN(n17804) );
  NAND2_X2 U12723 ( .A1(n11265), .A2(n17803), .ZN(n17736) );
  OR2_X2 U12724 ( .A1(n17537), .A2(n9782), .ZN(n10125) );
  INV_X2 U12725 ( .A(n11276), .ZN(n17553) );
  OR2_X2 U12726 ( .A1(n11275), .A2(n17918), .ZN(n11276) );
  NAND3_X1 U12727 ( .A1(n9934), .A2(n11272), .A3(n17925), .ZN(n9799) );
  NOR2_X2 U12728 ( .A1(n11155), .A2(n11151), .ZN(n17210) );
  NAND3_X1 U12729 ( .A1(n9803), .A2(n11153), .A3(
        P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n9801) );
  NAND3_X1 U12730 ( .A1(n9809), .A2(n11488), .A3(n9808), .ZN(P3_U2831) );
  AND2_X2 U12731 ( .A1(n13672), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11587) );
  NAND2_X1 U12732 ( .A1(n13561), .A2(n11610), .ZN(n9812) );
  NAND3_X1 U12733 ( .A1(n20256), .A2(n11704), .A3(n16055), .ZN(n9814) );
  NAND2_X1 U12734 ( .A1(n11682), .A2(n11683), .ZN(n20256) );
  NAND3_X1 U12735 ( .A1(n11686), .A2(n9819), .A3(n9815), .ZN(n11792) );
  OR2_X2 U12736 ( .A1(n11659), .A2(n9821), .ZN(n9815) );
  NAND2_X1 U12737 ( .A1(n11659), .A2(n9820), .ZN(n11686) );
  INV_X1 U12738 ( .A(n11674), .ZN(n9821) );
  INV_X1 U12739 ( .A(n14387), .ZN(n9824) );
  NAND2_X1 U12740 ( .A1(n9824), .A2(n9771), .ZN(n14375) );
  NAND3_X1 U12741 ( .A1(n9826), .A2(n9698), .A3(n9679), .ZN(n14124) );
  INV_X1 U12742 ( .A(n13964), .ZN(n9825) );
  NOR2_X1 U12743 ( .A1(n14297), .A2(n9827), .ZN(n12589) );
  NAND3_X1 U12744 ( .A1(n10064), .A2(n11586), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11724) );
  INV_X1 U12745 ( .A(n15837), .ZN(n15854) );
  NAND2_X1 U12746 ( .A1(n13326), .A2(n11611), .ZN(n13542) );
  AND2_X4 U12747 ( .A1(n20227), .A2(n9926), .ZN(n13412) );
  NAND2_X2 U12748 ( .A1(n9681), .A2(n9690), .ZN(n20227) );
  AND2_X1 U12749 ( .A1(n14793), .A2(n9843), .ZN(n9842) );
  NAND2_X2 U12750 ( .A1(n9990), .A2(n9841), .ZN(n14662) );
  NAND3_X1 U12751 ( .A1(n14697), .A2(n12505), .A3(n9842), .ZN(n9841) );
  NAND3_X1 U12752 ( .A1(n11812), .A2(n11825), .A3(n13866), .ZN(n9844) );
  NAND2_X1 U12753 ( .A1(n12577), .A2(n9692), .ZN(n9846) );
  NAND2_X1 U12754 ( .A1(n12577), .A2(n9848), .ZN(n9847) );
  OAI21_X2 U12755 ( .B1(n9918), .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n9847), .ZN(n13221) );
  NAND2_X1 U12756 ( .A1(n17285), .A2(n9790), .ZN(n17272) );
  NOR2_X1 U12757 ( .A1(n17299), .A2(n17345), .ZN(n17296) );
  INV_X1 U12758 ( .A(n17290), .ZN(n17295) );
  NAND4_X1 U12759 ( .A1(n9864), .A2(n9863), .A3(n9862), .A4(n9861), .ZN(n9860)
         );
  NAND2_X1 U12760 ( .A1(n13999), .A2(n9772), .ZN(n9867) );
  NAND2_X1 U12761 ( .A1(n9869), .A2(n16216), .ZN(n9868) );
  NAND2_X1 U12762 ( .A1(n9870), .A2(n9699), .ZN(n9869) );
  NAND2_X1 U12763 ( .A1(n13999), .A2(n9871), .ZN(n9870) );
  NAND3_X1 U12764 ( .A1(n10574), .A2(n10584), .A3(n9872), .ZN(n9875) );
  OAI211_X1 U12765 ( .C1(n10585), .C2(n9877), .A(n9876), .B(n9875), .ZN(n10586) );
  NAND2_X1 U12766 ( .A1(n13450), .A2(n9878), .ZN(n10585) );
  NAND3_X1 U12767 ( .A1(n9881), .A2(n9880), .A3(n9879), .ZN(n15269) );
  NAND3_X1 U12768 ( .A1(n9974), .A2(n9973), .A3(n10997), .ZN(n9879) );
  NAND2_X1 U12769 ( .A1(n15269), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11001) );
  AND2_X2 U12770 ( .A1(n9889), .A2(n10552), .ZN(n10593) );
  NAND2_X1 U12771 ( .A1(n15259), .A2(n10291), .ZN(n10028) );
  NAND2_X2 U12772 ( .A1(n10817), .A2(n9890), .ZN(n15259) );
  NAND2_X2 U12773 ( .A1(n11020), .A2(n9894), .ZN(n12910) );
  NAND3_X1 U12774 ( .A1(n10644), .A2(n10643), .A3(n10231), .ZN(n11020) );
  NAND2_X2 U12775 ( .A1(n10018), .A2(n10642), .ZN(n10643) );
  NAND2_X2 U12776 ( .A1(n10017), .A2(n10658), .ZN(n10644) );
  OR2_X1 U12777 ( .A1(n16153), .A2(n16151), .ZN(n9897) );
  INV_X1 U12778 ( .A(n9994), .ZN(n9992) );
  OAI211_X1 U12779 ( .C1(n9909), .C2(n9907), .A(n9906), .B(n9904), .ZN(n11678)
         );
  INV_X1 U12780 ( .A(n9905), .ZN(n9904) );
  OAI21_X1 U12781 ( .B1(n11619), .B2(n11514), .A(n11676), .ZN(n9905) );
  NAND2_X1 U12782 ( .A1(n11618), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9910) );
  INV_X1 U12783 ( .A(n9908), .ZN(n9907) );
  INV_X1 U12784 ( .A(n9957), .ZN(n9909) );
  NAND3_X1 U12785 ( .A1(n11677), .A2(n11619), .A3(n9910), .ZN(n11691) );
  NAND2_X1 U12786 ( .A1(n9912), .A2(n12517), .ZN(n12518) );
  NAND2_X2 U12787 ( .A1(n15896), .A2(n12558), .ZN(n15893) );
  NAND3_X1 U12788 ( .A1(n9915), .A2(n11705), .A3(n16055), .ZN(n10244) );
  XNOR2_X1 U12789 ( .A(n9915), .B(n20347), .ZN(n13800) );
  INV_X1 U12790 ( .A(n12577), .ZN(n14590) );
  INV_X2 U12791 ( .A(n9926), .ZN(n20220) );
  NAND2_X1 U12792 ( .A1(n9926), .A2(n20871), .ZN(n13772) );
  NAND2_X1 U12793 ( .A1(n9926), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n12458) );
  NAND2_X1 U12794 ( .A1(n20220), .A2(n20871), .ZN(n9923) );
  AND2_X1 U12795 ( .A1(n9926), .A2(n13654), .ZN(n13717) );
  NAND2_X1 U12796 ( .A1(n11600), .A2(n9926), .ZN(n9924) );
  NAND2_X1 U12797 ( .A1(n20212), .A2(n9926), .ZN(n13927) );
  NAND2_X1 U12798 ( .A1(n12335), .A2(n9926), .ZN(n12288) );
  NAND2_X1 U12799 ( .A1(n15752), .A2(n9926), .ZN(n9955) );
  NAND2_X1 U12800 ( .A1(n12342), .A2(n9926), .ZN(n9925) );
  OAI22_X1 U12801 ( .A1(n9958), .A2(n13336), .B1(n13420), .B2(n9926), .ZN(
        n13337) );
  XNOR2_X2 U12802 ( .A(n11719), .B(n11718), .ZN(n11812) );
  NAND2_X1 U12803 ( .A1(n9927), .A2(n10313), .ZN(n14637) );
  NOR2_X2 U12804 ( .A1(n15714), .A2(n16389), .ZN(n11469) );
  NAND2_X1 U12805 ( .A1(n17575), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9934) );
  NAND4_X1 U12806 ( .A1(n9940), .A2(n11220), .A3(n11219), .A4(n9737), .ZN(
        n9935) );
  NAND3_X1 U12807 ( .A1(n18056), .A2(n9943), .A3(n9942), .ZN(n9941) );
  NAND2_X2 U12808 ( .A1(n17810), .A2(n11261), .ZN(n11264) );
  XNOR2_X2 U12809 ( .A(n16374), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16846) );
  NAND4_X1 U12810 ( .A1(n17794), .A2(n9682), .A3(n9947), .A4(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17688) );
  NAND2_X1 U12811 ( .A1(n15752), .A2(n9743), .ZN(n9954) );
  NAND3_X1 U12812 ( .A1(n12594), .A2(n9954), .A3(n9958), .ZN(n9957) );
  NAND2_X1 U12814 ( .A1(n11606), .A2(n11576), .ZN(n11554) );
  NAND2_X1 U12815 ( .A1(n12922), .A2(n12921), .ZN(n9962) );
  NAND2_X1 U12816 ( .A1(n12922), .A2(n9963), .ZN(n9965) );
  INV_X1 U12817 ( .A(n12921), .ZN(n9964) );
  NAND2_X1 U12818 ( .A1(n15004), .A2(n9970), .ZN(n14985) );
  NAND2_X1 U12819 ( .A1(n16194), .A2(n9982), .ZN(n9981) );
  NAND2_X1 U12820 ( .A1(n14194), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9987) );
  NAND2_X2 U12821 ( .A1(n11600), .A2(n11622), .ZN(n12599) );
  NAND3_X1 U12822 ( .A1(n11602), .A2(n9995), .A3(n9996), .ZN(n11608) );
  NAND2_X1 U12823 ( .A1(n10141), .A2(n13906), .ZN(n9997) );
  NAND2_X1 U12824 ( .A1(n14153), .A2(n12532), .ZN(n13908) );
  OAI21_X1 U12825 ( .B1(n9664), .B2(n10003), .A(n10001), .ZN(n11659) );
  NAND3_X1 U12826 ( .A1(n10554), .A2(n10006), .A3(n10009), .ZN(n12692) );
  AND2_X2 U12827 ( .A1(n10008), .A2(n10007), .ZN(n10006) );
  NAND3_X1 U12828 ( .A1(n10011), .A2(n10366), .A3(n10367), .ZN(n10010) );
  NAND2_X1 U12829 ( .A1(n10015), .A2(n10012), .ZN(n10996) );
  NAND2_X1 U12830 ( .A1(n10014), .A2(n9697), .ZN(n10012) );
  INV_X1 U12831 ( .A(n10991), .ZN(n10014) );
  NAND3_X2 U12832 ( .A1(n10766), .A2(n10765), .A3(n10988), .ZN(n10991) );
  AND2_X2 U12833 ( .A1(n10675), .A2(n10676), .ZN(n10750) );
  AND2_X2 U12834 ( .A1(n10663), .A2(n10674), .ZN(n10749) );
  AOI21_X2 U12835 ( .B1(n15186), .B2(n15187), .A(n10305), .ZN(n15181) );
  NAND2_X1 U12836 ( .A1(n10028), .A2(n10029), .ZN(n16153) );
  INV_X1 U12837 ( .A(n12712), .ZN(n12847) );
  NAND2_X1 U12838 ( .A1(n13463), .A2(n12712), .ZN(n12698) );
  NOR2_X1 U12839 ( .A1(n10587), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12712) );
  NAND2_X1 U12840 ( .A1(n13260), .A2(n10044), .ZN(n15070) );
  INV_X1 U12841 ( .A(n16289), .ZN(n10047) );
  NAND2_X1 U12842 ( .A1(n10047), .A2(n10048), .ZN(n16254) );
  NOR3_X1 U12843 ( .A1(n15068), .A2(n14848), .A3(n13248), .ZN(n15048) );
  NAND3_X1 U12844 ( .A1(n10059), .A2(n10058), .A3(n15047), .ZN(n10057) );
  INV_X1 U12845 ( .A(n11759), .ZN(n11836) );
  OAI21_X1 U12846 ( .B1(n14578), .B2(n9791), .A(n10313), .ZN(n14581) );
  NAND4_X1 U12847 ( .A1(n10064), .A2(n11586), .A3(n9727), .A4(n9689), .ZN(
        n13417) );
  NAND2_X1 U12848 ( .A1(n10066), .A2(n13852), .ZN(n13853) );
  NAND2_X1 U12849 ( .A1(n13340), .A2(n12365), .ZN(n10066) );
  NAND2_X1 U12850 ( .A1(n14287), .A2(n9784), .ZN(n10067) );
  OR2_X1 U12851 ( .A1(n14287), .A2(n12360), .ZN(n10068) );
  NAND2_X1 U12852 ( .A1(n14287), .A2(n9775), .ZN(n14255) );
  INV_X1 U12853 ( .A(n10073), .ZN(n14460) );
  INV_X1 U12854 ( .A(n14349), .ZN(n10084) );
  NAND2_X1 U12855 ( .A1(n10086), .A2(n9741), .ZN(n10085) );
  NAND2_X1 U12856 ( .A1(n15258), .A2(n11003), .ZN(n10091) );
  AND2_X2 U12857 ( .A1(n10604), .A2(n10593), .ZN(n11028) );
  NAND3_X1 U12858 ( .A1(n10604), .A2(P2_REIP_REG_1__SCAN_IN), .A3(n10593), 
        .ZN(n10092) );
  NOR2_X1 U12859 ( .A1(n12910), .A2(n10686), .ZN(n10689) );
  CLKBUF_X1 U12860 ( .A(n12910), .Z(n10093) );
  NAND3_X1 U12861 ( .A1(n10102), .A2(n10273), .A3(n10099), .ZN(P2_U3015) );
  INV_X1 U12862 ( .A(n17575), .ZN(n11273) );
  OR3_X2 U12863 ( .A1(n17590), .A2(n17941), .A3(n17667), .ZN(n17575) );
  NAND3_X1 U12864 ( .A1(n11242), .A2(n10112), .A3(n10107), .ZN(n15800) );
  NAND3_X1 U12865 ( .A1(n11246), .A2(n11243), .A3(n10109), .ZN(n10108) );
  NAND2_X1 U12866 ( .A1(n10115), .A2(n17849), .ZN(n10114) );
  AOI21_X1 U12867 ( .B1(n17553), .B2(n11463), .A(n17920), .ZN(n10124) );
  INV_X2 U12868 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18887) );
  NAND3_X1 U12869 ( .A1(n11622), .A2(n11600), .A3(n11612), .ZN(n11555) );
  OAI21_X1 U12870 ( .B1(n15903), .B2(n9715), .A(n15897), .ZN(n10138) );
  INV_X1 U12871 ( .A(n10138), .ZN(n10137) );
  OAI21_X1 U12872 ( .B1(n13906), .B2(n10140), .A(n10139), .ZN(n15898) );
  AOI21_X1 U12873 ( .B1(n15903), .B2(n10142), .A(n9715), .ZN(n10139) );
  INV_X1 U12874 ( .A(n15903), .ZN(n10140) );
  NOR2_X1 U12875 ( .A1(n9715), .A2(n10142), .ZN(n10141) );
  NAND2_X1 U12876 ( .A1(n15904), .A2(n15903), .ZN(n15902) );
  INV_X1 U12877 ( .A(n13315), .ZN(n10144) );
  NAND4_X1 U12878 ( .A1(n10144), .A2(n13654), .A3(n11599), .A4(n10143), .ZN(
        n12341) );
  NAND2_X1 U12879 ( .A1(n10161), .A2(n10162), .ZN(n10831) );
  NAND2_X1 U12880 ( .A1(n10861), .A2(n9709), .ZN(n10916) );
  NAND2_X1 U12881 ( .A1(n10861), .A2(n10903), .ZN(n10908) );
  INV_X1 U12882 ( .A(n10169), .ZN(n10922) );
  NOR2_X2 U12883 ( .A1(n14905), .A2(n14906), .ZN(n14904) );
  AND2_X2 U12884 ( .A1(n9655), .A2(n10176), .ZN(n14905) );
  OR2_X2 U12885 ( .A1(n12619), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10178) );
  INV_X1 U12886 ( .A(n10183), .ZN(n12657) );
  AND3_X2 U12887 ( .A1(n9636), .A2(n10183), .A3(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12654) );
  NAND2_X1 U12888 ( .A1(n10186), .A2(n10187), .ZN(n13242) );
  AND2_X2 U12889 ( .A1(n10186), .A2(n10184), .ZN(n14843) );
  NAND2_X1 U12890 ( .A1(n10192), .A2(n10193), .ZN(n16088) );
  NAND3_X1 U12891 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10196) );
  NAND2_X1 U12892 ( .A1(n14909), .A2(n9706), .ZN(n13285) );
  INV_X1 U12893 ( .A(n13757), .ZN(n10200) );
  NAND2_X1 U12894 ( .A1(n10200), .A2(n9696), .ZN(n13880) );
  NAND2_X1 U12895 ( .A1(n13065), .A2(n10222), .ZN(n10221) );
  OR2_X2 U12896 ( .A1(n14977), .A2(n10219), .ZN(n10218) );
  NAND2_X1 U12897 ( .A1(n10218), .A2(n10221), .ZN(n14967) );
  NAND2_X1 U12898 ( .A1(n10228), .A2(n10227), .ZN(n10226) );
  NAND3_X1 U12899 ( .A1(n10644), .A2(n10643), .A3(n9704), .ZN(n10228) );
  INV_X1 U12900 ( .A(n13166), .ZN(n10240) );
  NAND2_X1 U12901 ( .A1(n10239), .A2(n14945), .ZN(n14941) );
  NAND2_X1 U12902 ( .A1(n10241), .A2(n10240), .ZN(n10239) );
  NAND2_X1 U12903 ( .A1(n10240), .A2(n10243), .ZN(n14951) );
  NAND2_X1 U12904 ( .A1(n13150), .A2(n13149), .ZN(n10243) );
  INV_X1 U12905 ( .A(n10245), .ZN(n14092) );
  NOR2_X1 U12906 ( .A1(n11835), .A2(n11781), .ZN(n10246) );
  AND2_X2 U12907 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13805) );
  NAND2_X1 U12908 ( .A1(n11813), .A2(n10248), .ZN(n11824) );
  OAI211_X1 U12909 ( .C1(n14148), .C2(n10251), .A(n11911), .B(n10249), .ZN(
        n14471) );
  NAND2_X1 U12910 ( .A1(n14148), .A2(n10250), .ZN(n11911) );
  NAND2_X1 U12911 ( .A1(n14557), .A2(n10259), .ZN(n14400) );
  NAND2_X1 U12912 ( .A1(n14282), .A2(n14283), .ZN(n14272) );
  NAND2_X1 U12913 ( .A1(n10996), .A2(n10899), .ZN(n10814) );
  NAND4_X1 U12914 ( .A1(n10275), .A2(n10276), .A3(n16309), .A4(n10274), .ZN(
        n10273) );
  NAND2_X1 U12915 ( .A1(n9738), .A2(n15136), .ZN(n10276) );
  NAND2_X1 U12916 ( .A1(n15136), .A2(n15134), .ZN(n15122) );
  NAND3_X1 U12917 ( .A1(n10276), .A2(n10274), .A3(n10275), .ZN(n15297) );
  INV_X1 U12918 ( .A(n10283), .ZN(n10282) );
  NOR2_X2 U12919 ( .A1(n10902), .A2(n15513), .ZN(n10285) );
  OAI21_X1 U12920 ( .B1(n15162), .B2(n10287), .A(n10935), .ZN(n10289) );
  NAND2_X1 U12921 ( .A1(n10289), .A2(n10937), .ZN(n10940) );
  CLKBUF_X1 U12922 ( .A(n10295), .Z(n10290) );
  OR2_X1 U12923 ( .A1(n13706), .A2(n13705), .ZN(n13707) );
  NOR2_X1 U12924 ( .A1(n11787), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11505) );
  INV_X1 U12925 ( .A(n12341), .ZN(n15752) );
  CLKBUF_X1 U12926 ( .A(n14977), .Z(n14980) );
  NAND2_X1 U12927 ( .A1(n14310), .A2(n14311), .ZN(n14297) );
  INV_X1 U12928 ( .A(n11846), .ZN(n12137) );
  NOR2_X1 U12929 ( .A1(n14957), .A2(n13127), .ZN(n13150) );
  AOI22_X1 U12930 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10524) );
  AOI22_X1 U12931 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9657), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10366) );
  AND2_X1 U12932 ( .A1(n19965), .A2(n12899), .ZN(n19031) );
  OR2_X1 U12933 ( .A1(n15027), .A2(n15005), .ZN(n10296) );
  AND2_X2 U12934 ( .A1(n20172), .A2(n12581), .ZN(n20152) );
  OR2_X1 U12935 ( .A1(n13650), .A2(n15741), .ZN(n20172) );
  NOR2_X1 U12936 ( .A1(n20512), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10297) );
  NAND2_X1 U12937 ( .A1(n12598), .A2(n19975), .ZN(n14528) );
  AND2_X1 U12938 ( .A1(n15123), .A2(n15135), .ZN(n10298) );
  INV_X1 U12939 ( .A(n17642), .ZN(n17614) );
  AND2_X1 U12940 ( .A1(n10620), .A2(n10619), .ZN(n10300) );
  INV_X1 U12941 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n14188) );
  OR2_X1 U12942 ( .A1(n11187), .A2(n11210), .ZN(n10301) );
  INV_X2 U12943 ( .A(n17257), .ZN(n17251) );
  INV_X1 U12944 ( .A(n14553), .ZN(n12600) );
  INV_X1 U12945 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n10595) );
  INV_X1 U12946 ( .A(n10319), .ZN(n10426) );
  AND3_X1 U12947 ( .A1(n10409), .A2(n10408), .A3(n10407), .ZN(n10303) );
  AND3_X1 U12948 ( .A1(n10324), .A2(n10323), .A3(n10322), .ZN(n10304) );
  NAND2_X1 U12949 ( .A1(n10940), .A2(n9731), .ZN(n15136) );
  INV_X1 U12950 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12312) );
  NOR3_X1 U12951 ( .A1(n13283), .A2(n10899), .A3(n15388), .ZN(n10305) );
  AND2_X1 U12952 ( .A1(n14543), .A2(DATAI_29_), .ZN(n10306) );
  INV_X1 U12953 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19922) );
  AND2_X1 U12954 ( .A1(n13125), .A2(n13147), .ZN(n10307) );
  INV_X1 U12955 ( .A(n15026), .ZN(n15040) );
  INV_X1 U12956 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20210) );
  AND3_X1 U12957 ( .A1(n10393), .A2(n10392), .A3(n10391), .ZN(n10308) );
  INV_X1 U12958 ( .A(n13850), .ZN(n11809) );
  AND2_X1 U12959 ( .A1(n10901), .A2(n15198), .ZN(n10310) );
  AND3_X1 U12960 ( .A1(n10369), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10368), .ZN(n10311) );
  INV_X1 U12961 ( .A(n12669), .ZN(n12846) );
  INV_X1 U12962 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19931) );
  AND4_X1 U12963 ( .A1(n10754), .A2(n10753), .A3(n10752), .A4(n10751), .ZN(
        n10312) );
  AND2_X4 U12964 ( .A1(n12549), .A2(n12498), .ZN(n10313) );
  AND4_X1 U12965 ( .A1(n11559), .A2(n11558), .A3(n11557), .A4(n11556), .ZN(
        n10314) );
  AND2_X2 U12966 ( .A1(n11503), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11993) );
  AND2_X1 U12967 ( .A1(n11578), .A2(n11577), .ZN(n10315) );
  NAND2_X1 U12968 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10594) );
  NAND2_X1 U12969 ( .A1(n10737), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10701) );
  AOI22_X1 U12970 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10741), .B1(
        n19446), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10691) );
  OR2_X1 U12971 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n12312), .ZN(
        n12310) );
  INV_X1 U12972 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11514) );
  OR2_X1 U12973 ( .A1(n11757), .A2(n11756), .ZN(n12550) );
  AND2_X1 U12974 ( .A1(n10757), .A2(n10756), .ZN(n10758) );
  INV_X1 U12975 ( .A(n12258), .ZN(n12231) );
  INV_X1 U12976 ( .A(n11835), .ZN(n11758) );
  OR2_X1 U12977 ( .A1(n11745), .A2(n11744), .ZN(n12542) );
  INV_X1 U12978 ( .A(n12496), .ZN(n11684) );
  XNOR2_X1 U12979 ( .A(n10510), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10418) );
  INV_X1 U12980 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10317) );
  INV_X1 U12981 ( .A(n14388), .ZN(n11992) );
  NOR2_X1 U12982 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13674) );
  OR2_X1 U12983 ( .A1(n11770), .A2(n11769), .ZN(n12560) );
  INV_X1 U12984 ( .A(n12326), .ZN(n12315) );
  OR2_X1 U12985 ( .A1(n12886), .A2(n10588), .ZN(n10589) );
  INV_X1 U12986 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10325) );
  AND2_X1 U12987 ( .A1(n13126), .A2(n10307), .ZN(n13127) );
  INV_X1 U12988 ( .A(n10559), .ZN(n12911) );
  INV_X1 U12989 ( .A(n15169), .ZN(n10926) );
  AND2_X1 U12990 ( .A1(n11135), .A2(n13617), .ZN(n11137) );
  NAND2_X1 U12991 ( .A1(n10664), .A2(n13613), .ZN(n10678) );
  AND2_X1 U12992 ( .A1(n17805), .A2(n17926), .ZN(n11271) );
  INV_X1 U12993 ( .A(n14374), .ZN(n12008) );
  NOR2_X1 U12994 ( .A1(n12129), .A2(n14328), .ZN(n12130) );
  NAND2_X1 U12995 ( .A1(n14474), .A2(n11911), .ZN(n14557) );
  NAND2_X1 U12996 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11816) );
  INV_X1 U12997 ( .A(n11656), .ZN(n12513) );
  AOI22_X1 U12998 ( .A1(n11588), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11587), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11540) );
  OR2_X1 U12999 ( .A1(n10954), .A2(n10953), .ZN(n10956) );
  AND2_X1 U13000 ( .A1(n11093), .A2(n11092), .ZN(n14971) );
  NOR2_X1 U13001 ( .A1(n10469), .A2(n10468), .ZN(n10470) );
  INV_X1 U13002 ( .A(n13862), .ZN(n12938) );
  INV_X1 U13003 ( .A(n10524), .ZN(n10529) );
  NOR2_X1 U13004 ( .A1(n18266), .A2(n17418), .ZN(n11393) );
  BUF_X1 U13005 ( .A(n11287), .Z(n17053) );
  AND2_X1 U13006 ( .A1(n17697), .A2(n18072), .ZN(n11265) );
  NOR2_X1 U13007 ( .A1(n17416), .A2(n16526), .ZN(n11398) );
  NAND2_X1 U13008 ( .A1(n12326), .A2(n13305), .ZN(n12336) );
  OR2_X1 U13009 ( .A1(n12274), .A2(n12273), .ZN(n12353) );
  INV_X1 U13010 ( .A(n12271), .ZN(n12245) );
  AND2_X1 U13011 ( .A1(n12593), .A2(n13675), .ZN(n13554) );
  NAND2_X1 U13012 ( .A1(n13547), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12271) );
  NAND2_X1 U13013 ( .A1(n12010), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12040) );
  OR2_X1 U13014 ( .A1(n11937), .A2(n15841), .ZN(n11942) );
  INV_X1 U13015 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11886) );
  NAND2_X1 U13016 ( .A1(n11723), .A2(n11722), .ZN(n20347) );
  AND2_X1 U13017 ( .A1(n13287), .A2(n13290), .ZN(n12861) );
  INV_X1 U13018 ( .A(n12663), .ZN(n12666) );
  AND2_X1 U13019 ( .A1(n11088), .A2(n11087), .ZN(n13286) );
  OR2_X1 U13020 ( .A1(n12927), .A2(n12926), .ZN(n12932) );
  INV_X1 U13021 ( .A(n12927), .ZN(n13147) );
  OR2_X1 U13022 ( .A1(n12877), .A2(n19846), .ZN(n12713) );
  NAND2_X1 U13023 ( .A1(n15292), .A2(n15291), .ZN(n15293) );
  OR2_X1 U13024 ( .A1(n10906), .A2(n15403), .ZN(n15395) );
  OR3_X1 U13025 ( .A1(n14921), .A2(n10899), .A3(n16229), .ZN(n16113) );
  INV_X1 U13026 ( .A(n15513), .ZN(n10857) );
  OR2_X1 U13027 ( .A1(n14139), .A2(n10899), .ZN(n10845) );
  OR3_X1 U13028 ( .A1(n13394), .A2(n13596), .A3(n13390), .ZN(n13593) );
  INV_X1 U13029 ( .A(n10734), .ZN(n12700) );
  XNOR2_X1 U13030 ( .A(n15579), .B(n12932), .ZN(n13469) );
  NOR2_X1 U13031 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17805), .ZN(
        n17665) );
  INV_X2 U13032 ( .A(n17135), .ZN(n17184) );
  NAND2_X1 U13033 ( .A1(n12339), .A2(n12348), .ZN(n12340) );
  INV_X1 U13034 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14383) );
  INV_X1 U13035 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14405) );
  NOR2_X1 U13036 ( .A1(n13224), .A2(n16053), .ZN(n12356) );
  NAND2_X1 U13037 ( .A1(n12462), .A2(n12461), .ZN(n20054) );
  AND2_X1 U13038 ( .A1(n12387), .A2(n12386), .ZN(n14150) );
  NOR2_X1 U13039 ( .A1(n11974), .A2(n15821), .ZN(n11975) );
  NAND2_X1 U13040 ( .A1(n11861), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11887) );
  NOR2_X1 U13041 ( .A1(n11782), .A2(n11775), .ZN(n11861) );
  AND2_X1 U13042 ( .A1(n13913), .A2(n20200), .ZN(n15980) );
  OAI21_X1 U13043 ( .B1(n20879), .B2(n13838), .A(n13837), .ZN(n14103) );
  INV_X1 U13044 ( .A(n20314), .ZN(n20326) );
  OR2_X1 U13045 ( .A1(n14089), .A2(n12521), .ZN(n20554) );
  AND2_X1 U13046 ( .A1(n11720), .A2(n20708), .ZN(n20456) );
  NAND3_X1 U13047 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n16055), .A3(n14103), 
        .ZN(n20235) );
  INV_X1 U13048 ( .A(n13108), .ZN(n13105) );
  AND2_X1 U13049 ( .A1(n12845), .A2(n12844), .ZN(n14922) );
  AND3_X1 U13050 ( .A1(n12681), .A2(n12680), .A3(n12679), .ZN(n13946) );
  OR2_X1 U13051 ( .A1(n15375), .A2(n15374), .ZN(n15348) );
  AND3_X1 U13052 ( .A1(n12826), .A2(n12825), .A3(n12824), .ZN(n15500) );
  AND2_X1 U13053 ( .A1(n10895), .A2(n15525), .ZN(n15513) );
  AND2_X1 U13054 ( .A1(n16160), .A2(n10846), .ZN(n15202) );
  AND2_X1 U13055 ( .A1(n13592), .A2(n19819), .ZN(n13618) );
  INV_X1 U13056 ( .A(n19899), .ZN(n19589) );
  OR2_X1 U13057 ( .A1(n19662), .A2(n19656), .ZN(n19706) );
  OAI21_X1 U13058 ( .B1(n11432), .B2(n11449), .A(n11431), .ZN(n11450) );
  NOR2_X1 U13059 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16668), .ZN(n16660) );
  NOR2_X1 U13060 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16693), .ZN(n16681) );
  NOR2_X1 U13061 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16745), .ZN(n16725) );
  NOR2_X1 U13062 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16778), .ZN(n16777) );
  INV_X1 U13063 ( .A(n16905), .ZN(n16898) );
  NAND2_X1 U13064 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17340), .ZN(n17304) );
  INV_X1 U13065 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16999) );
  AOI21_X1 U13066 ( .B1(n15709), .B2(n15612), .A(n18747), .ZN(n15797) );
  NAND2_X1 U13067 ( .A1(n17725), .A2(n17897), .ZN(n17642) );
  NOR2_X1 U13068 ( .A1(n18021), .A2(n17760), .ZN(n17969) );
  AND3_X1 U13069 ( .A1(n17784), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17755) );
  NOR2_X1 U13070 ( .A1(n17859), .A2(n17857), .ZN(n17822) );
  NAND2_X1 U13071 ( .A1(n18914), .A2(n15609), .ZN(n18188) );
  INV_X1 U13072 ( .A(n18074), .ZN(n18092) );
  INV_X1 U13073 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18709) );
  AOI22_X1 U13074 ( .A1(n18727), .A2(n18722), .B1(n11489), .B2(n18728), .ZN(
        n18733) );
  OAI21_X1 U13075 ( .B1(n14706), .B2(n20014), .A(n12475), .ZN(n12476) );
  INV_X1 U13076 ( .A(n14480), .ZN(n20071) );
  NOR2_X1 U13077 ( .A1(n14532), .A2(n16409), .ZN(n13214) );
  INV_X1 U13078 ( .A(n14532), .ZN(n14542) );
  INV_X1 U13079 ( .A(n20148), .ZN(n20131) );
  NAND2_X1 U13080 ( .A1(n11975), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12009) );
  AND2_X1 U13081 ( .A1(n11829), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11839) );
  INV_X1 U13082 ( .A(n20172), .ZN(n20156) );
  AND3_X1 U13083 ( .A1(n13869), .A2(P1_STATE2_REG_1__SCAN_IN), .A3(n16055), 
        .ZN(n20167) );
  INV_X1 U13084 ( .A(n14784), .ZN(n20185) );
  NOR2_X1 U13085 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20857) );
  AND2_X1 U13086 ( .A1(n20314), .A2(n20453), .ZN(n20279) );
  INV_X1 U13087 ( .A(n20296), .ZN(n20308) );
  NOR2_X2 U13088 ( .A1(n20326), .A2(n20670), .ZN(n20342) );
  NOR2_X2 U13089 ( .A1(n20326), .A2(n20553), .ZN(n20371) );
  NOR2_X2 U13090 ( .A1(n20426), .A2(n20641), .ZN(n20421) );
  NOR2_X2 U13091 ( .A1(n20426), .A2(n20670), .ZN(n20449) );
  INV_X1 U13092 ( .A(n20459), .ZN(n20480) );
  NOR2_X1 U13093 ( .A1(n20283), .A2(n14090), .ZN(n20453) );
  NOR2_X2 U13094 ( .A1(n20554), .A2(n20641), .ZN(n20541) );
  AND2_X1 U13095 ( .A1(n20283), .A2(n12509), .ZN(n20508) );
  NOR2_X2 U13096 ( .A1(n20554), .A2(n20553), .ZN(n20628) );
  INV_X1 U13097 ( .A(n20353), .ZN(n20261) );
  NOR2_X1 U13098 ( .A1(n20353), .A2(n20228), .ZN(n20738) );
  INV_X1 U13099 ( .A(n20773), .ZN(n20759) );
  INV_X1 U13100 ( .A(n19055), .ZN(n19017) );
  NOR2_X1 U13101 ( .A1(n19054), .A2(n19931), .ZN(n18996) );
  AND2_X1 U13102 ( .A1(n19965), .A2(n12667), .ZN(n19062) );
  OR2_X1 U13103 ( .A1(n12822), .A2(n12821), .ZN(n15042) );
  INV_X1 U13104 ( .A(n19121), .ZN(n19130) );
  AND2_X1 U13105 ( .A1(n13355), .A2(n13380), .ZN(n13532) );
  AND2_X1 U13106 ( .A1(n15496), .A2(n15495), .ZN(n16141) );
  AND2_X1 U13107 ( .A1(n11018), .A2(n19959), .ZN(n19174) );
  INV_X1 U13108 ( .A(n19206), .ZN(n16303) );
  NOR2_X1 U13109 ( .A1(n15548), .A2(n15549), .ZN(n16294) );
  AND2_X1 U13110 ( .A1(n13618), .A2(n16336), .ZN(n14012) );
  AND2_X1 U13111 ( .A1(n13618), .A2(n13608), .ZN(n19202) );
  OAI21_X1 U13112 ( .B1(n19230), .B2(n19229), .A(n19228), .ZN(n19265) );
  INV_X1 U13113 ( .A(n19291), .ZN(n19294) );
  INV_X1 U13114 ( .A(n19300), .ZN(n19323) );
  AND2_X1 U13115 ( .A1(n19454), .A2(n19899), .ZN(n19384) );
  AND2_X1 U13116 ( .A1(n19454), .A2(n19661), .ZN(n19440) );
  INV_X1 U13117 ( .A(n19466), .ZN(n19474) );
  INV_X1 U13118 ( .A(n19478), .ZN(n19512) );
  NOR2_X2 U13119 ( .A1(n19480), .A2(n19520), .ZN(n19544) );
  INV_X1 U13120 ( .A(n19554), .ZN(n19576) );
  INV_X1 U13121 ( .A(n19651), .ZN(n19661) );
  INV_X1 U13122 ( .A(n19766), .ZN(n19714) );
  INV_X1 U13123 ( .A(n19745), .ZN(n19747) );
  AND2_X1 U13124 ( .A1(n19242), .A2(n19261), .ZN(n19777) );
  INV_X1 U13125 ( .A(n19905), .ZN(n19756) );
  AND2_X1 U13126 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10976), .ZN(n19819) );
  XNOR2_X1 U13127 ( .A(n16530), .B(n17418), .ZN(n18914) );
  NOR3_X1 U13128 ( .A1(n17416), .A2(n16526), .A3(n16525), .ZN(n18724) );
  NOR2_X1 U13129 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16765), .ZN(n16749) );
  NOR2_X1 U13130 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16820), .ZN(n16794) );
  INV_X1 U13131 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16866) );
  INV_X1 U13132 ( .A(n16878), .ZN(n16891) );
  NOR2_X1 U13133 ( .A1(n16670), .A2(n17043), .ZN(n17044) );
  OR3_X1 U13134 ( .A1(n17231), .A2(n17235), .A3(n17232), .ZN(n17224) );
  NAND3_X1 U13135 ( .A1(n15797), .A2(n16530), .A3(n17418), .ZN(n17079) );
  AND2_X1 U13136 ( .A1(n17306), .A2(n17338), .ZN(n17326) );
  OAI211_X1 U13137 ( .C1(n17223), .C2(n16999), .A(n11175), .B(n11174), .ZN(
        n11361) );
  NOR2_X2 U13138 ( .A1(n18702), .A2(n17406), .ZN(n17410) );
  CLKBUF_X1 U13139 ( .A(n17515), .Z(n17519) );
  OAI21_X1 U13140 ( .B1(n11499), .B2(n17901), .A(n11498), .ZN(n11500) );
  INV_X1 U13141 ( .A(n18474), .ZN(n18525) );
  AND2_X1 U13142 ( .A1(n18196), .A2(n17942), .ZN(n17984) );
  INV_X1 U13143 ( .A(n18218), .ZN(n18196) );
  NOR2_X1 U13144 ( .A1(n9647), .A2(n18196), .ZN(n18186) );
  INV_X1 U13145 ( .A(n18175), .ZN(n18214) );
  INV_X1 U13146 ( .A(n18471), .ZN(n18464) );
  NAND2_X1 U13147 ( .A1(n16528), .A2(n18232), .ZN(n18474) );
  INV_X1 U13148 ( .A(n18613), .ZN(n18615) );
  INV_X1 U13149 ( .A(n18481), .ZN(n18633) );
  INV_X1 U13150 ( .A(n18621), .ZN(n18672) );
  INV_X1 U13151 ( .A(n12476), .ZN(n12477) );
  INV_X1 U13152 ( .A(n12492), .ZN(n12493) );
  INV_X1 U13153 ( .A(n20047), .ZN(n20014) );
  INV_X1 U13154 ( .A(n20041), .ZN(n14414) );
  INV_X1 U13155 ( .A(n20046), .ZN(n14040) );
  OR2_X1 U13156 ( .A1(n12615), .A2(n14547), .ZN(n14524) );
  NOR2_X1 U13157 ( .A1(n20076), .A2(n20872), .ZN(n15781) );
  INV_X1 U13158 ( .A(n20076), .ZN(n20104) );
  OR2_X1 U13159 ( .A1(n13773), .A2(n13772), .ZN(n20150) );
  NAND2_X1 U13160 ( .A1(n13338), .A2(n13337), .ZN(n16014) );
  INV_X1 U13161 ( .A(n20188), .ZN(n20208) );
  AND2_X1 U13162 ( .A1(n13568), .A2(n13567), .ZN(n20860) );
  INV_X1 U13163 ( .A(n14825), .ZN(n20254) );
  NAND2_X1 U13164 ( .A1(n20314), .A2(n20255), .ZN(n20296) );
  AOI22_X1 U13165 ( .A1(n20286), .A2(n20288), .B1(n20514), .B2(n10297), .ZN(
        n20312) );
  OR2_X1 U13166 ( .A1(n20426), .A2(n20575), .ZN(n20398) );
  AOI22_X1 U13167 ( .A1(n20404), .A2(n20401), .B1(n20581), .B2(n10297), .ZN(
        n20425) );
  OR2_X1 U13168 ( .A1(n20426), .A2(n20553), .ZN(n20459) );
  NAND2_X1 U13169 ( .A1(n20509), .A2(n20453), .ZN(n20507) );
  AOI22_X1 U13170 ( .A1(n20519), .A2(n20515), .B1(n20514), .B2(n20513), .ZN(
        n20545) );
  NAND2_X1 U13171 ( .A1(n20509), .A2(n20508), .ZN(n20574) );
  AOI22_X1 U13172 ( .A1(n20588), .A2(n20585), .B1(n20581), .B2(n20580), .ZN(
        n20633) );
  OR2_X1 U13173 ( .A1(n20716), .A2(n20575), .ZN(n20668) );
  OR2_X1 U13174 ( .A1(n20716), .A2(n20670), .ZN(n20762) );
  AND2_X1 U13175 ( .A1(n15750), .A2(n15749), .ZN(n15763) );
  INV_X1 U13176 ( .A(n20854), .ZN(n20850) );
  INV_X1 U13177 ( .A(n20840), .ZN(n20883) );
  INV_X1 U13178 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19827) );
  AND2_X1 U13179 ( .A1(n12901), .A2(n12900), .ZN(n12902) );
  INV_X1 U13180 ( .A(n19056), .ZN(n19053) );
  XNOR2_X1 U13181 ( .A(n12663), .B(n11123), .ZN(n15281) );
  AND2_X1 U13182 ( .A1(n13208), .A2(n19819), .ZN(n15036) );
  OAI21_X1 U13183 ( .B1(n13647), .B2(n13646), .A(n13645), .ZN(n19913) );
  AND2_X1 U13184 ( .A1(n13453), .A2(n19819), .ZN(n19121) );
  NAND2_X1 U13185 ( .A1(n19121), .A2(n13463), .ZN(n19135) );
  INV_X1 U13186 ( .A(n19107), .ZN(n19139) );
  INV_X1 U13187 ( .A(n19140), .ZN(n19172) );
  CLKBUF_X1 U13188 ( .A(n13499), .Z(n13625) );
  INV_X1 U13189 ( .A(n13532), .ZN(n13626) );
  INV_X1 U13190 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16150) );
  INV_X1 U13191 ( .A(n11014), .ZN(n16207) );
  NAND2_X1 U13192 ( .A1(n13352), .A2(n11016), .ZN(n16227) );
  INV_X1 U13193 ( .A(n16309), .ZN(n19209) );
  INV_X1 U13194 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19912) );
  AND2_X1 U13195 ( .A1(n13401), .A2(n13400), .ZN(n15607) );
  NAND2_X1 U13196 ( .A1(n19276), .A2(n19415), .ZN(n19291) );
  NAND2_X1 U13197 ( .A1(n19415), .A2(n19899), .ZN(n19346) );
  NAND2_X1 U13198 ( .A1(n19415), .A2(n19661), .ZN(n19403) );
  INV_X1 U13199 ( .A(n19440), .ZN(n19437) );
  NAND2_X1 U13200 ( .A1(n19415), .A2(n19756), .ZN(n19466) );
  AND2_X1 U13201 ( .A1(n19449), .A2(n19448), .ZN(n19472) );
  AOI211_X2 U13202 ( .C1(n19484), .C2(n19485), .A(n19483), .B(n19618), .ZN(
        n19517) );
  OR2_X1 U13203 ( .A1(n19652), .A2(n19520), .ZN(n19554) );
  NAND2_X1 U13204 ( .A1(n19712), .A2(n19899), .ZN(n19600) );
  NAND2_X1 U13205 ( .A1(n19712), .A2(n19661), .ZN(n19690) );
  OR2_X1 U13206 ( .A1(n19652), .A2(n19651), .ZN(n19745) );
  NOR2_X1 U13207 ( .A1(n18724), .A2(n17479), .ZN(n18921) );
  INV_X1 U13208 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18905) );
  INV_X1 U13209 ( .A(n16906), .ZN(n16894) );
  INV_X1 U13210 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17842) );
  AND2_X1 U13211 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n16976), .ZN(n16970) );
  NOR2_X1 U13212 ( .A1(n16914), .A2(n16982), .ZN(n16996) );
  AND2_X1 U13213 ( .A1(n17260), .A2(n17130), .ZN(n17242) );
  INV_X1 U13214 ( .A(n17079), .ZN(n17260) );
  NAND2_X1 U13215 ( .A1(n18702), .A2(n17376), .ZN(n17405) );
  INV_X1 U13216 ( .A(n17446), .ZN(n17475) );
  INV_X1 U13217 ( .A(n17528), .ZN(n17521) );
  INV_X1 U13218 ( .A(n17515), .ZN(n17530) );
  INV_X1 U13219 ( .A(n17644), .ZN(n17746) );
  INV_X1 U13220 ( .A(n17806), .ZN(n17780) );
  OAI21_X2 U13221 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18900), .A(n16511), 
        .ZN(n17897) );
  OR2_X1 U13222 ( .A1(n11465), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11466) );
  INV_X1 U13223 ( .A(n18134), .ZN(n18109) );
  INV_X1 U13224 ( .A(n18186), .ZN(n18203) );
  INV_X1 U13225 ( .A(n18216), .ZN(n18210) );
  INV_X1 U13226 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18717) );
  INV_X1 U13227 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18735) );
  INV_X1 U13228 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18557) );
  INV_X1 U13229 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18574) );
  INV_X1 U13230 ( .A(n18901), .ZN(n18747) );
  INV_X1 U13231 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18854) );
  INV_X1 U13232 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18771) );
  NAND2_X1 U13233 ( .A1(n12618), .A2(n12617), .ZN(P1_U2875) );
  INV_X1 U13234 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n14044) );
  AND2_X4 U13235 ( .A1(n10328), .A2(n10639), .ZN(n13046) );
  AND2_X2 U13236 ( .A1(n9650), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13029) );
  AND2_X4 U13237 ( .A1(n14180), .A2(n10639), .ZN(n10546) );
  AND2_X2 U13238 ( .A1(n13116), .A2(n10517), .ZN(n10726) );
  AOI22_X1 U13239 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10726), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10327) );
  NAND2_X1 U13240 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13049) );
  INV_X1 U13241 ( .A(n13049), .ZN(n10318) );
  NAND3_X1 U13242 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10963) );
  INV_X1 U13243 ( .A(n10963), .ZN(n10320) );
  AOI22_X1 U13244 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n13036), .ZN(n10324) );
  AND2_X2 U13246 ( .A1(n10330), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13030) );
  NAND2_X1 U13247 ( .A1(n13030), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10323) );
  NAND2_X1 U13248 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10322) );
  AOI22_X1 U13249 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10721), .B1(
        n10421), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10326) );
  NAND3_X1 U13250 ( .A1(n10327), .A2(n10304), .A3(n10326), .ZN(n10336) );
  AOI22_X1 U13251 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10720), .B1(
        n10381), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10334) );
  BUF_X1 U13252 ( .A(n13066), .Z(n10329) );
  AND2_X2 U13253 ( .A1(n10329), .A2(n10510), .ZN(n12723) );
  AOI22_X1 U13254 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10380), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10333) );
  AOI22_X1 U13255 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10332) );
  AND2_X2 U13256 ( .A1(n10330), .A2(n10510), .ZN(n10383) );
  AND2_X4 U13257 ( .A1(n14181), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10543) );
  INV_X1 U13258 ( .A(n10543), .ZN(n13048) );
  AOI22_X1 U13259 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10383), .B1(
        n13039), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10331) );
  NAND4_X1 U13260 ( .A1(n10334), .A2(n10333), .A3(n10332), .A4(n10331), .ZN(
        n10335) );
  MUX2_X1 U13261 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n19922), .S(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n10340) );
  INV_X1 U13262 ( .A(n10340), .ZN(n10339) );
  NAND2_X1 U13263 ( .A1(n19929), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10338) );
  NAND2_X1 U13264 ( .A1(n14182), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10337) );
  NAND2_X1 U13265 ( .A1(n10338), .A2(n10337), .ZN(n11127) );
  NAND2_X1 U13266 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19939), .ZN(
        n10957) );
  NAND2_X1 U13267 ( .A1(n10958), .A2(n10338), .ZN(n10402) );
  MUX2_X1 U13268 ( .A(n10340), .B(n10339), .S(n10402), .Z(n10952) );
  AOI22_X1 U13269 ( .A1(n13046), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10344) );
  AOI22_X1 U13270 ( .A1(n13066), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9651), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10343) );
  BUF_X4 U13271 ( .A(n10478), .Z(n13187) );
  AOI22_X1 U13272 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10342) );
  AOI22_X1 U13273 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9637), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10341) );
  NAND2_X1 U13274 ( .A1(n10345), .A2(n10510), .ZN(n10352) );
  AOI22_X1 U13275 ( .A1(n13046), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10349) );
  AOI22_X1 U13276 ( .A1(n13066), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9652), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10348) );
  AOI22_X1 U13277 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9657), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10347) );
  AOI22_X1 U13278 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13047), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10346) );
  NAND2_X1 U13279 ( .A1(n10350), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10351) );
  AOI22_X1 U13280 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10356) );
  AOI22_X1 U13281 ( .A1(n13066), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9651), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10355) );
  AOI22_X1 U13282 ( .A1(n13046), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10354) );
  AOI22_X1 U13283 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9637), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10353) );
  NAND4_X1 U13284 ( .A1(n10356), .A2(n10355), .A3(n10354), .A4(n10353), .ZN(
        n10362) );
  AOI22_X1 U13285 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10360) );
  AOI22_X1 U13286 ( .A1(n13066), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9653), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10359) );
  AOI22_X1 U13287 ( .A1(n13046), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10358) );
  AOI22_X1 U13288 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13047), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10357) );
  NAND4_X1 U13289 ( .A1(n10360), .A2(n10359), .A3(n10358), .A4(n10357), .ZN(
        n10361) );
  MUX2_X2 U13290 ( .A(n10362), .B(n10361), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n19220) );
  MUX2_X1 U13291 ( .A(n10734), .B(n11131), .S(n13617), .Z(n10968) );
  AOI22_X1 U13292 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9637), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10363) );
  AOI22_X1 U13293 ( .A1(n13046), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10364) );
  AOI22_X1 U13294 ( .A1(n13046), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10369) );
  AOI22_X1 U13295 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9637), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10368) );
  AOI22_X1 U13296 ( .A1(n9656), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10478), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10371) );
  AOI22_X1 U13297 ( .A1(n13066), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9653), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10370) );
  MUX2_X1 U13298 ( .A(n14044), .B(n10968), .S(n10770), .Z(n10774) );
  AOI22_X1 U13299 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10720), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10379) );
  AOI22_X1 U13300 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n12716), .ZN(n10378) );
  AOI22_X1 U13301 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n13036), .ZN(n10375) );
  NAND2_X1 U13302 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10374) );
  AND2_X1 U13303 ( .A1(n10375), .A2(n10374), .ZN(n10377) );
  NAND2_X1 U13304 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10376) );
  NAND4_X1 U13305 ( .A1(n10379), .A2(n10378), .A3(n10377), .A4(n10376), .ZN(
        n10389) );
  AOI22_X1 U13306 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10726), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10387) );
  AOI22_X1 U13307 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U13308 ( .A1(n10381), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10385) );
  AOI22_X1 U13309 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10383), .B1(
        n13030), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10384) );
  NAND4_X1 U13310 ( .A1(n10387), .A2(n10386), .A3(n10385), .A4(n10384), .ZN(
        n10388) );
  INV_X1 U13311 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n14070) );
  NOR2_X1 U13312 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n10390) );
  MUX2_X1 U13313 ( .A(n10981), .B(n10390), .S(n19251), .Z(n10773) );
  NAND2_X1 U13314 ( .A1(n10774), .A2(n10773), .ZN(n10779) );
  AOI22_X1 U13315 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10720), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10395) );
  AOI22_X1 U13316 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n13036), .ZN(n10393) );
  NAND2_X1 U13317 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10392) );
  NAND2_X1 U13318 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10391) );
  AOI22_X1 U13319 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_11__3__SCAN_IN), .B2(n12716), .ZN(n10394) );
  NAND3_X1 U13320 ( .A1(n10395), .A2(n10308), .A3(n10394), .ZN(n10401) );
  AOI22_X1 U13321 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10726), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10399) );
  AOI22_X1 U13322 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10398) );
  AOI22_X1 U13323 ( .A1(n10381), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10397) );
  AOI22_X1 U13324 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10383), .B1(
        n13030), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10396) );
  NAND4_X1 U13325 ( .A1(n10399), .A2(n10398), .A3(n10397), .A4(n10396), .ZN(
        n10400) );
  INV_X1 U13326 ( .A(n10402), .ZN(n10404) );
  NAND2_X1 U13327 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19922), .ZN(
        n10403) );
  NAND2_X1 U13328 ( .A1(n10404), .A2(n10403), .ZN(n10406) );
  NAND2_X1 U13329 ( .A1(n10639), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10405) );
  XNOR2_X1 U13330 ( .A(n10419), .B(n10418), .ZN(n10949) );
  NOR2_X2 U13331 ( .A1(n10779), .A2(n10780), .ZN(n10788) );
  INV_X1 U13332 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n14061) );
  AOI22_X1 U13333 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__4__SCAN_IN), .B2(n10421), .ZN(n10411) );
  AOI22_X1 U13334 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10410) );
  AOI22_X1 U13335 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n13036), .ZN(n10409) );
  NAND2_X1 U13336 ( .A1(n13030), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10408) );
  NAND2_X1 U13337 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10407) );
  NAND3_X1 U13338 ( .A1(n10411), .A2(n10410), .A3(n10303), .ZN(n10417) );
  AOI22_X1 U13339 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10720), .B1(
        n10381), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10415) );
  AOI22_X1 U13340 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10726), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10414) );
  AOI22_X1 U13341 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10413) );
  AOI22_X1 U13342 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10383), .B1(
        n13039), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10412) );
  NAND4_X1 U13343 ( .A1(n10415), .A2(n10414), .A3(n10413), .A4(n10412), .ZN(
        n10416) );
  NAND2_X1 U13344 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16351), .ZN(
        n10955) );
  MUX2_X1 U13345 ( .A(n10988), .B(n10951), .S(n13617), .Z(n10420) );
  MUX2_X1 U13346 ( .A(n14061), .B(n10420), .S(n10770), .Z(n10787) );
  NAND2_X1 U13347 ( .A1(n10788), .A2(n10787), .ZN(n10763) );
  AOI22_X1 U13348 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10720), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U13349 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12716), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10431) );
  INV_X1 U13350 ( .A(n10421), .ZN(n10422) );
  INV_X1 U13351 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10738) );
  NOR2_X1 U13352 ( .A1(n10422), .A2(n10738), .ZN(n10428) );
  INV_X1 U13353 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10425) );
  INV_X1 U13354 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10424) );
  OAI22_X1 U13355 ( .A1(n10426), .A2(n10425), .B1(n10424), .B2(n10423), .ZN(
        n10427) );
  NOR2_X1 U13356 ( .A1(n10428), .A2(n10427), .ZN(n10430) );
  NAND2_X1 U13357 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10429) );
  NAND4_X1 U13358 ( .A1(n10432), .A2(n10431), .A3(n10430), .A4(n10429), .ZN(
        n10438) );
  AOI22_X1 U13359 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10726), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10436) );
  AOI22_X1 U13360 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10435) );
  AOI22_X1 U13361 ( .A1(n10381), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10434) );
  AOI22_X1 U13362 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13030), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10433) );
  NAND4_X1 U13363 ( .A1(n10436), .A2(n10435), .A3(n10434), .A4(n10433), .ZN(
        n10437) );
  MUX2_X1 U13364 ( .A(n12676), .B(P2_EBX_REG_5__SCAN_IN), .S(n19251), .Z(
        n10762) );
  AOI22_X1 U13365 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10720), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10444) );
  AOI22_X1 U13366 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_11__6__SCAN_IN), .B2(n12716), .ZN(n10443) );
  AOI22_X1 U13367 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n13036), .ZN(n10440) );
  NAND2_X1 U13368 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n10439) );
  AND2_X1 U13369 ( .A1(n10440), .A2(n10439), .ZN(n10442) );
  NAND2_X1 U13370 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10441) );
  NAND4_X1 U13371 ( .A1(n10444), .A2(n10443), .A3(n10442), .A4(n10441), .ZN(
        n10450) );
  AOI22_X1 U13372 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10726), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10448) );
  AOI22_X1 U13373 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10447) );
  AOI22_X1 U13374 ( .A1(n10381), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10446) );
  AOI22_X1 U13375 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10383), .B1(
        n13030), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10445) );
  NAND4_X1 U13376 ( .A1(n10448), .A2(n10447), .A3(n10446), .A4(n10445), .ZN(
        n10449) );
  MUX2_X1 U13377 ( .A(n10810), .B(P2_EBX_REG_6__SCAN_IN), .S(n19251), .Z(
        n10813) );
  NAND2_X1 U13378 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10454) );
  NAND2_X1 U13379 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10453) );
  NAND2_X1 U13380 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10452) );
  NAND2_X1 U13381 ( .A1(n10381), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10451) );
  NAND4_X1 U13382 ( .A1(n10454), .A2(n10453), .A3(n10452), .A4(n10451), .ZN(
        n10460) );
  NAND2_X1 U13383 ( .A1(n10721), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10458) );
  NAND2_X1 U13384 ( .A1(n13030), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10457) );
  NAND2_X1 U13385 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10456) );
  NAND2_X1 U13386 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10455) );
  NAND4_X1 U13387 ( .A1(n10458), .A2(n10457), .A3(n10456), .A4(n10455), .ZN(
        n10459) );
  NOR2_X1 U13388 ( .A1(n10460), .A2(n10459), .ZN(n10471) );
  NAND2_X1 U13389 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10464) );
  NAND2_X1 U13390 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10463) );
  NAND2_X1 U13391 ( .A1(n10720), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10462) );
  NAND2_X1 U13392 ( .A1(n10726), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10461) );
  NAND4_X1 U13393 ( .A1(n10464), .A2(n10463), .A3(n10462), .A4(n10461), .ZN(
        n10469) );
  AOI22_X1 U13394 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n13036), .ZN(n10467) );
  NAND2_X1 U13395 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10466) );
  NAND2_X1 U13396 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10465) );
  NAND3_X1 U13397 ( .A1(n10467), .A2(n10466), .A3(n10465), .ZN(n10468) );
  INV_X2 U13398 ( .A(n10947), .ZN(n10899) );
  MUX2_X1 U13399 ( .A(P2_EBX_REG_7__SCAN_IN), .B(n9665), .S(n10770), .Z(n10820) );
  NOR2_X1 U13400 ( .A1(n10813), .A2(n10820), .ZN(n10472) );
  INV_X1 U13401 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n14142) );
  NAND2_X1 U13402 ( .A1(n19251), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10847) );
  INV_X1 U13403 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10474) );
  NOR2_X1 U13404 ( .A1(n10770), .A2(n10474), .ZN(n10854) );
  INV_X1 U13405 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n11053) );
  NOR2_X1 U13406 ( .A1(n10770), .A2(n11053), .ZN(n10882) );
  NAND2_X1 U13407 ( .A1(n19251), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10880) );
  AND2_X1 U13408 ( .A1(n19251), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10475) );
  NAND2_X1 U13409 ( .A1(n19251), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10873) );
  AND2_X1 U13410 ( .A1(n19251), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10869) );
  AND2_X1 U13411 ( .A1(n19251), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10866) );
  OR2_X2 U13412 ( .A1(n10871), .A2(n10866), .ZN(n10868) );
  INV_X1 U13413 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n13256) );
  NAND2_X1 U13414 ( .A1(n10864), .A2(n13256), .ZN(n10904) );
  NAND2_X2 U13415 ( .A1(n10904), .A2(n10924), .ZN(n10861) );
  NAND2_X1 U13416 ( .A1(n19251), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10903) );
  AND2_X1 U13417 ( .A1(n19251), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10907) );
  INV_X1 U13418 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n11096) );
  NAND2_X1 U13419 ( .A1(n19251), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10929) );
  INV_X1 U13420 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n10476) );
  NOR2_X1 U13421 ( .A1(n10770), .A2(n10476), .ZN(n10933) );
  NAND2_X1 U13422 ( .A1(n19251), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U13423 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9657), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10479) );
  AOI22_X1 U13424 ( .A1(n13066), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9652), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10482) );
  AOI22_X1 U13425 ( .A1(n13046), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10481) );
  AOI22_X1 U13426 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13047), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10480) );
  NAND3_X1 U13427 ( .A1(n10482), .A2(n10481), .A3(n10480), .ZN(n10483) );
  AOI22_X1 U13428 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9657), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U13429 ( .A1(n13066), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9651), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13430 ( .A1(n13046), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13431 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13047), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10485) );
  NAND4_X1 U13432 ( .A1(n10488), .A2(n10487), .A3(n10486), .A4(n10485), .ZN(
        n10489) );
  XNOR2_X1 U13433 ( .A(n10559), .B(n10558), .ZN(n13387) );
  NAND2_X1 U13434 ( .A1(n13066), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10493) );
  NAND2_X1 U13435 ( .A1(n13046), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10492) );
  NAND2_X1 U13436 ( .A1(n9651), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10491) );
  NAND2_X1 U13437 ( .A1(n10546), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10490) );
  NAND4_X1 U13438 ( .A1(n10493), .A2(n10492), .A3(n10491), .A4(n10490), .ZN(
        n10499) );
  NAND2_X1 U13439 ( .A1(n9656), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10497) );
  NAND2_X1 U13440 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10496) );
  NAND2_X1 U13441 ( .A1(n9637), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10495) );
  NAND2_X1 U13442 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10494) );
  NAND4_X1 U13443 ( .A1(n10497), .A2(n10496), .A3(n10495), .A4(n10494), .ZN(
        n10498) );
  NAND2_X1 U13444 ( .A1(n10578), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10512) );
  NAND2_X1 U13445 ( .A1(n13047), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10503) );
  NAND2_X1 U13446 ( .A1(n9656), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10502) );
  NAND2_X1 U13447 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10501) );
  NAND2_X1 U13448 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10500) );
  NAND4_X1 U13449 ( .A1(n10503), .A2(n10502), .A3(n10501), .A4(n10500), .ZN(
        n10509) );
  NAND2_X1 U13450 ( .A1(n13066), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10507) );
  NAND2_X1 U13451 ( .A1(n13046), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10506) );
  NAND2_X1 U13452 ( .A1(n9645), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10505) );
  NAND2_X1 U13453 ( .A1(n10546), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10504) );
  NAND4_X1 U13454 ( .A1(n10507), .A2(n10506), .A3(n10505), .A4(n10504), .ZN(
        n10508) );
  NAND2_X1 U13455 ( .A1(n10581), .A2(n10510), .ZN(n10511) );
  NAND2_X2 U13456 ( .A1(n10512), .A2(n10511), .ZN(n10553) );
  INV_X1 U13457 ( .A(n10553), .ZN(n13379) );
  NAND2_X1 U13458 ( .A1(n12692), .A2(n13379), .ZN(n13383) );
  AOI22_X1 U13459 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9657), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10516) );
  AOI22_X1 U13460 ( .A1(n13066), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n9645), .ZN(n10515) );
  AOI22_X1 U13461 ( .A1(n13046), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10514) );
  AOI22_X1 U13462 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13047), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10513) );
  NAND4_X1 U13463 ( .A1(n10516), .A2(n10515), .A3(n10514), .A4(n10513), .ZN(
        n10576) );
  NAND2_X1 U13464 ( .A1(n10576), .A2(n10517), .ZN(n10523) );
  AOI22_X1 U13465 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10521) );
  AOI22_X1 U13466 ( .A1(n13066), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9653), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10520) );
  AOI22_X1 U13467 ( .A1(n13046), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10519) );
  AOI22_X1 U13468 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13047), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10518) );
  NAND4_X1 U13469 ( .A1(n10521), .A2(n10520), .A3(n10519), .A4(n10518), .ZN(
        n10577) );
  NAND2_X1 U13470 ( .A1(n10577), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10522) );
  NAND3_X1 U13473 ( .A1(n13392), .A2(n13383), .A3(n19262), .ZN(n13595) );
  INV_X1 U13474 ( .A(n10556), .ZN(n13465) );
  AOI22_X1 U13475 ( .A1(n13066), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9652), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10527) );
  AOI22_X1 U13476 ( .A1(n13046), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10526) );
  NAND3_X1 U13477 ( .A1(n10527), .A2(n10526), .A3(n10525), .ZN(n10528) );
  AOI22_X1 U13478 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9657), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10533) );
  AOI22_X1 U13479 ( .A1(n13066), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10532) );
  AOI22_X1 U13480 ( .A1(n13046), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10531) );
  AOI22_X1 U13481 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9637), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10530) );
  NAND4_X1 U13482 ( .A1(n10533), .A2(n10532), .A3(n10531), .A4(n10530), .ZN(
        n10534) );
  NAND2_X1 U13483 ( .A1(n10534), .A2(n10510), .ZN(n10535) );
  NAND2_X2 U13484 ( .A1(n10536), .A2(n10535), .ZN(n19242) );
  INV_X2 U13485 ( .A(n19242), .ZN(n10569) );
  MUX2_X1 U13486 ( .A(n13595), .B(n13448), .S(n10569), .Z(n10623) );
  AOI22_X1 U13487 ( .A1(n13066), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10538) );
  AOI22_X1 U13488 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13047), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10537) );
  AND3_X1 U13489 ( .A1(n10538), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10537), .ZN(n10541) );
  AOI22_X1 U13490 ( .A1(n13046), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10540) );
  AOI22_X1 U13491 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9657), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10539) );
  NAND3_X1 U13492 ( .A1(n10541), .A2(n10540), .A3(n10539), .ZN(n10551) );
  AOI22_X1 U13493 ( .A1(n13066), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10545) );
  AOI22_X1 U13494 ( .A1(n10478), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9657), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10548) );
  AOI22_X1 U13495 ( .A1(n13046), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10547) );
  NAND2_X1 U13496 ( .A1(n10556), .A2(n10558), .ZN(n12671) );
  NAND2_X1 U13497 ( .A1(n13206), .A2(n19220), .ZN(n10567) );
  NAND4_X1 U13498 ( .A1(n13586), .A2(n10569), .A3(n10554), .A4(n10553), .ZN(
        n10555) );
  NOR2_X2 U13499 ( .A1(n10555), .A2(n13455), .ZN(n10568) );
  INV_X1 U13500 ( .A(n10568), .ZN(n10565) );
  NAND2_X1 U13501 ( .A1(n19237), .A2(n10556), .ZN(n10557) );
  AOI21_X1 U13502 ( .B1(n12692), .B2(n19242), .A(n10557), .ZN(n10563) );
  NAND2_X1 U13503 ( .A1(n10561), .A2(n10560), .ZN(n10562) );
  NAND2_X1 U13504 ( .A1(n10563), .A2(n10562), .ZN(n10564) );
  NAND2_X1 U13505 ( .A1(n10565), .A2(n10564), .ZN(n13594) );
  AND2_X1 U13506 ( .A1(n12692), .A2(n10587), .ZN(n10621) );
  OAI21_X2 U13507 ( .B1(n10623), .B2(n10567), .A(n10566), .ZN(n10638) );
  NAND2_X2 U13508 ( .A1(n10593), .A2(n19220), .ZN(n12886) );
  NAND2_X2 U13509 ( .A1(n13347), .A2(n12886), .ZN(n16335) );
  INV_X1 U13510 ( .A(n16335), .ZN(n10570) );
  AND2_X1 U13511 ( .A1(n10574), .A2(n10603), .ZN(n13450) );
  NAND2_X2 U13512 ( .A1(n10570), .A2(n10585), .ZN(n13609) );
  NAND2_X1 U13513 ( .A1(n9877), .A2(n14188), .ZN(n19964) );
  NOR2_X1 U13514 ( .A1(n19964), .A2(n19929), .ZN(n10571) );
  AOI21_X1 U13515 ( .B1(n13609), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10571), 
        .ZN(n10572) );
  OAI21_X1 U13516 ( .B1(n14182), .B2(n10638), .A(n10572), .ZN(n10599) );
  INV_X1 U13517 ( .A(n10574), .ZN(n10575) );
  NAND3_X1 U13518 ( .A1(n10576), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10510), 
        .ZN(n10582) );
  NAND3_X1 U13519 ( .A1(n10577), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n10579) );
  OR2_X1 U13520 ( .A1(n10579), .A2(n10578), .ZN(n10580) );
  OAI21_X1 U13521 ( .B1(n10582), .B2(n10581), .A(n10580), .ZN(n10583) );
  AND2_X1 U13522 ( .A1(n10569), .A2(n10583), .ZN(n10584) );
  INV_X1 U13523 ( .A(n10586), .ZN(n10590) );
  NAND2_X1 U13524 ( .A1(n10587), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10588) );
  NAND2_X4 U13525 ( .A1(n10590), .A2(n10589), .ZN(n11112) );
  NAND2_X1 U13526 ( .A1(n10631), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10596) );
  NAND2_X1 U13527 ( .A1(n10596), .A2(n9732), .ZN(n10597) );
  INV_X1 U13528 ( .A(n10600), .ZN(n10598) );
  NAND2_X1 U13529 ( .A1(n10599), .A2(n10598), .ZN(n10602) );
  INV_X1 U13530 ( .A(n10599), .ZN(n10601) );
  NAND2_X1 U13531 ( .A1(n10604), .A2(n10603), .ZN(n10605) );
  NAND2_X1 U13532 ( .A1(n10638), .A2(n10605), .ZN(n10607) );
  NAND2_X1 U13533 ( .A1(n10607), .A2(n10606), .ZN(n10615) );
  INV_X1 U13534 ( .A(n12692), .ZN(n13463) );
  MUX2_X1 U13535 ( .A(n10608), .B(n13463), .S(n19242), .Z(n10612) );
  NOR2_X1 U13536 ( .A1(n13465), .A2(n10553), .ZN(n10610) );
  AND2_X1 U13537 ( .A1(n10609), .A2(n10610), .ZN(n10611) );
  NAND2_X1 U13538 ( .A1(n10612), .A2(n10611), .ZN(n14178) );
  NOR2_X1 U13539 ( .A1(n19964), .A2(n19939), .ZN(n10613) );
  AOI21_X1 U13540 ( .B1(n15585), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10613), 
        .ZN(n10614) );
  NAND2_X1 U13541 ( .A1(n10615), .A2(n10614), .ZN(n10660) );
  NAND2_X1 U13542 ( .A1(n11112), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10629) );
  INV_X1 U13543 ( .A(n13206), .ZN(n10616) );
  AND2_X1 U13544 ( .A1(n19220), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13476) );
  AOI22_X1 U13545 ( .A1(n10616), .A2(n13476), .B1(n10631), .B2(
        P2_EBX_REG_0__SCAN_IN), .ZN(n10620) );
  NAND2_X1 U13546 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10617) );
  NAND2_X1 U13547 ( .A1(n19964), .A2(n10617), .ZN(n10618) );
  AOI21_X1 U13548 ( .B1(n11028), .B2(P2_REIP_REG_0__SCAN_IN), .A(n10618), .ZN(
        n10619) );
  INV_X1 U13549 ( .A(n10621), .ZN(n10622) );
  NAND2_X1 U13550 ( .A1(n10623), .A2(n10622), .ZN(n13600) );
  INV_X1 U13551 ( .A(n10624), .ZN(n10625) );
  NAND2_X1 U13552 ( .A1(n10625), .A2(n16342), .ZN(n10626) );
  NAND2_X1 U13553 ( .A1(n13600), .A2(n10626), .ZN(n10627) );
  NAND2_X1 U13554 ( .A1(n10627), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10628) );
  NAND3_X1 U13555 ( .A1(n10629), .A2(n10300), .A3(n10628), .ZN(n10661) );
  NAND2_X2 U13556 ( .A1(n10653), .A2(n10630), .ZN(n10657) );
  INV_X1 U13557 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13491) );
  NAND2_X1 U13558 ( .A1(n11113), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10633) );
  NAND2_X1 U13559 ( .A1(n11028), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10632) );
  OAI211_X1 U13560 ( .C1(n14188), .C2(n13491), .A(n10633), .B(n10632), .ZN(
        n10634) );
  INV_X1 U13561 ( .A(n10634), .ZN(n10637) );
  NAND2_X1 U13562 ( .A1(n11112), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10636) );
  OR2_X1 U13563 ( .A1(n10638), .A2(n10639), .ZN(n10641) );
  AOI21_X1 U13564 ( .B1(n9877), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10640) );
  INV_X1 U13565 ( .A(n10659), .ZN(n10642) );
  OR2_X1 U13566 ( .A1(n10638), .A2(n10517), .ZN(n10646) );
  OR2_X1 U13567 ( .A1(n19964), .A2(n19912), .ZN(n10645) );
  AOI22_X1 U13568 ( .A1(n11105), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10647) );
  NAND2_X1 U13569 ( .A1(n10648), .A2(n10649), .ZN(n11019) );
  INV_X1 U13570 ( .A(n10648), .ZN(n10651) );
  NAND2_X1 U13571 ( .A1(n10651), .A2(n10650), .ZN(n10652) );
  INV_X1 U13572 ( .A(n10654), .ZN(n10670) );
  INV_X1 U13573 ( .A(n10662), .ZN(n10655) );
  NAND2_X1 U13574 ( .A1(n10670), .A2(n10655), .ZN(n10656) );
  AND2_X2 U13575 ( .A1(n12910), .A2(n19207), .ZN(n10663) );
  INV_X1 U13576 ( .A(n19063), .ZN(n13613) );
  INV_X1 U13577 ( .A(n10678), .ZN(n10674) );
  INV_X2 U13578 ( .A(n10664), .ZN(n10688) );
  INV_X1 U13579 ( .A(n10665), .ZN(n10666) );
  NOR2_X1 U13580 ( .A1(n10653), .A2(n10666), .ZN(n10668) );
  AND2_X1 U13581 ( .A1(n10688), .A2(n10668), .ZN(n10667) );
  INV_X1 U13582 ( .A(n10668), .ZN(n10687) );
  NOR2_X1 U13583 ( .A1(n10688), .A2(n10687), .ZN(n10669) );
  NAND2_X1 U13584 ( .A1(n10670), .A2(n19063), .ZN(n10686) );
  NOR2_X1 U13585 ( .A1(n10688), .A2(n10686), .ZN(n10671) );
  INV_X1 U13586 ( .A(n10686), .ZN(n10672) );
  AND2_X1 U13587 ( .A1(n10688), .A2(n10672), .ZN(n10673) );
  INV_X1 U13588 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10679) );
  NAND2_X1 U13589 ( .A1(n10681), .A2(n19207), .ZN(n10798) );
  NOR2_X1 U13590 ( .A1(n12910), .A2(n10678), .ZN(n10680) );
  NAND2_X1 U13591 ( .A1(n10680), .A2(n19207), .ZN(n10755) );
  INV_X1 U13592 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12913) );
  OAI22_X1 U13593 ( .A1(n10679), .A2(n10798), .B1(n10755), .B2(n12913), .ZN(
        n10685) );
  INV_X1 U13594 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10683) );
  NAND2_X1 U13595 ( .A1(n10680), .A2(n19193), .ZN(n10802) );
  NAND2_X1 U13596 ( .A1(n10681), .A2(n19193), .ZN(n10801) );
  INV_X1 U13597 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10682) );
  OAI22_X1 U13598 ( .A1(n10683), .A2(n10802), .B1(n10801), .B2(n10682), .ZN(
        n10684) );
  NOR2_X1 U13599 ( .A1(n10685), .A2(n10684), .ZN(n10693) );
  NOR2_X1 U13600 ( .A1(n12910), .A2(n10687), .ZN(n10690) );
  AOI22_X1 U13601 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10742), .B1(
        n10737), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10692) );
  NAND4_X1 U13602 ( .A1(n10694), .A2(n10693), .A3(n10692), .A4(n10691), .ZN(
        n10695) );
  INV_X2 U13603 ( .A(n12670), .ZN(n13380) );
  NAND2_X1 U13604 ( .A1(n10695), .A2(n19956), .ZN(n10698) );
  NAND2_X1 U13605 ( .A1(n10696), .A2(n13380), .ZN(n10697) );
  INV_X1 U13606 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12926) );
  INV_X1 U13607 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10699) );
  OAI22_X1 U13608 ( .A1(n12926), .A2(n10755), .B1(n10801), .B2(n10699), .ZN(
        n10704) );
  INV_X1 U13609 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10702) );
  NAND2_X1 U13610 ( .A1(n19613), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10700) );
  OAI211_X1 U13611 ( .C1(n10798), .C2(n10702), .A(n10701), .B(n10700), .ZN(
        n10703) );
  NOR2_X1 U13612 ( .A1(n10704), .A2(n10703), .ZN(n10719) );
  AOI22_X1 U13613 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10742), .B1(
        n19446), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10718) );
  INV_X1 U13614 ( .A(n19752), .ZN(n10706) );
  INV_X1 U13615 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10705) );
  OAI21_X1 U13616 ( .B1(n10706), .B2(n10705), .A(n19956), .ZN(n10707) );
  AOI21_X1 U13617 ( .B1(n10741), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A(
        n10707), .ZN(n10717) );
  AOI22_X1 U13618 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19525), .B1(
        n19584), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10710) );
  NAND2_X1 U13619 ( .A1(n19552), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10709) );
  NAND2_X1 U13620 ( .A1(n19654), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10708) );
  NAND3_X1 U13621 ( .A1(n10710), .A2(n10709), .A3(n10708), .ZN(n10715) );
  INV_X1 U13622 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10713) );
  NAND2_X1 U13623 ( .A1(n10750), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10712) );
  NAND2_X1 U13624 ( .A1(n10749), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10711) );
  OAI211_X1 U13625 ( .C1(n10802), .C2(n10713), .A(n10712), .B(n10711), .ZN(
        n10714) );
  NOR2_X1 U13626 ( .A1(n10715), .A2(n10714), .ZN(n10716) );
  NAND4_X1 U13627 ( .A1(n10719), .A2(n10718), .A3(n10717), .A4(n10716), .ZN(
        n10736) );
  AOI22_X1 U13628 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13030), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10725) );
  AOI22_X1 U13629 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10421), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10724) );
  AOI22_X1 U13630 ( .A1(n10720), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12716), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10723) );
  AOI22_X1 U13631 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10722) );
  NAND4_X1 U13632 ( .A1(n10725), .A2(n10724), .A3(n10723), .A4(n10722), .ZN(
        n10733) );
  AOI22_X1 U13633 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10726), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10731) );
  AOI22_X1 U13634 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10319), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10730) );
  AOI22_X1 U13635 ( .A1(n10381), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13039), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10729) );
  AOI22_X1 U13636 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13036), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10728) );
  NAND4_X1 U13637 ( .A1(n10731), .A2(n10730), .A3(n10729), .A4(n10728), .ZN(
        n10732) );
  NOR2_X1 U13638 ( .A1(n10733), .A2(n10732), .ZN(n12682) );
  OR2_X1 U13639 ( .A1(n12682), .A2(n19956), .ZN(n10980) );
  INV_X1 U13640 ( .A(n10980), .ZN(n13482) );
  NAND2_X1 U13641 ( .A1(n13482), .A2(n10981), .ZN(n10979) );
  NAND2_X1 U13642 ( .A1(n10979), .A2(n12700), .ZN(n10735) );
  AND2_X2 U13643 ( .A1(n10736), .A2(n10735), .ZN(n10766) );
  INV_X1 U13644 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10740) );
  INV_X1 U13645 ( .A(n19446), .ZN(n10739) );
  INV_X1 U13646 ( .A(n10737), .ZN(n19330) );
  OAI22_X1 U13647 ( .A1(n10740), .A2(n10739), .B1(n19330), .B2(n10738), .ZN(
        n10748) );
  INV_X1 U13648 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10746) );
  INV_X1 U13649 ( .A(n10741), .ZN(n10745) );
  INV_X1 U13650 ( .A(n10742), .ZN(n10744) );
  INV_X1 U13651 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10743) );
  OAI22_X1 U13652 ( .A1(n10746), .A2(n10745), .B1(n10744), .B2(n10743), .ZN(
        n10747) );
  NOR2_X1 U13653 ( .A1(n10748), .A2(n10747), .ZN(n10759) );
  AOI22_X1 U13654 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n10749), .B1(
        n10750), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10754) );
  AOI22_X1 U13655 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19613), .B1(
        n19552), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10753) );
  AOI22_X1 U13656 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19654), .B1(
        n19752), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10752) );
  AOI22_X1 U13657 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19525), .B1(
        n19584), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10751) );
  INV_X1 U13658 ( .A(n10755), .ZN(n19227) );
  INV_X1 U13659 ( .A(n10801), .ZN(n19417) );
  AOI22_X1 U13660 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19227), .B1(
        n19417), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10757) );
  INV_X1 U13661 ( .A(n10798), .ZN(n19359) );
  INV_X1 U13662 ( .A(n10802), .ZN(n19303) );
  AOI22_X1 U13663 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19359), .B1(
        n19303), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10756) );
  NAND3_X1 U13664 ( .A1(n10759), .A2(n10312), .A3(n10758), .ZN(n10761) );
  NAND2_X1 U13665 ( .A1(n12676), .A2(n13380), .ZN(n10760) );
  XNOR2_X1 U13666 ( .A(n10991), .B(n10792), .ZN(n10992) );
  NAND2_X1 U13667 ( .A1(n10992), .A2(n10899), .ZN(n10764) );
  XNOR2_X1 U13668 ( .A(n10763), .B(n10762), .ZN(n19043) );
  INV_X1 U13669 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10994) );
  INV_X1 U13670 ( .A(n10765), .ZN(n10768) );
  INV_X1 U13671 ( .A(n10766), .ZN(n10767) );
  NAND2_X1 U13672 ( .A1(n10768), .A2(n10767), .ZN(n10769) );
  NAND2_X1 U13673 ( .A1(n16218), .A2(n10899), .ZN(n16221) );
  INV_X1 U13674 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19191) );
  OAI21_X1 U13675 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19939), .A(
        n10957), .ZN(n11128) );
  MUX2_X1 U13676 ( .A(n12682), .B(n11128), .S(n13617), .Z(n10971) );
  INV_X1 U13677 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13410) );
  MUX2_X1 U13678 ( .A(n10971), .B(n13410), .S(n19251), .Z(n19060) );
  INV_X1 U13679 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13483) );
  NOR2_X1 U13680 ( .A1(n19060), .A2(n13483), .ZN(n19185) );
  NOR3_X1 U13681 ( .A1(n10770), .A2(n14070), .A3(n13410), .ZN(n10771) );
  NOR2_X1 U13682 ( .A1(n10771), .A2(n10773), .ZN(n19184) );
  NAND2_X1 U13683 ( .A1(n19185), .A2(n19184), .ZN(n10772) );
  NOR2_X1 U13684 ( .A1(n19185), .A2(n19184), .ZN(n19183) );
  AOI21_X1 U13685 ( .B1(n19191), .B2(n10772), .A(n19183), .ZN(n13496) );
  OR2_X1 U13686 ( .A1(n10774), .A2(n10773), .ZN(n10775) );
  NAND2_X1 U13687 ( .A1(n10779), .A2(n10775), .ZN(n14048) );
  XNOR2_X1 U13688 ( .A(n14048), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13494) );
  NAND2_X1 U13689 ( .A1(n13496), .A2(n13494), .ZN(n10778) );
  INV_X1 U13690 ( .A(n14048), .ZN(n10776) );
  NAND2_X1 U13691 ( .A1(n10776), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10777) );
  NAND2_X1 U13692 ( .A1(n10778), .A2(n10777), .ZN(n16222) );
  INV_X1 U13693 ( .A(n10779), .ZN(n10782) );
  INV_X1 U13694 ( .A(n10780), .ZN(n10781) );
  NOR2_X1 U13695 ( .A1(n10782), .A2(n10781), .ZN(n10783) );
  NOR2_X1 U13696 ( .A1(n10783), .A2(n10788), .ZN(n14083) );
  AOI21_X1 U13697 ( .B1(n16222), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n14083), .ZN(n10784) );
  NAND2_X1 U13698 ( .A1(n16221), .A2(n10784), .ZN(n10786) );
  OR2_X1 U13699 ( .A1(n16222), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10785) );
  NAND2_X1 U13700 ( .A1(n10786), .A2(n10785), .ZN(n14003) );
  XNOR2_X1 U13701 ( .A(n10788), .B(n10787), .ZN(n14056) );
  INV_X1 U13702 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14014) );
  XNOR2_X1 U13703 ( .A(n14056), .B(n14014), .ZN(n14002) );
  NAND2_X1 U13704 ( .A1(n15558), .A2(n15557), .ZN(n10791) );
  NAND2_X1 U13705 ( .A1(n10789), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10790) );
  NAND2_X1 U13706 ( .A1(n10791), .A2(n10790), .ZN(n15271) );
  AOI22_X1 U13707 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19552), .B1(
        n10749), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10796) );
  AOI22_X1 U13708 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19613), .B1(
        n10750), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10795) );
  AOI22_X1 U13709 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19525), .B1(
        n19752), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10794) );
  AOI22_X1 U13710 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19654), .B1(
        n19584), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10793) );
  INV_X1 U13711 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10799) );
  INV_X1 U13712 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10797) );
  OAI22_X1 U13713 ( .A1(n10799), .A2(n10798), .B1(n10755), .B2(n10797), .ZN(
        n10805) );
  INV_X1 U13714 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10803) );
  INV_X1 U13715 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10800) );
  OAI22_X1 U13716 ( .A1(n10803), .A2(n10802), .B1(n10801), .B2(n10800), .ZN(
        n10804) );
  NOR2_X1 U13717 ( .A1(n10805), .A2(n10804), .ZN(n10808) );
  AOI22_X1 U13718 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19446), .B1(
        n10737), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10807) );
  AOI22_X1 U13719 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10742), .B1(
        n10741), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10806) );
  NAND4_X1 U13720 ( .A1(n10809), .A2(n10808), .A3(n10807), .A4(n10806), .ZN(
        n10812) );
  NAND2_X1 U13721 ( .A1(n10810), .A2(n13380), .ZN(n10811) );
  INV_X1 U13722 ( .A(n10813), .ZN(n10818) );
  XNOR2_X1 U13723 ( .A(n10819), .B(n10818), .ZN(n13998) );
  NAND2_X1 U13724 ( .A1(n10814), .A2(n13998), .ZN(n10815) );
  INV_X1 U13725 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15548) );
  XNOR2_X1 U13726 ( .A(n10815), .B(n15548), .ZN(n15270) );
  NAND2_X1 U13727 ( .A1(n15271), .A2(n15270), .ZN(n10817) );
  NAND2_X1 U13728 ( .A1(n10815), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10816) );
  NAND2_X1 U13729 ( .A1(n10819), .A2(n10818), .ZN(n10822) );
  INV_X1 U13730 ( .A(n10820), .ZN(n10821) );
  XNOR2_X1 U13731 ( .A(n10822), .B(n10821), .ZN(n19032) );
  AND2_X1 U13732 ( .A1(n19032), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15261) );
  INV_X1 U13733 ( .A(n15261), .ZN(n10823) );
  NAND2_X1 U13734 ( .A1(n10825), .A2(n10824), .ZN(n10826) );
  AND2_X1 U13735 ( .A1(n10831), .A2(n10826), .ZN(n14110) );
  NAND2_X1 U13736 ( .A1(n14110), .A2(n10947), .ZN(n10828) );
  INV_X1 U13737 ( .A(n10828), .ZN(n10827) );
  AND2_X1 U13738 ( .A1(n10827), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16198) );
  INV_X1 U13739 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11007) );
  NAND2_X1 U13740 ( .A1(n10828), .A2(n11007), .ZN(n16196) );
  INV_X1 U13741 ( .A(n19032), .ZN(n10829) );
  INV_X1 U13742 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16293) );
  NAND2_X1 U13743 ( .A1(n10829), .A2(n16293), .ZN(n16195) );
  AND2_X1 U13744 ( .A1(n16196), .A2(n16195), .ZN(n10830) );
  AND2_X1 U13745 ( .A1(n19251), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10832) );
  MUX2_X1 U13746 ( .A(n10770), .B(n10832), .S(n10831), .Z(n10833) );
  NOR2_X1 U13747 ( .A1(n10833), .A2(n10834), .ZN(n19015) );
  AOI21_X1 U13748 ( .B1(n19015), .B2(n10947), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15530) );
  NOR2_X1 U13749 ( .A1(n10834), .A2(n14142), .ZN(n10835) );
  NAND2_X1 U13750 ( .A1(n19251), .A2(n10835), .ZN(n10836) );
  AND2_X1 U13751 ( .A1(n10924), .A2(n10836), .ZN(n10837) );
  NAND2_X1 U13752 ( .A1(n10838), .A2(n10837), .ZN(n14139) );
  INV_X1 U13753 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16269) );
  AND3_X1 U13754 ( .A1(n19251), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n10838), .ZN(
        n10839) );
  OR2_X1 U13755 ( .A1(n10840), .A2(n10839), .ZN(n19004) );
  INV_X1 U13756 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16166) );
  OAI21_X1 U13757 ( .B1(n19004), .B2(n10899), .A(n16166), .ZN(n16161) );
  INV_X1 U13758 ( .A(n19004), .ZN(n10842) );
  NOR2_X1 U13759 ( .A1(n10899), .A2(n16166), .ZN(n10841) );
  NAND2_X1 U13760 ( .A1(n10842), .A2(n10841), .ZN(n16160) );
  INV_X1 U13761 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10843) );
  NOR2_X1 U13762 ( .A1(n10899), .A2(n10843), .ZN(n10844) );
  NAND2_X1 U13763 ( .A1(n19015), .A2(n10844), .ZN(n16172) );
  OR2_X1 U13764 ( .A1(n16269), .A2(n10845), .ZN(n16174) );
  NAND2_X1 U13765 ( .A1(n16172), .A2(n16174), .ZN(n16158) );
  INV_X1 U13766 ( .A(n16158), .ZN(n10846) );
  INV_X1 U13767 ( .A(n10847), .ZN(n10849) );
  NAND2_X1 U13768 ( .A1(n10849), .A2(n10848), .ZN(n10850) );
  NAND2_X1 U13769 ( .A1(n10855), .A2(n10850), .ZN(n18998) );
  INV_X1 U13770 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11046) );
  OR2_X1 U13771 ( .A1(n10899), .A2(n11046), .ZN(n10851) );
  NOR2_X1 U13772 ( .A1(n18998), .A2(n10851), .ZN(n16151) );
  INV_X1 U13773 ( .A(n16151), .ZN(n10852) );
  OR2_X1 U13774 ( .A1(n18998), .A2(n10899), .ZN(n10853) );
  NAND2_X1 U13775 ( .A1(n10853), .A2(n11046), .ZN(n15200) );
  NAND2_X1 U13776 ( .A1(n10855), .A2(n10854), .ZN(n10856) );
  AND2_X1 U13777 ( .A1(n10884), .A2(n10856), .ZN(n18981) );
  NAND2_X1 U13778 ( .A1(n18981), .A2(n10947), .ZN(n10895) );
  INV_X1 U13779 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15525) );
  NAND2_X1 U13780 ( .A1(n19251), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10859) );
  NOR2_X1 U13781 ( .A1(n10864), .A2(n10859), .ZN(n10860) );
  OR2_X1 U13782 ( .A1(n10861), .A2(n10860), .ZN(n13257) );
  OR2_X1 U13783 ( .A1(n13257), .A2(n10899), .ZN(n10862) );
  INV_X1 U13784 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15415) );
  NAND2_X1 U13785 ( .A1(n10862), .A2(n15415), .ZN(n15199) );
  NAND3_X1 U13786 ( .A1(n10868), .A2(P2_EBX_REG_20__SCAN_IN), .A3(n19251), 
        .ZN(n10863) );
  NAND2_X1 U13787 ( .A1(n10863), .A2(n10924), .ZN(n10865) );
  OR2_X1 U13788 ( .A1(n10865), .A2(n10864), .ZN(n14889) );
  INV_X1 U13789 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15232) );
  OAI21_X1 U13790 ( .B1(n14889), .B2(n10899), .A(n15232), .ZN(n15224) );
  NAND2_X1 U13791 ( .A1(n10871), .A2(n10866), .ZN(n10867) );
  NAND2_X1 U13792 ( .A1(n10868), .A2(n10867), .ZN(n14903) );
  OR2_X1 U13793 ( .A1(n14903), .A2(n10899), .ZN(n10889) );
  INV_X1 U13794 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15442) );
  NAND2_X1 U13795 ( .A1(n10889), .A2(n15442), .ZN(n15236) );
  NAND2_X1 U13796 ( .A1(n10875), .A2(n10869), .ZN(n10870) );
  NAND2_X1 U13797 ( .A1(n10871), .A2(n10870), .ZN(n14921) );
  OR2_X1 U13798 ( .A1(n14921), .A2(n10899), .ZN(n10872) );
  INV_X1 U13799 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16229) );
  NAND2_X1 U13800 ( .A1(n10872), .A2(n16229), .ZN(n16114) );
  AND2_X1 U13801 ( .A1(n15236), .A2(n16114), .ZN(n15221) );
  AND2_X1 U13802 ( .A1(n15224), .A2(n15221), .ZN(n15212) );
  OR2_X1 U13803 ( .A1(n9739), .A2(n10873), .ZN(n10874) );
  NAND2_X1 U13804 ( .A1(n10875), .A2(n10874), .ZN(n18947) );
  OR2_X1 U13805 ( .A1(n18947), .A2(n10899), .ZN(n10876) );
  INV_X1 U13806 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10893) );
  NAND2_X1 U13807 ( .A1(n10876), .A2(n10893), .ZN(n15211) );
  NAND3_X1 U13808 ( .A1(n10878), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n19251), 
        .ZN(n10877) );
  OAI211_X1 U13809 ( .C1(n10878), .C2(P2_EBX_REG_16__SCAN_IN), .A(n10877), .B(
        n10924), .ZN(n14930) );
  OR2_X1 U13810 ( .A1(n14930), .A2(n10899), .ZN(n10879) );
  XNOR2_X1 U13811 ( .A(n10879), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15246) );
  XNOR2_X1 U13812 ( .A(n10881), .B(n10158), .ZN(n18956) );
  AOI21_X1 U13813 ( .B1(n18956), .B2(n10947), .A(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15473) );
  INV_X1 U13814 ( .A(n15473), .ZN(n10886) );
  INV_X1 U13815 ( .A(n10882), .ZN(n10883) );
  XNOR2_X1 U13816 ( .A(n10884), .B(n10883), .ZN(n18974) );
  NAND2_X1 U13817 ( .A1(n18974), .A2(n10947), .ZN(n10885) );
  INV_X1 U13818 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15494) );
  NAND2_X1 U13819 ( .A1(n10885), .A2(n15494), .ZN(n15477) );
  AND4_X1 U13820 ( .A1(n15211), .A2(n15246), .A3(n10886), .A4(n15477), .ZN(
        n10887) );
  NAND3_X1 U13821 ( .A1(n15199), .A2(n15212), .A3(n10887), .ZN(n10902) );
  OR2_X1 U13822 ( .A1(n10899), .A2(n15232), .ZN(n10888) );
  NOR2_X1 U13823 ( .A1(n14889), .A2(n10888), .ZN(n15223) );
  INV_X1 U13824 ( .A(n10889), .ZN(n10890) );
  NAND2_X1 U13825 ( .A1(n10890), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15237) );
  INV_X1 U13826 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15482) );
  NOR2_X1 U13827 ( .A1(n10899), .A2(n15482), .ZN(n10891) );
  AND2_X1 U13828 ( .A1(n18956), .A2(n10891), .ZN(n15472) );
  NOR2_X1 U13829 ( .A1(n10899), .A2(n15494), .ZN(n10892) );
  AND2_X1 U13830 ( .A1(n18974), .A2(n10892), .ZN(n15475) );
  NOR2_X1 U13831 ( .A1(n15472), .A2(n15475), .ZN(n15205) );
  OR3_X1 U13832 ( .A1(n18947), .A2(n10899), .A3(n10893), .ZN(n15210) );
  INV_X1 U13833 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15463) );
  OR2_X1 U13834 ( .A1(n10899), .A2(n15463), .ZN(n10894) );
  OR2_X1 U13835 ( .A1(n14930), .A2(n10894), .ZN(n15207) );
  INV_X1 U13836 ( .A(n10895), .ZN(n10896) );
  NAND2_X1 U13837 ( .A1(n10896), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15511) );
  AND3_X1 U13838 ( .A1(n15210), .A2(n15207), .A3(n15511), .ZN(n10897) );
  NAND4_X1 U13839 ( .A1(n15237), .A2(n15205), .A3(n10897), .A4(n16113), .ZN(
        n10898) );
  NOR2_X1 U13840 ( .A1(n15223), .A2(n10898), .ZN(n10901) );
  OR2_X1 U13841 ( .A1(n10899), .A2(n15415), .ZN(n10900) );
  OR2_X1 U13842 ( .A1(n13257), .A2(n10900), .ZN(n15198) );
  NAND2_X1 U13843 ( .A1(n10904), .A2(n10168), .ZN(n10905) );
  NAND2_X1 U13844 ( .A1(n10908), .A2(n10905), .ZN(n13272) );
  NAND2_X1 U13845 ( .A1(n10906), .A2(n15403), .ZN(n15394) );
  NAND2_X1 U13846 ( .A1(n10908), .A2(n10907), .ZN(n10909) );
  NAND2_X1 U13847 ( .A1(n10911), .A2(n10909), .ZN(n13283) );
  OR2_X1 U13848 ( .A1(n13283), .A2(n10899), .ZN(n10910) );
  XNOR2_X1 U13849 ( .A(n10910), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15187) );
  INV_X1 U13850 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15388) );
  INV_X1 U13851 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15374) );
  NAND2_X1 U13852 ( .A1(n19251), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10912) );
  MUX2_X1 U13853 ( .A(P2_EBX_REG_24__SCAN_IN), .B(n10912), .S(n10911), .Z(
        n10913) );
  NAND2_X1 U13854 ( .A1(n10913), .A2(n10924), .ZN(n16083) );
  NOR2_X1 U13855 ( .A1(n16083), .A2(n10899), .ZN(n15179) );
  INV_X1 U13856 ( .A(n15181), .ZN(n10914) );
  AND3_X1 U13857 ( .A1(n19251), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n10916), .ZN(
        n10917) );
  NOR2_X1 U13858 ( .A1(n10918), .A2(n10917), .ZN(n10920) );
  INV_X1 U13859 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15350) );
  NOR2_X1 U13860 ( .A1(n10899), .A2(n15350), .ZN(n10919) );
  NAND2_X1 U13861 ( .A1(n10920), .A2(n10919), .ZN(n10939) );
  INV_X1 U13862 ( .A(n10920), .ZN(n16078) );
  OAI21_X1 U13863 ( .B1(n16078), .B2(n10899), .A(n15350), .ZN(n10921) );
  NAND2_X1 U13864 ( .A1(n10939), .A2(n10921), .ZN(n15163) );
  INV_X1 U13865 ( .A(n15163), .ZN(n10927) );
  NOR2_X1 U13866 ( .A1(n10922), .A2(n11096), .ZN(n10923) );
  NAND2_X1 U13867 ( .A1(n19251), .A2(n10923), .ZN(n10925) );
  OAI211_X1 U13868 ( .C1(n10169), .C2(P2_EBX_REG_25__SCAN_IN), .A(n10925), .B(
        n10924), .ZN(n14871) );
  NOR2_X1 U13869 ( .A1(n14871), .A2(n10899), .ZN(n10938) );
  NOR2_X1 U13870 ( .A1(n10938), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15169) );
  INV_X1 U13871 ( .A(n10929), .ZN(n10930) );
  NAND2_X1 U13872 ( .A1(n10930), .A2(n9716), .ZN(n10931) );
  NAND2_X1 U13873 ( .A1(n10932), .A2(n10931), .ZN(n13244) );
  AOI21_X1 U13874 ( .B1(n10933), .B2(n10932), .A(n10942), .ZN(n10934) );
  INV_X1 U13875 ( .A(n10934), .ZN(n14856) );
  OAI21_X1 U13876 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n15145), .ZN(n10935) );
  INV_X1 U13877 ( .A(n15145), .ZN(n10936) );
  INV_X1 U13878 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15327) );
  NAND2_X1 U13879 ( .A1(n10936), .A2(n15327), .ZN(n10937) );
  NAND2_X1 U13880 ( .A1(n10938), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15170) );
  XNOR2_X1 U13881 ( .A(n10942), .B(n10941), .ZN(n16064) );
  INV_X1 U13882 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15314) );
  OAI21_X1 U13883 ( .B1(n16064), .B2(n10899), .A(n15314), .ZN(n15134) );
  INV_X1 U13884 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n10943) );
  NOR2_X1 U13885 ( .A1(n10770), .A2(n10943), .ZN(n10944) );
  XNOR2_X1 U13886 ( .A(n10945), .B(n10944), .ZN(n12896) );
  INV_X1 U13887 ( .A(n12896), .ZN(n10946) );
  AOI21_X1 U13888 ( .B1(n10946), .B2(n10947), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15125) );
  INV_X1 U13889 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15280) );
  INV_X1 U13890 ( .A(n16064), .ZN(n10948) );
  NAND3_X1 U13891 ( .A1(n10948), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n10947), .ZN(n15135) );
  INV_X1 U13892 ( .A(n10949), .ZN(n10950) );
  INV_X1 U13893 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16329) );
  AND2_X1 U13894 ( .A1(n16329), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10953) );
  NAND2_X1 U13895 ( .A1(n11127), .A2(n10957), .ZN(n10967) );
  AND2_X1 U13896 ( .A1(n10958), .A2(n10967), .ZN(n11124) );
  INV_X1 U13897 ( .A(n10961), .ZN(n10959) );
  NAND2_X1 U13898 ( .A1(n11124), .A2(n10959), .ZN(n10960) );
  OAI21_X1 U13899 ( .B1(n11128), .B2(n10961), .A(n16333), .ZN(n10962) );
  INV_X1 U13900 ( .A(n10962), .ZN(n10964) );
  NAND2_X1 U13901 ( .A1(n16351), .A2(n10963), .ZN(n16341) );
  INV_X1 U13902 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n13353) );
  OAI21_X1 U13903 ( .B1(n10319), .B2(n16341), .A(n13353), .ZN(n19935) );
  MUX2_X1 U13904 ( .A(n10964), .B(n19935), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n19948) );
  NOR2_X1 U13905 ( .A1(n16343), .A2(n13380), .ZN(n10966) );
  NAND2_X1 U13906 ( .A1(n19948), .A2(n10966), .ZN(n10975) );
  INV_X1 U13907 ( .A(n10967), .ZN(n10970) );
  INV_X1 U13908 ( .A(n10968), .ZN(n10969) );
  OAI21_X1 U13909 ( .B1(n10971), .B2(n10970), .A(n10969), .ZN(n10973) );
  INV_X1 U13910 ( .A(n11135), .ZN(n10972) );
  AOI21_X1 U13911 ( .B1(n10973), .B2(n10972), .A(n11140), .ZN(n19946) );
  AND2_X1 U13912 ( .A1(n13380), .A2(n19220), .ZN(n12882) );
  INV_X1 U13913 ( .A(n12882), .ZN(n13388) );
  NOR2_X1 U13914 ( .A1(n16343), .A2(n13388), .ZN(n19944) );
  NAND2_X1 U13915 ( .A1(n19946), .A2(n19944), .ZN(n10974) );
  NAND2_X1 U13916 ( .A1(n10975), .A2(n10974), .ZN(n13584) );
  NAND2_X1 U13917 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14188), .ZN(n12883) );
  INV_X1 U13918 ( .A(n12883), .ZN(n10976) );
  AND2_X1 U13919 ( .A1(n19220), .A2(n19819), .ZN(n10977) );
  NAND2_X1 U13920 ( .A1(n13584), .A2(n10977), .ZN(n13352) );
  INV_X1 U13921 ( .A(n13352), .ZN(n10978) );
  NAND2_X1 U13922 ( .A1(n10978), .A2(n19956), .ZN(n16209) );
  XOR2_X1 U13923 ( .A(n12700), .B(n10979), .Z(n13490) );
  INV_X1 U13924 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14009) );
  NAND2_X1 U13925 ( .A1(n10980), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13480) );
  INV_X1 U13926 ( .A(n10981), .ZN(n12691) );
  XNOR2_X1 U13927 ( .A(n12682), .B(n12691), .ZN(n10982) );
  NOR2_X1 U13928 ( .A1(n13480), .A2(n10982), .ZN(n10983) );
  XNOR2_X1 U13929 ( .A(n13480), .B(n10982), .ZN(n19190) );
  NOR2_X1 U13930 ( .A1(n19191), .A2(n19190), .ZN(n19189) );
  NOR2_X1 U13931 ( .A1(n10983), .A2(n19189), .ZN(n10984) );
  XNOR2_X1 U13932 ( .A(n14009), .B(n10984), .ZN(n13489) );
  NOR2_X1 U13933 ( .A1(n13490), .A2(n13489), .ZN(n13488) );
  NOR2_X1 U13934 ( .A1(n10984), .A2(n14009), .ZN(n10985) );
  OR2_X1 U13935 ( .A1(n13488), .A2(n10985), .ZN(n10986) );
  XNOR2_X1 U13936 ( .A(n10986), .B(n10175), .ZN(n16217) );
  NAND2_X1 U13937 ( .A1(n16218), .A2(n16217), .ZN(n16216) );
  NAND2_X1 U13938 ( .A1(n10986), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10987) );
  INV_X1 U13939 ( .A(n10988), .ZN(n12678) );
  NAND2_X1 U13940 ( .A1(n10989), .A2(n12678), .ZN(n10990) );
  NAND2_X1 U13941 ( .A1(n10991), .A2(n10990), .ZN(n13999) );
  BUF_X1 U13942 ( .A(n10992), .Z(n10993) );
  INV_X1 U13943 ( .A(n10993), .ZN(n10995) );
  INV_X1 U13944 ( .A(n10996), .ZN(n10997) );
  INV_X1 U13945 ( .A(n10998), .ZN(n15569) );
  NAND2_X1 U13946 ( .A1(n10999), .A2(n10996), .ZN(n11000) );
  NAND2_X1 U13947 ( .A1(n15256), .A2(n16293), .ZN(n11003) );
  INV_X1 U13948 ( .A(n15256), .ZN(n11004) );
  NAND2_X1 U13949 ( .A1(n11004), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11005) );
  XNOR2_X1 U13950 ( .A(n11006), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16192) );
  NAND2_X1 U13951 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16119) );
  OR2_X1 U13952 ( .A1(n15482), .A2(n16119), .ZN(n16234) );
  INV_X1 U13953 ( .A(n16234), .ZN(n15196) );
  NAND2_X1 U13954 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15501) );
  NOR2_X1 U13955 ( .A1(n15494), .A2(n15501), .ZN(n15423) );
  NOR3_X1 U13956 ( .A1(n10843), .A2(n16269), .A3(n16166), .ZN(n15411) );
  AND3_X1 U13957 ( .A1(n15196), .A2(n15423), .A3(n15411), .ZN(n11010) );
  AND3_X1 U13958 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(n11010), .ZN(n11012) );
  AND2_X1 U13959 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11011) );
  NAND2_X1 U13960 ( .A1(n11012), .A2(n11011), .ZN(n15284) );
  NOR2_X1 U13961 ( .A1(n15284), .A2(n15403), .ZN(n11013) );
  INV_X1 U13962 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15365) );
  INV_X1 U13963 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15311) );
  NAND2_X1 U13964 ( .A1(n12654), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12650) );
  NAND2_X1 U13965 ( .A1(n12652), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12648) );
  INV_X1 U13966 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16191) );
  NAND2_X1 U13967 ( .A1(n12646), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12643) );
  INV_X1 U13968 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18960) );
  NAND2_X1 U13969 ( .A1(n12645), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12640) );
  INV_X1 U13970 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12642) );
  NAND2_X1 U13971 ( .A1(n12639), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12637) );
  INV_X1 U13972 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15240) );
  NAND2_X1 U13973 ( .A1(n12636), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12634) );
  INV_X1 U13974 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15215) );
  NAND2_X1 U13975 ( .A1(n12633), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12631) );
  INV_X1 U13976 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15188) );
  NAND2_X1 U13977 ( .A1(n12629), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12627) );
  INV_X1 U13978 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14863) );
  NAND2_X1 U13979 ( .A1(n12625), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12622) );
  INV_X1 U13980 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13243) );
  INV_X1 U13981 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15149) );
  INV_X1 U13982 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15128) );
  NOR2_X2 U13983 ( .A1(n12621), .A2(n15128), .ZN(n11015) );
  XNOR2_X1 U13984 ( .A(n11015), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12619) );
  NOR2_X2 U13985 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19902) );
  NOR2_X1 U13986 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19900) );
  OR2_X1 U13987 ( .A1(n19902), .A2(n19900), .ZN(n19930) );
  NAND2_X1 U13988 ( .A1(n19930), .A2(n9877), .ZN(n11016) );
  INV_X1 U13989 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19553) );
  NAND2_X1 U13990 ( .A1(n19553), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11017) );
  NAND2_X1 U13991 ( .A1(n10230), .A2(n11017), .ZN(n13485) );
  INV_X1 U13992 ( .A(n19900), .ZN(n19816) );
  NOR2_X1 U13993 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19816), .ZN(n11018) );
  INV_X2 U13994 ( .A(n19174), .ZN(n19033) );
  INV_X2 U13995 ( .A(n19033), .ZN(n19192) );
  AND2_X1 U13996 ( .A1(n19192), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n15290) );
  AOI21_X1 U13997 ( .B1(n19187), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15290), .ZN(n11145) );
  NAND2_X1 U13998 ( .A1(n11118), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11022) );
  AOI22_X1 U13999 ( .A1(n9643), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11021) );
  OAI211_X1 U14000 ( .C1(n11121), .C2(n14061), .A(n11022), .B(n11021), .ZN(
        n13754) );
  AOI22_X1 U14001 ( .A1(n9643), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11024) );
  NAND2_X1 U14002 ( .A1(n11113), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11023) );
  NAND2_X1 U14003 ( .A1(n11024), .A2(n11023), .ZN(n11025) );
  AOI21_X1 U14004 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n11118), .A(
        n11025), .ZN(n13758) );
  AOI22_X1 U14005 ( .A1(n11105), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11027) );
  NAND2_X1 U14006 ( .A1(n11113), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n11026) );
  OAI211_X1 U14007 ( .C1(n10635), .C2(n15548), .A(n11027), .B(n11026), .ZN(
        n13784) );
  AOI22_X1 U14008 ( .A1(n9643), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11030) );
  NAND2_X1 U14009 ( .A1(n11113), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n11029) );
  OAI211_X1 U14010 ( .C1(n10635), .C2(n16293), .A(n11030), .B(n11029), .ZN(
        n13765) );
  INV_X1 U14011 ( .A(n13765), .ZN(n11031) );
  INV_X1 U14012 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n14118) );
  NAND2_X1 U14013 ( .A1(n11112), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11033) );
  AOI22_X1 U14014 ( .A1(n9643), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11032) );
  OAI211_X1 U14015 ( .C1(n11121), .C2(n14118), .A(n11033), .B(n11032), .ZN(
        n13858) );
  AOI22_X1 U14016 ( .A1(n11105), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11035) );
  NAND2_X1 U14017 ( .A1(n11113), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11034) );
  OAI211_X1 U14018 ( .C1(n10635), .C2(n10843), .A(n11035), .B(n11034), .ZN(
        n11036) );
  INV_X1 U14019 ( .A(n11036), .ZN(n13881) );
  NOR2_X2 U14020 ( .A1(n13880), .A2(n13881), .ZN(n13901) );
  NAND2_X1 U14021 ( .A1(n11112), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11041) );
  NAND2_X1 U14022 ( .A1(n11113), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11039) );
  AND2_X1 U14023 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11037) );
  AOI21_X1 U14024 ( .B1(n9643), .B2(P2_REIP_REG_10__SCAN_IN), .A(n11037), .ZN(
        n11038) );
  AND2_X1 U14025 ( .A1(n11039), .A2(n11038), .ZN(n11040) );
  NAND2_X1 U14026 ( .A1(n11041), .A2(n11040), .ZN(n13902) );
  INV_X1 U14027 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n19005) );
  NAND2_X1 U14028 ( .A1(n11112), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11043) );
  AOI22_X1 U14029 ( .A1(n9643), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11042) );
  OAI211_X1 U14030 ( .C1(n11121), .C2(n19005), .A(n11043), .B(n11042), .ZN(
        n13920) );
  AOI22_X1 U14031 ( .A1(n9643), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11045) );
  NAND2_X1 U14032 ( .A1(n11113), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11044) );
  OAI211_X1 U14033 ( .C1(n10635), .C2(n11046), .A(n11045), .B(n11044), .ZN(
        n14020) );
  AOI22_X1 U14034 ( .A1(n11105), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11048) );
  NAND2_X1 U14035 ( .A1(n11113), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11047) );
  AND2_X1 U14036 ( .A1(n11048), .A2(n11047), .ZN(n11050) );
  NAND2_X1 U14037 ( .A1(n11118), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11049) );
  NAND2_X1 U14038 ( .A1(n11112), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11052) );
  AOI22_X1 U14039 ( .A1(n11105), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11051) );
  OAI211_X1 U14040 ( .C1(n11121), .C2(n11053), .A(n11052), .B(n11051), .ZN(
        n15037) );
  NAND2_X1 U14041 ( .A1(n11118), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11057) );
  AOI22_X1 U14042 ( .A1(n9643), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11055) );
  NAND2_X1 U14043 ( .A1(n11113), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11054) );
  AND2_X1 U14044 ( .A1(n11055), .A2(n11054), .ZN(n11056) );
  NAND2_X1 U14045 ( .A1(n11118), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11062) );
  NAND2_X1 U14046 ( .A1(n11113), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11060) );
  AND2_X1 U14047 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11058) );
  AOI21_X1 U14048 ( .B1(n11105), .B2(P2_REIP_REG_16__SCAN_IN), .A(n11058), 
        .ZN(n11059) );
  AND2_X1 U14049 ( .A1(n11060), .A2(n11059), .ZN(n11061) );
  NAND2_X1 U14050 ( .A1(n11062), .A2(n11061), .ZN(n14925) );
  NAND2_X1 U14051 ( .A1(n11112), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11066) );
  AOI22_X1 U14052 ( .A1(n11105), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11064) );
  NAND2_X1 U14053 ( .A1(n11113), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11063) );
  AND2_X1 U14054 ( .A1(n11064), .A2(n11063), .ZN(n11065) );
  NAND2_X1 U14055 ( .A1(n11112), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11070) );
  AOI22_X1 U14056 ( .A1(n9643), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11068) );
  NAND2_X1 U14057 ( .A1(n11113), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11067) );
  AND2_X1 U14058 ( .A1(n11068), .A2(n11067), .ZN(n11069) );
  NOR2_X2 U14059 ( .A1(n15013), .A2(n14908), .ZN(n14909) );
  INV_X1 U14060 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n11073) );
  NAND2_X1 U14061 ( .A1(n11118), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11072) );
  AOI22_X1 U14062 ( .A1(n9643), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11071) );
  OAI211_X1 U14063 ( .C1(n11121), .C2(n11073), .A(n11072), .B(n11071), .ZN(
        n14893) );
  NAND2_X1 U14064 ( .A1(n11112), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11077) );
  AOI22_X1 U14065 ( .A1(n9643), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n11075) );
  NAND2_X1 U14066 ( .A1(n11113), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11074) );
  AND2_X1 U14067 ( .A1(n11075), .A2(n11074), .ZN(n11076) );
  NAND2_X1 U14068 ( .A1(n11118), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11081) );
  AOI22_X1 U14069 ( .A1(n11105), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n11079) );
  NAND2_X1 U14070 ( .A1(n11113), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11078) );
  AND2_X1 U14071 ( .A1(n11079), .A2(n11078), .ZN(n11080) );
  INV_X1 U14072 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n11084) );
  NAND2_X1 U14073 ( .A1(n11112), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11083) );
  AOI22_X1 U14074 ( .A1(n11105), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11082) );
  OAI211_X1 U14075 ( .C1(n11121), .C2(n11084), .A(n11083), .B(n11082), .ZN(
        n13273) );
  NAND2_X1 U14076 ( .A1(n11118), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11088) );
  AOI22_X1 U14077 ( .A1(n11028), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11086) );
  NAND2_X1 U14078 ( .A1(n11113), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11085) );
  AND2_X1 U14079 ( .A1(n11086), .A2(n11085), .ZN(n11087) );
  NAND2_X1 U14080 ( .A1(n11112), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11093) );
  NAND2_X1 U14081 ( .A1(n9643), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11090) );
  NAND2_X1 U14082 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11089) );
  OAI211_X1 U14083 ( .C1(n11121), .C2(n10166), .A(n11090), .B(n11089), .ZN(
        n11091) );
  INV_X1 U14084 ( .A(n11091), .ZN(n11092) );
  NAND2_X1 U14085 ( .A1(n11118), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11095) );
  AOI22_X1 U14086 ( .A1(n11105), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11094) );
  OAI211_X1 U14087 ( .C1(n11121), .C2(n11096), .A(n11095), .B(n11094), .ZN(
        n14865) );
  NAND2_X1 U14088 ( .A1(n11112), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11100) );
  AOI22_X1 U14089 ( .A1(n9643), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11098) );
  NAND2_X1 U14090 ( .A1(n11113), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n11097) );
  AND2_X1 U14091 ( .A1(n11098), .A2(n11097), .ZN(n11099) );
  AND2_X1 U14092 ( .A1(n11100), .A2(n11099), .ZN(n14954) );
  NAND2_X1 U14093 ( .A1(n11118), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11104) );
  AOI22_X1 U14094 ( .A1(n9643), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11102) );
  NAND2_X1 U14095 ( .A1(n11113), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11101) );
  AND2_X1 U14096 ( .A1(n11102), .A2(n11101), .ZN(n11103) );
  AND2_X1 U14097 ( .A1(n11104), .A2(n11103), .ZN(n13246) );
  NAND2_X1 U14098 ( .A1(n11112), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11109) );
  AOI22_X1 U14099 ( .A1(n11028), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11107) );
  NAND2_X1 U14100 ( .A1(n11113), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11106) );
  AND2_X1 U14101 ( .A1(n11107), .A2(n11106), .ZN(n11108) );
  AND2_X1 U14102 ( .A1(n11109), .A2(n11108), .ZN(n14845) );
  INV_X1 U14103 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n16060) );
  NAND2_X1 U14104 ( .A1(n11118), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11111) );
  AOI22_X1 U14105 ( .A1(n11028), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11110) );
  OAI211_X1 U14106 ( .C1(n11121), .C2(n16060), .A(n11111), .B(n11110), .ZN(
        n14935) );
  NAND2_X1 U14107 ( .A1(n14936), .A2(n14935), .ZN(n14938) );
  NAND2_X1 U14108 ( .A1(n11112), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11117) );
  AOI22_X1 U14109 ( .A1(n11028), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11115) );
  NAND2_X1 U14110 ( .A1(n11113), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11114) );
  AND2_X1 U14111 ( .A1(n11115), .A2(n11114), .ZN(n11116) );
  AND2_X1 U14112 ( .A1(n11117), .A2(n11116), .ZN(n12664) );
  INV_X1 U14113 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n12890) );
  NAND2_X1 U14114 ( .A1(n11118), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11120) );
  AOI22_X1 U14115 ( .A1(n11028), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11119) );
  OAI211_X1 U14116 ( .C1(n11121), .C2(n12890), .A(n11120), .B(n11119), .ZN(
        n11122) );
  INV_X1 U14117 ( .A(n11122), .ZN(n11123) );
  NAND2_X1 U14118 ( .A1(n13380), .A2(n11128), .ZN(n11125) );
  AOI22_X1 U14119 ( .A1(n11125), .A2(n11124), .B1(n13380), .B2(n11131), .ZN(
        n11130) );
  OAI21_X1 U14120 ( .B1(n11128), .B2(n11127), .A(n11126), .ZN(n11129) );
  OAI21_X1 U14121 ( .B1(n11130), .B2(n19220), .A(n11129), .ZN(n11134) );
  NAND2_X1 U14122 ( .A1(n19956), .A2(n16342), .ZN(n11132) );
  MUX2_X1 U14123 ( .A(n11132), .B(n13617), .S(n11131), .Z(n11133) );
  AOI21_X1 U14124 ( .B1(n11134), .B2(n11133), .A(n11135), .ZN(n11138) );
  OAI21_X1 U14125 ( .B1(n11138), .B2(n11137), .A(n11136), .ZN(n11139) );
  MUX2_X1 U14126 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n11139), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n13578) );
  NAND2_X1 U14127 ( .A1(n11140), .A2(n13476), .ZN(n11141) );
  INV_X1 U14128 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19959) );
  NOR2_X1 U14129 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19961) );
  NOR2_X1 U14130 ( .A1(n19959), .A2(n14188), .ZN(n19936) );
  NOR2_X1 U14131 ( .A1(n19961), .A2(n19936), .ZN(n11142) );
  NAND2_X1 U14132 ( .A1(n15281), .A2(n19194), .ZN(n11144) );
  OAI211_X1 U14133 ( .C1(n12619), .C2(n19182), .A(n11145), .B(n11144), .ZN(
        n11146) );
  AOI21_X1 U14134 ( .B1(n15296), .B2(n11014), .A(n11146), .ZN(n11147) );
  OAI21_X1 U14135 ( .B1(n15297), .B2(n16209), .A(n11147), .ZN(P2_U2983) );
  INV_X1 U14136 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17918) );
  INV_X1 U14137 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18580) );
  NAND3_X1 U14138 ( .A1(n18880), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11156) );
  OR2_X2 U14139 ( .A1(n18860), .A2(n11156), .ZN(n17116) );
  NOR2_X2 U14140 ( .A1(n11151), .A2(n18690), .ZN(n11148) );
  AOI22_X1 U14141 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11148), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11165) );
  OR2_X2 U14142 ( .A1(n18860), .A2(n18686), .ZN(n11186) );
  INV_X1 U14143 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17105) );
  AOI22_X1 U14144 ( .A1(n11217), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11150) );
  INV_X2 U14145 ( .A(n17188), .ZN(n17211) );
  AOI22_X1 U14146 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17210), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11149) );
  OAI211_X1 U14147 ( .C1(n11186), .C2(n17105), .A(n11150), .B(n11149), .ZN(
        n11163) );
  AOI22_X1 U14148 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11161) );
  NOR2_X1 U14149 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11152) );
  NAND2_X1 U14150 ( .A1(n11153), .A2(n11152), .ZN(n17040) );
  AOI22_X1 U14151 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11160) );
  OR2_X2 U14152 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11156), .ZN(
        n11187) );
  AOI22_X1 U14153 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11159) );
  NOR3_X1 U14154 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18887), .ZN(n11157) );
  NAND2_X1 U14155 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11157), .ZN(
        n11287) );
  NAND2_X1 U14156 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11158) );
  NAND4_X1 U14157 ( .A1(n11161), .A2(n11160), .A3(n11159), .A4(n11158), .ZN(
        n11162) );
  AOI211_X1 U14158 ( .C1(n11202), .C2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n11163), .B(n11162), .ZN(n11164) );
  AOI22_X1 U14159 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11148), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11175) );
  INV_X1 U14160 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17236) );
  AOI22_X1 U14161 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11167) );
  INV_X2 U14162 ( .A(n9713), .ZN(n17185) );
  AOI22_X1 U14163 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11166) );
  OAI211_X1 U14164 ( .C1(n11186), .C2(n17236), .A(n11167), .B(n11166), .ZN(
        n11173) );
  AOI22_X1 U14165 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11171) );
  AOI22_X1 U14166 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17210), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11170) );
  AOI22_X1 U14167 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11169) );
  NAND2_X1 U14168 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11168) );
  NAND4_X1 U14169 ( .A1(n11171), .A2(n11170), .A3(n11169), .A4(n11168), .ZN(
        n11172) );
  AOI211_X1 U14170 ( .C1(n11202), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n11173), .B(n11172), .ZN(n11174) );
  INV_X1 U14171 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17031) );
  AOI22_X1 U14172 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17210), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11185) );
  INV_X1 U14173 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17244) );
  AOI22_X1 U14174 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11177) );
  AOI22_X1 U14175 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11176) );
  OAI211_X1 U14176 ( .C1(n11186), .C2(n17244), .A(n11177), .B(n11176), .ZN(
        n11183) );
  AOI22_X1 U14177 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17167), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11181) );
  AOI22_X1 U14178 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11180) );
  AOI22_X1 U14179 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11179) );
  NAND2_X1 U14180 ( .A1(n11202), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11178) );
  NAND4_X1 U14181 ( .A1(n11181), .A2(n11180), .A3(n11179), .A4(n11178), .ZN(
        n11182) );
  AOI211_X1 U14182 ( .C1(n17049), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n11183), .B(n11182), .ZN(n11184) );
  INV_X1 U14183 ( .A(n11364), .ZN(n17397) );
  INV_X1 U14184 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17170) );
  AOI22_X1 U14185 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11195) );
  INV_X1 U14186 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17250) );
  INV_X2 U14187 ( .A(n11187), .ZN(n17150) );
  AOI22_X1 U14188 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11188) );
  OAI21_X1 U14189 ( .B1(n11186), .B2(n17250), .A(n11188), .ZN(n11193) );
  INV_X1 U14190 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17048) );
  AOI22_X1 U14191 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11148), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11190) );
  OAI211_X1 U14192 ( .C1(n11287), .C2(n17048), .A(n11191), .B(n11190), .ZN(
        n11192) );
  AOI211_X1 U14193 ( .C1(n11202), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n11193), .B(n11192), .ZN(n11194) );
  OAI211_X1 U14194 ( .C1(n17040), .C2(n17170), .A(n11195), .B(n11194), .ZN(
        n11201) );
  INV_X1 U14195 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18560) );
  AOI22_X1 U14196 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11196) );
  OAI21_X1 U14197 ( .B1(n17015), .B2(n18560), .A(n11196), .ZN(n11197) );
  INV_X1 U14198 ( .A(n11197), .ZN(n11199) );
  INV_X2 U14199 ( .A(n17133), .ZN(n17189) );
  AOI22_X1 U14200 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17211), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n17189), .ZN(n11206) );
  AOI22_X1 U14201 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n17210), .ZN(n11205) );
  AOI22_X1 U14202 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11202), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11204) );
  NAND2_X1 U14203 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11203) );
  NAND4_X1 U14204 ( .A1(n11206), .A2(n11205), .A3(n11204), .A4(n11203), .ZN(
        n11215) );
  AOI22_X1 U14205 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n9649), .ZN(n11209) );
  AOI22_X1 U14206 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17167), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11208) );
  OAI211_X1 U14207 ( .C1(n17252), .C2(n11186), .A(n11209), .B(n11208), .ZN(
        n11214) );
  AOI22_X1 U14208 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n11217), .ZN(n11212) );
  INV_X1 U14209 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11210) );
  NAND3_X1 U14210 ( .A1(n11212), .A2(n11211), .A3(n10301), .ZN(n11213) );
  INV_X1 U14211 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n18565) );
  AOI22_X1 U14212 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17210), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11216) );
  OAI21_X1 U14213 ( .B1(n17015), .B2(n18565), .A(n11216), .ZN(n11224) );
  INV_X1 U14214 ( .A(n11217), .ZN(n16983) );
  INV_X1 U14215 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17134) );
  AOI22_X1 U14216 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11223) );
  INV_X1 U14217 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17240) );
  AOI22_X1 U14218 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11218) );
  OAI21_X1 U14219 ( .B1(n11186), .B2(n17240), .A(n11218), .ZN(n11222) );
  INV_X1 U14220 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11221) );
  AOI22_X1 U14221 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11220) );
  AOI22_X1 U14222 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11219) );
  NAND2_X1 U14223 ( .A1(n11252), .A2(n9935), .ZN(n11255) );
  AOI22_X1 U14224 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n9649), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11225) );
  OAI21_X1 U14225 ( .B1(n17015), .B2(n18574), .A(n11225), .ZN(n11234) );
  INV_X1 U14226 ( .A(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17123) );
  AOI22_X1 U14227 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11232) );
  INV_X1 U14228 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18493) );
  AOI22_X1 U14229 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11226) );
  OAI21_X1 U14230 ( .B1(n17053), .B2(n18493), .A(n11226), .ZN(n11230) );
  INV_X1 U14231 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17119) );
  AOI22_X1 U14232 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11228) );
  AOI22_X1 U14233 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17210), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11227) );
  OAI211_X1 U14234 ( .C1(n11186), .C2(n17119), .A(n11228), .B(n11227), .ZN(
        n11229) );
  AOI211_X1 U14235 ( .C1(n11202), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n11230), .B(n11229), .ZN(n11231) );
  OAI211_X1 U14236 ( .C1(n9746), .C2(n17123), .A(n11232), .B(n11231), .ZN(
        n11233) );
  INV_X1 U14237 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18008) );
  NAND2_X1 U14238 ( .A1(n17665), .A2(n18008), .ZN(n11235) );
  NOR2_X1 U14239 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n11235), .ZN(
        n17628) );
  INV_X1 U14240 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17630) );
  NAND2_X1 U14241 ( .A1(n17628), .A2(n17630), .ZN(n17610) );
  NOR3_X1 U14242 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17610), .ZN(n11269) );
  NOR4_X1 U14243 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11263) );
  OAI21_X1 U14244 ( .B1(n17381), .B2(n11463), .A(n17737), .ZN(n11259) );
  INV_X1 U14245 ( .A(n11259), .ZN(n11258) );
  NAND2_X1 U14246 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n11256), .ZN(
        n11257) );
  INV_X1 U14247 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17837) );
  INV_X1 U14248 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18194) );
  OR2_X1 U14249 ( .A1(n18194), .A2(n11239), .ZN(n11248) );
  XNOR2_X1 U14250 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11239), .ZN(
        n17880) );
  NAND2_X1 U14251 ( .A1(n11369), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11247) );
  XNOR2_X1 U14252 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n17409), .ZN(
        n17886) );
  INV_X1 U14253 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17209) );
  AOI22_X1 U14254 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11246) );
  INV_X1 U14255 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17090) );
  AOI22_X1 U14256 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11241) );
  AOI22_X1 U14257 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17210), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11240) );
  OAI211_X1 U14258 ( .C1(n11186), .C2(n17090), .A(n11241), .B(n11240), .ZN(
        n11245) );
  AOI22_X1 U14259 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n9649), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11244) );
  AOI22_X1 U14260 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11148), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11243) );
  AOI22_X1 U14261 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11242) );
  INV_X1 U14262 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18884) );
  NOR2_X1 U14263 ( .A1(n17895), .A2(n18884), .ZN(n17894) );
  NAND2_X1 U14264 ( .A1(n17886), .A2(n17894), .ZN(n17885) );
  NAND2_X1 U14265 ( .A1(n11250), .A2(n11249), .ZN(n11251) );
  NAND2_X1 U14266 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17866), .ZN(
        n17865) );
  NAND2_X1 U14267 ( .A1(n11251), .A2(n17865), .ZN(n17850) );
  INV_X1 U14268 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18171) );
  XOR2_X1 U14269 ( .A(n9935), .B(n11252), .Z(n11253) );
  XNOR2_X1 U14270 ( .A(n18171), .B(n11253), .ZN(n17851) );
  NAND2_X1 U14271 ( .A1(n17850), .A2(n17851), .ZN(n17849) );
  NAND2_X1 U14272 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11253), .ZN(
        n11254) );
  INV_X1 U14273 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18150) );
  NAND2_X1 U14274 ( .A1(n11258), .A2(n11260), .ZN(n11261) );
  AOI21_X1 U14275 ( .B1(n11263), .B2(n11262), .A(n17805), .ZN(n11268) );
  NAND2_X1 U14276 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18096) );
  INV_X1 U14277 ( .A(n18096), .ZN(n17763) );
  NAND2_X1 U14278 ( .A1(n17763), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18082) );
  INV_X1 U14279 ( .A(n18082), .ZN(n18072) );
  INV_X1 U14280 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18084) );
  NAND2_X1 U14281 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17716) );
  INV_X1 U14282 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18056) );
  NOR3_X1 U14283 ( .A1(n18084), .A2(n17716), .A3(n18056), .ZN(n16380) );
  INV_X1 U14284 ( .A(n16380), .ZN(n11266) );
  NOR2_X2 U14285 ( .A1(n17736), .A2(n11266), .ZN(n11267) );
  NOR2_X2 U14286 ( .A1(n11268), .A2(n11267), .ZN(n17684) );
  NAND2_X1 U14287 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18012) );
  NOR2_X1 U14288 ( .A1(n17684), .A2(n18012), .ZN(n17627) );
  INV_X1 U14289 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17956) );
  INV_X1 U14290 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17671) );
  INV_X1 U14291 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17966) );
  NOR2_X1 U14292 ( .A1(n18008), .A2(n17966), .ZN(n17981) );
  NAND2_X1 U14293 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17981), .ZN(
        n17905) );
  NOR2_X1 U14294 ( .A1(n17671), .A2(n17905), .ZN(n17963) );
  NAND2_X1 U14295 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17963), .ZN(
        n17598) );
  NOR2_X1 U14296 ( .A1(n17956), .A2(n17598), .ZN(n11270) );
  INV_X1 U14297 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18040) );
  INV_X1 U14298 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18016) );
  OAI221_X1 U14299 ( .B1(n11269), .B2(n17627), .C1(n11269), .C2(n11270), .A(
        n17636), .ZN(n17591) );
  INV_X1 U14300 ( .A(n17636), .ZN(n17609) );
  INV_X1 U14301 ( .A(n11270), .ZN(n17941) );
  NOR2_X1 U14302 ( .A1(n17805), .A2(n17590), .ZN(n17574) );
  INV_X1 U14303 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17926) );
  INV_X1 U14304 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17925) );
  NOR2_X1 U14305 ( .A1(n17926), .A2(n17925), .ZN(n17908) );
  AOI21_X1 U14306 ( .B1(n11273), .B2(n17908), .A(n17737), .ZN(n11274) );
  NOR2_X1 U14307 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17805), .ZN(
        n11468) );
  AND2_X2 U14308 ( .A1(n17918), .A2(n11275), .ZN(n17552) );
  AOI21_X1 U14309 ( .B1(n17805), .B2(n11276), .A(n17552), .ZN(n17537) );
  AOI22_X1 U14310 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11277) );
  OAI21_X1 U14311 ( .B1(n17040), .B2(n17252), .A(n11277), .ZN(n11286) );
  AOI22_X1 U14312 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11284) );
  INV_X1 U14313 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17065) );
  AOI22_X1 U14314 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11278) );
  OAI21_X1 U14315 ( .B1(n17191), .B2(n17065), .A(n11278), .ZN(n11282) );
  INV_X1 U14316 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17187) );
  AOI22_X1 U14317 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11280) );
  AOI22_X1 U14318 ( .A1(n11217), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11279) );
  OAI211_X1 U14319 ( .C1(n11287), .C2(n17187), .A(n11280), .B(n11279), .ZN(
        n11281) );
  AOI211_X1 U14320 ( .C1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .C2(n17158), .A(
        n11282), .B(n11281), .ZN(n11283) );
  OAI211_X1 U14321 ( .C1(n17116), .C2(n18557), .A(n11284), .B(n11283), .ZN(
        n11285) );
  AOI211_X4 U14322 ( .C1(n17212), .C2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A(
        n11286), .B(n11285), .ZN(n18906) );
  INV_X1 U14323 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17179) );
  AOI22_X1 U14324 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11297) );
  INV_X1 U14325 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17058) );
  AOI22_X1 U14326 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11289) );
  AOI22_X1 U14327 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11148), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11288) );
  OAI211_X1 U14328 ( .C1(n17053), .C2(n17058), .A(n11289), .B(n11288), .ZN(
        n11295) );
  AOI22_X1 U14329 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11293) );
  AOI22_X1 U14330 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11292) );
  AOI22_X1 U14331 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17158), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11291) );
  NAND2_X1 U14332 ( .A1(n11202), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11290) );
  NAND4_X1 U14333 ( .A1(n11293), .A2(n11292), .A3(n11291), .A4(n11290), .ZN(
        n11294) );
  NOR2_X1 U14334 ( .A1(n18906), .A2(n11454), .ZN(n11440) );
  AOI22_X1 U14335 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11307) );
  INV_X1 U14336 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17115) );
  AOI22_X1 U14337 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11299) );
  AOI22_X1 U14338 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11298) );
  OAI211_X1 U14339 ( .C1(n11186), .C2(n17115), .A(n11299), .B(n11298), .ZN(
        n11305) );
  AOI22_X1 U14340 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11303) );
  AOI22_X1 U14341 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11302) );
  AOI22_X1 U14342 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11301) );
  NAND2_X1 U14343 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11300) );
  NAND4_X1 U14344 ( .A1(n11303), .A2(n11302), .A3(n11301), .A4(n11300), .ZN(
        n11304) );
  AOI211_X1 U14345 ( .C1(n11202), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n11305), .B(n11304), .ZN(n11306) );
  OAI211_X1 U14346 ( .C1(n17116), .C2(n18574), .A(n11307), .B(n11306), .ZN(
        n11391) );
  NAND2_X1 U14347 ( .A1(n11440), .A2(n11391), .ZN(n11445) );
  INV_X1 U14348 ( .A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15655) );
  AOI22_X1 U14349 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11317) );
  AOI22_X1 U14350 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11309) );
  AOI22_X1 U14351 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11308) );
  OAI211_X1 U14352 ( .C1(n17155), .C2(n17209), .A(n11309), .B(n11308), .ZN(
        n11315) );
  AOI22_X1 U14353 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11313) );
  AOI22_X1 U14354 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11312) );
  AOI22_X1 U14355 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17158), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11311) );
  NAND2_X1 U14356 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11310) );
  NAND4_X1 U14357 ( .A1(n11313), .A2(n11312), .A3(n11311), .A4(n11310), .ZN(
        n11314) );
  AOI211_X1 U14358 ( .C1(n11202), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n11315), .B(n11314), .ZN(n11316) );
  AOI21_X1 U14359 ( .B1(n18234), .B2(n16530), .A(n11454), .ZN(n11404) );
  INV_X1 U14360 ( .A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17026) );
  AOI22_X1 U14361 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11318) );
  OAI21_X1 U14362 ( .B1(n17223), .B2(n17026), .A(n11318), .ZN(n11328) );
  INV_X1 U14363 ( .A(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11326) );
  AOI22_X1 U14364 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11325) );
  INV_X1 U14365 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17136) );
  AOI22_X1 U14366 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11319) );
  OAI21_X1 U14367 ( .B1(n11186), .B2(n17136), .A(n11319), .ZN(n11323) );
  INV_X1 U14368 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17016) );
  AOI22_X1 U14369 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11321) );
  AOI22_X1 U14370 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11320) );
  OAI211_X1 U14371 ( .C1(n17053), .C2(n17016), .A(n11321), .B(n11320), .ZN(
        n11322) );
  AOI211_X1 U14372 ( .C1(n11202), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n11323), .B(n11322), .ZN(n11324) );
  OAI211_X1 U14373 ( .C1(n9746), .C2(n11326), .A(n11325), .B(n11324), .ZN(
        n11327) );
  INV_X1 U14374 ( .A(n9677), .ZN(n15611) );
  INV_X1 U14375 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17000) );
  AOI22_X1 U14376 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11329) );
  OAI21_X1 U14377 ( .B1(n17015), .B2(n17000), .A(n11329), .ZN(n11338) );
  INV_X1 U14378 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15691) );
  AOI22_X1 U14379 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11336) );
  AOI22_X1 U14380 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11330) );
  OAI21_X1 U14381 ( .B1(n11287), .B2(n16999), .A(n11330), .ZN(n11334) );
  INV_X1 U14382 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16998) );
  AOI22_X1 U14383 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U14384 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11331) );
  OAI211_X1 U14385 ( .C1(n11186), .C2(n16998), .A(n11332), .B(n11331), .ZN(
        n11333) );
  AOI211_X1 U14386 ( .C1(n11202), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n11334), .B(n11333), .ZN(n11335) );
  OAI211_X1 U14387 ( .C1(n17133), .C2(n15691), .A(n11336), .B(n11335), .ZN(
        n11337) );
  NOR2_X1 U14388 ( .A1(n18259), .A2(n17266), .ZN(n11394) );
  INV_X1 U14389 ( .A(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11340) );
  AOI22_X1 U14390 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11339) );
  OAI21_X1 U14391 ( .B1(n16983), .B2(n11340), .A(n11339), .ZN(n11349) );
  INV_X1 U14392 ( .A(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17096) );
  AOI22_X1 U14393 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11347) );
  INV_X1 U14394 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16935) );
  AOI22_X1 U14395 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11341) );
  OAI21_X1 U14396 ( .B1(n17053), .B2(n16935), .A(n11341), .ZN(n11345) );
  INV_X1 U14397 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17097) );
  AOI22_X1 U14398 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U14399 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11342) );
  OAI211_X1 U14400 ( .C1(n11186), .C2(n17097), .A(n11343), .B(n11342), .ZN(
        n11344) );
  AOI211_X1 U14401 ( .C1(n11202), .C2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n11345), .B(n11344), .ZN(n11346) );
  OAI211_X1 U14402 ( .C1(n17015), .C2(n17096), .A(n11347), .B(n11346), .ZN(
        n11348) );
  AOI211_X4 U14403 ( .C1(n17211), .C2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n11349), .B(n11348), .ZN(n18266) );
  AOI22_X1 U14404 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11350) );
  OAI21_X1 U14405 ( .B1(n17040), .B2(n17244), .A(n11350), .ZN(n11359) );
  INV_X1 U14406 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17032) );
  AOI22_X1 U14407 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11357) );
  INV_X1 U14408 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17148) );
  OAI22_X1 U14409 ( .A1(n17191), .A2(n17031), .B1(n11186), .B2(n17148), .ZN(
        n11355) );
  AOI22_X1 U14410 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U14411 ( .A1(n11217), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11352) );
  AOI22_X1 U14412 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11351) );
  NAND3_X1 U14413 ( .A1(n11353), .A2(n11352), .A3(n11351), .ZN(n11354) );
  AOI211_X1 U14414 ( .C1(n17214), .C2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n11355), .B(n11354), .ZN(n11356) );
  OAI211_X1 U14415 ( .C1(n17015), .C2(n17032), .A(n11357), .B(n11356), .ZN(
        n11358) );
  AOI211_X1 U14416 ( .C1(n15611), .C2(n18702), .A(n11394), .B(n11392), .ZN(
        n11360) );
  NAND2_X1 U14417 ( .A1(n11404), .A2(n11360), .ZN(n11434) );
  NAND2_X1 U14418 ( .A1(n11489), .A2(n17381), .ZN(n17920) );
  NAND2_X1 U14419 ( .A1(n15800), .A2(n17409), .ZN(n11366) );
  NAND2_X1 U14420 ( .A1(n11237), .A2(n11366), .ZN(n11365) );
  NAND2_X1 U14421 ( .A1(n11365), .A2(n11364), .ZN(n11374) );
  NOR2_X1 U14422 ( .A1(n17394), .A2(n11374), .ZN(n11362) );
  NAND2_X1 U14423 ( .A1(n11362), .A2(n11361), .ZN(n11377) );
  NOR2_X1 U14424 ( .A1(n17387), .A2(n11377), .ZN(n11381) );
  NAND2_X1 U14425 ( .A1(n11381), .A2(n17381), .ZN(n11382) );
  XOR2_X1 U14426 ( .A(n11362), .B(n11361), .Z(n11363) );
  XNOR2_X1 U14427 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n11363), .ZN(
        n17841) );
  XOR2_X1 U14428 ( .A(n11365), .B(n11364), .Z(n11372) );
  AND2_X1 U14429 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n11372), .ZN(
        n11373) );
  XOR2_X1 U14430 ( .A(n11237), .B(n11366), .Z(n11367) );
  NOR2_X1 U14431 ( .A1(n11367), .A2(n18194), .ZN(n11371) );
  XNOR2_X1 U14432 ( .A(n18194), .B(n11367), .ZN(n17877) );
  NOR2_X1 U14433 ( .A1(n11369), .A2(n18884), .ZN(n11370) );
  NAND3_X1 U14434 ( .A1(n17895), .A2(n11369), .A3(n18884), .ZN(n11368) );
  OAI221_X1 U14435 ( .B1(n11370), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n17895), .C2(n11369), .A(n11368), .ZN(n17876) );
  NOR2_X1 U14436 ( .A1(n17877), .A2(n17876), .ZN(n17875) );
  NOR2_X1 U14437 ( .A1(n11371), .A2(n17875), .ZN(n17869) );
  XNOR2_X1 U14438 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n11372), .ZN(
        n17868) );
  NOR2_X1 U14439 ( .A1(n17869), .A2(n17868), .ZN(n17867) );
  NOR2_X1 U14440 ( .A1(n11373), .A2(n17867), .ZN(n11376) );
  XOR2_X1 U14441 ( .A(n11374), .B(n9935), .Z(n11375) );
  NOR2_X1 U14442 ( .A1(n11376), .A2(n11375), .ZN(n17853) );
  NAND2_X1 U14443 ( .A1(n11376), .A2(n11375), .ZN(n17852) );
  OAI21_X1 U14444 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n17853), .A(
        n17852), .ZN(n17840) );
  XNOR2_X1 U14445 ( .A(n11377), .B(n17387), .ZN(n11379) );
  NOR2_X1 U14446 ( .A1(n11378), .A2(n11379), .ZN(n11380) );
  NOR2_X1 U14447 ( .A1(n11380), .A2(n17829), .ZN(n11383) );
  INV_X1 U14448 ( .A(n17381), .ZN(n15720) );
  XOR2_X1 U14449 ( .A(n11381), .B(n15720), .Z(n11384) );
  NAND2_X1 U14450 ( .A1(n11383), .A2(n11384), .ZN(n17815) );
  NAND2_X1 U14451 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17815), .ZN(
        n11386) );
  NOR2_X1 U14452 ( .A1(n11382), .A2(n11386), .ZN(n11388) );
  INV_X1 U14453 ( .A(n11382), .ZN(n11387) );
  OR2_X1 U14454 ( .A1(n11384), .A2(n11383), .ZN(n17816) );
  OAI21_X1 U14455 ( .B1(n11387), .B2(n11386), .A(n17816), .ZN(n11385) );
  INV_X1 U14456 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18130) );
  NAND2_X1 U14457 ( .A1(n18072), .A2(n16380), .ZN(n18021) );
  NOR2_X1 U14458 ( .A1(n18012), .A2(n17671), .ZN(n17904) );
  INV_X1 U14459 ( .A(n17905), .ZN(n11389) );
  NAND2_X1 U14460 ( .A1(n17904), .A2(n11389), .ZN(n17965) );
  INV_X1 U14461 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17974) );
  OR2_X1 U14462 ( .A1(n17965), .A2(n17974), .ZN(n16381) );
  NOR2_X1 U14463 ( .A1(n17956), .A2(n16381), .ZN(n11413) );
  NAND2_X1 U14464 ( .A1(n17968), .A2(n11413), .ZN(n17945) );
  INV_X1 U14465 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17592) );
  NOR2_X1 U14466 ( .A1(n17945), .A2(n17592), .ZN(n17577) );
  INV_X1 U14467 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17534) );
  NOR2_X1 U14468 ( .A1(n17918), .A2(n17534), .ZN(n16383) );
  INV_X1 U14469 ( .A(n16383), .ZN(n11390) );
  NOR2_X1 U14470 ( .A1(n17911), .A2(n11390), .ZN(n16402) );
  NAND2_X1 U14471 ( .A1(n17266), .A2(n18241), .ZN(n11443) );
  NAND2_X1 U14472 ( .A1(n15611), .A2(n18259), .ZN(n18683) );
  NAND2_X1 U14473 ( .A1(n18245), .A2(n18241), .ZN(n18682) );
  NOR4_X4 U14474 ( .A1(n18234), .A2(n11392), .A3(n17266), .A4(n11400), .ZN(
        n17478) );
  NOR2_X1 U14475 ( .A1(n18254), .A2(n18259), .ZN(n11405) );
  NAND4_X1 U14476 ( .A1(n18245), .A2(n9677), .A3(n11393), .A4(n11405), .ZN(
        n11412) );
  NOR2_X1 U14477 ( .A1(n18241), .A2(n11412), .ZN(n11435) );
  INV_X1 U14478 ( .A(n11393), .ZN(n11408) );
  INV_X1 U14479 ( .A(n18682), .ZN(n11395) );
  NAND2_X1 U14480 ( .A1(n11395), .A2(n11394), .ZN(n15610) );
  INV_X1 U14481 ( .A(n15610), .ZN(n11396) );
  NAND3_X1 U14482 ( .A1(n11393), .A2(n18906), .A3(n11396), .ZN(n11397) );
  NOR2_X1 U14483 ( .A1(n11399), .A2(n17416), .ZN(n11410) );
  AOI211_X1 U14484 ( .C1(n17345), .C2(n18702), .A(n18234), .B(n16530), .ZN(
        n11439) );
  AOI21_X1 U14485 ( .B1(n11443), .B2(n11400), .A(n11439), .ZN(n11409) );
  INV_X1 U14486 ( .A(n11405), .ZN(n11453) );
  AOI21_X1 U14487 ( .B1(n17345), .B2(n11453), .A(n9677), .ZN(n11407) );
  OAI21_X1 U14488 ( .B1(n11405), .B2(n11402), .A(n11401), .ZN(n11403) );
  OAI21_X1 U14489 ( .B1(n11405), .B2(n11404), .A(n11403), .ZN(n11406) );
  INV_X1 U14490 ( .A(n18722), .ZN(n18091) );
  NAND2_X1 U14491 ( .A1(n11413), .A2(n17969), .ZN(n17947) );
  NOR2_X1 U14492 ( .A1(n17592), .A2(n17947), .ZN(n17578) );
  NAND2_X1 U14493 ( .A1(n17908), .A2(n17578), .ZN(n17545) );
  INV_X1 U14494 ( .A(n17545), .ZN(n17903) );
  NAND2_X1 U14495 ( .A1(n16383), .A2(n17903), .ZN(n16388) );
  INV_X1 U14496 ( .A(n11489), .ZN(n18729) );
  NOR2_X1 U14497 ( .A1(n18729), .A2(n17381), .ZN(n18074) );
  INV_X1 U14498 ( .A(n18703), .ZN(n18219) );
  NOR2_X1 U14499 ( .A1(n18723), .A2(n18219), .ZN(n18105) );
  INV_X1 U14500 ( .A(n18021), .ZN(n17685) );
  NAND3_X1 U14501 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11414) );
  INV_X1 U14502 ( .A(n11414), .ZN(n18018) );
  NAND3_X1 U14503 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n18018), .ZN(n18122) );
  INV_X1 U14504 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18142) );
  NOR3_X1 U14505 ( .A1(n18142), .A2(n18150), .A3(n18130), .ZN(n11415) );
  INV_X1 U14506 ( .A(n11415), .ZN(n18019) );
  NOR2_X1 U14507 ( .A1(n18122), .A2(n18019), .ZN(n18032) );
  NAND2_X1 U14508 ( .A1(n17685), .A2(n18032), .ZN(n18009) );
  NOR2_X1 U14509 ( .A1(n16381), .A2(n18009), .ZN(n17906) );
  NAND2_X1 U14510 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17906), .ZN(
        n11417) );
  NAND2_X1 U14511 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17927) );
  INV_X1 U14512 ( .A(n17927), .ZN(n17929) );
  NAND2_X1 U14513 ( .A1(n17908), .A2(n17929), .ZN(n17902) );
  INV_X1 U14514 ( .A(n17902), .ZN(n17558) );
  NAND2_X1 U14515 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17558), .ZN(
        n17549) );
  INV_X1 U14516 ( .A(n17598), .ZN(n11461) );
  AOI21_X1 U14517 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18165) );
  NOR2_X1 U14518 ( .A1(n18165), .A2(n11414), .ZN(n18124) );
  NAND2_X1 U14519 ( .A1(n11415), .A2(n18124), .ZN(n18034) );
  NOR3_X1 U14520 ( .A1(n18021), .A2(n18012), .A3(n18034), .ZN(n18010) );
  NAND2_X1 U14521 ( .A1(n11461), .A2(n18010), .ZN(n17950) );
  OAI21_X1 U14522 ( .B1(n17902), .B2(n17950), .A(n18723), .ZN(n17907) );
  OAI221_X1 U14523 ( .B1(n18703), .B2(n17906), .C1(n18703), .C2(n17558), .A(
        n17907), .ZN(n11416) );
  AOI221_X1 U14524 ( .B1(n11417), .B2(n9640), .C1(n17549), .C2(n9640), .A(
        n11416), .ZN(n11484) );
  NOR2_X1 U14525 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18883) );
  INV_X1 U14526 ( .A(n18883), .ZN(n18868) );
  NOR2_X1 U14527 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18868), .ZN(n18918) );
  INV_X1 U14528 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n16528) );
  NAND2_X1 U14529 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18707), .ZN(
        n11424) );
  OAI21_X1 U14530 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18707), .A(
        n11424), .ZN(n11448) );
  INV_X1 U14531 ( .A(n11448), .ZN(n11433) );
  AOI22_X1 U14532 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n18709), .B2(n18880), .ZN(
        n11447) );
  INV_X1 U14533 ( .A(n11447), .ZN(n11425) );
  INV_X1 U14534 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18718) );
  NOR2_X1 U14535 ( .A1(n11447), .A2(n11424), .ZN(n11418) );
  OAI22_X1 U14536 ( .A1(n18872), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18714), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11426) );
  NOR2_X1 U14537 ( .A1(n11420), .A2(n18860), .ZN(n11429) );
  AOI22_X1 U14538 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18735), .B1(
        n11420), .B2(n18860), .ZN(n11430) );
  OAI21_X1 U14539 ( .B1(n18717), .B2(n11429), .A(n11430), .ZN(n11421) );
  INV_X1 U14540 ( .A(n11421), .ZN(n11422) );
  NAND2_X1 U14541 ( .A1(n11425), .A2(n11424), .ZN(n11423) );
  OAI211_X1 U14542 ( .C1(n11425), .C2(n11424), .A(n11431), .B(n11423), .ZN(
        n11442) );
  XNOR2_X1 U14543 ( .A(n11427), .B(n11426), .ZN(n11432) );
  NAND2_X1 U14544 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18735), .ZN(
        n11428) );
  OAI22_X1 U14545 ( .A1(n11430), .A2(n18717), .B1(n11429), .B2(n11428), .ZN(
        n11449) );
  OAI21_X1 U14546 ( .B1(n11433), .B2(n11442), .A(n11450), .ZN(n18728) );
  INV_X1 U14547 ( .A(n18728), .ZN(n11446) );
  INV_X1 U14548 ( .A(n11434), .ZN(n11437) );
  AOI21_X1 U14549 ( .B1(n11437), .B2(n11436), .A(n11435), .ZN(n11438) );
  NOR2_X1 U14550 ( .A1(n11439), .A2(n11438), .ZN(n15710) );
  NAND2_X1 U14551 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n18907) );
  INV_X1 U14552 ( .A(n18907), .ZN(n18766) );
  NAND2_X1 U14553 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18771), .ZN(n18896) );
  NAND2_X1 U14554 ( .A1(n18830), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18840) );
  NOR2_X1 U14555 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18760) );
  INV_X1 U14556 ( .A(n18760), .ZN(n16507) );
  NAND3_X1 U14557 ( .A1(n18771), .A2(n18833), .A3(n16507), .ZN(n18904) );
  AOI211_X1 U14558 ( .C1(n18906), .C2(n11454), .A(n11440), .B(n17415), .ZN(
        n11441) );
  NOR2_X1 U14559 ( .A1(n18766), .A2(n11441), .ZN(n16508) );
  NAND3_X1 U14560 ( .A1(n16508), .A2(n11443), .A3(n18725), .ZN(n11444) );
  OAI211_X1 U14561 ( .C1(n11446), .C2(n11445), .A(n15710), .B(n11444), .ZN(
        n11456) );
  NOR2_X1 U14562 ( .A1(n11448), .A2(n11447), .ZN(n11452) );
  INV_X1 U14563 ( .A(n11449), .ZN(n11451) );
  OAI21_X1 U14564 ( .B1(n11454), .B2(n11453), .A(n9677), .ZN(n11455) );
  INV_X1 U14565 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18865) );
  NAND2_X1 U14566 ( .A1(n18865), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18752) );
  OAI211_X1 U14567 ( .C1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n18105), .A(
        n11484), .B(n18203), .ZN(n15721) );
  AOI21_X1 U14568 ( .B1(n16388), .B2(n18074), .A(n15721), .ZN(n11457) );
  OAI21_X1 U14569 ( .B1(n16402), .B2(n18091), .A(n11457), .ZN(n11458) );
  NOR2_X2 U14570 ( .A1(n18218), .A2(n17920), .ZN(n18134) );
  AOI22_X1 U14571 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n11459), .B1(
        n17552), .B2(n11464), .ZN(n11467) );
  NAND2_X1 U14572 ( .A1(n9647), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17540) );
  INV_X1 U14573 ( .A(n9640), .ZN(n18701) );
  OAI21_X1 U14574 ( .B1(n18701), .B2(n18884), .A(n18703), .ZN(n18187) );
  OAI22_X1 U14575 ( .A1(n17762), .A2(n18091), .B1(n17760), .B2(n18092), .ZN(
        n18020) );
  AOI21_X1 U14576 ( .B1(n18032), .B2(n18187), .A(n18020), .ZN(n11460) );
  OR2_X1 U14577 ( .A1(n18021), .A2(n18012), .ZN(n17589) );
  NAND2_X1 U14578 ( .A1(n18723), .A2(n18010), .ZN(n11477) );
  OAI21_X1 U14579 ( .B1(n11460), .B2(n17589), .A(n11477), .ZN(n17942) );
  NAND2_X1 U14580 ( .A1(n11461), .A2(n17942), .ZN(n17957) );
  NOR3_X1 U14581 ( .A1(n18218), .A2(n17549), .A3(n17957), .ZN(n11462) );
  NAND3_X1 U14582 ( .A1(n11467), .A2(n17540), .A3(n11466), .ZN(P3_U2834) );
  INV_X1 U14583 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16389) );
  NAND3_X1 U14584 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17805), .A3(
        n17553), .ZN(n15714) );
  NAND2_X1 U14585 ( .A1(n17552), .A2(n11468), .ZN(n15715) );
  NOR2_X1 U14586 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15715), .ZN(
        n11472) );
  NOR2_X1 U14587 ( .A1(n11469), .A2(n11472), .ZN(n15773) );
  NOR2_X1 U14588 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15773), .ZN(
        n15772) );
  INV_X1 U14589 ( .A(n11471), .ZN(n11470) );
  INV_X1 U14590 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18863) );
  AOI22_X1 U14591 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17805), .B1(
        n17737), .B2(n18863), .ZN(n11473) );
  NAND2_X1 U14592 ( .A1(n11470), .A2(n11473), .ZN(n11474) );
  NAND2_X1 U14593 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18863), .ZN(
        n11478) );
  NOR2_X1 U14594 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18863), .ZN(
        n11485) );
  NAND2_X1 U14595 ( .A1(n16383), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11482) );
  NOR2_X1 U14596 ( .A1(n11482), .A2(n17545), .ZN(n16387) );
  NAND2_X1 U14597 ( .A1(n16387), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11475) );
  XNOR2_X1 U14598 ( .A(n11475), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11495) );
  OAI221_X1 U14599 ( .B1(n18219), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C1(
        n18219), .C2(n9640), .A(n17906), .ZN(n11476) );
  OAI21_X1 U14600 ( .B1(n17598), .B2(n11477), .A(n11476), .ZN(n17928) );
  NAND3_X1 U14601 ( .A1(n16383), .A2(n17558), .A3(n17928), .ZN(n15717) );
  NOR3_X1 U14602 ( .A1(n16389), .A2(n11478), .A3(n15717), .ZN(n11480) );
  NOR2_X1 U14603 ( .A1(n18091), .A2(n11499), .ZN(n11479) );
  AOI211_X1 U14604 ( .C1(n11495), .C2(n18074), .A(n11480), .B(n11479), .ZN(
        n11481) );
  INV_X1 U14605 ( .A(n18125), .ZN(n18059) );
  NOR2_X1 U14606 ( .A1(n18059), .A2(n18218), .ZN(n18126) );
  AOI21_X1 U14607 ( .B1(n18126), .B2(n11482), .A(n18186), .ZN(n11483) );
  OAI21_X1 U14608 ( .B1(n11484), .B2(n18218), .A(n11483), .ZN(n15776) );
  INV_X1 U14609 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18837) );
  NOR2_X1 U14610 ( .A1(n18837), .A2(n18217), .ZN(n11494) );
  AOI21_X1 U14611 ( .B1(n11485), .B2(n18126), .A(n11494), .ZN(n11486) );
  INV_X1 U14612 ( .A(n11486), .ZN(n11487) );
  AOI21_X1 U14613 ( .B1(n15776), .B2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n11487), .ZN(n11488) );
  NAND2_X1 U14614 ( .A1(n11490), .A2(n16530), .ZN(n17900) );
  NOR2_X1 U14615 ( .A1(n18865), .A2(n18905), .ZN(n17859) );
  NAND2_X1 U14616 ( .A1(n18749), .A2(n18854), .ZN(n16505) );
  AND2_X1 U14617 ( .A1(n18868), .A2(n16505), .ZN(n18900) );
  NOR2_X4 U14618 ( .A1(n18865), .A2(n17891), .ZN(n17644) );
  INV_X1 U14619 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17889) );
  NAND2_X1 U14620 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17858) );
  INV_X1 U14621 ( .A(n17858), .ZN(n16844) );
  NAND2_X1 U14622 ( .A1(n16844), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17843) );
  NAND2_X1 U14623 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17796) );
  INV_X1 U14624 ( .A(n17796), .ZN(n17784) );
  NAND2_X1 U14625 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17730) );
  NAND2_X1 U14626 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17689) );
  NAND2_X1 U14627 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17652) );
  NAND2_X1 U14628 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17616) );
  NAND2_X1 U14629 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17581) );
  NAND2_X1 U14630 ( .A1(n17563), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17538) );
  NAND2_X1 U14631 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17539) );
  INV_X1 U14632 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16574) );
  NOR2_X1 U14633 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18749), .ZN(n17725) );
  NOR2_X1 U14634 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18854), .ZN(
        n18881) );
  INV_X1 U14635 ( .A(n18881), .ZN(n18867) );
  OAI221_X1 U14636 ( .B1(n18749), .B2(P3_STATE2_REG_1__SCAN_IN), .C1(
        P3_STATE2_REG_2__SCAN_IN), .C2(n18865), .A(n18867), .ZN(n18232) );
  NOR3_X2 U14637 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n18905), .ZN(n18585) );
  INV_X2 U14638 ( .A(n18263), .ZN(n18257) );
  OR2_X1 U14639 ( .A1(n11491), .A2(n17729), .ZN(n16376) );
  INV_X1 U14640 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16532) );
  XOR2_X1 U14641 ( .A(n16532), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n11492) );
  NOR2_X1 U14642 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17642), .ZN(
        n16392) );
  AND2_X1 U14643 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17563), .ZN(
        n17532) );
  NAND2_X1 U14644 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17532), .ZN(
        n16541) );
  NOR2_X1 U14645 ( .A1(n17539), .A2(n16541), .ZN(n16390) );
  INV_X1 U14646 ( .A(n17725), .ZN(n17896) );
  NAND2_X1 U14647 ( .A1(n18257), .A2(n11491), .ZN(n16396) );
  OAI211_X1 U14648 ( .C1(n16390), .C2(n17896), .A(n17897), .B(n16396), .ZN(
        n16399) );
  NOR2_X1 U14649 ( .A1(n16392), .A2(n16399), .ZN(n16375) );
  OAI22_X1 U14650 ( .A1(n16376), .A2(n11492), .B1(n16375), .B2(n16532), .ZN(
        n11493) );
  AOI211_X1 U14651 ( .C1(n17644), .C2(n16846), .A(n11494), .B(n11493), .ZN(
        n11497) );
  NOR2_X2 U14652 ( .A1(n17381), .A2(n17900), .ZN(n17761) );
  NAND2_X1 U14653 ( .A1(n11495), .A2(n17761), .ZN(n11496) );
  AOI21_X1 U14654 ( .B1(n11501), .B2(n17806), .A(n11500), .ZN(n11502) );
  INV_X1 U14655 ( .A(n11502), .ZN(P3_U2799) );
  AOI22_X1 U14656 ( .A1(n11588), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11587), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11509) );
  AOI22_X1 U14657 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11993), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11508) );
  AOI22_X1 U14658 ( .A1(n12260), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11846), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11507) );
  AND2_X4 U14659 ( .A1(n11513), .A2(n11505), .ZN(n11631) );
  AOI22_X1 U14660 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12259), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11506) );
  AOI22_X1 U14661 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11664), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11520) );
  INV_X2 U14662 ( .A(n12141), .ZN(n11930) );
  AOI22_X1 U14663 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11879), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11519) );
  AOI22_X1 U14664 ( .A1(n12232), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9661), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11518) );
  AOI22_X1 U14665 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11517) );
  AOI22_X1 U14666 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11993), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11524) );
  AOI22_X1 U14667 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U14668 ( .A1(n12260), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11846), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11522) );
  NAND4_X1 U14669 ( .A1(n11524), .A2(n11523), .A3(n11522), .A4(n11521), .ZN(
        n11530) );
  AOI22_X1 U14670 ( .A1(n9660), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11528) );
  AOI22_X1 U14671 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11664), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U14672 ( .A1(n12232), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11570), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U14673 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11879), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11525) );
  NAND4_X1 U14674 ( .A1(n11528), .A2(n11527), .A3(n11526), .A4(n11525), .ZN(
        n11529) );
  AOI22_X1 U14675 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U14676 ( .A1(n9659), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11879), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11534) );
  AOI22_X1 U14677 ( .A1(n12261), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11570), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11533) );
  AOI22_X1 U14678 ( .A1(n9673), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11664), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11532) );
  AOI22_X1 U14679 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12259), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11539) );
  AOI22_X1 U14680 ( .A1(n12260), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11846), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11538) );
  NAND2_X1 U14681 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11537) );
  NAND2_X1 U14682 ( .A1(n11993), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11536) );
  AND3_X4 U14683 ( .A1(n11542), .A2(n11541), .A3(n11540), .ZN(n11612) );
  AOI22_X1 U14684 ( .A1(n9639), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11587), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11547) );
  AOI22_X1 U14685 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11993), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U14686 ( .A1(n9671), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11846), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11545) );
  AOI22_X1 U14687 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11544) );
  NAND4_X1 U14688 ( .A1(n11547), .A2(n11546), .A3(n11545), .A4(n11544), .ZN(
        n11553) );
  AOI22_X1 U14689 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11570), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U14690 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11550) );
  AOI22_X1 U14691 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11664), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U14692 ( .A1(n9661), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11879), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11548) );
  NAND4_X1 U14693 ( .A1(n11551), .A2(n11550), .A3(n11549), .A4(n11548), .ZN(
        n11552) );
  NAND2_X1 U14694 ( .A1(n11555), .A2(n11614), .ZN(n13315) );
  AOI22_X1 U14695 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11559) );
  AOI22_X1 U14696 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11846), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11558) );
  NAND2_X1 U14697 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n11557) );
  NAND2_X1 U14698 ( .A1(n11993), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11556) );
  AOI22_X1 U14699 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11570), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U14700 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11562) );
  AOI22_X1 U14701 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11664), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U14702 ( .A1(n9659), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11879), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11560) );
  AOI22_X1 U14703 ( .A1(n9639), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11587), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U14704 ( .A1(n11588), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11587), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U14705 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11993), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11568) );
  AOI22_X1 U14706 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11846), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11567) );
  AOI22_X1 U14707 ( .A1(n12089), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11566) );
  AOI22_X1 U14708 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11570), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11575) );
  AOI22_X1 U14709 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11574) );
  AOI22_X1 U14710 ( .A1(n9673), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11664), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11573) );
  AOI22_X1 U14711 ( .A1(n9659), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11879), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11572) );
  NAND2_X1 U14712 ( .A1(n13336), .A2(n13725), .ZN(n11597) );
  NAND2_X1 U14713 ( .A1(n11993), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11578) );
  AOI22_X1 U14714 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11581) );
  NAND2_X1 U14715 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11580) );
  AOI22_X1 U14716 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11846), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U14717 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11570), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11585) );
  INV_X4 U14718 ( .A(n12184), .ZN(n12213) );
  AOI22_X1 U14719 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14720 ( .A1(n9673), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11664), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U14721 ( .A1(n9660), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11879), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U14722 ( .A1(n11588), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11587), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11592) );
  AOI22_X1 U14723 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11993), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11591) );
  AOI22_X1 U14724 ( .A1(n9671), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11846), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11590) );
  AOI22_X1 U14725 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11589) );
  AOI22_X1 U14726 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11664), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U14727 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9660), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U14728 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11879), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11594) );
  AOI22_X1 U14729 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11593) );
  INV_X1 U14730 ( .A(n11597), .ZN(n11598) );
  INV_X1 U14731 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n11603) );
  XNOR2_X1 U14732 ( .A(n11603), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n12454) );
  NAND2_X1 U14733 ( .A1(n11605), .A2(n20220), .ZN(n11609) );
  INV_X1 U14734 ( .A(n11724), .ZN(n11717) );
  OAI21_X1 U14735 ( .B1(n11608), .B2(n11609), .A(n11717), .ZN(n11619) );
  NAND2_X1 U14736 ( .A1(n13654), .A2(n13561), .ZN(n11611) );
  NOR2_X1 U14737 ( .A1(n13770), .A2(n11612), .ZN(n11613) );
  INV_X1 U14738 ( .A(n11614), .ZN(n11623) );
  NAND2_X1 U14739 ( .A1(n12599), .A2(n11612), .ZN(n11615) );
  INV_X1 U14740 ( .A(n11629), .ZN(n11616) );
  NAND2_X1 U14741 ( .A1(n12446), .A2(n12592), .ZN(n13322) );
  NAND2_X1 U14742 ( .A1(n11617), .A2(n13322), .ZN(n11618) );
  NAND2_X1 U14743 ( .A1(n16053), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20775) );
  INV_X1 U14744 ( .A(n20775), .ZN(n11620) );
  NAND2_X1 U14745 ( .A1(n20857), .A2(n16055), .ZN(n12580) );
  MUX2_X1 U14746 ( .A(n11620), .B(n12580), .S(n20634), .Z(n11621) );
  NAND2_X1 U14747 ( .A1(n13804), .A2(n11622), .ZN(n13328) );
  NAND2_X1 U14748 ( .A1(n11623), .A2(n20873), .ZN(n11624) );
  AND2_X1 U14749 ( .A1(n20857), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19978) );
  NAND4_X1 U14750 ( .A1(n13328), .A2(n11624), .A3(n19978), .A4(n13927), .ZN(
        n11625) );
  NAND3_X1 U14751 ( .A1(n13417), .A2(n12599), .A3(n20227), .ZN(n11626) );
  NAND2_X1 U14752 ( .A1(n11608), .A2(n11626), .ZN(n11627) );
  INV_X1 U14753 ( .A(n11679), .ZN(n11630) );
  AOI22_X1 U14754 ( .A1(n12237), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11631), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U14755 ( .A1(n12094), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9661), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11634) );
  AOI22_X1 U14756 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11633) );
  AOI22_X1 U14757 ( .A1(n12232), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11632) );
  AND4_X1 U14758 ( .A1(n11635), .A2(n11634), .A3(n11633), .A4(n11632), .ZN(
        n11642) );
  AOI22_X1 U14759 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12259), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11639) );
  AOI22_X1 U14760 ( .A1(n9671), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11846), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11638) );
  NAND2_X1 U14761 ( .A1(n12208), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11637) );
  NAND2_X1 U14762 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11636) );
  AOI22_X1 U14763 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n12231), .B1(
        n11643), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11640) );
  AOI22_X1 U14764 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U14765 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14766 ( .A1(n9671), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11846), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14767 ( .A1(n12237), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12094), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11644) );
  NAND4_X1 U14768 ( .A1(n11647), .A2(n11646), .A3(n11645), .A4(n11644), .ZN(
        n11653) );
  AOI22_X1 U14769 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14770 ( .A1(n9659), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11650) );
  AOI22_X1 U14771 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11649) );
  AOI22_X1 U14772 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11648) );
  NAND4_X1 U14773 ( .A1(n11651), .A2(n11650), .A3(n11649), .A4(n11648), .ZN(
        n11652) );
  XNOR2_X1 U14774 ( .A(n11656), .B(n12569), .ZN(n11654) );
  NAND2_X1 U14775 ( .A1(n11654), .A2(n11684), .ZN(n11655) );
  INV_X1 U14776 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20218) );
  AOI21_X1 U14777 ( .B1(n20212), .B2(n12513), .A(n16055), .ZN(n11658) );
  NAND2_X1 U14778 ( .A1(n11612), .A2(n12569), .ZN(n11657) );
  INV_X1 U14779 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11673) );
  AOI22_X1 U14780 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11663) );
  AOI22_X1 U14781 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11662) );
  AOI22_X1 U14782 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11661) );
  AOI22_X1 U14783 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12259), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11660) );
  NAND4_X1 U14784 ( .A1(n11663), .A2(n11662), .A3(n11661), .A4(n11660), .ZN(
        n11670) );
  AOI22_X1 U14785 ( .A1(n12237), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11668) );
  AOI22_X1 U14786 ( .A1(n12232), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11631), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U14787 ( .A1(n12094), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11666) );
  AOI22_X1 U14788 ( .A1(n9660), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11665) );
  NAND4_X1 U14789 ( .A1(n11668), .A2(n11667), .A3(n11666), .A4(n11665), .ZN(
        n11669) );
  NAND2_X1 U14790 ( .A1(n11717), .A2(n12514), .ZN(n11672) );
  OR2_X1 U14791 ( .A1(n12496), .A2(n12569), .ZN(n11671) );
  OAI211_X1 U14792 ( .C1(n12315), .C2(n11673), .A(n11672), .B(n11671), .ZN(
        n11674) );
  NAND2_X1 U14793 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11695) );
  OAI21_X1 U14794 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11695), .ZN(n20512) );
  NAND2_X1 U14795 ( .A1(n20775), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11688) );
  OAI21_X1 U14796 ( .B1(n12580), .B2(n20512), .A(n11688), .ZN(n11675) );
  INV_X1 U14797 ( .A(n11675), .ZN(n11676) );
  AND2_X2 U14798 ( .A1(n11680), .A2(n11679), .ZN(n11681) );
  INV_X1 U14799 ( .A(n20315), .ZN(n11683) );
  INV_X1 U14800 ( .A(n11681), .ZN(n11682) );
  NAND2_X1 U14801 ( .A1(n11684), .A2(n12514), .ZN(n11685) );
  INV_X1 U14802 ( .A(n11677), .ZN(n11690) );
  NAND2_X1 U14803 ( .A1(n11688), .A2(n11514), .ZN(n11689) );
  NAND2_X1 U14804 ( .A1(n11690), .A2(n11689), .ZN(n11702) );
  NAND2_X1 U14805 ( .A1(n11691), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11693) );
  NAND2_X1 U14806 ( .A1(n20775), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11692) );
  INV_X1 U14807 ( .A(n12580), .ZN(n11721) );
  INV_X1 U14808 ( .A(n11695), .ZN(n11694) );
  NAND2_X1 U14809 ( .A1(n11694), .A2(n12312), .ZN(n20547) );
  NAND2_X1 U14810 ( .A1(n11695), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11696) );
  NAND2_X1 U14811 ( .A1(n20547), .A2(n11696), .ZN(n14097) );
  AND2_X1 U14812 ( .A1(n11721), .A2(n14097), .ZN(n11700) );
  INV_X1 U14813 ( .A(n11699), .ZN(n11703) );
  INV_X1 U14814 ( .A(n11700), .ZN(n11701) );
  NAND4_X1 U14815 ( .A1(n11704), .A2(n11703), .A3(n11702), .A4(n11701), .ZN(
        n11705) );
  AOI22_X1 U14816 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U14817 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11708) );
  AOI22_X1 U14818 ( .A1(n9671), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11707) );
  AOI22_X1 U14819 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11706) );
  NAND4_X1 U14820 ( .A1(n11709), .A2(n11708), .A3(n11707), .A4(n11706), .ZN(
        n11715) );
  AOI22_X1 U14821 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12237), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U14822 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U14823 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12094), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14824 ( .A1(n9661), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11710) );
  NAND4_X1 U14825 ( .A1(n11713), .A2(n11712), .A3(n11711), .A4(n11710), .ZN(
        n11714) );
  AOI22_X1 U14826 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11717), .B2(n11716), .ZN(n11718) );
  NAND2_X1 U14827 ( .A1(n11691), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11723) );
  INV_X1 U14828 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20546) );
  NOR3_X1 U14829 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12312), .A3(
        n20582), .ZN(n20431) );
  NAND2_X1 U14830 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20431), .ZN(
        n20427) );
  NAND2_X1 U14831 ( .A1(n20546), .A2(n20427), .ZN(n11720) );
  NAND3_X1 U14832 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20711) );
  INV_X1 U14833 ( .A(n20711), .ZN(n20720) );
  NAND2_X1 U14834 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20720), .ZN(
        n20708) );
  AOI22_X1 U14835 ( .A1(n11721), .A2(n20456), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20775), .ZN(n11722) );
  AOI22_X1 U14836 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11728) );
  AOI22_X1 U14837 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11727) );
  AOI22_X1 U14838 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11726) );
  AOI22_X1 U14839 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11725) );
  NAND4_X1 U14840 ( .A1(n11728), .A2(n11727), .A3(n11726), .A4(n11725), .ZN(
        n11734) );
  AOI22_X1 U14841 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12237), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11732) );
  AOI22_X1 U14842 ( .A1(n12094), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9661), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11731) );
  AOI22_X1 U14843 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11730) );
  AOI22_X1 U14844 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11729) );
  NAND4_X1 U14845 ( .A1(n11732), .A2(n11731), .A3(n11730), .A4(n11729), .ZN(
        n11733) );
  AOI22_X1 U14846 ( .A1(n12335), .A2(n12534), .B1(n12326), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11735) );
  AOI22_X1 U14847 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11739) );
  AOI22_X1 U14848 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11738) );
  AOI22_X1 U14849 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U14850 ( .A1(n12237), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9667), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11736) );
  NAND4_X1 U14851 ( .A1(n11739), .A2(n11738), .A3(n11737), .A4(n11736), .ZN(
        n11745) );
  AOI22_X1 U14852 ( .A1(n12094), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9659), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11743) );
  AOI22_X1 U14853 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11742) );
  AOI22_X1 U14854 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11741) );
  AOI22_X1 U14855 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11740) );
  NAND4_X1 U14856 ( .A1(n11743), .A2(n11742), .A3(n11741), .A4(n11740), .ZN(
        n11744) );
  NAND2_X1 U14857 ( .A1(n12335), .A2(n12542), .ZN(n11747) );
  NAND2_X1 U14858 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11746) );
  INV_X1 U14859 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20242) );
  AOI22_X1 U14860 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U14861 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11750) );
  AOI22_X1 U14862 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11749) );
  AOI22_X1 U14863 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12259), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11748) );
  NAND4_X1 U14864 ( .A1(n11751), .A2(n11750), .A3(n11749), .A4(n11748), .ZN(
        n11757) );
  AOI22_X1 U14865 ( .A1(n12232), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12237), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11755) );
  AOI22_X1 U14866 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11754) );
  AOI22_X1 U14867 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12094), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11753) );
  AOI22_X1 U14868 ( .A1(n9660), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11752) );
  NAND4_X1 U14869 ( .A1(n11755), .A2(n11754), .A3(n11753), .A4(n11752), .ZN(
        n11756) );
  AOI22_X1 U14870 ( .A1(n12335), .A2(n12550), .B1(n12326), .B2(
        P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11835) );
  AOI22_X1 U14871 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U14872 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11763) );
  AOI22_X1 U14873 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11762) );
  AOI22_X1 U14874 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11631), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11761) );
  NAND4_X1 U14875 ( .A1(n11764), .A2(n11763), .A3(n11762), .A4(n11761), .ZN(
        n11770) );
  AOI22_X1 U14876 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12237), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11768) );
  AOI22_X1 U14877 ( .A1(n9673), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11767) );
  AOI22_X1 U14878 ( .A1(n12094), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9659), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11766) );
  AOI22_X1 U14879 ( .A1(n12160), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11765) );
  NAND4_X1 U14880 ( .A1(n11768), .A2(n11767), .A3(n11766), .A4(n11765), .ZN(
        n11769) );
  AOI22_X1 U14881 ( .A1(n12335), .A2(n12560), .B1(n12326), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11781) );
  INV_X1 U14882 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14107) );
  NAND2_X1 U14883 ( .A1(n12335), .A2(n12569), .ZN(n11771) );
  OAI21_X1 U14884 ( .B1(n14107), .B2(n12315), .A(n11771), .ZN(n11772) );
  INV_X2 U14885 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n11773) );
  INV_X1 U14886 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11779) );
  NOR2_X1 U14887 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12275) );
  INV_X1 U14888 ( .A(n11816), .ZN(n11774) );
  INV_X1 U14889 ( .A(n11782), .ZN(n11777) );
  INV_X1 U14890 ( .A(n11861), .ZN(n11776) );
  OAI21_X1 U14891 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n11777), .A(
        n11776), .ZN(n20025) );
  AOI22_X1 U14892 ( .A1(n12350), .A2(n20025), .B1(n12277), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11778) );
  OAI21_X1 U14893 ( .B1(n10316), .B2(n11779), .A(n11778), .ZN(n11780) );
  INV_X1 U14894 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11784) );
  OAI21_X1 U14895 ( .B1(n11839), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n11782), .ZN(n20032) );
  AOI22_X1 U14896 ( .A1(n20032), .A2(n12350), .B1(n12277), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11783) );
  OAI21_X1 U14897 ( .B1(n10316), .B2(n11784), .A(n11783), .ZN(n11785) );
  NAND2_X1 U14898 ( .A1(n9956), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11828) );
  XNOR2_X1 U14899 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13967) );
  AOI21_X1 U14900 ( .B1(n12350), .B2(n13967), .A(n12277), .ZN(n11789) );
  NAND2_X1 U14901 ( .A1(n11987), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11788) );
  OAI211_X1 U14902 ( .C1(n11828), .C2(n11787), .A(n11789), .B(n11788), .ZN(
        n11790) );
  INV_X1 U14903 ( .A(n11790), .ZN(n11791) );
  NAND2_X1 U14904 ( .A1(n12277), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11811) );
  INV_X1 U14905 ( .A(n13849), .ZN(n11810) );
  NAND2_X1 U14906 ( .A1(n11792), .A2(n12512), .ZN(n11793) );
  NAND2_X1 U14907 ( .A1(n20283), .A2(n11971), .ZN(n11799) );
  AOI22_X1 U14908 ( .A1(n11987), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n11773), .ZN(n11797) );
  INV_X1 U14909 ( .A(n11828), .ZN(n11795) );
  NAND2_X1 U14910 ( .A1(n11795), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11796) );
  AND2_X1 U14911 ( .A1(n11797), .A2(n11796), .ZN(n11798) );
  NAND2_X1 U14912 ( .A1(n11799), .A2(n11798), .ZN(n13728) );
  NAND2_X1 U14913 ( .A1(n12509), .A2(n11622), .ZN(n11802) );
  NAND2_X1 U14914 ( .A1(n11802), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13723) );
  INV_X1 U14915 ( .A(n9664), .ZN(n13846) );
  NAND2_X1 U14916 ( .A1(n11773), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11805) );
  NAND2_X1 U14917 ( .A1(n11987), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11804) );
  OAI211_X1 U14918 ( .C1(n11828), .C2(n13576), .A(n11805), .B(n11804), .ZN(
        n11806) );
  AOI21_X1 U14919 ( .B1(n9664), .B2(n11971), .A(n11806), .ZN(n13724) );
  OR2_X1 U14920 ( .A1(n13723), .A2(n13724), .ZN(n13721) );
  INV_X1 U14921 ( .A(n13724), .ZN(n11807) );
  NAND2_X1 U14922 ( .A1(n13721), .A2(n11808), .ZN(n13727) );
  NAND2_X1 U14923 ( .A1(n13728), .A2(n13727), .ZN(n13850) );
  NAND2_X1 U14924 ( .A1(n11810), .A2(n11809), .ZN(n13851) );
  INV_X1 U14925 ( .A(n13866), .ZN(n13868) );
  INV_X1 U14926 ( .A(n14089), .ZN(n11814) );
  INV_X1 U14927 ( .A(n11815), .ZN(n11831) );
  INV_X1 U14928 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11817) );
  NAND2_X1 U14929 ( .A1(n11817), .A2(n11816), .ZN(n11818) );
  NAND2_X1 U14930 ( .A1(n11831), .A2(n11818), .ZN(n14157) );
  AOI22_X1 U14931 ( .A1(n14157), .A2(n12350), .B1(n12277), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11820) );
  NAND2_X1 U14932 ( .A1(n11987), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11819) );
  OAI211_X1 U14933 ( .C1(n11828), .C2(n13807), .A(n11820), .B(n11819), .ZN(
        n11821) );
  INV_X1 U14934 ( .A(n11821), .ZN(n11822) );
  INV_X1 U14935 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12327) );
  NAND2_X1 U14936 ( .A1(n11773), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11827) );
  NAND2_X1 U14937 ( .A1(n11987), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11826) );
  OAI211_X1 U14938 ( .C1(n11828), .C2(n12327), .A(n11827), .B(n11826), .ZN(
        n11833) );
  INV_X1 U14939 ( .A(n11829), .ZN(n11841) );
  INV_X1 U14940 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11830) );
  NAND2_X1 U14941 ( .A1(n11831), .A2(n11830), .ZN(n11832) );
  NAND2_X1 U14942 ( .A1(n11841), .A2(n11832), .ZN(n20160) );
  MUX2_X1 U14943 ( .A(n11833), .B(n20160), .S(n12350), .Z(n11834) );
  NAND2_X1 U14944 ( .A1(n11836), .A2(n11835), .ZN(n11837) );
  NAND2_X1 U14945 ( .A1(n11838), .A2(n11837), .ZN(n12546) );
  INV_X1 U14946 ( .A(n11839), .ZN(n11843) );
  INV_X1 U14947 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11840) );
  NAND2_X1 U14948 ( .A1(n11841), .A2(n11840), .ZN(n11842) );
  NAND2_X1 U14949 ( .A1(n11843), .A2(n11842), .ZN(n20052) );
  AOI22_X1 U14950 ( .A1(n20052), .A2(n12275), .B1(n12277), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11845) );
  NAND2_X1 U14951 ( .A1(n11987), .A2(P1_EAX_REG_5__SCAN_IN), .ZN(n11844) );
  NAND2_X1 U14952 ( .A1(n11987), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11860) );
  XNOR2_X1 U14953 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n11861), .ZN(
        n20009) );
  AOI22_X1 U14954 ( .A1(n12350), .A2(n20009), .B1(n12277), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11859) );
  AOI22_X1 U14955 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n11643), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U14956 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n11543), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U14957 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U14958 ( .A1(n12094), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12259), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11847) );
  NAND4_X1 U14959 ( .A1(n11850), .A2(n11849), .A3(n11848), .A4(n11847), .ZN(
        n11856) );
  AOI22_X1 U14960 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n12237), .B1(
        n9659), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11854) );
  AOI22_X1 U14961 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11631), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11853) );
  AOI22_X1 U14962 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11852) );
  AOI22_X1 U14963 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11851) );
  NAND4_X1 U14964 ( .A1(n11854), .A2(n11853), .A3(n11852), .A4(n11851), .ZN(
        n11855) );
  NOR2_X1 U14965 ( .A1(n11856), .A2(n11855), .ZN(n11857) );
  OR2_X1 U14966 ( .A1(n11955), .A2(n11857), .ZN(n11858) );
  XNOR2_X1 U14967 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11887), .ZN(
        n20002) );
  AOI22_X1 U14968 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11865) );
  AOI22_X1 U14969 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11864) );
  AOI22_X1 U14970 ( .A1(n9671), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11863) );
  AOI22_X1 U14971 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12259), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11862) );
  NAND4_X1 U14972 ( .A1(n11865), .A2(n11864), .A3(n11863), .A4(n11862), .ZN(
        n11871) );
  AOI22_X1 U14973 ( .A1(n12237), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11631), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11869) );
  AOI22_X1 U14974 ( .A1(n12094), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9660), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11868) );
  AOI22_X1 U14975 ( .A1(n9673), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11867) );
  AOI22_X1 U14976 ( .A1(n12232), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11866) );
  NAND4_X1 U14977 ( .A1(n11869), .A2(n11868), .A3(n11867), .A4(n11866), .ZN(
        n11870) );
  OR2_X1 U14978 ( .A1(n11871), .A2(n11870), .ZN(n11872) );
  AOI22_X1 U14979 ( .A1(n11971), .A2(n11872), .B1(n12277), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11874) );
  NAND2_X1 U14980 ( .A1(n11987), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11873) );
  OAI211_X1 U14981 ( .C1(n20002), .C2(n12056), .A(n11874), .B(n11873), .ZN(
        n14193) );
  AOI22_X1 U14982 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U14983 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U14984 ( .A1(n12260), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11876) );
  AOI22_X1 U14985 ( .A1(n12232), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11631), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11875) );
  NAND4_X1 U14986 ( .A1(n11878), .A2(n11877), .A3(n11876), .A4(n11875), .ZN(
        n11885) );
  AOI22_X1 U14987 ( .A1(n12237), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9667), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11883) );
  AOI22_X1 U14988 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9661), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11882) );
  AOI22_X1 U14989 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11881) );
  AOI22_X1 U14990 ( .A1(n12094), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11880) );
  NAND4_X1 U14991 ( .A1(n11883), .A2(n11882), .A3(n11881), .A4(n11880), .ZN(
        n11884) );
  NOR2_X1 U14992 ( .A1(n11885), .A2(n11884), .ZN(n11890) );
  XNOR2_X1 U14993 ( .A(n11891), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14700) );
  NAND2_X1 U14994 ( .A1(n14700), .A2(n12275), .ZN(n11889) );
  AOI22_X1 U14995 ( .A1(n11987), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n12277), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11888) );
  OAI211_X1 U14996 ( .C1(n11890), .C2(n11955), .A(n11889), .B(n11888), .ZN(
        n14209) );
  INV_X1 U14997 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11895) );
  INV_X1 U14998 ( .A(n12277), .ZN(n11894) );
  OAI21_X1 U14999 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11892), .A(
        n11937), .ZN(n15890) );
  NAND2_X1 U15000 ( .A1(n15890), .A2(n12275), .ZN(n11893) );
  OAI21_X1 U15001 ( .B1(n11895), .B2(n11894), .A(n11893), .ZN(n11896) );
  AOI21_X1 U15002 ( .B1(n11987), .B2(P1_EAX_REG_11__SCAN_IN), .A(n11896), .ZN(
        n11897) );
  INV_X1 U15003 ( .A(n14471), .ZN(n11910) );
  AOI22_X1 U15004 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11901) );
  AOI22_X1 U15005 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11900) );
  AOI22_X1 U15006 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11899) );
  AOI22_X1 U15007 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11898) );
  NAND4_X1 U15008 ( .A1(n11901), .A2(n11900), .A3(n11899), .A4(n11898), .ZN(
        n11907) );
  AOI22_X1 U15009 ( .A1(n9673), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9667), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U15010 ( .A1(n12237), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12094), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U15011 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11903) );
  AOI22_X1 U15012 ( .A1(n9661), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11902) );
  NAND4_X1 U15013 ( .A1(n11905), .A2(n11904), .A3(n11903), .A4(n11902), .ZN(
        n11906) );
  NOR2_X1 U15014 ( .A1(n11907), .A2(n11906), .ZN(n11908) );
  OR2_X1 U15015 ( .A1(n11955), .A2(n11908), .ZN(n14472) );
  NAND2_X1 U15016 ( .A1(n11910), .A2(n11909), .ZN(n14474) );
  AOI22_X1 U15017 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11915) );
  AOI22_X1 U15018 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U15019 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11913) );
  AOI22_X1 U15020 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11912) );
  NAND4_X1 U15021 ( .A1(n11915), .A2(n11914), .A3(n11913), .A4(n11912), .ZN(
        n11921) );
  AOI22_X1 U15022 ( .A1(n12237), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11631), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11919) );
  AOI22_X1 U15023 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12094), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11918) );
  AOI22_X1 U15024 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9659), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11917) );
  AOI22_X1 U15025 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11916) );
  NAND4_X1 U15026 ( .A1(n11919), .A2(n11918), .A3(n11917), .A4(n11916), .ZN(
        n11920) );
  NOR2_X1 U15027 ( .A1(n11921), .A2(n11920), .ZN(n11925) );
  NAND2_X1 U15028 ( .A1(n11987), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11924) );
  XNOR2_X1 U15029 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11937), .ZN(
        n15879) );
  INV_X1 U15030 ( .A(n15879), .ZN(n11922) );
  AOI22_X1 U15031 ( .A1(n12277), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n12350), .B2(n11922), .ZN(n11923) );
  OAI211_X1 U15032 ( .C1(n11955), .C2(n11925), .A(n11924), .B(n11923), .ZN(
        n14558) );
  AOI22_X1 U15033 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11929) );
  AOI22_X1 U15034 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11928) );
  AOI22_X1 U15035 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11927) );
  AOI22_X1 U15036 ( .A1(n12232), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12259), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11926) );
  NAND4_X1 U15037 ( .A1(n11929), .A2(n11928), .A3(n11927), .A4(n11926), .ZN(
        n11936) );
  AOI22_X1 U15038 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11631), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11934) );
  AOI22_X1 U15039 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12094), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U15040 ( .A1(n9661), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11932) );
  AOI22_X1 U15041 ( .A1(n12237), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11931) );
  NAND4_X1 U15042 ( .A1(n11934), .A2(n11933), .A3(n11932), .A4(n11931), .ZN(
        n11935) );
  NOR2_X1 U15043 ( .A1(n11936), .A2(n11935), .ZN(n11941) );
  NAND2_X1 U15044 ( .A1(n11987), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11940) );
  INV_X1 U15045 ( .A(n11942), .ZN(n11938) );
  XNOR2_X1 U15046 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n11938), .ZN(
        n14692) );
  AOI22_X1 U15047 ( .A1(n12275), .A2(n14692), .B1(n12277), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11939) );
  OAI211_X1 U15048 ( .C1(n11955), .C2(n11941), .A(n11940), .B(n11939), .ZN(
        n14401) );
  INV_X1 U15049 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15830) );
  XNOR2_X1 U15050 ( .A(n15830), .B(n11959), .ZN(n15868) );
  INV_X1 U15051 ( .A(n15868), .ZN(n11958) );
  AOI22_X1 U15052 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11946) );
  AOI22_X1 U15053 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11945) );
  AOI22_X1 U15054 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11944) );
  AOI22_X1 U15055 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11631), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11943) );
  NAND4_X1 U15056 ( .A1(n11946), .A2(n11945), .A3(n11944), .A4(n11943), .ZN(
        n11952) );
  AOI22_X1 U15057 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12237), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U15058 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U15059 ( .A1(n12094), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9660), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U15060 ( .A1(n12160), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11947) );
  NAND4_X1 U15061 ( .A1(n11950), .A2(n11949), .A3(n11948), .A4(n11947), .ZN(
        n11951) );
  NOR2_X1 U15062 ( .A1(n11952), .A2(n11951), .ZN(n11956) );
  NAND2_X1 U15063 ( .A1(n11987), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11954) );
  NAND2_X1 U15064 ( .A1(n12277), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11953) );
  OAI211_X1 U15065 ( .C1(n11956), .C2(n11955), .A(n11954), .B(n11953), .ZN(
        n11957) );
  AOI21_X1 U15066 ( .B1(n11958), .B2(n12275), .A(n11957), .ZN(n14463) );
  XNOR2_X1 U15067 ( .A(n11974), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15819) );
  AOI22_X1 U15068 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11963) );
  AOI22_X1 U15069 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U15070 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11961) );
  AOI22_X1 U15071 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11960) );
  NAND4_X1 U15072 ( .A1(n11963), .A2(n11962), .A3(n11961), .A4(n11960), .ZN(
        n11969) );
  AOI22_X1 U15073 ( .A1(n12237), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9674), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11967) );
  AOI22_X1 U15074 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11631), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11966) );
  AOI22_X1 U15075 ( .A1(n12094), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11965) );
  AOI22_X1 U15076 ( .A1(n9659), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11964) );
  NAND4_X1 U15077 ( .A1(n11967), .A2(n11966), .A3(n11965), .A4(n11964), .ZN(
        n11968) );
  OR2_X1 U15078 ( .A1(n11969), .A2(n11968), .ZN(n11970) );
  AOI22_X1 U15079 ( .A1(n11971), .A2(n11970), .B1(n12277), .B2(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11973) );
  NAND2_X1 U15080 ( .A1(n11987), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11972) );
  OAI211_X1 U15081 ( .C1(n15819), .C2(n12056), .A(n11973), .B(n11972), .ZN(
        n14459) );
  OR2_X1 U15082 ( .A1(n11975), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11976) );
  NAND2_X1 U15083 ( .A1(n11976), .A2(n12009), .ZN(n15867) );
  INV_X1 U15084 ( .A(n13571), .ZN(n13547) );
  AOI22_X1 U15085 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11587), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11980) );
  AOI22_X1 U15086 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n12208), .B1(
        n11543), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11979) );
  AOI22_X1 U15087 ( .A1(n9671), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11978) );
  AOI22_X1 U15088 ( .A1(n12237), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11977) );
  NAND4_X1 U15089 ( .A1(n11980), .A2(n11979), .A3(n11978), .A4(n11977), .ZN(
        n11986) );
  AOI22_X1 U15090 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11984) );
  AOI22_X1 U15091 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11983) );
  AOI22_X1 U15092 ( .A1(n12094), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11982) );
  AOI22_X1 U15093 ( .A1(n9661), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11981) );
  NAND4_X1 U15094 ( .A1(n11984), .A2(n11983), .A3(n11982), .A4(n11981), .ZN(
        n11985) );
  NOR2_X1 U15095 ( .A1(n11986), .A2(n11985), .ZN(n11990) );
  INV_X1 U15096 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20874) );
  OAI21_X1 U15097 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20874), .A(
        n11773), .ZN(n11989) );
  NAND2_X1 U15098 ( .A1(n11987), .A2(P1_EAX_REG_16__SCAN_IN), .ZN(n11988) );
  OAI211_X1 U15099 ( .C1(n12271), .C2(n11990), .A(n11989), .B(n11988), .ZN(
        n11991) );
  OAI21_X1 U15100 ( .B1(n15867), .B2(n12056), .A(n11991), .ZN(n14388) );
  AOI22_X1 U15101 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11997) );
  AOI22_X1 U15102 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11993), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11996) );
  AOI22_X1 U15103 ( .A1(n9671), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11995) );
  AOI22_X1 U15104 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11994) );
  NAND4_X1 U15105 ( .A1(n11997), .A2(n11996), .A3(n11995), .A4(n11994), .ZN(
        n12003) );
  AOI22_X1 U15106 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9661), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U15107 ( .A1(n12237), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12094), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U15108 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U15109 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11998) );
  NAND4_X1 U15110 ( .A1(n12001), .A2(n12000), .A3(n11999), .A4(n11998), .ZN(
        n12002) );
  OR2_X1 U15111 ( .A1(n12003), .A2(n12002), .ZN(n12007) );
  INV_X1 U15112 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14535) );
  INV_X1 U15113 ( .A(n12009), .ZN(n12004) );
  XNOR2_X1 U15114 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12004), .ZN(
        n14676) );
  AOI22_X1 U15115 ( .A1(n12275), .A2(n14676), .B1(n12277), .B2(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12005) );
  OAI21_X1 U15116 ( .B1(n10316), .B2(n14535), .A(n12005), .ZN(n12006) );
  AOI21_X1 U15117 ( .B1(n12245), .B2(n12007), .A(n12006), .ZN(n14374) );
  OR2_X1 U15118 ( .A1(n12010), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12011) );
  NAND2_X1 U15119 ( .A1(n12011), .A2(n12040), .ZN(n15813) );
  AOI22_X1 U15120 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11587), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U15121 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U15122 ( .A1(n9671), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U15123 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12012) );
  NAND4_X1 U15124 ( .A1(n12015), .A2(n12014), .A3(n12013), .A4(n12012), .ZN(
        n12021) );
  AOI22_X1 U15125 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12237), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U15126 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9667), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U15127 ( .A1(n12094), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9659), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U15128 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12016) );
  NAND4_X1 U15129 ( .A1(n12019), .A2(n12018), .A3(n12017), .A4(n12016), .ZN(
        n12020) );
  NOR2_X1 U15130 ( .A1(n12021), .A2(n12020), .ZN(n12023) );
  AOI22_X1 U15131 ( .A1(n11987), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n11773), .ZN(n12022) );
  OAI21_X1 U15132 ( .B1(n12271), .B2(n12023), .A(n12022), .ZN(n12024) );
  MUX2_X1 U15133 ( .A(n15813), .B(n12024), .S(n12056), .Z(n12025) );
  AOI22_X1 U15134 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11587), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12029) );
  AOI22_X1 U15135 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U15136 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U15137 ( .A1(n12237), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12026) );
  NAND4_X1 U15138 ( .A1(n12029), .A2(n12028), .A3(n12027), .A4(n12026), .ZN(
        n12035) );
  AOI22_X1 U15139 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12094), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12033) );
  AOI22_X1 U15140 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9661), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U15141 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12031) );
  AOI22_X1 U15142 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12030) );
  NAND4_X1 U15143 ( .A1(n12033), .A2(n12032), .A3(n12031), .A4(n12030), .ZN(
        n12034) );
  NOR2_X1 U15144 ( .A1(n12035), .A2(n12034), .ZN(n12037) );
  AOI22_X1 U15145 ( .A1(n11987), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n11773), .ZN(n12036) );
  OAI21_X1 U15146 ( .B1(n12271), .B2(n12037), .A(n12036), .ZN(n12039) );
  INV_X1 U15147 ( .A(n12040), .ZN(n12038) );
  XNOR2_X1 U15148 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n12038), .ZN(
        n14656) );
  MUX2_X1 U15149 ( .A(n12039), .B(n14656), .S(n12350), .Z(n14362) );
  NAND2_X1 U15150 ( .A1(n14360), .A2(n14362), .ZN(n14361) );
  INV_X1 U15151 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14369) );
  OR2_X1 U15152 ( .A1(n12041), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12042) );
  NAND2_X1 U15153 ( .A1(n12042), .A2(n12069), .ZN(n15857) );
  INV_X1 U15154 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14519) );
  AOI22_X1 U15155 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12094), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U15156 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12045) );
  AOI22_X1 U15157 ( .A1(n9659), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12044) );
  AOI22_X1 U15158 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12043) );
  NAND4_X1 U15159 ( .A1(n12046), .A2(n12045), .A3(n12044), .A4(n12043), .ZN(
        n12052) );
  AOI22_X1 U15160 ( .A1(n9658), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11587), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U15161 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12049) );
  AOI22_X1 U15162 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12048) );
  AOI22_X1 U15163 ( .A1(n12237), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12047) );
  NAND4_X1 U15164 ( .A1(n12050), .A2(n12049), .A3(n12048), .A4(n12047), .ZN(
        n12051) );
  OAI21_X1 U15165 ( .B1(n12052), .B2(n12051), .A(n12245), .ZN(n12054) );
  OAI21_X1 U15166 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20874), .A(
        n11773), .ZN(n12053) );
  OAI211_X1 U15167 ( .C1(n10316), .C2(n14519), .A(n12054), .B(n12053), .ZN(
        n12055) );
  OAI21_X1 U15168 ( .B1(n15857), .B2(n12056), .A(n12055), .ZN(n14444) );
  AOI22_X1 U15169 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12060) );
  AOI22_X1 U15170 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12059) );
  AOI22_X1 U15171 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12058) );
  AOI22_X1 U15172 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12094), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12057) );
  NAND4_X1 U15173 ( .A1(n12060), .A2(n12059), .A3(n12058), .A4(n12057), .ZN(
        n12066) );
  AOI22_X1 U15174 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9661), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U15175 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12063) );
  AOI22_X1 U15176 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U15177 ( .A1(n12237), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12061) );
  NAND4_X1 U15178 ( .A1(n12064), .A2(n12063), .A3(n12062), .A4(n12061), .ZN(
        n12065) );
  NOR2_X1 U15179 ( .A1(n12066), .A2(n12065), .ZN(n12068) );
  AOI22_X1 U15180 ( .A1(n11987), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n11773), .ZN(n12067) );
  OAI21_X1 U15181 ( .B1(n12271), .B2(n12068), .A(n12067), .ZN(n12070) );
  XNOR2_X1 U15182 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n12083), .ZN(
        n14647) );
  MUX2_X1 U15183 ( .A(n12070), .B(n14647), .S(n12350), .Z(n14348) );
  AOI22_X1 U15184 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11587), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12074) );
  AOI22_X1 U15185 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12073) );
  AOI22_X1 U15186 ( .A1(n9671), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12072) );
  AOI22_X1 U15187 ( .A1(n12237), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12071) );
  NAND4_X1 U15188 ( .A1(n12074), .A2(n12073), .A3(n12072), .A4(n12071), .ZN(
        n12080) );
  AOI22_X1 U15189 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11930), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15190 ( .A1(n12094), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9660), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12077) );
  AOI22_X1 U15191 ( .A1(n9673), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11631), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12076) );
  AOI22_X1 U15192 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12075) );
  NAND4_X1 U15193 ( .A1(n12078), .A2(n12077), .A3(n12076), .A4(n12075), .ZN(
        n12079) );
  NOR2_X1 U15194 ( .A1(n12080), .A2(n12079), .ZN(n12082) );
  AOI22_X1 U15195 ( .A1(n11987), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n11773), .ZN(n12081) );
  OAI21_X1 U15196 ( .B1(n12271), .B2(n12082), .A(n12081), .ZN(n12088) );
  INV_X1 U15197 ( .A(n12084), .ZN(n12086) );
  INV_X1 U15198 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12085) );
  NAND2_X1 U15199 ( .A1(n12086), .A2(n12085), .ZN(n12087) );
  NAND2_X1 U15200 ( .A1(n12129), .A2(n12087), .ZN(n14640) );
  MUX2_X1 U15201 ( .A(n12088), .B(n14640), .S(n12350), .Z(n14338) );
  AOI22_X1 U15202 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12093) );
  AOI22_X1 U15203 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12092) );
  AOI22_X1 U15204 ( .A1(n12259), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12091) );
  AOI22_X1 U15205 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11631), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12090) );
  NAND4_X1 U15206 ( .A1(n12093), .A2(n12092), .A3(n12091), .A4(n12090), .ZN(
        n12100) );
  AOI22_X1 U15207 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11760), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12098) );
  AOI22_X1 U15208 ( .A1(n12237), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12094), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U15209 ( .A1(n12208), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U15210 ( .A1(n9673), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9660), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12095) );
  NAND4_X1 U15211 ( .A1(n12098), .A2(n12097), .A3(n12096), .A4(n12095), .ZN(
        n12099) );
  NOR2_X1 U15212 ( .A1(n12100), .A2(n12099), .ZN(n12114) );
  AOI22_X1 U15213 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n11643), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12104) );
  AOI22_X1 U15214 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n12116), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12103) );
  AOI22_X1 U15215 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U15216 ( .A1(n12237), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12101) );
  NAND4_X1 U15217 ( .A1(n12104), .A2(n12103), .A3(n12102), .A4(n12101), .ZN(
        n12110) );
  AOI22_X1 U15218 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n11760), .B1(
        n11631), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12108) );
  AOI22_X1 U15219 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n12094), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12107) );
  AOI22_X1 U15220 ( .A1(n12232), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9661), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12106) );
  AOI22_X1 U15221 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12105) );
  NAND4_X1 U15222 ( .A1(n12108), .A2(n12107), .A3(n12106), .A4(n12105), .ZN(
        n12109) );
  NOR2_X1 U15223 ( .A1(n12110), .A2(n12109), .ZN(n12115) );
  XOR2_X1 U15224 ( .A(n12114), .B(n12115), .Z(n12112) );
  INV_X1 U15225 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14506) );
  INV_X1 U15226 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14328) );
  OAI22_X1 U15227 ( .A1(n10316), .A2(n14506), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14328), .ZN(n12111) );
  AOI21_X1 U15228 ( .B1(n12112), .B2(n12245), .A(n12111), .ZN(n12113) );
  XNOR2_X1 U15229 ( .A(n12129), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14327) );
  MUX2_X1 U15230 ( .A(n12113), .B(n14327), .S(n12350), .Z(n14323) );
  NOR2_X1 U15231 ( .A1(n12115), .A2(n12114), .ZN(n12135) );
  AOI22_X1 U15232 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12120) );
  AOI22_X1 U15233 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U15234 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12118) );
  AOI22_X1 U15235 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12259), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12117) );
  NAND4_X1 U15236 ( .A1(n12120), .A2(n12119), .A3(n12118), .A4(n12117), .ZN(
        n12126) );
  AOI22_X1 U15237 ( .A1(n12232), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12237), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12124) );
  AOI22_X1 U15238 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12123) );
  AOI22_X1 U15239 ( .A1(n9673), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12094), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U15240 ( .A1(n9660), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12121) );
  NAND4_X1 U15241 ( .A1(n12124), .A2(n12123), .A3(n12122), .A4(n12121), .ZN(
        n12125) );
  OR2_X1 U15242 ( .A1(n12126), .A2(n12125), .ZN(n12134) );
  XNOR2_X1 U15243 ( .A(n12135), .B(n12134), .ZN(n12128) );
  AOI22_X1 U15244 ( .A1(n11987), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n11773), .ZN(n12127) );
  OAI21_X1 U15245 ( .B1(n12128), .B2(n12271), .A(n12127), .ZN(n12133) );
  INV_X1 U15246 ( .A(n12130), .ZN(n12131) );
  INV_X1 U15247 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14618) );
  NAND2_X1 U15248 ( .A1(n12131), .A2(n14618), .ZN(n12132) );
  NAND2_X1 U15249 ( .A1(n12174), .A2(n12132), .ZN(n14315) );
  MUX2_X1 U15250 ( .A(n12133), .B(n14315), .S(n12350), .Z(n14311) );
  NAND2_X1 U15251 ( .A1(n12135), .A2(n12134), .ZN(n12158) );
  INV_X1 U15252 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12147) );
  INV_X1 U15253 ( .A(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12138) );
  INV_X1 U15254 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12136) );
  OAI22_X1 U15255 ( .A1(n12139), .A2(n12138), .B1(n12137), .B2(n12136), .ZN(
        n12144) );
  INV_X1 U15256 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12142) );
  INV_X1 U15257 ( .A(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12140) );
  OAI22_X1 U15258 ( .A1(n12188), .A2(n12142), .B1(n12141), .B2(n12140), .ZN(
        n12143) );
  AOI211_X1 U15259 ( .C1(n9658), .C2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n12144), .B(n12143), .ZN(n12146) );
  AOI22_X1 U15260 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12145) );
  OAI211_X1 U15261 ( .C1(n12258), .C2(n12147), .A(n12146), .B(n12145), .ZN(
        n12153) );
  AOI22_X1 U15262 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12151) );
  AOI22_X1 U15263 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12150) );
  AOI22_X1 U15264 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9659), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12149) );
  AOI22_X1 U15265 ( .A1(n12094), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12148) );
  NAND4_X1 U15266 ( .A1(n12151), .A2(n12150), .A3(n12149), .A4(n12148), .ZN(
        n12152) );
  NOR2_X1 U15267 ( .A1(n12153), .A2(n12152), .ZN(n12159) );
  XOR2_X1 U15268 ( .A(n12158), .B(n12159), .Z(n12156) );
  INV_X1 U15269 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n14497) );
  INV_X1 U15270 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12154) );
  OAI22_X1 U15271 ( .A1(n10316), .A2(n14497), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12154), .ZN(n12155) );
  AOI21_X1 U15272 ( .B1(n12156), .B2(n12245), .A(n12155), .ZN(n12157) );
  XNOR2_X1 U15273 ( .A(n12174), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14300) );
  MUX2_X1 U15274 ( .A(n12157), .B(n14300), .S(n12350), .Z(n14299) );
  NOR2_X1 U15275 ( .A1(n12159), .A2(n12158), .ZN(n12182) );
  AOI22_X1 U15276 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12164) );
  AOI22_X1 U15277 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12163) );
  AOI22_X1 U15278 ( .A1(n9671), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12162) );
  AOI22_X1 U15279 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12161) );
  NAND4_X1 U15280 ( .A1(n12164), .A2(n12163), .A3(n12162), .A4(n12161), .ZN(
        n12171) );
  AOI22_X1 U15281 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12237), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U15282 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U15283 ( .A1(n9673), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12094), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12167) );
  AOI22_X1 U15284 ( .A1(n9660), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12166) );
  NAND4_X1 U15285 ( .A1(n12169), .A2(n12168), .A3(n12167), .A4(n12166), .ZN(
        n12170) );
  OR2_X1 U15286 ( .A1(n12171), .A2(n12170), .ZN(n12181) );
  XNOR2_X1 U15287 ( .A(n12182), .B(n12181), .ZN(n12173) );
  AOI22_X1 U15288 ( .A1(n11987), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n11773), .ZN(n12172) );
  OAI21_X1 U15289 ( .B1(n12173), .B2(n12271), .A(n12172), .ZN(n12180) );
  INV_X1 U15290 ( .A(n12174), .ZN(n12175) );
  INV_X1 U15291 ( .A(n12176), .ZN(n12178) );
  INV_X1 U15292 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12177) );
  NAND2_X1 U15293 ( .A1(n12178), .A2(n12177), .ZN(n12179) );
  NAND2_X1 U15294 ( .A1(n12222), .A2(n12179), .ZN(n14603) );
  MUX2_X1 U15295 ( .A(n12180), .B(n14603), .S(n12350), .Z(n14283) );
  NAND2_X1 U15296 ( .A1(n12182), .A2(n12181), .ZN(n12206) );
  INV_X1 U15297 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12195) );
  INV_X1 U15298 ( .A(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12185) );
  INV_X1 U15299 ( .A(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12183) );
  OAI22_X1 U15300 ( .A1(n12186), .A2(n12185), .B1(n12184), .B2(n12183), .ZN(
        n12192) );
  INV_X1 U15301 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12189) );
  INV_X1 U15302 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12187) );
  OAI22_X1 U15303 ( .A1(n12190), .A2(n12189), .B1(n12188), .B2(n12187), .ZN(
        n12191) );
  AOI211_X1 U15304 ( .C1(n12231), .C2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n12192), .B(n12191), .ZN(n12194) );
  AOI22_X1 U15305 ( .A1(n9659), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12193) );
  OAI211_X1 U15306 ( .C1(n13803), .C2(n12195), .A(n12194), .B(n12193), .ZN(
        n12201) );
  AOI22_X1 U15307 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12199) );
  AOI22_X1 U15308 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12198) );
  AOI22_X1 U15309 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11631), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12197) );
  AOI22_X1 U15310 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12094), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12196) );
  NAND4_X1 U15311 ( .A1(n12199), .A2(n12198), .A3(n12197), .A4(n12196), .ZN(
        n12200) );
  NOR2_X1 U15312 ( .A1(n12201), .A2(n12200), .ZN(n12207) );
  XOR2_X1 U15313 ( .A(n12206), .B(n12207), .Z(n12204) );
  INV_X1 U15314 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14488) );
  INV_X1 U15315 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12202) );
  OAI22_X1 U15316 ( .A1(n10316), .A2(n14488), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12202), .ZN(n12203) );
  AOI21_X1 U15317 ( .B1(n12204), .B2(n12245), .A(n12203), .ZN(n12205) );
  XNOR2_X1 U15318 ( .A(n12222), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14592) );
  MUX2_X1 U15319 ( .A(n12205), .B(n14592), .S(n12350), .Z(n14273) );
  NOR2_X1 U15320 ( .A1(n12207), .A2(n12206), .ZN(n12230) );
  AOI22_X1 U15321 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U15322 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12211) );
  AOI22_X1 U15323 ( .A1(n9671), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U15324 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12209) );
  NAND4_X1 U15325 ( .A1(n12212), .A2(n12211), .A3(n12210), .A4(n12209), .ZN(
        n12219) );
  AOI22_X1 U15326 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12237), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12217) );
  AOI22_X1 U15327 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U15328 ( .A1(n9673), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12094), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12215) );
  AOI22_X1 U15329 ( .A1(n9660), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12214) );
  NAND4_X1 U15330 ( .A1(n12217), .A2(n12216), .A3(n12215), .A4(n12214), .ZN(
        n12218) );
  OR2_X1 U15331 ( .A1(n12219), .A2(n12218), .ZN(n12229) );
  XNOR2_X1 U15332 ( .A(n12230), .B(n12229), .ZN(n12221) );
  AOI22_X1 U15333 ( .A1(n11987), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n11773), .ZN(n12220) );
  OAI21_X1 U15334 ( .B1(n12221), .B2(n12271), .A(n12220), .ZN(n12228) );
  INV_X1 U15335 ( .A(n12222), .ZN(n12223) );
  INV_X1 U15336 ( .A(n12224), .ZN(n12226) );
  INV_X1 U15337 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12225) );
  NAND2_X1 U15338 ( .A1(n12226), .A2(n12225), .ZN(n12227) );
  NAND2_X1 U15339 ( .A1(n12274), .A2(n12227), .ZN(n14585) );
  MUX2_X1 U15340 ( .A(n12228), .B(n14585), .S(n12350), .Z(n14258) );
  NAND2_X1 U15341 ( .A1(n12230), .A2(n12229), .ZN(n12248) );
  AOI22_X1 U15342 ( .A1(n11643), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12236) );
  AOI22_X1 U15343 ( .A1(n12208), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12235) );
  AOI22_X1 U15344 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12260), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12234) );
  AOI22_X1 U15345 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12233) );
  NAND4_X1 U15346 ( .A1(n12236), .A2(n12235), .A3(n12234), .A4(n12233), .ZN(
        n12243) );
  AOI22_X1 U15347 ( .A1(n12237), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12241) );
  AOI22_X1 U15348 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12094), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12240) );
  AOI22_X1 U15349 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9660), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12239) );
  AOI22_X1 U15350 ( .A1(n12160), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12238) );
  NAND4_X1 U15351 ( .A1(n12241), .A2(n12240), .A3(n12239), .A4(n12238), .ZN(
        n12242) );
  NOR2_X1 U15352 ( .A1(n12243), .A2(n12242), .ZN(n12249) );
  XOR2_X1 U15353 ( .A(n12248), .B(n12249), .Z(n12246) );
  INV_X1 U15354 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n12612) );
  INV_X1 U15355 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12273) );
  OAI22_X1 U15356 ( .A1(n10316), .A2(n12612), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12273), .ZN(n12244) );
  AOI21_X1 U15357 ( .B1(n12246), .B2(n12245), .A(n12244), .ZN(n12247) );
  XNOR2_X1 U15358 ( .A(n12274), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14249) );
  MUX2_X1 U15359 ( .A(n12247), .B(n14249), .S(n12350), .Z(n12590) );
  NOR2_X1 U15360 ( .A1(n12249), .A2(n12248), .ZN(n12269) );
  INV_X1 U15361 ( .A(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12257) );
  INV_X1 U15362 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15363 ( .A1(n11631), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12250), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15364 ( .A1(n12094), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12251) );
  OAI211_X1 U15365 ( .C1(n13803), .C2(n12253), .A(n12252), .B(n12251), .ZN(
        n12254) );
  INV_X1 U15366 ( .A(n12254), .ZN(n12256) );
  AOI22_X1 U15367 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12255) );
  OAI211_X1 U15368 ( .C1(n12258), .C2(n12257), .A(n12256), .B(n12255), .ZN(
        n12267) );
  AOI22_X1 U15369 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12208), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15370 ( .A1(n9671), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12264) );
  AOI22_X1 U15371 ( .A1(n12237), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12263) );
  AOI22_X1 U15372 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9659), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12262) );
  NAND4_X1 U15373 ( .A1(n12265), .A2(n12264), .A3(n12263), .A4(n12262), .ZN(
        n12266) );
  NOR2_X1 U15374 ( .A1(n12267), .A2(n12266), .ZN(n12268) );
  XOR2_X1 U15375 ( .A(n12269), .B(n12268), .Z(n12272) );
  AOI22_X1 U15376 ( .A1(n11987), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n11773), .ZN(n12270) );
  OAI21_X1 U15377 ( .B1(n12272), .B2(n12271), .A(n12270), .ZN(n12276) );
  INV_X1 U15378 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12485) );
  XNOR2_X1 U15379 ( .A(n12353), .B(n12485), .ZN(n12583) );
  MUX2_X1 U15380 ( .A(n12276), .B(n12583), .S(n12275), .Z(n12479) );
  AOI22_X1 U15381 ( .A1(n11987), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n12277), .ZN(n12278) );
  INV_X1 U15382 ( .A(n12278), .ZN(n12279) );
  NAND2_X1 U15383 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20634), .ZN(
        n12290) );
  OAI21_X1 U15384 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20634), .A(
        n12290), .ZN(n12281) );
  INV_X1 U15385 ( .A(n12281), .ZN(n12284) );
  NAND2_X1 U15386 ( .A1(n12335), .A2(n12284), .ZN(n12282) );
  NAND2_X1 U15387 ( .A1(n12282), .A2(n12336), .ZN(n12286) );
  NAND2_X1 U15388 ( .A1(n11606), .A2(n13654), .ZN(n12283) );
  NAND2_X1 U15389 ( .A1(n12283), .A2(n20220), .ZN(n12305) );
  OAI211_X1 U15390 ( .C1(n13319), .C2(n20212), .A(n12305), .B(n12284), .ZN(
        n12285) );
  NAND2_X1 U15391 ( .A1(n12286), .A2(n12285), .ZN(n12295) );
  NAND2_X1 U15392 ( .A1(n11606), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12287) );
  INV_X1 U15393 ( .A(n12294), .ZN(n12293) );
  NAND2_X1 U15394 ( .A1(n20582), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12297) );
  NAND2_X1 U15395 ( .A1(n11687), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12289) );
  NAND2_X1 U15396 ( .A1(n12297), .A2(n12289), .ZN(n12291) );
  NAND2_X1 U15397 ( .A1(n12291), .A2(n12290), .ZN(n12292) );
  NAND2_X1 U15398 ( .A1(n12298), .A2(n12292), .ZN(n12343) );
  OAI211_X1 U15399 ( .C1(n12295), .C2(n12293), .A(n12343), .B(n12329), .ZN(
        n12304) );
  NOR2_X1 U15400 ( .A1(n12343), .A2(n12294), .ZN(n12296) );
  NAND2_X1 U15401 ( .A1(n12296), .A2(n12295), .ZN(n12303) );
  NAND2_X1 U15402 ( .A1(n12298), .A2(n12297), .ZN(n12311) );
  MUX2_X1 U15403 ( .A(n12312), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n12299) );
  XNOR2_X1 U15404 ( .A(n12311), .B(n12299), .ZN(n12345) );
  INV_X1 U15405 ( .A(n12345), .ZN(n12306) );
  NAND2_X1 U15406 ( .A1(n12335), .A2(n12306), .ZN(n12301) );
  NAND2_X1 U15407 ( .A1(n12326), .A2(n12345), .ZN(n12300) );
  NAND3_X1 U15408 ( .A1(n12301), .A2(n12305), .A3(n12300), .ZN(n12302) );
  NAND3_X1 U15409 ( .A1(n12304), .A2(n12303), .A3(n12302), .ZN(n12309) );
  INV_X1 U15410 ( .A(n12305), .ZN(n12307) );
  NAND3_X1 U15411 ( .A1(n12307), .A2(n12306), .A3(n12335), .ZN(n12308) );
  NAND2_X1 U15412 ( .A1(n12309), .A2(n12308), .ZN(n12317) );
  NAND2_X1 U15413 ( .A1(n12311), .A2(n12310), .ZN(n12314) );
  NAND2_X1 U15414 ( .A1(n12312), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12313) );
  NAND2_X1 U15415 ( .A1(n12314), .A2(n12313), .ZN(n12321) );
  XNOR2_X1 U15416 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12320) );
  XNOR2_X1 U15417 ( .A(n12321), .B(n12320), .ZN(n12344) );
  NAND2_X1 U15418 ( .A1(n12315), .A2(n12344), .ZN(n12316) );
  NAND2_X1 U15419 ( .A1(n12317), .A2(n12316), .ZN(n12325) );
  INV_X1 U15420 ( .A(n12336), .ZN(n12318) );
  NAND2_X1 U15421 ( .A1(n12318), .A2(n12344), .ZN(n12324) );
  NOR2_X1 U15422 ( .A1(n13807), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12319) );
  AOI21_X1 U15423 ( .B1(n12321), .B2(n12320), .A(n12319), .ZN(n12334) );
  NOR2_X1 U15424 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20210), .ZN(
        n12332) );
  AND2_X1 U15425 ( .A1(n12334), .A2(n12332), .ZN(n12346) );
  INV_X1 U15426 ( .A(n12346), .ZN(n12322) );
  NOR2_X1 U15427 ( .A1(n12326), .A2(n12322), .ZN(n12323) );
  AOI21_X1 U15428 ( .B1(n12325), .B2(n12324), .A(n12323), .ZN(n12331) );
  NAND2_X1 U15429 ( .A1(n12326), .A2(n12346), .ZN(n12328) );
  OAI22_X1 U15430 ( .A1(n12329), .A2(n12328), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n12327), .ZN(n12330) );
  NAND2_X1 U15431 ( .A1(n20210), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12333) );
  AOI21_X1 U15432 ( .B1(n12334), .B2(n12333), .A(n12332), .ZN(n12338) );
  AND2_X1 U15433 ( .A1(n12335), .A2(n12338), .ZN(n12337) );
  INV_X1 U15434 ( .A(n12338), .ZN(n12348) );
  OR4_X1 U15435 ( .A1(n12346), .A2(n12345), .A3(n12344), .A4(n12343), .ZN(
        n12347) );
  NAND2_X1 U15436 ( .A1(n12342), .A2(n13422), .ZN(n13415) );
  NOR2_X1 U15437 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20879) );
  NAND2_X1 U15438 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20879), .ZN(n15757) );
  AND2_X1 U15439 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n16055), .ZN(n12349) );
  NAND2_X1 U15440 ( .A1(n12350), .A2(n12349), .ZN(n12351) );
  OAI211_X1 U15441 ( .C1(n15757), .C2(n16055), .A(n20170), .B(n12351), .ZN(
        n12352) );
  INV_X1 U15442 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12354) );
  NAND2_X1 U15443 ( .A1(n13218), .A2(n20041), .ZN(n12478) );
  AOI22_X1 U15444 ( .A1(P1_EBX_REG_31__SCAN_IN), .A2(n12446), .B1(n12361), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12450) );
  NAND2_X1 U15445 ( .A1(n12446), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n12358) );
  NAND2_X1 U15446 ( .A1(n12361), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12357) );
  NAND2_X1 U15447 ( .A1(n12358), .A2(n12357), .ZN(n12482) );
  OR2_X1 U15448 ( .A1(n12443), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n12363) );
  INV_X1 U15449 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13911) );
  NAND2_X1 U15450 ( .A1(n9638), .A2(n13911), .ZN(n12359) );
  OAI211_X1 U15451 ( .C1(n12361), .C2(P1_EBX_REG_1__SCAN_IN), .A(n12360), .B(
        n12359), .ZN(n12362) );
  NAND2_X1 U15452 ( .A1(n12363), .A2(n12362), .ZN(n12365) );
  NAND2_X1 U15453 ( .A1(n9638), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12364) );
  OAI21_X1 U15454 ( .B1(n13412), .B2(P1_EBX_REG_0__SCAN_IN), .A(n12364), .ZN(
        n13711) );
  XNOR2_X1 U15455 ( .A(n12365), .B(n13711), .ZN(n13339) );
  NAND2_X1 U15456 ( .A1(n13339), .A2(n13717), .ZN(n13340) );
  OR2_X1 U15457 ( .A1(n12443), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n12368) );
  INV_X1 U15458 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20191) );
  NAND2_X1 U15459 ( .A1(n9638), .A2(n20191), .ZN(n12366) );
  OAI211_X1 U15460 ( .C1(n12361), .C2(P1_EBX_REG_2__SCAN_IN), .A(n12360), .B(
        n12366), .ZN(n12367) );
  MUX2_X1 U15461 ( .A(n12439), .B(n13412), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12371) );
  INV_X1 U15462 ( .A(n12371), .ZN(n12372) );
  OAI21_X1 U15463 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n12446), .A(
        n12372), .ZN(n13888) );
  MUX2_X1 U15464 ( .A(n12443), .B(n9638), .S(P1_EBX_REG_4__SCAN_IN), .Z(n12376) );
  INV_X1 U15465 ( .A(n9638), .ZN(n12373) );
  NAND2_X1 U15466 ( .A1(n12373), .A2(n12361), .ZN(n12415) );
  NAND2_X1 U15467 ( .A1(n12361), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12374) );
  AND2_X1 U15468 ( .A1(n12415), .A2(n12374), .ZN(n12375) );
  NAND2_X1 U15469 ( .A1(n12376), .A2(n12375), .ZN(n13909) );
  INV_X1 U15470 ( .A(n12439), .ZN(n12434) );
  NAND2_X1 U15471 ( .A1(n12360), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12377) );
  OAI211_X1 U15472 ( .C1(n12361), .C2(P1_EBX_REG_5__SCAN_IN), .A(n9638), .B(
        n12377), .ZN(n12378) );
  OAI21_X1 U15473 ( .B1(n12434), .B2(P1_EBX_REG_5__SCAN_IN), .A(n12378), .ZN(
        n16039) );
  INV_X1 U15474 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20033) );
  MUX2_X1 U15475 ( .A(n9638), .B(n12443), .S(n20033), .Z(n12381) );
  NAND2_X1 U15476 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12361), .ZN(
        n12379) );
  AND2_X1 U15477 ( .A1(n12415), .A2(n12379), .ZN(n12380) );
  NAND2_X1 U15478 ( .A1(n12381), .A2(n12380), .ZN(n16021) );
  INV_X1 U15479 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20068) );
  NAND2_X1 U15480 ( .A1(n12439), .A2(n20068), .ZN(n12384) );
  NAND2_X1 U15481 ( .A1(n12360), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12382) );
  OAI211_X1 U15482 ( .C1(n12361), .C2(P1_EBX_REG_7__SCAN_IN), .A(n9638), .B(
        n12382), .ZN(n12383) );
  INV_X1 U15483 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n20010) );
  MUX2_X1 U15484 ( .A(n9638), .B(n12443), .S(n20010), .Z(n12387) );
  NAND2_X1 U15485 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n12361), .ZN(
        n12385) );
  AND2_X1 U15486 ( .A1(n12415), .A2(n12385), .ZN(n12386) );
  INV_X1 U15487 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20064) );
  NAND2_X1 U15488 ( .A1(n12439), .A2(n20064), .ZN(n12390) );
  NAND2_X1 U15489 ( .A1(n12360), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12388) );
  OAI211_X1 U15490 ( .C1(n12361), .C2(P1_EBX_REG_9__SCAN_IN), .A(n9638), .B(
        n12388), .ZN(n12389) );
  AND2_X1 U15491 ( .A1(n12390), .A2(n12389), .ZN(n16010) );
  NAND2_X1 U15492 ( .A1(n16011), .A2(n16010), .ZN(n16013) );
  OR2_X1 U15493 ( .A1(n12443), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n12394) );
  INV_X1 U15494 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12391) );
  NAND2_X1 U15495 ( .A1(n9638), .A2(n12391), .ZN(n12392) );
  OAI211_X1 U15496 ( .C1(n12361), .C2(P1_EBX_REG_10__SCAN_IN), .A(n12360), .B(
        n12392), .ZN(n12393) );
  MUX2_X1 U15497 ( .A(n12439), .B(n13412), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12395) );
  INV_X1 U15498 ( .A(n12395), .ZN(n12396) );
  OAI21_X1 U15499 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n12446), .A(
        n12396), .ZN(n14475) );
  MUX2_X1 U15500 ( .A(n12439), .B(n13412), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n12398) );
  NOR2_X1 U15501 ( .A1(n12446), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12397) );
  NOR2_X1 U15502 ( .A1(n12398), .A2(n12397), .ZN(n14402) );
  OR2_X1 U15503 ( .A1(n12443), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n12401) );
  INV_X1 U15504 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14804) );
  NAND2_X1 U15505 ( .A1(n9638), .A2(n14804), .ZN(n12399) );
  OAI211_X1 U15506 ( .C1(n12361), .C2(P1_EBX_REG_12__SCAN_IN), .A(n12360), .B(
        n12399), .ZN(n12400) );
  NAND2_X1 U15507 ( .A1(n12401), .A2(n12400), .ZN(n15838) );
  AND2_X1 U15508 ( .A1(n14402), .A2(n15838), .ZN(n12402) );
  OR2_X1 U15509 ( .A1(n12443), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n12405) );
  INV_X1 U15510 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12501) );
  NAND2_X1 U15511 ( .A1(n9638), .A2(n12501), .ZN(n12403) );
  OAI211_X1 U15512 ( .C1(n12361), .C2(P1_EBX_REG_14__SCAN_IN), .A(n12360), .B(
        n12403), .ZN(n12404) );
  NAND2_X1 U15513 ( .A1(n12405), .A2(n12404), .ZN(n14464) );
  MUX2_X1 U15514 ( .A(n12439), .B(n13412), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12406) );
  INV_X1 U15515 ( .A(n12406), .ZN(n12408) );
  INV_X1 U15516 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14790) );
  INV_X1 U15517 ( .A(n12446), .ZN(n13713) );
  NAND2_X1 U15518 ( .A1(n14790), .A2(n13713), .ZN(n12407) );
  NAND2_X1 U15519 ( .A1(n12408), .A2(n12407), .ZN(n14461) );
  OR2_X1 U15520 ( .A1(n12443), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n12411) );
  INV_X1 U15521 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14802) );
  NAND2_X1 U15522 ( .A1(n9638), .A2(n14802), .ZN(n12409) );
  OAI211_X1 U15523 ( .C1(n12361), .C2(P1_EBX_REG_16__SCAN_IN), .A(n12360), .B(
        n12409), .ZN(n12410) );
  MUX2_X1 U15524 ( .A(n12439), .B(n13412), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12413) );
  NOR2_X1 U15525 ( .A1(n12446), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12412) );
  NOR2_X1 U15526 ( .A1(n12413), .A2(n12412), .ZN(n14380) );
  MUX2_X1 U15527 ( .A(n12443), .B(n9638), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n12417) );
  NAND2_X1 U15528 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n12361), .ZN(
        n12414) );
  AND2_X1 U15529 ( .A1(n12415), .A2(n12414), .ZN(n12416) );
  NAND2_X1 U15530 ( .A1(n12417), .A2(n12416), .ZN(n14449) );
  MUX2_X1 U15531 ( .A(n12439), .B(n13412), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12418) );
  INV_X1 U15532 ( .A(n12418), .ZN(n12419) );
  OAI21_X1 U15533 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n12446), .A(
        n12419), .ZN(n14364) );
  INV_X1 U15534 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n12420) );
  MUX2_X1 U15535 ( .A(n9638), .B(n12443), .S(n12420), .Z(n12422) );
  NAND2_X1 U15536 ( .A1(n12361), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12421) );
  AND2_X1 U15537 ( .A1(n12422), .A2(n12421), .ZN(n14440) );
  MUX2_X1 U15538 ( .A(n12439), .B(n13412), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12424) );
  NOR2_X1 U15539 ( .A1(n12446), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12423) );
  NOR2_X1 U15540 ( .A1(n12424), .A2(n12423), .ZN(n14349) );
  MUX2_X1 U15541 ( .A(n12443), .B(n9638), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n12426) );
  NAND2_X1 U15542 ( .A1(n12361), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12425) );
  NAND2_X1 U15543 ( .A1(n12426), .A2(n12425), .ZN(n14335) );
  MUX2_X1 U15544 ( .A(n12439), .B(n13412), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n12427) );
  INV_X1 U15545 ( .A(n12427), .ZN(n12428) );
  OAI21_X1 U15546 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n12446), .A(
        n12428), .ZN(n14324) );
  OR2_X1 U15547 ( .A1(n12443), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n12431) );
  INV_X1 U15548 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14609) );
  NAND2_X1 U15549 ( .A1(n9638), .A2(n14609), .ZN(n12429) );
  OAI211_X1 U15550 ( .C1(n12361), .C2(P1_EBX_REG_24__SCAN_IN), .A(n12360), .B(
        n12429), .ZN(n12430) );
  AND2_X1 U15551 ( .A1(n12431), .A2(n12430), .ZN(n14314) );
  NAND2_X1 U15552 ( .A1(n12360), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12432) );
  OAI211_X1 U15553 ( .C1(n12361), .C2(P1_EBX_REG_25__SCAN_IN), .A(n9638), .B(
        n12432), .ZN(n12433) );
  OAI21_X1 U15554 ( .B1(n12434), .B2(P1_EBX_REG_25__SCAN_IN), .A(n12433), .ZN(
        n14294) );
  OR2_X1 U15555 ( .A1(n12443), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n12438) );
  INV_X1 U15556 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12435) );
  NAND2_X1 U15557 ( .A1(n9638), .A2(n12435), .ZN(n12436) );
  OAI211_X1 U15558 ( .C1(n12361), .C2(P1_EBX_REG_26__SCAN_IN), .A(n12360), .B(
        n12436), .ZN(n12437) );
  NAND2_X1 U15559 ( .A1(n12438), .A2(n12437), .ZN(n14289) );
  MUX2_X1 U15560 ( .A(n12439), .B(n13412), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12441) );
  NOR2_X1 U15561 ( .A1(n12446), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12440) );
  NOR2_X1 U15562 ( .A1(n12441), .A2(n12440), .ZN(n14269) );
  MUX2_X1 U15563 ( .A(n12443), .B(n9638), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n12445) );
  NAND2_X1 U15564 ( .A1(n12361), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12444) );
  NAND2_X1 U15565 ( .A1(n12445), .A2(n12444), .ZN(n14253) );
  OR2_X1 U15566 ( .A1(n12361), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n12448) );
  OR2_X1 U15567 ( .A1(n12446), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12447) );
  NAND2_X1 U15568 ( .A1(n12448), .A2(n12447), .ZN(n12481) );
  MUX2_X1 U15569 ( .A(n12481), .B(n12448), .S(n13412), .Z(n14248) );
  NAND2_X1 U15570 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20871) );
  AND2_X1 U15571 ( .A1(n20871), .A2(n20874), .ZN(n12451) );
  NOR2_X1 U15572 ( .A1(n12458), .A2(n12451), .ZN(n12452) );
  INV_X1 U15573 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n12453) );
  NAND2_X1 U15574 ( .A1(n12454), .A2(n12453), .ZN(n20875) );
  INV_X1 U15575 ( .A(n20871), .ZN(n13769) );
  OR2_X1 U15576 ( .A1(n20875), .A2(n13769), .ZN(n13553) );
  NAND2_X1 U15577 ( .A1(n13772), .A2(n13553), .ZN(n13300) );
  AND2_X1 U15578 ( .A1(n13300), .A2(n20874), .ZN(n12460) );
  NAND2_X1 U15579 ( .A1(n14416), .A2(n14217), .ZN(n20021) );
  INV_X1 U15580 ( .A(n20021), .ZN(n14377) );
  INV_X1 U15581 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n21017) );
  INV_X1 U15582 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20963) );
  NOR2_X1 U15583 ( .A1(n21017), .A2(n20963), .ZN(n12470) );
  AND2_X1 U15584 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14326) );
  NAND2_X1 U15585 ( .A1(n14326), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14304) );
  NAND3_X1 U15586 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n12466) );
  INV_X1 U15587 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20811) );
  NAND2_X1 U15588 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14406) );
  NOR2_X1 U15589 ( .A1(n20811), .A2(n14406), .ZN(n12465) );
  INV_X1 U15590 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20806) );
  INV_X1 U15591 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20804) );
  INV_X1 U15592 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20802) );
  INV_X1 U15593 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20800) );
  NAND2_X1 U15594 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20023) );
  OR2_X1 U15595 ( .A1(n20800), .A2(n20023), .ZN(n12464) );
  AND4_X1 U15596 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n12463)
         );
  NAND2_X1 U15597 ( .A1(n14217), .A2(n12463), .ZN(n20022) );
  NOR3_X1 U15598 ( .A1(n20806), .A2(n20804), .A3(n19998), .ZN(n14215) );
  NAND3_X1 U15599 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n12465), .A3(n14215), 
        .ZN(n14389) );
  NOR2_X1 U15600 ( .A1(n12466), .A2(n14389), .ZN(n14378) );
  NAND4_X1 U15601 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .A3(P1_REIP_REG_18__SCAN_IN), .A4(n14378), .ZN(n14339) );
  NOR2_X1 U15602 ( .A1(n14304), .A2(n14339), .ZN(n14303) );
  NAND2_X1 U15603 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n12468) );
  INV_X1 U15604 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21010) );
  NOR2_X1 U15605 ( .A1(n12468), .A2(n21010), .ZN(n12455) );
  NAND2_X1 U15606 ( .A1(n14303), .A2(n12455), .ZN(n14274) );
  NAND2_X1 U15607 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n12456) );
  OR2_X1 U15608 ( .A1(n14274), .A2(n12456), .ZN(n12457) );
  NAND2_X1 U15609 ( .A1(n20021), .A2(n12457), .ZN(n14259) );
  OAI21_X1 U15610 ( .B1(n14377), .B2(n12470), .A(n14259), .ZN(n12486) );
  INV_X1 U15611 ( .A(n12458), .ZN(n12459) );
  NOR2_X1 U15612 ( .A1(n12460), .A2(n12459), .ZN(n12461) );
  INV_X1 U15613 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14428) );
  NAND2_X1 U15614 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20016), .ZN(n20008) );
  NAND3_X1 U15615 ( .A1(n15815), .A2(P1_REIP_REG_19__SCAN_IN), .A3(
        P1_REIP_REG_18__SCAN_IN), .ZN(n15809) );
  INV_X1 U15616 ( .A(n15809), .ZN(n12467) );
  INV_X1 U15617 ( .A(n12468), .ZN(n12469) );
  INV_X1 U15618 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20948) );
  INV_X1 U15619 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20835) );
  INV_X1 U15620 ( .A(n12470), .ZN(n12471) );
  NOR2_X1 U15621 ( .A1(n12471), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n12472) );
  AOI22_X1 U15622 ( .A1(n20048), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B1(
        n14250), .B2(n12472), .ZN(n12473) );
  OAI21_X1 U15623 ( .B1(n20054), .B2(n14428), .A(n12473), .ZN(n12474) );
  AOI21_X1 U15624 ( .B1(n12486), .B2(P1_REIP_REG_31__SCAN_IN), .A(n12474), 
        .ZN(n12475) );
  NAND2_X1 U15625 ( .A1(n12478), .A2(n12477), .ZN(P1_U2809) );
  NAND2_X1 U15626 ( .A1(n12480), .A2(n20041), .ZN(n12494) );
  OAI22_X1 U15627 ( .A1(n9718), .A2(n12360), .B1(n12481), .B2(n14255), .ZN(
        n12483) );
  XNOR2_X1 U15628 ( .A(n12483), .B(n12482), .ZN(n14735) );
  AND2_X1 U15629 ( .A1(n13224), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12484) );
  OAI22_X1 U15630 ( .A1(n12485), .A2(n20000), .B1(n20053), .B2(n12583), .ZN(
        n12490) );
  INV_X1 U15631 ( .A(n12486), .ZN(n12488) );
  AOI21_X1 U15632 ( .B1(n14250), .B2(P1_REIP_REG_29__SCAN_IN), .A(
        P1_REIP_REG_30__SCAN_IN), .ZN(n12487) );
  NOR2_X1 U15633 ( .A1(n12488), .A2(n12487), .ZN(n12489) );
  AOI211_X1 U15634 ( .C1(n15848), .C2(P1_EBX_REG_30__SCAN_IN), .A(n12490), .B(
        n12489), .ZN(n12491) );
  OAI21_X1 U15635 ( .B1(n14735), .B2(n20014), .A(n12491), .ZN(n12492) );
  NAND2_X1 U15636 ( .A1(n12494), .A2(n12493), .ZN(P1_U2810) );
  INV_X1 U15637 ( .A(n20167), .ZN(n12495) );
  OR2_X1 U15638 ( .A1(n14241), .A2(n12495), .ZN(n12588) );
  NAND2_X1 U15639 ( .A1(n13305), .A2(n12569), .ZN(n12497) );
  NOR2_X1 U15640 ( .A1(n12497), .A2(n12496), .ZN(n12498) );
  AOI21_X1 U15641 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n10313), .ZN(n14688) );
  NOR2_X1 U15642 ( .A1(n10313), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15873) );
  INV_X1 U15643 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12499) );
  NAND2_X1 U15644 ( .A1(n15883), .A2(n12501), .ZN(n12500) );
  NAND2_X1 U15645 ( .A1(n14809), .A2(n12500), .ZN(n14680) );
  OR2_X1 U15646 ( .A1(n15883), .A2(n12501), .ZN(n12502) );
  NAND2_X1 U15647 ( .A1(n14806), .A2(n12502), .ZN(n14681) );
  NOR2_X1 U15648 ( .A1(n15883), .A2(n14790), .ZN(n12503) );
  NAND2_X1 U15649 ( .A1(n14680), .A2(n14788), .ZN(n12505) );
  AOI22_X1 U15650 ( .A1(n10313), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n14802), .B2(n15883), .ZN(n14791) );
  INV_X1 U15651 ( .A(n14791), .ZN(n12504) );
  AOI21_X1 U15652 ( .B1(n15883), .B2(n14790), .A(n12504), .ZN(n14793) );
  NAND2_X1 U15653 ( .A1(n12513), .A2(n12514), .ZN(n12523) );
  NAND2_X1 U15654 ( .A1(n12523), .A2(n12522), .ZN(n12535) );
  INV_X1 U15655 ( .A(n12534), .ZN(n12506) );
  XNOR2_X1 U15656 ( .A(n12535), .B(n12506), .ZN(n12507) );
  NAND2_X1 U15657 ( .A1(n12507), .A2(n20873), .ZN(n12508) );
  INV_X1 U15658 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20179) );
  XNOR2_X1 U15659 ( .A(n12531), .B(n20179), .ZN(n14155) );
  NAND2_X1 U15660 ( .A1(n20212), .A2(n20227), .ZN(n12524) );
  OAI21_X1 U15661 ( .B1(n13770), .B2(n12513), .A(n12524), .ZN(n12510) );
  INV_X1 U15662 ( .A(n12510), .ZN(n12511) );
  OAI211_X1 U15663 ( .C1(n12514), .C2(n12513), .A(n20873), .B(n12523), .ZN(
        n12516) );
  NOR2_X1 U15664 ( .A1(n12592), .A2(n11606), .ZN(n12515) );
  AND2_X1 U15665 ( .A1(n12516), .A2(n12515), .ZN(n12517) );
  INV_X1 U15666 ( .A(n20162), .ZN(n12519) );
  NAND2_X1 U15667 ( .A1(n12519), .A2(n12518), .ZN(n12520) );
  NAND2_X1 U15668 ( .A1(n12521), .A2(n13305), .ZN(n12528) );
  XNOR2_X1 U15669 ( .A(n12523), .B(n12522), .ZN(n12526) );
  INV_X1 U15670 ( .A(n12524), .ZN(n12525) );
  AOI21_X1 U15671 ( .B1(n12526), .B2(n20873), .A(n12525), .ZN(n12527) );
  NAND2_X1 U15672 ( .A1(n12528), .A2(n12527), .ZN(n13893) );
  NAND2_X1 U15673 ( .A1(n13894), .A2(n13893), .ZN(n13892) );
  NAND2_X1 U15674 ( .A1(n12529), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12530) );
  NAND2_X1 U15675 ( .A1(n13892), .A2(n12530), .ZN(n14154) );
  NAND2_X1 U15676 ( .A1(n14155), .A2(n14154), .ZN(n14153) );
  NAND2_X1 U15677 ( .A1(n12531), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12532) );
  NAND2_X1 U15678 ( .A1(n12533), .A2(n13305), .ZN(n12539) );
  AND2_X1 U15679 ( .A1(n12535), .A2(n12534), .ZN(n12543) );
  INV_X1 U15680 ( .A(n12542), .ZN(n12536) );
  XNOR2_X1 U15681 ( .A(n12543), .B(n12536), .ZN(n12537) );
  NAND2_X1 U15682 ( .A1(n12537), .A2(n20873), .ZN(n12538) );
  NAND2_X1 U15683 ( .A1(n12539), .A2(n12538), .ZN(n12540) );
  INV_X1 U15684 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13915) );
  NAND2_X1 U15685 ( .A1(n12540), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12541) );
  NAND2_X1 U15686 ( .A1(n12543), .A2(n12542), .ZN(n12551) );
  XNOR2_X1 U15687 ( .A(n12550), .B(n12551), .ZN(n12544) );
  NAND2_X1 U15688 ( .A1(n20873), .A2(n12544), .ZN(n12545) );
  OAI21_X1 U15689 ( .B1(n12546), .B2(n9924), .A(n12545), .ZN(n12547) );
  INV_X1 U15690 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16045) );
  XNOR2_X1 U15691 ( .A(n12547), .B(n16045), .ZN(n15903) );
  NAND3_X1 U15692 ( .A1(n12549), .A2(n13305), .A3(n12548), .ZN(n12556) );
  INV_X1 U15693 ( .A(n12550), .ZN(n12552) );
  NOR2_X1 U15694 ( .A1(n12552), .A2(n12551), .ZN(n12561) );
  INV_X1 U15695 ( .A(n12561), .ZN(n12553) );
  XNOR2_X1 U15696 ( .A(n12560), .B(n12553), .ZN(n12554) );
  NAND2_X1 U15697 ( .A1(n20873), .A2(n12554), .ZN(n12555) );
  NAND2_X1 U15698 ( .A1(n12556), .A2(n12555), .ZN(n12557) );
  INV_X1 U15699 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14197) );
  XNOR2_X1 U15700 ( .A(n12557), .B(n14197), .ZN(n15897) );
  NAND2_X1 U15701 ( .A1(n12557), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12558) );
  NAND2_X1 U15702 ( .A1(n12559), .A2(n13305), .ZN(n12564) );
  NAND2_X1 U15703 ( .A1(n12561), .A2(n12560), .ZN(n12567) );
  XNOR2_X1 U15704 ( .A(n12569), .B(n12567), .ZN(n12562) );
  NAND2_X1 U15705 ( .A1(n20873), .A2(n12562), .ZN(n12563) );
  NAND2_X1 U15706 ( .A1(n12564), .A2(n12563), .ZN(n15891) );
  OR2_X1 U15707 ( .A1(n15891), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12565) );
  NAND2_X1 U15708 ( .A1(n15891), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12566) );
  INV_X1 U15709 ( .A(n12567), .ZN(n12568) );
  INV_X1 U15710 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16019) );
  NAND2_X1 U15711 ( .A1(n15883), .A2(n16019), .ZN(n12571) );
  INV_X1 U15712 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14672) );
  INV_X1 U15713 ( .A(n14788), .ZN(n12573) );
  NOR2_X1 U15714 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15875) );
  AND2_X1 U15715 ( .A1(n15875), .A2(n14804), .ZN(n12572) );
  NOR2_X1 U15716 ( .A1(n15883), .A2(n12572), .ZN(n14668) );
  XNOR2_X1 U15717 ( .A(n15883), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14661) );
  NAND2_X1 U15718 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15921) );
  INV_X1 U15719 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15950) );
  INV_X1 U15720 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15936) );
  NAND2_X1 U15721 ( .A1(n15950), .A2(n15936), .ZN(n12574) );
  INV_X1 U15722 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15791) );
  INV_X1 U15723 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14629) );
  INV_X1 U15724 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15910) );
  NAND3_X1 U15725 ( .A1(n14629), .A2(n15910), .A3(n14609), .ZN(n14577) );
  NAND2_X1 U15726 ( .A1(n14608), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12576) );
  NOR2_X1 U15727 ( .A1(n15883), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14566) );
  NAND3_X1 U15728 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14718) );
  NAND2_X1 U15729 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14724) );
  AND2_X1 U15730 ( .A1(n15883), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14565) );
  AOI21_X1 U15731 ( .B1(n9745), .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n13221), .ZN(n14743) );
  NAND2_X1 U15732 ( .A1(n13571), .A2(n20212), .ZN(n12578) );
  NAND2_X1 U15733 ( .A1(n12579), .A2(n12578), .ZN(n13308) );
  OR2_X1 U15734 ( .A1(n13308), .A2(n13319), .ZN(n15741) );
  NAND2_X1 U15735 ( .A1(n12580), .A2(n20719), .ZN(n20870) );
  NAND2_X1 U15736 ( .A1(n20870), .A2(n16055), .ZN(n12581) );
  NOR2_X1 U15737 ( .A1(n20170), .A2(n21017), .ZN(n14740) );
  NAND2_X1 U15738 ( .A1(n16055), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15753) );
  NAND2_X1 U15739 ( .A1(n20874), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12582) );
  AND2_X1 U15740 ( .A1(n15753), .A2(n12582), .ZN(n20164) );
  OR2_X2 U15741 ( .A1(n20152), .A2(n20164), .ZN(n20161) );
  NOR2_X1 U15742 ( .A1(n20161), .A2(n12583), .ZN(n12584) );
  AOI211_X1 U15743 ( .C1(n20152), .C2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14740), .B(n12584), .ZN(n12585) );
  NAND2_X1 U15744 ( .A1(n12588), .A2(n12587), .ZN(P1_U2969) );
  NOR2_X2 U15745 ( .A1(n9641), .A2(n12591), .ZN(n14575) );
  OR2_X1 U15746 ( .A1(n13420), .A2(n13772), .ZN(n12593) );
  NOR2_X1 U15747 ( .A1(n13571), .A2(n12592), .ZN(n13314) );
  NAND2_X1 U15748 ( .A1(n13314), .A2(n11607), .ZN(n13675) );
  NAND2_X1 U15749 ( .A1(n13422), .A2(n20871), .ZN(n12595) );
  OR2_X1 U15750 ( .A1(n12594), .A2(n12595), .ZN(n13560) );
  INV_X1 U15751 ( .A(n13725), .ZN(n14104) );
  NAND2_X1 U15752 ( .A1(n9953), .A2(n13716), .ZN(n12596) );
  AND2_X1 U15753 ( .A1(n13560), .A2(n12596), .ZN(n12597) );
  OAI21_X1 U15754 ( .B1(n13715), .B2(n13554), .A(n12597), .ZN(n12598) );
  NAND2_X1 U15755 ( .A1(n12599), .A2(n13725), .ZN(n13742) );
  NAND2_X2 U15756 ( .A1(n14550), .A2(n13742), .ZN(n14553) );
  NAND2_X1 U15757 ( .A1(n14575), .A2(n12600), .ZN(n12618) );
  OR2_X1 U15758 ( .A1(n14528), .A2(n13298), .ZN(n12615) );
  NOR4_X1 U15759 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12604) );
  NOR4_X1 U15760 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12603) );
  NOR4_X1 U15761 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12602) );
  NOR4_X1 U15762 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12601) );
  AND4_X1 U15763 ( .A1(n12604), .A2(n12603), .A3(n12602), .A4(n12601), .ZN(
        n12609) );
  NOR4_X1 U15764 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12607) );
  NOR4_X1 U15765 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12606) );
  NOR4_X1 U15766 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12605) );
  INV_X1 U15767 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20791) );
  AND4_X1 U15768 ( .A1(n12607), .A2(n12606), .A3(n12605), .A4(n20791), .ZN(
        n12608) );
  NAND2_X1 U15769 ( .A1(n12609), .A2(n12608), .ZN(n12610) );
  AND2_X2 U15770 ( .A1(n12610), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14547)
         );
  INV_X1 U15771 ( .A(n14547), .ZN(n14481) );
  NOR3_X1 U15772 ( .A1(n14528), .A2(n14104), .A3(n11600), .ZN(n14530) );
  INV_X1 U15773 ( .A(DATAI_13_), .ZN(n20953) );
  NAND2_X1 U15774 ( .A1(n14547), .A2(BUF1_REG_13__SCAN_IN), .ZN(n12611) );
  OAI21_X1 U15775 ( .B1(n14547), .B2(n20953), .A(n12611), .ZN(n20140) );
  INV_X1 U15776 ( .A(n20140), .ZN(n14555) );
  INV_X2 U15777 ( .A(n14528), .ZN(n14550) );
  OAI22_X1 U15778 ( .A1(n14540), .A2(n14555), .B1(n14550), .B2(n12612), .ZN(
        n12613) );
  AOI21_X1 U15779 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n14542), .A(n12613), .ZN(
        n12614) );
  INV_X1 U15780 ( .A(n12614), .ZN(n12616) );
  NOR2_X1 U15781 ( .A1(n12616), .A2(n10306), .ZN(n12617) );
  INV_X1 U15782 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15289) );
  OAI21_X1 U15783 ( .B1(n12620), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n12621), .ZN(n15141) );
  INV_X1 U15784 ( .A(n15141), .ZN(n16057) );
  AOI21_X1 U15785 ( .B1(n15149), .B2(n9781), .A(n12620), .ZN(n15153) );
  NAND2_X1 U15786 ( .A1(n12623), .A2(n13243), .ZN(n12624) );
  AND2_X1 U15787 ( .A1(n9781), .A2(n12624), .ZN(n15159) );
  OAI21_X1 U15788 ( .B1(n12625), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n12623), .ZN(n12626) );
  INV_X1 U15789 ( .A(n12626), .ZN(n16071) );
  AOI21_X1 U15790 ( .B1(n12628), .B2(n14863), .A(n12625), .ZN(n15174) );
  OAI21_X1 U15791 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n12629), .A(
        n12628), .ZN(n12630) );
  INV_X1 U15792 ( .A(n12630), .ZN(n16089) );
  AOI21_X1 U15793 ( .B1(n15188), .B2(n12632), .A(n12629), .ZN(n15192) );
  OAI21_X1 U15794 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12633), .A(
        n12632), .ZN(n16112) );
  INV_X1 U15795 ( .A(n16112), .ZN(n13270) );
  AOI21_X1 U15796 ( .B1(n15215), .B2(n12635), .A(n12633), .ZN(n15218) );
  OAI21_X1 U15797 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12636), .A(
        n12635), .ZN(n15229) );
  INV_X1 U15798 ( .A(n15229), .ZN(n14874) );
  AOI21_X1 U15799 ( .B1(n12638), .B2(n15240), .A(n12636), .ZN(n15243) );
  OAI21_X1 U15800 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12639), .A(
        n12638), .ZN(n16124) );
  INV_X1 U15801 ( .A(n16124), .ZN(n14906) );
  AOI21_X1 U15802 ( .B1(n12642), .B2(n12641), .A(n12639), .ZN(n18951) );
  AOI21_X1 U15803 ( .B1(n18960), .B2(n12644), .A(n12645), .ZN(n18963) );
  AOI21_X1 U15804 ( .B1(n16150), .B2(n12660), .A(n12646), .ZN(n18987) );
  AOI21_X1 U15805 ( .B1(n16171), .B2(n9683), .A(n12647), .ZN(n19010) );
  AOI21_X1 U15806 ( .B1(n16191), .B2(n12659), .A(n12649), .ZN(n19023) );
  AOI21_X1 U15807 ( .B1(n15264), .B2(n12651), .A(n12652), .ZN(n19029) );
  AOI21_X1 U15808 ( .B1(n16214), .B2(n12653), .A(n12655), .ZN(n19047) );
  AOI21_X1 U15809 ( .B1(n12656), .B2(n12657), .A(n12658), .ZN(n16215) );
  OAI22_X1 U15810 ( .A1(n9877), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n19072) );
  INV_X1 U15811 ( .A(n19072), .ZN(n14187) );
  AOI22_X1 U15812 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19191), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n9877), .ZN(n14068) );
  NOR2_X1 U15813 ( .A1(n14187), .A2(n14068), .ZN(n14067) );
  OAI21_X1 U15814 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n12657), .ZN(n14041) );
  NAND2_X1 U15815 ( .A1(n14067), .A2(n14041), .ZN(n14080) );
  NOR2_X1 U15816 ( .A1(n16215), .A2(n14080), .ZN(n14052) );
  OAI21_X1 U15817 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12658), .A(
        n12653), .ZN(n19181) );
  NAND2_X1 U15818 ( .A1(n14052), .A2(n19181), .ZN(n19045) );
  NOR2_X1 U15819 ( .A1(n19047), .A2(n19045), .ZN(n13986) );
  OAI21_X1 U15820 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n12655), .A(
        n12651), .ZN(n15272) );
  NAND2_X1 U15821 ( .A1(n13986), .A2(n15272), .ZN(n19028) );
  NOR2_X1 U15822 ( .A1(n19029), .A2(n19028), .ZN(n14111) );
  OAI21_X1 U15823 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n12652), .A(
        n12659), .ZN(n16206) );
  NAND2_X1 U15824 ( .A1(n14111), .A2(n16206), .ZN(n19021) );
  NOR2_X1 U15825 ( .A1(n19023), .A2(n19021), .ZN(n14135) );
  OAI21_X1 U15826 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12649), .A(
        n9683), .ZN(n16185) );
  NAND2_X1 U15827 ( .A1(n14135), .A2(n16185), .ZN(n19008) );
  NOR2_X1 U15828 ( .A1(n19010), .A2(n19008), .ZN(n18992) );
  OAI21_X1 U15829 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n12647), .A(
        n12660), .ZN(n18994) );
  NAND2_X1 U15830 ( .A1(n18992), .A2(n18994), .ZN(n18985) );
  NOR2_X1 U15831 ( .A1(n18987), .A2(n18985), .ZN(n18970) );
  OAI21_X1 U15832 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n12646), .A(
        n12644), .ZN(n18972) );
  NAND2_X1 U15833 ( .A1(n18970), .A2(n18972), .ZN(n18955) );
  NOR2_X1 U15834 ( .A1(n18963), .A2(n18955), .ZN(n14923) );
  OAI21_X1 U15835 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12645), .A(
        n12641), .ZN(n15248) );
  NAND2_X1 U15836 ( .A1(n14923), .A2(n15248), .ZN(n18945) );
  NOR2_X1 U15837 ( .A1(n18951), .A2(n18945), .ZN(n18944) );
  NOR2_X1 U15838 ( .A1(n15243), .A2(n14891), .ZN(n14890) );
  NOR2_X1 U15839 ( .A1(n18993), .A2(n14890), .ZN(n14873) );
  NOR2_X1 U15840 ( .A1(n14874), .A2(n14873), .ZN(n14872) );
  NOR2_X1 U15841 ( .A1(n18993), .A2(n14872), .ZN(n13255) );
  NOR2_X1 U15842 ( .A1(n13270), .A2(n13269), .ZN(n13268) );
  NOR2_X1 U15843 ( .A1(n18993), .A2(n13268), .ZN(n13282) );
  NOR2_X1 U15844 ( .A1(n18993), .A2(n14857), .ZN(n16070) );
  NOR2_X1 U15845 ( .A1(n18993), .A2(n14842), .ZN(n16058) );
  NOR2_X1 U15846 ( .A1(n16057), .A2(n16058), .ZN(n16056) );
  XOR2_X1 U15847 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n12621), .Z(
        n15131) );
  XNOR2_X1 U15848 ( .A(n12661), .B(n15131), .ZN(n12662) );
  NOR3_X1 U15849 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15796) );
  NAND2_X1 U15850 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15796), .ZN(n19822) );
  NAND2_X1 U15851 ( .A1(n12662), .A2(n19049), .ZN(n12903) );
  NAND2_X1 U15852 ( .A1(n14938), .A2(n12664), .ZN(n12665) );
  NAND2_X1 U15853 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19967) );
  INV_X1 U15854 ( .A(n19967), .ZN(n19960) );
  OR2_X1 U15855 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19960), .ZN(n12897) );
  NOR2_X1 U15856 ( .A1(n13617), .A2(n12897), .ZN(n12667) );
  NOR2_X1 U15857 ( .A1(n19262), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12669) );
  INV_X1 U15858 ( .A(n12846), .ZN(n12764) );
  AOI22_X1 U15859 ( .A1(n12764), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12871), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12675) );
  INV_X1 U15860 ( .A(n12671), .ZN(n13454) );
  INV_X1 U15861 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n12673) );
  OR2_X1 U15862 ( .A1(n12877), .A2(n12673), .ZN(n12674) );
  OAI211_X1 U15863 ( .C1(n12676), .C2(n12842), .A(n12675), .B(n12674), .ZN(
        n15561) );
  INV_X1 U15864 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12677) );
  OR2_X1 U15865 ( .A1(n12877), .A2(n12677), .ZN(n12681) );
  AOI22_X1 U15866 ( .A1(n12764), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12871), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12680) );
  OR2_X1 U15867 ( .A1(n12842), .A2(n12678), .ZN(n12679) );
  OR2_X1 U15868 ( .A1(n12682), .A2(n12842), .ZN(n12686) );
  OAI22_X1 U15869 ( .A1(n19262), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n19939), 
        .B2(n19931), .ZN(n12683) );
  INV_X1 U15870 ( .A(n12683), .ZN(n12684) );
  AND2_X1 U15871 ( .A1(n12698), .A2(n12684), .ZN(n12685) );
  INV_X1 U15872 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19173) );
  AOI21_X1 U15873 ( .B1(n19956), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12687) );
  OAI211_X1 U15874 ( .C1(n19173), .C2(n19262), .A(n12688), .B(n12687), .ZN(
        n13458) );
  AOI22_X1 U15875 ( .A1(n12669), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12712), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12690) );
  NAND2_X1 U15876 ( .A1(n12690), .A2(n12689), .ZN(n12695) );
  XNOR2_X1 U15877 ( .A(n13456), .B(n12695), .ZN(n13732) );
  OR2_X1 U15878 ( .A1(n12842), .A2(n12691), .ZN(n12694) );
  NAND3_X1 U15879 ( .A1(n12692), .A2(n19931), .A3(n19262), .ZN(n12693) );
  OAI211_X1 U15880 ( .C1(n19931), .C2(n19929), .A(n12694), .B(n12693), .ZN(
        n13731) );
  NOR2_X1 U15881 ( .A1(n13732), .A2(n13731), .ZN(n12697) );
  NOR2_X1 U15882 ( .A1(n13456), .A2(n12695), .ZN(n12696) );
  NAND2_X1 U15883 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12699) );
  OAI211_X1 U15884 ( .C1(n12842), .C2(n12700), .A(n12699), .B(n12698), .ZN(
        n12701) );
  XNOR2_X1 U15885 ( .A(n12702), .B(n12701), .ZN(n13630) );
  INV_X1 U15886 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19167) );
  INV_X1 U15887 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19841) );
  OAI222_X1 U15888 ( .A1(n12847), .A2(n14009), .B1(n12846), .B2(n19167), .C1(
        n12877), .C2(n19841), .ZN(n13629) );
  NOR2_X1 U15889 ( .A1(n13630), .A2(n13629), .ZN(n13628) );
  NOR2_X1 U15890 ( .A1(n12702), .A2(n12701), .ZN(n12703) );
  INV_X1 U15891 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n12705) );
  AOI22_X1 U15892 ( .A1(n12871), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12704) );
  OAI21_X1 U15893 ( .B1(n12877), .B2(n12705), .A(n12704), .ZN(n12709) );
  NAND2_X1 U15894 ( .A1(n12764), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12706) );
  OAI21_X1 U15895 ( .B1(n12842), .B2(n12707), .A(n12706), .ZN(n12708) );
  INV_X1 U15896 ( .A(n12842), .ZN(n12711) );
  AOI22_X1 U15897 ( .A1(n12764), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12871), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12714) );
  INV_X1 U15898 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19846) );
  NAND2_X1 U15899 ( .A1(n12714), .A2(n12713), .ZN(n13988) );
  INV_X1 U15900 ( .A(n13988), .ZN(n12715) );
  INV_X1 U15901 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19158) );
  INV_X1 U15902 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19848) );
  OAI222_X1 U15903 ( .A1(n16293), .A2(n12847), .B1(n12846), .B2(n19158), .C1(
        n12877), .C2(n19848), .ZN(n16290) );
  AOI22_X1 U15904 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10726), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12722) );
  AOI22_X1 U15905 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13036), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12718) );
  NAND2_X1 U15906 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12717) );
  AND2_X1 U15907 ( .A1(n12718), .A2(n12717), .ZN(n12721) );
  AOI22_X1 U15908 ( .A1(n10720), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10421), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12720) );
  NAND2_X1 U15909 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12719) );
  NAND4_X1 U15910 ( .A1(n12722), .A2(n12721), .A3(n12720), .A4(n12719), .ZN(
        n12729) );
  AOI22_X1 U15911 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10381), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12727) );
  AOI22_X1 U15912 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12726) );
  AOI22_X1 U15913 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12725) );
  AOI22_X1 U15914 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13030), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12724) );
  NAND4_X1 U15915 ( .A1(n12727), .A2(n12726), .A3(n12725), .A4(n12724), .ZN(
        n12728) );
  AOI22_X1 U15916 ( .A1(n12764), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12871), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12730) );
  OAI21_X1 U15917 ( .B1(n12938), .B2(n12842), .A(n12730), .ZN(n12731) );
  AOI21_X1 U15918 ( .B1(n12794), .B2(P2_REIP_REG_8__SCAN_IN), .A(n12731), .ZN(
        n14114) );
  AOI22_X1 U15919 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10720), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12737) );
  AOI22_X1 U15920 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n12716), .ZN(n12736) );
  AOI22_X1 U15921 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n13036), .ZN(n12733) );
  NAND2_X1 U15922 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12732) );
  AND2_X1 U15923 ( .A1(n12733), .A2(n12732), .ZN(n12735) );
  NAND2_X1 U15924 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12734) );
  NAND4_X1 U15925 ( .A1(n12737), .A2(n12736), .A3(n12735), .A4(n12734), .ZN(
        n12743) );
  AOI22_X1 U15926 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10726), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12741) );
  AOI22_X1 U15927 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12740) );
  AOI22_X1 U15928 ( .A1(n10381), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12739) );
  AOI22_X1 U15929 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10383), .B1(
        n13030), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12738) );
  NAND4_X1 U15930 ( .A1(n12741), .A2(n12740), .A3(n12739), .A4(n12738), .ZN(
        n12742) );
  AOI22_X1 U15931 ( .A1(n12764), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12871), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12746) );
  INV_X1 U15932 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n12744) );
  OR2_X1 U15933 ( .A1(n12877), .A2(n12744), .ZN(n12745) );
  OAI211_X1 U15934 ( .C1(n12939), .C2(n12842), .A(n12746), .B(n12745), .ZN(
        n15539) );
  INV_X1 U15935 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n12747) );
  OR2_X1 U15936 ( .A1(n12877), .A2(n12747), .ZN(n12763) );
  AOI22_X1 U15937 ( .A1(n12764), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12871), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12762) );
  AOI22_X1 U15938 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12723), .B1(
        n13029), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12751) );
  AOI22_X1 U15939 ( .A1(n10720), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12750) );
  AOI22_X1 U15940 ( .A1(n10381), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U15941 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10383), .B1(
        n13039), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12748) );
  NAND4_X1 U15942 ( .A1(n12751), .A2(n12750), .A3(n12749), .A4(n12748), .ZN(
        n12759) );
  AOI22_X1 U15943 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10726), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12757) );
  AOI22_X1 U15944 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n13036), .ZN(n12753) );
  NAND2_X1 U15945 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n12752) );
  AND2_X1 U15946 ( .A1(n12753), .A2(n12752), .ZN(n12756) );
  AOI22_X1 U15947 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10421), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12755) );
  NAND2_X1 U15948 ( .A1(n13030), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n12754) );
  NAND4_X1 U15949 ( .A1(n12757), .A2(n12756), .A3(n12755), .A4(n12754), .ZN(
        n12758) );
  INV_X1 U15950 ( .A(n13900), .ZN(n12760) );
  OR2_X1 U15951 ( .A1(n12842), .A2(n12760), .ZN(n12761) );
  AOI22_X1 U15952 ( .A1(n12794), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n12764), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n12779) );
  AOI22_X1 U15953 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10720), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12770) );
  AOI22_X1 U15954 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__3__SCAN_IN), .B2(n12716), .ZN(n12769) );
  AOI22_X1 U15955 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n13036), .ZN(n12766) );
  NAND2_X1 U15956 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n12765) );
  AND2_X1 U15957 ( .A1(n12766), .A2(n12765), .ZN(n12768) );
  NAND2_X1 U15958 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12767) );
  NAND4_X1 U15959 ( .A1(n12770), .A2(n12769), .A3(n12768), .A4(n12767), .ZN(
        n12776) );
  AOI22_X1 U15960 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10726), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12774) );
  AOI22_X1 U15961 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12773) );
  AOI22_X1 U15962 ( .A1(n10381), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12772) );
  AOI22_X1 U15963 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10383), .B1(
        n13030), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12771) );
  NAND4_X1 U15964 ( .A1(n12774), .A2(n12773), .A3(n12772), .A4(n12771), .ZN(
        n12775) );
  NOR2_X1 U15965 ( .A1(n12776), .A2(n12775), .ZN(n14024) );
  OAI22_X1 U15966 ( .A1(n12842), .A2(n14024), .B1(n12847), .B2(n16166), .ZN(
        n12777) );
  INV_X1 U15967 ( .A(n12777), .ZN(n12778) );
  NAND2_X1 U15968 ( .A1(n12779), .A2(n12778), .ZN(n16255) );
  AOI22_X1 U15969 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10726), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12785) );
  AOI22_X1 U15970 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__4__SCAN_IN), .B2(n12716), .ZN(n12784) );
  AOI22_X1 U15971 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n13036), .ZN(n12781) );
  NAND2_X1 U15972 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12780) );
  AND2_X1 U15973 ( .A1(n12781), .A2(n12780), .ZN(n12783) );
  NAND2_X1 U15974 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12782) );
  NAND4_X1 U15975 ( .A1(n12785), .A2(n12784), .A3(n12783), .A4(n12782), .ZN(
        n12791) );
  AOI22_X1 U15976 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10720), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12789) );
  AOI22_X1 U15977 ( .A1(n10381), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12788) );
  AOI22_X1 U15978 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12787) );
  AOI22_X1 U15979 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10383), .B1(
        n13030), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12786) );
  NAND4_X1 U15980 ( .A1(n12789), .A2(n12788), .A3(n12787), .A4(n12786), .ZN(
        n12790) );
  NOR2_X1 U15981 ( .A1(n12791), .A2(n12790), .ZN(n14023) );
  AOI22_X1 U15982 ( .A1(n12669), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12871), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12792) );
  OAI21_X1 U15983 ( .B1(n14023), .B2(n12842), .A(n12792), .ZN(n12793) );
  AOI21_X1 U15984 ( .B1(n12794), .B2(P2_REIP_REG_12__SCAN_IN), .A(n12793), 
        .ZN(n16241) );
  AOI22_X1 U15985 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10720), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12800) );
  AOI22_X1 U15986 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12716), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12799) );
  AOI22_X1 U15987 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13036), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12796) );
  NAND2_X1 U15988 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n12795) );
  AND2_X1 U15989 ( .A1(n12796), .A2(n12795), .ZN(n12798) );
  NAND2_X1 U15990 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12797) );
  NAND4_X1 U15991 ( .A1(n12800), .A2(n12799), .A3(n12798), .A4(n12797), .ZN(
        n12806) );
  AOI22_X1 U15992 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10726), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12804) );
  AOI22_X1 U15993 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12803) );
  AOI22_X1 U15994 ( .A1(n10381), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12802) );
  AOI22_X1 U15995 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13030), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12801) );
  NAND4_X1 U15996 ( .A1(n12804), .A2(n12803), .A3(n12802), .A4(n12801), .ZN(
        n12805) );
  AOI22_X1 U15997 ( .A1(n12669), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12871), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12809) );
  INV_X1 U15998 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n12807) );
  OR2_X1 U15999 ( .A1(n12877), .A2(n12807), .ZN(n12808) );
  OAI211_X1 U16000 ( .C1(n12940), .C2(n12842), .A(n12809), .B(n12808), .ZN(
        n15519) );
  INV_X1 U16001 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n12810) );
  OR2_X1 U16002 ( .A1(n12877), .A2(n12810), .ZN(n12826) );
  AOI22_X1 U16003 ( .A1(n12669), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12871), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12825) );
  AOI22_X1 U16004 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10381), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12814) );
  AOI22_X1 U16005 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10720), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12813) );
  AOI22_X1 U16006 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12812) );
  AOI22_X1 U16007 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10383), .B1(
        n13039), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12811) );
  NAND4_X1 U16008 ( .A1(n12814), .A2(n12813), .A3(n12812), .A4(n12811), .ZN(
        n12822) );
  AOI22_X1 U16009 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n12716), .ZN(n12820) );
  AOI22_X1 U16010 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n13036), .ZN(n12816) );
  NAND2_X1 U16011 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12815) );
  AND2_X1 U16012 ( .A1(n12816), .A2(n12815), .ZN(n12819) );
  AOI22_X1 U16013 ( .A1(n10726), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12818) );
  NAND2_X1 U16014 ( .A1(n13030), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12817) );
  NAND4_X1 U16015 ( .A1(n12820), .A2(n12819), .A3(n12818), .A4(n12817), .ZN(
        n12821) );
  INV_X1 U16016 ( .A(n15042), .ZN(n12823) );
  OR2_X1 U16017 ( .A1(n12842), .A2(n12823), .ZN(n12824) );
  AOI22_X1 U16018 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10720), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12832) );
  AOI22_X1 U16019 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n12716), .ZN(n12831) );
  AOI22_X1 U16020 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n13036), .ZN(n12828) );
  NAND2_X1 U16021 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12827) );
  AND2_X1 U16022 ( .A1(n12828), .A2(n12827), .ZN(n12830) );
  NAND2_X1 U16023 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12829) );
  NAND4_X1 U16024 ( .A1(n12832), .A2(n12831), .A3(n12830), .A4(n12829), .ZN(
        n12838) );
  AOI22_X1 U16025 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10726), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12836) );
  AOI22_X1 U16026 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12835) );
  AOI22_X1 U16027 ( .A1(n10381), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12834) );
  AOI22_X1 U16028 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10383), .B1(
        n13030), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12833) );
  NAND4_X1 U16029 ( .A1(n12836), .A2(n12835), .A3(n12834), .A4(n12833), .ZN(
        n12837) );
  AOI22_X1 U16030 ( .A1(n12669), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12871), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12841) );
  INV_X1 U16031 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n12839) );
  OR2_X1 U16032 ( .A1(n12877), .A2(n12839), .ZN(n12840) );
  OAI211_X1 U16033 ( .C1(n12941), .C2(n12842), .A(n12841), .B(n12840), .ZN(
        n15486) );
  INV_X1 U16034 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n12843) );
  OR2_X1 U16035 ( .A1(n12877), .A2(n12843), .ZN(n12845) );
  AOI22_X1 U16036 ( .A1(n12669), .A2(P2_EAX_REG_16__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n12871), .ZN(n12844) );
  INV_X1 U16037 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19862) );
  INV_X1 U16038 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n15115) );
  OAI222_X1 U16039 ( .A1(n12877), .A2(n19862), .B1(n12847), .B2(n10893), .C1(
        n12846), .C2(n15115), .ZN(n15114) );
  AOI22_X1 U16040 ( .A1(n12669), .A2(P2_EAX_REG_18__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n12871), .ZN(n12849) );
  INV_X1 U16041 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n14914) );
  OR2_X1 U16042 ( .A1(n12877), .A2(n14914), .ZN(n12848) );
  INV_X1 U16043 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19865) );
  OR2_X1 U16044 ( .A1(n12877), .A2(n19865), .ZN(n12851) );
  AOI22_X1 U16045 ( .A1(n12764), .A2(P2_EAX_REG_19__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n12871), .ZN(n12850) );
  AOI22_X1 U16046 ( .A1(n12764), .A2(P2_EAX_REG_20__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n12871), .ZN(n12853) );
  INV_X1 U16047 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19867) );
  OR2_X1 U16048 ( .A1(n12877), .A2(n19867), .ZN(n12852) );
  NAND2_X1 U16049 ( .A1(n12853), .A2(n12852), .ZN(n14881) );
  AOI22_X1 U16050 ( .A1(n12669), .A2(P2_EAX_REG_21__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n12871), .ZN(n12855) );
  INV_X1 U16051 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19869) );
  OR2_X1 U16052 ( .A1(n12877), .A2(n19869), .ZN(n12854) );
  NAND2_X1 U16053 ( .A1(n12855), .A2(n12854), .ZN(n13261) );
  AOI22_X1 U16054 ( .A1(n12669), .A2(P2_EAX_REG_22__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n12871), .ZN(n12858) );
  INV_X1 U16055 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n12856) );
  OR2_X1 U16056 ( .A1(n12877), .A2(n12856), .ZN(n12857) );
  NAND2_X1 U16057 ( .A1(n12858), .A2(n12857), .ZN(n13287) );
  AOI22_X1 U16058 ( .A1(n12669), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12871), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12860) );
  INV_X1 U16059 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19872) );
  OR2_X1 U16060 ( .A1(n12877), .A2(n19872), .ZN(n12859) );
  NAND2_X1 U16061 ( .A1(n12860), .A2(n12859), .ZN(n13290) );
  INV_X1 U16062 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19874) );
  OR2_X1 U16063 ( .A1(n12877), .A2(n19874), .ZN(n12863) );
  AOI22_X1 U16064 ( .A1(n12764), .A2(P2_EAX_REG_24__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n12871), .ZN(n12862) );
  AND2_X1 U16065 ( .A1(n12863), .A2(n12862), .ZN(n15081) );
  AOI22_X1 U16066 ( .A1(n12764), .A2(P2_EAX_REG_25__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n12871), .ZN(n12865) );
  INV_X1 U16067 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19876) );
  OR2_X1 U16068 ( .A1(n12877), .A2(n19876), .ZN(n12864) );
  NAND2_X1 U16069 ( .A1(n12865), .A2(n12864), .ZN(n14860) );
  INV_X1 U16070 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n16073) );
  OR2_X1 U16071 ( .A1(n12877), .A2(n16073), .ZN(n12867) );
  AOI22_X1 U16072 ( .A1(n12764), .A2(P2_EAX_REG_26__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n12871), .ZN(n12866) );
  AND2_X1 U16073 ( .A1(n12867), .A2(n12866), .ZN(n15071) );
  INV_X1 U16074 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19880) );
  OR2_X1 U16075 ( .A1(n12877), .A2(n19880), .ZN(n12869) );
  AOI22_X1 U16076 ( .A1(n12764), .A2(P2_EAX_REG_27__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n12871), .ZN(n12868) );
  AND2_X1 U16077 ( .A1(n12869), .A2(n12868), .ZN(n13248) );
  INV_X1 U16078 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n12870) );
  OR2_X1 U16079 ( .A1(n12877), .A2(n12870), .ZN(n12873) );
  AOI22_X1 U16080 ( .A1(n12764), .A2(P2_EAX_REG_28__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n12871), .ZN(n12872) );
  AND2_X1 U16081 ( .A1(n12873), .A2(n12872), .ZN(n14848) );
  AOI22_X1 U16082 ( .A1(n12764), .A2(P2_EAX_REG_29__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n12871), .ZN(n12875) );
  INV_X1 U16083 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19882) );
  OR2_X1 U16084 ( .A1(n12877), .A2(n19882), .ZN(n12874) );
  NAND2_X1 U16085 ( .A1(n12875), .A2(n12874), .ZN(n15047) );
  INV_X1 U16086 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n12876) );
  OR2_X1 U16087 ( .A1(n12877), .A2(n12876), .ZN(n12879) );
  AOI22_X1 U16088 ( .A1(n12764), .A2(P2_EAX_REG_30__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n12871), .ZN(n12878) );
  AND2_X1 U16089 ( .A1(n12879), .A2(n12878), .ZN(n12880) );
  NAND2_X1 U16090 ( .A1(n9730), .A2(n12880), .ZN(n12881) );
  NAND2_X1 U16091 ( .A1(n19827), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19971) );
  INV_X2 U16092 ( .A(n19971), .ZN(n19974) );
  OR2_X1 U16093 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19833) );
  NAND3_X1 U16094 ( .A1(n19827), .A2(n19884), .A3(n19833), .ZN(n19830) );
  NOR2_X1 U16095 ( .A1(n19960), .A2(n19830), .ZN(n13587) );
  INV_X1 U16096 ( .A(n13587), .ZN(n13378) );
  NOR2_X1 U16097 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n13378), .ZN(n12888) );
  AND2_X1 U16098 ( .A1(n12882), .A2(n12888), .ZN(n16361) );
  NAND2_X1 U16099 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19959), .ZN(n19269) );
  NOR2_X1 U16100 ( .A1(n12883), .A2(n19269), .ZN(n16359) );
  NAND2_X1 U16101 ( .A1(n19033), .A2(n19822), .ZN(n12884) );
  OR2_X1 U16102 ( .A1(n16359), .A2(n12884), .ZN(n12885) );
  AOI22_X1 U16103 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n18996), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19054), .ZN(n12894) );
  INV_X1 U16104 ( .A(n12886), .ZN(n12887) );
  INV_X1 U16105 ( .A(n12888), .ZN(n12889) );
  NAND2_X1 U16106 ( .A1(n13532), .A2(n12889), .ZN(n14836) );
  INV_X1 U16107 ( .A(n13355), .ZN(n13354) );
  NAND2_X1 U16108 ( .A1(n12890), .A2(n12897), .ZN(n12891) );
  OR2_X1 U16109 ( .A1(n13354), .A2(n12891), .ZN(n12892) );
  NAND2_X1 U16110 ( .A1(n14836), .A2(n12892), .ZN(n19055) );
  NAND2_X1 U16111 ( .A1(n19055), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12893) );
  OAI211_X1 U16112 ( .C1(n15300), .C2(n19053), .A(n12894), .B(n12893), .ZN(
        n12895) );
  AOI21_X1 U16113 ( .B1(n15301), .B2(n19062), .A(n12895), .ZN(n12901) );
  NAND2_X1 U16114 ( .A1(n12897), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12898) );
  NOR2_X1 U16115 ( .A1(n13617), .A2(n12898), .ZN(n12899) );
  NAND2_X1 U16116 ( .A1(n10946), .A2(n19031), .ZN(n12900) );
  NAND2_X1 U16117 ( .A1(n12903), .A2(n12902), .ZN(P2_U2825) );
  NAND2_X1 U16118 ( .A1(n12904), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12905) );
  NAND2_X1 U16119 ( .A1(n12928), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12909) );
  NOR2_X1 U16120 ( .A1(n19922), .A2(n19929), .ZN(n19713) );
  NAND2_X1 U16121 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19713), .ZN(
        n12918) );
  INV_X1 U16122 ( .A(n12918), .ZN(n12907) );
  INV_X1 U16123 ( .A(n19804), .ZN(n12906) );
  OAI211_X1 U16124 ( .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n12907), .A(
        n12906), .B(n19902), .ZN(n12908) );
  INV_X1 U16125 ( .A(n12916), .ZN(n12936) );
  INV_X1 U16126 ( .A(n12915), .ZN(n12914) );
  NAND2_X1 U16127 ( .A1(n12936), .A2(n12914), .ZN(n13749) );
  NAND2_X1 U16128 ( .A1(n12916), .A2(n12915), .ZN(n12917) );
  NAND2_X1 U16129 ( .A1(n10688), .A2(n12931), .ZN(n12922) );
  INV_X1 U16130 ( .A(n19902), .ZN(n19906) );
  NAND2_X1 U16131 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19581) );
  NAND2_X1 U16132 ( .A1(n19581), .A2(n19922), .ZN(n12919) );
  NAND2_X1 U16133 ( .A1(n12919), .A2(n12918), .ZN(n19358) );
  NOR2_X1 U16134 ( .A1(n19906), .A2(n19358), .ZN(n12920) );
  AOI21_X1 U16135 ( .B1(n12928), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12920), .ZN(n12921) );
  AOI22_X1 U16136 ( .A1(n12928), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19902), .B2(n19939), .ZN(n12924) );
  NAND2_X1 U16137 ( .A1(n12928), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12929) );
  XNOR2_X1 U16138 ( .A(n19929), .B(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19357) );
  NAND2_X1 U16139 ( .A1(n19357), .A2(n19902), .ZN(n19551) );
  NAND2_X1 U16140 ( .A1(n12929), .A2(n19551), .ZN(n12930) );
  NAND2_X1 U16141 ( .A1(n13409), .A2(n12932), .ZN(n12933) );
  NAND2_X1 U16142 ( .A1(n13706), .A2(n13705), .ZN(n13704) );
  NAND2_X1 U16143 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n12904), .ZN(
        n12935) );
  AND2_X1 U16144 ( .A1(n12936), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12937) );
  NAND2_X1 U16145 ( .A1(n14164), .A2(n15042), .ZN(n15025) );
  AOI22_X1 U16146 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10720), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12947) );
  AOI22_X1 U16147 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__3__SCAN_IN), .B2(n12716), .ZN(n12946) );
  AOI22_X1 U16148 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n13036), .ZN(n12943) );
  NAND2_X1 U16149 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n12942) );
  AND2_X1 U16150 ( .A1(n12943), .A2(n12942), .ZN(n12945) );
  NAND2_X1 U16151 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12944) );
  NAND4_X1 U16152 ( .A1(n12947), .A2(n12946), .A3(n12945), .A4(n12944), .ZN(
        n12953) );
  AOI22_X1 U16153 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10726), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12951) );
  AOI22_X1 U16154 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12950) );
  AOI22_X1 U16155 ( .A1(n10381), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12949) );
  AOI22_X1 U16156 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10383), .B1(
        n13030), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12948) );
  NAND4_X1 U16157 ( .A1(n12951), .A2(n12950), .A3(n12949), .A4(n12948), .ZN(
        n12952) );
  OR2_X1 U16158 ( .A1(n12953), .A2(n12952), .ZN(n15001) );
  AOI22_X1 U16159 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10720), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12959) );
  AOI22_X1 U16160 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__2__SCAN_IN), .B2(n12716), .ZN(n12958) );
  AOI22_X1 U16161 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n13036), .ZN(n12955) );
  NAND2_X1 U16162 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12954) );
  AND2_X1 U16163 ( .A1(n12955), .A2(n12954), .ZN(n12957) );
  NAND2_X1 U16164 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12956) );
  NAND4_X1 U16165 ( .A1(n12959), .A2(n12958), .A3(n12957), .A4(n12956), .ZN(
        n12965) );
  AOI22_X1 U16166 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10726), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12963) );
  AOI22_X1 U16167 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12962) );
  AOI22_X1 U16168 ( .A1(n10381), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12961) );
  AOI22_X1 U16169 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10383), .B1(
        n13030), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12960) );
  NAND4_X1 U16170 ( .A1(n12963), .A2(n12962), .A3(n12961), .A4(n12960), .ZN(
        n12964) );
  NOR2_X1 U16171 ( .A1(n12965), .A2(n12964), .ZN(n15007) );
  AOI22_X1 U16172 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10720), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12971) );
  AOI22_X1 U16173 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n12716), .ZN(n12970) );
  AOI22_X1 U16174 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n13036), .ZN(n12967) );
  NAND2_X1 U16175 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12966) );
  AND2_X1 U16176 ( .A1(n12967), .A2(n12966), .ZN(n12969) );
  NAND2_X1 U16177 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12968) );
  NAND4_X1 U16178 ( .A1(n12971), .A2(n12970), .A3(n12969), .A4(n12968), .ZN(
        n12977) );
  AOI22_X1 U16179 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10726), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12975) );
  AOI22_X1 U16180 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12974) );
  AOI22_X1 U16181 ( .A1(n10381), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12973) );
  AOI22_X1 U16182 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10383), .B1(
        n13030), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12972) );
  NAND4_X1 U16183 ( .A1(n12975), .A2(n12974), .A3(n12973), .A4(n12972), .ZN(
        n12976) );
  OR2_X1 U16184 ( .A1(n12977), .A2(n12976), .ZN(n15011) );
  INV_X1 U16185 ( .A(n15011), .ZN(n12990) );
  AOI22_X1 U16186 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10720), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12983) );
  AOI22_X1 U16187 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12716), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12982) );
  AOI22_X1 U16188 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13036), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12979) );
  NAND2_X1 U16189 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12978) );
  AND2_X1 U16190 ( .A1(n12979), .A2(n12978), .ZN(n12981) );
  NAND2_X1 U16191 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12980) );
  NAND4_X1 U16192 ( .A1(n12983), .A2(n12982), .A3(n12981), .A4(n12980), .ZN(
        n12989) );
  AOI22_X1 U16193 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10726), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12987) );
  AOI22_X1 U16194 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12986) );
  AOI22_X1 U16195 ( .A1(n10381), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12985) );
  AOI22_X1 U16196 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13030), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12984) );
  NAND4_X1 U16197 ( .A1(n12987), .A2(n12986), .A3(n12985), .A4(n12984), .ZN(
        n12988) );
  NOR2_X1 U16198 ( .A1(n12989), .A2(n12988), .ZN(n15020) );
  OR2_X1 U16199 ( .A1(n12990), .A2(n15020), .ZN(n15005) );
  NOR2_X1 U16200 ( .A1(n15007), .A2(n15005), .ZN(n15000) );
  AND2_X1 U16201 ( .A1(n15001), .A2(n15000), .ZN(n12991) );
  AOI22_X1 U16202 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10720), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12997) );
  AOI22_X1 U16203 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__4__SCAN_IN), .B2(n12716), .ZN(n12996) );
  AOI22_X1 U16204 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n13036), .ZN(n12993) );
  NAND2_X1 U16205 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12992) );
  AND2_X1 U16206 ( .A1(n12993), .A2(n12992), .ZN(n12995) );
  NAND2_X1 U16207 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12994) );
  NAND4_X1 U16208 ( .A1(n12997), .A2(n12996), .A3(n12995), .A4(n12994), .ZN(
        n13003) );
  AOI22_X1 U16209 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10726), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13001) );
  AOI22_X1 U16210 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13000) );
  AOI22_X1 U16211 ( .A1(n10381), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12999) );
  AOI22_X1 U16212 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10383), .B1(
        n13030), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12998) );
  NAND4_X1 U16213 ( .A1(n13001), .A2(n13000), .A3(n12999), .A4(n12998), .ZN(
        n13002) );
  NOR2_X1 U16214 ( .A1(n13003), .A2(n13002), .ZN(n14996) );
  INV_X1 U16215 ( .A(n14996), .ZN(n13004) );
  AOI22_X1 U16216 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10726), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13008) );
  AOI22_X1 U16217 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13007) );
  AOI22_X1 U16218 ( .A1(n10381), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13006) );
  AOI22_X1 U16219 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13030), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13005) );
  NAND4_X1 U16220 ( .A1(n13008), .A2(n13007), .A3(n13006), .A4(n13005), .ZN(
        n13016) );
  AOI22_X1 U16221 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10720), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13014) );
  AOI22_X1 U16222 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12716), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13013) );
  AOI22_X1 U16223 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13036), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13010) );
  NAND2_X1 U16224 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n13009) );
  AND2_X1 U16225 ( .A1(n13010), .A2(n13009), .ZN(n13012) );
  NAND2_X1 U16226 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n13011) );
  NAND4_X1 U16227 ( .A1(n13014), .A2(n13013), .A3(n13012), .A4(n13011), .ZN(
        n13015) );
  NOR2_X1 U16228 ( .A1(n13016), .A2(n13015), .ZN(n14991) );
  AOI22_X1 U16229 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10720), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13022) );
  AOI22_X1 U16230 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__6__SCAN_IN), .B2(n12716), .ZN(n13021) );
  AOI22_X1 U16231 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n13036), .ZN(n13018) );
  NAND2_X1 U16232 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n13017) );
  AND2_X1 U16233 ( .A1(n13018), .A2(n13017), .ZN(n13020) );
  NAND2_X1 U16234 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n13019) );
  NAND4_X1 U16235 ( .A1(n13022), .A2(n13021), .A3(n13020), .A4(n13019), .ZN(
        n13028) );
  AOI22_X1 U16236 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10726), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13026) );
  AOI22_X1 U16237 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13025) );
  AOI22_X1 U16238 ( .A1(n10381), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13024) );
  AOI22_X1 U16239 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10383), .B1(
        n13030), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13023) );
  NAND4_X1 U16240 ( .A1(n13026), .A2(n13025), .A3(n13024), .A4(n13023), .ZN(
        n13027) );
  OR2_X1 U16241 ( .A1(n13028), .A2(n13027), .ZN(n14986) );
  AOI22_X1 U16242 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10381), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13034) );
  AOI22_X1 U16243 ( .A1(n13029), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10720), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13033) );
  AOI22_X1 U16244 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10721), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13032) );
  AOI22_X1 U16245 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10383), .B1(
        n13030), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13031) );
  NAND4_X1 U16246 ( .A1(n13034), .A2(n13033), .A3(n13032), .A4(n13031), .ZN(
        n13045) );
  AOI22_X1 U16247 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13043) );
  AOI22_X1 U16248 ( .A1(n10319), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n13036), .ZN(n13038) );
  NAND2_X1 U16249 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n13037) );
  AND2_X1 U16250 ( .A1(n13038), .A2(n13037), .ZN(n13042) );
  AOI22_X1 U16251 ( .A1(n10726), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10421), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13041) );
  NAND2_X1 U16252 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n13040) );
  NAND4_X1 U16253 ( .A1(n13043), .A2(n13042), .A3(n13041), .A4(n13040), .ZN(
        n13044) );
  NOR2_X1 U16254 ( .A1(n13045), .A2(n13044), .ZN(n13081) );
  AOI22_X1 U16255 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9650), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13055) );
  AOI22_X1 U16256 ( .A1(n13187), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13116), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13054) );
  AOI22_X1 U16257 ( .A1(n10330), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13053) );
  INV_X1 U16258 ( .A(n13048), .ZN(n15598) );
  NAND2_X1 U16259 ( .A1(n15598), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n13051) );
  NAND2_X1 U16260 ( .A1(n9653), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13050) );
  OAI21_X1 U16261 ( .B1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n13049), .ZN(n13195) );
  AND3_X1 U16262 ( .A1(n13051), .A2(n13050), .A3(n13195), .ZN(n13052) );
  NAND4_X1 U16263 ( .A1(n13055), .A2(n13054), .A3(n13053), .A4(n13052), .ZN(
        n13063) );
  AOI22_X1 U16264 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9650), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13061) );
  AOI22_X1 U16265 ( .A1(n13187), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13116), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13060) );
  AOI22_X1 U16266 ( .A1(n10330), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9657), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13059) );
  NAND2_X1 U16267 ( .A1(n15598), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13057) );
  NAND2_X1 U16268 ( .A1(n9645), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13056) );
  INV_X1 U16269 ( .A(n13195), .ZN(n13174) );
  AND3_X1 U16270 ( .A1(n13057), .A2(n13056), .A3(n13174), .ZN(n13058) );
  NAND4_X1 U16271 ( .A1(n13061), .A2(n13060), .A3(n13059), .A4(n13058), .ZN(
        n13062) );
  NAND2_X1 U16272 ( .A1(n13063), .A2(n13062), .ZN(n13086) );
  NOR2_X1 U16273 ( .A1(n13380), .A2(n13086), .ZN(n13064) );
  XOR2_X1 U16274 ( .A(n13081), .B(n13064), .Z(n13087) );
  XNOR2_X1 U16275 ( .A(n14985), .B(n13087), .ZN(n14977) );
  INV_X1 U16276 ( .A(n13086), .ZN(n13082) );
  NAND2_X1 U16277 ( .A1(n13380), .A2(n13082), .ZN(n14979) );
  AOI22_X1 U16278 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9650), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13072) );
  AOI22_X1 U16279 ( .A1(n13187), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13116), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13071) );
  AOI22_X1 U16280 ( .A1(n10330), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13070) );
  NAND2_X1 U16281 ( .A1(n15598), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n13068) );
  NAND2_X1 U16282 ( .A1(n9645), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n13067) );
  AND3_X1 U16283 ( .A1(n13068), .A2(n13067), .A3(n13195), .ZN(n13069) );
  NAND4_X1 U16284 ( .A1(n13072), .A2(n13071), .A3(n13070), .A4(n13069), .ZN(
        n13080) );
  AOI22_X1 U16285 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9650), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13078) );
  AOI22_X1 U16286 ( .A1(n13187), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13116), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13077) );
  AOI22_X1 U16287 ( .A1(n10330), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9657), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13076) );
  NAND2_X1 U16288 ( .A1(n15598), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13074) );
  NAND2_X1 U16289 ( .A1(n9651), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13073) );
  AND3_X1 U16290 ( .A1(n13074), .A2(n13073), .A3(n13174), .ZN(n13075) );
  NAND4_X1 U16291 ( .A1(n13078), .A2(n13077), .A3(n13076), .A4(n13075), .ZN(
        n13079) );
  NAND2_X1 U16292 ( .A1(n13080), .A2(n13079), .ZN(n13088) );
  INV_X1 U16293 ( .A(n13081), .ZN(n13083) );
  NAND2_X1 U16294 ( .A1(n13083), .A2(n13082), .ZN(n13089) );
  XOR2_X1 U16295 ( .A(n13088), .B(n13089), .Z(n13084) );
  NAND2_X1 U16296 ( .A1(n13084), .A2(n13147), .ZN(n14968) );
  INV_X1 U16297 ( .A(n13088), .ZN(n13085) );
  NAND2_X1 U16298 ( .A1(n13380), .A2(n13085), .ZN(n14970) );
  NOR2_X1 U16299 ( .A1(n13089), .A2(n13088), .ZN(n13104) );
  AOI22_X1 U16300 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9650), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13095) );
  AOI22_X1 U16301 ( .A1(n13187), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13116), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13094) );
  AOI22_X1 U16302 ( .A1(n10330), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9657), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13093) );
  NAND2_X1 U16303 ( .A1(n15598), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n13091) );
  NAND2_X1 U16304 ( .A1(n9645), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n13090) );
  AND3_X1 U16305 ( .A1(n13091), .A2(n13090), .A3(n13195), .ZN(n13092) );
  NAND4_X1 U16306 ( .A1(n13095), .A2(n13094), .A3(n13093), .A4(n13092), .ZN(
        n13103) );
  AOI22_X1 U16307 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9650), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13101) );
  AOI22_X1 U16308 ( .A1(n13187), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13116), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13100) );
  AOI22_X1 U16309 ( .A1(n10330), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9657), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13099) );
  NAND2_X1 U16310 ( .A1(n15598), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13097) );
  NAND2_X1 U16311 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n13096) );
  AND3_X1 U16312 ( .A1(n13097), .A2(n13096), .A3(n13174), .ZN(n13098) );
  NAND4_X1 U16313 ( .A1(n13101), .A2(n13100), .A3(n13099), .A4(n13098), .ZN(
        n13102) );
  AND2_X1 U16314 ( .A1(n13103), .A2(n13102), .ZN(n13106) );
  NAND2_X1 U16315 ( .A1(n13104), .A2(n13106), .ZN(n13144) );
  OAI211_X1 U16316 ( .C1(n13104), .C2(n13106), .A(n13147), .B(n13144), .ZN(
        n13108) );
  XNOR2_X1 U16317 ( .A(n9691), .B(n13105), .ZN(n14964) );
  INV_X1 U16318 ( .A(n13106), .ZN(n13107) );
  NOR2_X1 U16319 ( .A1(n19956), .A2(n13107), .ZN(n14963) );
  NAND2_X1 U16320 ( .A1(n14964), .A2(n14963), .ZN(n14962) );
  OR2_X1 U16321 ( .A1(n9691), .A2(n13108), .ZN(n13109) );
  NAND2_X1 U16322 ( .A1(n14962), .A2(n13109), .ZN(n13126) );
  AOI22_X1 U16323 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9650), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13115) );
  AOI22_X1 U16324 ( .A1(n13187), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13116), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13114) );
  AOI22_X1 U16325 ( .A1(n10330), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13113) );
  NAND2_X1 U16326 ( .A1(n15598), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n13111) );
  NAND2_X1 U16327 ( .A1(n9651), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n13110) );
  AND3_X1 U16328 ( .A1(n13111), .A2(n13110), .A3(n13195), .ZN(n13112) );
  NAND4_X1 U16329 ( .A1(n13115), .A2(n13114), .A3(n13113), .A4(n13112), .ZN(
        n13124) );
  AOI22_X1 U16330 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9650), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13122) );
  AOI22_X1 U16331 ( .A1(n13187), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13116), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13121) );
  AOI22_X1 U16332 ( .A1(n10330), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13120) );
  NAND2_X1 U16333 ( .A1(n15598), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n13118) );
  NAND2_X1 U16334 ( .A1(n9653), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n13117) );
  AND3_X1 U16335 ( .A1(n13118), .A2(n13117), .A3(n13174), .ZN(n13119) );
  NAND4_X1 U16336 ( .A1(n13122), .A2(n13121), .A3(n13120), .A4(n13119), .ZN(
        n13123) );
  AND2_X1 U16337 ( .A1(n13124), .A2(n13123), .ZN(n13142) );
  XNOR2_X1 U16338 ( .A(n13144), .B(n13142), .ZN(n13125) );
  XNOR2_X1 U16339 ( .A(n13126), .B(n10307), .ZN(n14959) );
  NAND2_X1 U16340 ( .A1(n13380), .A2(n13142), .ZN(n14958) );
  NOR2_X1 U16341 ( .A1(n14959), .A2(n14958), .ZN(n14957) );
  AOI22_X1 U16342 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9650), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13133) );
  AOI22_X1 U16343 ( .A1(n13187), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13116), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13132) );
  AOI22_X1 U16344 ( .A1(n10330), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9657), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13131) );
  NAND2_X1 U16345 ( .A1(n15598), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n13129) );
  NAND2_X1 U16346 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n13128) );
  AND3_X1 U16347 ( .A1(n13129), .A2(n13128), .A3(n13195), .ZN(n13130) );
  NAND4_X1 U16348 ( .A1(n13133), .A2(n13132), .A3(n13131), .A4(n13130), .ZN(
        n13141) );
  AOI22_X1 U16349 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9650), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13139) );
  AOI22_X1 U16350 ( .A1(n13187), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13116), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13138) );
  AOI22_X1 U16351 ( .A1(n10330), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9657), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13137) );
  NAND2_X1 U16352 ( .A1(n15598), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n13135) );
  NAND2_X1 U16353 ( .A1(n9645), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n13134) );
  AND3_X1 U16354 ( .A1(n13135), .A2(n13134), .A3(n13174), .ZN(n13136) );
  NAND4_X1 U16355 ( .A1(n13139), .A2(n13138), .A3(n13137), .A4(n13136), .ZN(
        n13140) );
  NAND2_X1 U16356 ( .A1(n13141), .A2(n13140), .ZN(n13145) );
  INV_X1 U16357 ( .A(n13145), .ZN(n13151) );
  INV_X1 U16358 ( .A(n13142), .ZN(n13143) );
  OR2_X1 U16359 ( .A1(n13144), .A2(n13143), .ZN(n13146) );
  INV_X1 U16360 ( .A(n13146), .ZN(n13148) );
  OR2_X1 U16361 ( .A1(n13146), .A2(n13145), .ZN(n14944) );
  OAI211_X1 U16362 ( .C1(n13151), .C2(n13148), .A(n14944), .B(n13147), .ZN(
        n13149) );
  NOR2_X1 U16363 ( .A1(n13150), .A2(n13149), .ZN(n13166) );
  NAND2_X1 U16364 ( .A1(n13380), .A2(n13151), .ZN(n14950) );
  AOI22_X1 U16365 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9650), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13157) );
  AOI22_X1 U16366 ( .A1(n13187), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13116), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13156) );
  AOI22_X1 U16367 ( .A1(n10330), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13155) );
  NAND2_X1 U16368 ( .A1(n15598), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n13153) );
  NAND2_X1 U16369 ( .A1(n9653), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n13152) );
  AND3_X1 U16370 ( .A1(n13153), .A2(n13152), .A3(n13195), .ZN(n13154) );
  NAND4_X1 U16371 ( .A1(n13157), .A2(n13156), .A3(n13155), .A4(n13154), .ZN(
        n13165) );
  AOI22_X1 U16372 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9650), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13163) );
  AOI22_X1 U16373 ( .A1(n13187), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13116), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13162) );
  AOI22_X1 U16374 ( .A1(n10330), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13161) );
  NAND2_X1 U16375 ( .A1(n15598), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n13159) );
  NAND2_X1 U16376 ( .A1(n9645), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n13158) );
  AND3_X1 U16377 ( .A1(n13159), .A2(n13158), .A3(n13174), .ZN(n13160) );
  NAND4_X1 U16378 ( .A1(n13163), .A2(n13162), .A3(n13161), .A4(n13160), .ZN(
        n13164) );
  AND2_X1 U16379 ( .A1(n13165), .A2(n13164), .ZN(n14945) );
  NAND2_X1 U16380 ( .A1(n19956), .A2(n14945), .ZN(n13167) );
  NOR2_X1 U16381 ( .A1(n14944), .A2(n13167), .ZN(n13184) );
  AOI22_X1 U16382 ( .A1(n9650), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13116), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13173) );
  AOI22_X1 U16383 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13187), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13172) );
  AOI22_X1 U16384 ( .A1(n10330), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13171) );
  NAND2_X1 U16385 ( .A1(n15598), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n13169) );
  NAND2_X1 U16386 ( .A1(n9645), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n13168) );
  AND3_X1 U16387 ( .A1(n13169), .A2(n13168), .A3(n13195), .ZN(n13170) );
  NAND4_X1 U16388 ( .A1(n13173), .A2(n13172), .A3(n13171), .A4(n13170), .ZN(
        n13182) );
  AOI22_X1 U16389 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13116), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13180) );
  AOI22_X1 U16390 ( .A1(n9650), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9657), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13179) );
  INV_X1 U16391 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n19509) );
  AOI22_X1 U16392 ( .A1(n13187), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10330), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13178) );
  NAND2_X1 U16393 ( .A1(n15598), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n13176) );
  NAND2_X1 U16394 ( .A1(n9651), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n13175) );
  AND3_X1 U16395 ( .A1(n13176), .A2(n13175), .A3(n13174), .ZN(n13177) );
  NAND4_X1 U16396 ( .A1(n13180), .A2(n13179), .A3(n13178), .A4(n13177), .ZN(
        n13181) );
  AND2_X1 U16397 ( .A1(n13182), .A2(n13181), .ZN(n13183) );
  NAND2_X1 U16398 ( .A1(n13184), .A2(n13183), .ZN(n13185) );
  OAI21_X1 U16399 ( .B1(n13184), .B2(n13183), .A(n13185), .ZN(n14940) );
  NOR2_X1 U16400 ( .A1(n14941), .A2(n14940), .ZN(n14939) );
  INV_X1 U16401 ( .A(n13185), .ZN(n13186) );
  NOR2_X1 U16402 ( .A1(n14939), .A2(n13186), .ZN(n13204) );
  AOI22_X1 U16403 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13116), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13189) );
  AOI22_X1 U16404 ( .A1(n9650), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13187), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13188) );
  NAND2_X1 U16405 ( .A1(n13189), .A2(n13188), .ZN(n13202) );
  INV_X1 U16406 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13192) );
  AOI22_X1 U16407 ( .A1(n10330), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9657), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13191) );
  AOI21_X1 U16408 ( .B1(n9652), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n13195), .ZN(n13190) );
  OAI211_X1 U16409 ( .C1(n13048), .C2(n13192), .A(n13191), .B(n13190), .ZN(
        n13201) );
  AOI22_X1 U16410 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13187), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13194) );
  AOI22_X1 U16411 ( .A1(n9650), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n9657), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13193) );
  NAND2_X1 U16412 ( .A1(n13194), .A2(n13193), .ZN(n13200) );
  AOI22_X1 U16413 ( .A1(n13116), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n15598), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13198) );
  NAND2_X1 U16414 ( .A1(n9645), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n13197) );
  NAND2_X1 U16415 ( .A1(n10330), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n13196) );
  NAND4_X1 U16416 ( .A1(n13198), .A2(n13197), .A3(n13196), .A4(n13195), .ZN(
        n13199) );
  OAI22_X1 U16417 ( .A1(n13202), .A2(n13201), .B1(n13200), .B2(n13199), .ZN(
        n13203) );
  XNOR2_X1 U16418 ( .A(n13204), .B(n13203), .ZN(n14247) );
  INV_X1 U16419 ( .A(n14178), .ZN(n13205) );
  AND2_X1 U16420 ( .A1(n13206), .A2(n13205), .ZN(n15586) );
  NAND2_X1 U16421 ( .A1(n16340), .A2(n15586), .ZN(n13396) );
  INV_X1 U16422 ( .A(n15584), .ZN(n13604) );
  NAND2_X1 U16423 ( .A1(n13396), .A2(n13604), .ZN(n13208) );
  NAND2_X1 U16424 ( .A1(n15036), .A2(n19262), .ZN(n15019) );
  NAND2_X1 U16425 ( .A1(n15301), .A2(n15036), .ZN(n13210) );
  NAND2_X1 U16426 ( .A1(n14987), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13209) );
  OAI21_X1 U16427 ( .B1(n14247), .B2(n15019), .A(n13211), .ZN(P2_U2857) );
  AND2_X1 U16428 ( .A1(n14550), .A2(n14104), .ZN(n13212) );
  NAND2_X1 U16429 ( .A1(n13218), .A2(n13212), .ZN(n13217) );
  AOI22_X1 U16430 ( .A1(n14543), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14528), .ZN(n13213) );
  INV_X1 U16431 ( .A(n13213), .ZN(n13215) );
  INV_X1 U16432 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16409) );
  NOR2_X1 U16433 ( .A1(n13215), .A2(n13214), .ZN(n13216) );
  NAND2_X1 U16434 ( .A1(n13217), .A2(n13216), .ZN(P1_U2873) );
  NAND2_X1 U16435 ( .A1(n13218), .A2(n20154), .ZN(n13227) );
  INV_X1 U16436 ( .A(n14565), .ZN(n13219) );
  INV_X1 U16437 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14737) );
  NOR2_X1 U16438 ( .A1(n13219), .A2(n14737), .ZN(n13220) );
  AOI22_X1 U16439 ( .A1(n13221), .A2(n10313), .B1(n14567), .B2(n13220), .ZN(
        n13222) );
  INV_X1 U16440 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20839) );
  NOR2_X1 U16441 ( .A1(n20170), .A2(n20839), .ZN(n14730) );
  AOI21_X1 U16442 ( .B1(n20152), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14730), .ZN(n13223) );
  OAI21_X1 U16443 ( .B1(n20161), .B2(n13224), .A(n13223), .ZN(n13225) );
  NAND2_X1 U16444 ( .A1(n13227), .A2(n13226), .ZN(P1_U2968) );
  NOR2_X1 U16445 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13229) );
  NOR4_X1 U16446 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13228) );
  NAND4_X1 U16447 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13229), .A4(n13228), .ZN(n13241) );
  NOR2_X1 U16448 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13241), .ZN(n16481)
         );
  INV_X1 U16449 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n21002) );
  NOR3_X1 U16450 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        n21002), .ZN(n13231) );
  NOR4_X1 U16451 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n13230)
         );
  NAND4_X1 U16452 ( .A1(n14547), .A2(P1_W_R_N_REG_SCAN_IN), .A3(n13231), .A4(
        n13230), .ZN(U214) );
  NOR4_X1 U16453 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13235) );
  NOR4_X1 U16454 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n13234) );
  NOR4_X1 U16455 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13233) );
  NOR4_X1 U16456 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n13232) );
  NAND4_X1 U16457 ( .A1(n13235), .A2(n13234), .A3(n13233), .A4(n13232), .ZN(
        n13240) );
  NOR4_X1 U16458 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n13238) );
  NOR4_X1 U16459 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13237) );
  NOR4_X1 U16460 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13236) );
  INV_X1 U16461 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19843) );
  NAND4_X1 U16462 ( .A1(n13238), .A2(n13237), .A3(n13236), .A4(n19843), .ZN(
        n13239) );
  NOR2_X1 U16463 ( .A1(n13525), .A2(n13241), .ZN(n16408) );
  NAND2_X1 U16464 ( .A1(n16408), .A2(U214), .ZN(U212) );
  AOI211_X1 U16465 ( .C1(n15159), .C2(n9742), .A(n13242), .B(n19822), .ZN(
        n13253) );
  INV_X1 U16466 ( .A(n18996), .ZN(n19006) );
  OAI22_X1 U16467 ( .A1(n13244), .A2(n9646), .B1(n13243), .B2(n19006), .ZN(
        n13252) );
  INV_X1 U16468 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n13245) );
  OAI22_X1 U16469 ( .A1(n19017), .A2(n13245), .B1(n19880), .B2(n19035), .ZN(
        n13251) );
  NAND2_X1 U16470 ( .A1(n14956), .A2(n13246), .ZN(n13247) );
  NAND2_X1 U16471 ( .A1(n14846), .A2(n13247), .ZN(n15341) );
  INV_X1 U16472 ( .A(n19062), .ZN(n19036) );
  NAND2_X1 U16473 ( .A1(n15068), .A2(n13248), .ZN(n13249) );
  NAND2_X1 U16474 ( .A1(n9729), .A2(n13249), .ZN(n15061) );
  OAI22_X1 U16475 ( .A1(n15341), .A2(n19036), .B1(n15061), .B2(n19053), .ZN(
        n13250) );
  OR4_X1 U16476 ( .A1(n13253), .A2(n13252), .A3(n13251), .A4(n13250), .ZN(
        P2_U2828) );
  AOI211_X1 U16477 ( .C1(n15218), .C2(n13255), .A(n13254), .B(n19822), .ZN(
        n13267) );
  OAI22_X1 U16478 ( .A1(n15215), .A2(n19006), .B1(n19869), .B2(n19035), .ZN(
        n13266) );
  OAI22_X1 U16479 ( .A1(n13257), .A2(n9646), .B1(n13256), .B2(n19017), .ZN(
        n13265) );
  AND2_X1 U16480 ( .A1(n14877), .A2(n13258), .ZN(n13259) );
  OR2_X1 U16481 ( .A1(n13259), .A2(n9750), .ZN(n15414) );
  OR2_X1 U16482 ( .A1(n13260), .A2(n13261), .ZN(n13262) );
  AND2_X1 U16483 ( .A1(n13262), .A2(n13288), .ZN(n15419) );
  INV_X1 U16484 ( .A(n15419), .ZN(n13263) );
  OAI22_X1 U16485 ( .A1(n15414), .A2(n19036), .B1(n19053), .B2(n13263), .ZN(
        n13264) );
  OR4_X1 U16486 ( .A1(n13267), .A2(n13266), .A3(n13265), .A4(n13264), .ZN(
        P2_U2834) );
  AOI211_X1 U16487 ( .C1(n13270), .C2(n13269), .A(n13268), .B(n19822), .ZN(
        n13280) );
  INV_X1 U16488 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n13271) );
  OAI22_X1 U16489 ( .A1(n13271), .A2(n19006), .B1(n12856), .B2(n19035), .ZN(
        n13279) );
  OAI22_X1 U16490 ( .A1(n13272), .A2(n9646), .B1(n19017), .B2(n11084), .ZN(
        n13278) );
  OR2_X1 U16491 ( .A1(n9750), .A2(n13273), .ZN(n13274) );
  AND2_X1 U16492 ( .A1(n13285), .A2(n13274), .ZN(n16108) );
  INV_X1 U16493 ( .A(n16108), .ZN(n13276) );
  XNOR2_X1 U16494 ( .A(n13287), .B(n13275), .ZN(n15400) );
  OAI22_X1 U16495 ( .A1(n13276), .A2(n19036), .B1(n19053), .B2(n15400), .ZN(
        n13277) );
  OR4_X1 U16496 ( .A1(n13280), .A2(n13279), .A3(n13278), .A4(n13277), .ZN(
        P2_U2833) );
  AOI211_X1 U16497 ( .C1(n15192), .C2(n13282), .A(n13281), .B(n19822), .ZN(
        n13295) );
  OAI22_X1 U16498 ( .A1(n15188), .A2(n19006), .B1(n19872), .B2(n19035), .ZN(
        n13294) );
  INV_X1 U16499 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n14982) );
  OAI22_X1 U16500 ( .A1(n13283), .A2(n9646), .B1(n19017), .B2(n14982), .ZN(
        n13293) );
  INV_X1 U16501 ( .A(n14972), .ZN(n13284) );
  AOI21_X1 U16502 ( .B1(n13286), .B2(n13285), .A(n13284), .ZN(n15382) );
  INV_X1 U16503 ( .A(n15382), .ZN(n15189) );
  INV_X1 U16504 ( .A(n13287), .ZN(n13289) );
  NOR2_X1 U16505 ( .A1(n13289), .A2(n13288), .ZN(n13291) );
  OAI21_X1 U16506 ( .B1(n13291), .B2(n13290), .A(n15082), .ZN(n15384) );
  OAI22_X1 U16507 ( .A1(n15189), .A2(n19036), .B1(n19053), .B2(n15384), .ZN(
        n13292) );
  OR4_X1 U16508 ( .A1(n13295), .A2(n13294), .A3(n13293), .A4(n13292), .ZN(
        P2_U2832) );
  NAND2_X1 U16509 ( .A1(n13422), .A2(n13296), .ZN(n13304) );
  INV_X1 U16510 ( .A(n13297), .ZN(n13301) );
  NAND2_X1 U16511 ( .A1(n13654), .A2(n13298), .ZN(n13299) );
  AOI21_X1 U16512 ( .B1(n13301), .B2(n13300), .A(n13299), .ZN(n13302) );
  OR2_X1 U16513 ( .A1(n13715), .A2(n13302), .ZN(n13303) );
  MUX2_X1 U16514 ( .A(n13304), .B(n13303), .S(n14820), .Z(n13311) );
  AOI21_X1 U16515 ( .B1(n13305), .B2(n11622), .A(n20212), .ZN(n13306) );
  AND2_X1 U16516 ( .A1(n13307), .A2(n13306), .ZN(n13316) );
  NOR2_X1 U16517 ( .A1(n13308), .A2(n13316), .ZN(n13309) );
  OR2_X1 U16518 ( .A1(n13309), .A2(n12342), .ZN(n13559) );
  NAND3_X1 U16519 ( .A1(n13311), .A2(n13559), .A3(n13310), .ZN(n13312) );
  INV_X1 U16520 ( .A(n13338), .ZN(n13313) );
  NAND2_X1 U16521 ( .A1(n13313), .A2(n20170), .ZN(n20200) );
  INV_X1 U16522 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20198) );
  AND2_X1 U16523 ( .A1(n13314), .A2(n13717), .ZN(n13714) );
  NAND2_X1 U16524 ( .A1(n13338), .A2(n13714), .ZN(n14784) );
  AND2_X1 U16525 ( .A1(n13315), .A2(n13412), .ZN(n13317) );
  NOR2_X1 U16526 ( .A1(n13317), .A2(n13316), .ZN(n13325) );
  NAND2_X1 U16527 ( .A1(n11608), .A2(n11607), .ZN(n13324) );
  INV_X1 U16528 ( .A(n13927), .ZN(n13318) );
  OAI21_X1 U16529 ( .B1(n13804), .B2(n13319), .A(n13318), .ZN(n13321) );
  AOI21_X1 U16530 ( .B1(n13561), .B2(n11622), .A(n14104), .ZN(n13320) );
  AND3_X1 U16531 ( .A1(n13322), .A2(n13321), .A3(n13320), .ZN(n13323) );
  AND3_X1 U16532 ( .A1(n13325), .A2(n13324), .A3(n13323), .ZN(n13546) );
  MUX2_X1 U16533 ( .A(n13326), .B(n14820), .S(n13654), .Z(n13327) );
  NAND3_X1 U16534 ( .A1(n13546), .A2(n13328), .A3(n13327), .ZN(n13329) );
  NAND2_X1 U16535 ( .A1(n13338), .A2(n13329), .ZN(n14716) );
  NAND2_X1 U16536 ( .A1(n14784), .A2(n14716), .ZN(n13334) );
  NAND2_X1 U16537 ( .A1(n20198), .A2(n13334), .ZN(n20205) );
  AOI21_X1 U16538 ( .B1(n20200), .B2(n20205), .A(n13911), .ZN(n13346) );
  NOR2_X1 U16539 ( .A1(n13330), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13956) );
  INV_X1 U16540 ( .A(n13331), .ZN(n13955) );
  NAND2_X1 U16541 ( .A1(n13335), .A2(n13336), .ZN(n13332) );
  NAND4_X1 U16542 ( .A1(n9788), .A2(n13675), .A3(n15741), .A4(n13332), .ZN(
        n13333) );
  NOR3_X1 U16543 ( .A1(n13956), .A2(n13955), .A3(n20208), .ZN(n13345) );
  NAND2_X1 U16544 ( .A1(n13338), .A2(n15727), .ZN(n20199) );
  INV_X1 U16545 ( .A(n20199), .ZN(n15785) );
  AOI211_X1 U16546 ( .C1(n20198), .C2(n20199), .A(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n14787), .ZN(n13344) );
  OR2_X1 U16547 ( .A1(n13339), .A2(n13717), .ZN(n13341) );
  AND2_X1 U16548 ( .A1(n13341), .A2(n13340), .ZN(n13729) );
  INV_X1 U16549 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n13342) );
  OR2_X1 U16550 ( .A1(n20170), .A2(n13342), .ZN(n13952) );
  OAI21_X1 U16551 ( .B1(n16014), .B2(n13729), .A(n13952), .ZN(n13343) );
  OR4_X1 U16552 ( .A1(n13346), .A2(n13345), .A3(n13344), .A4(n13343), .ZN(
        P1_U3030) );
  INV_X1 U16553 ( .A(n13347), .ZN(n13402) );
  AND2_X1 U16554 ( .A1(n13402), .A2(n13348), .ZN(n14076) );
  INV_X1 U16555 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n19973) );
  NAND2_X1 U16556 ( .A1(n19902), .A2(n14188), .ZN(n18923) );
  OAI211_X1 U16557 ( .C1(n14076), .C2(n19973), .A(n13354), .B(n18923), .ZN(
        P2_U2814) );
  NOR2_X1 U16558 ( .A1(n19965), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n13349)
         );
  INV_X1 U16559 ( .A(n10609), .ZN(n19958) );
  AOI22_X1 U16560 ( .A1(n13349), .A2(n18923), .B1(n19958), .B2(n19965), .ZN(
        P2_U3612) );
  NAND2_X1 U16561 ( .A1(n10609), .A2(n19967), .ZN(n13350) );
  AND3_X1 U16562 ( .A1(n16333), .A2(n13350), .A3(n13378), .ZN(n13351) );
  NAND2_X1 U16563 ( .A1(n16335), .A2(n13351), .ZN(n16348) );
  AND2_X1 U16564 ( .A1(n16348), .A2(n19819), .ZN(n19942) );
  OAI21_X1 U16565 ( .B1(n13353), .B2(n19942), .A(n13352), .ZN(P2_U2819) );
  OAI21_X1 U16566 ( .B1(n19960), .B2(n13354), .A(n13626), .ZN(n13499) );
  INV_X1 U16567 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n13357) );
  NAND3_X1 U16568 ( .A1(n13355), .A2(n19956), .A3(n19967), .ZN(n13627) );
  AOI22_X1 U16569 ( .A1(n19219), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13525), .ZN(n19243) );
  NOR2_X1 U16570 ( .A1(n13627), .A2(n19243), .ZN(n13508) );
  AOI21_X1 U16571 ( .B1(P2_EAX_REG_3__SCAN_IN), .B2(n13532), .A(n13508), .ZN(
        n13356) );
  OAI21_X1 U16572 ( .B1(n13499), .B2(n13357), .A(n13356), .ZN(P2_U2970) );
  INV_X1 U16573 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n13362) );
  INV_X1 U16574 ( .A(n13627), .ZN(n13441) );
  INV_X1 U16575 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16433) );
  OR2_X1 U16576 ( .A1(n19217), .A2(n16433), .ZN(n13359) );
  NAND2_X1 U16577 ( .A1(n19217), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13358) );
  AND2_X1 U16578 ( .A1(n13359), .A2(n13358), .ZN(n19092) );
  INV_X1 U16579 ( .A(n19092), .ZN(n13360) );
  NAND2_X1 U16580 ( .A1(n13441), .A2(n13360), .ZN(n13431) );
  NAND2_X1 U16581 ( .A1(n13532), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n13361) );
  OAI211_X1 U16582 ( .C1(n13499), .C2(n13362), .A(n13431), .B(n13361), .ZN(
        P2_U2980) );
  INV_X1 U16583 ( .A(P2_LWORD_REG_9__SCAN_IN), .ZN(n13367) );
  INV_X1 U16584 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16441) );
  OR2_X1 U16585 ( .A1(n13525), .A2(n16441), .ZN(n13364) );
  NAND2_X1 U16586 ( .A1(n19217), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13363) );
  AND2_X1 U16587 ( .A1(n13364), .A2(n13363), .ZN(n19104) );
  INV_X1 U16588 ( .A(n19104), .ZN(n13365) );
  NAND2_X1 U16589 ( .A1(n13441), .A2(n13365), .ZN(n13439) );
  NAND2_X1 U16590 ( .A1(n13532), .A2(P2_EAX_REG_9__SCAN_IN), .ZN(n13366) );
  OAI211_X1 U16591 ( .C1(n13499), .C2(n13367), .A(n13439), .B(n13366), .ZN(
        P2_U2976) );
  INV_X1 U16592 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n13372) );
  INV_X1 U16593 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16437) );
  OR2_X1 U16594 ( .A1(n19217), .A2(n16437), .ZN(n13369) );
  NAND2_X1 U16595 ( .A1(n19217), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13368) );
  AND2_X1 U16596 ( .A1(n13369), .A2(n13368), .ZN(n19098) );
  INV_X1 U16597 ( .A(n19098), .ZN(n13370) );
  NAND2_X1 U16598 ( .A1(n13441), .A2(n13370), .ZN(n13428) );
  NAND2_X1 U16599 ( .A1(n13532), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n13371) );
  OAI211_X1 U16600 ( .C1(n13499), .C2(n13372), .A(n13428), .B(n13371), .ZN(
        P2_U2978) );
  INV_X1 U16601 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13374) );
  AOI22_X1 U16602 ( .A1(n19219), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19217), .ZN(n19086) );
  INV_X1 U16603 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13373) );
  OAI222_X1 U16604 ( .A1(n13374), .A2(n13499), .B1(n13627), .B2(n19086), .C1(
        n13626), .C2(n13373), .ZN(P2_U2982) );
  NOR2_X1 U16605 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20719), .ZN(n14216) );
  AOI21_X1 U16606 ( .B1(n13375), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n14216), 
        .ZN(n13376) );
  NAND2_X1 U16607 ( .A1(n13773), .A2(n13376), .ZN(P1_U2801) );
  INV_X1 U16608 ( .A(n16340), .ZN(n13377) );
  NAND2_X1 U16609 ( .A1(n13377), .A2(n19956), .ZN(n13585) );
  OR2_X1 U16610 ( .A1(n13347), .A2(n13378), .ZN(n13399) );
  NAND2_X1 U16611 ( .A1(n13379), .A2(n13380), .ZN(n13390) );
  NAND2_X1 U16612 ( .A1(n13390), .A2(n16342), .ZN(n13381) );
  NAND2_X1 U16613 ( .A1(n13381), .A2(n19262), .ZN(n13382) );
  AOI21_X1 U16614 ( .B1(n13382), .B2(n19237), .A(n10603), .ZN(n13386) );
  NAND2_X1 U16615 ( .A1(n13383), .A2(n19237), .ZN(n13384) );
  NAND2_X1 U16616 ( .A1(n13347), .A2(n13384), .ZN(n13385) );
  NAND2_X1 U16617 ( .A1(n13386), .A2(n13385), .ZN(n13394) );
  INV_X1 U16618 ( .A(n13387), .ZN(n13389) );
  AOI21_X1 U16619 ( .B1(n13389), .B2(n19262), .A(n13388), .ZN(n13596) );
  NAND4_X1 U16620 ( .A1(n16335), .A2(n16333), .A3(n10609), .A4(n19967), .ZN(
        n13391) );
  OAI21_X1 U16621 ( .B1(n16340), .B2(n13593), .A(n13391), .ZN(n13452) );
  INV_X1 U16622 ( .A(n13452), .ZN(n13398) );
  NAND3_X1 U16623 ( .A1(n10593), .A2(n16333), .A3(n13587), .ZN(n13393) );
  NAND2_X1 U16624 ( .A1(n13393), .A2(n13392), .ZN(n13395) );
  NOR3_X1 U16625 ( .A1(n13395), .A2(n13596), .A3(n13394), .ZN(n13581) );
  AND2_X1 U16626 ( .A1(n13396), .A2(n13581), .ZN(n13397) );
  OAI211_X1 U16627 ( .C1(n13585), .C2(n13399), .A(n13398), .B(n13397), .ZN(
        n16352) );
  NAND2_X1 U16628 ( .A1(n16352), .A2(n19819), .ZN(n13401) );
  NAND2_X1 U16629 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19936), .ZN(n16369) );
  INV_X1 U16630 ( .A(n16369), .ZN(n16371) );
  AOI22_X1 U16631 ( .A1(n16371), .A2(P2_FLUSH_REG_SCAN_IN), .B1(
        P2_STATE2_REG_3__SCAN_IN), .B2(n9877), .ZN(n13400) );
  NAND4_X1 U16632 ( .A1(n13402), .A2(n13380), .A3(n19900), .A4(n16341), .ZN(
        n13404) );
  NAND2_X1 U16633 ( .A1(n15607), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13403) );
  OAI21_X1 U16634 ( .B1(n15607), .B2(n13404), .A(n13403), .ZN(P2_U3595) );
  INV_X1 U16635 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13407) );
  NAND2_X1 U16636 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19931), .ZN(n13405) );
  NOR2_X1 U16637 ( .A1(n12904), .A2(n13405), .ZN(n13406) );
  OAI21_X1 U16638 ( .B1(n13380), .B2(n13407), .A(n13406), .ZN(n13408) );
  MUX2_X1 U16639 ( .A(n13613), .B(n13410), .S(n14987), .Z(n13411) );
  OAI21_X1 U16640 ( .B1(n19933), .B2(n15019), .A(n13411), .ZN(P2_U2887) );
  NOR2_X1 U16641 ( .A1(P1_READREQUEST_REG_SCAN_IN), .A2(n14216), .ZN(n13414)
         );
  OAI21_X1 U16642 ( .B1(n11607), .B2(n13412), .A(n20869), .ZN(n13413) );
  OAI21_X1 U16643 ( .B1(n13414), .B2(n20869), .A(n13413), .ZN(P1_U3487) );
  AND2_X1 U16644 ( .A1(n13415), .A2(n13420), .ZN(n13416) );
  AOI21_X1 U16645 ( .B1(n13715), .B2(n13417), .A(n13416), .ZN(n19976) );
  INV_X1 U16646 ( .A(n13553), .ZN(n15751) );
  NAND2_X1 U16647 ( .A1(n13927), .A2(n20871), .ZN(n13418) );
  NAND2_X1 U16648 ( .A1(n13418), .A2(n13553), .ZN(n20877) );
  OAI21_X1 U16649 ( .B1(n15751), .B2(n13770), .A(n20877), .ZN(n13419) );
  AND2_X1 U16650 ( .A1(n19976), .A2(n13419), .ZN(n15744) );
  NOR2_X1 U16651 ( .A1(n15744), .A2(n15762), .ZN(n19984) );
  INV_X1 U16652 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n20919) );
  INV_X1 U16653 ( .A(n13714), .ZN(n13557) );
  AND3_X1 U16654 ( .A1(n13420), .A2(n15741), .A3(n13675), .ZN(n13421) );
  MUX2_X1 U16655 ( .A(n13557), .B(n13421), .S(n13715), .Z(n13425) );
  INV_X1 U16656 ( .A(n13422), .ZN(n13423) );
  NAND2_X1 U16657 ( .A1(n12342), .A2(n13423), .ZN(n13424) );
  AND2_X1 U16658 ( .A1(n13425), .A2(n13424), .ZN(n15747) );
  INV_X1 U16659 ( .A(n15747), .ZN(n13426) );
  NAND2_X1 U16660 ( .A1(n19984), .A2(n13426), .ZN(n13427) );
  OAI21_X1 U16661 ( .B1(n19984), .B2(n20919), .A(n13427), .ZN(P1_U3484) );
  INV_X1 U16662 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n15062) );
  INV_X1 U16663 ( .A(n13499), .ZN(n13445) );
  NAND2_X1 U16664 ( .A1(n13445), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13429) );
  OAI211_X1 U16665 ( .C1(n13626), .C2(n15062), .A(n13429), .B(n13428), .ZN(
        P2_U2963) );
  INV_X1 U16666 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13538) );
  NAND2_X1 U16667 ( .A1(n13445), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13430) );
  MUX2_X1 U16668 ( .A(BUF1_REG_8__SCAN_IN), .B(BUF2_REG_8__SCAN_IN), .S(n13525), .Z(n19108) );
  NAND2_X1 U16669 ( .A1(n13441), .A2(n19108), .ZN(n13435) );
  OAI211_X1 U16670 ( .C1(n13538), .C2(n13626), .A(n13430), .B(n13435), .ZN(
        P2_U2960) );
  INV_X1 U16671 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n15050) );
  NAND2_X1 U16672 ( .A1(n13445), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13432) );
  OAI211_X1 U16673 ( .C1(n13626), .C2(n15050), .A(n13432), .B(n13431), .ZN(
        P2_U2965) );
  INV_X1 U16674 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13540) );
  NAND2_X1 U16675 ( .A1(n13445), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13433) );
  MUX2_X1 U16676 ( .A(BUF1_REG_12__SCAN_IN), .B(BUF2_REG_12__SCAN_IN), .S(
        n13525), .Z(n19095) );
  NAND2_X1 U16677 ( .A1(n13441), .A2(n19095), .ZN(n13446) );
  OAI211_X1 U16678 ( .C1(n13540), .C2(n13626), .A(n13433), .B(n13446), .ZN(
        P2_U2964) );
  INV_X1 U16679 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13699) );
  NAND2_X1 U16680 ( .A1(n13445), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13434) );
  MUX2_X1 U16681 ( .A(BUF1_REG_10__SCAN_IN), .B(BUF2_REG_10__SCAN_IN), .S(
        n19217), .Z(n19101) );
  NAND2_X1 U16682 ( .A1(n13441), .A2(n19101), .ZN(n13437) );
  OAI211_X1 U16683 ( .C1(n13699), .C2(n13626), .A(n13434), .B(n13437), .ZN(
        P2_U2962) );
  INV_X1 U16684 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19156) );
  NAND2_X1 U16685 ( .A1(n13445), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13436) );
  OAI211_X1 U16686 ( .C1(n19156), .C2(n13626), .A(n13436), .B(n13435), .ZN(
        P2_U2975) );
  INV_X1 U16687 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19151) );
  NAND2_X1 U16688 ( .A1(n13445), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13438) );
  OAI211_X1 U16689 ( .C1(n19151), .C2(n13626), .A(n13438), .B(n13437), .ZN(
        P2_U2977) );
  INV_X1 U16690 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n15076) );
  NAND2_X1 U16691 ( .A1(n13445), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13440) );
  OAI211_X1 U16692 ( .C1(n13626), .C2(n15076), .A(n13440), .B(n13439), .ZN(
        P2_U2961) );
  INV_X1 U16693 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19143) );
  NAND2_X1 U16694 ( .A1(n13445), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13442) );
  MUX2_X1 U16695 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n13525), .Z(n19089) );
  NAND2_X1 U16696 ( .A1(n13441), .A2(n19089), .ZN(n13443) );
  OAI211_X1 U16697 ( .C1(n19143), .C2(n13626), .A(n13442), .B(n13443), .ZN(
        P2_U2981) );
  INV_X1 U16698 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13479) );
  NAND2_X1 U16699 ( .A1(n13445), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13444) );
  OAI211_X1 U16700 ( .C1(n13479), .C2(n13626), .A(n13444), .B(n13443), .ZN(
        P2_U2966) );
  INV_X1 U16701 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19147) );
  NAND2_X1 U16702 ( .A1(n13445), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13447) );
  OAI211_X1 U16703 ( .C1(n19147), .C2(n13626), .A(n13447), .B(n13446), .ZN(
        P2_U2979) );
  INV_X1 U16704 ( .A(n13448), .ZN(n13449) );
  AND2_X1 U16705 ( .A1(n13450), .A2(n13449), .ZN(n13451) );
  AND2_X1 U16706 ( .A1(n19121), .A2(n13454), .ZN(n19077) );
  NAND2_X1 U16707 ( .A1(n19121), .A2(n9887), .ZN(n14242) );
  NAND2_X1 U16708 ( .A1(n15116), .A2(n14242), .ZN(n19107) );
  INV_X1 U16709 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16462) );
  INV_X1 U16710 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18230) );
  AOI22_X1 U16711 ( .A1(n19219), .A2(n16462), .B1(n18230), .B2(n19217), .ZN(
        n19076) );
  INV_X1 U16712 ( .A(n19076), .ZN(n19225) );
  INV_X1 U16713 ( .A(n13456), .ZN(n13462) );
  INV_X1 U16714 ( .A(n13457), .ZN(n13460) );
  INV_X1 U16715 ( .A(n13458), .ZN(n13459) );
  NAND2_X1 U16716 ( .A1(n13460), .A2(n13459), .ZN(n13461) );
  NAND2_X1 U16717 ( .A1(n13462), .A2(n13461), .ZN(n13614) );
  INV_X1 U16718 ( .A(n13614), .ZN(n19057) );
  NOR2_X1 U16719 ( .A1(n19933), .A2(n13614), .ZN(n19134) );
  INV_X1 U16720 ( .A(n19134), .ZN(n13464) );
  OAI211_X1 U16721 ( .C1(n19479), .C2(n19057), .A(n13464), .B(n19085), .ZN(
        n13467) );
  NAND2_X1 U16722 ( .A1(n19121), .A2(n13465), .ZN(n19122) );
  AOI22_X1 U16723 ( .A1(n19131), .A2(n19057), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19130), .ZN(n13466) );
  OAI211_X1 U16724 ( .C1(n19139), .C2(n19225), .A(n13467), .B(n13466), .ZN(
        P2_U2919) );
  MUX2_X1 U16725 ( .A(n19207), .B(n14070), .S(n14987), .Z(n13472) );
  OAI21_X1 U16726 ( .B1(n19903), .B2(n15019), .A(n13472), .ZN(P2_U2886) );
  INV_X1 U16727 ( .A(n19819), .ZN(n13473) );
  OR2_X1 U16728 ( .A1(n13347), .A2(n13473), .ZN(n13474) );
  OAI21_X1 U16729 ( .B1(n13585), .B2(n13474), .A(n13626), .ZN(n13475) );
  INV_X1 U16730 ( .A(n19830), .ZN(n19955) );
  NAND2_X1 U16731 ( .A1(n19140), .A2(n13476), .ZN(n13703) );
  INV_X1 U16732 ( .A(n19936), .ZN(n13477) );
  NOR2_X1 U16733 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13477), .ZN(n13701) );
  AOI22_X1 U16734 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n19154), .B1(n13701), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13478) );
  OAI21_X1 U16735 ( .B1(n13479), .B2(n13703), .A(n13478), .ZN(P2_U2921) );
  XOR2_X1 U16736 ( .A(n19060), .B(n13483), .Z(n13620) );
  AND2_X1 U16737 ( .A1(n19192), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13616) );
  INV_X1 U16738 ( .A(n13480), .ZN(n13481) );
  AOI21_X1 U16739 ( .B1(n13483), .B2(n13482), .A(n13481), .ZN(n13619) );
  AND2_X1 U16740 ( .A1(n11014), .A2(n13619), .ZN(n13484) );
  AOI211_X1 U16741 ( .C1(n19188), .C2(n13620), .A(n13616), .B(n13484), .ZN(
        n13487) );
  OAI21_X1 U16742 ( .B1(n19187), .B2(n13485), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13486) );
  OAI211_X1 U16743 ( .C1(n19218), .C2(n13613), .A(n13487), .B(n13486), .ZN(
        P2_U3014) );
  AOI21_X1 U16744 ( .B1(n13490), .B2(n13489), .A(n13488), .ZN(n13632) );
  OAI22_X1 U16745 ( .A1(n16227), .A2(n13491), .B1(n19841), .B2(n19033), .ZN(
        n13493) );
  NOR2_X1 U16746 ( .A1(n19182), .A2(n14041), .ZN(n13492) );
  AOI211_X1 U16747 ( .C1(n13632), .C2(n11014), .A(n13493), .B(n13492), .ZN(
        n13498) );
  INV_X1 U16748 ( .A(n13494), .ZN(n13495) );
  XNOR2_X1 U16749 ( .A(n13496), .B(n13495), .ZN(n13640) );
  NAND2_X1 U16750 ( .A1(n13640), .A2(n19188), .ZN(n13497) );
  OAI211_X1 U16751 ( .C1(n19218), .C2(n13648), .A(n13498), .B(n13497), .ZN(
        P2_U3012) );
  INV_X1 U16752 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n13501) );
  AOI22_X1 U16753 ( .A1(n19219), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19217), .ZN(n19264) );
  NOR2_X1 U16754 ( .A1(n13627), .A2(n19264), .ZN(n13522) );
  AOI21_X1 U16755 ( .B1(n13532), .B2(P2_EAX_REG_7__SCAN_IN), .A(n13522), .ZN(
        n13500) );
  OAI21_X1 U16756 ( .B1(n13625), .B2(n13501), .A(n13500), .ZN(P2_U2974) );
  INV_X1 U16757 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n13503) );
  INV_X1 U16758 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16452) );
  INV_X1 U16759 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18249) );
  AOI22_X1 U16760 ( .A1(n19219), .A2(n16452), .B1(n18249), .B2(n19217), .ZN(
        n16095) );
  INV_X1 U16761 ( .A(n16095), .ZN(n19246) );
  NOR2_X1 U16762 ( .A1(n13627), .A2(n19246), .ZN(n13514) );
  AOI21_X1 U16763 ( .B1(P2_EAX_REG_4__SCAN_IN), .B2(n13532), .A(n13514), .ZN(
        n13502) );
  OAI21_X1 U16764 ( .B1(n13625), .B2(n13503), .A(n13502), .ZN(P2_U2971) );
  INV_X1 U16765 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n13505) );
  AOI22_X1 U16766 ( .A1(n19219), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13525), .ZN(n19252) );
  NOR2_X1 U16767 ( .A1(n13627), .A2(n19252), .ZN(n13517) );
  AOI21_X1 U16768 ( .B1(P2_EAX_REG_5__SCAN_IN), .B2(n13532), .A(n13517), .ZN(
        n13504) );
  OAI21_X1 U16769 ( .B1(n13625), .B2(n13505), .A(n13504), .ZN(P2_U2972) );
  INV_X1 U16770 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n13507) );
  AOI22_X1 U16771 ( .A1(n19219), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13525), .ZN(n19233) );
  NOR2_X1 U16772 ( .A1(n13627), .A2(n19233), .ZN(n13511) );
  AOI21_X1 U16773 ( .B1(P2_EAX_REG_1__SCAN_IN), .B2(n13532), .A(n13511), .ZN(
        n13506) );
  OAI21_X1 U16774 ( .B1(n13625), .B2(n13507), .A(n13506), .ZN(P2_U2968) );
  INV_X1 U16775 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n13510) );
  AOI21_X1 U16776 ( .B1(n13532), .B2(P2_EAX_REG_19__SCAN_IN), .A(n13508), .ZN(
        n13509) );
  OAI21_X1 U16777 ( .B1(n13625), .B2(n13510), .A(n13509), .ZN(P2_U2955) );
  INV_X1 U16778 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n13513) );
  AOI21_X1 U16779 ( .B1(n13532), .B2(P2_EAX_REG_17__SCAN_IN), .A(n13511), .ZN(
        n13512) );
  OAI21_X1 U16780 ( .B1(n13625), .B2(n13513), .A(n13512), .ZN(P2_U2953) );
  INV_X1 U16781 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n13516) );
  AOI21_X1 U16782 ( .B1(P2_EAX_REG_20__SCAN_IN), .B2(n13532), .A(n13514), .ZN(
        n13515) );
  OAI21_X1 U16783 ( .B1(n13625), .B2(n13516), .A(n13515), .ZN(P2_U2956) );
  INV_X1 U16784 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n13519) );
  AOI21_X1 U16785 ( .B1(n13532), .B2(P2_EAX_REG_21__SCAN_IN), .A(n13517), .ZN(
        n13518) );
  OAI21_X1 U16786 ( .B1(n13625), .B2(n13519), .A(n13518), .ZN(P2_U2957) );
  INV_X1 U16787 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n13521) );
  INV_X1 U16788 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16456) );
  INV_X1 U16789 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18240) );
  AOI22_X1 U16790 ( .A1(n19219), .A2(n16456), .B1(n18240), .B2(n19217), .ZN(
        n16102) );
  INV_X1 U16791 ( .A(n16102), .ZN(n19238) );
  NOR2_X1 U16792 ( .A1(n13627), .A2(n19238), .ZN(n13531) );
  AOI21_X1 U16793 ( .B1(P2_EAX_REG_2__SCAN_IN), .B2(n13532), .A(n13531), .ZN(
        n13520) );
  OAI21_X1 U16794 ( .B1(n13625), .B2(n13521), .A(n13520), .ZN(P2_U2969) );
  INV_X1 U16795 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n13524) );
  AOI21_X1 U16796 ( .B1(n13532), .B2(P2_EAX_REG_23__SCAN_IN), .A(n13522), .ZN(
        n13523) );
  OAI21_X1 U16797 ( .B1(n13625), .B2(n13524), .A(n13523), .ZN(P2_U2959) );
  INV_X1 U16798 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n13527) );
  AOI22_X1 U16799 ( .A1(n19219), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13525), .ZN(n19255) );
  NOR2_X1 U16800 ( .A1(n13627), .A2(n19255), .ZN(n13528) );
  AOI21_X1 U16801 ( .B1(n13532), .B2(P2_EAX_REG_6__SCAN_IN), .A(n13528), .ZN(
        n13526) );
  OAI21_X1 U16802 ( .B1(n13625), .B2(n13527), .A(n13526), .ZN(P2_U2973) );
  INV_X1 U16803 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n13530) );
  AOI21_X1 U16804 ( .B1(n13532), .B2(P2_EAX_REG_22__SCAN_IN), .A(n13528), .ZN(
        n13529) );
  OAI21_X1 U16805 ( .B1(n13625), .B2(n13530), .A(n13529), .ZN(P2_U2958) );
  INV_X1 U16806 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n13534) );
  AOI21_X1 U16807 ( .B1(P2_EAX_REG_18__SCAN_IN), .B2(n13532), .A(n13531), .ZN(
        n13533) );
  OAI21_X1 U16808 ( .B1(n13625), .B2(n13534), .A(n13533), .ZN(P2_U2954) );
  INV_X1 U16809 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n15089) );
  AOI22_X1 U16810 ( .A1(n13701), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19154), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13535) );
  OAI21_X1 U16811 ( .B1(n15089), .B2(n13703), .A(n13535), .ZN(P2_U2928) );
  AOI22_X1 U16812 ( .A1(n13701), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19154), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13536) );
  OAI21_X1 U16813 ( .B1(n15076), .B2(n13703), .A(n13536), .ZN(P2_U2926) );
  AOI22_X1 U16814 ( .A1(n13701), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19154), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13537) );
  OAI21_X1 U16815 ( .B1(n13538), .B2(n13703), .A(n13537), .ZN(P2_U2927) );
  AOI22_X1 U16816 ( .A1(n13701), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19154), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13539) );
  OAI21_X1 U16817 ( .B1(n13540), .B2(n13703), .A(n13539), .ZN(P2_U2923) );
  AOI22_X1 U16818 ( .A1(n13701), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19154), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13541) );
  OAI21_X1 U16819 ( .B1(n15062), .B2(n13703), .A(n13541), .ZN(P2_U2924) );
  INV_X1 U16820 ( .A(n13542), .ZN(n13544) );
  AND3_X1 U16821 ( .A1(n13297), .A2(n13544), .A3(n13543), .ZN(n13545) );
  NAND3_X1 U16822 ( .A1(n12594), .A2(n13546), .A3(n13545), .ZN(n13817) );
  INV_X1 U16823 ( .A(n13817), .ZN(n13671) );
  NOR2_X1 U16824 ( .A1(n11513), .A2(n13810), .ZN(n13549) );
  AOI22_X1 U16825 ( .A1(n15727), .A2(n11687), .B1(n13549), .B2(n13547), .ZN(
        n13548) );
  OAI21_X1 U16826 ( .B1(n20455), .B2(n13671), .A(n13548), .ZN(n15730) );
  INV_X1 U16827 ( .A(n13549), .ZN(n13551) );
  INV_X1 U16828 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14727) );
  AOI22_X1 U16829 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n13911), .B2(n14727), .ZN(
        n13686) );
  NOR2_X1 U16830 ( .A1(n16053), .A2(n20198), .ZN(n13685) );
  INV_X1 U16831 ( .A(n13685), .ZN(n13550) );
  OAI22_X1 U16832 ( .A1(n13837), .A2(n13551), .B1(n13686), .B2(n13550), .ZN(
        n13552) );
  AOI21_X1 U16833 ( .B1(n15730), .B2(n20857), .A(n13552), .ZN(n13570) );
  NAND2_X1 U16834 ( .A1(n13297), .A2(n13675), .ZN(n13556) );
  NAND2_X1 U16835 ( .A1(n13554), .A2(n13553), .ZN(n13555) );
  OAI21_X1 U16836 ( .B1(n15727), .B2(n13556), .A(n13555), .ZN(n13558) );
  MUX2_X1 U16837 ( .A(n13558), .B(n13557), .S(n13715), .Z(n13564) );
  OAI211_X1 U16838 ( .C1(n13927), .C2(n13561), .A(n13560), .B(n13559), .ZN(
        n13562) );
  INV_X1 U16839 ( .A(n13562), .ZN(n13563) );
  NAND2_X1 U16840 ( .A1(n13564), .A2(n13563), .ZN(n15725) );
  NAND2_X1 U16841 ( .A1(n15725), .A2(n19975), .ZN(n13568) );
  INV_X1 U16842 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19983) );
  NAND2_X1 U16843 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16054) );
  NOR3_X1 U16844 ( .A1(n16055), .A2(n19983), .A3(n16054), .ZN(n13566) );
  NOR2_X1 U16845 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20590), .ZN(n13565) );
  NOR2_X1 U16846 ( .A1(n13566), .A2(n13565), .ZN(n13567) );
  NAND2_X1 U16847 ( .A1(n20860), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13569) );
  OAI21_X1 U16848 ( .B1(n13570), .B2(n20860), .A(n13569), .ZN(P1_U3473) );
  AOI21_X1 U16849 ( .B1(n15727), .B2(n20857), .A(n20860), .ZN(n13577) );
  NOR2_X1 U16850 ( .A1(n13571), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13572) );
  AOI21_X1 U16851 ( .B1(n9664), .B2(n13817), .A(n13572), .ZN(n15729) );
  INV_X1 U16852 ( .A(n15729), .ZN(n13574) );
  OAI22_X1 U16853 ( .A1(n13837), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n16053), .ZN(n13573) );
  AOI21_X1 U16854 ( .B1(n13574), .B2(n20857), .A(n13573), .ZN(n13575) );
  OAI22_X1 U16855 ( .A1(n13577), .A2(n13576), .B1(n13575), .B2(n20860), .ZN(
        P1_U3474) );
  AOI21_X1 U16856 ( .B1(n13578), .B2(n16342), .A(n10553), .ZN(n13583) );
  MUX2_X1 U16857 ( .A(n10593), .B(n13586), .S(n13380), .Z(n13579) );
  NAND3_X1 U16858 ( .A1(n13579), .A2(n16333), .A3(n19967), .ZN(n13580) );
  NAND2_X1 U16859 ( .A1(n13581), .A2(n13580), .ZN(n13582) );
  AOI21_X1 U16860 ( .B1(n13585), .B2(n13583), .A(n13582), .ZN(n13591) );
  INV_X1 U16861 ( .A(n13584), .ZN(n13590) );
  INV_X1 U16862 ( .A(n13585), .ZN(n13588) );
  NAND3_X1 U16863 ( .A1(n13588), .A2(n13587), .A3(n13586), .ZN(n13589) );
  NAND3_X1 U16864 ( .A1(n13591), .A2(n13590), .A3(n13589), .ZN(n13592) );
  INV_X1 U16865 ( .A(n13593), .ZN(n16336) );
  INV_X1 U16866 ( .A(n14012), .ZN(n15455) );
  MUX2_X1 U16867 ( .A(n13594), .B(n19237), .S(n19220), .Z(n13599) );
  AND2_X1 U16868 ( .A1(n13595), .A2(n19956), .ZN(n14177) );
  OAI21_X1 U16869 ( .B1(n14177), .B2(n13596), .A(n19242), .ZN(n13598) );
  OAI21_X1 U16870 ( .B1(n10603), .B2(n13379), .A(n19958), .ZN(n13597) );
  AND3_X1 U16871 ( .A1(n13599), .A2(n13598), .A3(n13597), .ZN(n13603) );
  INV_X1 U16872 ( .A(n13600), .ZN(n13601) );
  NAND2_X1 U16873 ( .A1(n13601), .A2(n10603), .ZN(n13602) );
  AND2_X1 U16874 ( .A1(n13603), .A2(n13602), .ZN(n14176) );
  NAND2_X1 U16875 ( .A1(n14176), .A2(n13604), .ZN(n13605) );
  NAND2_X1 U16876 ( .A1(n13618), .A2(n13605), .ZN(n15456) );
  NAND2_X1 U16877 ( .A1(n15455), .A2(n15456), .ZN(n19201) );
  INV_X1 U16878 ( .A(n19201), .ZN(n15427) );
  INV_X1 U16879 ( .A(n13618), .ZN(n13606) );
  NAND2_X1 U16880 ( .A1(n13606), .A2(n19033), .ZN(n13634) );
  INV_X1 U16881 ( .A(n13634), .ZN(n19212) );
  INV_X1 U16882 ( .A(n15586), .ZN(n16339) );
  NAND2_X1 U16883 ( .A1(n16335), .A2(n19956), .ZN(n13607) );
  NAND2_X1 U16884 ( .A1(n16339), .A2(n13607), .ZN(n13608) );
  INV_X1 U16885 ( .A(n15585), .ZN(n13611) );
  NAND2_X1 U16886 ( .A1(n13609), .A2(n13380), .ZN(n13610) );
  NAND2_X1 U16887 ( .A1(n13611), .A2(n13610), .ZN(n13612) );
  NAND2_X1 U16888 ( .A1(n13618), .A2(n13612), .ZN(n19206) );
  OAI22_X1 U16889 ( .A1(n16306), .A2(n13614), .B1(n13613), .B2(n19206), .ZN(
        n13615) );
  AOI211_X1 U16890 ( .C1(n19212), .C2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13616), .B(n13615), .ZN(n13622) );
  NOR2_X1 U16891 ( .A1(n16343), .A2(n13617), .ZN(n19943) );
  AOI22_X1 U16892 ( .A1(n16309), .A2(n13620), .B1(n19204), .B2(n13619), .ZN(
        n13621) );
  OAI211_X1 U16893 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n15427), .A(
        n13622), .B(n13621), .ZN(P2_U3046) );
  INV_X1 U16894 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n13623) );
  OAI222_X1 U16895 ( .A1(n13623), .A2(n13625), .B1(n13627), .B2(n19225), .C1(
        n13626), .C2(n19173), .ZN(P2_U2967) );
  INV_X1 U16896 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13694) );
  INV_X1 U16897 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13624) );
  OAI222_X1 U16898 ( .A1(n13627), .A2(n19225), .B1(n13626), .B2(n13694), .C1(
        n13625), .C2(n13624), .ZN(P2_U2952) );
  AOI21_X1 U16899 ( .B1(n13630), .B2(n13629), .A(n13628), .ZN(n19915) );
  NOR2_X1 U16900 ( .A1(n13648), .A2(n19206), .ZN(n13639) );
  NOR2_X1 U16901 ( .A1(n15456), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14008) );
  AND2_X1 U16902 ( .A1(n14012), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13631) );
  NAND2_X1 U16903 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14010) );
  INV_X1 U16904 ( .A(n14010), .ZN(n19216) );
  OAI21_X1 U16905 ( .B1(n14008), .B2(n13631), .A(n19216), .ZN(n13637) );
  AOI22_X1 U16906 ( .A1(P2_REIP_REG_2__SCAN_IN), .A2(n19192), .B1(n19204), 
        .B2(n13632), .ZN(n13636) );
  NOR2_X1 U16907 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19216), .ZN(
        n13633) );
  NAND2_X1 U16908 ( .A1(n14012), .A2(n13633), .ZN(n14005) );
  OAI21_X1 U16909 ( .B1(n15456), .B2(n19216), .A(n13634), .ZN(n14004) );
  NAND2_X1 U16910 ( .A1(n14004), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13635) );
  NAND4_X1 U16911 ( .A1(n13637), .A2(n13636), .A3(n14005), .A4(n13635), .ZN(
        n13638) );
  AOI211_X1 U16912 ( .C1(n16309), .C2(n13640), .A(n13639), .B(n13638), .ZN(
        n13641) );
  OAI21_X1 U16913 ( .B1(n19915), .B2(n16306), .A(n13641), .ZN(P2_U3044) );
  INV_X1 U16914 ( .A(n20860), .ZN(n13644) );
  INV_X1 U16915 ( .A(n20347), .ZN(n20579) );
  XNOR2_X1 U16916 ( .A(n13642), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14423) );
  INV_X1 U16917 ( .A(n12594), .ZN(n13830) );
  NAND4_X1 U16918 ( .A1(n14423), .A2(n20857), .A3(n13830), .A4(n13644), .ZN(
        n13643) );
  OAI21_X1 U16919 ( .B1(n12327), .B2(n13644), .A(n13643), .ZN(P1_U3468) );
  MUX2_X1 U16920 ( .A(n13648), .B(n14044), .S(n14987), .Z(n13649) );
  OAI21_X1 U16921 ( .B1(n19913), .B2(n15019), .A(n13649), .ZN(P2_U2885) );
  INV_X1 U16922 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13656) );
  INV_X1 U16923 ( .A(n20875), .ZN(n13652) );
  AND2_X1 U16924 ( .A1(n13653), .A2(n13652), .ZN(n20076) );
  NAND2_X1 U16925 ( .A1(n20076), .A2(n13654), .ZN(n13798) );
  NOR2_X1 U16926 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16054), .ZN(n20102) );
  AOI22_X1 U16927 ( .A1(n20872), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n15781), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13655) );
  OAI21_X1 U16928 ( .B1(n13656), .B2(n13798), .A(n13655), .ZN(P1_U2915) );
  INV_X1 U16929 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13658) );
  AOI22_X1 U16930 ( .A1(n20872), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n15781), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13657) );
  OAI21_X1 U16931 ( .B1(n13658), .B2(n13798), .A(n13657), .ZN(P1_U2914) );
  INV_X1 U16932 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13660) );
  AOI22_X1 U16933 ( .A1(n20872), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n15781), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13659) );
  OAI21_X1 U16934 ( .B1(n13660), .B2(n13798), .A(n13659), .ZN(P1_U2908) );
  INV_X1 U16935 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13662) );
  AOI22_X1 U16936 ( .A1(n20872), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n15781), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13661) );
  OAI21_X1 U16937 ( .B1(n13662), .B2(n13798), .A(n13661), .ZN(P1_U2917) );
  AOI22_X1 U16938 ( .A1(n20872), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n15781), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13663) );
  OAI21_X1 U16939 ( .B1(n14497), .B2(n13798), .A(n13663), .ZN(P1_U2911) );
  AOI22_X1 U16940 ( .A1(n20872), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n15781), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13664) );
  OAI21_X1 U16941 ( .B1(n14488), .B2(n13798), .A(n13664), .ZN(P1_U2909) );
  INV_X1 U16942 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13666) );
  AOI22_X1 U16943 ( .A1(n20872), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n15781), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13665) );
  OAI21_X1 U16944 ( .B1(n13666), .B2(n13798), .A(n13665), .ZN(P1_U2918) );
  INV_X1 U16945 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13668) );
  AOI22_X1 U16946 ( .A1(n20872), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n15781), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13667) );
  OAI21_X1 U16947 ( .B1(n13668), .B2(n13798), .A(n13667), .ZN(P1_U2912) );
  AOI22_X1 U16948 ( .A1(n20872), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n15781), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13669) );
  OAI21_X1 U16949 ( .B1(n14506), .B2(n13798), .A(n13669), .ZN(P1_U2913) );
  AOI22_X1 U16950 ( .A1(n20872), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n15781), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13670) );
  OAI21_X1 U16951 ( .B1(n14519), .B2(n13798), .A(n13670), .ZN(P1_U2916) );
  OR2_X1 U16952 ( .A1(n10245), .A2(n13671), .ZN(n13683) );
  INV_X1 U16953 ( .A(n13672), .ZN(n13801) );
  INV_X1 U16954 ( .A(n13810), .ZN(n13673) );
  NAND2_X1 U16955 ( .A1(n13673), .A2(n11787), .ZN(n13808) );
  NAND2_X1 U16956 ( .A1(n13801), .A2(n13808), .ZN(n13677) );
  INV_X1 U16957 ( .A(n13677), .ZN(n13684) );
  NAND2_X1 U16958 ( .A1(n13804), .A2(n13684), .ZN(n13680) );
  NOR2_X1 U16959 ( .A1(n13674), .A2(n13805), .ZN(n13678) );
  INV_X1 U16960 ( .A(n13675), .ZN(n13676) );
  OR2_X1 U16961 ( .A1(n13676), .A2(n13714), .ZN(n13813) );
  AOI22_X1 U16962 ( .A1(n15727), .A2(n13678), .B1(n13813), .B2(n13677), .ZN(
        n13679) );
  OAI21_X1 U16963 ( .B1(n13817), .B2(n13680), .A(n13679), .ZN(n13681) );
  INV_X1 U16964 ( .A(n13681), .ZN(n13682) );
  NAND2_X1 U16965 ( .A1(n13683), .A2(n13682), .ZN(n15726) );
  INV_X1 U16966 ( .A(n13837), .ZN(n20856) );
  AOI222_X1 U16967 ( .A1(n15726), .A2(n20857), .B1(n13686), .B2(n13685), .C1(
        n13684), .C2(n20856), .ZN(n13688) );
  NAND2_X1 U16968 ( .A1(n20860), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13687) );
  OAI21_X1 U16969 ( .B1(n13688), .B2(n20860), .A(n13687), .ZN(P1_U3472) );
  INV_X1 U16970 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13690) );
  AOI22_X1 U16971 ( .A1(n19968), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19170), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13689) );
  OAI21_X1 U16972 ( .B1(n13690), .B2(n13703), .A(n13689), .ZN(P2_U2933) );
  AOI22_X1 U16973 ( .A1(n19968), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19170), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13691) );
  OAI21_X1 U16974 ( .B1(n15115), .B2(n13703), .A(n13691), .ZN(P2_U2934) );
  INV_X1 U16975 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n15107) );
  AOI22_X1 U16976 ( .A1(n19968), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19170), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13692) );
  OAI21_X1 U16977 ( .B1(n15107), .B2(n13703), .A(n13692), .ZN(P2_U2932) );
  AOI22_X1 U16978 ( .A1(n19968), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19170), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13693) );
  OAI21_X1 U16979 ( .B1(n13694), .B2(n13703), .A(n13693), .ZN(P2_U2935) );
  INV_X1 U16980 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15102) );
  AOI22_X1 U16981 ( .A1(n13701), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19170), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13695) );
  OAI21_X1 U16982 ( .B1(n15102), .B2(n13703), .A(n13695), .ZN(P2_U2930) );
  INV_X1 U16983 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13697) );
  AOI22_X1 U16984 ( .A1(n13701), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19170), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13696) );
  OAI21_X1 U16985 ( .B1(n13697), .B2(n13703), .A(n13696), .ZN(P2_U2931) );
  AOI22_X1 U16986 ( .A1(n13701), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19170), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13698) );
  OAI21_X1 U16987 ( .B1(n13699), .B2(n13703), .A(n13698), .ZN(P2_U2925) );
  AOI22_X1 U16988 ( .A1(n13701), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19170), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13700) );
  OAI21_X1 U16989 ( .B1(n15050), .B2(n13703), .A(n13700), .ZN(P2_U2922) );
  INV_X1 U16990 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n15095) );
  AOI22_X1 U16991 ( .A1(n13701), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19170), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13702) );
  OAI21_X1 U16992 ( .B1(n15095), .B2(n13703), .A(n13702), .ZN(P2_U2929) );
  INV_X1 U16993 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13708) );
  MUX2_X1 U16994 ( .A(n13709), .B(n13708), .S(n14987), .Z(n13710) );
  OAI21_X1 U16995 ( .B1(n19904), .B2(n15019), .A(n13710), .ZN(P2_U2884) );
  INV_X1 U16996 ( .A(n13711), .ZN(n13712) );
  AOI21_X1 U16997 ( .B1(n13713), .B2(n20198), .A(n13712), .ZN(n20204) );
  INV_X1 U16998 ( .A(n20204), .ZN(n13726) );
  NAND2_X1 U16999 ( .A1(n13715), .A2(n13714), .ZN(n13719) );
  NAND3_X1 U17000 ( .A1(n10309), .A2(n13717), .A3(n13716), .ZN(n13718) );
  NAND2_X1 U17001 ( .A1(n13719), .A2(n13718), .ZN(n13720) );
  INV_X1 U17002 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13938) );
  INV_X1 U17003 ( .A(n13721), .ZN(n13722) );
  AOI21_X1 U17004 ( .B1(n13724), .B2(n13723), .A(n13722), .ZN(n20168) );
  INV_X1 U17005 ( .A(n20168), .ZN(n13942) );
  OAI222_X1 U17006 ( .A1(n13726), .A2(n14467), .B1(n13938), .B2(n20075), .C1(
        n13942), .C2(n14480), .ZN(P1_U2872) );
  OAI21_X1 U17007 ( .B1(n13728), .B2(n13727), .A(n13850), .ZN(n13951) );
  INV_X1 U17008 ( .A(n13729), .ZN(n13933) );
  INV_X1 U17009 ( .A(n20075), .ZN(n14478) );
  AOI22_X1 U17010 ( .A1(n20070), .A2(n13933), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n14478), .ZN(n13730) );
  OAI21_X1 U17011 ( .B1(n13951), .B2(n14480), .A(n13730), .ZN(P1_U2871) );
  XNOR2_X1 U17012 ( .A(n19913), .B(n19915), .ZN(n13737) );
  XNOR2_X1 U17013 ( .A(n13732), .B(n13731), .ZN(n19927) );
  INV_X1 U17014 ( .A(n19927), .ZN(n13733) );
  NAND2_X1 U17015 ( .A1(n19903), .A2(n13733), .ZN(n13734) );
  OAI21_X1 U17016 ( .B1(n19903), .B2(n13733), .A(n13734), .ZN(n19133) );
  NOR2_X1 U17017 ( .A1(n19133), .A2(n19134), .ZN(n19132) );
  INV_X1 U17018 ( .A(n13734), .ZN(n13735) );
  NOR2_X1 U17019 ( .A1(n19132), .A2(n13735), .ZN(n13736) );
  NOR2_X1 U17020 ( .A1(n13736), .A2(n13737), .ZN(n13945) );
  AOI21_X1 U17021 ( .B1(n13737), .B2(n13736), .A(n13945), .ZN(n13741) );
  AOI22_X1 U17022 ( .A1(n19107), .A2(n16102), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19130), .ZN(n13740) );
  INV_X1 U17023 ( .A(n19915), .ZN(n13738) );
  NAND2_X1 U17024 ( .A1(n13738), .A2(n19131), .ZN(n13739) );
  OAI211_X1 U17025 ( .C1(n13741), .C2(n19135), .A(n13740), .B(n13739), .ZN(
        P2_U2917) );
  INV_X1 U17026 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20105) );
  INV_X1 U17027 ( .A(n13742), .ZN(n13743) );
  NAND2_X1 U17028 ( .A1(n14481), .A2(DATAI_0_), .ZN(n13745) );
  NAND2_X1 U17029 ( .A1(n14547), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13744) );
  AND2_X1 U17030 ( .A1(n13745), .A2(n13744), .ZN(n20214) );
  OAI222_X1 U17031 ( .A1(n14553), .A2(n13942), .B1(n14550), .B2(n20105), .C1(
        n14562), .C2(n20214), .ZN(P1_U2904) );
  INV_X1 U17032 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20100) );
  INV_X1 U17033 ( .A(DATAI_1_), .ZN(n20950) );
  NAND2_X1 U17034 ( .A1(n14481), .A2(n20950), .ZN(n13747) );
  INV_X1 U17035 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16458) );
  NAND2_X1 U17036 ( .A1(n14547), .A2(n16458), .ZN(n13746) );
  AND2_X1 U17037 ( .A1(n13747), .A2(n13746), .ZN(n20222) );
  INV_X1 U17038 ( .A(n20222), .ZN(n20118) );
  OAI222_X1 U17039 ( .A1(n13951), .A2(n14553), .B1(n14550), .B2(n20100), .C1(
        n14562), .C2(n20118), .ZN(P1_U2903) );
  INV_X1 U17040 ( .A(n13750), .ZN(n13751) );
  NAND2_X1 U17041 ( .A1(n13749), .A2(n13751), .ZN(n13753) );
  OAI21_X1 U17042 ( .B1(n13748), .B2(n13753), .A(n13752), .ZN(n19114) );
  OAI21_X1 U17043 ( .B1(n13755), .B2(n13754), .A(n13757), .ZN(n19175) );
  MUX2_X1 U17044 ( .A(n19175), .B(n14061), .S(n14987), .Z(n13756) );
  OAI21_X1 U17045 ( .B1(n19114), .B2(n15019), .A(n13756), .ZN(P2_U2883) );
  XOR2_X1 U17046 ( .A(n13752), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13761)
         );
  INV_X1 U17047 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13759) );
  AOI21_X1 U17048 ( .B1(n13758), .B2(n13757), .A(n13783), .ZN(n19048) );
  INV_X1 U17049 ( .A(n19048), .ZN(n15565) );
  MUX2_X1 U17050 ( .A(n13759), .B(n15565), .S(n15036), .Z(n13760) );
  OAI21_X1 U17051 ( .B1(n13761), .B2(n15019), .A(n13760), .ZN(P2_U2882) );
  XNOR2_X1 U17052 ( .A(n13762), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13768) );
  INV_X1 U17053 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13766) );
  INV_X1 U17054 ( .A(n13782), .ZN(n13764) );
  INV_X1 U17055 ( .A(n13857), .ZN(n13763) );
  OAI21_X1 U17056 ( .B1(n13765), .B2(n13764), .A(n13763), .ZN(n19037) );
  MUX2_X1 U17057 ( .A(n13766), .B(n19037), .S(n15036), .Z(n13767) );
  OAI21_X1 U17058 ( .B1(n13768), .B2(n15019), .A(n13767), .ZN(P2_U2880) );
  AND2_X1 U17059 ( .A1(n13770), .A2(n13769), .ZN(n13771) );
  OR2_X2 U17060 ( .A1(n13773), .A2(n13771), .ZN(n20147) );
  INV_X1 U17061 ( .A(n20150), .ZN(n20144) );
  AOI22_X1 U17062 ( .A1(n20144), .A2(n20140), .B1(P1_UWORD_REG_13__SCAN_IN), 
        .B2(n20147), .ZN(n13774) );
  OAI21_X1 U17063 ( .B1(n20148), .B2(n12612), .A(n13774), .ZN(P1_U2950) );
  INV_X1 U17064 ( .A(DATAI_11_), .ZN(n20947) );
  NAND2_X1 U17065 ( .A1(n14547), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13775) );
  OAI21_X1 U17066 ( .B1(n14547), .B2(n20947), .A(n13775), .ZN(n20135) );
  AOI22_X1 U17067 ( .A1(n20144), .A2(n20135), .B1(P1_UWORD_REG_11__SCAN_IN), 
        .B2(n20147), .ZN(n13776) );
  OAI21_X1 U17068 ( .B1(n20148), .B2(n14488), .A(n13776), .ZN(P1_U2948) );
  INV_X1 U17069 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13799) );
  INV_X1 U17070 ( .A(DATAI_14_), .ZN(n21024) );
  NAND2_X1 U17071 ( .A1(n14547), .A2(BUF1_REG_14__SCAN_IN), .ZN(n13777) );
  OAI21_X1 U17072 ( .B1(n14547), .B2(n21024), .A(n13777), .ZN(n20143) );
  AOI22_X1 U17073 ( .A1(n20144), .A2(n20143), .B1(P1_UWORD_REG_14__SCAN_IN), 
        .B2(n20147), .ZN(n13778) );
  OAI21_X1 U17074 ( .B1(n20148), .B2(n13799), .A(n13778), .ZN(P1_U2951) );
  INV_X1 U17075 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13795) );
  INV_X1 U17076 ( .A(DATAI_10_), .ZN(n13780) );
  NAND2_X1 U17077 ( .A1(n14547), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13779) );
  OAI21_X1 U17078 ( .B1(n14547), .B2(n13780), .A(n13779), .ZN(n20132) );
  AOI22_X1 U17079 ( .A1(n20144), .A2(n20132), .B1(P1_UWORD_REG_10__SCAN_IN), 
        .B2(n20147), .ZN(n13781) );
  OAI21_X1 U17080 ( .B1(n20148), .B2(n13795), .A(n13781), .ZN(P1_U2947) );
  OAI21_X1 U17081 ( .B1(n13784), .B2(n13783), .A(n13782), .ZN(n15551) );
  NOR2_X1 U17082 ( .A1(n13752), .A2(n10424), .ZN(n13786) );
  INV_X1 U17083 ( .A(n13762), .ZN(n13785) );
  OAI211_X1 U17084 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13786), .A(
        n13785), .B(n15041), .ZN(n13788) );
  NAND2_X1 U17085 ( .A1(n14987), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13787) );
  OAI211_X1 U17086 ( .C1(n15551), .C2(n14987), .A(n13788), .B(n13787), .ZN(
        P2_U2881) );
  INV_X1 U17087 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14539) );
  AOI22_X1 U17088 ( .A1(n20102), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n20101), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13789) );
  OAI21_X1 U17089 ( .B1(n14539), .B2(n13798), .A(n13789), .ZN(P1_U2920) );
  INV_X1 U17090 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20086) );
  INV_X1 U17091 ( .A(DATAI_9_), .ZN(n20968) );
  MUX2_X1 U17092 ( .A(n20968), .B(n16441), .S(n14547), .Z(n14498) );
  NOR2_X1 U17093 ( .A1(n20150), .A2(n14498), .ZN(n13792) );
  AOI21_X1 U17094 ( .B1(P1_LWORD_REG_9__SCAN_IN), .B2(n20147), .A(n13792), 
        .ZN(n13790) );
  OAI21_X1 U17095 ( .B1(n20086), .B2(n20148), .A(n13790), .ZN(P1_U2961) );
  AOI22_X1 U17096 ( .A1(n20102), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20101), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13791) );
  OAI21_X1 U17097 ( .B1(n14535), .B2(n13798), .A(n13791), .ZN(P1_U2919) );
  AOI21_X1 U17098 ( .B1(P1_UWORD_REG_9__SCAN_IN), .B2(n20147), .A(n13792), 
        .ZN(n13793) );
  OAI21_X1 U17099 ( .B1(n14497), .B2(n20148), .A(n13793), .ZN(P1_U2946) );
  AOI22_X1 U17100 ( .A1(n20872), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20101), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13794) );
  OAI21_X1 U17101 ( .B1(n13795), .B2(n13798), .A(n13794), .ZN(P1_U2910) );
  AOI22_X1 U17102 ( .A1(n20872), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20101), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13796) );
  OAI21_X1 U17103 ( .B1(n12612), .B2(n13798), .A(n13796), .ZN(P1_U2907) );
  AOI22_X1 U17104 ( .A1(n20872), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n20101), .ZN(n13797) );
  OAI21_X1 U17105 ( .B1(n13799), .B2(n13798), .A(n13797), .ZN(P1_U2906) );
  NAND2_X1 U17106 ( .A1(n20454), .A2(n13817), .ZN(n13820) );
  NAND2_X1 U17107 ( .A1(n13801), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13802) );
  NAND2_X1 U17108 ( .A1(n13803), .A2(n13802), .ZN(n20855) );
  NAND2_X1 U17109 ( .A1(n13804), .A2(n20855), .ZN(n13816) );
  XNOR2_X1 U17110 ( .A(n13805), .B(n13807), .ZN(n13814) );
  INV_X1 U17111 ( .A(n13806), .ZN(n13811) );
  NAND2_X1 U17112 ( .A1(n13808), .A2(n13807), .ZN(n13809) );
  OAI21_X1 U17113 ( .B1(n13811), .B2(n13810), .A(n13809), .ZN(n13812) );
  AOI22_X1 U17114 ( .A1(n15727), .A2(n13814), .B1(n13813), .B2(n13812), .ZN(
        n13815) );
  OAI21_X1 U17115 ( .B1(n13817), .B2(n13816), .A(n13815), .ZN(n13818) );
  INV_X1 U17116 ( .A(n13818), .ZN(n13819) );
  NAND2_X1 U17117 ( .A1(n13820), .A2(n13819), .ZN(n20858) );
  MUX2_X1 U17118 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20858), .S(
        n15725), .Z(n15739) );
  NAND2_X1 U17119 ( .A1(n15739), .A2(n16053), .ZN(n13823) );
  NAND2_X1 U17120 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n19983), .ZN(n13824) );
  INV_X1 U17121 ( .A(n13824), .ZN(n13821) );
  NAND2_X1 U17122 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13821), .ZN(
        n13822) );
  NAND2_X1 U17123 ( .A1(n13823), .A2(n13822), .ZN(n13829) );
  NAND2_X1 U17124 ( .A1(n13824), .A2(n15725), .ZN(n13826) );
  NAND2_X1 U17125 ( .A1(n15725), .A2(n16053), .ZN(n13831) );
  INV_X1 U17126 ( .A(n13831), .ZN(n13825) );
  OAI22_X1 U17127 ( .A1(n15726), .A2(n13826), .B1(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n13825), .ZN(n13827) );
  INV_X1 U17128 ( .A(n13827), .ZN(n13828) );
  NAND2_X1 U17129 ( .A1(n13829), .A2(n13828), .ZN(n15748) );
  AOI21_X1 U17130 ( .B1(n14423), .B2(n13830), .A(n13831), .ZN(n13835) );
  NAND2_X1 U17131 ( .A1(n12327), .A2(n13831), .ZN(n13833) );
  NAND2_X1 U17132 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_FLUSH_REG_SCAN_IN), 
        .ZN(n13832) );
  NAND2_X1 U17133 ( .A1(n13833), .A2(n13832), .ZN(n13834) );
  OR2_X1 U17134 ( .A1(n13835), .A2(n13834), .ZN(n15745) );
  OAI21_X1 U17135 ( .B1(n15748), .B2(n11513), .A(n15745), .ZN(n13844) );
  NOR2_X1 U17136 ( .A1(n16055), .A2(n16054), .ZN(n13836) );
  OAI21_X1 U17137 ( .B1(n13844), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13836), .ZN(
        n13839) );
  INV_X1 U17138 ( .A(n16054), .ZN(n13838) );
  NAND2_X1 U17139 ( .A1(n13839), .A2(n20353), .ZN(n20209) );
  INV_X1 U17140 ( .A(n13869), .ZN(n13840) );
  NOR2_X1 U17141 ( .A1(n20283), .A2(n13840), .ZN(n13867) );
  NOR2_X1 U17142 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20719), .ZN(n13870) );
  NAND2_X1 U17143 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20590), .ZN(n13845) );
  AOI22_X1 U17144 ( .A1(n20283), .A2(n13870), .B1(n20674), .B2(n13845), .ZN(
        n13841) );
  INV_X1 U17145 ( .A(n13841), .ZN(n13842) );
  OAI21_X1 U17146 ( .B1(n13867), .B2(n13842), .A(n20209), .ZN(n13843) );
  OAI21_X1 U17147 ( .B1(n20209), .B2(n20582), .A(n13843), .ZN(P1_U3477) );
  NOR2_X1 U17148 ( .A1(n13844), .A2(n16054), .ZN(n15760) );
  INV_X1 U17149 ( .A(n13845), .ZN(n14817) );
  OAI22_X1 U17150 ( .A1(n12509), .A2(n20719), .B1(n13846), .B2(n14817), .ZN(
        n13847) );
  OAI21_X1 U17151 ( .B1(n15760), .B2(n13847), .A(n20209), .ZN(n13848) );
  OAI21_X1 U17152 ( .B1(n20209), .B2(n20634), .A(n13848), .ZN(P1_U3478) );
  OAI21_X1 U17153 ( .B1(n11810), .B2(n11809), .A(n13851), .ZN(n13978) );
  AND2_X1 U17154 ( .A1(n13889), .A2(n13853), .ZN(n20183) );
  AOI22_X1 U17155 ( .A1(n20070), .A2(n20183), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n14478), .ZN(n13854) );
  OAI21_X1 U17156 ( .B1(n13978), .B2(n14480), .A(n13854), .ZN(P1_U2870) );
  INV_X1 U17157 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20098) );
  NAND2_X1 U17158 ( .A1(n14481), .A2(DATAI_2_), .ZN(n13856) );
  NAND2_X1 U17159 ( .A1(n14547), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13855) );
  AND2_X1 U17160 ( .A1(n13856), .A2(n13855), .ZN(n20120) );
  OAI222_X1 U17161 ( .A1(n14553), .A2(n13978), .B1(n14550), .B2(n20098), .C1(
        n14562), .C2(n20120), .ZN(P1_U2902) );
  OR2_X1 U17162 ( .A1(n13858), .A2(n13857), .ZN(n13859) );
  NAND2_X1 U17163 ( .A1(n13859), .A2(n13880), .ZN(n16280) );
  INV_X1 U17164 ( .A(n13860), .ZN(n13863) );
  OAI211_X1 U17165 ( .C1(n13863), .C2(n13862), .A(n15041), .B(n13861), .ZN(
        n13865) );
  NAND2_X1 U17166 ( .A1(n14987), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13864) );
  OAI211_X1 U17167 ( .C1(n16280), .C2(n14987), .A(n13865), .B(n13864), .ZN(
        P2_U2879) );
  NOR2_X1 U17168 ( .A1(n20554), .A2(n20719), .ZN(n13873) );
  NAND2_X1 U17169 ( .A1(n12521), .A2(n13866), .ZN(n20716) );
  INV_X1 U17170 ( .A(n13867), .ZN(n20260) );
  NOR2_X1 U17171 ( .A1(n20716), .A2(n20260), .ZN(n20639) );
  NAND2_X1 U17172 ( .A1(n20283), .A2(n13869), .ZN(n20551) );
  NOR2_X1 U17173 ( .A1(n20426), .A2(n20551), .ZN(n20432) );
  INV_X1 U17174 ( .A(n13870), .ZN(n20577) );
  INV_X1 U17175 ( .A(n20454), .ZN(n13871) );
  OAI22_X1 U17176 ( .A1(n14089), .A2(n20577), .B1(n13871), .B2(n14817), .ZN(
        n13872) );
  NOR4_X1 U17177 ( .A1(n13873), .A2(n20639), .A3(n20432), .A4(n13872), .ZN(
        n13876) );
  INV_X1 U17178 ( .A(n20209), .ZN(n13875) );
  NAND2_X1 U17179 ( .A1(n13875), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13874) );
  OAI21_X1 U17180 ( .B1(n13876), .B2(n13875), .A(n13874), .ZN(P1_U3475) );
  INV_X1 U17181 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n19016) );
  INV_X1 U17182 ( .A(n13861), .ZN(n13879) );
  INV_X1 U17183 ( .A(n9773), .ZN(n13877) );
  OAI211_X1 U17184 ( .C1(n13879), .C2(n13878), .A(n13877), .B(n15041), .ZN(
        n13883) );
  AOI21_X1 U17185 ( .B1(n13881), .B2(n13880), .A(n13901), .ZN(n19024) );
  NAND2_X1 U17186 ( .A1(n19024), .A2(n15036), .ZN(n13882) );
  OAI211_X1 U17187 ( .C1(n15036), .C2(n19016), .A(n13883), .B(n13882), .ZN(
        P2_U2878) );
  OAI21_X1 U17188 ( .B1(n13884), .B2(n13885), .A(n13963), .ZN(n14161) );
  INV_X1 U17189 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20096) );
  NAND2_X1 U17190 ( .A1(n14481), .A2(DATAI_3_), .ZN(n13887) );
  NAND2_X1 U17191 ( .A1(n14547), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13886) );
  AND2_X1 U17192 ( .A1(n13887), .A2(n13886), .ZN(n20228) );
  OAI222_X1 U17193 ( .A1(n14553), .A2(n14161), .B1(n14550), .B2(n20096), .C1(
        n14562), .C2(n20228), .ZN(P1_U2901) );
  AND2_X1 U17194 ( .A1(n13889), .A2(n13888), .ZN(n13890) );
  NOR2_X1 U17195 ( .A1(n13910), .A2(n13890), .ZN(n20174) );
  INV_X1 U17196 ( .A(n20174), .ZN(n13891) );
  INV_X1 U17197 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n14035) );
  OAI222_X1 U17198 ( .A1(n13891), .A2(n14467), .B1(n14035), .B2(n20075), .C1(
        n14161), .C2(n14480), .ZN(P1_U2869) );
  OAI21_X1 U17199 ( .B1(n13894), .B2(n13893), .A(n13892), .ZN(n20186) );
  INV_X1 U17200 ( .A(n13978), .ZN(n13897) );
  INV_X2 U17201 ( .A(n20170), .ZN(n20190) );
  AOI22_X1 U17202 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20190), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13895) );
  OAI21_X1 U17203 ( .B1(n20161), .B2(n13967), .A(n13895), .ZN(n13896) );
  AOI21_X1 U17204 ( .B1(n13897), .B2(n20167), .A(n13896), .ZN(n13898) );
  OAI21_X1 U17205 ( .B1(n20172), .B2(n20186), .A(n13898), .ZN(P1_U2997) );
  OAI211_X1 U17206 ( .C1(n9773), .C2(n13900), .A(n13899), .B(n15041), .ZN(
        n13905) );
  NOR2_X1 U17207 ( .A1(n13902), .A2(n13901), .ZN(n13903) );
  OR2_X1 U17208 ( .A1(n13921), .A2(n13903), .ZN(n14146) );
  INV_X1 U17209 ( .A(n14146), .ZN(n16272) );
  NAND2_X1 U17210 ( .A1(n15036), .A2(n16272), .ZN(n13904) );
  OAI211_X1 U17211 ( .C1(n15036), .C2(n14142), .A(n13905), .B(n13904), .ZN(
        P2_U2877) );
  OAI21_X1 U17212 ( .B1(n13908), .B2(n13907), .A(n13906), .ZN(n20153) );
  OAI21_X1 U17213 ( .B1(n13910), .B2(n13909), .A(n16040), .ZN(n14420) );
  NOR2_X1 U17214 ( .A1(n16014), .A2(n14420), .ZN(n13918) );
  NOR2_X1 U17215 ( .A1(n13915), .A2(n20179), .ZN(n16046) );
  OAI21_X1 U17216 ( .B1(n20198), .B2(n13911), .A(n20191), .ZN(n20181) );
  INV_X1 U17217 ( .A(n20181), .ZN(n13914) );
  NOR2_X1 U17218 ( .A1(n20191), .A2(n13911), .ZN(n14708) );
  OAI21_X1 U17219 ( .B1(n14716), .B2(n20198), .A(n20199), .ZN(n20192) );
  AOI21_X1 U17220 ( .B1(n14708), .B2(n20192), .A(n20185), .ZN(n15975) );
  NOR2_X1 U17221 ( .A1(n13914), .A2(n15975), .ZN(n20176) );
  OAI21_X1 U17222 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20176), .ZN(n13916) );
  NAND2_X1 U17223 ( .A1(n20199), .A2(n14716), .ZN(n15976) );
  INV_X1 U17224 ( .A(n15976), .ZN(n15998) );
  INV_X1 U17225 ( .A(n14716), .ZN(n13912) );
  NAND2_X1 U17226 ( .A1(n13912), .A2(n20198), .ZN(n13913) );
  OAI21_X1 U17227 ( .B1(n15998), .B2(n14708), .A(n15980), .ZN(n20187) );
  AOI21_X1 U17228 ( .B1(n20185), .B2(n13914), .A(n20187), .ZN(n20180) );
  OAI22_X1 U17229 ( .A1(n16046), .A2(n13916), .B1(n20180), .B2(n13915), .ZN(
        n13917) );
  AOI211_X1 U17230 ( .C1(n20190), .C2(P1_REIP_REG_4__SCAN_IN), .A(n13918), .B(
        n13917), .ZN(n13919) );
  OAI21_X1 U17231 ( .B1(n20208), .B2(n20153), .A(n13919), .ZN(P1_U3027) );
  XNOR2_X1 U17232 ( .A(n13899), .B(n14024), .ZN(n13924) );
  NOR2_X1 U17233 ( .A1(n13921), .A2(n13920), .ZN(n13922) );
  OR2_X1 U17234 ( .A1(n14021), .A2(n13922), .ZN(n16261) );
  MUX2_X1 U17235 ( .A(n19005), .B(n16261), .S(n15036), .Z(n13923) );
  OAI21_X1 U17236 ( .B1(n13924), .B2(n15019), .A(n13923), .ZN(P2_U2876) );
  INV_X1 U17237 ( .A(n13928), .ZN(n13925) );
  NAND2_X1 U17238 ( .A1(n13925), .A2(n11607), .ZN(n13926) );
  NAND2_X1 U17239 ( .A1(n13926), .A2(n14414), .ZN(n20046) );
  AOI22_X1 U17240 ( .A1(n13342), .A2(n14407), .B1(n15848), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13935) );
  INV_X1 U17241 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13931) );
  NOR2_X1 U17242 ( .A1(n13928), .A2(n13927), .ZN(n14422) );
  NAND2_X1 U17243 ( .A1(n14422), .A2(n20674), .ZN(n13930) );
  INV_X1 U17244 ( .A(n14217), .ZN(n13972) );
  AOI22_X1 U17245 ( .A1(n20027), .A2(n13931), .B1(n13972), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n13929) );
  OAI211_X1 U17246 ( .C1(n20000), .C2(n13931), .A(n13930), .B(n13929), .ZN(
        n13932) );
  AOI21_X1 U17247 ( .B1(n20047), .B2(n13933), .A(n13932), .ZN(n13934) );
  OAI211_X1 U17248 ( .C1(n13951), .C2(n14040), .A(n13935), .B(n13934), .ZN(
        P1_U2839) );
  NAND2_X1 U17249 ( .A1(n14422), .A2(n9664), .ZN(n13937) );
  OAI21_X1 U17250 ( .B1(n20048), .B2(n20027), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13936) );
  OAI211_X1 U17251 ( .C1(n20054), .C2(n13938), .A(n13937), .B(n13936), .ZN(
        n13939) );
  AOI21_X1 U17252 ( .B1(n20047), .B2(n20204), .A(n13939), .ZN(n13941) );
  NAND2_X1 U17253 ( .A1(n20021), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13940) );
  OAI211_X1 U17254 ( .C1(n13942), .C2(n14040), .A(n13941), .B(n13940), .ZN(
        P1_U2840) );
  XNOR2_X1 U17255 ( .A(n13944), .B(n13943), .ZN(n19898) );
  AOI21_X1 U17256 ( .B1(n19915), .B2(n19913), .A(n13945), .ZN(n19125) );
  XNOR2_X1 U17257 ( .A(n19898), .B(n19904), .ZN(n19126) );
  NOR2_X1 U17258 ( .A1(n19125), .A2(n19126), .ZN(n19124) );
  AOI21_X1 U17259 ( .B1(n19898), .B2(n19904), .A(n19124), .ZN(n13947) );
  XNOR2_X1 U17260 ( .A(n13946), .B(n9776), .ZN(n14058) );
  NOR2_X1 U17261 ( .A1(n13947), .A2(n14058), .ZN(n19115) );
  XNOR2_X1 U17262 ( .A(n19115), .B(n19114), .ZN(n13950) );
  AOI22_X1 U17263 ( .A1(n19131), .A2(n14058), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19130), .ZN(n13949) );
  NAND2_X1 U17264 ( .A1(n19107), .A2(n16095), .ZN(n13948) );
  OAI211_X1 U17265 ( .C1(n13950), .C2(n19135), .A(n13949), .B(n13948), .ZN(
        P2_U2915) );
  INV_X1 U17266 ( .A(n13951), .ZN(n13959) );
  INV_X1 U17267 ( .A(n13952), .ZN(n13953) );
  AOI21_X1 U17268 ( .B1(n20152), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13953), .ZN(n13954) );
  OAI21_X1 U17269 ( .B1(n20161), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13954), .ZN(n13958) );
  NOR3_X1 U17270 ( .A1(n13956), .A2(n13955), .A3(n20172), .ZN(n13957) );
  AOI211_X1 U17271 ( .C1(n20154), .C2(n13959), .A(n13958), .B(n13957), .ZN(
        n13960) );
  INV_X1 U17272 ( .A(n13960), .ZN(P1_U2998) );
  INV_X1 U17273 ( .A(DATAI_4_), .ZN(n20923) );
  NAND2_X1 U17274 ( .A1(n14481), .A2(n20923), .ZN(n13962) );
  NAND2_X1 U17275 ( .A1(n14547), .A2(n16452), .ZN(n13961) );
  AND2_X1 U17276 ( .A1(n13962), .A2(n13961), .ZN(n14826) );
  INV_X1 U17277 ( .A(n14826), .ZN(n20123) );
  INV_X1 U17278 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20094) );
  XOR2_X1 U17279 ( .A(n13964), .B(n13963), .Z(n20155) );
  INV_X1 U17280 ( .A(n20155), .ZN(n13965) );
  OAI222_X1 U17281 ( .A1(n20123), .A2(n14562), .B1(n14550), .B2(n20094), .C1(
        n14553), .C2(n13965), .ZN(P1_U2900) );
  INV_X1 U17282 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13966) );
  OAI222_X1 U17283 ( .A1(n14420), .A2(n14467), .B1(n20075), .B2(n13966), .C1(
        n14480), .C2(n13965), .ZN(P1_U2868) );
  INV_X1 U17284 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13971) );
  NAND2_X1 U17285 ( .A1(n20047), .A2(n20183), .ZN(n13970) );
  INV_X1 U17286 ( .A(n13967), .ZN(n13968) );
  AOI22_X1 U17287 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n20048), .B1(
        n20027), .B2(n13968), .ZN(n13969) );
  OAI211_X1 U17288 ( .C1(n13971), .C2(n20054), .A(n13970), .B(n13969), .ZN(
        n13976) );
  NAND2_X1 U17289 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n13973) );
  AOI21_X1 U17290 ( .B1(n14407), .B2(n13973), .A(n13972), .ZN(n14036) );
  AOI21_X1 U17291 ( .B1(n14407), .B2(P1_REIP_REG_1__SCAN_IN), .A(
        P1_REIP_REG_2__SCAN_IN), .ZN(n13974) );
  NOR2_X1 U17292 ( .A1(n14036), .A2(n13974), .ZN(n13975) );
  AOI211_X1 U17293 ( .C1(n14422), .C2(n14092), .A(n13976), .B(n13975), .ZN(
        n13977) );
  OAI21_X1 U17294 ( .B1(n14040), .B2(n13978), .A(n13977), .ZN(P1_U2838) );
  OR2_X1 U17295 ( .A1(n13981), .A2(n13980), .ZN(n13982) );
  AND2_X1 U17296 ( .A1(n13979), .A2(n13982), .ZN(n20072) );
  INV_X1 U17297 ( .A(n20072), .ZN(n13985) );
  INV_X1 U17298 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20092) );
  INV_X1 U17299 ( .A(DATAI_5_), .ZN(n13984) );
  NAND2_X1 U17300 ( .A1(n14547), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13983) );
  OAI21_X1 U17301 ( .B1(n14547), .B2(n13984), .A(n13983), .ZN(n20237) );
  INV_X1 U17302 ( .A(n20237), .ZN(n20125) );
  OAI222_X1 U17303 ( .A1(n14553), .A2(n13985), .B1(n14550), .B2(n20092), .C1(
        n14562), .C2(n20125), .ZN(P1_U2899) );
  NOR2_X1 U17304 ( .A1(n18993), .A2(n13986), .ZN(n13987) );
  XNOR2_X1 U17305 ( .A(n13987), .B(n15272), .ZN(n13990) );
  XNOR2_X1 U17306 ( .A(n13989), .B(n13988), .ZN(n15550) );
  AOI22_X1 U17307 ( .A1(n19049), .A2(n13990), .B1(n19056), .B2(n15550), .ZN(
        n13997) );
  INV_X1 U17308 ( .A(n15551), .ZN(n13995) );
  INV_X1 U17309 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13993) );
  OAI21_X1 U17310 ( .B1(n19846), .B2(n19035), .A(n19033), .ZN(n13991) );
  AOI21_X1 U17311 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19068), .A(
        n13991), .ZN(n13992) );
  OAI21_X1 U17312 ( .B1(n19017), .B2(n13993), .A(n13992), .ZN(n13994) );
  AOI21_X1 U17313 ( .B1(n13995), .B2(n19062), .A(n13994), .ZN(n13996) );
  OAI211_X1 U17314 ( .C1(n13998), .C2(n9646), .A(n13997), .B(n13996), .ZN(
        P2_U2849) );
  XNOR2_X1 U17315 ( .A(n13999), .B(n14014), .ZN(n14001) );
  XNOR2_X1 U17316 ( .A(n14001), .B(n14000), .ZN(n19178) );
  INV_X1 U17317 ( .A(n19178), .ZN(n14019) );
  XOR2_X1 U17318 ( .A(n14003), .B(n14002), .Z(n19176) );
  INV_X1 U17319 ( .A(n14004), .ZN(n14006) );
  NAND2_X1 U17320 ( .A1(n14006), .A2(n14005), .ZN(n14007) );
  INV_X1 U17321 ( .A(n16257), .ZN(n16277) );
  NOR3_X1 U17322 ( .A1(n14008), .A2(n14007), .A3(n10175), .ZN(n16312) );
  NOR2_X1 U17323 ( .A1(n16277), .A2(n16312), .ZN(n15573) );
  NOR3_X1 U17324 ( .A1(n15456), .A2(n14010), .A3(n14009), .ZN(n14011) );
  OAI22_X1 U17325 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19216), .B1(
        n14012), .B2(n14011), .ZN(n16311) );
  NOR2_X1 U17326 ( .A1(n10175), .A2(n16311), .ZN(n15560) );
  NOR2_X1 U17327 ( .A1(n12677), .A2(n19033), .ZN(n14013) );
  AOI221_X1 U17328 ( .B1(n15573), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(
        n15560), .C2(n14014), .A(n14013), .ZN(n14016) );
  NAND2_X1 U17329 ( .A1(n19202), .A2(n14058), .ZN(n14015) );
  OAI211_X1 U17330 ( .C1(n19175), .C2(n19206), .A(n14016), .B(n14015), .ZN(
        n14017) );
  AOI21_X1 U17331 ( .B1(n19176), .B2(n16309), .A(n14017), .ZN(n14018) );
  OAI21_X1 U17332 ( .B1(n14019), .B2(n16301), .A(n14018), .ZN(P2_U3042) );
  OAI21_X1 U17333 ( .B1(n14021), .B2(n14020), .A(n14169), .ZN(n16248) );
  OAI21_X1 U17334 ( .B1(n13899), .B2(n14024), .A(n14023), .ZN(n14025) );
  NAND3_X1 U17335 ( .A1(n14022), .A2(n15041), .A3(n14025), .ZN(n14027) );
  NAND2_X1 U17336 ( .A1(n14987), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14026) );
  OAI211_X1 U17337 ( .C1(n16248), .C2(n14987), .A(n14027), .B(n14026), .ZN(
        P2_U2875) );
  NAND2_X1 U17338 ( .A1(n20047), .A2(n20174), .ZN(n14034) );
  NAND3_X1 U17339 ( .A1(n14407), .A2(P1_REIP_REG_1__SCAN_IN), .A3(
        P1_REIP_REG_2__SCAN_IN), .ZN(n14031) );
  NAND2_X1 U17340 ( .A1(n20048), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14030) );
  INV_X1 U17341 ( .A(n14157), .ZN(n14028) );
  NAND2_X1 U17342 ( .A1(n20027), .A2(n14028), .ZN(n14029) );
  OAI211_X1 U17343 ( .C1(P1_REIP_REG_3__SCAN_IN), .C2(n14031), .A(n14030), .B(
        n14029), .ZN(n14032) );
  INV_X1 U17344 ( .A(n14032), .ZN(n14033) );
  OAI211_X1 U17345 ( .C1(n14035), .C2(n20054), .A(n14034), .B(n14033), .ZN(
        n14038) );
  INV_X1 U17346 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20792) );
  NOR2_X1 U17347 ( .A1(n14036), .A2(n20792), .ZN(n14037) );
  AOI211_X1 U17348 ( .C1(n14422), .C2(n20454), .A(n14038), .B(n14037), .ZN(
        n14039) );
  OAI21_X1 U17349 ( .B1(n14040), .B2(n14161), .A(n14039), .ZN(P1_U2837) );
  INV_X1 U17350 ( .A(n14076), .ZN(n19065) );
  NOR2_X1 U17351 ( .A1(n18993), .A2(n14067), .ZN(n14042) );
  XNOR2_X1 U17352 ( .A(n14042), .B(n14041), .ZN(n14043) );
  NAND2_X1 U17353 ( .A1(n14043), .A2(n19049), .ZN(n14051) );
  OAI22_X1 U17354 ( .A1(n19017), .A2(n14044), .B1(n19915), .B2(n19053), .ZN(
        n14046) );
  NOR2_X1 U17355 ( .A1(n19035), .A2(n19841), .ZN(n14045) );
  AOI211_X1 U17356 ( .C1(n19068), .C2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n14046), .B(n14045), .ZN(n14047) );
  OAI21_X1 U17357 ( .B1(n14048), .B2(n9646), .A(n14047), .ZN(n14049) );
  AOI21_X1 U17358 ( .B1(n10688), .B2(n19062), .A(n14049), .ZN(n14050) );
  OAI211_X1 U17359 ( .C1(n19065), .C2(n19913), .A(n14051), .B(n14050), .ZN(
        P2_U2853) );
  INV_X1 U17360 ( .A(n19181), .ZN(n14055) );
  NOR2_X1 U17361 ( .A1(n18993), .A2(n14052), .ZN(n14054) );
  AOI21_X1 U17362 ( .B1(n14055), .B2(n14054), .A(n19822), .ZN(n14053) );
  OAI21_X1 U17363 ( .B1(n14055), .B2(n14054), .A(n14053), .ZN(n14066) );
  INV_X1 U17364 ( .A(n14056), .ZN(n14064) );
  NOR2_X1 U17365 ( .A1(n19035), .A2(n12677), .ZN(n14057) );
  AOI211_X1 U17366 ( .C1(n19068), .C2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n19192), .B(n14057), .ZN(n14060) );
  NAND2_X1 U17367 ( .A1(n19056), .A2(n14058), .ZN(n14059) );
  OAI211_X1 U17368 ( .C1(n14061), .C2(n19017), .A(n14060), .B(n14059), .ZN(
        n14063) );
  NOR2_X1 U17369 ( .A1(n19175), .A2(n19036), .ZN(n14062) );
  AOI211_X1 U17370 ( .C1(n19031), .C2(n14064), .A(n14063), .B(n14062), .ZN(
        n14065) );
  OAI211_X1 U17371 ( .C1(n19065), .C2(n19114), .A(n14066), .B(n14065), .ZN(
        P2_U2851) );
  INV_X1 U17372 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14073) );
  AOI211_X1 U17373 ( .C1(n14187), .C2(n14068), .A(n18993), .B(n14067), .ZN(
        n14186) );
  AOI21_X1 U17374 ( .B1(n18993), .B2(n14073), .A(n14186), .ZN(n14078) );
  INV_X1 U17375 ( .A(n19184), .ZN(n14069) );
  OAI22_X1 U17376 ( .A1(n19017), .A2(n14070), .B1(n14069), .B2(n9646), .ZN(
        n14071) );
  AOI21_X1 U17377 ( .B1(n19056), .B2(n19927), .A(n14071), .ZN(n14072) );
  OAI21_X1 U17378 ( .B1(n19207), .B2(n19036), .A(n14072), .ZN(n14075) );
  OAI22_X1 U17379 ( .A1(n14073), .A2(n19006), .B1(n10595), .B2(n19035), .ZN(
        n14074) );
  AOI211_X1 U17380 ( .C1(n14076), .C2(n19923), .A(n14075), .B(n14074), .ZN(
        n14077) );
  OAI21_X1 U17381 ( .B1(n14078), .B2(n19822), .A(n14077), .ZN(P2_U2854) );
  NAND2_X1 U17382 ( .A1(n14079), .A2(n14080), .ZN(n14081) );
  XNOR2_X1 U17383 ( .A(n16215), .B(n14081), .ZN(n14082) );
  NAND2_X1 U17384 ( .A1(n14082), .A2(n19049), .ZN(n14087) );
  INV_X1 U17385 ( .A(n14083), .ZN(n16220) );
  AOI22_X1 U17386 ( .A1(n19055), .A2(P2_EBX_REG_3__SCAN_IN), .B1(n19054), .B2(
        P2_REIP_REG_3__SCAN_IN), .ZN(n14084) );
  OAI21_X1 U17387 ( .B1(n16220), .B2(n9646), .A(n14084), .ZN(n14086) );
  OAI22_X1 U17388 ( .A1(n12656), .A2(n19006), .B1(n19053), .B2(n19898), .ZN(
        n14085) );
  OAI211_X1 U17389 ( .C1(n19904), .C2(n19065), .A(n14087), .B(n9783), .ZN(
        P2_U2852) );
  XOR2_X1 U17390 ( .A(n13979), .B(n14125), .Z(n20042) );
  INV_X1 U17391 ( .A(n20042), .ZN(n14133) );
  XNOR2_X1 U17392 ( .A(n16042), .B(n16021), .ZN(n20035) );
  AOI22_X1 U17393 ( .A1(n20070), .A2(n20035), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14478), .ZN(n14088) );
  OAI21_X1 U17394 ( .B1(n14133), .B2(n14480), .A(n14088), .ZN(P1_U2866) );
  INV_X1 U17395 ( .A(n12521), .ZN(n14816) );
  OAI21_X1 U17396 ( .B1(n20279), .B2(n20759), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14091) );
  NAND2_X1 U17397 ( .A1(n14091), .A2(n20721), .ZN(n14101) );
  OR2_X1 U17398 ( .A1(n20454), .A2(n14092), .ZN(n20318) );
  OR2_X1 U17399 ( .A1(n20318), .A2(n20674), .ZN(n14096) );
  INV_X1 U17400 ( .A(n20456), .ZN(n14093) );
  NAND2_X1 U17401 ( .A1(n14093), .A2(n20512), .ZN(n20349) );
  NOR2_X1 U17402 ( .A1(n14097), .A2(n11773), .ZN(n20514) );
  INV_X1 U17403 ( .A(n20514), .ZN(n20457) );
  OAI22_X1 U17404 ( .A1(n14101), .A2(n14096), .B1(n20349), .B2(n20457), .ZN(
        n20250) );
  INV_X1 U17405 ( .A(DATAI_7_), .ZN(n14095) );
  NAND2_X1 U17406 ( .A1(n14547), .A2(BUF1_REG_7__SCAN_IN), .ZN(n14094) );
  OAI21_X1 U17407 ( .B1(n14547), .B2(n14095), .A(n14094), .ZN(n14129) );
  NAND2_X1 U17408 ( .A1(n20261), .A2(n14129), .ZN(n20632) );
  INV_X1 U17409 ( .A(n20632), .ZN(n20764) );
  INV_X1 U17410 ( .A(n14096), .ZN(n14100) );
  NAND3_X1 U17411 ( .A1(n20546), .A2(n12312), .A3(n20582), .ZN(n20259) );
  NOR2_X1 U17412 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20259), .ZN(
        n20236) );
  INV_X1 U17413 ( .A(n20236), .ZN(n20244) );
  NAND2_X1 U17414 ( .A1(n14097), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20672) );
  NAND2_X1 U17415 ( .A1(n20261), .A2(n20672), .ZN(n20458) );
  AOI21_X1 U17416 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20244), .A(n20458), 
        .ZN(n14099) );
  NAND2_X1 U17417 ( .A1(n20349), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14098) );
  OAI211_X1 U17418 ( .C1(n14101), .C2(n14100), .A(n14099), .B(n14098), .ZN(
        n14825) );
  INV_X1 U17419 ( .A(DATAI_23_), .ZN(n14102) );
  INV_X1 U17420 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16419) );
  OAI22_X1 U17421 ( .A1(n14102), .A2(n20247), .B1(n16419), .B2(n20248), .ZN(
        n20664) );
  NOR2_X2 U17422 ( .A1(n20235), .A2(n14104), .ZN(n20767) );
  AOI22_X1 U17423 ( .A1(n20279), .A2(n20664), .B1(n20236), .B2(n20767), .ZN(
        n14106) );
  INV_X1 U17424 ( .A(DATAI_31_), .ZN(n21000) );
  OAI22_X2 U17425 ( .A1(n21000), .A2(n20247), .B1(n16409), .B2(n20248), .ZN(
        n20768) );
  NAND2_X1 U17426 ( .A1(n20759), .A2(n20768), .ZN(n14105) );
  OAI211_X1 U17427 ( .C1(n20254), .C2(n14107), .A(n14106), .B(n14105), .ZN(
        n14108) );
  AOI21_X1 U17428 ( .B1(n20250), .B2(n20764), .A(n14108), .ZN(n14109) );
  INV_X1 U17429 ( .A(n14109), .ZN(P1_U3040) );
  INV_X1 U17430 ( .A(n14110), .ZN(n14123) );
  NOR2_X1 U17431 ( .A1(n18993), .A2(n14111), .ZN(n14112) );
  XNOR2_X1 U17432 ( .A(n14112), .B(n16206), .ZN(n14115) );
  AOI21_X1 U17433 ( .B1(n14114), .B2(n16289), .A(n14113), .ZN(n19106) );
  AOI22_X1 U17434 ( .A1(n19049), .A2(n14115), .B1(n19056), .B2(n19106), .ZN(
        n14122) );
  INV_X1 U17435 ( .A(n16280), .ZN(n14120) );
  AOI21_X1 U17436 ( .B1(n18996), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n19192), .ZN(n14117) );
  NAND2_X1 U17437 ( .A1(n19054), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n14116) );
  OAI211_X1 U17438 ( .C1(n19017), .C2(n14118), .A(n14117), .B(n14116), .ZN(
        n14119) );
  AOI21_X1 U17439 ( .B1(n19062), .B2(n14120), .A(n14119), .ZN(n14121) );
  OAI211_X1 U17440 ( .C1(n14123), .C2(n9646), .A(n14122), .B(n14121), .ZN(
        P2_U2847) );
  OR2_X1 U17441 ( .A1(n13979), .A2(n14125), .ZN(n14127) );
  NAND2_X1 U17442 ( .A1(n14127), .A2(n14126), .ZN(n14128) );
  AND2_X1 U17443 ( .A1(n14124), .A2(n14128), .ZN(n20066) );
  INV_X1 U17444 ( .A(n20066), .ZN(n14130) );
  INV_X1 U17445 ( .A(n14129), .ZN(n20128) );
  OAI222_X1 U17446 ( .A1(n14553), .A2(n14130), .B1(n14550), .B2(n11779), .C1(
        n14562), .C2(n20128), .ZN(P1_U2897) );
  NAND2_X1 U17447 ( .A1(n14481), .A2(DATAI_6_), .ZN(n14132) );
  NAND2_X1 U17448 ( .A1(n14547), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14131) );
  AND2_X1 U17449 ( .A1(n14132), .A2(n14131), .ZN(n20246) );
  OAI222_X1 U17450 ( .A1(n14562), .A2(n20246), .B1(n14553), .B2(n14133), .C1(
        n11784), .C2(n14550), .ZN(P1_U2898) );
  AOI21_X1 U17451 ( .B1(n14134), .B2(n15538), .A(n16256), .ZN(n19100) );
  NOR2_X1 U17452 ( .A1(n18993), .A2(n14135), .ZN(n14136) );
  XNOR2_X1 U17453 ( .A(n14136), .B(n16185), .ZN(n14137) );
  AOI22_X1 U17454 ( .A1(n19100), .A2(n19056), .B1(n19049), .B2(n14137), .ZN(
        n14145) );
  INV_X1 U17455 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n14138) );
  OAI22_X1 U17456 ( .A1(n14139), .A2(n9646), .B1(n19006), .B2(n14138), .ZN(
        n14140) );
  INV_X1 U17457 ( .A(n14140), .ZN(n14141) );
  OAI21_X1 U17458 ( .B1(n19017), .B2(n14142), .A(n14141), .ZN(n14143) );
  AOI211_X1 U17459 ( .C1(n19054), .C2(P2_REIP_REG_10__SCAN_IN), .A(n19192), 
        .B(n14143), .ZN(n14144) );
  OAI211_X1 U17460 ( .C1(n19036), .C2(n14146), .A(n14145), .B(n14144), .ZN(
        P2_U2845) );
  AND2_X1 U17461 ( .A1(n14124), .A2(n14147), .ZN(n14149) );
  OR2_X1 U17462 ( .A1(n14149), .A2(n14148), .ZN(n14203) );
  INV_X1 U17463 ( .A(n16011), .ZN(n14152) );
  NAND2_X1 U17464 ( .A1(n16026), .A2(n14150), .ZN(n14151) );
  NAND2_X1 U17465 ( .A1(n14152), .A2(n14151), .ZN(n20013) );
  OAI222_X1 U17466 ( .A1(n14203), .A2(n14480), .B1(n20075), .B2(n20010), .C1(
        n20013), .C2(n14467), .ZN(P1_U2864) );
  OAI21_X1 U17467 ( .B1(n14155), .B2(n14154), .A(n14153), .ZN(n14156) );
  INV_X1 U17468 ( .A(n14156), .ZN(n20175) );
  NAND2_X1 U17469 ( .A1(n20175), .A2(n20156), .ZN(n14160) );
  NOR2_X1 U17470 ( .A1(n20170), .A2(n20792), .ZN(n20173) );
  NOR2_X1 U17471 ( .A1(n20161), .A2(n14157), .ZN(n14158) );
  AOI211_X1 U17472 ( .C1(n20152), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20173), .B(n14158), .ZN(n14159) );
  OAI211_X1 U17473 ( .C1(n12495), .C2(n14161), .A(n14160), .B(n14159), .ZN(
        P1_U2996) );
  INV_X1 U17474 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20088) );
  NAND2_X1 U17475 ( .A1(n14481), .A2(DATAI_8_), .ZN(n14163) );
  NAND2_X1 U17476 ( .A1(n14547), .A2(BUF1_REG_8__SCAN_IN), .ZN(n14162) );
  AND2_X1 U17477 ( .A1(n14163), .A2(n14162), .ZN(n20130) );
  OAI222_X1 U17478 ( .A1(n14553), .A2(n14203), .B1(n14550), .B2(n20088), .C1(
        n14562), .C2(n20130), .ZN(P1_U2896) );
  INV_X1 U17479 ( .A(n14022), .ZN(n14168) );
  INV_X1 U17480 ( .A(n14165), .ZN(n14166) );
  OAI211_X1 U17481 ( .C1(n14168), .C2(n14167), .A(n14166), .B(n15041), .ZN(
        n14175) );
  NAND2_X1 U17482 ( .A1(n14170), .A2(n14169), .ZN(n14173) );
  INV_X1 U17483 ( .A(n14171), .ZN(n14172) );
  AND2_X1 U17484 ( .A1(n14173), .A2(n14172), .ZN(n18988) );
  NAND2_X1 U17485 ( .A1(n15036), .A2(n18988), .ZN(n14174) );
  OAI211_X1 U17486 ( .C1(n15036), .C2(n10474), .A(n14175), .B(n14174), .ZN(
        P2_U2874) );
  INV_X1 U17487 ( .A(n14176), .ZN(n15605) );
  NAND2_X1 U17488 ( .A1(n19193), .A2(n15605), .ZN(n14185) );
  INV_X1 U17489 ( .A(n14177), .ZN(n14179) );
  NAND2_X1 U17490 ( .A1(n14179), .A2(n14178), .ZN(n15575) );
  NOR2_X1 U17491 ( .A1(n14180), .A2(n14181), .ZN(n14183) );
  AOI22_X1 U17492 ( .A1(n15575), .A2(n14183), .B1(n14182), .B2(n13609), .ZN(
        n14184) );
  NAND2_X1 U17493 ( .A1(n14185), .A2(n14184), .ZN(n16321) );
  AOI21_X1 U17494 ( .B1(n18993), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n14186), .ZN(n15593) );
  OAI22_X1 U17495 ( .A1(n14079), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n14187), .B2(n18993), .ZN(n15577) );
  NOR2_X1 U17496 ( .A1(n14188), .A2(n15577), .ZN(n15581) );
  AOI222_X1 U17497 ( .A1(n16321), .A2(n19900), .B1(n15593), .B2(n15581), .C1(
        n19923), .C2(n16362), .ZN(n14190) );
  NAND2_X1 U17498 ( .A1(n15607), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14189) );
  OAI21_X1 U17499 ( .B1(n14190), .B2(n15607), .A(n14189), .ZN(P2_U3600) );
  INV_X1 U17500 ( .A(n14191), .ZN(n14192) );
  OAI21_X1 U17501 ( .B1(n14148), .B2(n14193), .A(n14192), .ZN(n19999) );
  OAI222_X1 U17502 ( .A1(n19999), .A2(n14553), .B1(n20086), .B2(n14550), .C1(
        n14562), .C2(n14498), .ZN(P1_U2895) );
  XOR2_X1 U17503 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n14194), .Z(
        n14195) );
  XNOR2_X1 U17504 ( .A(n14196), .B(n14195), .ZN(n14208) );
  INV_X1 U17505 ( .A(n20013), .ZN(n14201) );
  NOR2_X1 U17506 ( .A1(n20170), .A2(n20802), .ZN(n14204) );
  INV_X1 U17507 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14198) );
  INV_X1 U17508 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16031) );
  NOR2_X1 U17509 ( .A1(n14198), .A2(n16031), .ZN(n16003) );
  AND2_X1 U17510 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n16046), .ZN(
        n14707) );
  NAND2_X1 U17511 ( .A1(n14707), .A2(n20181), .ZN(n14709) );
  NOR3_X1 U17512 ( .A1(n15975), .A2(n14709), .A3(n14197), .ZN(n16027) );
  OAI21_X1 U17513 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16027), .ZN(n14199) );
  OAI21_X1 U17514 ( .B1(n14707), .B2(n14787), .A(n20180), .ZN(n16043) );
  AOI21_X1 U17515 ( .B1(n14197), .B2(n16001), .A(n16043), .ZN(n16032) );
  OAI22_X1 U17516 ( .A1(n16003), .A2(n14199), .B1(n16032), .B2(n14198), .ZN(
        n14200) );
  AOI211_X1 U17517 ( .C1(n20203), .C2(n14201), .A(n14204), .B(n14200), .ZN(
        n14202) );
  OAI21_X1 U17518 ( .B1(n14208), .B2(n20208), .A(n14202), .ZN(P1_U3023) );
  INV_X1 U17519 ( .A(n14203), .ZN(n20017) );
  AOI21_X1 U17520 ( .B1(n20152), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n14204), .ZN(n14205) );
  OAI21_X1 U17521 ( .B1(n20161), .B2(n20009), .A(n14205), .ZN(n14206) );
  AOI21_X1 U17522 ( .B1(n20017), .B2(n20167), .A(n14206), .ZN(n14207) );
  OAI21_X1 U17523 ( .B1(n14208), .B2(n20172), .A(n14207), .ZN(P1_U2991) );
  XOR2_X1 U17524 ( .A(n14209), .B(n14191), .Z(n14702) );
  NAND2_X1 U17525 ( .A1(n16013), .A2(n14210), .ZN(n14211) );
  NAND2_X1 U17526 ( .A1(n14476), .A2(n14211), .ZN(n16004) );
  INV_X1 U17527 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14212) );
  OAI22_X1 U17528 ( .A1(n16004), .A2(n14467), .B1(n14212), .B2(n20075), .ZN(
        n14213) );
  AOI21_X1 U17529 ( .B1(n14702), .B2(n20071), .A(n14213), .ZN(n14214) );
  INV_X1 U17530 ( .A(n14214), .ZN(P1_U2862) );
  INV_X1 U17531 ( .A(n14702), .ZN(n14225) );
  NOR2_X1 U17532 ( .A1(n14215), .A2(n14377), .ZN(n15851) );
  NAND2_X1 U17533 ( .A1(n14217), .A2(n14216), .ZN(n20049) );
  AOI21_X1 U17534 ( .B1(n20048), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20040), .ZN(n14220) );
  OAI22_X1 U17535 ( .A1(n20054), .A2(n14212), .B1(n14700), .B2(n20053), .ZN(
        n14218) );
  INV_X1 U17536 ( .A(n14218), .ZN(n14219) );
  OAI211_X1 U17537 ( .C1(n20014), .C2(n16004), .A(n14220), .B(n14219), .ZN(
        n14221) );
  AOI221_X1 U17538 ( .B1(n15851), .B2(P1_REIP_REG_10__SCAN_IN), .C1(n14222), 
        .C2(n20806), .A(n14221), .ZN(n14223) );
  OAI21_X1 U17539 ( .B1(n14225), .B2(n14414), .A(n14223), .ZN(P1_U2830) );
  INV_X1 U17540 ( .A(n20132), .ZN(n14226) );
  INV_X1 U17541 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14224) );
  OAI222_X1 U17542 ( .A1(n14562), .A2(n14226), .B1(n14553), .B2(n14225), .C1(
        n14224), .C2(n14550), .ZN(P1_U2894) );
  XNOR2_X1 U17543 ( .A(n15883), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14227) );
  XNOR2_X1 U17544 ( .A(n14228), .B(n14227), .ZN(n16017) );
  NAND2_X1 U17545 ( .A1(n16017), .A2(n20156), .ZN(n14231) );
  INV_X1 U17546 ( .A(n20161), .ZN(n15878) );
  INV_X1 U17547 ( .A(n20152), .ZN(n20165) );
  OAI22_X1 U17548 ( .A1(n20165), .A2(n11886), .B1(n20170), .B2(n20804), .ZN(
        n14229) );
  AOI21_X1 U17549 ( .B1(n15878), .B2(n20002), .A(n14229), .ZN(n14230) );
  OAI211_X1 U17550 ( .C1(n12495), .C2(n19999), .A(n14231), .B(n14230), .ZN(
        P1_U2990) );
  AOI21_X1 U17551 ( .B1(n18691), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15712) );
  NAND2_X1 U17552 ( .A1(n15712), .A2(n17116), .ZN(n18223) );
  NOR2_X1 U17553 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18223), .ZN(n14232) );
  NAND3_X1 U17554 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18852)
         );
  OAI21_X1 U17555 ( .B1(n14232), .B2(n18852), .A(n18474), .ZN(n18229) );
  INV_X1 U17556 ( .A(n18229), .ZN(n14233) );
  NOR2_X1 U17557 ( .A1(n17859), .A2(n18900), .ZN(n15704) );
  AOI21_X1 U17558 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15704), .ZN(n15705) );
  NOR2_X1 U17559 ( .A1(n14233), .A2(n15705), .ZN(n14235) );
  NOR2_X1 U17560 ( .A1(n18854), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18270) );
  OR2_X1 U17561 ( .A1(n18270), .A2(n14233), .ZN(n15703) );
  OR2_X1 U17562 ( .A1(n18585), .A2(n15703), .ZN(n14234) );
  MUX2_X1 U17563 ( .A(n14235), .B(n14234), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  INV_X1 U17564 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n14237) );
  AOI22_X1 U17565 ( .A1(n14530), .A2(n20143), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n14528), .ZN(n14236) );
  OAI21_X1 U17566 ( .B1(n14237), .B2(n14532), .A(n14236), .ZN(n14238) );
  AOI21_X1 U17567 ( .B1(n14543), .B2(DATAI_30_), .A(n14238), .ZN(n14239) );
  OAI21_X1 U17568 ( .B1(n14241), .B2(n14553), .A(n14239), .ZN(P1_U2874) );
  INV_X1 U17569 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14240) );
  OAI222_X1 U17570 ( .A1(n14467), .A2(n14735), .B1(n14480), .B2(n14241), .C1(
        n14240), .C2(n20075), .ZN(P1_U2842) );
  NOR2_X2 U17571 ( .A1(n14242), .A2(n19217), .ZN(n19079) );
  NOR2_X2 U17572 ( .A1(n14242), .A2(n19219), .ZN(n19078) );
  AOI22_X1 U17573 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19079), .B1(n19078), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n14244) );
  AOI22_X1 U17574 ( .A1(n19077), .A2(n19089), .B1(n19130), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n14243) );
  OAI211_X1 U17575 ( .C1(n15300), .C2(n19122), .A(n14244), .B(n14243), .ZN(
        n14245) );
  INV_X1 U17576 ( .A(n14245), .ZN(n14246) );
  OAI21_X1 U17577 ( .B1(n14247), .B2(n19135), .A(n14246), .ZN(P2_U2889) );
  INV_X1 U17578 ( .A(n14575), .ZN(n14430) );
  AOI21_X1 U17579 ( .B1(n14248), .B2(n14255), .A(n9718), .ZN(n14747) );
  INV_X1 U17580 ( .A(n14249), .ZN(n14573) );
  AOI22_X1 U17581 ( .A1(n20048), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B1(
        n14250), .B2(n20963), .ZN(n14251) );
  OAI21_X1 U17582 ( .B1(n14430), .B2(n14414), .A(n14252), .ZN(P1_U2811) );
  OR2_X1 U17583 ( .A1(n14271), .A2(n14253), .ZN(n14254) );
  NAND2_X1 U17584 ( .A1(n14255), .A2(n14254), .ZN(n14754) );
  OAI21_X1 U17585 ( .B1(n14256), .B2(n14258), .A(n14257), .ZN(n14487) );
  INV_X1 U17586 ( .A(n14487), .ZN(n14587) );
  NAND2_X1 U17587 ( .A1(n14587), .A2(n20041), .ZN(n14268) );
  INV_X1 U17588 ( .A(n14259), .ZN(n14266) );
  INV_X1 U17589 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14431) );
  NAND2_X1 U17590 ( .A1(n20835), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14260) );
  NOR2_X1 U17591 ( .A1(n14275), .A2(n14260), .ZN(n14261) );
  AOI21_X1 U17592 ( .B1(n20048), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14261), .ZN(n14264) );
  INV_X1 U17593 ( .A(n14585), .ZN(n14262) );
  NAND2_X1 U17594 ( .A1(n20027), .A2(n14262), .ZN(n14263) );
  OAI211_X1 U17595 ( .C1(n20054), .C2(n14431), .A(n14264), .B(n14263), .ZN(
        n14265) );
  AOI21_X1 U17596 ( .B1(n14266), .B2(P1_REIP_REG_28__SCAN_IN), .A(n14265), 
        .ZN(n14267) );
  OAI211_X1 U17597 ( .C1(n14754), .C2(n20014), .A(n14268), .B(n14267), .ZN(
        P1_U2812) );
  NOR2_X1 U17598 ( .A1(n14287), .A2(n14269), .ZN(n14270) );
  OR2_X1 U17599 ( .A1(n14271), .A2(n14270), .ZN(n14761) );
  AOI21_X1 U17600 ( .B1(n14273), .B2(n14272), .A(n14256), .ZN(n14596) );
  NAND2_X1 U17601 ( .A1(n14596), .A2(n20041), .ZN(n14281) );
  AND2_X1 U17602 ( .A1(n20021), .A2(n14274), .ZN(n14292) );
  INV_X1 U17603 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14432) );
  NOR2_X1 U17604 ( .A1(n14275), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14276) );
  AOI21_X1 U17605 ( .B1(n20048), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14276), .ZN(n14278) );
  NAND2_X1 U17606 ( .A1(n20027), .A2(n14592), .ZN(n14277) );
  OAI211_X1 U17607 ( .C1(n20054), .C2(n14432), .A(n14278), .B(n14277), .ZN(
        n14279) );
  AOI21_X1 U17608 ( .B1(n14292), .B2(P1_REIP_REG_27__SCAN_IN), .A(n14279), 
        .ZN(n14280) );
  OAI211_X1 U17609 ( .C1(n14761), .C2(n20014), .A(n14281), .B(n14280), .ZN(
        P1_U2813) );
  OAI21_X1 U17610 ( .B1(n14282), .B2(n14283), .A(n14272), .ZN(n14601) );
  NAND2_X1 U17611 ( .A1(n15848), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n14286) );
  INV_X1 U17612 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21011) );
  NOR2_X1 U17613 ( .A1(n21011), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14284) );
  AOI22_X1 U17614 ( .A1(n20048), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n14301), .B2(n14284), .ZN(n14285) );
  OAI211_X1 U17615 ( .C1(n20053), .C2(n14603), .A(n14286), .B(n14285), .ZN(
        n14291) );
  INV_X1 U17616 ( .A(n14287), .ZN(n14288) );
  OAI21_X1 U17617 ( .B1(n14295), .B2(n14289), .A(n14288), .ZN(n14766) );
  NOR2_X1 U17618 ( .A1(n14766), .A2(n20014), .ZN(n14290) );
  AOI211_X1 U17619 ( .C1(n14292), .C2(P1_REIP_REG_26__SCAN_IN), .A(n14291), 
        .B(n14290), .ZN(n14293) );
  OAI21_X1 U17620 ( .B1(n14601), .B2(n14414), .A(n14293), .ZN(P1_U2814) );
  AND2_X1 U17621 ( .A1(n14312), .A2(n14294), .ZN(n14296) );
  OR2_X1 U17622 ( .A1(n14296), .A2(n14295), .ZN(n15912) );
  XOR2_X1 U17623 ( .A(n14299), .B(n14298), .Z(n14614) );
  NAND2_X1 U17624 ( .A1(n14614), .A2(n20041), .ZN(n14309) );
  INV_X1 U17625 ( .A(n14300), .ZN(n14612) );
  AOI22_X1 U17626 ( .A1(n20048), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        n14301), .B2(n21011), .ZN(n14302) );
  OAI21_X1 U17627 ( .B1(n20053), .B2(n14612), .A(n14302), .ZN(n14307) );
  OR2_X1 U17628 ( .A1(n14377), .A2(n14303), .ZN(n14332) );
  INV_X1 U17629 ( .A(n14304), .ZN(n14305) );
  NAND3_X1 U17630 ( .A1(n14305), .A2(n14355), .A3(n21010), .ZN(n14317) );
  AOI21_X1 U17631 ( .B1(n14332), .B2(n14317), .A(n21011), .ZN(n14306) );
  AOI211_X1 U17632 ( .C1(P1_EBX_REG_25__SCAN_IN), .C2(n15848), .A(n14307), .B(
        n14306), .ZN(n14308) );
  OAI211_X1 U17633 ( .C1(n15912), .C2(n20014), .A(n14309), .B(n14308), .ZN(
        P1_U2815) );
  OAI21_X1 U17634 ( .B1(n14310), .B2(n14311), .A(n14298), .ZN(n14623) );
  INV_X1 U17635 ( .A(n14312), .ZN(n14313) );
  AOI21_X1 U17636 ( .B1(n14314), .B2(n9714), .A(n14313), .ZN(n15917) );
  INV_X1 U17637 ( .A(n14315), .ZN(n14620) );
  NAND2_X1 U17638 ( .A1(n20027), .A2(n14620), .ZN(n14316) );
  OAI211_X1 U17639 ( .C1(n20000), .C2(n14618), .A(n14317), .B(n14316), .ZN(
        n14318) );
  AOI21_X1 U17640 ( .B1(n15848), .B2(P1_EBX_REG_24__SCAN_IN), .A(n14318), .ZN(
        n14319) );
  OAI21_X1 U17641 ( .B1(n14332), .B2(n21010), .A(n14319), .ZN(n14320) );
  AOI21_X1 U17642 ( .B1(n15917), .B2(n20047), .A(n14320), .ZN(n14321) );
  OAI21_X1 U17643 ( .B1(n14623), .B2(n14414), .A(n14321), .ZN(P1_U2816) );
  AOI21_X1 U17644 ( .B1(n14323), .B2(n14322), .A(n14310), .ZN(n14634) );
  INV_X1 U17645 ( .A(n14634), .ZN(n14510) );
  NAND2_X1 U17646 ( .A1(n9753), .A2(n14324), .ZN(n14325) );
  NAND2_X1 U17647 ( .A1(n9714), .A2(n14325), .ZN(n14436) );
  INV_X1 U17648 ( .A(n14436), .ZN(n15930) );
  AOI21_X1 U17649 ( .B1(n14355), .B2(n14326), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n14331) );
  INV_X1 U17650 ( .A(n14327), .ZN(n14632) );
  OAI22_X1 U17651 ( .A1(n14328), .A2(n20000), .B1(n20053), .B2(n14632), .ZN(
        n14329) );
  AOI21_X1 U17652 ( .B1(P1_EBX_REG_23__SCAN_IN), .B2(n15848), .A(n14329), .ZN(
        n14330) );
  OAI21_X1 U17653 ( .B1(n14332), .B2(n14331), .A(n14330), .ZN(n14333) );
  AOI21_X1 U17654 ( .B1(n15930), .B2(n20047), .A(n14333), .ZN(n14334) );
  OAI21_X1 U17655 ( .B1(n14510), .B2(n14414), .A(n14334), .ZN(P1_U2817) );
  OR2_X1 U17656 ( .A1(n14351), .A2(n14335), .ZN(n14336) );
  NAND2_X1 U17657 ( .A1(n9753), .A2(n14336), .ZN(n14774) );
  OAI21_X1 U17658 ( .B1(n14337), .B2(n14338), .A(n14322), .ZN(n14514) );
  INV_X1 U17659 ( .A(n14514), .ZN(n14642) );
  NAND2_X1 U17660 ( .A1(n14642), .A2(n20041), .ZN(n14347) );
  NAND2_X1 U17661 ( .A1(n20021), .A2(n14339), .ZN(n15810) );
  INV_X1 U17662 ( .A(n15810), .ZN(n14345) );
  INV_X1 U17663 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14438) );
  INV_X1 U17664 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21023) );
  XNOR2_X1 U17665 ( .A(n21023), .B(P1_REIP_REG_21__SCAN_IN), .ZN(n14340) );
  AOI22_X1 U17666 ( .A1(n20048), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n14355), .B2(n14340), .ZN(n14343) );
  INV_X1 U17667 ( .A(n14640), .ZN(n14341) );
  NAND2_X1 U17668 ( .A1(n20027), .A2(n14341), .ZN(n14342) );
  OAI211_X1 U17669 ( .C1(n20054), .C2(n14438), .A(n14343), .B(n14342), .ZN(
        n14344) );
  AOI21_X1 U17670 ( .B1(n14345), .B2(P1_REIP_REG_22__SCAN_IN), .A(n14344), 
        .ZN(n14346) );
  OAI211_X1 U17671 ( .C1(n14774), .C2(n20014), .A(n14347), .B(n14346), .ZN(
        P1_U2818) );
  OAI21_X1 U17672 ( .B1(n9684), .B2(n14348), .A(n10268), .ZN(n14518) );
  INV_X1 U17673 ( .A(n14518), .ZN(n14649) );
  NOR2_X1 U17674 ( .A1(n14442), .A2(n14349), .ZN(n14350) );
  OR2_X1 U17675 ( .A1(n14351), .A2(n14350), .ZN(n15766) );
  INV_X1 U17676 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20985) );
  INV_X1 U17677 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14439) );
  OAI22_X1 U17678 ( .A1(n20054), .A2(n14439), .B1(n14647), .B2(n20053), .ZN(
        n14352) );
  INV_X1 U17679 ( .A(n14352), .ZN(n14353) );
  OAI21_X1 U17680 ( .B1(n20985), .B2(n15810), .A(n14353), .ZN(n14354) );
  AOI21_X1 U17681 ( .B1(n14355), .B2(n20985), .A(n14354), .ZN(n14357) );
  NAND2_X1 U17682 ( .A1(n20048), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14356) );
  OAI211_X1 U17683 ( .C1(n15766), .C2(n20014), .A(n14357), .B(n14356), .ZN(
        n14358) );
  AOI21_X1 U17684 ( .B1(n14649), .B2(n20041), .A(n14358), .ZN(n14359) );
  INV_X1 U17685 ( .A(n14359), .ZN(P1_U2819) );
  OAI21_X1 U17686 ( .B1(n14360), .B2(n14362), .A(n14361), .ZN(n14654) );
  NAND2_X1 U17687 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n14363) );
  OAI211_X1 U17688 ( .C1(P1_REIP_REG_19__SCAN_IN), .C2(P1_REIP_REG_18__SCAN_IN), .A(n15815), .B(n14363), .ZN(n14373) );
  NAND2_X1 U17689 ( .A1(n14448), .A2(n14364), .ZN(n14365) );
  AND2_X1 U17690 ( .A1(n14441), .A2(n14365), .ZN(n15938) );
  INV_X1 U17691 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14366) );
  OAI22_X1 U17692 ( .A1(n20054), .A2(n14366), .B1(n14656), .B2(n20053), .ZN(
        n14367) );
  INV_X1 U17693 ( .A(n14367), .ZN(n14368) );
  OAI211_X1 U17694 ( .C1(n20000), .C2(n14369), .A(n14368), .B(n20049), .ZN(
        n14371) );
  INV_X1 U17695 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20823) );
  NOR3_X1 U17696 ( .A1(n14377), .A2(n14378), .A3(n20823), .ZN(n14370) );
  AOI211_X1 U17697 ( .C1(n15938), .C2(n20047), .A(n14371), .B(n14370), .ZN(
        n14372) );
  OAI211_X1 U17698 ( .C1(n14654), .C2(n14414), .A(n14373), .B(n14372), .ZN(
        P1_U2821) );
  OAI21_X1 U17699 ( .B1(n9685), .B2(n12008), .A(n14376), .ZN(n14674) );
  INV_X1 U17700 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20814) );
  NOR2_X1 U17701 ( .A1(n15828), .A2(n20814), .ZN(n14397) );
  NOR2_X1 U17702 ( .A1(n14378), .A2(n14377), .ZN(n15811) );
  OAI221_X1 U17703 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(P1_REIP_REG_16__SCAN_IN), .C1(P1_REIP_REG_17__SCAN_IN), .C2(n14397), .A(n15811), .ZN(n14386) );
  INV_X1 U17704 ( .A(n14450), .ZN(n14379) );
  OAI21_X1 U17705 ( .B1(n14380), .B2(n14392), .A(n14379), .ZN(n14452) );
  INV_X1 U17706 ( .A(n14452), .ZN(n15954) );
  INV_X1 U17707 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14453) );
  OAI22_X1 U17708 ( .A1(n20054), .A2(n14453), .B1(n14676), .B2(n20053), .ZN(
        n14381) );
  INV_X1 U17709 ( .A(n14381), .ZN(n14382) );
  OAI211_X1 U17710 ( .C1(n20000), .C2(n14383), .A(n14382), .B(n20049), .ZN(
        n14384) );
  AOI21_X1 U17711 ( .B1(n15954), .B2(n20047), .A(n14384), .ZN(n14385) );
  OAI211_X1 U17712 ( .C1(n14674), .C2(n14414), .A(n14386), .B(n14385), .ZN(
        P1_U2823) );
  AOI21_X1 U17713 ( .B1(n14388), .B2(n14387), .A(n9685), .ZN(n15864) );
  INV_X1 U17714 ( .A(n15864), .ZN(n14546) );
  INV_X1 U17715 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20817) );
  NAND2_X1 U17716 ( .A1(n20021), .A2(n14389), .ZN(n15835) );
  OAI21_X1 U17717 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n15828), .A(n15835), 
        .ZN(n14396) );
  AND2_X1 U17718 ( .A1(n14460), .A2(n14390), .ZN(n14391) );
  NOR2_X1 U17719 ( .A1(n14392), .A2(n14391), .ZN(n14454) );
  INV_X1 U17720 ( .A(n14454), .ZN(n14795) );
  INV_X1 U17721 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14457) );
  OAI22_X1 U17722 ( .A1(n14795), .A2(n20014), .B1(n14457), .B2(n20054), .ZN(
        n14393) );
  AOI211_X1 U17723 ( .C1(n20048), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n20040), .B(n14393), .ZN(n14394) );
  OAI21_X1 U17724 ( .B1(n15867), .B2(n20053), .A(n14394), .ZN(n14395) );
  AOI221_X1 U17725 ( .B1(n14397), .B2(n20817), .C1(n14396), .C2(
        P1_REIP_REG_16__SCAN_IN), .A(n14395), .ZN(n14398) );
  OAI21_X1 U17726 ( .B1(n14546), .B2(n14414), .A(n14398), .ZN(P1_U2824) );
  OAI21_X1 U17727 ( .B1(n14399), .B2(n14401), .A(n14400), .ZN(n14696) );
  INV_X1 U17728 ( .A(n14692), .ZN(n14412) );
  AOI21_X1 U17729 ( .B1(n15840), .B2(n15838), .A(n14402), .ZN(n14403) );
  NOR2_X1 U17730 ( .A1(n14403), .A2(n14465), .ZN(n15969) );
  AOI22_X1 U17731 ( .A1(n15969), .A2(n20047), .B1(n15848), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14404) );
  OAI211_X1 U17732 ( .C1(n20000), .C2(n14405), .A(n14404), .B(n20049), .ZN(
        n14411) );
  NOR2_X1 U17733 ( .A1(n15854), .A2(n14406), .ZN(n14409) );
  AOI21_X1 U17734 ( .B1(n14407), .B2(n14406), .A(n15851), .ZN(n15847) );
  INV_X1 U17735 ( .A(n15847), .ZN(n14408) );
  MUX2_X1 U17736 ( .A(n14409), .B(n14408), .S(P1_REIP_REG_13__SCAN_IN), .Z(
        n14410) );
  AOI211_X1 U17737 ( .C1(n20027), .C2(n14412), .A(n14411), .B(n14410), .ZN(
        n14413) );
  OAI21_X1 U17738 ( .B1(n14696), .B2(n14414), .A(n14413), .ZN(P1_U2827) );
  NAND3_X1 U17739 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n14415) );
  NOR3_X1 U17740 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n14416), .A3(n14415), .ZN(
        n14426) );
  NAND2_X1 U17741 ( .A1(n20022), .A2(n20021), .ZN(n20060) );
  INV_X1 U17742 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20793) );
  AOI21_X1 U17743 ( .B1(n20048), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20040), .ZN(n14417) );
  OAI21_X1 U17744 ( .B1(n20160), .B2(n20053), .A(n14417), .ZN(n14418) );
  AOI21_X1 U17745 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(n15848), .A(n14418), .ZN(
        n14419) );
  OAI21_X1 U17746 ( .B1(n20014), .B2(n14420), .A(n14419), .ZN(n14421) );
  AOI21_X1 U17747 ( .B1(n14423), .B2(n14422), .A(n14421), .ZN(n14424) );
  OAI21_X1 U17748 ( .B1(n20060), .B2(n20793), .A(n14424), .ZN(n14425) );
  AOI211_X1 U17749 ( .C1(n20155), .C2(n20046), .A(n14426), .B(n14425), .ZN(
        n14427) );
  INV_X1 U17750 ( .A(n14427), .ZN(P1_U2836) );
  OAI22_X1 U17751 ( .A1(n14706), .A2(n14467), .B1(n20075), .B2(n14428), .ZN(
        P1_U2841) );
  AOI22_X1 U17752 ( .A1(n14747), .A2(n20070), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14478), .ZN(n14429) );
  OAI21_X1 U17753 ( .B1(n14430), .B2(n14480), .A(n14429), .ZN(P1_U2843) );
  OAI222_X1 U17754 ( .A1(n14480), .A2(n14487), .B1(n14431), .B2(n20075), .C1(
        n14754), .C2(n14467), .ZN(P1_U2844) );
  INV_X1 U17755 ( .A(n14596), .ZN(n14492) );
  OAI222_X1 U17756 ( .A1(n14480), .A2(n14492), .B1(n14432), .B2(n20075), .C1(
        n14761), .C2(n14467), .ZN(P1_U2845) );
  INV_X1 U17757 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14433) );
  OAI222_X1 U17758 ( .A1(n14601), .A2(n14480), .B1(n14433), .B2(n20075), .C1(
        n14766), .C2(n14467), .ZN(P1_U2846) );
  INV_X1 U17759 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14434) );
  INV_X1 U17760 ( .A(n14614), .ZN(n14502) );
  OAI222_X1 U17761 ( .A1(n15912), .A2(n14467), .B1(n14434), .B2(n20075), .C1(
        n14480), .C2(n14502), .ZN(P1_U2847) );
  AOI22_X1 U17762 ( .A1(n15917), .A2(n20070), .B1(P1_EBX_REG_24__SCAN_IN), 
        .B2(n14478), .ZN(n14435) );
  OAI21_X1 U17763 ( .B1(n14623), .B2(n14480), .A(n14435), .ZN(P1_U2848) );
  INV_X1 U17764 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14437) );
  OAI222_X1 U17765 ( .A1(n14510), .A2(n14480), .B1(n20075), .B2(n14437), .C1(
        n14436), .C2(n14467), .ZN(P1_U2849) );
  OAI222_X1 U17766 ( .A1(n14514), .A2(n14480), .B1(n14438), .B2(n20075), .C1(
        n14774), .C2(n14467), .ZN(P1_U2850) );
  OAI222_X1 U17767 ( .A1(n14518), .A2(n14480), .B1(n14439), .B2(n20075), .C1(
        n15766), .C2(n14467), .ZN(P1_U2851) );
  AND2_X1 U17768 ( .A1(n14441), .A2(n14440), .ZN(n14443) );
  OR2_X1 U17769 ( .A1(n14443), .A2(n14442), .ZN(n15805) );
  AOI21_X1 U17770 ( .B1(n14444), .B2(n14361), .A(n9684), .ZN(n15807) );
  INV_X1 U17771 ( .A(n15807), .ZN(n15858) );
  OAI222_X1 U17772 ( .A1(n15805), .A2(n14467), .B1(n20075), .B2(n12420), .C1(
        n15858), .C2(n14480), .ZN(P1_U2852) );
  AOI22_X1 U17773 ( .A1(n15938), .A2(n20070), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14478), .ZN(n14445) );
  OAI21_X1 U17774 ( .B1(n14654), .B2(n14480), .A(n14445), .ZN(P1_U2853) );
  AND2_X1 U17775 ( .A1(n14376), .A2(n14446), .ZN(n14447) );
  OR2_X1 U17776 ( .A1(n14447), .A2(n14360), .ZN(n14663) );
  INV_X1 U17777 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14451) );
  OAI21_X1 U17778 ( .B1(n14450), .B2(n14449), .A(n14448), .ZN(n15944) );
  OAI222_X1 U17779 ( .A1(n14663), .A2(n14480), .B1(n14451), .B2(n20075), .C1(
        n15944), .C2(n14467), .ZN(P1_U2854) );
  OAI222_X1 U17780 ( .A1(n14674), .A2(n14480), .B1(n14453), .B2(n20075), .C1(
        n14452), .C2(n14467), .ZN(P1_U2855) );
  NAND2_X1 U17781 ( .A1(n15864), .A2(n20071), .ZN(n14456) );
  NAND2_X1 U17782 ( .A1(n14454), .A2(n20070), .ZN(n14455) );
  OAI211_X1 U17783 ( .C1(n14457), .C2(n20075), .A(n14456), .B(n14455), .ZN(
        P1_U2856) );
  OAI21_X1 U17784 ( .B1(n14458), .B2(n14459), .A(n14387), .ZN(n15820) );
  AOI21_X1 U17785 ( .B1(n14461), .B2(n9703), .A(n10073), .ZN(n15962) );
  AOI22_X1 U17786 ( .A1(n15962), .A2(n20070), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n14478), .ZN(n14462) );
  OAI21_X1 U17787 ( .B1(n15820), .B2(n14480), .A(n14462), .ZN(P1_U2857) );
  AOI21_X1 U17788 ( .B1(n14463), .B2(n14400), .A(n14458), .ZN(n15869) );
  OAI21_X1 U17789 ( .B1(n14465), .B2(n14464), .A(n9703), .ZN(n15829) );
  INV_X1 U17790 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14466) );
  OAI22_X1 U17791 ( .A1(n15829), .A2(n14467), .B1(n14466), .B2(n20075), .ZN(
        n14468) );
  AOI21_X1 U17792 ( .B1(n15869), .B2(n20071), .A(n14468), .ZN(n14469) );
  INV_X1 U17793 ( .A(n14469), .ZN(P1_U2858) );
  AOI22_X1 U17794 ( .A1(n15969), .A2(n20070), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14478), .ZN(n14470) );
  OAI21_X1 U17795 ( .B1(n14696), .B2(n14480), .A(n14470), .ZN(P1_U2859) );
  NAND2_X1 U17796 ( .A1(n14471), .A2(n14472), .ZN(n14473) );
  AND2_X1 U17797 ( .A1(n14474), .A2(n14473), .ZN(n15887) );
  INV_X1 U17798 ( .A(n15887), .ZN(n14564) );
  AND2_X1 U17799 ( .A1(n14476), .A2(n14475), .ZN(n14477) );
  NOR2_X1 U17800 ( .A1(n15840), .A2(n14477), .ZN(n15991) );
  AOI22_X1 U17801 ( .A1(n15991), .A2(n20070), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n14478), .ZN(n14479) );
  OAI21_X1 U17802 ( .B1(n14564), .B2(n14480), .A(n14479), .ZN(P1_U2861) );
  NAND2_X1 U17803 ( .A1(n14481), .A2(DATAI_12_), .ZN(n14483) );
  NAND2_X1 U17804 ( .A1(n14547), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14482) );
  AND2_X1 U17805 ( .A1(n14483), .A2(n14482), .ZN(n20139) );
  OAI22_X1 U17806 ( .A1(n14540), .A2(n20139), .B1(n14550), .B2(n13660), .ZN(
        n14484) );
  AOI21_X1 U17807 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n14542), .A(n14484), .ZN(
        n14486) );
  NAND2_X1 U17808 ( .A1(n14543), .A2(DATAI_28_), .ZN(n14485) );
  OAI211_X1 U17809 ( .C1(n14487), .C2(n14553), .A(n14486), .B(n14485), .ZN(
        P1_U2876) );
  INV_X1 U17810 ( .A(n20135), .ZN(n14561) );
  OAI22_X1 U17811 ( .A1(n14540), .A2(n14561), .B1(n14550), .B2(n14488), .ZN(
        n14489) );
  AOI21_X1 U17812 ( .B1(BUF1_REG_27__SCAN_IN), .B2(n14542), .A(n14489), .ZN(
        n14491) );
  NAND2_X1 U17813 ( .A1(n14543), .A2(DATAI_27_), .ZN(n14490) );
  OAI211_X1 U17814 ( .C1(n14492), .C2(n14553), .A(n14491), .B(n14490), .ZN(
        P1_U2877) );
  INV_X1 U17815 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n14494) );
  AOI22_X1 U17816 ( .A1(n14530), .A2(n20132), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n14528), .ZN(n14493) );
  OAI21_X1 U17817 ( .B1(n14532), .B2(n14494), .A(n14493), .ZN(n14495) );
  AOI21_X1 U17818 ( .B1(n14543), .B2(DATAI_26_), .A(n14495), .ZN(n14496) );
  OAI21_X1 U17819 ( .B1(n14601), .B2(n14553), .A(n14496), .ZN(P1_U2878) );
  INV_X1 U17820 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20219) );
  NOR2_X1 U17821 ( .A1(n14532), .A2(n20219), .ZN(n14500) );
  OAI22_X1 U17822 ( .A1(n14540), .A2(n14498), .B1(n14550), .B2(n14497), .ZN(
        n14499) );
  AOI211_X1 U17823 ( .C1(DATAI_25_), .C2(n14543), .A(n14500), .B(n14499), .ZN(
        n14501) );
  OAI21_X1 U17824 ( .B1(n14502), .B2(n14553), .A(n14501), .ZN(P1_U2879) );
  OAI22_X1 U17825 ( .A1(n14540), .A2(n20130), .B1(n14550), .B2(n13668), .ZN(
        n14503) );
  AOI21_X1 U17826 ( .B1(n14542), .B2(BUF1_REG_24__SCAN_IN), .A(n14503), .ZN(
        n14505) );
  NAND2_X1 U17827 ( .A1(n14543), .A2(DATAI_24_), .ZN(n14504) );
  OAI211_X1 U17828 ( .C1(n14623), .C2(n14553), .A(n14505), .B(n14504), .ZN(
        P1_U2880) );
  OAI22_X1 U17829 ( .A1(n14540), .A2(n20128), .B1(n14550), .B2(n14506), .ZN(
        n14507) );
  AOI21_X1 U17830 ( .B1(n14542), .B2(BUF1_REG_23__SCAN_IN), .A(n14507), .ZN(
        n14509) );
  NAND2_X1 U17831 ( .A1(n14543), .A2(DATAI_23_), .ZN(n14508) );
  OAI211_X1 U17832 ( .C1(n14510), .C2(n14553), .A(n14509), .B(n14508), .ZN(
        P1_U2881) );
  OAI22_X1 U17833 ( .A1(n14540), .A2(n20246), .B1(n14550), .B2(n13658), .ZN(
        n14511) );
  AOI21_X1 U17834 ( .B1(n14542), .B2(BUF1_REG_22__SCAN_IN), .A(n14511), .ZN(
        n14513) );
  NAND2_X1 U17835 ( .A1(n14543), .A2(DATAI_22_), .ZN(n14512) );
  OAI211_X1 U17836 ( .C1(n14514), .C2(n14553), .A(n14513), .B(n14512), .ZN(
        P1_U2882) );
  OAI22_X1 U17837 ( .A1(n14540), .A2(n20125), .B1(n14550), .B2(n13656), .ZN(
        n14515) );
  AOI21_X1 U17838 ( .B1(n14542), .B2(BUF1_REG_21__SCAN_IN), .A(n14515), .ZN(
        n14517) );
  NAND2_X1 U17839 ( .A1(n14543), .A2(DATAI_21_), .ZN(n14516) );
  OAI211_X1 U17840 ( .C1(n14518), .C2(n14553), .A(n14517), .B(n14516), .ZN(
        P1_U2883) );
  INV_X1 U17841 ( .A(DATAI_20_), .ZN(n14523) );
  NAND2_X1 U17842 ( .A1(n15807), .A2(n12600), .ZN(n14522) );
  OAI22_X1 U17843 ( .A1(n14540), .A2(n20123), .B1(n14550), .B2(n14519), .ZN(
        n14520) );
  AOI21_X1 U17844 ( .B1(n14542), .B2(BUF1_REG_20__SCAN_IN), .A(n14520), .ZN(
        n14521) );
  OAI211_X1 U17845 ( .C1(n14524), .C2(n14523), .A(n14522), .B(n14521), .ZN(
        P1_U2884) );
  OAI22_X1 U17846 ( .A1(n14540), .A2(n20228), .B1(n14550), .B2(n13662), .ZN(
        n14525) );
  AOI21_X1 U17847 ( .B1(n14542), .B2(BUF1_REG_19__SCAN_IN), .A(n14525), .ZN(
        n14527) );
  NAND2_X1 U17848 ( .A1(n14543), .A2(DATAI_19_), .ZN(n14526) );
  OAI211_X1 U17849 ( .C1(n14654), .C2(n14553), .A(n14527), .B(n14526), .ZN(
        P1_U2885) );
  INV_X1 U17850 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16426) );
  INV_X1 U17851 ( .A(n20120), .ZN(n14529) );
  AOI22_X1 U17852 ( .A1(n14530), .A2(n14529), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n14528), .ZN(n14531) );
  OAI21_X1 U17853 ( .B1(n16426), .B2(n14532), .A(n14531), .ZN(n14533) );
  AOI21_X1 U17854 ( .B1(n14543), .B2(DATAI_18_), .A(n14533), .ZN(n14534) );
  OAI21_X1 U17855 ( .B1(n14663), .B2(n14553), .A(n14534), .ZN(P1_U2886) );
  OAI22_X1 U17856 ( .A1(n14540), .A2(n20118), .B1(n14550), .B2(n14535), .ZN(
        n14536) );
  AOI21_X1 U17857 ( .B1(n14542), .B2(BUF1_REG_17__SCAN_IN), .A(n14536), .ZN(
        n14538) );
  NAND2_X1 U17858 ( .A1(n14543), .A2(DATAI_17_), .ZN(n14537) );
  OAI211_X1 U17859 ( .C1(n14674), .C2(n14553), .A(n14538), .B(n14537), .ZN(
        P1_U2887) );
  OAI22_X1 U17860 ( .A1(n14540), .A2(n20214), .B1(n14550), .B2(n14539), .ZN(
        n14541) );
  AOI21_X1 U17861 ( .B1(n14542), .B2(BUF1_REG_16__SCAN_IN), .A(n14541), .ZN(
        n14545) );
  NAND2_X1 U17862 ( .A1(n14543), .A2(DATAI_16_), .ZN(n14544) );
  OAI211_X1 U17863 ( .C1(n14546), .C2(n14553), .A(n14545), .B(n14544), .ZN(
        P1_U2888) );
  INV_X1 U17864 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20078) );
  INV_X1 U17865 ( .A(DATAI_15_), .ZN(n14549) );
  INV_X1 U17866 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n14548) );
  MUX2_X1 U17867 ( .A(n14549), .B(n14548), .S(n14547), .Z(n20151) );
  OAI222_X1 U17868 ( .A1(n14553), .A2(n15820), .B1(n14550), .B2(n20078), .C1(
        n14562), .C2(n20151), .ZN(P1_U2889) );
  INV_X1 U17869 ( .A(n15869), .ZN(n14554) );
  INV_X1 U17870 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14552) );
  INV_X1 U17871 ( .A(n20143), .ZN(n14551) );
  OAI222_X1 U17872 ( .A1(n14554), .A2(n14553), .B1(n14552), .B2(n14550), .C1(
        n14562), .C2(n14551), .ZN(P1_U2890) );
  INV_X1 U17873 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14556) );
  OAI222_X1 U17874 ( .A1(n14696), .A2(n14553), .B1(n14556), .B2(n14550), .C1(
        n14562), .C2(n14555), .ZN(P1_U2891) );
  NOR2_X1 U17875 ( .A1(n14557), .A2(n14558), .ZN(n14559) );
  NOR2_X1 U17876 ( .A1(n14399), .A2(n14559), .ZN(n15880) );
  INV_X1 U17877 ( .A(n15880), .ZN(n14560) );
  INV_X1 U17878 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20082) );
  OAI222_X1 U17879 ( .A1(n14553), .A2(n14560), .B1(n14550), .B2(n20082), .C1(
        n14562), .C2(n20139), .ZN(P1_U2892) );
  INV_X1 U17880 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14563) );
  OAI222_X1 U17881 ( .A1(n14564), .A2(n14553), .B1(n14563), .B2(n14550), .C1(
        n14562), .C2(n14561), .ZN(P1_U2893) );
  NOR2_X1 U17882 ( .A1(n14566), .A2(n14565), .ZN(n14571) );
  INV_X1 U17883 ( .A(n14567), .ZN(n14569) );
  XOR2_X1 U17884 ( .A(n14571), .B(n14570), .Z(n14751) );
  NOR2_X1 U17885 ( .A1(n20170), .A2(n20963), .ZN(n14746) );
  AOI21_X1 U17886 ( .B1(n20152), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14746), .ZN(n14572) );
  OAI21_X1 U17887 ( .B1(n20161), .B2(n14573), .A(n14572), .ZN(n14574) );
  AOI21_X1 U17888 ( .B1(n14575), .B2(n20154), .A(n14574), .ZN(n14576) );
  OAI21_X1 U17889 ( .B1(n14751), .B2(n20172), .A(n14576), .ZN(P1_U2970) );
  NAND3_X1 U17890 ( .A1(n14578), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14579) );
  INV_X1 U17891 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14582) );
  NOR2_X1 U17892 ( .A1(n20170), .A2(n20835), .ZN(n14752) );
  AOI21_X1 U17893 ( .B1(n20152), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14752), .ZN(n14584) );
  OAI21_X1 U17894 ( .B1(n20161), .B2(n14585), .A(n14584), .ZN(n14586) );
  AOI21_X1 U17895 ( .B1(n14587), .B2(n20154), .A(n14586), .ZN(n14588) );
  OAI21_X1 U17896 ( .B1(n20172), .B2(n14755), .A(n14588), .ZN(P1_U2971) );
  MUX2_X1 U17897 ( .A(n14590), .B(n14589), .S(n10313), .Z(n14591) );
  INV_X1 U17898 ( .A(n14592), .ZN(n14594) );
  AOI22_X1 U17899 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B1(
        n20190), .B2(P1_REIP_REG_27__SCAN_IN), .ZN(n14593) );
  OAI21_X1 U17900 ( .B1(n20161), .B2(n14594), .A(n14593), .ZN(n14595) );
  AOI21_X1 U17901 ( .B1(n14596), .B2(n20167), .A(n14595), .ZN(n14597) );
  OAI21_X1 U17902 ( .B1(n20172), .B2(n14762), .A(n14597), .ZN(P1_U2972) );
  INV_X1 U17903 ( .A(n14625), .ZN(n14607) );
  NOR2_X1 U17904 ( .A1(n14607), .A2(n14718), .ZN(n14598) );
  MUX2_X1 U17905 ( .A(n14599), .B(n14598), .S(n15883), .Z(n14600) );
  XNOR2_X1 U17906 ( .A(n14600), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14773) );
  INV_X1 U17907 ( .A(n14601), .ZN(n14605) );
  AOI22_X1 U17908 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n20190), .B2(P1_REIP_REG_26__SCAN_IN), .ZN(n14602) );
  OAI21_X1 U17909 ( .B1(n20161), .B2(n14603), .A(n14602), .ZN(n14604) );
  AOI21_X1 U17910 ( .B1(n14605), .B2(n20167), .A(n14604), .ZN(n14606) );
  OAI21_X1 U17911 ( .B1(n20172), .B2(n14773), .A(n14606), .ZN(P1_U2973) );
  NAND2_X1 U17912 ( .A1(n14607), .A2(n10313), .ZN(n14624) );
  NAND2_X1 U17913 ( .A1(n14608), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14616) );
  OAI33_X1 U17914 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n14624), .B1(n14609), .B2(
        n10313), .B3(n14616), .ZN(n14610) );
  XNOR2_X1 U17915 ( .A(n14610), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15916) );
  AOI22_X1 U17916 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        n20190), .B2(P1_REIP_REG_25__SCAN_IN), .ZN(n14611) );
  OAI21_X1 U17917 ( .B1(n20161), .B2(n14612), .A(n14611), .ZN(n14613) );
  AOI21_X1 U17918 ( .B1(n14614), .B2(n20167), .A(n14613), .ZN(n14615) );
  OAI21_X1 U17919 ( .B1(n15916), .B2(n20172), .A(n14615), .ZN(P1_U2974) );
  MUX2_X1 U17920 ( .A(n10313), .B(n14624), .S(n14616), .Z(n14617) );
  XNOR2_X1 U17921 ( .A(n14617), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15918) );
  NAND2_X1 U17922 ( .A1(n15918), .A2(n20156), .ZN(n14622) );
  OAI22_X1 U17923 ( .A1(n20165), .A2(n14618), .B1(n20170), .B2(n21010), .ZN(
        n14619) );
  AOI21_X1 U17924 ( .B1(n14620), .B2(n15878), .A(n14619), .ZN(n14621) );
  OAI211_X1 U17925 ( .C1(n12495), .C2(n14623), .A(n14622), .B(n14621), .ZN(
        P1_U2975) );
  INV_X1 U17926 ( .A(n14624), .ZN(n14630) );
  NOR2_X1 U17927 ( .A1(n10313), .A2(n14629), .ZN(n14627) );
  MUX2_X1 U17928 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n14629), .S(
        n15883), .Z(n14626) );
  MUX2_X1 U17929 ( .A(n14627), .B(n14626), .S(n14625), .Z(n14628) );
  AOI21_X1 U17930 ( .B1(n14630), .B2(n14629), .A(n14628), .ZN(n15929) );
  AOI22_X1 U17931 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n20190), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n14631) );
  OAI21_X1 U17932 ( .B1(n20161), .B2(n14632), .A(n14631), .ZN(n14633) );
  AOI21_X1 U17933 ( .B1(n14634), .B2(n20167), .A(n14633), .ZN(n14635) );
  OAI21_X1 U17934 ( .B1(n15929), .B2(n20172), .A(n14635), .ZN(P1_U2976) );
  NAND2_X1 U17935 ( .A1(n14637), .A2(n14636), .ZN(n14638) );
  XOR2_X1 U17936 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n14638), .Z(
        n14782) );
  NOR2_X1 U17937 ( .A1(n20170), .A2(n21023), .ZN(n14776) );
  AOI21_X1 U17938 ( .B1(n20152), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n14776), .ZN(n14639) );
  OAI21_X1 U17939 ( .B1(n20161), .B2(n14640), .A(n14639), .ZN(n14641) );
  AOI21_X1 U17940 ( .B1(n14642), .B2(n20167), .A(n14641), .ZN(n14643) );
  OAI21_X1 U17941 ( .B1(n20172), .B2(n14782), .A(n14643), .ZN(P1_U2977) );
  MUX2_X1 U17942 ( .A(n14644), .B(n9695), .S(n10313), .Z(n14645) );
  XNOR2_X1 U17943 ( .A(n14645), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15765) );
  AOI22_X1 U17944 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n20190), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n14646) );
  OAI21_X1 U17945 ( .B1(n20161), .B2(n14647), .A(n14646), .ZN(n14648) );
  AOI21_X1 U17946 ( .B1(n14649), .B2(n20167), .A(n14648), .ZN(n14650) );
  OAI21_X1 U17947 ( .B1(n15765), .B2(n20172), .A(n14650), .ZN(P1_U2978) );
  NOR2_X1 U17948 ( .A1(n15883), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14652) );
  MUX2_X1 U17949 ( .A(n15883), .B(n14652), .S(n14651), .Z(n14653) );
  XNOR2_X1 U17950 ( .A(n14653), .B(n15936), .ZN(n15939) );
  INV_X1 U17951 ( .A(n15939), .ZN(n14660) );
  INV_X1 U17952 ( .A(n14654), .ZN(n14658) );
  AOI22_X1 U17953 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n20190), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n14655) );
  OAI21_X1 U17954 ( .B1(n20161), .B2(n14656), .A(n14655), .ZN(n14657) );
  AOI21_X1 U17955 ( .B1(n14658), .B2(n20167), .A(n14657), .ZN(n14659) );
  OAI21_X1 U17956 ( .B1(n14660), .B2(n20172), .A(n14659), .ZN(P1_U2980) );
  OAI21_X1 U17957 ( .B1(n14662), .B2(n14661), .A(n14651), .ZN(n15945) );
  INV_X1 U17958 ( .A(n14663), .ZN(n15816) );
  AOI22_X1 U17959 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n20190), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14664) );
  OAI21_X1 U17960 ( .B1(n20161), .B2(n15813), .A(n14664), .ZN(n14665) );
  AOI21_X1 U17961 ( .B1(n15816), .B2(n20167), .A(n14665), .ZN(n14666) );
  OAI21_X1 U17962 ( .B1(n20172), .B2(n15945), .A(n14666), .ZN(P1_U2981) );
  NAND2_X1 U17963 ( .A1(n10313), .A2(n14802), .ZN(n14671) );
  INV_X1 U17964 ( .A(n14668), .ZN(n14689) );
  AOI21_X1 U17965 ( .B1(n14788), .B2(n14805), .A(n14669), .ZN(n14670) );
  MUX2_X1 U17966 ( .A(n14671), .B(n10313), .S(n14670), .Z(n14673) );
  XNOR2_X1 U17967 ( .A(n14673), .B(n14672), .ZN(n15953) );
  INV_X1 U17968 ( .A(n14674), .ZN(n14678) );
  AOI22_X1 U17969 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n20190), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n14675) );
  OAI21_X1 U17970 ( .B1(n20161), .B2(n14676), .A(n14675), .ZN(n14677) );
  AOI21_X1 U17971 ( .B1(n14678), .B2(n20167), .A(n14677), .ZN(n14679) );
  OAI21_X1 U17972 ( .B1(n15953), .B2(n20172), .A(n14679), .ZN(P1_U2982) );
  OR2_X1 U17973 ( .A1(n14680), .A2(n14805), .ZN(n14789) );
  INV_X1 U17974 ( .A(n14681), .ZN(n14682) );
  NAND2_X1 U17975 ( .A1(n14789), .A2(n14682), .ZN(n14684) );
  AOI22_X1 U17976 ( .A1(n10313), .A2(n14790), .B1(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15883), .ZN(n14683) );
  XNOR2_X1 U17977 ( .A(n14684), .B(n14683), .ZN(n15963) );
  NAND2_X1 U17978 ( .A1(n15963), .A2(n20156), .ZN(n14687) );
  INV_X1 U17979 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15821) );
  NAND2_X1 U17980 ( .A1(n20190), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n15960) );
  OAI21_X1 U17981 ( .B1(n20165), .B2(n15821), .A(n15960), .ZN(n14685) );
  AOI21_X1 U17982 ( .B1(n15878), .B2(n15819), .A(n14685), .ZN(n14686) );
  OAI211_X1 U17983 ( .C1(n12495), .C2(n15820), .A(n14687), .B(n14686), .ZN(
        P1_U2984) );
  OR2_X1 U17984 ( .A1(n14667), .A2(n14688), .ZN(n15874) );
  AOI21_X1 U17985 ( .B1(n15874), .B2(n14689), .A(n15873), .ZN(n14691) );
  XNOR2_X1 U17986 ( .A(n14691), .B(n14690), .ZN(n15971) );
  NAND2_X1 U17987 ( .A1(n15971), .A2(n20156), .ZN(n14695) );
  NOR2_X1 U17988 ( .A1(n20170), .A2(n20811), .ZN(n15968) );
  NOR2_X1 U17989 ( .A1(n20161), .A2(n14692), .ZN(n14693) );
  AOI211_X1 U17990 ( .C1(n20152), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n15968), .B(n14693), .ZN(n14694) );
  OAI211_X1 U17991 ( .C1(n12495), .C2(n14696), .A(n14695), .B(n14694), .ZN(
        P1_U2986) );
  MUX2_X1 U17992 ( .A(n14697), .B(n14667), .S(n15883), .Z(n14698) );
  XOR2_X1 U17993 ( .A(n12391), .B(n14698), .Z(n16007) );
  INV_X1 U17994 ( .A(n16007), .ZN(n14704) );
  AOI22_X1 U17995 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20190), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14699) );
  OAI21_X1 U17996 ( .B1(n20161), .B2(n14700), .A(n14699), .ZN(n14701) );
  AOI21_X1 U17997 ( .B1(n14702), .B2(n20167), .A(n14701), .ZN(n14703) );
  OAI21_X1 U17998 ( .B1(n14704), .B2(n20172), .A(n14703), .ZN(P1_U2989) );
  NOR2_X1 U17999 ( .A1(n14706), .A2(n16014), .ZN(n14732) );
  INV_X1 U18000 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15981) );
  AND2_X1 U18001 ( .A1(n14708), .A2(n14707), .ZN(n15997) );
  NAND2_X1 U18002 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16003), .ZN(
        n16000) );
  NOR3_X1 U18003 ( .A1(n12391), .A2(n16019), .A3(n16000), .ZN(n14710) );
  NAND2_X1 U18004 ( .A1(n15997), .A2(n14710), .ZN(n15977) );
  NOR3_X1 U18005 ( .A1(n15981), .A2(n14804), .A3(n15977), .ZN(n14712) );
  INV_X1 U18006 ( .A(n14712), .ZN(n14786) );
  NOR2_X1 U18007 ( .A1(n14716), .A2(n14786), .ZN(n14711) );
  INV_X1 U18008 ( .A(n14709), .ZN(n16034) );
  AND2_X1 U18009 ( .A1(n14710), .A2(n16034), .ZN(n14803) );
  NAND2_X1 U18010 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14803), .ZN(
        n15978) );
  NOR2_X1 U18011 ( .A1(n14804), .A2(n15978), .ZN(n14783) );
  AOI22_X1 U18012 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n14711), .B1(
        n20185), .B2(n14783), .ZN(n15789) );
  OAI21_X1 U18013 ( .B1(n20199), .B2(n14786), .A(n15789), .ZN(n15970) );
  NAND3_X1 U18014 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n15970), .ZN(n15967) );
  NOR2_X1 U18015 ( .A1(n14790), .A2(n14802), .ZN(n15951) );
  NAND2_X1 U18016 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n15951), .ZN(
        n15943) );
  NOR2_X1 U18017 ( .A1(n15967), .A2(n15943), .ZN(n15948) );
  NAND2_X1 U18018 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15948), .ZN(
        n15942) );
  NOR2_X1 U18019 ( .A1(n15936), .A2(n15942), .ZN(n15792) );
  NAND2_X1 U18020 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15792), .ZN(
        n15771) );
  NAND2_X1 U18021 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15920) );
  NOR2_X1 U18022 ( .A1(n15771), .A2(n15920), .ZN(n15919) );
  NAND3_X1 U18023 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n15919), .ZN(n14767) );
  NAND2_X1 U18024 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14722) );
  NOR2_X1 U18025 ( .A1(n14767), .A2(n14722), .ZN(n14765) );
  NAND3_X1 U18026 ( .A1(n14765), .A2(n9920), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14738) );
  NOR3_X1 U18027 ( .A1(n14738), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14737), .ZN(n14731) );
  NOR4_X1 U18028 ( .A1(n15950), .A2(n12499), .A3(n12501), .A4(n15943), .ZN(
        n14713) );
  NAND2_X1 U18029 ( .A1(n14712), .A2(n14713), .ZN(n15788) );
  NAND2_X1 U18030 ( .A1(n14783), .A2(n14713), .ZN(n15784) );
  AOI211_X1 U18031 ( .C1(n15788), .C2(n15976), .A(n15921), .B(n15784), .ZN(
        n14714) );
  OAI21_X1 U18032 ( .B1(n14787), .B2(n14714), .A(n15980), .ZN(n15764) );
  AOI21_X1 U18033 ( .B1(n15920), .B2(n16001), .A(n15764), .ZN(n15934) );
  OAI21_X1 U18034 ( .B1(n14784), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15934), .ZN(n15922) );
  AND2_X1 U18035 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14715) );
  NOR2_X1 U18036 ( .A1(n14716), .A2(n14715), .ZN(n14717) );
  NOR2_X1 U18037 ( .A1(n15922), .A2(n14717), .ZN(n14728) );
  NAND2_X1 U18038 ( .A1(n15785), .A2(n14718), .ZN(n14719) );
  OAI21_X1 U18039 ( .B1(n14784), .B2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n14719), .ZN(n14720) );
  INV_X1 U18040 ( .A(n14720), .ZN(n14721) );
  NAND2_X1 U18041 ( .A1(n14728), .A2(n14721), .ZN(n15909) );
  AND2_X1 U18042 ( .A1(n16001), .A2(n14722), .ZN(n14723) );
  OR2_X1 U18043 ( .A1(n15909), .A2(n14723), .ZN(n14759) );
  AND2_X1 U18044 ( .A1(n16001), .A2(n14724), .ZN(n14725) );
  NOR2_X1 U18045 ( .A1(n14759), .A2(n14725), .ZN(n14744) );
  INV_X1 U18046 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14748) );
  AOI21_X1 U18047 ( .B1(n16001), .B2(n14748), .A(n14737), .ZN(n14726) );
  AND2_X1 U18048 ( .A1(n14744), .A2(n14726), .ZN(n14736) );
  AOI211_X1 U18049 ( .C1(n14787), .C2(n14728), .A(n14727), .B(n14736), .ZN(
        n14729) );
  NOR4_X1 U18050 ( .A1(n14732), .A2(n14731), .A3(n14730), .A4(n14729), .ZN(
        n14733) );
  OAI21_X1 U18051 ( .B1(n14734), .B2(n20208), .A(n14733), .ZN(P1_U3000) );
  INV_X1 U18052 ( .A(n14735), .ZN(n14741) );
  AOI21_X1 U18053 ( .B1(n14738), .B2(n14737), .A(n14736), .ZN(n14739) );
  AOI211_X1 U18054 ( .C1(n14741), .C2(n20203), .A(n14740), .B(n14739), .ZN(
        n14742) );
  OAI21_X1 U18055 ( .B1(n14743), .B2(n20208), .A(n14742), .ZN(P1_U3001) );
  NOR2_X1 U18056 ( .A1(n14744), .A2(n14748), .ZN(n14745) );
  AOI211_X1 U18057 ( .C1(n14747), .C2(n20203), .A(n14746), .B(n14745), .ZN(
        n14750) );
  NAND3_X1 U18058 ( .A1(n14765), .A2(n9920), .A3(n14748), .ZN(n14749) );
  OAI211_X1 U18059 ( .C1(n14751), .C2(n20208), .A(n14750), .B(n14749), .ZN(
        P1_U3002) );
  INV_X1 U18060 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14764) );
  XNOR2_X1 U18061 ( .A(n14764), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14757) );
  AOI21_X1 U18062 ( .B1(n14759), .B2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14752), .ZN(n14753) );
  OAI21_X1 U18063 ( .B1(n14754), .B2(n16014), .A(n14753), .ZN(n14756) );
  NOR2_X1 U18064 ( .A1(n20170), .A2(n20948), .ZN(n14758) );
  AOI21_X1 U18065 ( .B1(n14759), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14758), .ZN(n14760) );
  OAI21_X1 U18066 ( .B1(n14761), .B2(n16014), .A(n14760), .ZN(n14763) );
  NOR2_X1 U18067 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n14767), .ZN(
        n15908) );
  OAI21_X1 U18068 ( .B1(n15908), .B2(n15909), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14772) );
  INV_X1 U18069 ( .A(n14766), .ZN(n14770) );
  NOR3_X1 U18070 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n15910), .A3(
        n14767), .ZN(n14769) );
  INV_X1 U18071 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21013) );
  NOR2_X1 U18072 ( .A1(n20170), .A2(n21013), .ZN(n14768) );
  AOI211_X1 U18073 ( .C1(n14770), .C2(n20203), .A(n14769), .B(n14768), .ZN(
        n14771) );
  OAI211_X1 U18074 ( .C1(n14773), .C2(n20208), .A(n14772), .B(n14771), .ZN(
        P1_U3005) );
  NOR2_X1 U18075 ( .A1(n14774), .A2(n16014), .ZN(n14775) );
  AOI211_X1 U18076 ( .C1(n15764), .C2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n14776), .B(n14775), .ZN(n14781) );
  INV_X1 U18077 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14778) );
  INV_X1 U18078 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14777) );
  AOI21_X1 U18079 ( .B1(n14778), .B2(n14777), .A(n15771), .ZN(n14779) );
  NAND2_X1 U18080 ( .A1(n14779), .A2(n15920), .ZN(n14780) );
  OAI211_X1 U18081 ( .C1(n14782), .C2(n20208), .A(n14781), .B(n14780), .ZN(
        P1_U3009) );
  OAI221_X1 U18082 ( .B1(n14784), .B2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), 
        .C1(n14784), .C2(n14783), .A(n15980), .ZN(n14785) );
  AOI221_X1 U18083 ( .B1(n12499), .B2(n15976), .C1(n14786), .C2(n15976), .A(
        n14785), .ZN(n15974) );
  OAI21_X1 U18084 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n14787), .A(
        n15974), .ZN(n15964) );
  INV_X1 U18085 ( .A(n15964), .ZN(n14801) );
  NAND2_X1 U18086 ( .A1(n14789), .A2(n14788), .ZN(n14794) );
  NAND2_X1 U18087 ( .A1(n14790), .A2(n14802), .ZN(n14797) );
  AOI21_X1 U18088 ( .B1(n14797), .B2(n14794), .A(n14791), .ZN(n14792) );
  AOI21_X1 U18089 ( .B1(n14794), .B2(n14793), .A(n14792), .ZN(n15863) );
  NAND2_X1 U18090 ( .A1(n15863), .A2(n20188), .ZN(n14800) );
  NOR2_X1 U18091 ( .A1(n15951), .A2(n15967), .ZN(n14798) );
  OAI22_X1 U18092 ( .A1(n14795), .A2(n16014), .B1(n20170), .B2(n20817), .ZN(
        n14796) );
  AOI21_X1 U18093 ( .B1(n14798), .B2(n14797), .A(n14796), .ZN(n14799) );
  OAI211_X1 U18094 ( .C1(n14802), .C2(n14801), .A(n14800), .B(n14799), .ZN(
        P1_U3015) );
  INV_X1 U18095 ( .A(n15975), .ZN(n16033) );
  NAND2_X1 U18096 ( .A1(n14803), .A2(n16033), .ZN(n15996) );
  NOR4_X1 U18097 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n14804), .A3(
        n15981), .A4(n15996), .ZN(n14813) );
  INV_X1 U18098 ( .A(n14805), .ZN(n14808) );
  INV_X1 U18099 ( .A(n14806), .ZN(n14807) );
  AOI21_X1 U18100 ( .B1(n14809), .B2(n14808), .A(n14807), .ZN(n14811) );
  AOI22_X1 U18101 ( .A1(n10313), .A2(n12501), .B1(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15883), .ZN(n14810) );
  XNOR2_X1 U18102 ( .A(n14811), .B(n14810), .ZN(n15872) );
  OAI22_X1 U18103 ( .A1(n15974), .A2(n12501), .B1(n15872), .B2(n20208), .ZN(
        n14812) );
  AOI21_X1 U18104 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n14813), .A(
        n14812), .ZN(n14815) );
  NAND2_X1 U18105 ( .A1(n20190), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n14814) );
  OAI211_X1 U18106 ( .C1(n16014), .C2(n15829), .A(n14815), .B(n14814), .ZN(
        P1_U3017) );
  NAND2_X1 U18107 ( .A1(n20283), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20715) );
  XNOR2_X1 U18108 ( .A(n14816), .B(n20715), .ZN(n14818) );
  OAI22_X1 U18109 ( .A1(n14818), .A2(n20719), .B1(n10245), .B2(n14817), .ZN(
        n14819) );
  MUX2_X1 U18110 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n14819), .S(
        n20209), .Z(P1_U3476) );
  NAND2_X1 U18111 ( .A1(n14825), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14824) );
  NAND2_X1 U18112 ( .A1(n20250), .A2(n20732), .ZN(n14823) );
  INV_X1 U18113 ( .A(DATAI_18_), .ZN(n20959) );
  NOR2_X2 U18114 ( .A1(n20235), .A2(n14820), .ZN(n20733) );
  AOI22_X1 U18115 ( .A1(n20279), .A2(n20734), .B1(n20236), .B2(n20733), .ZN(
        n14822) );
  INV_X1 U18116 ( .A(DATAI_26_), .ZN(n21014) );
  NAND2_X1 U18117 ( .A1(n20759), .A2(n20684), .ZN(n14821) );
  NAND4_X1 U18118 ( .A1(n14824), .A2(n14823), .A3(n14822), .A4(n14821), .ZN(
        P1_U3035) );
  NAND2_X1 U18119 ( .A1(n14825), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14830) );
  NAND2_X1 U18120 ( .A1(n20261), .A2(n14826), .ZN(n20614) );
  INV_X1 U18121 ( .A(n20614), .ZN(n20744) );
  NAND2_X1 U18122 ( .A1(n20250), .A2(n20744), .ZN(n14829) );
  INV_X1 U18123 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16423) );
  OAI22_X1 U18124 ( .A1(n14523), .A2(n20247), .B1(n16423), .B2(n20248), .ZN(
        n20654) );
  NOR2_X2 U18125 ( .A1(n20235), .A2(n11612), .ZN(n20745) );
  AOI22_X1 U18126 ( .A1(n20279), .A2(n20654), .B1(n20236), .B2(n20745), .ZN(
        n14828) );
  INV_X1 U18127 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16413) );
  INV_X1 U18128 ( .A(DATAI_28_), .ZN(n20981) );
  OAI22_X2 U18129 ( .A1(n16413), .A2(n20248), .B1(n20981), .B2(n20247), .ZN(
        n20746) );
  NAND2_X1 U18130 ( .A1(n20759), .A2(n20746), .ZN(n14827) );
  NAND4_X1 U18131 ( .A1(n14830), .A2(n14829), .A3(n14828), .A4(n14827), .ZN(
        P1_U3037) );
  NAND4_X1 U18132 ( .A1(n16056), .A2(n19049), .A3(n14079), .A4(n15131), .ZN(
        n14840) );
  AOI22_X1 U18133 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n18996), .B1(
        P2_REIP_REG_31__SCAN_IN), .B2(n19054), .ZN(n14831) );
  INV_X1 U18134 ( .A(n14831), .ZN(n14838) );
  INV_X1 U18135 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n14833) );
  AOI22_X1 U18136 ( .A1(n12764), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n12871), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14832) );
  OAI21_X1 U18137 ( .B1(n12877), .B2(n14833), .A(n14832), .ZN(n14834) );
  INV_X1 U18138 ( .A(n14834), .ZN(n14835) );
  OAI22_X1 U18139 ( .A1(n15282), .A2(n19053), .B1(n12890), .B2(n14836), .ZN(
        n14837) );
  AOI211_X1 U18140 ( .C1(n15281), .C2(n19062), .A(n14838), .B(n14837), .ZN(
        n14839) );
  OAI211_X1 U18141 ( .C1(n9646), .C2(n14841), .A(n14840), .B(n14839), .ZN(
        P2_U2824) );
  AOI21_X1 U18142 ( .B1(n14843), .B2(n15153), .A(n14842), .ZN(n14844) );
  NAND2_X1 U18143 ( .A1(n14844), .A2(n19049), .ZN(n14855) );
  AND2_X1 U18144 ( .A1(n14846), .A2(n14845), .ZN(n14847) );
  NOR2_X1 U18145 ( .A1(n14936), .A2(n14847), .ZN(n15323) );
  INV_X1 U18146 ( .A(n15048), .ZN(n14850) );
  NAND2_X1 U18147 ( .A1(n9729), .A2(n14848), .ZN(n14849) );
  NAND2_X1 U18148 ( .A1(n14850), .A2(n14849), .ZN(n15321) );
  AOI22_X1 U18149 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19068), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19054), .ZN(n14852) );
  NAND2_X1 U18150 ( .A1(n19055), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n14851) );
  OAI211_X1 U18151 ( .C1(n15321), .C2(n19053), .A(n14852), .B(n14851), .ZN(
        n14853) );
  AOI21_X1 U18152 ( .B1(n15323), .B2(n19062), .A(n14853), .ZN(n14854) );
  OAI211_X1 U18153 ( .C1(n9646), .C2(n14856), .A(n14855), .B(n14854), .ZN(
        P2_U2827) );
  AOI211_X1 U18154 ( .C1(n14858), .C2(n15174), .A(n14857), .B(n19822), .ZN(
        n14859) );
  INV_X1 U18155 ( .A(n14859), .ZN(n14870) );
  OR2_X1 U18156 ( .A1(n9751), .A2(n14860), .ZN(n14861) );
  AND2_X1 U18157 ( .A1(n15070), .A2(n14861), .ZN(n15359) );
  AOI22_X1 U18158 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n19055), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19054), .ZN(n14862) );
  OAI21_X1 U18159 ( .B1(n14863), .B2(n19006), .A(n14862), .ZN(n14868) );
  OR2_X1 U18160 ( .A1(n14973), .A2(n14865), .ZN(n14866) );
  NAND2_X1 U18161 ( .A1(n14864), .A2(n14866), .ZN(n15362) );
  NOR2_X1 U18162 ( .A1(n15362), .A2(n19036), .ZN(n14867) );
  AOI211_X1 U18163 ( .C1(n15359), .C2(n19056), .A(n14868), .B(n14867), .ZN(
        n14869) );
  OAI211_X1 U18164 ( .C1(n9646), .C2(n14871), .A(n14870), .B(n14869), .ZN(
        P2_U2830) );
  AOI211_X1 U18165 ( .C1(n14874), .C2(n14873), .A(n14872), .B(n19822), .ZN(
        n14875) );
  INV_X1 U18166 ( .A(n14875), .ZN(n14888) );
  INV_X1 U18167 ( .A(n14877), .ZN(n14878) );
  AOI21_X1 U18168 ( .B1(n14879), .B2(n14876), .A(n14878), .ZN(n15432) );
  INV_X1 U18169 ( .A(n13260), .ZN(n14880) );
  OAI21_X1 U18170 ( .B1(n14882), .B2(n14881), .A(n14880), .ZN(n16096) );
  AOI22_X1 U18171 ( .A1(n19055), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19054), .ZN(n14883) );
  INV_X1 U18172 ( .A(n14883), .ZN(n14884) );
  AOI21_X1 U18173 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18996), .A(
        n14884), .ZN(n14885) );
  OAI21_X1 U18174 ( .B1(n16096), .B2(n19053), .A(n14885), .ZN(n14886) );
  AOI21_X1 U18175 ( .B1(n15432), .B2(n19062), .A(n14886), .ZN(n14887) );
  OAI211_X1 U18176 ( .C1(n9646), .C2(n14889), .A(n14888), .B(n14887), .ZN(
        P2_U2835) );
  AOI211_X1 U18177 ( .C1(n15243), .C2(n14891), .A(n14890), .B(n19822), .ZN(
        n14892) );
  INV_X1 U18178 ( .A(n14892), .ZN(n14902) );
  OR2_X1 U18179 ( .A1(n14909), .A2(n14893), .ZN(n14894) );
  NAND2_X1 U18180 ( .A1(n14876), .A2(n14894), .ZN(n15440) );
  INV_X1 U18181 ( .A(n15440), .ZN(n14900) );
  XNOR2_X1 U18182 ( .A(n14911), .B(n14895), .ZN(n15445) );
  AOI21_X1 U18183 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19068), .A(
        n19192), .ZN(n14896) );
  OAI21_X1 U18184 ( .B1(n19035), .B2(n19865), .A(n14896), .ZN(n14897) );
  AOI21_X1 U18185 ( .B1(n19055), .B2(P2_EBX_REG_19__SCAN_IN), .A(n14897), .ZN(
        n14898) );
  OAI21_X1 U18186 ( .B1(n15445), .B2(n19053), .A(n14898), .ZN(n14899) );
  AOI21_X1 U18187 ( .B1(n14900), .B2(n19062), .A(n14899), .ZN(n14901) );
  OAI211_X1 U18188 ( .C1(n9646), .C2(n14903), .A(n14902), .B(n14901), .ZN(
        P2_U2836) );
  AOI211_X1 U18189 ( .C1(n14906), .C2(n14905), .A(n14904), .B(n19822), .ZN(
        n14907) );
  INV_X1 U18190 ( .A(n14907), .ZN(n14920) );
  AND2_X1 U18191 ( .A1(n15013), .A2(n14908), .ZN(n14910) );
  OR2_X1 U18192 ( .A1(n14910), .A2(n14909), .ZN(n15010) );
  INV_X1 U18193 ( .A(n15010), .ZN(n16232) );
  INV_X1 U18194 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n14917) );
  NAND2_X1 U18195 ( .A1(n9786), .A2(n9758), .ZN(n14912) );
  AND2_X1 U18196 ( .A1(n14912), .A2(n14911), .ZN(n16228) );
  NAND2_X1 U18197 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18996), .ZN(
        n14913) );
  OAI211_X1 U18198 ( .C1(n19035), .C2(n14914), .A(n19033), .B(n14913), .ZN(
        n14915) );
  AOI21_X1 U18199 ( .B1(n19056), .B2(n16228), .A(n14915), .ZN(n14916) );
  OAI21_X1 U18200 ( .B1(n19017), .B2(n14917), .A(n14916), .ZN(n14918) );
  AOI21_X1 U18201 ( .B1(n16232), .B2(n19062), .A(n14918), .ZN(n14919) );
  OAI211_X1 U18202 ( .C1(n9646), .C2(n14921), .A(n14920), .B(n14919), .ZN(
        P2_U2837) );
  AOI21_X1 U18203 ( .B1(n14922), .B2(n15485), .A(n15113), .ZN(n19080) );
  NOR3_X1 U18204 ( .A1(n18993), .A2(n14923), .A3(n19822), .ZN(n18968) );
  AOI22_X1 U18205 ( .A1(n19080), .A2(n19056), .B1(n18968), .B2(n15248), .ZN(
        n14934) );
  NOR2_X1 U18206 ( .A1(n18993), .A2(n14923), .ZN(n14924) );
  NOR3_X1 U18207 ( .A1(n14924), .A2(n19822), .A3(n15248), .ZN(n14932) );
  OAI21_X1 U18208 ( .B1(n14925), .B2(n15030), .A(n15015), .ZN(n15466) );
  INV_X1 U18209 ( .A(n15466), .ZN(n15252) );
  INV_X1 U18210 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n14927) );
  AOI22_X1 U18211 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n19068), .B1(
        P2_REIP_REG_16__SCAN_IN), .B2(n19054), .ZN(n14926) );
  OAI211_X1 U18212 ( .C1(n19017), .C2(n14927), .A(n14926), .B(n19033), .ZN(
        n14928) );
  AOI21_X1 U18213 ( .B1(n19062), .B2(n15252), .A(n14928), .ZN(n14929) );
  OAI21_X1 U18214 ( .B1(n14930), .B2(n9646), .A(n14929), .ZN(n14931) );
  NOR2_X1 U18215 ( .A1(n14932), .A2(n14931), .ZN(n14933) );
  NAND2_X1 U18216 ( .A1(n14934), .A2(n14933), .ZN(P2_U2839) );
  MUX2_X1 U18217 ( .A(n15281), .B(P2_EBX_REG_31__SCAN_IN), .S(n14987), .Z(
        P2_U2856) );
  OR2_X1 U18218 ( .A1(n14936), .A2(n14935), .ZN(n14937) );
  INV_X1 U18219 ( .A(n14939), .ZN(n15046) );
  NAND2_X1 U18220 ( .A1(n14941), .A2(n14940), .ZN(n15045) );
  NAND3_X1 U18221 ( .A1(n15046), .A2(n15041), .A3(n15045), .ZN(n14943) );
  NAND2_X1 U18222 ( .A1(n14987), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14942) );
  OAI211_X1 U18223 ( .C1(n14987), .C2(n15308), .A(n14943), .B(n14942), .ZN(
        P2_U2858) );
  INV_X1 U18224 ( .A(n15323), .ZN(n14948) );
  NAND2_X1 U18225 ( .A1(n15058), .A2(n15041), .ZN(n14947) );
  NAND2_X1 U18226 ( .A1(n14987), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n14946) );
  OAI211_X1 U18227 ( .C1(n14948), .C2(n14987), .A(n14947), .B(n14946), .ZN(
        P2_U2859) );
  AOI21_X1 U18228 ( .B1(n14951), .B2(n14950), .A(n14949), .ZN(n15060) );
  NAND2_X1 U18229 ( .A1(n15060), .A2(n15041), .ZN(n14953) );
  NAND2_X1 U18230 ( .A1(n14987), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14952) );
  OAI211_X1 U18231 ( .C1(n15341), .C2(n14987), .A(n14953), .B(n14952), .ZN(
        P2_U2860) );
  NAND2_X1 U18232 ( .A1(n14864), .A2(n14954), .ZN(n14955) );
  NAND2_X1 U18233 ( .A1(n14956), .A2(n14955), .ZN(n16074) );
  AOI21_X1 U18234 ( .B1(n14959), .B2(n14958), .A(n14957), .ZN(n15067) );
  NAND2_X1 U18235 ( .A1(n15067), .A2(n15041), .ZN(n14961) );
  NAND2_X1 U18236 ( .A1(n14987), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14960) );
  OAI211_X1 U18237 ( .C1(n16074), .C2(n14987), .A(n14961), .B(n14960), .ZN(
        P2_U2861) );
  OAI21_X1 U18238 ( .B1(n14964), .B2(n14963), .A(n14962), .ZN(n15080) );
  NOR2_X1 U18239 ( .A1(n15362), .A2(n14987), .ZN(n14965) );
  AOI21_X1 U18240 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n14987), .A(n14965), .ZN(
        n14966) );
  OAI21_X1 U18241 ( .B1(n15080), .B2(n15019), .A(n14966), .ZN(P2_U2862) );
  AOI21_X1 U18242 ( .B1(n9755), .B2(n14968), .A(n14967), .ZN(n14969) );
  XOR2_X1 U18243 ( .A(n14970), .B(n14969), .Z(n15088) );
  AND2_X1 U18244 ( .A1(n14972), .A2(n14971), .ZN(n14974) );
  OR2_X1 U18245 ( .A1(n14974), .A2(n14973), .ZN(n16086) );
  NOR2_X1 U18246 ( .A1(n16086), .A2(n14987), .ZN(n14975) );
  AOI21_X1 U18247 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n14987), .A(n14975), .ZN(
        n14976) );
  OAI21_X1 U18248 ( .B1(n15088), .B2(n15019), .A(n14976), .ZN(P2_U2863) );
  AOI21_X1 U18249 ( .B1(n14980), .B2(n14979), .A(n14978), .ZN(n14981) );
  INV_X1 U18250 ( .A(n14981), .ZN(n15094) );
  MUX2_X1 U18251 ( .A(n14982), .B(n15189), .S(n15036), .Z(n14983) );
  OAI21_X1 U18252 ( .B1(n15094), .B2(n15019), .A(n14983), .ZN(P2_U2864) );
  OAI21_X1 U18253 ( .B1(n14984), .B2(n14986), .A(n14985), .ZN(n15100) );
  NAND2_X1 U18254 ( .A1(n14987), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n14989) );
  NAND2_X1 U18255 ( .A1(n16108), .A2(n15036), .ZN(n14988) );
  OAI211_X1 U18256 ( .C1(n15100), .C2(n15019), .A(n14989), .B(n14988), .ZN(
        P2_U2865) );
  AOI21_X1 U18257 ( .B1(n14991), .B2(n14990), .A(n14984), .ZN(n15101) );
  NAND2_X1 U18258 ( .A1(n15101), .A2(n15041), .ZN(n14993) );
  NAND2_X1 U18259 ( .A1(n14987), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n14992) );
  OAI211_X1 U18260 ( .C1(n15414), .C2(n14987), .A(n14993), .B(n14992), .ZN(
        P2_U2866) );
  INV_X1 U18261 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n14999) );
  INV_X1 U18262 ( .A(n14990), .ZN(n14995) );
  AOI21_X1 U18263 ( .B1(n14996), .B2(n14994), .A(n14995), .ZN(n16098) );
  NAND2_X1 U18264 ( .A1(n16098), .A2(n15041), .ZN(n14998) );
  NAND2_X1 U18265 ( .A1(n15432), .A2(n15036), .ZN(n14997) );
  OAI211_X1 U18266 ( .C1(n15036), .C2(n14999), .A(n14998), .B(n14997), .ZN(
        P2_U2867) );
  AND2_X1 U18267 ( .A1(n15004), .A2(n15000), .ZN(n15006) );
  OAI21_X1 U18268 ( .B1(n15006), .B2(n15001), .A(n14994), .ZN(n15112) );
  NOR2_X1 U18269 ( .A1(n15440), .A2(n14987), .ZN(n15002) );
  AOI21_X1 U18270 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n14987), .A(n15002), .ZN(
        n15003) );
  OAI21_X1 U18271 ( .B1(n15112), .B2(n15019), .A(n15003), .ZN(P2_U2868) );
  INV_X1 U18272 ( .A(n15004), .ZN(n15027) );
  AOI21_X1 U18273 ( .B1(n15007), .B2(n10296), .A(n15006), .ZN(n16103) );
  NAND2_X1 U18274 ( .A1(n16103), .A2(n15041), .ZN(n15009) );
  NAND2_X1 U18275 ( .A1(n14987), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n15008) );
  OAI211_X1 U18276 ( .C1(n15010), .C2(n14987), .A(n15009), .B(n15008), .ZN(
        P2_U2869) );
  OR2_X1 U18277 ( .A1(n15027), .A2(n15020), .ZN(n15022) );
  INV_X1 U18278 ( .A(n15022), .ZN(n15012) );
  OAI21_X1 U18279 ( .B1(n15012), .B2(n15011), .A(n10296), .ZN(n15121) );
  NAND2_X1 U18280 ( .A1(n14987), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15018) );
  INV_X1 U18281 ( .A(n15013), .ZN(n15014) );
  AOI21_X1 U18282 ( .B1(n15016), .B2(n15015), .A(n15014), .ZN(n18950) );
  NAND2_X1 U18283 ( .A1(n18950), .A2(n15036), .ZN(n15017) );
  OAI211_X1 U18284 ( .C1(n15121), .C2(n15019), .A(n15018), .B(n15017), .ZN(
        P2_U2870) );
  NAND2_X1 U18285 ( .A1(n15027), .A2(n15020), .ZN(n15021) );
  AND2_X1 U18286 ( .A1(n15022), .A2(n15021), .ZN(n19081) );
  NAND2_X1 U18287 ( .A1(n19081), .A2(n15041), .ZN(n15024) );
  NAND2_X1 U18288 ( .A1(n14987), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n15023) );
  OAI211_X1 U18289 ( .C1(n15466), .C2(n14987), .A(n15024), .B(n15023), .ZN(
        P2_U2871) );
  INV_X1 U18290 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n15035) );
  OAI211_X1 U18291 ( .C1(n15040), .C2(n15028), .A(n15027), .B(n15041), .ZN(
        n15034) );
  NAND2_X1 U18292 ( .A1(n15029), .A2(n15038), .ZN(n15032) );
  INV_X1 U18293 ( .A(n15030), .ZN(n15031) );
  NAND2_X1 U18294 ( .A1(n15036), .A2(n18957), .ZN(n15033) );
  OAI211_X1 U18295 ( .C1(n15036), .C2(n15035), .A(n15034), .B(n15033), .ZN(
        P2_U2872) );
  OR2_X1 U18296 ( .A1(n15037), .A2(n14171), .ZN(n15039) );
  NAND2_X1 U18297 ( .A1(n15039), .A2(n15038), .ZN(n16140) );
  OAI211_X1 U18298 ( .C1(n14165), .C2(n15042), .A(n15026), .B(n15041), .ZN(
        n15044) );
  NAND2_X1 U18299 ( .A1(n14987), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n15043) );
  OAI211_X1 U18300 ( .C1(n16140), .C2(n14987), .A(n15044), .B(n15043), .ZN(
        P2_U2873) );
  NAND3_X1 U18301 ( .A1(n15046), .A2(n19085), .A3(n15045), .ZN(n15054) );
  OR2_X1 U18302 ( .A1(n15048), .A2(n15047), .ZN(n15049) );
  NAND2_X1 U18303 ( .A1(n9730), .A2(n15049), .ZN(n16068) );
  INV_X1 U18304 ( .A(n16068), .ZN(n15310) );
  OAI22_X1 U18305 ( .A1(n15116), .A2(n19092), .B1(n19121), .B2(n15050), .ZN(
        n15051) );
  AOI21_X1 U18306 ( .B1(n19131), .B2(n15310), .A(n15051), .ZN(n15053) );
  AOI22_X1 U18307 ( .A1(n19079), .A2(BUF1_REG_29__SCAN_IN), .B1(n19078), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n15052) );
  NAND3_X1 U18308 ( .A1(n15054), .A2(n15053), .A3(n15052), .ZN(P2_U2890) );
  AOI22_X1 U18309 ( .A1(n19079), .A2(BUF1_REG_28__SCAN_IN), .B1(n19078), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n15056) );
  AOI22_X1 U18310 ( .A1(n19077), .A2(n19095), .B1(n19130), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n15055) );
  OAI211_X1 U18311 ( .C1(n19122), .C2(n15321), .A(n15056), .B(n15055), .ZN(
        n15057) );
  AOI21_X1 U18312 ( .B1(n15058), .B2(n19085), .A(n15057), .ZN(n15059) );
  INV_X1 U18313 ( .A(n15059), .ZN(P2_U2891) );
  INV_X1 U18314 ( .A(n15060), .ZN(n15066) );
  INV_X1 U18315 ( .A(n15061), .ZN(n15338) );
  OAI22_X1 U18316 ( .A1(n15116), .A2(n19098), .B1(n19121), .B2(n15062), .ZN(
        n15063) );
  AOI21_X1 U18317 ( .B1(n19131), .B2(n15338), .A(n15063), .ZN(n15065) );
  AOI22_X1 U18318 ( .A1(n19079), .A2(BUF1_REG_27__SCAN_IN), .B1(n19078), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n15064) );
  OAI211_X1 U18319 ( .C1(n15066), .C2(n19135), .A(n15065), .B(n15064), .ZN(
        P2_U2892) );
  NAND2_X1 U18320 ( .A1(n15067), .A2(n19085), .ZN(n15075) );
  AOI22_X1 U18321 ( .A1(n19077), .A2(n19101), .B1(n19130), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15074) );
  AOI22_X1 U18322 ( .A1(n19079), .A2(BUF1_REG_26__SCAN_IN), .B1(n19078), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n15073) );
  INV_X1 U18323 ( .A(n15068), .ZN(n15069) );
  AOI21_X1 U18324 ( .B1(n15071), .B2(n15070), .A(n15069), .ZN(n16081) );
  NAND2_X1 U18325 ( .A1(n19131), .A2(n16081), .ZN(n15072) );
  NAND4_X1 U18326 ( .A1(n15075), .A2(n15074), .A3(n15073), .A4(n15072), .ZN(
        P2_U2893) );
  OAI22_X1 U18327 ( .A1(n15116), .A2(n19104), .B1(n19121), .B2(n15076), .ZN(
        n15077) );
  AOI21_X1 U18328 ( .B1(n19131), .B2(n15359), .A(n15077), .ZN(n15079) );
  AOI22_X1 U18329 ( .A1(n19079), .A2(BUF1_REG_25__SCAN_IN), .B1(n19078), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n15078) );
  OAI211_X1 U18330 ( .C1(n15080), .C2(n19135), .A(n15079), .B(n15078), .ZN(
        P2_U2894) );
  AND2_X1 U18331 ( .A1(n15082), .A2(n15081), .ZN(n15083) );
  OR2_X1 U18332 ( .A1(n15083), .A2(n9751), .ZN(n16085) );
  AOI22_X1 U18333 ( .A1(n19079), .A2(BUF1_REG_24__SCAN_IN), .B1(n19078), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n15085) );
  AOI22_X1 U18334 ( .A1(n19077), .A2(n19108), .B1(n19130), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n15084) );
  OAI211_X1 U18335 ( .C1(n19122), .C2(n16085), .A(n15085), .B(n15084), .ZN(
        n15086) );
  INV_X1 U18336 ( .A(n15086), .ZN(n15087) );
  OAI21_X1 U18337 ( .B1(n15088), .B2(n19135), .A(n15087), .ZN(P2_U2895) );
  INV_X1 U18338 ( .A(n15384), .ZN(n15091) );
  OAI22_X1 U18339 ( .A1(n15116), .A2(n19264), .B1(n19121), .B2(n15089), .ZN(
        n15090) );
  AOI21_X1 U18340 ( .B1(n19131), .B2(n15091), .A(n15090), .ZN(n15093) );
  AOI22_X1 U18341 ( .A1(n19079), .A2(BUF1_REG_23__SCAN_IN), .B1(n19078), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n15092) );
  OAI211_X1 U18342 ( .C1(n15094), .C2(n19135), .A(n15093), .B(n15092), .ZN(
        P2_U2896) );
  INV_X1 U18343 ( .A(n15400), .ZN(n15097) );
  OAI22_X1 U18344 ( .A1(n15116), .A2(n19255), .B1(n19121), .B2(n15095), .ZN(
        n15096) );
  AOI21_X1 U18345 ( .B1(n19131), .B2(n15097), .A(n15096), .ZN(n15099) );
  AOI22_X1 U18346 ( .A1(n19079), .A2(BUF1_REG_22__SCAN_IN), .B1(n19078), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n15098) );
  OAI211_X1 U18347 ( .C1(n15100), .C2(n19135), .A(n15099), .B(n15098), .ZN(
        P2_U2897) );
  INV_X1 U18348 ( .A(n15101), .ZN(n15106) );
  OAI22_X1 U18349 ( .A1(n15116), .A2(n19252), .B1(n19121), .B2(n15102), .ZN(
        n15103) );
  AOI21_X1 U18350 ( .B1(n19131), .B2(n15419), .A(n15103), .ZN(n15105) );
  AOI22_X1 U18351 ( .A1(n19079), .A2(BUF1_REG_21__SCAN_IN), .B1(n19078), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n15104) );
  OAI211_X1 U18352 ( .C1(n15106), .C2(n19135), .A(n15105), .B(n15104), .ZN(
        P2_U2898) );
  INV_X1 U18353 ( .A(n15445), .ZN(n15109) );
  OAI22_X1 U18354 ( .A1(n15116), .A2(n19243), .B1(n19121), .B2(n15107), .ZN(
        n15108) );
  AOI21_X1 U18355 ( .B1(n19131), .B2(n15109), .A(n15108), .ZN(n15111) );
  AOI22_X1 U18356 ( .A1(n19079), .A2(BUF1_REG_19__SCAN_IN), .B1(n19078), .B2(
        BUF2_REG_19__SCAN_IN), .ZN(n15110) );
  OAI211_X1 U18357 ( .C1(n15112), .C2(n19135), .A(n15111), .B(n15110), .ZN(
        P2_U2900) );
  OAI21_X1 U18358 ( .B1(n15114), .B2(n15113), .A(n9758), .ZN(n18954) );
  INV_X1 U18359 ( .A(n18954), .ZN(n15118) );
  OAI22_X1 U18360 ( .A1(n15116), .A2(n19233), .B1(n19121), .B2(n15115), .ZN(
        n15117) );
  AOI21_X1 U18361 ( .B1(n19131), .B2(n15118), .A(n15117), .ZN(n15120) );
  AOI22_X1 U18362 ( .A1(n19079), .A2(BUF1_REG_17__SCAN_IN), .B1(n19078), .B2(
        BUF2_REG_17__SCAN_IN), .ZN(n15119) );
  OAI211_X1 U18363 ( .C1(n15121), .C2(n19135), .A(n15120), .B(n15119), .ZN(
        P2_U2902) );
  NAND2_X1 U18364 ( .A1(n15122), .A2(n15135), .ZN(n15127) );
  INV_X1 U18365 ( .A(n15123), .ZN(n15124) );
  NOR2_X1 U18366 ( .A1(n15125), .A2(n15124), .ZN(n15126) );
  XNOR2_X1 U18367 ( .A(n15127), .B(n15126), .ZN(n15307) );
  XOR2_X1 U18368 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n15138), .Z(
        n15305) );
  NAND2_X1 U18369 ( .A1(n19192), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15299) );
  OAI21_X1 U18370 ( .B1(n16227), .B2(n15128), .A(n15299), .ZN(n15129) );
  AOI21_X1 U18371 ( .B1(n15301), .B2(n19194), .A(n15129), .ZN(n15130) );
  OAI21_X1 U18372 ( .B1(n15131), .B2(n19182), .A(n15130), .ZN(n15132) );
  AOI21_X1 U18373 ( .B1(n15305), .B2(n11014), .A(n15132), .ZN(n15133) );
  OAI21_X1 U18374 ( .B1(n15307), .B2(n16209), .A(n15133), .ZN(P2_U2984) );
  NAND2_X1 U18375 ( .A1(n15135), .A2(n15134), .ZN(n15137) );
  XOR2_X1 U18376 ( .A(n15137), .B(n15136), .Z(n15318) );
  AOI21_X1 U18377 ( .B1(n15314), .B2(n15150), .A(n15138), .ZN(n15316) );
  NOR2_X1 U18378 ( .A1(n19033), .A2(n19882), .ZN(n15309) );
  NOR2_X1 U18379 ( .A1(n15308), .A2(n19218), .ZN(n15139) );
  AOI211_X1 U18380 ( .C1(n19187), .C2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15309), .B(n15139), .ZN(n15140) );
  OAI21_X1 U18381 ( .B1(n19182), .B2(n15141), .A(n15140), .ZN(n15142) );
  AOI21_X1 U18382 ( .B1(n15316), .B2(n11014), .A(n15142), .ZN(n15143) );
  OAI21_X1 U18383 ( .B1(n15318), .B2(n16209), .A(n15143), .ZN(P2_U2985) );
  XNOR2_X1 U18384 ( .A(n15145), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15146) );
  XNOR2_X1 U18385 ( .A(n15147), .B(n15146), .ZN(n15332) );
  NAND2_X1 U18386 ( .A1(n15323), .A2(n19194), .ZN(n15148) );
  NAND2_X1 U18387 ( .A1(n19192), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15320) );
  OAI211_X1 U18388 ( .C1(n16227), .C2(n15149), .A(n15148), .B(n15320), .ZN(
        n15152) );
  NOR2_X1 U18389 ( .A1(n15319), .A2(n16207), .ZN(n15151) );
  AOI211_X1 U18390 ( .C1(n19195), .C2(n15153), .A(n15152), .B(n15151), .ZN(
        n15154) );
  OAI21_X1 U18391 ( .B1(n15332), .B2(n16209), .A(n15154), .ZN(P2_U2986) );
  XNOR2_X1 U18392 ( .A(n15155), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15346) );
  NAND2_X1 U18393 ( .A1(n19192), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15336) );
  NAND2_X1 U18394 ( .A1(n19187), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15156) );
  OAI211_X1 U18395 ( .C1(n15341), .C2(n19218), .A(n15336), .B(n15156), .ZN(
        n15158) );
  NOR2_X1 U18396 ( .A1(n9882), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15334) );
  NOR3_X1 U18397 ( .A1(n15334), .A2(n15333), .A3(n16207), .ZN(n15157) );
  AOI211_X1 U18398 ( .C1(n19195), .C2(n15159), .A(n15158), .B(n15157), .ZN(
        n15160) );
  OAI21_X1 U18399 ( .B1(n15346), .B2(n16209), .A(n15160), .ZN(P2_U2987) );
  OAI21_X1 U18400 ( .B1(n15175), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15161), .ZN(n15358) );
  AOI21_X1 U18401 ( .B1(n15162), .B2(n15170), .A(n15169), .ZN(n15164) );
  XNOR2_X1 U18402 ( .A(n15164), .B(n15163), .ZN(n15347) );
  NAND2_X1 U18403 ( .A1(n15347), .A2(n19188), .ZN(n15168) );
  NAND2_X1 U18404 ( .A1(n19192), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15352) );
  NAND2_X1 U18405 ( .A1(n19187), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15165) );
  OAI211_X1 U18406 ( .C1(n16074), .C2(n19218), .A(n15352), .B(n15165), .ZN(
        n15166) );
  AOI21_X1 U18407 ( .B1(n16071), .B2(n19195), .A(n15166), .ZN(n15167) );
  OAI211_X1 U18408 ( .C1(n16207), .C2(n15358), .A(n15168), .B(n15167), .ZN(
        P2_U2988) );
  NAND2_X1 U18409 ( .A1(n10926), .A2(n15170), .ZN(n15171) );
  XNOR2_X1 U18410 ( .A(n15162), .B(n15171), .ZN(n15370) );
  NAND2_X1 U18411 ( .A1(n19192), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15361) );
  NAND2_X1 U18412 ( .A1(n19187), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15172) );
  OAI211_X1 U18413 ( .C1(n15362), .C2(n19218), .A(n15361), .B(n15172), .ZN(
        n15173) );
  AOI21_X1 U18414 ( .B1(n15174), .B2(n19195), .A(n15173), .ZN(n15177) );
  AOI21_X1 U18415 ( .B1(n15365), .B2(n15178), .A(n15175), .ZN(n15367) );
  NAND2_X1 U18416 ( .A1(n15367), .A2(n11014), .ZN(n15176) );
  OAI211_X1 U18417 ( .C1(n15370), .C2(n16209), .A(n15177), .B(n15176), .ZN(
        P2_U2989) );
  OAI21_X1 U18418 ( .B1(n15193), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15178), .ZN(n15381) );
  XOR2_X1 U18419 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n15179), .Z(
        n15180) );
  XNOR2_X1 U18420 ( .A(n15181), .B(n15180), .ZN(n15371) );
  NAND2_X1 U18421 ( .A1(n15371), .A2(n19188), .ZN(n15185) );
  NAND2_X1 U18422 ( .A1(n19192), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n15372) );
  NAND2_X1 U18423 ( .A1(n19187), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15182) );
  OAI211_X1 U18424 ( .C1(n16086), .C2(n19218), .A(n15372), .B(n15182), .ZN(
        n15183) );
  AOI21_X1 U18425 ( .B1(n16089), .B2(n19195), .A(n15183), .ZN(n15184) );
  OAI211_X1 U18426 ( .C1(n15381), .C2(n16207), .A(n15185), .B(n15184), .ZN(
        P2_U2990) );
  XNOR2_X1 U18427 ( .A(n15186), .B(n15187), .ZN(n15392) );
  OAI22_X1 U18428 ( .A1(n16227), .A2(n15188), .B1(n19872), .B2(n19033), .ZN(
        n15191) );
  NOR2_X1 U18429 ( .A1(n15189), .A2(n19218), .ZN(n15190) );
  AOI211_X1 U18430 ( .C1(n15192), .C2(n19195), .A(n15191), .B(n15190), .ZN(
        n15195) );
  AOI21_X1 U18431 ( .B1(n15388), .B2(n15398), .A(n15193), .ZN(n15390) );
  NAND2_X1 U18432 ( .A1(n15390), .A2(n11014), .ZN(n15194) );
  OAI211_X1 U18433 ( .C1(n15392), .C2(n16209), .A(n15195), .B(n15194), .ZN(
        P2_U2991) );
  AND2_X1 U18434 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15196), .ZN(
        n15426) );
  NAND2_X1 U18435 ( .A1(n16121), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15235) );
  NOR2_X1 U18436 ( .A1(n15235), .A2(n15232), .ZN(n15231) );
  INV_X1 U18437 ( .A(n15284), .ZN(n15197) );
  NAND2_X1 U18438 ( .A1(n15534), .A2(n15197), .ZN(n15397) );
  OAI21_X1 U18439 ( .B1(n15231), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15397), .ZN(n15422) );
  NAND2_X1 U18440 ( .A1(n15199), .A2(n15198), .ZN(n15214) );
  NOR2_X1 U18441 ( .A1(n15201), .A2(n9903), .ZN(n15204) );
  NAND3_X1 U18442 ( .A1(n15511), .A2(n15202), .A3(n10852), .ZN(n15203) );
  OAI211_X1 U18443 ( .C1(n15204), .C2(n15203), .A(n10857), .B(n15477), .ZN(
        n15206) );
  AOI21_X1 U18444 ( .B1(n15206), .B2(n15205), .A(n15473), .ZN(n15247) );
  INV_X1 U18445 ( .A(n15247), .ZN(n15209) );
  INV_X1 U18446 ( .A(n15246), .ZN(n15208) );
  NAND2_X1 U18447 ( .A1(n15211), .A2(n15210), .ZN(n15453) );
  NAND3_X1 U18448 ( .A1(n16115), .A2(n15237), .A3(n16113), .ZN(n15222) );
  AOI21_X1 U18449 ( .B1(n15222), .B2(n15212), .A(n15223), .ZN(n15213) );
  XOR2_X1 U18450 ( .A(n15214), .B(n15213), .Z(n15410) );
  NAND2_X1 U18451 ( .A1(n15410), .A2(n19188), .ZN(n15220) );
  NAND2_X1 U18452 ( .A1(n19192), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15413) );
  OAI21_X1 U18453 ( .B1(n16227), .B2(n15215), .A(n15413), .ZN(n15217) );
  NOR2_X1 U18454 ( .A1(n15414), .A2(n19218), .ZN(n15216) );
  AOI211_X1 U18455 ( .C1(n19195), .C2(n15218), .A(n15217), .B(n15216), .ZN(
        n15219) );
  OAI211_X1 U18456 ( .C1(n16207), .C2(n15422), .A(n15220), .B(n15219), .ZN(
        P2_U2993) );
  NAND2_X1 U18457 ( .A1(n15222), .A2(n15221), .ZN(n15227) );
  INV_X1 U18458 ( .A(n15223), .ZN(n15225) );
  NAND2_X1 U18459 ( .A1(n15225), .A2(n15224), .ZN(n15226) );
  XNOR2_X1 U18460 ( .A(n15227), .B(n15226), .ZN(n15438) );
  NAND2_X1 U18461 ( .A1(n19192), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n15428) );
  NAND2_X1 U18462 ( .A1(n19187), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15228) );
  OAI211_X1 U18463 ( .C1(n19182), .C2(n15229), .A(n15428), .B(n15228), .ZN(
        n15230) );
  AOI21_X1 U18464 ( .B1(n19194), .B2(n15432), .A(n15230), .ZN(n15234) );
  AOI21_X1 U18465 ( .B1(n15232), .B2(n15235), .A(n15231), .ZN(n15436) );
  NAND2_X1 U18466 ( .A1(n15436), .A2(n11014), .ZN(n15233) );
  OAI211_X1 U18467 ( .C1(n15438), .C2(n16209), .A(n15234), .B(n15233), .ZN(
        P2_U2994) );
  OAI21_X1 U18468 ( .B1(n16121), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15235), .ZN(n15451) );
  NAND2_X1 U18469 ( .A1(n15237), .A2(n15236), .ZN(n15239) );
  NAND2_X1 U18470 ( .A1(n16115), .A2(n16113), .ZN(n16118) );
  NAND2_X1 U18471 ( .A1(n16118), .A2(n16114), .ZN(n15238) );
  XOR2_X1 U18472 ( .A(n15239), .B(n15238), .Z(n15439) );
  NAND2_X1 U18473 ( .A1(n15439), .A2(n19188), .ZN(n15245) );
  NAND2_X1 U18474 ( .A1(n19192), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15444) );
  OAI21_X1 U18475 ( .B1(n16227), .B2(n15240), .A(n15444), .ZN(n15242) );
  NOR2_X1 U18476 ( .A1(n19218), .A2(n15440), .ZN(n15241) );
  AOI211_X1 U18477 ( .C1(n19195), .C2(n15243), .A(n15242), .B(n15241), .ZN(
        n15244) );
  OAI211_X1 U18478 ( .C1(n16207), .C2(n15451), .A(n15245), .B(n15244), .ZN(
        P2_U2995) );
  XNOR2_X1 U18479 ( .A(n15247), .B(n15246), .ZN(n15471) );
  NOR2_X1 U18480 ( .A1(n12843), .A2(n19033), .ZN(n15251) );
  INV_X1 U18481 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15249) );
  OAI22_X1 U18482 ( .A1(n16227), .A2(n15249), .B1(n19182), .B2(n15248), .ZN(
        n15250) );
  AOI211_X1 U18483 ( .C1(n19194), .C2(n15252), .A(n15251), .B(n15250), .ZN(
        n15255) );
  NAND2_X1 U18484 ( .A1(n15492), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16120) );
  XNOR2_X1 U18485 ( .A(n16120), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15253) );
  NAND2_X1 U18486 ( .A1(n15253), .A2(n11014), .ZN(n15254) );
  OAI211_X1 U18487 ( .C1(n15471), .C2(n16209), .A(n15255), .B(n15254), .ZN(
        P2_U2998) );
  XNOR2_X1 U18488 ( .A(n15256), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15257) );
  XNOR2_X1 U18489 ( .A(n15258), .B(n15257), .ZN(n16300) );
  INV_X1 U18490 ( .A(n16195), .ZN(n15263) );
  OAI21_X1 U18491 ( .B1(n15261), .B2(n15263), .A(n15260), .ZN(n15262) );
  OAI21_X1 U18492 ( .B1(n15259), .B2(n15263), .A(n15262), .ZN(n16297) );
  OAI22_X1 U18493 ( .A1(n16227), .A2(n15264), .B1(n19848), .B2(n19033), .ZN(
        n15267) );
  INV_X1 U18494 ( .A(n19029), .ZN(n15265) );
  OAI22_X1 U18495 ( .A1(n19182), .A2(n15265), .B1(n19218), .B2(n19037), .ZN(
        n15266) );
  AOI211_X1 U18496 ( .C1(n16297), .C2(n19188), .A(n15267), .B(n15266), .ZN(
        n15268) );
  OAI21_X1 U18497 ( .B1(n16207), .B2(n16300), .A(n15268), .ZN(P2_U3007) );
  XNOR2_X1 U18498 ( .A(n15269), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15556) );
  XOR2_X1 U18499 ( .A(n15270), .B(n15271), .Z(n15554) );
  OAI22_X1 U18500 ( .A1(n19846), .A2(n19033), .B1(n19182), .B2(n15272), .ZN(
        n15275) );
  INV_X1 U18501 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n15273) );
  OAI22_X1 U18502 ( .A1(n19218), .A2(n15551), .B1(n16227), .B2(n15273), .ZN(
        n15274) );
  AOI211_X1 U18503 ( .C1(n15554), .C2(n19188), .A(n15275), .B(n15274), .ZN(
        n15276) );
  OAI21_X1 U18504 ( .B1(n15556), .B2(n16207), .A(n15276), .ZN(P2_U3008) );
  NAND3_X1 U18505 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15288) );
  NAND2_X1 U18506 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16284) );
  INV_X1 U18507 ( .A(n16284), .ZN(n15283) );
  NAND3_X1 U18508 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n16312), .ZN(n15545) );
  NOR2_X1 U18509 ( .A1(n15548), .A2(n15545), .ZN(n16278) );
  NAND2_X1 U18510 ( .A1(n15283), .A2(n16278), .ZN(n16258) );
  OAI21_X1 U18511 ( .B1(n16258), .B2(n15284), .A(n16257), .ZN(n15416) );
  NAND2_X1 U18512 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15285) );
  NAND2_X1 U18513 ( .A1(n16257), .A2(n15285), .ZN(n15277) );
  NAND2_X1 U18514 ( .A1(n15416), .A2(n15277), .ZN(n15349) );
  NAND3_X1 U18515 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15278) );
  AND2_X1 U18516 ( .A1(n16257), .A2(n15278), .ZN(n15279) );
  OR2_X1 U18517 ( .A1(n15349), .A2(n15279), .ZN(n15335) );
  AOI211_X1 U18518 ( .C1(n16257), .C2(n15288), .A(n15280), .B(n15335), .ZN(
        n15303) );
  NOR3_X1 U18519 ( .A1(n15303), .A2(n16277), .A3(n15289), .ZN(n15295) );
  INV_X1 U18520 ( .A(n15281), .ZN(n15294) );
  INV_X1 U18521 ( .A(n15282), .ZN(n19073) );
  NAND3_X1 U18522 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n15560), .ZN(n15549) );
  NAND2_X1 U18523 ( .A1(n16294), .A2(n15283), .ZN(n15535) );
  NOR2_X1 U18524 ( .A1(n15284), .A2(n15535), .ZN(n15404) );
  INV_X1 U18525 ( .A(n15285), .ZN(n15286) );
  NAND2_X1 U18526 ( .A1(n15404), .A2(n15286), .ZN(n15375) );
  NAND2_X1 U18527 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15287) );
  NOR2_X1 U18528 ( .A1(n15348), .A2(n15287), .ZN(n15324) );
  INV_X1 U18529 ( .A(n15288), .ZN(n15298) );
  NAND4_X1 U18530 ( .A1(n15324), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15298), .A4(n15289), .ZN(n15292) );
  INV_X1 U18531 ( .A(n15290), .ZN(n15291) );
  AOI21_X1 U18532 ( .B1(n15324), .B2(n15298), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15302) );
  AOI21_X1 U18533 ( .B1(n15305), .B2(n19204), .A(n15304), .ZN(n15306) );
  OAI21_X1 U18534 ( .B1(n15307), .B2(n19209), .A(n15306), .ZN(P2_U3016) );
  AND2_X1 U18535 ( .A1(n15324), .A2(n15311), .ZN(n15343) );
  NOR2_X1 U18536 ( .A1(n15343), .A2(n15335), .ZN(n15328) );
  OAI21_X1 U18537 ( .B1(n15311), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15312) );
  OAI211_X1 U18538 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(n15324), .B(n15312), .ZN(
        n15313) );
  AOI21_X1 U18539 ( .B1(n15316), .B2(n19204), .A(n15315), .ZN(n15317) );
  OAI21_X1 U18540 ( .B1(n15318), .B2(n19209), .A(n15317), .ZN(P2_U3017) );
  INV_X1 U18541 ( .A(n15319), .ZN(n15330) );
  OAI21_X1 U18542 ( .B1(n16306), .B2(n15321), .A(n15320), .ZN(n15322) );
  AOI21_X1 U18543 ( .B1(n15323), .B2(n16303), .A(n15322), .ZN(n15326) );
  NAND3_X1 U18544 ( .A1(n15324), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n15327), .ZN(n15325) );
  OAI211_X1 U18545 ( .C1(n15328), .C2(n15327), .A(n15326), .B(n15325), .ZN(
        n15329) );
  AOI21_X1 U18546 ( .B1(n15330), .B2(n19204), .A(n15329), .ZN(n15331) );
  OAI21_X1 U18547 ( .B1(n15332), .B2(n19209), .A(n15331), .ZN(P2_U3018) );
  NOR3_X1 U18548 ( .A1(n15334), .A2(n15333), .A3(n16301), .ZN(n15344) );
  NAND2_X1 U18549 ( .A1(n15335), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15340) );
  INV_X1 U18550 ( .A(n15336), .ZN(n15337) );
  AOI21_X1 U18551 ( .B1(n19202), .B2(n15338), .A(n15337), .ZN(n15339) );
  OAI211_X1 U18552 ( .C1(n15341), .C2(n19206), .A(n15340), .B(n15339), .ZN(
        n15342) );
  NOR3_X1 U18553 ( .A1(n15344), .A2(n15343), .A3(n15342), .ZN(n15345) );
  OAI21_X1 U18554 ( .B1(n15346), .B2(n19209), .A(n15345), .ZN(P2_U3019) );
  NAND2_X1 U18555 ( .A1(n15347), .A2(n16309), .ZN(n15357) );
  INV_X1 U18556 ( .A(n15348), .ZN(n15366) );
  XNOR2_X1 U18557 ( .A(n15350), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15355) );
  NOR2_X1 U18558 ( .A1(n15349), .A2(n15374), .ZN(n15373) );
  NOR3_X1 U18559 ( .A1(n16277), .A2(n15373), .A3(n15350), .ZN(n15354) );
  NAND2_X1 U18560 ( .A1(n19202), .A2(n16081), .ZN(n15351) );
  OAI211_X1 U18561 ( .C1(n16074), .C2(n19206), .A(n15352), .B(n15351), .ZN(
        n15353) );
  AOI211_X1 U18562 ( .C1(n15366), .C2(n15355), .A(n15354), .B(n15353), .ZN(
        n15356) );
  OAI211_X1 U18563 ( .C1(n15358), .C2(n16301), .A(n15357), .B(n15356), .ZN(
        P2_U3020) );
  NOR3_X1 U18564 ( .A1(n16277), .A2(n15373), .A3(n15365), .ZN(n15364) );
  NAND2_X1 U18565 ( .A1(n19202), .A2(n15359), .ZN(n15360) );
  OAI211_X1 U18566 ( .C1(n15362), .C2(n19206), .A(n15361), .B(n15360), .ZN(
        n15363) );
  AOI211_X1 U18567 ( .C1(n15366), .C2(n15365), .A(n15364), .B(n15363), .ZN(
        n15369) );
  NAND2_X1 U18568 ( .A1(n15367), .A2(n19204), .ZN(n15368) );
  OAI211_X1 U18569 ( .C1(n15370), .C2(n19209), .A(n15369), .B(n15368), .ZN(
        P2_U3021) );
  NAND2_X1 U18570 ( .A1(n15371), .A2(n16309), .ZN(n15380) );
  INV_X1 U18571 ( .A(n16086), .ZN(n15378) );
  OAI21_X1 U18572 ( .B1(n16306), .B2(n16085), .A(n15372), .ZN(n15377) );
  AOI21_X1 U18573 ( .B1(n15375), .B2(n15374), .A(n15373), .ZN(n15376) );
  AOI211_X1 U18574 ( .C1(n16303), .C2(n15378), .A(n15377), .B(n15376), .ZN(
        n15379) );
  OAI211_X1 U18575 ( .C1(n16301), .C2(n15381), .A(n15380), .B(n15379), .ZN(
        P2_U3022) );
  XNOR2_X1 U18576 ( .A(n15403), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15386) );
  AOI22_X1 U18577 ( .A1(n15382), .A2(n16303), .B1(P2_REIP_REG_23__SCAN_IN), 
        .B2(n19192), .ZN(n15383) );
  OAI21_X1 U18578 ( .B1(n16306), .B2(n15384), .A(n15383), .ZN(n15385) );
  AOI21_X1 U18579 ( .B1(n15404), .B2(n15386), .A(n15385), .ZN(n15387) );
  OAI21_X1 U18580 ( .B1(n15416), .B2(n15388), .A(n15387), .ZN(n15389) );
  AOI21_X1 U18581 ( .B1(n15390), .B2(n19204), .A(n15389), .ZN(n15391) );
  OAI21_X1 U18582 ( .B1(n15392), .B2(n19209), .A(n15391), .ZN(P2_U3023) );
  NAND2_X1 U18583 ( .A1(n15395), .A2(n15394), .ZN(n15396) );
  XNOR2_X1 U18584 ( .A(n15393), .B(n15396), .ZN(n16109) );
  INV_X1 U18585 ( .A(n16109), .ZN(n15409) );
  NAND2_X1 U18586 ( .A1(n15397), .A2(n15403), .ZN(n15399) );
  AND2_X1 U18587 ( .A1(n15399), .A2(n15398), .ZN(n16107) );
  NOR2_X1 U18588 ( .A1(n12856), .A2(n19033), .ZN(n15402) );
  NOR2_X1 U18589 ( .A1(n16306), .A2(n15400), .ZN(n15401) );
  AOI211_X1 U18590 ( .C1(n16108), .C2(n16303), .A(n15402), .B(n15401), .ZN(
        n15406) );
  INV_X1 U18591 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15403) );
  NAND2_X1 U18592 ( .A1(n15404), .A2(n15403), .ZN(n15405) );
  OAI211_X1 U18593 ( .C1(n15416), .C2(n15403), .A(n15406), .B(n15405), .ZN(
        n15407) );
  AOI21_X1 U18594 ( .B1(n16107), .B2(n19204), .A(n15407), .ZN(n15408) );
  OAI21_X1 U18595 ( .B1(n15409), .B2(n19209), .A(n15408), .ZN(P2_U3024) );
  NAND2_X1 U18596 ( .A1(n15410), .A2(n16309), .ZN(n15421) );
  NOR2_X1 U18597 ( .A1(n9984), .A2(n15535), .ZN(n15516) );
  NAND2_X1 U18598 ( .A1(n15423), .A2(n15516), .ZN(n15480) );
  NOR2_X1 U18599 ( .A1(n16234), .A2(n15480), .ZN(n16230) );
  NAND2_X1 U18600 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16230), .ZN(
        n15430) );
  INV_X1 U18601 ( .A(n15430), .ZN(n15441) );
  NAND4_X1 U18602 ( .A1(n15415), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A4(n15441), .ZN(n15412) );
  OAI211_X1 U18603 ( .C1(n15414), .C2(n19206), .A(n15413), .B(n15412), .ZN(
        n15418) );
  NOR2_X1 U18604 ( .A1(n15416), .A2(n15415), .ZN(n15417) );
  AOI211_X1 U18605 ( .C1(n19202), .C2(n15419), .A(n15418), .B(n15417), .ZN(
        n15420) );
  OAI211_X1 U18606 ( .C1(n15422), .C2(n16301), .A(n15421), .B(n15420), .ZN(
        P2_U3025) );
  AOI22_X1 U18607 ( .A1(n9984), .A2(n19201), .B1(n16257), .B2(n16258), .ZN(
        n15502) );
  NAND2_X1 U18608 ( .A1(n16257), .A2(n9980), .ZN(n15424) );
  NAND2_X1 U18609 ( .A1(n15502), .A2(n15424), .ZN(n16235) );
  INV_X1 U18610 ( .A(n16235), .ZN(n15425) );
  OAI21_X1 U18611 ( .B1(n15427), .B2(n15426), .A(n15425), .ZN(n15448) );
  NAND2_X1 U18612 ( .A1(n15448), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15434) );
  XNOR2_X1 U18613 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15429) );
  OAI21_X1 U18614 ( .B1(n15430), .B2(n15429), .A(n15428), .ZN(n15431) );
  AOI21_X1 U18615 ( .B1(n15432), .B2(n16303), .A(n15431), .ZN(n15433) );
  OAI211_X1 U18616 ( .C1(n16306), .C2(n16096), .A(n15434), .B(n15433), .ZN(
        n15435) );
  AOI21_X1 U18617 ( .B1(n15436), .B2(n19204), .A(n15435), .ZN(n15437) );
  OAI21_X1 U18618 ( .B1(n15438), .B2(n19209), .A(n15437), .ZN(P2_U3026) );
  NAND2_X1 U18619 ( .A1(n15439), .A2(n16309), .ZN(n15450) );
  NOR2_X1 U18620 ( .A1(n19206), .A2(n15440), .ZN(n15447) );
  NAND2_X1 U18621 ( .A1(n15442), .A2(n15441), .ZN(n15443) );
  OAI211_X1 U18622 ( .C1(n16306), .C2(n15445), .A(n15444), .B(n15443), .ZN(
        n15446) );
  AOI211_X1 U18623 ( .C1(n15448), .C2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15447), .B(n15446), .ZN(n15449) );
  OAI211_X1 U18624 ( .C1(n15451), .C2(n16301), .A(n15450), .B(n15449), .ZN(
        P2_U3027) );
  XOR2_X1 U18625 ( .A(n15453), .B(n15452), .Z(n16131) );
  AND2_X1 U18626 ( .A1(n19192), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n16128) );
  INV_X1 U18627 ( .A(n16128), .ZN(n15454) );
  OAI21_X1 U18628 ( .B1(n16306), .B2(n18954), .A(n15454), .ZN(n15462) );
  OR2_X1 U18629 ( .A1(n16120), .A2(n15463), .ZN(n16127) );
  NAND2_X1 U18630 ( .A1(n16301), .A2(n15455), .ZN(n15459) );
  NOR2_X1 U18631 ( .A1(n15456), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15457) );
  OR2_X1 U18632 ( .A1(n16235), .A2(n15457), .ZN(n15458) );
  AOI21_X1 U18633 ( .B1(n19201), .B2(n15463), .A(n10893), .ZN(n15461) );
  OAI22_X1 U18634 ( .A1(n15482), .A2(n15480), .B1(n16301), .B2(n16120), .ZN(
        n15469) );
  AOI21_X1 U18635 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15469), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15460) );
  NOR2_X1 U18636 ( .A1(n15464), .A2(n15463), .ZN(n15468) );
  AOI22_X1 U18637 ( .A1(n19202), .A2(n19080), .B1(P2_REIP_REG_16__SCAN_IN), 
        .B2(n19192), .ZN(n15465) );
  OAI21_X1 U18638 ( .B1(n19206), .B2(n15466), .A(n15465), .ZN(n15467) );
  AOI211_X1 U18639 ( .C1(n15469), .C2(n15463), .A(n15468), .B(n15467), .ZN(
        n15470) );
  OAI21_X1 U18640 ( .B1(n19209), .B2(n15471), .A(n15470), .ZN(P2_U3030) );
  NOR2_X1 U18641 ( .A1(n15473), .A2(n15472), .ZN(n15479) );
  INV_X1 U18642 ( .A(n15477), .ZN(n15476) );
  NOR2_X1 U18643 ( .A1(n15476), .A2(n15475), .ZN(n15498) );
  NAND2_X1 U18644 ( .A1(n15499), .A2(n15498), .ZN(n15497) );
  NAND2_X1 U18645 ( .A1(n15497), .A2(n15477), .ZN(n15478) );
  XOR2_X1 U18646 ( .A(n15479), .B(n15478), .Z(n16136) );
  OAI21_X1 U18647 ( .B1(n15492), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n16120), .ZN(n16135) );
  INV_X1 U18648 ( .A(n15480), .ZN(n15483) );
  NOR2_X1 U18649 ( .A1(n12839), .A2(n19033), .ZN(n15481) );
  AOI221_X1 U18650 ( .B1(n15483), .B2(n15482), .C1(n16235), .C2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(n15481), .ZN(n15489) );
  OAI21_X1 U18651 ( .B1(n15486), .B2(n15484), .A(n15485), .ZN(n19087) );
  INV_X1 U18652 ( .A(n19087), .ZN(n15487) );
  AOI22_X1 U18653 ( .A1(n16303), .A2(n18957), .B1(n19202), .B2(n15487), .ZN(
        n15488) );
  OAI211_X1 U18654 ( .C1(n16135), .C2(n16301), .A(n15489), .B(n15488), .ZN(
        n15490) );
  INV_X1 U18655 ( .A(n15490), .ZN(n15491) );
  OAI21_X1 U18656 ( .B1(n16136), .B2(n19209), .A(n15491), .ZN(P2_U3031) );
  INV_X1 U18657 ( .A(n15492), .ZN(n15496) );
  INV_X1 U18658 ( .A(n15501), .ZN(n15493) );
  NAND2_X1 U18659 ( .A1(n16165), .A2(n15493), .ZN(n15526) );
  NAND2_X1 U18660 ( .A1(n15526), .A2(n15494), .ZN(n15495) );
  INV_X1 U18661 ( .A(n16141), .ZN(n15510) );
  OAI21_X1 U18662 ( .B1(n15499), .B2(n15498), .A(n15497), .ZN(n16142) );
  NAND2_X1 U18663 ( .A1(n16142), .A2(n16309), .ZN(n15509) );
  AOI21_X1 U18664 ( .B1(n15500), .B2(n15518), .A(n15484), .ZN(n19088) );
  OAI22_X1 U18665 ( .A1(n19206), .A2(n16140), .B1(n12810), .B2(n19033), .ZN(
        n15507) );
  INV_X1 U18666 ( .A(n15516), .ZN(n16244) );
  NOR2_X1 U18667 ( .A1(n15501), .A2(n16244), .ZN(n15505) );
  OAI21_X1 U18668 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16244), .A(
        n15502), .ZN(n16242) );
  AOI21_X1 U18669 ( .B1(n15516), .B2(n15525), .A(n16242), .ZN(n15503) );
  INV_X1 U18670 ( .A(n15503), .ZN(n15504) );
  MUX2_X1 U18671 ( .A(n15505), .B(n15504), .S(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n15506) );
  AOI211_X1 U18672 ( .C1(n19202), .C2(n19088), .A(n15507), .B(n15506), .ZN(
        n15508) );
  OAI211_X1 U18673 ( .C1(n15510), .C2(n16301), .A(n15509), .B(n15508), .ZN(
        P2_U3032) );
  INV_X1 U18674 ( .A(n15511), .ZN(n15515) );
  OAI21_X1 U18675 ( .B1(n15513), .B2(n15515), .A(n15512), .ZN(n15514) );
  OAI21_X1 U18676 ( .B1(n15474), .B2(n15515), .A(n15514), .ZN(n16146) );
  NAND2_X1 U18677 ( .A1(n15516), .A2(n15525), .ZN(n15523) );
  NOR2_X1 U18678 ( .A1(n12807), .A2(n19033), .ZN(n15517) );
  AOI21_X1 U18679 ( .B1(n16303), .B2(n18988), .A(n15517), .ZN(n15522) );
  OAI21_X1 U18680 ( .B1(n15519), .B2(n16240), .A(n15518), .ZN(n19093) );
  INV_X1 U18681 ( .A(n19093), .ZN(n15520) );
  NAND2_X1 U18682 ( .A1(n19202), .A2(n15520), .ZN(n15521) );
  OAI211_X1 U18683 ( .C1(n15523), .C2(n11046), .A(n15522), .B(n15521), .ZN(
        n15524) );
  AOI21_X1 U18684 ( .B1(n16242), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15524), .ZN(n15529) );
  NAND2_X1 U18685 ( .A1(n16165), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16154) );
  NAND2_X1 U18686 ( .A1(n16154), .A2(n15525), .ZN(n15527) );
  NAND2_X1 U18687 ( .A1(n15527), .A2(n15526), .ZN(n16145) );
  OR2_X1 U18688 ( .A1(n16145), .A2(n16301), .ZN(n15528) );
  OAI211_X1 U18689 ( .C1(n16146), .C2(n19209), .A(n15529), .B(n15528), .ZN(
        P2_U3033) );
  INV_X1 U18690 ( .A(n16172), .ZN(n15531) );
  OR2_X1 U18691 ( .A1(n15531), .A2(n15530), .ZN(n15532) );
  XNOR2_X1 U18692 ( .A(n15533), .B(n15532), .ZN(n16186) );
  AND2_X1 U18693 ( .A1(n15534), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16164) );
  INV_X1 U18694 ( .A(n16164), .ZN(n16179) );
  OAI21_X1 U18695 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15534), .A(
        n16179), .ZN(n16187) );
  AND2_X1 U18696 ( .A1(n16257), .A2(n16258), .ZN(n15537) );
  INV_X1 U18697 ( .A(n15535), .ZN(n16253) );
  NOR2_X1 U18698 ( .A1(n12744), .A2(n19033), .ZN(n15536) );
  AOI221_X1 U18699 ( .B1(n15537), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n16253), .C2(n10843), .A(n15536), .ZN(n15542) );
  OAI21_X1 U18700 ( .B1(n15539), .B2(n14113), .A(n15538), .ZN(n19105) );
  INV_X1 U18701 ( .A(n19105), .ZN(n15540) );
  AOI22_X1 U18702 ( .A1(n16303), .A2(n19024), .B1(n19202), .B2(n15540), .ZN(
        n15541) );
  OAI211_X1 U18703 ( .C1(n16187), .C2(n16301), .A(n15542), .B(n15541), .ZN(
        n15543) );
  INV_X1 U18704 ( .A(n15543), .ZN(n15544) );
  OAI21_X1 U18705 ( .B1(n19209), .B2(n16186), .A(n15544), .ZN(P2_U3037) );
  NAND2_X1 U18706 ( .A1(n16257), .A2(n15545), .ZN(n15547) );
  NAND2_X1 U18707 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n19192), .ZN(n15546) );
  OAI221_X1 U18708 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15549), .C1(
        n15548), .C2(n15547), .A(n15546), .ZN(n15553) );
  INV_X1 U18709 ( .A(n15550), .ZN(n19112) );
  OAI22_X1 U18710 ( .A1(n16306), .A2(n19112), .B1(n19206), .B2(n15551), .ZN(
        n15552) );
  AOI211_X1 U18711 ( .C1(n15554), .C2(n16309), .A(n15553), .B(n15552), .ZN(
        n15555) );
  OAI21_X1 U18712 ( .B1(n15556), .B2(n16301), .A(n15555), .ZN(P2_U3040) );
  XNOR2_X1 U18713 ( .A(n15558), .B(n15557), .ZN(n16210) );
  NAND2_X1 U18714 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15559) );
  OAI211_X1 U18715 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n15560), .B(n15559), .ZN(n15564) );
  XNOR2_X1 U18716 ( .A(n15561), .B(n9777), .ZN(n19118) );
  INV_X1 U18717 ( .A(n19118), .ZN(n15562) );
  AOI22_X1 U18718 ( .A1(n19202), .A2(n15562), .B1(n19192), .B2(
        P2_REIP_REG_5__SCAN_IN), .ZN(n15563) );
  OAI211_X1 U18719 ( .C1(n19206), .C2(n15565), .A(n15564), .B(n15563), .ZN(
        n15572) );
  OAI21_X1 U18720 ( .B1(n15569), .B2(n15567), .A(n15566), .ZN(n15568) );
  OAI21_X1 U18721 ( .B1(n15570), .B2(n15569), .A(n15568), .ZN(n16208) );
  NOR2_X1 U18722 ( .A1(n16208), .A2(n16301), .ZN(n15571) );
  AOI211_X1 U18723 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n15573), .A(
        n15572), .B(n15571), .ZN(n15574) );
  OAI21_X1 U18724 ( .B1(n19209), .B2(n16210), .A(n15574), .ZN(P2_U3041) );
  INV_X1 U18725 ( .A(n16362), .ZN(n15606) );
  MUX2_X1 U18726 ( .A(n15575), .B(n13609), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15576) );
  AOI21_X1 U18727 ( .B1(n19063), .B2(n15605), .A(n15576), .ZN(n16318) );
  INV_X1 U18728 ( .A(n15577), .ZN(n15578) );
  OAI222_X1 U18729 ( .A1(n15606), .A2(n15579), .B1(n19816), .B2(n16318), .C1(
        n14188), .C2(n15578), .ZN(n15580) );
  MUX2_X1 U18730 ( .A(n15580), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n15607), .Z(P2_U3601) );
  INV_X1 U18731 ( .A(n15581), .ZN(n15592) );
  NOR2_X1 U18732 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15590) );
  INV_X1 U18733 ( .A(n15582), .ZN(n15583) );
  NAND2_X1 U18734 ( .A1(n13609), .A2(n15583), .ZN(n15595) );
  OAI21_X1 U18735 ( .B1(n15585), .B2(n15584), .A(n13048), .ZN(n15597) );
  NOR2_X1 U18736 ( .A1(n14181), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15600) );
  NOR2_X1 U18737 ( .A1(n16336), .A2(n15586), .ZN(n15601) );
  OAI21_X1 U18738 ( .B1(n15597), .B2(n15600), .A(n15601), .ZN(n15588) );
  INV_X1 U18739 ( .A(n15600), .ZN(n15596) );
  NAND3_X1 U18740 ( .A1(n15597), .A2(n13048), .A3(n15596), .ZN(n15587) );
  NAND2_X1 U18741 ( .A1(n15588), .A2(n15587), .ZN(n15589) );
  OAI21_X1 U18742 ( .B1(n15590), .B2(n15595), .A(n15589), .ZN(n15591) );
  AOI21_X1 U18743 ( .B1(n10688), .B2(n15605), .A(n15591), .ZN(n16315) );
  OAI222_X1 U18744 ( .A1(n15606), .A2(n19913), .B1(n15593), .B2(n15592), .C1(
        n19816), .C2(n16315), .ZN(n15594) );
  MUX2_X1 U18745 ( .A(n15594), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15607), .Z(P2_U3599) );
  NAND3_X1 U18746 ( .A1(n15597), .A2(n15596), .A3(n15595), .ZN(n15603) );
  AOI21_X1 U18747 ( .B1(n13609), .B2(n15582), .A(n15598), .ZN(n15599) );
  OAI21_X1 U18748 ( .B1(n15601), .B2(n15600), .A(n15599), .ZN(n15602) );
  MUX2_X1 U18749 ( .A(n15603), .B(n15602), .S(n10510), .Z(n15604) );
  OAI22_X1 U18750 ( .A1(n19904), .A2(n15606), .B1(n16323), .B2(n19816), .ZN(
        n15608) );
  MUX2_X1 U18751 ( .A(n15608), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15607), .Z(P2_U3596) );
  INV_X1 U18752 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n16916) );
  INV_X1 U18753 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16914) );
  INV_X1 U18754 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16670) );
  NAND2_X1 U18755 ( .A1(n18727), .A2(n15609), .ZN(n15709) );
  INV_X1 U18756 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17094) );
  INV_X1 U18757 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16748) );
  INV_X1 U18758 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n15613) );
  NAND3_X1 U18759 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17239) );
  NOR3_X1 U18760 ( .A1(n15613), .A2(n16866), .A3(n17239), .ZN(n17130) );
  INV_X1 U18761 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17231) );
  INV_X1 U18762 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17235) );
  NAND4_X1 U18763 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(P3_EBX_REG_9__SCAN_IN), .A4(P3_EBX_REG_8__SCAN_IN), .ZN(n15614) );
  NOR3_X1 U18764 ( .A1(n17231), .A2(n17235), .A3(n15614), .ZN(n17131) );
  NAND4_X1 U18765 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(n17130), .A4(n17131), .ZN(n15700) );
  NOR2_X1 U18766 ( .A1(n16748), .A2(n15700), .ZN(n17108) );
  NAND3_X1 U18767 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(n17108), .ZN(n17091) );
  NOR2_X1 U18768 ( .A1(n17094), .A2(n17091), .ZN(n17076) );
  NAND2_X1 U18769 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17076), .ZN(n17075) );
  NOR2_X1 U18770 ( .A1(n17079), .A2(n17075), .ZN(n17061) );
  NAND2_X1 U18771 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17061), .ZN(n17043) );
  NAND2_X1 U18772 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17044), .ZN(n17027) );
  NOR2_X1 U18773 ( .A1(n17345), .A2(n17027), .ZN(n16997) );
  NAND2_X1 U18774 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16997), .ZN(n16982) );
  NAND2_X1 U18775 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n16996), .ZN(n16971) );
  NAND2_X1 U18776 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16970), .ZN(n16961) );
  INV_X1 U18777 ( .A(n16961), .ZN(n16966) );
  NAND2_X1 U18778 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16966), .ZN(n15688) );
  INV_X1 U18779 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n16918) );
  INV_X1 U18780 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16917) );
  NOR3_X1 U18781 ( .A1(n16918), .A2(n16917), .A3(n16961), .ZN(n16955) );
  NOR2_X1 U18782 ( .A1(n17257), .A2(n16955), .ZN(n16956) );
  AOI22_X1 U18783 ( .A1(n11217), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15615) );
  OAI21_X1 U18784 ( .B1(n17223), .B2(n17000), .A(n15615), .ZN(n15624) );
  AOI22_X1 U18785 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9663), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15622) );
  OAI22_X1 U18786 ( .A1(n17188), .A2(n15691), .B1(n17133), .B2(n16998), .ZN(
        n15620) );
  AOI22_X1 U18787 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15618) );
  AOI22_X1 U18788 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15617) );
  AOI22_X1 U18789 ( .A1(n11202), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15616) );
  NAND3_X1 U18790 ( .A1(n15618), .A2(n15617), .A3(n15616), .ZN(n15619) );
  AOI211_X1 U18791 ( .C1(n17214), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n15620), .B(n15619), .ZN(n15621) );
  OAI211_X1 U18792 ( .C1(n11187), .C2(n16999), .A(n15622), .B(n15621), .ZN(
        n15623) );
  AOI211_X1 U18793 ( .C1(n17184), .C2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n15624), .B(n15623), .ZN(n15686) );
  AOI22_X1 U18794 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15625) );
  OAI21_X1 U18795 ( .B1(n17223), .B2(n17032), .A(n15625), .ZN(n15634) );
  AOI22_X1 U18796 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15632) );
  INV_X1 U18797 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17147) );
  INV_X1 U18798 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17154) );
  OAI22_X1 U18799 ( .A1(n11187), .A2(n17147), .B1(n11186), .B2(n17154), .ZN(
        n15630) );
  AOI22_X1 U18800 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15628) );
  AOI22_X1 U18801 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15627) );
  AOI22_X1 U18802 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15626) );
  NAND3_X1 U18803 ( .A1(n15628), .A2(n15627), .A3(n15626), .ZN(n15629) );
  AOI211_X1 U18804 ( .C1(n11202), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n15630), .B(n15629), .ZN(n15631) );
  OAI211_X1 U18805 ( .C1(n17133), .C2(n17148), .A(n15632), .B(n15631), .ZN(
        n15633) );
  AOI211_X1 U18806 ( .C1(n11207), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n15634), .B(n15633), .ZN(n16963) );
  AOI22_X1 U18807 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9649), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17189), .ZN(n15635) );
  OAI21_X1 U18808 ( .B1(n17252), .B2(n9713), .A(n15635), .ZN(n15644) );
  INV_X1 U18809 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17200) );
  AOI22_X1 U18810 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15642) );
  AOI22_X1 U18811 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n9663), .B1(
        n11202), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15636) );
  OAI21_X1 U18812 ( .B1(n11187), .B2(n17187), .A(n15636), .ZN(n15640) );
  AOI22_X1 U18813 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17184), .ZN(n15638) );
  AOI22_X1 U18814 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11217), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17149), .ZN(n15637) );
  OAI211_X1 U18815 ( .C1(n18557), .C2(n17053), .A(n15638), .B(n15637), .ZN(
        n15639) );
  AOI211_X1 U18816 ( .C1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .C2(n17049), .A(
        n15640), .B(n15639), .ZN(n15641) );
  OAI211_X1 U18817 ( .C1(n17223), .C2(n17200), .A(n15642), .B(n15641), .ZN(
        n15643) );
  AOI211_X1 U18818 ( .C1(n17212), .C2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n15644), .B(n15643), .ZN(n16973) );
  AOI22_X1 U18819 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15654) );
  INV_X1 U18820 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18554) );
  AOI22_X1 U18821 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11148), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15646) );
  AOI22_X1 U18822 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17167), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15645) );
  OAI211_X1 U18823 ( .C1(n11287), .C2(n18554), .A(n15646), .B(n15645), .ZN(
        n15652) );
  AOI22_X1 U18824 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15650) );
  AOI22_X1 U18825 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15649) );
  AOI22_X1 U18826 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9663), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15648) );
  NAND2_X1 U18827 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n15647) );
  NAND4_X1 U18828 ( .A1(n15650), .A2(n15649), .A3(n15648), .A4(n15647), .ZN(
        n15651) );
  AOI211_X1 U18829 ( .C1(n11202), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n15652), .B(n15651), .ZN(n15653) );
  OAI211_X1 U18830 ( .C1(n16983), .C2(n15655), .A(n15654), .B(n15653), .ZN(
        n16978) );
  AOI22_X1 U18831 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15665) );
  AOI22_X1 U18832 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15657) );
  AOI22_X1 U18833 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15656) );
  OAI211_X1 U18834 ( .C1(n11287), .C2(n17096), .A(n15657), .B(n15656), .ZN(
        n15663) );
  AOI22_X1 U18835 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11148), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15661) );
  AOI22_X1 U18836 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15660) );
  AOI22_X1 U18837 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9663), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15659) );
  NAND2_X1 U18838 ( .A1(n11202), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n15658) );
  NAND4_X1 U18839 ( .A1(n15661), .A2(n15660), .A3(n15659), .A4(n15658), .ZN(
        n15662) );
  AOI211_X1 U18840 ( .C1(n17049), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n15663), .B(n15662), .ZN(n15664) );
  OAI211_X1 U18841 ( .C1(n9746), .C2(n16935), .A(n15665), .B(n15664), .ZN(
        n16979) );
  NAND2_X1 U18842 ( .A1(n16978), .A2(n16979), .ZN(n16977) );
  NOR2_X1 U18843 ( .A1(n16973), .A2(n16977), .ZN(n16972) );
  AOI22_X1 U18844 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15675) );
  AOI22_X1 U18845 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15666) );
  OAI21_X1 U18846 ( .B1(n17015), .B2(n17250), .A(n15666), .ZN(n15673) );
  OAI22_X1 U18847 ( .A1(n11187), .A2(n17058), .B1(n17053), .B2(n18560), .ZN(
        n15667) );
  AOI21_X1 U18848 ( .B1(n11202), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n15667), .ZN(n15671) );
  AOI22_X1 U18849 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17212), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15670) );
  AOI22_X1 U18850 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15669) );
  AOI22_X1 U18851 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9663), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15668) );
  NAND4_X1 U18852 ( .A1(n15671), .A2(n15670), .A3(n15669), .A4(n15668), .ZN(
        n15672) );
  AOI211_X1 U18853 ( .C1(n17167), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n15673), .B(n15672), .ZN(n15674) );
  OAI211_X1 U18854 ( .C1(n17116), .C2(n17170), .A(n15675), .B(n15674), .ZN(
        n16968) );
  NAND2_X1 U18855 ( .A1(n16972), .A2(n16968), .ZN(n16967) );
  NOR2_X1 U18856 ( .A1(n16963), .A2(n16967), .ZN(n16962) );
  AOI22_X1 U18857 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15685) );
  AOI22_X1 U18858 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15684) );
  OAI22_X1 U18859 ( .A1(n11187), .A2(n17016), .B1(n11287), .B2(n18565), .ZN(
        n15682) );
  AOI22_X1 U18860 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15680) );
  AOI22_X1 U18861 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11148), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15677) );
  AOI22_X1 U18862 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15676) );
  OAI211_X1 U18863 ( .C1(n17155), .C2(n17134), .A(n15677), .B(n15676), .ZN(
        n15678) );
  AOI21_X1 U18864 ( .B1(n9663), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(n15678), .ZN(n15679) );
  OAI211_X1 U18865 ( .C1(n16983), .C2(n17026), .A(n15680), .B(n15679), .ZN(
        n15681) );
  AOI211_X1 U18866 ( .C1(n11202), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n15682), .B(n15681), .ZN(n15683) );
  NAND3_X1 U18867 ( .A1(n15685), .A2(n15684), .A3(n15683), .ZN(n16959) );
  NAND2_X1 U18868 ( .A1(n16962), .A2(n16959), .ZN(n16958) );
  NOR2_X1 U18869 ( .A1(n15686), .A2(n16958), .ZN(n16953) );
  AOI21_X1 U18870 ( .B1(n15686), .B2(n16958), .A(n16953), .ZN(n17276) );
  AOI22_X1 U18871 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16956), .B1(n17276), 
        .B2(n17257), .ZN(n15687) );
  OAI21_X1 U18872 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n15688), .A(n15687), .ZN(
        P3_U2675) );
  AOI22_X1 U18873 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11148), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15699) );
  AOI22_X1 U18874 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17210), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15690) );
  AOI22_X1 U18875 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15689) );
  OAI211_X1 U18876 ( .C1(n17053), .C2(n15691), .A(n15690), .B(n15689), .ZN(
        n15697) );
  AOI22_X1 U18877 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15695) );
  AOI22_X1 U18878 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15694) );
  AOI22_X1 U18879 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15693) );
  NAND2_X1 U18880 ( .A1(n9663), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n15692) );
  NAND4_X1 U18881 ( .A1(n15695), .A2(n15694), .A3(n15693), .A4(n15692), .ZN(
        n15696) );
  AOI211_X1 U18882 ( .C1(n11202), .C2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n15697), .B(n15696), .ZN(n15698) );
  OAI211_X1 U18883 ( .C1(n17116), .C2(n16998), .A(n15699), .B(n15698), .ZN(
        n17356) );
  NAND2_X1 U18884 ( .A1(n18266), .A2(n17260), .ZN(n17255) );
  AOI211_X1 U18885 ( .C1(n16748), .C2(n15700), .A(n17108), .B(n17255), .ZN(
        n15701) );
  AOI21_X1 U18886 ( .B1(n17257), .B2(n17356), .A(n15701), .ZN(n15702) );
  OAI21_X1 U18887 ( .B1(n17260), .B2(n16748), .A(n15702), .ZN(P3_U2690) );
  NAND2_X1 U18888 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18401) );
  AOI221_X1 U18889 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18401), .C1(n15704), 
        .C2(n18401), .A(n15703), .ZN(n18228) );
  NOR2_X1 U18890 ( .A1(n15705), .A2(n18709), .ZN(n15706) );
  OAI21_X1 U18891 ( .B1(n15706), .B2(n18585), .A(n18229), .ZN(n18226) );
  AOI22_X1 U18892 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18228), .B1(
        n18226), .B2(n18714), .ZN(P3_U2865) );
  NAND4_X1 U18893 ( .A1(n17416), .A2(n17415), .A3(n18907), .A4(n18725), .ZN(
        n15708) );
  NAND4_X1 U18894 ( .A1(n15710), .A2(n15709), .A3(n15799), .A4(n15708), .ZN(
        n18734) );
  NOR2_X1 U18895 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18854), .ZN(n18233) );
  INV_X1 U18896 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18224) );
  NOR2_X1 U18897 ( .A1(n18224), .A2(n18852), .ZN(n15711) );
  INV_X1 U18898 ( .A(n18888), .ZN(n18885) );
  INV_X1 U18899 ( .A(n16525), .ZN(n18692) );
  NOR2_X1 U18900 ( .A1(n15712), .A2(n18692), .ZN(n18730) );
  NAND3_X1 U18901 ( .A1(n18885), .A2(n18883), .A3(n18730), .ZN(n15713) );
  OAI21_X1 U18902 ( .B1(n18885), .B2(n18735), .A(n15713), .ZN(P3_U3284) );
  NAND2_X1 U18903 ( .A1(n15715), .A2(n15714), .ZN(n15716) );
  XNOR2_X1 U18904 ( .A(n15716), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16405) );
  OAI21_X1 U18905 ( .B1(n18092), .B2(n16388), .A(n15717), .ZN(n15718) );
  AOI21_X1 U18906 ( .B1(n18722), .B2(n16402), .A(n15718), .ZN(n15719) );
  NOR2_X1 U18907 ( .A1(n15719), .A2(n18218), .ZN(n15774) );
  NOR2_X1 U18908 ( .A1(n18729), .A2(n18218), .ZN(n18216) );
  NAND2_X1 U18909 ( .A1(n15720), .A2(n18216), .ZN(n18137) );
  NAND2_X1 U18910 ( .A1(n18722), .A2(n18196), .ZN(n18175) );
  OAI22_X1 U18911 ( .A1(n16387), .A2(n18137), .B1(n16400), .B2(n18175), .ZN(
        n15775) );
  AOI22_X1 U18912 ( .A1(n18126), .A2(n17534), .B1(n18217), .B2(n15721), .ZN(
        n15722) );
  NAND2_X1 U18913 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15722), .ZN(
        n15723) );
  OAI22_X1 U18914 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15774), .B1(
        n15775), .B2(n15723), .ZN(n15724) );
  NAND2_X1 U18915 ( .A1(n9647), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16394) );
  OAI211_X1 U18916 ( .C1(n16405), .C2(n18109), .A(n15724), .B(n16394), .ZN(
        P3_U2833) );
  INV_X1 U18917 ( .A(n15725), .ZN(n15732) );
  NAND2_X1 U18918 ( .A1(n15725), .A2(n15726), .ZN(n15737) );
  AOI21_X1 U18919 ( .B1(n15727), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n20634), .ZN(n15728) );
  AND2_X1 U18920 ( .A1(n15729), .A2(n15728), .ZN(n15731) );
  INV_X1 U18921 ( .A(n15731), .ZN(n15735) );
  INV_X1 U18922 ( .A(n15730), .ZN(n15733) );
  OAI22_X1 U18923 ( .A1(n15733), .A2(n15732), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n15731), .ZN(n15734) );
  OAI21_X1 U18924 ( .B1(n15735), .B2(n20582), .A(n15734), .ZN(n15736) );
  AOI222_X1 U18925 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n15737), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15736), .C1(n15737), 
        .C2(n15736), .ZN(n15738) );
  AOI222_X1 U18926 ( .A1(n20546), .A2(n15739), .B1(n20546), .B2(n15738), .C1(
        n15739), .C2(n15738), .ZN(n15740) );
  OR2_X1 U18927 ( .A1(n15740), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n15750) );
  NAND2_X1 U18928 ( .A1(n20919), .A2(n19983), .ZN(n15743) );
  INV_X1 U18929 ( .A(n15741), .ZN(n15742) );
  AOI21_X1 U18930 ( .B1(n15744), .B2(n15743), .A(n15742), .ZN(n15746) );
  AND4_X1 U18931 ( .A1(n15748), .A2(n15747), .A3(n15746), .A4(n15745), .ZN(
        n15749) );
  INV_X1 U18932 ( .A(n15763), .ZN(n15756) );
  NAND4_X1 U18933 ( .A1(n15752), .A2(n20220), .A3(n15751), .A4(n20874), .ZN(
        n15755) );
  OAI21_X1 U18934 ( .B1(n15753), .B2(n20871), .A(n20775), .ZN(n15754) );
  NAND2_X1 U18935 ( .A1(n15755), .A2(n15754), .ZN(n16051) );
  AOI221_X1 U18936 ( .B1(n16055), .B2(n16053), .C1(n15756), .C2(n16053), .A(
        n16051), .ZN(n15758) );
  NOR2_X1 U18937 ( .A1(n15758), .A2(n16055), .ZN(n20776) );
  OAI211_X1 U18938 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20871), .A(n20776), 
        .B(n15757), .ZN(n16052) );
  AOI21_X1 U18939 ( .B1(n20879), .B2(n20856), .A(n15758), .ZN(n15759) );
  OAI22_X1 U18940 ( .A1(n15760), .A2(n16052), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n15759), .ZN(n15761) );
  OAI21_X1 U18941 ( .B1(n15763), .B2(n15762), .A(n15761), .ZN(P1_U3161) );
  AOI22_X1 U18942 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15764), .B1(
        n20190), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15770) );
  INV_X1 U18943 ( .A(n15765), .ZN(n15768) );
  INV_X1 U18944 ( .A(n15766), .ZN(n15767) );
  AOI22_X1 U18945 ( .A1(n15768), .A2(n20188), .B1(n20203), .B2(n15767), .ZN(
        n15769) );
  OAI211_X1 U18946 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15771), .A(
        n15770), .B(n15769), .ZN(P1_U3010) );
  AOI21_X1 U18947 ( .B1(n15773), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n15772), .ZN(n16386) );
  NOR2_X1 U18948 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16389), .ZN(
        n16382) );
  AOI22_X1 U18949 ( .A1(n9647), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n16382), 
        .B2(n15774), .ZN(n15778) );
  OAI21_X1 U18950 ( .B1(n15776), .B2(n15775), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15777) );
  OAI211_X1 U18951 ( .C1(n16386), .C2(n18109), .A(n15778), .B(n15777), .ZN(
        P3_U2832) );
  INV_X1 U18952 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20778) );
  INV_X1 U18953 ( .A(HOLD), .ZN(n21032) );
  INV_X1 U18954 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20967) );
  OAI22_X1 U18955 ( .A1(n20778), .A2(n21032), .B1(n12453), .B2(n20967), .ZN(
        n15779) );
  OAI21_X1 U18956 ( .B1(n21032), .B2(n11603), .A(n15779), .ZN(n15780) );
  OAI211_X1 U18957 ( .C1(n20871), .C2(n20778), .A(n20875), .B(n15780), .ZN(
        P1_U3195) );
  AND2_X1 U18958 ( .A1(n15781), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR2_X1 U18959 ( .A1(n14651), .A2(n15936), .ZN(n15782) );
  MUX2_X1 U18960 ( .A(n9740), .B(n15782), .S(n15883), .Z(n15783) );
  XNOR2_X1 U18961 ( .A(n15783), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15862) );
  INV_X1 U18962 ( .A(n15980), .ZN(n15999) );
  AOI22_X1 U18963 ( .A1(n15936), .A2(n15785), .B1(n15784), .B2(n20185), .ZN(
        n15786) );
  INV_X1 U18964 ( .A(n15786), .ZN(n15787) );
  AOI211_X1 U18965 ( .C1(n15788), .C2(n15976), .A(n15999), .B(n15787), .ZN(
        n15935) );
  OAI21_X1 U18966 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15789), .A(
        n15935), .ZN(n15790) );
  INV_X1 U18967 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20824) );
  NOR2_X1 U18968 ( .A1(n20170), .A2(n20824), .ZN(n15860) );
  AOI221_X1 U18969 ( .B1(n15792), .B2(n15791), .C1(n15790), .C2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(n15860), .ZN(n15795) );
  INV_X1 U18970 ( .A(n15805), .ZN(n15793) );
  NAND2_X1 U18971 ( .A1(n15793), .A2(n20203), .ZN(n15794) );
  OAI211_X1 U18972 ( .C1(n15862), .C2(n20208), .A(n15795), .B(n15794), .ZN(
        P1_U3011) );
  NOR3_X1 U18973 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n9877), .A3(n19967), 
        .ZN(n16358) );
  NOR4_X1 U18974 ( .A1(n15796), .A2(n19961), .A3(n16371), .A4(n16358), .ZN(
        P2_U3178) );
  INV_X1 U18975 ( .A(n19948), .ZN(n16370) );
  AOI221_X1 U18976 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16371), .C1(n16370), .C2(
        n16371), .A(n19761), .ZN(n19940) );
  INV_X1 U18977 ( .A(n19940), .ZN(n19937) );
  NOR2_X1 U18978 ( .A1(n16329), .A2(n19937), .ZN(P2_U3047) );
  NAND3_X1 U18979 ( .A1(n18906), .A2(n18234), .A3(n15797), .ZN(n15798) );
  NAND2_X1 U18980 ( .A1(n18266), .A2(n17262), .ZN(n17400) );
  INV_X1 U18981 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17476) );
  INV_X1 U18982 ( .A(n17262), .ZN(n17406) );
  AOI22_X1 U18983 ( .A1(n17411), .A2(BUF2_REG_0__SCAN_IN), .B1(n17410), .B2(
        n15800), .ZN(n15801) );
  OAI221_X1 U18984 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17400), .C1(n17476), 
        .C2(n17262), .A(n15801), .ZN(P3_U2735) );
  INV_X1 U18985 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15802) );
  OAI22_X1 U18986 ( .A1(n15802), .A2(n20000), .B1(n20053), .B2(n15857), .ZN(
        n15803) );
  AOI21_X1 U18987 ( .B1(P1_EBX_REG_20__SCAN_IN), .B2(n15848), .A(n15803), .ZN(
        n15804) );
  OAI21_X1 U18988 ( .B1(n15805), .B2(n20014), .A(n15804), .ZN(n15806) );
  AOI21_X1 U18989 ( .B1(n15807), .B2(n20041), .A(n15806), .ZN(n15808) );
  OAI221_X1 U18990 ( .B1(n15810), .B2(n20824), .C1(n15810), .C2(n15809), .A(
        n15808), .ZN(P1_U2820) );
  AOI22_X1 U18991 ( .A1(n15811), .A2(P1_REIP_REG_18__SCAN_IN), .B1(n15848), 
        .B2(P1_EBX_REG_18__SCAN_IN), .ZN(n15812) );
  OAI21_X1 U18992 ( .B1(n15813), .B2(n20053), .A(n15812), .ZN(n15814) );
  AOI211_X1 U18993 ( .C1(n20048), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20040), .B(n15814), .ZN(n15818) );
  INV_X1 U18994 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20821) );
  AOI22_X1 U18995 ( .A1(n15816), .A2(n20041), .B1(n20821), .B2(n15815), .ZN(
        n15817) );
  OAI211_X1 U18996 ( .C1(n20014), .C2(n15944), .A(n15818), .B(n15817), .ZN(
        P1_U2822) );
  AOI22_X1 U18997 ( .A1(n15819), .A2(n20027), .B1(n20047), .B2(n15962), .ZN(
        n15827) );
  INV_X1 U18998 ( .A(n15820), .ZN(n15825) );
  OAI21_X1 U18999 ( .B1(n20000), .B2(n15821), .A(n20049), .ZN(n15822) );
  AOI21_X1 U19000 ( .B1(n15848), .B2(P1_EBX_REG_15__SCAN_IN), .A(n15822), .ZN(
        n15823) );
  OAI21_X1 U19001 ( .B1(n15835), .B2(n20814), .A(n15823), .ZN(n15824) );
  AOI21_X1 U19002 ( .B1(n15825), .B2(n20041), .A(n15824), .ZN(n15826) );
  OAI211_X1 U19003 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n15828), .A(n15827), 
        .B(n15826), .ZN(P1_U2825) );
  NOR2_X1 U19004 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n9722), .ZN(n15836) );
  AOI22_X1 U19005 ( .A1(n15848), .A2(P1_EBX_REG_14__SCAN_IN), .B1(n20027), 
        .B2(n15868), .ZN(n15834) );
  NOR2_X1 U19006 ( .A1(n15829), .A2(n20014), .ZN(n15832) );
  OAI21_X1 U19007 ( .B1(n20000), .B2(n15830), .A(n20049), .ZN(n15831) );
  AOI211_X1 U19008 ( .C1(n15869), .C2(n20041), .A(n15832), .B(n15831), .ZN(
        n15833) );
  OAI211_X1 U19009 ( .C1(n15836), .C2(n15835), .A(n15834), .B(n15833), .ZN(
        P1_U2826) );
  AOI21_X1 U19010 ( .B1(n15837), .B2(P1_REIP_REG_11__SCAN_IN), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15846) );
  INV_X1 U19011 ( .A(n15838), .ZN(n15839) );
  XNOR2_X1 U19012 ( .A(n15840), .B(n15839), .ZN(n15985) );
  AOI22_X1 U19013 ( .A1(n15879), .A2(n20027), .B1(n20047), .B2(n15985), .ZN(
        n15845) );
  INV_X1 U19014 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15856) );
  NOR2_X1 U19015 ( .A1(n20054), .A2(n15856), .ZN(n15843) );
  OAI21_X1 U19016 ( .B1(n20000), .B2(n15841), .A(n20049), .ZN(n15842) );
  AOI211_X1 U19017 ( .C1(n15880), .C2(n20041), .A(n15843), .B(n15842), .ZN(
        n15844) );
  OAI211_X1 U19018 ( .C1(n15847), .C2(n15846), .A(n15845), .B(n15844), .ZN(
        P1_U2828) );
  AOI22_X1 U19019 ( .A1(n15991), .A2(n20047), .B1(n15848), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n15849) );
  OAI21_X1 U19020 ( .B1(n15890), .B2(n20053), .A(n15849), .ZN(n15850) );
  AOI211_X1 U19021 ( .C1(n20048), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20040), .B(n15850), .ZN(n15853) );
  AOI22_X1 U19022 ( .A1(n15887), .A2(n20041), .B1(P1_REIP_REG_11__SCAN_IN), 
        .B2(n15851), .ZN(n15852) );
  OAI211_X1 U19023 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n15854), .A(n15853), 
        .B(n15852), .ZN(P1_U2829) );
  AOI22_X1 U19024 ( .A1(n15880), .A2(n20071), .B1(n20070), .B2(n15985), .ZN(
        n15855) );
  OAI21_X1 U19025 ( .B1(n20075), .B2(n15856), .A(n15855), .ZN(P1_U2860) );
  OAI22_X1 U19026 ( .A1(n15858), .A2(n12495), .B1(n15857), .B2(n20161), .ZN(
        n15859) );
  AOI211_X1 U19027 ( .C1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n20152), .A(
        n15860), .B(n15859), .ZN(n15861) );
  OAI21_X1 U19028 ( .B1(n15862), .B2(n20172), .A(n15861), .ZN(P1_U2979) );
  AOI22_X1 U19029 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20190), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15866) );
  AOI22_X1 U19030 ( .A1(n15864), .A2(n20167), .B1(n20156), .B2(n15863), .ZN(
        n15865) );
  OAI211_X1 U19031 ( .C1(n20161), .C2(n15867), .A(n15866), .B(n15865), .ZN(
        P1_U2983) );
  AOI22_X1 U19032 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20190), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15871) );
  AOI22_X1 U19033 ( .A1(n15869), .A2(n20167), .B1(n15878), .B2(n15868), .ZN(
        n15870) );
  OAI211_X1 U19034 ( .C1(n15872), .C2(n20172), .A(n15871), .B(n15870), .ZN(
        P1_U2985) );
  AOI21_X1 U19035 ( .B1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n10313), .A(
        n15873), .ZN(n15877) );
  OAI21_X1 U19036 ( .B1(n15875), .B2(n15883), .A(n15874), .ZN(n15876) );
  XNOR2_X1 U19037 ( .A(n15877), .B(n15876), .ZN(n15990) );
  AOI22_X1 U19038 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20190), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15882) );
  AOI22_X1 U19039 ( .A1(n15880), .A2(n20167), .B1(n15879), .B2(n15878), .ZN(
        n15881) );
  OAI211_X1 U19040 ( .C1(n15990), .C2(n20172), .A(n15882), .B(n15881), .ZN(
        P1_U2987) );
  AOI22_X1 U19041 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20190), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15889) );
  NOR2_X1 U19042 ( .A1(n14697), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15885) );
  NOR2_X1 U19043 ( .A1(n14667), .A2(n12391), .ZN(n15884) );
  MUX2_X1 U19044 ( .A(n15885), .B(n15884), .S(n15883), .Z(n15886) );
  XNOR2_X1 U19045 ( .A(n15886), .B(n15981), .ZN(n15992) );
  AOI22_X1 U19046 ( .A1(n15992), .A2(n20156), .B1(n20154), .B2(n15887), .ZN(
        n15888) );
  OAI211_X1 U19047 ( .C1(n20161), .C2(n15890), .A(n15889), .B(n15888), .ZN(
        P1_U2988) );
  AOI22_X1 U19048 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20190), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15895) );
  XNOR2_X1 U19049 ( .A(n15891), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15892) );
  XNOR2_X1 U19050 ( .A(n15893), .B(n15892), .ZN(n16028) );
  AOI22_X1 U19051 ( .A1(n16028), .A2(n20156), .B1(n20154), .B2(n20066), .ZN(
        n15894) );
  OAI211_X1 U19052 ( .C1(n20161), .C2(n20025), .A(n15895), .B(n15894), .ZN(
        P1_U2992) );
  AOI22_X1 U19053 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20190), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15901) );
  OAI21_X1 U19054 ( .B1(n15898), .B2(n15897), .A(n15896), .ZN(n15899) );
  INV_X1 U19055 ( .A(n15899), .ZN(n16035) );
  AOI22_X1 U19056 ( .A1(n16035), .A2(n20156), .B1(n20154), .B2(n20042), .ZN(
        n15900) );
  OAI211_X1 U19057 ( .C1(n20161), .C2(n20032), .A(n15901), .B(n15900), .ZN(
        P1_U2993) );
  AOI22_X1 U19058 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20190), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15907) );
  OAI21_X1 U19059 ( .B1(n15904), .B2(n15903), .A(n15902), .ZN(n15905) );
  INV_X1 U19060 ( .A(n15905), .ZN(n16044) );
  AOI22_X1 U19061 ( .A1(n16044), .A2(n20156), .B1(n20154), .B2(n20072), .ZN(
        n15906) );
  OAI211_X1 U19062 ( .C1(n20161), .C2(n20052), .A(n15907), .B(n15906), .ZN(
        P1_U2994) );
  AOI21_X1 U19063 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n20190), .A(n15908), 
        .ZN(n15915) );
  INV_X1 U19064 ( .A(n15909), .ZN(n15911) );
  OAI22_X1 U19065 ( .A1(n15912), .A2(n16014), .B1(n15911), .B2(n15910), .ZN(
        n15913) );
  INV_X1 U19066 ( .A(n15913), .ZN(n15914) );
  OAI211_X1 U19067 ( .C1(n20208), .C2(n15916), .A(n15915), .B(n15914), .ZN(
        P1_U3006) );
  AOI22_X1 U19068 ( .A1(n15918), .A2(n20188), .B1(n20203), .B2(n15917), .ZN(
        n15926) );
  NAND2_X1 U19069 ( .A1(n20190), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15925) );
  NAND3_X1 U19070 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n15919), .A3(
        n14609), .ZN(n15924) );
  NOR3_X1 U19071 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n15921), .A3(
        n15920), .ZN(n15927) );
  OAI221_X1 U19072 ( .B1(n15922), .B2(n20192), .C1(n15922), .C2(n15927), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15923) );
  NAND4_X1 U19073 ( .A1(n15926), .A2(n15925), .A3(n15924), .A4(n15923), .ZN(
        P1_U3007) );
  INV_X1 U19074 ( .A(n15942), .ZN(n15928) );
  AOI22_X1 U19075 ( .A1(n20190), .A2(P1_REIP_REG_23__SCAN_IN), .B1(n15928), 
        .B2(n15927), .ZN(n15933) );
  INV_X1 U19076 ( .A(n15929), .ZN(n15931) );
  AOI22_X1 U19077 ( .A1(n15931), .A2(n20188), .B1(n20203), .B2(n15930), .ZN(
        n15932) );
  OAI211_X1 U19078 ( .C1(n15934), .C2(n14629), .A(n15933), .B(n15932), .ZN(
        P1_U3008) );
  OAI22_X1 U19079 ( .A1(n15936), .A2(n15935), .B1(n20170), .B2(n20823), .ZN(
        n15937) );
  INV_X1 U19080 ( .A(n15937), .ZN(n15941) );
  AOI22_X1 U19081 ( .A1(n15939), .A2(n20188), .B1(n20203), .B2(n15938), .ZN(
        n15940) );
  OAI211_X1 U19082 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15942), .A(
        n15941), .B(n15940), .ZN(P1_U3012) );
  AOI21_X1 U19083 ( .B1(n15943), .B2(n16001), .A(n15964), .ZN(n15959) );
  NOR2_X1 U19084 ( .A1(n20170), .A2(n20821), .ZN(n15947) );
  OAI22_X1 U19085 ( .A1(n15945), .A2(n20208), .B1(n16014), .B2(n15944), .ZN(
        n15946) );
  AOI211_X1 U19086 ( .C1(n15948), .C2(n15950), .A(n15947), .B(n15946), .ZN(
        n15949) );
  OAI21_X1 U19087 ( .B1(n15959), .B2(n15950), .A(n15949), .ZN(P1_U3013) );
  INV_X1 U19088 ( .A(n15967), .ZN(n15952) );
  AOI21_X1 U19089 ( .B1(n15952), .B2(n15951), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15958) );
  INV_X1 U19090 ( .A(n15953), .ZN(n15955) );
  AOI22_X1 U19091 ( .A1(n15955), .A2(n20188), .B1(n20203), .B2(n15954), .ZN(
        n15957) );
  NAND2_X1 U19092 ( .A1(n20190), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15956) );
  OAI211_X1 U19093 ( .C1(n15959), .C2(n15958), .A(n15957), .B(n15956), .ZN(
        P1_U3014) );
  INV_X1 U19094 ( .A(n15960), .ZN(n15961) );
  AOI21_X1 U19095 ( .B1(n15962), .B2(n20203), .A(n15961), .ZN(n15966) );
  AOI22_X1 U19096 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n15964), .B1(
        n20188), .B2(n15963), .ZN(n15965) );
  OAI211_X1 U19097 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15967), .A(
        n15966), .B(n15965), .ZN(P1_U3016) );
  AOI21_X1 U19098 ( .B1(n15969), .B2(n20203), .A(n15968), .ZN(n15973) );
  AOI22_X1 U19099 ( .A1(n15971), .A2(n20188), .B1(n12499), .B2(n15970), .ZN(
        n15972) );
  OAI211_X1 U19100 ( .C1(n15974), .C2(n12499), .A(n15973), .B(n15972), .ZN(
        P1_U3018) );
  NOR2_X1 U19101 ( .A1(n15975), .A2(n15978), .ZN(n15984) );
  AOI22_X1 U19102 ( .A1(n20185), .A2(n15978), .B1(n15977), .B2(n15976), .ZN(
        n15979) );
  NAND2_X1 U19103 ( .A1(n15980), .A2(n15979), .ZN(n15993) );
  AOI21_X1 U19104 ( .B1(n20192), .B2(n15981), .A(n15993), .ZN(n15982) );
  INV_X1 U19105 ( .A(n15982), .ZN(n15983) );
  MUX2_X1 U19106 ( .A(n15984), .B(n15983), .S(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n15988) );
  INV_X1 U19107 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20809) );
  NAND2_X1 U19108 ( .A1(n15985), .A2(n20203), .ZN(n15986) );
  OAI21_X1 U19109 ( .B1(n20809), .B2(n20170), .A(n15986), .ZN(n15987) );
  NOR2_X1 U19110 ( .A1(n15988), .A2(n15987), .ZN(n15989) );
  OAI21_X1 U19111 ( .B1(n15990), .B2(n20208), .A(n15989), .ZN(P1_U3019) );
  AOI22_X1 U19112 ( .A1(n15991), .A2(n20203), .B1(n20190), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n15995) );
  AOI22_X1 U19113 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15993), .B1(
        n20188), .B2(n15992), .ZN(n15994) );
  OAI211_X1 U19114 ( .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15996), .A(
        n15995), .B(n15994), .ZN(P1_U3020) );
  AOI21_X1 U19115 ( .B1(n16034), .B2(n15998), .A(n15997), .ZN(n16002) );
  AOI221_X1 U19116 ( .B1(n16002), .B2(n16001), .C1(n16000), .C2(n16001), .A(
        n15999), .ZN(n16020) );
  NAND2_X1 U19117 ( .A1(n16003), .A2(n16027), .ZN(n16009) );
  AOI221_X1 U19118 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n12391), .C2(n16019), .A(
        n16009), .ZN(n16006) );
  OAI22_X1 U19119 ( .A1(n16004), .A2(n16014), .B1(n20806), .B2(n20170), .ZN(
        n16005) );
  AOI211_X1 U19120 ( .C1(n16007), .C2(n20188), .A(n16006), .B(n16005), .ZN(
        n16008) );
  OAI21_X1 U19121 ( .B1(n16020), .B2(n12391), .A(n16008), .ZN(P1_U3021) );
  NOR2_X1 U19122 ( .A1(n16009), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16016) );
  OR2_X1 U19123 ( .A1(n16011), .A2(n16010), .ZN(n16012) );
  NAND2_X1 U19124 ( .A1(n16013), .A2(n16012), .ZN(n20003) );
  OAI22_X1 U19125 ( .A1(n20003), .A2(n16014), .B1(n20804), .B2(n20170), .ZN(
        n16015) );
  AOI211_X1 U19126 ( .C1(n16017), .C2(n20188), .A(n16016), .B(n16015), .ZN(
        n16018) );
  OAI21_X1 U19127 ( .B1(n16020), .B2(n16019), .A(n16018), .ZN(P1_U3022) );
  INV_X1 U19128 ( .A(n16021), .ZN(n16024) );
  INV_X1 U19129 ( .A(n16022), .ZN(n16023) );
  OAI21_X1 U19130 ( .B1(n16042), .B2(n16024), .A(n16023), .ZN(n16025) );
  AND2_X1 U19131 ( .A1(n16026), .A2(n16025), .ZN(n20065) );
  AOI22_X1 U19132 ( .A1(n20203), .A2(n20065), .B1(n20190), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16030) );
  AOI22_X1 U19133 ( .A1(n16028), .A2(n20188), .B1(n16031), .B2(n16027), .ZN(
        n16029) );
  OAI211_X1 U19134 ( .C1(n16032), .C2(n16031), .A(n16030), .B(n16029), .ZN(
        P1_U3024) );
  NAND2_X1 U19135 ( .A1(n16034), .A2(n16033), .ZN(n16038) );
  AOI22_X1 U19136 ( .A1(n20203), .A2(n20035), .B1(n20190), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n16037) );
  AOI22_X1 U19137 ( .A1(n16035), .A2(n20188), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16043), .ZN(n16036) );
  OAI211_X1 U19138 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16038), .A(
        n16037), .B(n16036), .ZN(P1_U3025) );
  NAND2_X1 U19139 ( .A1(n16040), .A2(n16039), .ZN(n16041) );
  AND2_X1 U19140 ( .A1(n16042), .A2(n16041), .ZN(n20069) );
  AOI22_X1 U19141 ( .A1(n20203), .A2(n20069), .B1(n20190), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n16049) );
  AOI22_X1 U19142 ( .A1(n16044), .A2(n20188), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16043), .ZN(n16048) );
  NAND3_X1 U19143 ( .A1(n16046), .A2(n20176), .A3(n16045), .ZN(n16047) );
  NAND3_X1 U19144 ( .A1(n16049), .A2(n16048), .A3(n16047), .ZN(P1_U3026) );
  OAI221_X1 U19145 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATEBS16_REG_SCAN_IN), .C1(n16055), .C2(n20871), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n20777) );
  NAND2_X1 U19146 ( .A1(n16054), .A2(n20777), .ZN(n16050) );
  AOI22_X1 U19147 ( .A1(n16053), .A2(n16052), .B1(n16051), .B2(n16050), .ZN(
        P1_U3162) );
  OAI22_X1 U19148 ( .A1(n20776), .A2(n20590), .B1(n16055), .B2(n16054), .ZN(
        P1_U3466) );
  AOI21_X1 U19149 ( .B1(n16058), .B2(n16057), .A(n16056), .ZN(n16066) );
  INV_X1 U19150 ( .A(n15308), .ZN(n16062) );
  AOI22_X1 U19151 ( .A1(n19054), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19068), .ZN(n16059) );
  OAI21_X1 U19152 ( .B1(n19017), .B2(n16060), .A(n16059), .ZN(n16061) );
  AOI21_X1 U19153 ( .B1(n16062), .B2(n19062), .A(n16061), .ZN(n16063) );
  OAI21_X1 U19154 ( .B1(n16064), .B2(n9646), .A(n16063), .ZN(n16065) );
  AOI21_X1 U19155 ( .B1(n19049), .B2(n16066), .A(n16065), .ZN(n16067) );
  OAI21_X1 U19156 ( .B1(n16068), .B2(n19053), .A(n16067), .ZN(P2_U2826) );
  AOI211_X1 U19157 ( .C1(n16071), .C2(n16070), .A(n16069), .B(n19822), .ZN(
        n16080) );
  INV_X1 U19158 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16072) );
  OAI22_X1 U19159 ( .A1(n19035), .A2(n16073), .B1(n16072), .B2(n19006), .ZN(
        n16076) );
  NOR2_X1 U19160 ( .A1(n16074), .A2(n19036), .ZN(n16075) );
  AOI211_X1 U19161 ( .C1(P2_EBX_REG_26__SCAN_IN), .C2(n19055), .A(n16076), .B(
        n16075), .ZN(n16077) );
  OAI21_X1 U19162 ( .B1(n16078), .B2(n9646), .A(n16077), .ZN(n16079) );
  AOI211_X1 U19163 ( .C1(n19056), .C2(n16081), .A(n16080), .B(n16079), .ZN(
        n16082) );
  INV_X1 U19164 ( .A(n16082), .ZN(P2_U2829) );
  AOI22_X1 U19165 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19068), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19054), .ZN(n16094) );
  INV_X1 U19166 ( .A(n16083), .ZN(n16084) );
  AOI22_X1 U19167 ( .A1(n16084), .A2(n19031), .B1(P2_EBX_REG_24__SCAN_IN), 
        .B2(n19055), .ZN(n16093) );
  OAI22_X1 U19168 ( .A1(n16086), .A2(n19036), .B1(n19053), .B2(n16085), .ZN(
        n16087) );
  INV_X1 U19169 ( .A(n16087), .ZN(n16092) );
  AOI21_X1 U19170 ( .B1(n16089), .B2(n9765), .A(n16088), .ZN(n16090) );
  NAND2_X1 U19171 ( .A1(n19049), .A2(n16090), .ZN(n16091) );
  NAND4_X1 U19172 ( .A1(n16094), .A2(n16093), .A3(n16092), .A4(n16091), .ZN(
        P2_U2831) );
  AOI22_X1 U19173 ( .A1(n19077), .A2(n16095), .B1(n19130), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16101) );
  AOI22_X1 U19174 ( .A1(n19079), .A2(BUF1_REG_20__SCAN_IN), .B1(n19078), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16100) );
  INV_X1 U19175 ( .A(n16096), .ZN(n16097) );
  AOI22_X1 U19176 ( .A1(n16098), .A2(n19085), .B1(n19131), .B2(n16097), .ZN(
        n16099) );
  NAND3_X1 U19177 ( .A1(n16101), .A2(n16100), .A3(n16099), .ZN(P2_U2899) );
  AOI22_X1 U19178 ( .A1(n19077), .A2(n16102), .B1(n19130), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16106) );
  AOI22_X1 U19179 ( .A1(n19079), .A2(BUF1_REG_18__SCAN_IN), .B1(n19078), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16105) );
  AOI22_X1 U19180 ( .A1(n16103), .A2(n19085), .B1(n19131), .B2(n16228), .ZN(
        n16104) );
  NAND3_X1 U19181 ( .A1(n16106), .A2(n16105), .A3(n16104), .ZN(P2_U2901) );
  AOI22_X1 U19182 ( .A1(n19187), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19192), .ZN(n16111) );
  AOI222_X1 U19183 ( .A1(n16109), .A2(n19188), .B1(n19194), .B2(n16108), .C1(
        n11014), .C2(n16107), .ZN(n16110) );
  OAI211_X1 U19184 ( .C1(n19182), .C2(n16112), .A(n16111), .B(n16110), .ZN(
        P2_U2992) );
  AOI22_X1 U19185 ( .A1(n19187), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19192), .ZN(n16123) );
  INV_X1 U19186 ( .A(n16114), .ZN(n16117) );
  AND2_X1 U19187 ( .A1(n16114), .A2(n16113), .ZN(n16116) );
  OAI22_X1 U19188 ( .A1(n16118), .A2(n16117), .B1(n16116), .B2(n16115), .ZN(
        n16233) );
  OR2_X1 U19189 ( .A1(n16120), .A2(n16119), .ZN(n16125) );
  AOI21_X1 U19190 ( .B1(n16125), .B2(n16229), .A(n16121), .ZN(n16231) );
  AOI222_X1 U19191 ( .A1(n16233), .A2(n19188), .B1(n19194), .B2(n16232), .C1(
        n11014), .C2(n16231), .ZN(n16122) );
  OAI211_X1 U19192 ( .C1(n19182), .C2(n16124), .A(n16123), .B(n16122), .ZN(
        P2_U2996) );
  INV_X1 U19193 ( .A(n16125), .ZN(n16126) );
  AOI211_X1 U19194 ( .C1(n10893), .C2(n16127), .A(n16207), .B(n16126), .ZN(
        n16133) );
  AOI21_X1 U19195 ( .B1(n19187), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n16128), .ZN(n16130) );
  NAND2_X1 U19196 ( .A1(n18951), .A2(n19195), .ZN(n16129) );
  OAI211_X1 U19197 ( .C1(n16131), .C2(n16209), .A(n16130), .B(n16129), .ZN(
        n16132) );
  AOI211_X1 U19198 ( .C1(n18950), .C2(n19194), .A(n16133), .B(n16132), .ZN(
        n16134) );
  INV_X1 U19199 ( .A(n16134), .ZN(P2_U2997) );
  AOI22_X1 U19200 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19192), .B1(n19195), 
        .B2(n18963), .ZN(n16139) );
  OAI22_X1 U19201 ( .A1(n16136), .A2(n16209), .B1(n16207), .B2(n16135), .ZN(
        n16137) );
  AOI21_X1 U19202 ( .B1(n19194), .B2(n18957), .A(n16137), .ZN(n16138) );
  OAI211_X1 U19203 ( .C1(n16227), .C2(n18960), .A(n16139), .B(n16138), .ZN(
        P2_U2999) );
  AOI22_X1 U19204 ( .A1(n19187), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19192), .ZN(n16144) );
  INV_X1 U19205 ( .A(n16140), .ZN(n18977) );
  AOI222_X1 U19206 ( .A1(n16142), .A2(n19188), .B1(n19194), .B2(n18977), .C1(
        n11014), .C2(n16141), .ZN(n16143) );
  OAI211_X1 U19207 ( .C1(n19182), .C2(n18972), .A(n16144), .B(n16143), .ZN(
        P2_U3000) );
  AOI22_X1 U19208 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19192), .B1(n19195), 
        .B2(n18987), .ZN(n16149) );
  OAI22_X1 U19209 ( .A1(n16146), .A2(n16209), .B1(n16207), .B2(n16145), .ZN(
        n16147) );
  AOI21_X1 U19210 ( .B1(n19194), .B2(n18988), .A(n16147), .ZN(n16148) );
  OAI211_X1 U19211 ( .C1(n16227), .C2(n16150), .A(n16149), .B(n16148), .ZN(
        P2_U3001) );
  AOI22_X1 U19212 ( .A1(n19187), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19174), .ZN(n16157) );
  NOR2_X1 U19213 ( .A1(n9903), .A2(n16151), .ZN(n16152) );
  XNOR2_X1 U19214 ( .A(n16153), .B(n16152), .ZN(n16252) );
  OAI21_X1 U19215 ( .B1(n16165), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n16154), .ZN(n16247) );
  OAI222_X1 U19216 ( .A1(n16248), .A2(n19218), .B1(n16209), .B2(n16252), .C1(
        n16207), .C2(n16247), .ZN(n16155) );
  INV_X1 U19217 ( .A(n16155), .ZN(n16156) );
  OAI211_X1 U19218 ( .C1(n19182), .C2(n18994), .A(n16157), .B(n16156), .ZN(
        P2_U3002) );
  AOI22_X1 U19219 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19192), .B1(n19195), 
        .B2(n19010), .ZN(n16170) );
  INV_X1 U19220 ( .A(n16261), .ZN(n19011) );
  NOR2_X1 U19221 ( .A1(n16159), .A2(n16158), .ZN(n16163) );
  NAND2_X1 U19222 ( .A1(n16161), .A2(n16160), .ZN(n16162) );
  XNOR2_X1 U19223 ( .A(n16163), .B(n16162), .ZN(n16266) );
  NAND2_X1 U19224 ( .A1(n16164), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16181) );
  AOI21_X1 U19225 ( .B1(n16181), .B2(n16166), .A(n16165), .ZN(n16263) );
  INV_X1 U19226 ( .A(n16263), .ZN(n16167) );
  OAI22_X1 U19227 ( .A1(n16266), .A2(n16209), .B1(n16167), .B2(n16207), .ZN(
        n16168) );
  AOI21_X1 U19228 ( .B1(n19194), .B2(n19011), .A(n16168), .ZN(n16169) );
  OAI211_X1 U19229 ( .C1(n16227), .C2(n16171), .A(n16170), .B(n16169), .ZN(
        P2_U3003) );
  AOI22_X1 U19230 ( .A1(n19187), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19192), .ZN(n16184) );
  NAND2_X1 U19231 ( .A1(n16173), .A2(n16172), .ZN(n16178) );
  INV_X1 U19232 ( .A(n16174), .ZN(n16175) );
  NOR2_X1 U19233 ( .A1(n16176), .A2(n16175), .ZN(n16177) );
  XNOR2_X1 U19234 ( .A(n16178), .B(n16177), .ZN(n16276) );
  INV_X1 U19235 ( .A(n16276), .ZN(n16182) );
  NAND2_X1 U19236 ( .A1(n16179), .A2(n16269), .ZN(n16180) );
  AOI222_X1 U19237 ( .A1(n16182), .A2(n19188), .B1(n19194), .B2(n16272), .C1(
        n11014), .C2(n16273), .ZN(n16183) );
  OAI211_X1 U19238 ( .C1(n19182), .C2(n16185), .A(n16184), .B(n16183), .ZN(
        P2_U3004) );
  AOI22_X1 U19239 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19192), .B1(n19195), 
        .B2(n19023), .ZN(n16190) );
  OAI22_X1 U19240 ( .A1(n16187), .A2(n16207), .B1(n16209), .B2(n16186), .ZN(
        n16188) );
  AOI21_X1 U19241 ( .B1(n19194), .B2(n19024), .A(n16188), .ZN(n16189) );
  OAI211_X1 U19242 ( .C1(n16227), .C2(n16191), .A(n16190), .B(n16189), .ZN(
        P2_U3005) );
  AOI22_X1 U19243 ( .A1(n19187), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19192), .ZN(n16205) );
  INV_X1 U19244 ( .A(n16192), .ZN(n16193) );
  XNOR2_X1 U19245 ( .A(n16194), .B(n16193), .ZN(n16279) );
  NAND2_X1 U19246 ( .A1(n16279), .A2(n11014), .ZN(n16202) );
  NAND2_X1 U19247 ( .A1(n15259), .A2(n16195), .ZN(n16200) );
  INV_X1 U19248 ( .A(n16196), .ZN(n16197) );
  NOR2_X1 U19249 ( .A1(n16198), .A2(n16197), .ZN(n16199) );
  XNOR2_X1 U19250 ( .A(n16200), .B(n16199), .ZN(n16283) );
  NAND2_X1 U19251 ( .A1(n16283), .A2(n19188), .ZN(n16201) );
  OAI211_X1 U19252 ( .C1(n19218), .C2(n16280), .A(n16202), .B(n16201), .ZN(
        n16203) );
  INV_X1 U19253 ( .A(n16203), .ZN(n16204) );
  OAI211_X1 U19254 ( .C1(n19182), .C2(n16206), .A(n16205), .B(n16204), .ZN(
        P2_U3006) );
  AOI22_X1 U19255 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19192), .B1(n19195), 
        .B2(n19047), .ZN(n16213) );
  OAI22_X1 U19256 ( .A1(n16210), .A2(n16209), .B1(n16208), .B2(n16207), .ZN(
        n16211) );
  AOI21_X1 U19257 ( .B1(n19194), .B2(n19048), .A(n16211), .ZN(n16212) );
  OAI211_X1 U19258 ( .C1(n16227), .C2(n16214), .A(n16213), .B(n16212), .ZN(
        P2_U3009) );
  AOI22_X1 U19259 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n19192), .B1(n19195), 
        .B2(n16215), .ZN(n16226) );
  OAI21_X1 U19260 ( .B1(n16218), .B2(n16217), .A(n16216), .ZN(n16219) );
  INV_X1 U19261 ( .A(n16219), .ZN(n16302) );
  NAND2_X1 U19262 ( .A1(n16221), .A2(n16220), .ZN(n16224) );
  XNOR2_X1 U19263 ( .A(n16222), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n16223) );
  XNOR2_X1 U19264 ( .A(n16224), .B(n16223), .ZN(n16308) );
  OAI211_X1 U19265 ( .C1(n12656), .C2(n16227), .A(n16226), .B(n16225), .ZN(
        P2_U3011) );
  AOI22_X1 U19266 ( .A1(n16230), .A2(n16229), .B1(n16228), .B2(n19202), .ZN(
        n16239) );
  AOI222_X1 U19267 ( .A1(n16233), .A2(n16309), .B1(n16303), .B2(n16232), .C1(
        n19204), .C2(n16231), .ZN(n16238) );
  NAND2_X1 U19268 ( .A1(P2_REIP_REG_18__SCAN_IN), .A2(n19192), .ZN(n16237) );
  OAI221_X1 U19269 ( .B1(n16235), .B2(n16234), .C1(n16235), .C2(n19201), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16236) );
  NAND4_X1 U19270 ( .A1(n16239), .A2(n16238), .A3(n16237), .A4(n16236), .ZN(
        P2_U3028) );
  AOI21_X1 U19271 ( .B1(n16254), .B2(n16241), .A(n16240), .ZN(n19094) );
  INV_X1 U19272 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19856) );
  NOR2_X1 U19273 ( .A1(n19033), .A2(n19856), .ZN(n16246) );
  INV_X1 U19274 ( .A(n16242), .ZN(n16243) );
  AOI21_X1 U19275 ( .B1(n11046), .B2(n16244), .A(n16243), .ZN(n16245) );
  AOI211_X1 U19276 ( .C1(n19202), .C2(n19094), .A(n16246), .B(n16245), .ZN(
        n16251) );
  INV_X1 U19277 ( .A(n16247), .ZN(n16249) );
  INV_X1 U19278 ( .A(n16248), .ZN(n19000) );
  AOI22_X1 U19279 ( .A1(n16249), .A2(n19204), .B1(n16303), .B2(n19000), .ZN(
        n16250) );
  OAI211_X1 U19280 ( .C1(n16252), .C2(n19209), .A(n16251), .B(n16250), .ZN(
        P2_U3034) );
  NAND2_X1 U19281 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16253), .ZN(
        n16270) );
  AOI221_X1 U19282 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C1(n16269), .C2(n16166), .A(
        n16270), .ZN(n16260) );
  OAI21_X1 U19283 ( .B1(n16256), .B2(n16255), .A(n16254), .ZN(n19099) );
  OAI21_X1 U19284 ( .B1(n16258), .B2(n10843), .A(n16257), .ZN(n16268) );
  OAI22_X1 U19285 ( .A1(n19099), .A2(n16306), .B1(n16166), .B2(n16268), .ZN(
        n16259) );
  AOI211_X1 U19286 ( .C1(n19174), .C2(P2_REIP_REG_11__SCAN_IN), .A(n16260), 
        .B(n16259), .ZN(n16265) );
  NOR2_X1 U19287 ( .A1(n19206), .A2(n16261), .ZN(n16262) );
  AOI21_X1 U19288 ( .B1(n16263), .B2(n19204), .A(n16262), .ZN(n16264) );
  OAI211_X1 U19289 ( .C1(n16266), .C2(n19209), .A(n16265), .B(n16264), .ZN(
        P2_U3035) );
  NAND2_X1 U19290 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19192), .ZN(n16267) );
  OAI221_X1 U19291 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16270), 
        .C1(n16269), .C2(n16268), .A(n16267), .ZN(n16271) );
  AOI21_X1 U19292 ( .B1(n19202), .B2(n19100), .A(n16271), .ZN(n16275) );
  AOI22_X1 U19293 ( .A1(n16273), .A2(n19204), .B1(n16303), .B2(n16272), .ZN(
        n16274) );
  OAI211_X1 U19294 ( .C1(n16276), .C2(n19209), .A(n16275), .B(n16274), .ZN(
        P2_U3036) );
  NOR2_X1 U19295 ( .A1(n16278), .A2(n16277), .ZN(n16295) );
  AOI22_X1 U19296 ( .A1(n16295), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19202), .B2(n19106), .ZN(n16288) );
  INV_X1 U19297 ( .A(n16279), .ZN(n16281) );
  OAI22_X1 U19298 ( .A1(n16281), .A2(n16301), .B1(n19206), .B2(n16280), .ZN(
        n16282) );
  AOI21_X1 U19299 ( .B1(n16309), .B2(n16283), .A(n16282), .ZN(n16287) );
  NAND2_X1 U19300 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19192), .ZN(n16286) );
  OAI211_X1 U19301 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16294), .B(n16284), .ZN(n16285) );
  NAND4_X1 U19302 ( .A1(n16288), .A2(n16287), .A3(n16286), .A4(n16285), .ZN(
        P2_U3038) );
  OAI21_X1 U19303 ( .B1(n16291), .B2(n16290), .A(n16289), .ZN(n19111) );
  OAI22_X1 U19304 ( .A1(n16306), .A2(n19111), .B1(n19848), .B2(n19033), .ZN(
        n16292) );
  AOI221_X1 U19305 ( .B1(n16295), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(
        n16294), .C2(n16293), .A(n16292), .ZN(n16299) );
  INV_X1 U19306 ( .A(n19037), .ZN(n16296) );
  AOI22_X1 U19307 ( .A1(n16297), .A2(n16309), .B1(n16303), .B2(n16296), .ZN(
        n16298) );
  OAI211_X1 U19308 ( .C1(n16301), .C2(n16300), .A(n16299), .B(n16298), .ZN(
        P2_U3039) );
  NAND2_X1 U19309 ( .A1(n16302), .A2(n19204), .ZN(n16305) );
  OAI211_X1 U19310 ( .C1(n19898), .C2(n16306), .A(n16305), .B(n16304), .ZN(
        n16307) );
  AOI21_X1 U19311 ( .B1(n16309), .B2(n16308), .A(n16307), .ZN(n16310) );
  OAI221_X1 U19312 ( .B1(n16312), .B2(n10175), .C1(n16312), .C2(n16311), .A(
        n16310), .ZN(P2_U3043) );
  NAND2_X1 U19313 ( .A1(n16323), .A2(n16352), .ZN(n16314) );
  OR2_X1 U19314 ( .A1(n16352), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16313) );
  NAND2_X1 U19315 ( .A1(n16314), .A2(n16313), .ZN(n16331) );
  NAND2_X1 U19316 ( .A1(n16315), .A2(n16352), .ZN(n16317) );
  OR2_X1 U19317 ( .A1(n16352), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16316) );
  NAND2_X1 U19318 ( .A1(n16317), .A2(n16316), .ZN(n16332) );
  OR2_X1 U19319 ( .A1(n16332), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n16324) );
  OR2_X1 U19320 ( .A1(n16324), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n16328) );
  NAND2_X1 U19321 ( .A1(n16321), .A2(n19929), .ZN(n16319) );
  NAND3_X1 U19322 ( .A1(n16319), .A2(n16318), .A3(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n16320) );
  OAI211_X1 U19323 ( .C1(n19929), .C2(n16321), .A(n16320), .B(n16352), .ZN(
        n16322) );
  AOI21_X1 U19324 ( .B1(n16323), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n16322), .ZN(n16326) );
  NAND2_X1 U19325 ( .A1(n16324), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n16325) );
  NAND2_X1 U19326 ( .A1(n16326), .A2(n16325), .ZN(n16327) );
  OAI211_X1 U19327 ( .C1(n16331), .C2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n16328), .B(n16327), .ZN(n16330) );
  NAND2_X1 U19328 ( .A1(n16330), .A2(n16329), .ZN(n16357) );
  INV_X1 U19329 ( .A(n16331), .ZN(n16355) );
  INV_X1 U19330 ( .A(n16332), .ZN(n16354) );
  INV_X1 U19331 ( .A(n16333), .ZN(n16334) );
  NAND2_X1 U19332 ( .A1(n16335), .A2(n16334), .ZN(n16338) );
  NAND2_X1 U19333 ( .A1(n16340), .A2(n16336), .ZN(n16337) );
  OAI211_X1 U19334 ( .C1(n16340), .C2(n16339), .A(n16338), .B(n16337), .ZN(
        n19950) );
  NOR2_X1 U19335 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P2_MORE_REG_SCAN_IN), .ZN(
        n16347) );
  NAND2_X1 U19336 ( .A1(n13380), .A2(n16341), .ZN(n16344) );
  OAI22_X1 U19337 ( .A1(n13347), .A2(n16344), .B1(n16343), .B2(n16342), .ZN(
        n16345) );
  INV_X1 U19338 ( .A(n16345), .ZN(n16346) );
  OAI21_X1 U19339 ( .B1(n16348), .B2(n16347), .A(n16346), .ZN(n16349) );
  NOR2_X1 U19340 ( .A1(n19950), .A2(n16349), .ZN(n16350) );
  OAI21_X1 U19341 ( .B1(n16352), .B2(n16351), .A(n16350), .ZN(n16353) );
  AOI21_X1 U19342 ( .B1(n16355), .B2(n16354), .A(n16353), .ZN(n16356) );
  NAND2_X1 U19343 ( .A1(n16357), .A2(n16356), .ZN(n16363) );
  AOI211_X1 U19344 ( .C1(n19819), .C2(n16363), .A(n16359), .B(n16358), .ZN(
        n16368) );
  NAND2_X1 U19345 ( .A1(n19964), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16360) );
  AOI21_X1 U19346 ( .B1(n10593), .B2(n16361), .A(n16360), .ZN(n16364) );
  AOI22_X1 U19347 ( .A1(n16362), .A2(n19961), .B1(n19960), .B2(n16364), .ZN(
        n16366) );
  OAI21_X1 U19348 ( .B1(n16363), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n16365) );
  AND2_X1 U19349 ( .A1(n16365), .A2(n16364), .ZN(n19815) );
  INV_X1 U19350 ( .A(n19815), .ZN(n19817) );
  NAND2_X1 U19351 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19817), .ZN(n16372) );
  OAI21_X1 U19352 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16366), .A(n16372), 
        .ZN(n16367) );
  OAI211_X1 U19353 ( .C1(n16370), .C2(n16369), .A(n16368), .B(n16367), .ZN(
        P2_U3176) );
  AOI21_X1 U19354 ( .B1(n16372), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n16371), 
        .ZN(n16373) );
  INV_X1 U19355 ( .A(n16373), .ZN(P2_U3593) );
  OAI22_X1 U19356 ( .A1(n16400), .A2(n17901), .B1(n16387), .B2(n17809), .ZN(
        n16379) );
  INV_X1 U19357 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16555) );
  OAI21_X1 U19358 ( .B1(n16391), .B2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n16374), .ZN(n16553) );
  OAI22_X1 U19359 ( .A1(n16375), .A2(n16555), .B1(n17746), .B2(n16553), .ZN(
        n16378) );
  INV_X1 U19360 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18839) );
  OAI22_X1 U19361 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16376), .B1(
        n18217), .B2(n18839), .ZN(n16377) );
  AOI211_X1 U19362 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n16379), .A(
        n16378), .B(n16377), .ZN(n16385) );
  NAND3_X1 U19363 ( .A1(n16380), .A2(n18072), .A3(n17773), .ZN(n17696) );
  NOR2_X1 U19364 ( .A1(n16381), .A2(n17696), .ZN(n17562) );
  NAND4_X1 U19365 ( .A1(n16383), .A2(n17558), .A3(n16382), .A4(n17562), .ZN(
        n16384) );
  OAI211_X1 U19366 ( .C1(n16386), .C2(n17780), .A(n16385), .B(n16384), .ZN(
        P3_U2800) );
  AOI211_X1 U19367 ( .C1(n16389), .C2(n16388), .A(n16387), .B(n17809), .ZN(
        n16398) );
  INV_X1 U19368 ( .A(n16390), .ZN(n16539) );
  AOI21_X1 U19369 ( .B1(n16574), .B2(n16539), .A(n16391), .ZN(n16568) );
  OAI21_X1 U19370 ( .B1(n17644), .B2(n16392), .A(n16568), .ZN(n16393) );
  OAI211_X1 U19371 ( .C1(n16396), .C2(n16395), .A(n16394), .B(n16393), .ZN(
        n16397) );
  AOI211_X1 U19372 ( .C1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n16399), .A(
        n16398), .B(n16397), .ZN(n16404) );
  NOR2_X1 U19373 ( .A1(n16400), .A2(n17901), .ZN(n16401) );
  OAI21_X1 U19374 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16402), .A(
        n16401), .ZN(n16403) );
  OAI211_X1 U19375 ( .C1(n16405), .C2(n17780), .A(n16404), .B(n16403), .ZN(
        P3_U2801) );
  NOR3_X1 U19376 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16407) );
  NOR4_X1 U19377 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16406) );
  NAND4_X1 U19378 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16407), .A3(n16406), .A4(
        U215), .ZN(U213) );
  INV_X1 U19379 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16497) );
  INV_X2 U19380 ( .A(U214), .ZN(n16459) );
  INV_X1 U19381 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16498) );
  OAI222_X1 U19382 ( .A1(U212), .A2(n16497), .B1(n16461), .B2(n16409), .C1(
        U214), .C2(n16498), .ZN(U216) );
  AOI22_X1 U19383 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16446), .ZN(n16410) );
  OAI21_X1 U19384 ( .B1(n14237), .B2(n16461), .A(n16410), .ZN(U217) );
  INV_X1 U19385 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20234) );
  AOI22_X1 U19386 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16446), .ZN(n16411) );
  OAI21_X1 U19387 ( .B1(n20234), .B2(n16461), .A(n16411), .ZN(U218) );
  AOI22_X1 U19388 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16446), .ZN(n16412) );
  OAI21_X1 U19389 ( .B1(n16413), .B2(n16461), .A(n16412), .ZN(U219) );
  INV_X1 U19390 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20226) );
  AOI22_X1 U19391 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16446), .ZN(n16414) );
  OAI21_X1 U19392 ( .B1(n20226), .B2(n16461), .A(n16414), .ZN(U220) );
  AOI22_X1 U19393 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16446), .ZN(n16415) );
  OAI21_X1 U19394 ( .B1(n14494), .B2(n16461), .A(n16415), .ZN(U221) );
  AOI22_X1 U19395 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16446), .ZN(n16416) );
  OAI21_X1 U19396 ( .B1(n20219), .B2(n16461), .A(n16416), .ZN(U222) );
  INV_X1 U19397 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20211) );
  AOI22_X1 U19398 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16446), .ZN(n16417) );
  OAI21_X1 U19399 ( .B1(n20211), .B2(n16461), .A(n16417), .ZN(U223) );
  AOI22_X1 U19400 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16446), .ZN(n16418) );
  OAI21_X1 U19401 ( .B1(n16419), .B2(n16461), .A(n16418), .ZN(U224) );
  INV_X1 U19402 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20249) );
  AOI22_X1 U19403 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16446), .ZN(n16420) );
  OAI21_X1 U19404 ( .B1(n20249), .B2(n16461), .A(n16420), .ZN(U225) );
  INV_X1 U19405 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20238) );
  AOI22_X1 U19406 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16446), .ZN(n16421) );
  OAI21_X1 U19407 ( .B1(n20238), .B2(n16461), .A(n16421), .ZN(U226) );
  AOI22_X1 U19408 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16446), .ZN(n16422) );
  OAI21_X1 U19409 ( .B1(n16423), .B2(n16461), .A(n16422), .ZN(U227) );
  INV_X1 U19410 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20229) );
  AOI22_X1 U19411 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16446), .ZN(n16424) );
  OAI21_X1 U19412 ( .B1(n20229), .B2(n16461), .A(n16424), .ZN(U228) );
  AOI22_X1 U19413 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16446), .ZN(n16425) );
  OAI21_X1 U19414 ( .B1(n16426), .B2(n16461), .A(n16425), .ZN(U229) );
  INV_X1 U19415 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20223) );
  AOI22_X1 U19416 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16446), .ZN(n16427) );
  OAI21_X1 U19417 ( .B1(n20223), .B2(n16461), .A(n16427), .ZN(U230) );
  INV_X1 U19418 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20215) );
  AOI22_X1 U19419 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16446), .ZN(n16428) );
  OAI21_X1 U19420 ( .B1(n20215), .B2(n16461), .A(n16428), .ZN(U231) );
  AOI22_X1 U19421 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16446), .ZN(n16429) );
  OAI21_X1 U19422 ( .B1(n14548), .B2(n16461), .A(n16429), .ZN(U232) );
  INV_X1 U19423 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16431) );
  AOI22_X1 U19424 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16446), .ZN(n16430) );
  OAI21_X1 U19425 ( .B1(n16431), .B2(n16461), .A(n16430), .ZN(U233) );
  AOI22_X1 U19426 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16446), .ZN(n16432) );
  OAI21_X1 U19427 ( .B1(n16433), .B2(n16461), .A(n16432), .ZN(U234) );
  INV_X1 U19428 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16435) );
  AOI22_X1 U19429 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16446), .ZN(n16434) );
  OAI21_X1 U19430 ( .B1(n16435), .B2(n16461), .A(n16434), .ZN(U235) );
  AOI22_X1 U19431 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16446), .ZN(n16436) );
  OAI21_X1 U19432 ( .B1(n16437), .B2(n16461), .A(n16436), .ZN(U236) );
  INV_X1 U19433 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16439) );
  AOI22_X1 U19434 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16446), .ZN(n16438) );
  OAI21_X1 U19435 ( .B1(n16439), .B2(n16461), .A(n16438), .ZN(U237) );
  AOI22_X1 U19436 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16446), .ZN(n16440) );
  OAI21_X1 U19437 ( .B1(n16441), .B2(n16461), .A(n16440), .ZN(U238) );
  INV_X1 U19438 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16443) );
  AOI22_X1 U19439 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16446), .ZN(n16442) );
  OAI21_X1 U19440 ( .B1(n16443), .B2(n16461), .A(n16442), .ZN(U239) );
  INV_X1 U19441 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16445) );
  AOI22_X1 U19442 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16446), .ZN(n16444) );
  OAI21_X1 U19443 ( .B1(n16445), .B2(n16461), .A(n16444), .ZN(U240) );
  INV_X1 U19444 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16448) );
  AOI22_X1 U19445 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16446), .ZN(n16447) );
  OAI21_X1 U19446 ( .B1(n16448), .B2(n16461), .A(n16447), .ZN(U241) );
  INV_X1 U19447 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16450) );
  AOI22_X1 U19448 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16446), .ZN(n16449) );
  OAI21_X1 U19449 ( .B1(n16450), .B2(n16461), .A(n16449), .ZN(U242) );
  AOI22_X1 U19450 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16446), .ZN(n16451) );
  OAI21_X1 U19451 ( .B1(n16452), .B2(n16461), .A(n16451), .ZN(U243) );
  INV_X1 U19452 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16454) );
  AOI22_X1 U19453 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16446), .ZN(n16453) );
  OAI21_X1 U19454 ( .B1(n16454), .B2(n16461), .A(n16453), .ZN(U244) );
  AOI22_X1 U19455 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16446), .ZN(n16455) );
  OAI21_X1 U19456 ( .B1(n16456), .B2(n16461), .A(n16455), .ZN(U245) );
  AOI22_X1 U19457 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16446), .ZN(n16457) );
  OAI21_X1 U19458 ( .B1(n16458), .B2(n16461), .A(n16457), .ZN(U246) );
  AOI22_X1 U19459 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16459), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16446), .ZN(n16460) );
  OAI21_X1 U19460 ( .B1(n16462), .B2(n16461), .A(n16460), .ZN(U247) );
  INV_X1 U19461 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16463) );
  AOI22_X1 U19462 ( .A1(n16495), .A2(n16463), .B1(n18230), .B2(U215), .ZN(U251) );
  OAI22_X1 U19463 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16495), .ZN(n16464) );
  INV_X1 U19464 ( .A(n16464), .ZN(U252) );
  INV_X1 U19465 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16465) );
  AOI22_X1 U19466 ( .A1(n16495), .A2(n16465), .B1(n18240), .B2(U215), .ZN(U253) );
  INV_X1 U19467 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16466) );
  INV_X1 U19468 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18244) );
  AOI22_X1 U19469 ( .A1(n16495), .A2(n16466), .B1(n18244), .B2(U215), .ZN(U254) );
  INV_X1 U19470 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16467) );
  AOI22_X1 U19471 ( .A1(n16495), .A2(n16467), .B1(n18249), .B2(U215), .ZN(U255) );
  INV_X1 U19472 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16468) );
  INV_X1 U19473 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18253) );
  AOI22_X1 U19474 ( .A1(n16481), .A2(n16468), .B1(n18253), .B2(U215), .ZN(U256) );
  INV_X1 U19475 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16469) );
  INV_X1 U19476 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18258) );
  AOI22_X1 U19477 ( .A1(n16495), .A2(n16469), .B1(n18258), .B2(U215), .ZN(U257) );
  OAI22_X1 U19478 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16495), .ZN(n16470) );
  INV_X1 U19479 ( .A(n16470), .ZN(U258) );
  INV_X1 U19480 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16471) );
  INV_X1 U19481 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17510) );
  AOI22_X1 U19482 ( .A1(n16495), .A2(n16471), .B1(n17510), .B2(U215), .ZN(U259) );
  INV_X1 U19483 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16472) );
  INV_X1 U19484 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17512) );
  AOI22_X1 U19485 ( .A1(n16481), .A2(n16472), .B1(n17512), .B2(U215), .ZN(U260) );
  INV_X1 U19486 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16473) );
  INV_X1 U19487 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17514) );
  AOI22_X1 U19488 ( .A1(n16495), .A2(n16473), .B1(n17514), .B2(U215), .ZN(U261) );
  INV_X1 U19489 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16474) );
  INV_X1 U19490 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17517) );
  AOI22_X1 U19491 ( .A1(n16481), .A2(n16474), .B1(n17517), .B2(U215), .ZN(U262) );
  INV_X1 U19492 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16475) );
  INV_X1 U19493 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17522) );
  AOI22_X1 U19494 ( .A1(n16481), .A2(n16475), .B1(n17522), .B2(U215), .ZN(U263) );
  OAI22_X1 U19495 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16481), .ZN(n16476) );
  INV_X1 U19496 ( .A(n16476), .ZN(U264) );
  OAI22_X1 U19497 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16481), .ZN(n16477) );
  INV_X1 U19498 ( .A(n16477), .ZN(U265) );
  OAI22_X1 U19499 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16481), .ZN(n16478) );
  INV_X1 U19500 ( .A(n16478), .ZN(U266) );
  OAI22_X1 U19501 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16481), .ZN(n16479) );
  INV_X1 U19502 ( .A(n16479), .ZN(U267) );
  OAI22_X1 U19503 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16481), .ZN(n16480) );
  INV_X1 U19504 ( .A(n16480), .ZN(U268) );
  OAI22_X1 U19505 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16481), .ZN(n16482) );
  INV_X1 U19506 ( .A(n16482), .ZN(U269) );
  OAI22_X1 U19507 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16495), .ZN(n16483) );
  INV_X1 U19508 ( .A(n16483), .ZN(U270) );
  OAI22_X1 U19509 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16495), .ZN(n16484) );
  INV_X1 U19510 ( .A(n16484), .ZN(U271) );
  OAI22_X1 U19511 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16495), .ZN(n16485) );
  INV_X1 U19512 ( .A(n16485), .ZN(U272) );
  OAI22_X1 U19513 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16495), .ZN(n16486) );
  INV_X1 U19514 ( .A(n16486), .ZN(U273) );
  OAI22_X1 U19515 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16495), .ZN(n16487) );
  INV_X1 U19516 ( .A(n16487), .ZN(U274) );
  OAI22_X1 U19517 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16495), .ZN(n16488) );
  INV_X1 U19518 ( .A(n16488), .ZN(U275) );
  OAI22_X1 U19519 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16495), .ZN(n16489) );
  INV_X1 U19520 ( .A(n16489), .ZN(U276) );
  INV_X1 U19521 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n16490) );
  INV_X1 U19522 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n18239) );
  AOI22_X1 U19523 ( .A1(n16495), .A2(n16490), .B1(n18239), .B2(U215), .ZN(U277) );
  OAI22_X1 U19524 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16495), .ZN(n16491) );
  INV_X1 U19525 ( .A(n16491), .ZN(U278) );
  INV_X1 U19526 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n16492) );
  INV_X1 U19527 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n18248) );
  AOI22_X1 U19528 ( .A1(n16495), .A2(n16492), .B1(n18248), .B2(U215), .ZN(U279) );
  OAI22_X1 U19529 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16495), .ZN(n16493) );
  INV_X1 U19530 ( .A(n16493), .ZN(U280) );
  OAI22_X1 U19531 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16495), .ZN(n16494) );
  INV_X1 U19532 ( .A(n16494), .ZN(U281) );
  INV_X1 U19533 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18262) );
  AOI22_X1 U19534 ( .A1(n16495), .A2(n16497), .B1(n18262), .B2(U215), .ZN(U282) );
  INV_X1 U19535 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16496) );
  AOI222_X1 U19536 ( .A1(n16498), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16497), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16496), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16499) );
  INV_X2 U19537 ( .A(n16501), .ZN(n16500) );
  INV_X1 U19538 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18794) );
  INV_X1 U19539 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19853) );
  AOI22_X1 U19540 ( .A1(n16500), .A2(n18794), .B1(n19853), .B2(n16501), .ZN(
        U347) );
  INV_X1 U19541 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18792) );
  INV_X1 U19542 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19852) );
  AOI22_X1 U19543 ( .A1(n16500), .A2(n18792), .B1(n19852), .B2(n16501), .ZN(
        U348) );
  INV_X1 U19544 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18789) );
  INV_X1 U19545 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19851) );
  AOI22_X1 U19546 ( .A1(n16500), .A2(n18789), .B1(n19851), .B2(n16501), .ZN(
        U349) );
  INV_X1 U19547 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18788) );
  INV_X1 U19548 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19849) );
  AOI22_X1 U19549 ( .A1(n16500), .A2(n18788), .B1(n19849), .B2(n16501), .ZN(
        U350) );
  INV_X1 U19550 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18786) );
  INV_X1 U19551 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19847) );
  AOI22_X1 U19552 ( .A1(n16500), .A2(n18786), .B1(n19847), .B2(n16501), .ZN(
        U351) );
  INV_X1 U19553 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18784) );
  INV_X1 U19554 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19845) );
  AOI22_X1 U19555 ( .A1(n16500), .A2(n18784), .B1(n19845), .B2(n16501), .ZN(
        U352) );
  INV_X1 U19556 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18782) );
  INV_X1 U19557 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19844) );
  AOI22_X1 U19558 ( .A1(n16500), .A2(n18782), .B1(n19844), .B2(n16501), .ZN(
        U353) );
  INV_X1 U19559 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18780) );
  AOI22_X1 U19560 ( .A1(n16500), .A2(n18780), .B1(n19843), .B2(n16501), .ZN(
        U354) );
  INV_X1 U19561 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18835) );
  INV_X1 U19562 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19883) );
  AOI22_X1 U19563 ( .A1(n16500), .A2(n18835), .B1(n19883), .B2(n16501), .ZN(
        U356) );
  INV_X1 U19564 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18831) );
  INV_X1 U19565 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19881) );
  AOI22_X1 U19566 ( .A1(n16500), .A2(n18831), .B1(n19881), .B2(n16501), .ZN(
        U357) );
  INV_X1 U19567 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18829) );
  INV_X1 U19568 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19879) );
  AOI22_X1 U19569 ( .A1(n16500), .A2(n18829), .B1(n19879), .B2(n16501), .ZN(
        U358) );
  INV_X1 U19570 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18826) );
  INV_X1 U19571 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19878) );
  AOI22_X1 U19572 ( .A1(n16500), .A2(n18826), .B1(n19878), .B2(n16501), .ZN(
        U359) );
  INV_X1 U19573 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18824) );
  INV_X1 U19574 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19877) );
  AOI22_X1 U19575 ( .A1(n16500), .A2(n18824), .B1(n19877), .B2(n16501), .ZN(
        U360) );
  INV_X1 U19576 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18822) );
  INV_X1 U19577 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19875) );
  AOI22_X1 U19578 ( .A1(n16500), .A2(n18822), .B1(n19875), .B2(n16501), .ZN(
        U361) );
  INV_X1 U19579 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18819) );
  INV_X1 U19580 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19873) );
  AOI22_X1 U19581 ( .A1(n16500), .A2(n18819), .B1(n19873), .B2(n16501), .ZN(
        U362) );
  INV_X1 U19582 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18818) );
  INV_X1 U19583 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19871) );
  AOI22_X1 U19584 ( .A1(n16500), .A2(n18818), .B1(n19871), .B2(n16501), .ZN(
        U363) );
  INV_X1 U19585 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18816) );
  INV_X1 U19586 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19870) );
  AOI22_X1 U19587 ( .A1(n16500), .A2(n18816), .B1(n19870), .B2(n16501), .ZN(
        U364) );
  INV_X1 U19588 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18778) );
  INV_X1 U19589 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19842) );
  AOI22_X1 U19590 ( .A1(n16500), .A2(n18778), .B1(n19842), .B2(n16501), .ZN(
        U365) );
  INV_X1 U19591 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18813) );
  INV_X1 U19592 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19868) );
  AOI22_X1 U19593 ( .A1(n16500), .A2(n18813), .B1(n19868), .B2(n16501), .ZN(
        U366) );
  INV_X1 U19594 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18812) );
  INV_X1 U19595 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19866) );
  AOI22_X1 U19596 ( .A1(n16500), .A2(n18812), .B1(n19866), .B2(n16501), .ZN(
        U367) );
  INV_X1 U19597 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18810) );
  INV_X1 U19598 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19864) );
  AOI22_X1 U19599 ( .A1(n16500), .A2(n18810), .B1(n19864), .B2(n16501), .ZN(
        U368) );
  INV_X1 U19600 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18808) );
  INV_X1 U19601 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19863) );
  AOI22_X1 U19602 ( .A1(n16500), .A2(n18808), .B1(n19863), .B2(n16501), .ZN(
        U369) );
  INV_X1 U19603 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18806) );
  INV_X1 U19604 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19861) );
  AOI22_X1 U19605 ( .A1(n16500), .A2(n18806), .B1(n19861), .B2(n16501), .ZN(
        U370) );
  INV_X1 U19606 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18804) );
  INV_X1 U19607 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19860) );
  AOI22_X1 U19608 ( .A1(n16500), .A2(n18804), .B1(n19860), .B2(n16501), .ZN(
        U371) );
  INV_X1 U19609 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18801) );
  INV_X1 U19610 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19859) );
  AOI22_X1 U19611 ( .A1(n16500), .A2(n18801), .B1(n19859), .B2(n16501), .ZN(
        U372) );
  INV_X1 U19612 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18800) );
  INV_X1 U19613 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19858) );
  AOI22_X1 U19614 ( .A1(n16500), .A2(n18800), .B1(n19858), .B2(n16501), .ZN(
        U373) );
  INV_X1 U19615 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18798) );
  INV_X1 U19616 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19857) );
  AOI22_X1 U19617 ( .A1(n16500), .A2(n18798), .B1(n19857), .B2(n16501), .ZN(
        U374) );
  INV_X1 U19618 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18796) );
  INV_X1 U19619 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19855) );
  AOI22_X1 U19620 ( .A1(n16500), .A2(n18796), .B1(n19855), .B2(n16501), .ZN(
        U375) );
  INV_X1 U19621 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18775) );
  INV_X1 U19622 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19840) );
  AOI22_X1 U19623 ( .A1(n16500), .A2(n18775), .B1(n19840), .B2(n16501), .ZN(
        U376) );
  INV_X1 U19624 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16503) );
  INV_X1 U19625 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18774) );
  NAND2_X1 U19626 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18774), .ZN(n16502) );
  AOI22_X1 U19627 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n16502), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18771), .ZN(n18851) );
  OAI21_X1 U19628 ( .B1(n18771), .B2(n16503), .A(n9631), .ZN(P3_U2633) );
  OAI21_X1 U19629 ( .B1(n16510), .B2(n17479), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16504) );
  OAI21_X1 U19630 ( .B1(n16505), .B2(n18752), .A(n16504), .ZN(P3_U2634) );
  AOI21_X1 U19631 ( .B1(n18771), .B2(n18774), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16506) );
  AOI22_X1 U19632 ( .A1(n18830), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16506), 
        .B2(n18896), .ZN(P3_U2635) );
  INV_X1 U19633 ( .A(BS16), .ZN(n21030) );
  AOI21_X1 U19634 ( .B1(n16507), .B2(n21030), .A(n9631), .ZN(n18847) );
  INV_X1 U19635 ( .A(n18847), .ZN(n18849) );
  OAI21_X1 U19636 ( .B1(n18851), .B2(n18905), .A(n18849), .ZN(P3_U2636) );
  INV_X1 U19637 ( .A(n18725), .ZN(n16509) );
  NOR3_X1 U19638 ( .A1(n16510), .A2(n16509), .A3(n16508), .ZN(n18731) );
  NOR2_X1 U19639 ( .A1(n18731), .A2(n18747), .ZN(n18898) );
  OAI21_X1 U19640 ( .B1(n18898), .B2(n18224), .A(n16511), .ZN(P3_U2637) );
  NOR4_X1 U19641 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16515) );
  NOR4_X1 U19642 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16514) );
  NOR4_X1 U19643 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16513) );
  NOR4_X1 U19644 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16512) );
  NAND4_X1 U19645 ( .A1(n16515), .A2(n16514), .A3(n16513), .A4(n16512), .ZN(
        n16521) );
  NOR4_X1 U19646 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16519) );
  AOI211_X1 U19647 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16518) );
  NOR4_X1 U19648 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16517) );
  NOR4_X1 U19649 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16516) );
  NAND4_X1 U19650 ( .A1(n16519), .A2(n16518), .A3(n16517), .A4(n16516), .ZN(
        n16520) );
  NOR2_X1 U19651 ( .A1(n16521), .A2(n16520), .ZN(n18895) );
  INV_X1 U19652 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18845) );
  NOR3_X1 U19653 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16523) );
  OAI21_X1 U19654 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16523), .A(n18895), .ZN(
        n16522) );
  OAI21_X1 U19655 ( .B1(n18895), .B2(n18845), .A(n16522), .ZN(P3_U2638) );
  INV_X1 U19656 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18776) );
  INV_X1 U19657 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18850) );
  AOI21_X1 U19658 ( .B1(n18776), .B2(n18850), .A(n16523), .ZN(n16524) );
  INV_X1 U19659 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18842) );
  INV_X1 U19660 ( .A(n18895), .ZN(n18892) );
  AOI22_X1 U19661 ( .A1(n18895), .A2(n16524), .B1(n18842), .B2(n18892), .ZN(
        P3_U2639) );
  NAND2_X1 U19662 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n16530), .ZN(n16527) );
  AOI211_X4 U19663 ( .C1(n18905), .C2(n18907), .A(n18919), .B(n16527), .ZN(
        n16905) );
  NOR3_X1 U19664 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16872) );
  NAND2_X1 U19665 ( .A1(n16872), .A2(n16866), .ZN(n16865) );
  NOR2_X1 U19666 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16865), .ZN(n16849) );
  INV_X1 U19667 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16840) );
  NAND2_X1 U19668 ( .A1(n16849), .A2(n16840), .ZN(n16839) );
  NOR2_X1 U19669 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16839), .ZN(n16823) );
  NAND2_X1 U19670 ( .A1(n16823), .A2(n17231), .ZN(n16820) );
  INV_X1 U19671 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16787) );
  NAND2_X1 U19672 ( .A1(n16794), .A2(n16787), .ZN(n16778) );
  INV_X1 U19673 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16773) );
  NAND2_X1 U19674 ( .A1(n16777), .A2(n16773), .ZN(n16765) );
  NAND2_X1 U19675 ( .A1(n16749), .A2(n16748), .ZN(n16745) );
  INV_X1 U19676 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16718) );
  NAND2_X1 U19677 ( .A1(n16725), .A2(n16718), .ZN(n16715) );
  INV_X1 U19678 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16695) );
  NAND2_X1 U19679 ( .A1(n16704), .A2(n16695), .ZN(n16693) );
  NAND2_X1 U19680 ( .A1(n16681), .A2(n16670), .ZN(n16668) );
  INV_X1 U19681 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16913) );
  NAND2_X1 U19682 ( .A1(n16660), .A2(n16913), .ZN(n16652) );
  NOR2_X1 U19683 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16652), .ZN(n16639) );
  INV_X1 U19684 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16915) );
  NAND2_X1 U19685 ( .A1(n16639), .A2(n16915), .ZN(n16633) );
  NOR2_X1 U19686 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16633), .ZN(n16619) );
  INV_X1 U19687 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16613) );
  NAND2_X1 U19688 ( .A1(n16619), .A2(n16613), .ZN(n16612) );
  NOR2_X1 U19689 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16612), .ZN(n16594) );
  NAND2_X1 U19690 ( .A1(n16594), .A2(n16917), .ZN(n16590) );
  NOR2_X1 U19691 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16590), .ZN(n16575) );
  INV_X1 U19692 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16954) );
  NAND2_X1 U19693 ( .A1(n16575), .A2(n16954), .ZN(n16552) );
  NOR2_X1 U19694 ( .A1(n16898), .A2(n16552), .ZN(n16560) );
  INV_X1 U19695 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16924) );
  NAND3_X1 U19696 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(P3_REIP_REG_24__SCAN_IN), .ZN(n16537) );
  OAI211_X1 U19697 ( .C1(n17415), .C2(n16530), .A(n18907), .B(n18905), .ZN(
        n18741) );
  INV_X1 U19698 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18811) );
  INV_X1 U19699 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18809) );
  INV_X1 U19700 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18802) );
  INV_X1 U19701 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18799) );
  INV_X1 U19702 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18795) );
  INV_X1 U19703 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18787) );
  INV_X1 U19704 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18785) );
  INV_X1 U19705 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18779) );
  NAND2_X1 U19706 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16875) );
  NOR2_X1 U19707 ( .A1(n18779), .A2(n16875), .ZN(n16853) );
  NAND3_X1 U19708 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(P3_REIP_REG_4__SCAN_IN), 
        .A3(n16853), .ZN(n16815) );
  NOR3_X1 U19709 ( .A1(n18787), .A2(n18785), .A3(n16815), .ZN(n16800) );
  NAND2_X1 U19710 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16800), .ZN(n16783) );
  NAND2_X1 U19711 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16761) );
  NOR3_X1 U19712 ( .A1(n18795), .A2(n16783), .A3(n16761), .ZN(n16752) );
  NAND2_X1 U19713 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16752), .ZN(n16738) );
  NOR3_X1 U19714 ( .A1(n18802), .A2(n18799), .A3(n16738), .ZN(n16701) );
  NAND4_X1 U19715 ( .A1(n16701), .A2(P3_REIP_REG_17__SCAN_IN), .A3(
        P3_REIP_REG_16__SCAN_IN), .A4(P3_REIP_REG_15__SCAN_IN), .ZN(n16671) );
  NOR3_X1 U19716 ( .A1(n18811), .A2(n18809), .A3(n16671), .ZN(n16657) );
  NAND2_X1 U19717 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16657), .ZN(n16636) );
  NAND3_X1 U19718 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .A3(P3_REIP_REG_21__SCAN_IN), .ZN(n16536) );
  NOR2_X1 U19719 ( .A1(n16636), .A2(n16536), .ZN(n16618) );
  NAND2_X1 U19720 ( .A1(n16874), .A2(n16618), .ZN(n16607) );
  NOR2_X1 U19721 ( .A1(n16537), .A2(n16607), .ZN(n16589) );
  NAND4_X1 U19722 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16589), .ZN(n16535) );
  NOR3_X1 U19723 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18839), .A3(n16535), 
        .ZN(n16534) );
  NAND3_X1 U19724 ( .A1(n16528), .A2(n18749), .A3(n18905), .ZN(n18757) );
  NOR2_X2 U19725 ( .A1(n18865), .A2(n18757), .ZN(n16893) );
  NOR2_X1 U19726 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18854), .ZN(n18750) );
  INV_X1 U19727 ( .A(n18750), .ZN(n18622) );
  OR2_X1 U19728 ( .A1(n18752), .A2(n18622), .ZN(n18745) );
  INV_X1 U19729 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n16531) );
  INV_X1 U19730 ( .A(n18741), .ZN(n16529) );
  AOI211_X4 U19731 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n16530), .A(n16529), .B(
        n18919), .ZN(n16906) );
  OAI22_X1 U19732 ( .A1(n16532), .A2(n16878), .B1(n16531), .B2(n16894), .ZN(
        n16533) );
  AOI211_X1 U19733 ( .C1(n16560), .C2(n16924), .A(n16534), .B(n16533), .ZN(
        n16551) );
  NOR2_X1 U19734 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16535), .ZN(n16558) );
  NAND3_X1 U19735 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16538) );
  INV_X1 U19736 ( .A(n16636), .ZN(n16626) );
  NAND2_X1 U19737 ( .A1(n16626), .A2(n16909), .ZN(n16646) );
  OR2_X1 U19738 ( .A1(n16646), .A2(n16536), .ZN(n16604) );
  NAND2_X1 U19739 ( .A1(n16909), .A2(n16895), .ZN(n16908) );
  OAI21_X1 U19740 ( .B1(n16604), .B2(n16537), .A(n16908), .ZN(n16593) );
  INV_X1 U19741 ( .A(n16593), .ZN(n16600) );
  AOI21_X1 U19742 ( .B1(n16874), .B2(n16538), .A(n16600), .ZN(n16556) );
  INV_X1 U19743 ( .A(n16556), .ZN(n16571) );
  OAI21_X1 U19744 ( .B1(n16558), .B2(n16571), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n16550) );
  INV_X1 U19745 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17555) );
  NOR2_X1 U19746 ( .A1(n17555), .A2(n16541), .ZN(n16540) );
  OAI21_X1 U19747 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16540), .A(
        n16539), .ZN(n17542) );
  INV_X1 U19748 ( .A(n17542), .ZN(n16578) );
  AOI21_X1 U19749 ( .B1(n17555), .B2(n16541), .A(n16540), .ZN(n17551) );
  OAI21_X1 U19750 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17532), .A(
        n16541), .ZN(n17566) );
  INV_X1 U19751 ( .A(n17566), .ZN(n16597) );
  INV_X1 U19752 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16608) );
  NOR2_X1 U19753 ( .A1(n17889), .A2(n17580), .ZN(n16544) );
  NAND2_X1 U19754 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16544), .ZN(
        n16542) );
  AOI21_X1 U19755 ( .B1(n16608), .B2(n16542), .A(n17532), .ZN(n17573) );
  INV_X1 U19756 ( .A(n16544), .ZN(n16543) );
  INV_X1 U19757 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17587) );
  AOI22_X1 U19758 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16544), .B1(
        n16543), .B2(n17587), .ZN(n17585) );
  NAND2_X1 U19759 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9774), .ZN(
        n16545) );
  AOI21_X1 U19760 ( .B1(n9952), .B2(n16545), .A(n16544), .ZN(n17601) );
  INV_X1 U19761 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17620) );
  INV_X1 U19762 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16688) );
  NAND2_X1 U19763 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17672), .ZN(
        n16689) );
  NOR2_X1 U19764 ( .A1(n16688), .A2(n16689), .ZN(n17650) );
  INV_X1 U19765 ( .A(n17650), .ZN(n16677) );
  NOR2_X1 U19766 ( .A1(n17652), .A2(n16677), .ZN(n16548) );
  INV_X1 U19767 ( .A(n16548), .ZN(n17612) );
  NOR2_X1 U19768 ( .A1(n9951), .A2(n17612), .ZN(n16547) );
  NAND2_X1 U19769 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16547), .ZN(
        n16546) );
  AOI22_X1 U19770 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9774), .B1(
        n17620), .B2(n16546), .ZN(n17618) );
  INV_X1 U19771 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17625) );
  XNOR2_X1 U19772 ( .A(n17625), .B(n16547), .ZN(n17634) );
  AOI21_X1 U19773 ( .B1(n9951), .B2(n17612), .A(n16547), .ZN(n17643) );
  INV_X1 U19774 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16890) );
  NOR2_X1 U19775 ( .A1(n17643), .A2(n16659), .ZN(n16658) );
  NOR2_X1 U19776 ( .A1(n16658), .A2(n16858), .ZN(n16649) );
  NOR2_X1 U19777 ( .A1(n17634), .A2(n16649), .ZN(n16648) );
  NOR2_X1 U19778 ( .A1(n16648), .A2(n16858), .ZN(n16638) );
  NOR2_X1 U19779 ( .A1(n17618), .A2(n16638), .ZN(n16637) );
  NOR2_X1 U19780 ( .A1(n16637), .A2(n16858), .ZN(n16628) );
  NOR2_X1 U19781 ( .A1(n17601), .A2(n16628), .ZN(n16627) );
  NOR2_X1 U19782 ( .A1(n16627), .A2(n16858), .ZN(n16621) );
  NOR2_X1 U19783 ( .A1(n17585), .A2(n16621), .ZN(n16620) );
  NOR2_X1 U19784 ( .A1(n16620), .A2(n16858), .ZN(n16606) );
  NOR2_X1 U19785 ( .A1(n17573), .A2(n16606), .ZN(n16605) );
  NOR2_X1 U19786 ( .A1(n16605), .A2(n16858), .ZN(n16596) );
  NOR2_X1 U19787 ( .A1(n16597), .A2(n16596), .ZN(n16595) );
  NOR2_X1 U19788 ( .A1(n16595), .A2(n16858), .ZN(n16586) );
  NOR2_X1 U19789 ( .A1(n17551), .A2(n16586), .ZN(n16585) );
  NOR2_X1 U19790 ( .A1(n16585), .A2(n16858), .ZN(n16577) );
  NOR2_X1 U19791 ( .A1(n16578), .A2(n16577), .ZN(n16576) );
  NOR2_X1 U19792 ( .A1(n16576), .A2(n16858), .ZN(n16567) );
  NOR2_X1 U19793 ( .A1(n16568), .A2(n16567), .ZN(n16566) );
  NAND4_X1 U19794 ( .A1(n16846), .A2(n16893), .A3(n16566), .A4(n16553), .ZN(
        n16549) );
  NAND3_X1 U19795 ( .A1(n16551), .A2(n16550), .A3(n16549), .ZN(P3_U2640) );
  NAND2_X1 U19796 ( .A1(n16905), .A2(n16552), .ZN(n16564) );
  NOR2_X1 U19797 ( .A1(n16566), .A2(n16858), .ZN(n16554) );
  XNOR2_X1 U19798 ( .A(n16554), .B(n16553), .ZN(n16559) );
  OAI22_X1 U19799 ( .A1(n16556), .A2(n18839), .B1(n16555), .B2(n16878), .ZN(
        n16557) );
  AOI211_X1 U19800 ( .C1(n16559), .C2(n16893), .A(n16558), .B(n16557), .ZN(
        n16562) );
  OAI21_X1 U19801 ( .B1(n16906), .B2(n16560), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16561) );
  OAI211_X1 U19802 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16564), .A(n16562), .B(
        n16561), .ZN(P3_U2641) );
  NAND2_X1 U19803 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16581) );
  NOR2_X1 U19804 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16581), .ZN(n16563) );
  AOI22_X1 U19805 ( .A1(n16906), .A2(P3_EBX_REG_29__SCAN_IN), .B1(n16589), 
        .B2(n16563), .ZN(n16573) );
  INV_X1 U19806 ( .A(n16575), .ZN(n16565) );
  AOI21_X1 U19807 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16565), .A(n16564), .ZN(
        n16570) );
  AOI211_X1 U19808 ( .C1(n16568), .C2(n16567), .A(n16566), .B(n18755), .ZN(
        n16569) );
  AOI211_X1 U19809 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n16571), .A(n16570), 
        .B(n16569), .ZN(n16572) );
  OAI211_X1 U19810 ( .C1(n16574), .C2(n16878), .A(n16573), .B(n16572), .ZN(
        P3_U2642) );
  AOI22_X1 U19811 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16891), .B1(
        n16906), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16584) );
  AOI211_X1 U19812 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16590), .A(n16575), .B(
        n16898), .ZN(n16580) );
  AOI211_X1 U19813 ( .C1(n16578), .C2(n16577), .A(n16576), .B(n18755), .ZN(
        n16579) );
  AOI211_X1 U19814 ( .C1(n16600), .C2(P3_REIP_REG_28__SCAN_IN), .A(n16580), 
        .B(n16579), .ZN(n16583) );
  OAI211_X1 U19815 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16589), .B(n16581), .ZN(n16582) );
  NAND3_X1 U19816 ( .A1(n16584), .A2(n16583), .A3(n16582), .ZN(P3_U2643) );
  INV_X1 U19817 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18828) );
  AOI211_X1 U19818 ( .C1(n17551), .C2(n16586), .A(n16585), .B(n18755), .ZN(
        n16588) );
  OAI22_X1 U19819 ( .A1(n17555), .A2(n16878), .B1(n16894), .B2(n16917), .ZN(
        n16587) );
  AOI211_X1 U19820 ( .C1(n16589), .C2(n18828), .A(n16588), .B(n16587), .ZN(
        n16592) );
  OAI211_X1 U19821 ( .C1(n16594), .C2(n16917), .A(n16905), .B(n16590), .ZN(
        n16591) );
  OAI211_X1 U19822 ( .C1(n16593), .C2(n18828), .A(n16592), .B(n16591), .ZN(
        P3_U2644) );
  INV_X1 U19823 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18825) );
  NAND3_X1 U19824 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(P3_REIP_REG_24__SCAN_IN), 
        .A3(n18825), .ZN(n16603) );
  AOI22_X1 U19825 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16891), .B1(
        n16906), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16602) );
  AOI211_X1 U19826 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16612), .A(n16594), .B(
        n16898), .ZN(n16599) );
  AOI211_X1 U19827 ( .C1(n16597), .C2(n16596), .A(n16595), .B(n18755), .ZN(
        n16598) );
  AOI211_X1 U19828 ( .C1(n16600), .C2(P3_REIP_REG_26__SCAN_IN), .A(n16599), 
        .B(n16598), .ZN(n16601) );
  OAI211_X1 U19829 ( .C1(n16607), .C2(n16603), .A(n16602), .B(n16601), .ZN(
        P3_U2645) );
  INV_X1 U19830 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18821) );
  AND2_X1 U19831 ( .A1(n16908), .A2(n16604), .ZN(n16632) );
  AOI21_X1 U19832 ( .B1(n16874), .B2(n18821), .A(n16632), .ZN(n16616) );
  INV_X1 U19833 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18823) );
  AOI211_X1 U19834 ( .C1(n17573), .C2(n16606), .A(n16605), .B(n18755), .ZN(
        n16611) );
  NOR3_X1 U19835 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n18821), .A3(n16607), 
        .ZN(n16610) );
  OAI22_X1 U19836 ( .A1(n16608), .A2(n16878), .B1(n16894), .B2(n16613), .ZN(
        n16609) );
  NOR3_X1 U19837 ( .A1(n16611), .A2(n16610), .A3(n16609), .ZN(n16615) );
  OAI211_X1 U19838 ( .C1(n16619), .C2(n16613), .A(n16905), .B(n16612), .ZN(
        n16614) );
  OAI211_X1 U19839 ( .C1(n16616), .C2(n18823), .A(n16615), .B(n16614), .ZN(
        P3_U2646) );
  NOR2_X1 U19840 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16895), .ZN(n16617) );
  AOI22_X1 U19841 ( .A1(n16906), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16618), 
        .B2(n16617), .ZN(n16625) );
  AOI211_X1 U19842 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16633), .A(n16619), .B(
        n16898), .ZN(n16623) );
  AOI211_X1 U19843 ( .C1(n17585), .C2(n16621), .A(n16620), .B(n18755), .ZN(
        n16622) );
  AOI211_X1 U19844 ( .C1(n16632), .C2(P3_REIP_REG_24__SCAN_IN), .A(n16623), 
        .B(n16622), .ZN(n16624) );
  OAI211_X1 U19845 ( .C1(n17587), .C2(n16878), .A(n16625), .B(n16624), .ZN(
        P3_U2647) );
  INV_X1 U19846 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18817) );
  NAND3_X1 U19847 ( .A1(n16874), .A2(n16626), .A3(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n16645) );
  INV_X1 U19848 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18820) );
  OAI21_X1 U19849 ( .B1(n18817), .B2(n16645), .A(n18820), .ZN(n16631) );
  AOI211_X1 U19850 ( .C1(n17601), .C2(n16628), .A(n16627), .B(n18755), .ZN(
        n16630) );
  OAI22_X1 U19851 ( .A1(n9952), .A2(n16878), .B1(n16894), .B2(n16915), .ZN(
        n16629) );
  AOI211_X1 U19852 ( .C1(n16632), .C2(n16631), .A(n16630), .B(n16629), .ZN(
        n16635) );
  OAI211_X1 U19853 ( .C1(n16639), .C2(n16915), .A(n16905), .B(n16633), .ZN(
        n16634) );
  NAND2_X1 U19854 ( .A1(n16635), .A2(n16634), .ZN(P3_U2648) );
  NOR3_X1 U19855 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16636), .A3(n16895), 
        .ZN(n16650) );
  AOI21_X1 U19856 ( .B1(n16908), .B2(n16646), .A(n16650), .ZN(n16644) );
  AOI211_X1 U19857 ( .C1(n17618), .C2(n16638), .A(n16637), .B(n18755), .ZN(
        n16642) );
  AOI211_X1 U19858 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16652), .A(n16639), .B(
        n16898), .ZN(n16641) );
  OAI22_X1 U19859 ( .A1(n17620), .A2(n16878), .B1(n16894), .B2(n16914), .ZN(
        n16640) );
  NOR3_X1 U19860 ( .A1(n16642), .A2(n16641), .A3(n16640), .ZN(n16643) );
  OAI221_X1 U19861 ( .B1(P3_REIP_REG_22__SCAN_IN), .B2(n16645), .C1(n18817), 
        .C2(n16644), .A(n16643), .ZN(P3_U2649) );
  INV_X1 U19862 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18815) );
  NAND2_X1 U19863 ( .A1(n16908), .A2(n16646), .ZN(n16665) );
  AOI22_X1 U19864 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16891), .B1(
        n16906), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n16655) );
  INV_X1 U19865 ( .A(n16660), .ZN(n16647) );
  AOI21_X1 U19866 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n16647), .A(n16898), .ZN(
        n16653) );
  AOI211_X1 U19867 ( .C1(n17634), .C2(n16649), .A(n16648), .B(n18755), .ZN(
        n16651) );
  AOI211_X1 U19868 ( .C1(n16653), .C2(n16652), .A(n16651), .B(n16650), .ZN(
        n16654) );
  OAI211_X1 U19869 ( .C1(n18815), .C2(n16665), .A(n16655), .B(n16654), .ZN(
        P3_U2650) );
  INV_X1 U19870 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18814) );
  NOR2_X1 U19871 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16895), .ZN(n16656) );
  AOI22_X1 U19872 ( .A1(n16906), .A2(P3_EBX_REG_20__SCAN_IN), .B1(n16657), 
        .B2(n16656), .ZN(n16664) );
  AOI211_X1 U19873 ( .C1(n17643), .C2(n16659), .A(n16658), .B(n18755), .ZN(
        n16662) );
  AOI211_X1 U19874 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16668), .A(n16660), .B(
        n16898), .ZN(n16661) );
  AOI211_X1 U19875 ( .C1(n16891), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16662), .B(n16661), .ZN(n16663) );
  OAI211_X1 U19876 ( .C1(n18814), .C2(n16665), .A(n16664), .B(n16663), .ZN(
        P3_U2651) );
  INV_X1 U19877 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17663) );
  NOR2_X1 U19878 ( .A1(n17663), .A2(n16677), .ZN(n16666) );
  OAI21_X1 U19879 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16666), .A(
        n17612), .ZN(n17655) );
  NOR2_X1 U19880 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16677), .ZN(
        n16678) );
  AOI21_X1 U19881 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n16678), .A(
        n16858), .ZN(n16667) );
  XOR2_X1 U19882 ( .A(n17655), .B(n16667), .Z(n16676) );
  OAI211_X1 U19883 ( .C1(n16681), .C2(n16670), .A(n16905), .B(n16668), .ZN(
        n16669) );
  OAI211_X1 U19884 ( .C1(n16894), .C2(n16670), .A(n18217), .B(n16669), .ZN(
        n16674) );
  NOR4_X1 U19885 ( .A1(n16895), .A2(n18802), .A3(n18799), .A4(n16738), .ZN(
        n16714) );
  NAND4_X1 U19886 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .A4(n16714), .ZN(n16687) );
  XNOR2_X1 U19887 ( .A(n18811), .B(n18809), .ZN(n16672) );
  INV_X1 U19888 ( .A(n16909), .ZN(n16901) );
  AOI21_X1 U19889 ( .B1(n16874), .B2(n16671), .A(n16901), .ZN(n16699) );
  OAI22_X1 U19890 ( .A1(n16687), .A2(n16672), .B1(n18811), .B2(n16699), .ZN(
        n16673) );
  AOI211_X1 U19891 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n16891), .A(
        n16674), .B(n16673), .ZN(n16675) );
  OAI21_X1 U19892 ( .B1(n18755), .B2(n16676), .A(n16675), .ZN(P3_U2652) );
  AOI22_X1 U19893 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16677), .B1(
        n17650), .B2(n17663), .ZN(n17660) );
  OR2_X1 U19894 ( .A1(n16678), .A2(n16858), .ZN(n16680) );
  OAI21_X1 U19895 ( .B1(n17660), .B2(n16680), .A(n16893), .ZN(n16679) );
  AOI21_X1 U19896 ( .B1(n17660), .B2(n16680), .A(n16679), .ZN(n16685) );
  AOI211_X1 U19897 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16693), .A(n16681), .B(
        n16898), .ZN(n16684) );
  INV_X1 U19898 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n16682) );
  OAI22_X1 U19899 ( .A1(n17663), .A2(n16878), .B1(n16894), .B2(n16682), .ZN(
        n16683) );
  NOR4_X1 U19900 ( .A1(n9647), .A2(n16685), .A3(n16684), .A4(n16683), .ZN(
        n16686) );
  OAI221_X1 U19901 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16687), .C1(n18809), 
        .C2(n16699), .A(n16686), .ZN(P3_U2653) );
  NAND3_X1 U19902 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .A3(n16714), .ZN(n16700) );
  INV_X1 U19903 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18807) );
  AOI21_X1 U19904 ( .B1(n16688), .B2(n16689), .A(n17650), .ZN(n17674) );
  INV_X1 U19905 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17704) );
  NOR2_X1 U19906 ( .A1(n17889), .A2(n17728), .ZN(n17727) );
  INV_X1 U19907 ( .A(n17727), .ZN(n16733) );
  NOR2_X1 U19908 ( .A1(n17730), .A2(n16733), .ZN(n16734) );
  NAND2_X1 U19909 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16734), .ZN(
        n16724) );
  NOR2_X1 U19910 ( .A1(n17704), .A2(n16724), .ZN(n16690) );
  INV_X1 U19911 ( .A(n16690), .ZN(n16711) );
  NOR2_X1 U19912 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16711), .ZN(
        n16723) );
  OAI21_X1 U19913 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16690), .A(
        n16689), .ZN(n17692) );
  AOI21_X1 U19914 ( .B1(n16723), .B2(n17692), .A(n16858), .ZN(n16692) );
  OAI21_X1 U19915 ( .B1(n17674), .B2(n16692), .A(n16893), .ZN(n16691) );
  AOI21_X1 U19916 ( .B1(n17674), .B2(n16692), .A(n16691), .ZN(n16697) );
  OAI211_X1 U19917 ( .C1(n16704), .C2(n16695), .A(n16905), .B(n16693), .ZN(
        n16694) );
  OAI211_X1 U19918 ( .C1(n16894), .C2(n16695), .A(n18217), .B(n16694), .ZN(
        n16696) );
  AOI211_X1 U19919 ( .C1(n16891), .C2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n16697), .B(n16696), .ZN(n16698) );
  OAI221_X1 U19920 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n16700), .C1(n18807), 
        .C2(n16699), .A(n16698), .ZN(P3_U2654) );
  NAND2_X1 U19921 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16714), .ZN(n16710) );
  INV_X1 U19922 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18805) );
  INV_X1 U19923 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18803) );
  NAND2_X1 U19924 ( .A1(n16701), .A2(n16909), .ZN(n16726) );
  OAI21_X1 U19925 ( .B1(n18803), .B2(n16726), .A(n16908), .ZN(n16712) );
  OAI21_X1 U19926 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16711), .A(
        n16846), .ZN(n16703) );
  OAI21_X1 U19927 ( .B1(n17692), .B2(n16703), .A(n16893), .ZN(n16702) );
  AOI21_X1 U19928 ( .B1(n17692), .B2(n16703), .A(n16702), .ZN(n16708) );
  AOI211_X1 U19929 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16715), .A(n16704), .B(
        n16898), .ZN(n16707) );
  INV_X1 U19930 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16705) );
  OAI22_X1 U19931 ( .A1(n16705), .A2(n16878), .B1(n16894), .B2(n17094), .ZN(
        n16706) );
  NOR4_X1 U19932 ( .A1(n9647), .A2(n16708), .A3(n16707), .A4(n16706), .ZN(
        n16709) );
  OAI221_X1 U19933 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(n16710), .C1(n18805), 
        .C2(n16712), .A(n16709), .ZN(P3_U2655) );
  NOR2_X1 U19934 ( .A1(n16858), .A2(n18755), .ZN(n16885) );
  INV_X1 U19935 ( .A(n16724), .ZN(n17687) );
  OAI21_X1 U19936 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17687), .A(
        n16711), .ZN(n17701) );
  NAND2_X1 U19937 ( .A1(n16885), .A2(n17701), .ZN(n16722) );
  OAI21_X1 U19938 ( .B1(n16858), .B2(n16890), .A(n16893), .ZN(n16904) );
  AOI211_X1 U19939 ( .C1(n16846), .C2(n16724), .A(n17701), .B(n16904), .ZN(
        n16720) );
  INV_X1 U19940 ( .A(n16712), .ZN(n16713) );
  OAI21_X1 U19941 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16714), .A(n16713), 
        .ZN(n16717) );
  OAI211_X1 U19942 ( .C1(n16725), .C2(n16718), .A(n16905), .B(n16715), .ZN(
        n16716) );
  OAI211_X1 U19943 ( .C1(n16718), .C2(n16894), .A(n16717), .B(n16716), .ZN(
        n16719) );
  AOI211_X1 U19944 ( .C1(n16891), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16720), .B(n16719), .ZN(n16721) );
  OAI211_X1 U19945 ( .C1(n16723), .C2(n16722), .A(n16721), .B(n18217), .ZN(
        P3_U2656) );
  OAI21_X1 U19946 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16734), .A(
        n16724), .ZN(n17712) );
  NOR2_X1 U19947 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17889), .ZN(
        n16886) );
  INV_X1 U19948 ( .A(n16886), .ZN(n16845) );
  OR2_X1 U19949 ( .A1(n17728), .A2(n16845), .ZN(n16754) );
  OAI21_X1 U19950 ( .B1(n17730), .B2(n16754), .A(n16846), .ZN(n16737) );
  XNOR2_X1 U19951 ( .A(n17712), .B(n16737), .ZN(n16732) );
  AOI211_X1 U19952 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16745), .A(n16725), .B(
        n16898), .ZN(n16730) );
  INV_X1 U19953 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17113) );
  NOR3_X1 U19954 ( .A1(n16895), .A2(n18799), .A3(n16738), .ZN(n16727) );
  OAI211_X1 U19955 ( .C1(P3_REIP_REG_14__SCAN_IN), .C2(n16727), .A(n16908), 
        .B(n16726), .ZN(n16728) );
  OAI211_X1 U19956 ( .C1(n16894), .C2(n17113), .A(n18217), .B(n16728), .ZN(
        n16729) );
  AOI211_X1 U19957 ( .C1(n16891), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16730), .B(n16729), .ZN(n16731) );
  OAI21_X1 U19958 ( .B1(n18755), .B2(n16732), .A(n16731), .ZN(P3_U2657) );
  INV_X1 U19959 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17749) );
  NOR2_X1 U19960 ( .A1(n17749), .A2(n16733), .ZN(n16736) );
  INV_X1 U19961 ( .A(n16736), .ZN(n16753) );
  INV_X1 U19962 ( .A(n16734), .ZN(n16735) );
  OAI21_X1 U19963 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16736), .A(
        n16735), .ZN(n17733) );
  AOI211_X1 U19964 ( .C1(n16846), .C2(n16753), .A(n17733), .B(n16904), .ZN(
        n16744) );
  INV_X1 U19965 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18797) );
  OAI21_X1 U19966 ( .B1(n16752), .B2(n16895), .A(n16909), .ZN(n16771) );
  AOI21_X1 U19967 ( .B1(n16874), .B2(n18797), .A(n16771), .ZN(n16742) );
  NOR2_X1 U19968 ( .A1(n18755), .A2(n16737), .ZN(n16740) );
  NOR2_X1 U19969 ( .A1(n16895), .A2(n16738), .ZN(n16739) );
  AOI22_X1 U19970 ( .A1(n16740), .A2(n17733), .B1(n16739), .B2(n18799), .ZN(
        n16741) );
  OAI211_X1 U19971 ( .C1(n16742), .C2(n18799), .A(n16741), .B(n18217), .ZN(
        n16743) );
  AOI211_X1 U19972 ( .C1(n16891), .C2(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16744), .B(n16743), .ZN(n16747) );
  OAI211_X1 U19973 ( .C1(n16749), .C2(n16748), .A(n16905), .B(n16745), .ZN(
        n16746) );
  OAI211_X1 U19974 ( .C1(n16748), .C2(n16894), .A(n16747), .B(n16746), .ZN(
        P3_U2658) );
  AOI211_X1 U19975 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16765), .A(n16749), .B(
        n16898), .ZN(n16750) );
  AOI21_X1 U19976 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n16906), .A(n16750), .ZN(
        n16759) );
  NOR2_X1 U19977 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16895), .ZN(n16751) );
  AOI22_X1 U19978 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16891), .B1(
        n16752), .B2(n16751), .ZN(n16758) );
  OAI21_X1 U19979 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17727), .A(
        n16753), .ZN(n17745) );
  NAND2_X1 U19980 ( .A1(n16846), .A2(n16754), .ZN(n16755) );
  XOR2_X1 U19981 ( .A(n17745), .B(n16755), .Z(n16756) );
  AOI22_X1 U19982 ( .A1(n16893), .A2(n16756), .B1(P3_REIP_REG_12__SCAN_IN), 
        .B2(n16771), .ZN(n16757) );
  NAND4_X1 U19983 ( .A1(n16759), .A2(n16758), .A3(n16757), .A4(n18217), .ZN(
        P3_U2659) );
  NOR2_X1 U19984 ( .A1(n16895), .A2(n16783), .ZN(n16779) );
  INV_X1 U19985 ( .A(n16779), .ZN(n16760) );
  OAI21_X1 U19986 ( .B1(n16761), .B2(n16760), .A(n18795), .ZN(n16770) );
  INV_X1 U19987 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16768) );
  INV_X1 U19988 ( .A(n17794), .ZN(n17795) );
  NOR2_X1 U19989 ( .A1(n17889), .A2(n17795), .ZN(n16774) );
  NAND2_X1 U19990 ( .A1(n17755), .A2(n16774), .ZN(n16762) );
  AOI21_X1 U19991 ( .B1(n16768), .B2(n16762), .A(n17727), .ZN(n17759) );
  INV_X1 U19992 ( .A(n16762), .ZN(n16775) );
  AOI21_X1 U19993 ( .B1(n16775), .B2(n16890), .A(n16858), .ZN(n16764) );
  AOI21_X1 U19994 ( .B1(n17759), .B2(n16764), .A(n18755), .ZN(n16763) );
  OAI21_X1 U19995 ( .B1(n17759), .B2(n16764), .A(n16763), .ZN(n16767) );
  OAI211_X1 U19996 ( .C1(n16777), .C2(n16773), .A(n16905), .B(n16765), .ZN(
        n16766) );
  OAI211_X1 U19997 ( .C1(n16878), .C2(n16768), .A(n16767), .B(n16766), .ZN(
        n16769) );
  AOI21_X1 U19998 ( .B1(n16771), .B2(n16770), .A(n16769), .ZN(n16772) );
  OAI211_X1 U19999 ( .C1(n16894), .C2(n16773), .A(n16772), .B(n18217), .ZN(
        P3_U2660) );
  INV_X1 U20000 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17770) );
  INV_X1 U20001 ( .A(n16774), .ZN(n16824) );
  NOR2_X1 U20002 ( .A1(n17796), .A2(n16824), .ZN(n16803) );
  NAND2_X1 U20003 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16803), .ZN(
        n16788) );
  AOI21_X1 U20004 ( .B1(n17770), .B2(n16788), .A(n16775), .ZN(n17775) );
  NOR3_X1 U20005 ( .A1(n17795), .A2(n17796), .A3(n16845), .ZN(n16789) );
  AOI21_X1 U20006 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16789), .A(
        n16858), .ZN(n16776) );
  INV_X1 U20007 ( .A(n16776), .ZN(n16791) );
  XOR2_X1 U20008 ( .A(n17775), .B(n16791), .Z(n16786) );
  AOI211_X1 U20009 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16778), .A(n16777), .B(
        n16898), .ZN(n16782) );
  INV_X1 U20010 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18793) );
  NAND3_X1 U20011 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16779), .A3(n18793), 
        .ZN(n16780) );
  OAI211_X1 U20012 ( .C1(n17770), .C2(n16878), .A(n18217), .B(n16780), .ZN(
        n16781) );
  AOI211_X1 U20013 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16906), .A(n16782), .B(
        n16781), .ZN(n16785) );
  NOR3_X1 U20014 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16783), .A3(n16895), .ZN(
        n16793) );
  NAND2_X1 U20015 ( .A1(n16874), .A2(n16783), .ZN(n16798) );
  NAND2_X1 U20016 ( .A1(n16909), .A2(n16798), .ZN(n16806) );
  OAI21_X1 U20017 ( .B1(n16793), .B2(n16806), .A(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n16784) );
  OAI211_X1 U20018 ( .C1(n18755), .C2(n16786), .A(n16785), .B(n16784), .ZN(
        P3_U2661) );
  NOR2_X1 U20019 ( .A1(n16794), .A2(n16898), .ZN(n16802) );
  AOI22_X1 U20020 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16891), .B1(
        n16802), .B2(n16787), .ZN(n16797) );
  OAI21_X1 U20021 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16803), .A(
        n16788), .ZN(n17788) );
  NAND2_X1 U20022 ( .A1(n16893), .A2(n16858), .ZN(n16889) );
  OAI21_X1 U20023 ( .B1(n16789), .B2(n17788), .A(n16893), .ZN(n16790) );
  AOI22_X1 U20024 ( .A1(n17788), .A2(n16791), .B1(n16889), .B2(n16790), .ZN(
        n16792) );
  AOI211_X1 U20025 ( .C1(P3_REIP_REG_9__SCAN_IN), .C2(n16806), .A(n16793), .B(
        n16792), .ZN(n16796) );
  OAI221_X1 U20026 ( .B1(n16906), .B2(n16905), .C1(n16906), .C2(n16794), .A(
        P3_EBX_REG_9__SCAN_IN), .ZN(n16795) );
  NAND4_X1 U20027 ( .A1(n16797), .A2(n16796), .A3(n18217), .A4(n16795), .ZN(
        P3_U2662) );
  INV_X1 U20028 ( .A(n16798), .ZN(n16799) );
  AOI22_X1 U20029 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16891), .B1(
        n16800), .B2(n16799), .ZN(n16810) );
  NAND2_X1 U20030 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16820), .ZN(n16801) );
  AOI22_X1 U20031 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16906), .B1(n16802), .B2(
        n16801), .ZN(n16809) );
  INV_X1 U20032 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17812) );
  NOR3_X1 U20033 ( .A1(n17889), .A2(n17795), .A3(n17812), .ZN(n16812) );
  INV_X1 U20034 ( .A(n16803), .ZN(n16804) );
  OAI21_X1 U20035 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16812), .A(
        n16804), .ZN(n17799) );
  INV_X1 U20036 ( .A(n16812), .ZN(n16805) );
  OAI21_X1 U20037 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16805), .A(
        n16846), .ZN(n16814) );
  XOR2_X1 U20038 ( .A(n17799), .B(n16814), .Z(n16807) );
  AOI22_X1 U20039 ( .A1(n16893), .A2(n16807), .B1(P3_REIP_REG_8__SCAN_IN), 
        .B2(n16806), .ZN(n16808) );
  NAND4_X1 U20040 ( .A1(n16810), .A2(n16809), .A3(n16808), .A4(n18217), .ZN(
        P3_U2663) );
  AOI21_X1 U20041 ( .B1(n16874), .B2(n16815), .A(n16901), .ZN(n16836) );
  NOR2_X1 U20042 ( .A1(n16895), .A2(n16815), .ZN(n16811) );
  NAND2_X1 U20043 ( .A1(n16811), .A2(n18785), .ZN(n16828) );
  AOI21_X1 U20044 ( .B1(n16836), .B2(n16828), .A(n18787), .ZN(n16819) );
  AOI21_X1 U20045 ( .B1(n17794), .B2(n16886), .A(n16858), .ZN(n16826) );
  AOI21_X1 U20046 ( .B1(n17812), .B2(n16824), .A(n16812), .ZN(n17818) );
  INV_X1 U20047 ( .A(n17818), .ZN(n16813) );
  AOI221_X1 U20048 ( .B1(n16826), .B2(n17818), .C1(n16814), .C2(n16813), .A(
        n18755), .ZN(n16818) );
  NOR4_X1 U20049 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n16895), .A3(n18785), .A4(
        n16815), .ZN(n16817) );
  OAI21_X1 U20050 ( .B1(n16894), .B2(n17231), .A(n18217), .ZN(n16816) );
  NOR4_X1 U20051 ( .A1(n16819), .A2(n16818), .A3(n16817), .A4(n16816), .ZN(
        n16822) );
  OAI211_X1 U20052 ( .C1(n16823), .C2(n17231), .A(n16905), .B(n16820), .ZN(
        n16821) );
  OAI211_X1 U20053 ( .C1(n16878), .C2(n17812), .A(n16822), .B(n16821), .ZN(
        P3_U2664) );
  AOI211_X1 U20054 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16839), .A(n16823), .B(
        n16898), .ZN(n16831) );
  NOR2_X1 U20055 ( .A1(n17889), .A2(n17821), .ZN(n16833) );
  OAI21_X1 U20056 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16833), .A(
        n16824), .ZN(n17833) );
  AOI211_X1 U20057 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n16846), .A(
        n17833), .B(n16904), .ZN(n16825) );
  AOI21_X1 U20058 ( .B1(n16891), .B2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16825), .ZN(n16829) );
  NAND3_X1 U20059 ( .A1(n16893), .A2(n16826), .A3(n17833), .ZN(n16827) );
  NAND4_X1 U20060 ( .A1(n16829), .A2(n18217), .A3(n16828), .A4(n16827), .ZN(
        n16830) );
  AOI211_X1 U20061 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16906), .A(n16831), .B(
        n16830), .ZN(n16832) );
  OAI21_X1 U20062 ( .B1(n18785), .B2(n16836), .A(n16832), .ZN(P3_U2665) );
  NOR3_X1 U20063 ( .A1(n16895), .A2(n18779), .A3(n16875), .ZN(n16854) );
  AOI21_X1 U20064 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n16854), .A(
        P3_REIP_REG_5__SCAN_IN), .ZN(n16837) );
  NOR2_X1 U20065 ( .A1(n17889), .A2(n17843), .ZN(n16834) );
  INV_X1 U20066 ( .A(n16834), .ZN(n16843) );
  AOI21_X1 U20067 ( .B1(n17842), .B2(n16843), .A(n16833), .ZN(n17844) );
  AOI21_X1 U20068 ( .B1(n16890), .B2(n16834), .A(n16858), .ZN(n16848) );
  XNOR2_X1 U20069 ( .A(n17844), .B(n16848), .ZN(n16835) );
  OAI22_X1 U20070 ( .A1(n16837), .A2(n16836), .B1(n18755), .B2(n16835), .ZN(
        n16838) );
  AOI211_X1 U20071 ( .C1(n16906), .C2(P3_EBX_REG_5__SCAN_IN), .A(n9647), .B(
        n16838), .ZN(n16842) );
  OAI211_X1 U20072 ( .C1(n16849), .C2(n16840), .A(n16905), .B(n16839), .ZN(
        n16841) );
  OAI211_X1 U20073 ( .C1(n16878), .C2(n17842), .A(n16842), .B(n16841), .ZN(
        P3_U2666) );
  NOR2_X1 U20074 ( .A1(n17889), .A2(n17858), .ZN(n16859) );
  OAI21_X1 U20075 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16859), .A(
        n16843), .ZN(n17861) );
  INV_X1 U20076 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17860) );
  NAND2_X1 U20077 ( .A1(n16844), .A2(n17860), .ZN(n17856) );
  OAI22_X1 U20078 ( .A1(n16846), .A2(n17861), .B1(n16845), .B2(n17856), .ZN(
        n16847) );
  AOI21_X1 U20079 ( .B1(n16848), .B2(n17861), .A(n16847), .ZN(n16857) );
  AOI211_X1 U20080 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16865), .A(n16849), .B(
        n16898), .ZN(n16852) );
  NOR2_X1 U20081 ( .A1(n17418), .A2(n18916), .ZN(n16907) );
  OAI21_X1 U20082 ( .B1(n9663), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16907), .ZN(n16850) );
  OAI211_X1 U20083 ( .C1(n17860), .C2(n16878), .A(n18217), .B(n16850), .ZN(
        n16851) );
  AOI211_X1 U20084 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16906), .A(n16852), .B(
        n16851), .ZN(n16856) );
  OAI21_X1 U20085 ( .B1(n16853), .B2(n16895), .A(n16909), .ZN(n16863) );
  INV_X1 U20086 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18781) );
  AOI22_X1 U20087 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16863), .B1(n16854), 
        .B2(n18781), .ZN(n16855) );
  OAI211_X1 U20088 ( .C1(n16857), .C2(n18755), .A(n16856), .B(n16855), .ZN(
        P3_U2667) );
  AOI22_X1 U20089 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n16891), .B1(
        n16906), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n16870) );
  INV_X1 U20090 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17884) );
  NOR2_X1 U20091 ( .A1(n17889), .A2(n17884), .ZN(n16883) );
  AOI21_X1 U20092 ( .B1(n16883), .B2(n16890), .A(n16858), .ZN(n16861) );
  INV_X1 U20093 ( .A(n16859), .ZN(n16860) );
  OAI21_X1 U20094 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n16883), .A(
        n16860), .ZN(n17872) );
  XNOR2_X1 U20095 ( .A(n16861), .B(n17872), .ZN(n16864) );
  OAI21_X1 U20096 ( .B1(n16895), .B2(n16875), .A(n18779), .ZN(n16862) );
  AOI22_X1 U20097 ( .A1(n16893), .A2(n16864), .B1(n16863), .B2(n16862), .ZN(
        n16869) );
  OAI211_X1 U20098 ( .C1(n16872), .C2(n16866), .A(n16905), .B(n16865), .ZN(
        n16868) );
  AOI21_X1 U20099 ( .B1(n18860), .B2(n18686), .A(n9663), .ZN(n18857) );
  NAND2_X1 U20100 ( .A1(n16907), .A2(n18857), .ZN(n16867) );
  NAND4_X1 U20101 ( .A1(n16870), .A2(n16869), .A3(n16868), .A4(n16867), .ZN(
        P3_U2668) );
  AOI21_X1 U20102 ( .B1(n17889), .B2(n17884), .A(n16883), .ZN(n16871) );
  INV_X1 U20103 ( .A(n16871), .ZN(n17881) );
  INV_X1 U20104 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17259) );
  INV_X1 U20105 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17253) );
  NAND2_X1 U20106 ( .A1(n17259), .A2(n17253), .ZN(n16873) );
  AOI211_X1 U20107 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16873), .A(n16872), .B(
        n16898), .ZN(n16882) );
  OAI211_X1 U20108 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16875), .B(n16874), .ZN(n16876) );
  INV_X1 U20109 ( .A(n16876), .ZN(n16881) );
  INV_X1 U20110 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n16877) );
  OAI22_X1 U20111 ( .A1(n17884), .A2(n16878), .B1(n16894), .B2(n16877), .ZN(
        n16880) );
  INV_X1 U20112 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18777) );
  NAND2_X1 U20113 ( .A1(n18872), .A2(n18690), .ZN(n18684) );
  NAND2_X1 U20114 ( .A1(n18686), .A2(n18684), .ZN(n18866) );
  INV_X1 U20115 ( .A(n16907), .ZN(n16897) );
  OAI22_X1 U20116 ( .A1(n16909), .A2(n18777), .B1(n18866), .B2(n16897), .ZN(
        n16879) );
  NOR4_X1 U20117 ( .A1(n16882), .A2(n16881), .A3(n16880), .A4(n16879), .ZN(
        n16888) );
  NAND2_X1 U20118 ( .A1(n16883), .A2(n16890), .ZN(n16884) );
  OAI211_X1 U20119 ( .C1(n16886), .C2(n17881), .A(n16885), .B(n16884), .ZN(
        n16887) );
  OAI211_X1 U20120 ( .C1(n16889), .C2(n17881), .A(n16888), .B(n16887), .ZN(
        P3_U2669) );
  NOR2_X1 U20121 ( .A1(n16858), .A2(n16890), .ZN(n16892) );
  AOI21_X1 U20122 ( .B1(n16893), .B2(n16892), .A(n16891), .ZN(n16903) );
  OAI22_X1 U20123 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16895), .B1(n16894), 
        .B2(n17253), .ZN(n16900) );
  NAND2_X1 U20124 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17246) );
  OAI21_X1 U20125 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17246), .ZN(n17254) );
  NAND2_X1 U20126 ( .A1(n16896), .A2(n18690), .ZN(n18873) );
  OAI22_X1 U20127 ( .A1(n16898), .A2(n17254), .B1(n18873), .B2(n16897), .ZN(
        n16899) );
  AOI211_X1 U20128 ( .C1(n16901), .C2(P3_REIP_REG_1__SCAN_IN), .A(n16900), .B(
        n16899), .ZN(n16902) );
  OAI221_X1 U20129 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16904), .C1(
        n17889), .C2(n16903), .A(n16902), .ZN(P3_U2670) );
  NOR2_X1 U20130 ( .A1(n16906), .A2(n16905), .ZN(n16912) );
  AOI22_X1 U20131 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n16908), .B1(n16907), 
        .B2(n18887), .ZN(n16911) );
  NAND3_X1 U20132 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18868), .A3(
        n16909), .ZN(n16910) );
  OAI211_X1 U20133 ( .C1(n16912), .C2(n17259), .A(n16911), .B(n16910), .ZN(
        P3_U2671) );
  NOR4_X1 U20134 ( .A1(n16916), .A2(n16915), .A3(n16914), .A4(n16913), .ZN(
        n16920) );
  NOR4_X1 U20135 ( .A1(n16954), .A2(n16918), .A3(n16917), .A4(n17027), .ZN(
        n16919) );
  NAND4_X1 U20136 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n16920), .A4(n16919), .ZN(n16923) );
  NOR2_X1 U20137 ( .A1(n16924), .A2(n16923), .ZN(n16950) );
  NAND2_X1 U20138 ( .A1(n17251), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16922) );
  NAND2_X1 U20139 ( .A1(n16950), .A2(n18266), .ZN(n16921) );
  OAI22_X1 U20140 ( .A1(n16950), .A2(n16922), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16921), .ZN(P3_U2672) );
  NAND2_X1 U20141 ( .A1(n16924), .A2(n16923), .ZN(n16925) );
  NAND2_X1 U20142 ( .A1(n16925), .A2(n17251), .ZN(n16949) );
  AOI22_X1 U20143 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17210), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16926) );
  OAI21_X1 U20144 ( .B1(n9713), .B2(n17105), .A(n16926), .ZN(n16937) );
  AOI22_X1 U20145 ( .A1(n11217), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16934) );
  INV_X1 U20146 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16927) );
  OAI22_X1 U20147 ( .A1(n17155), .A2(n16927), .B1(n11287), .B2(n18580), .ZN(
        n16932) );
  AOI22_X1 U20148 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16930) );
  AOI22_X1 U20149 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16929) );
  AOI22_X1 U20150 ( .A1(n11202), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9663), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16928) );
  NAND3_X1 U20151 ( .A1(n16930), .A2(n16929), .A3(n16928), .ZN(n16931) );
  AOI211_X1 U20152 ( .C1(n17214), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n16932), .B(n16931), .ZN(n16933) );
  OAI211_X1 U20153 ( .C1(n11187), .C2(n16935), .A(n16934), .B(n16933), .ZN(
        n16936) );
  AOI211_X1 U20154 ( .C1(n17212), .C2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n16937), .B(n16936), .ZN(n16948) );
  INV_X1 U20155 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17114) );
  AOI22_X1 U20156 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16947) );
  AOI22_X1 U20157 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16939) );
  AOI22_X1 U20158 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16938) );
  OAI211_X1 U20159 ( .C1(n17053), .C2(n18574), .A(n16939), .B(n16938), .ZN(
        n16945) );
  AOI22_X1 U20160 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17210), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16943) );
  AOI22_X1 U20161 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16942) );
  AOI22_X1 U20162 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16941) );
  NAND2_X1 U20163 ( .A1(n11202), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n16940) );
  NAND4_X1 U20164 ( .A1(n16943), .A2(n16942), .A3(n16941), .A4(n16940), .ZN(
        n16944) );
  AOI211_X1 U20165 ( .C1(n9663), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n16945), .B(n16944), .ZN(n16946) );
  OAI211_X1 U20166 ( .C1(n17116), .C2(n17114), .A(n16947), .B(n16946), .ZN(
        n16952) );
  NAND2_X1 U20167 ( .A1(n16953), .A2(n16952), .ZN(n16951) );
  XNOR2_X1 U20168 ( .A(n16948), .B(n16951), .ZN(n17271) );
  OAI22_X1 U20169 ( .A1(n16950), .A2(n16949), .B1(n17271), .B2(n17251), .ZN(
        P3_U2673) );
  OAI21_X1 U20170 ( .B1(n16953), .B2(n16952), .A(n16951), .ZN(n17275) );
  AOI22_X1 U20171 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16956), .B1(n16955), 
        .B2(n16954), .ZN(n16957) );
  OAI21_X1 U20172 ( .B1(n17275), .B2(n17251), .A(n16957), .ZN(P3_U2674) );
  OAI21_X1 U20173 ( .B1(n16962), .B2(n16959), .A(n16958), .ZN(n17283) );
  NAND3_X1 U20174 ( .A1(n16961), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17251), 
        .ZN(n16960) );
  OAI221_X1 U20175 ( .B1(n16961), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17251), 
        .C2(n17283), .A(n16960), .ZN(P3_U2676) );
  AOI21_X1 U20176 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17251), .A(n16970), .ZN(
        n16965) );
  AOI21_X1 U20177 ( .B1(n16963), .B2(n16967), .A(n16962), .ZN(n17284) );
  INV_X1 U20178 ( .A(n17284), .ZN(n16964) );
  OAI22_X1 U20179 ( .A1(n16966), .A2(n16965), .B1(n16964), .B2(n17251), .ZN(
        P3_U2677) );
  AOI21_X1 U20180 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17251), .A(n16976), .ZN(
        n16969) );
  OAI21_X1 U20181 ( .B1(n16972), .B2(n16968), .A(n16967), .ZN(n17293) );
  OAI22_X1 U20182 ( .A1(n16970), .A2(n16969), .B1(n17293), .B2(n17251), .ZN(
        P3_U2678) );
  INV_X1 U20183 ( .A(n16971), .ZN(n16981) );
  AOI21_X1 U20184 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17251), .A(n16981), .ZN(
        n16975) );
  AOI21_X1 U20185 ( .B1(n16973), .B2(n16977), .A(n16972), .ZN(n17294) );
  INV_X1 U20186 ( .A(n17294), .ZN(n16974) );
  OAI22_X1 U20187 ( .A1(n16976), .A2(n16975), .B1(n17251), .B2(n16974), .ZN(
        P3_U2679) );
  AOI21_X1 U20188 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17251), .A(n16996), .ZN(
        n16980) );
  OAI21_X1 U20189 ( .B1(n16979), .B2(n16978), .A(n16977), .ZN(n17303) );
  OAI22_X1 U20190 ( .A1(n16981), .A2(n16980), .B1(n17251), .B2(n17303), .ZN(
        P3_U2680) );
  INV_X1 U20191 ( .A(n16982), .ZN(n17013) );
  AOI21_X1 U20192 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17251), .A(n17013), .ZN(
        n16995) );
  AOI22_X1 U20193 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16993) );
  AOI22_X1 U20194 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16992) );
  OAI22_X1 U20195 ( .A1(n9713), .A2(n17115), .B1(n16983), .B2(n17123), .ZN(
        n16990) );
  AOI22_X1 U20196 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16988) );
  AOI22_X1 U20197 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16985) );
  AOI22_X1 U20198 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16984) );
  OAI211_X1 U20199 ( .C1(n17191), .C2(n17114), .A(n16985), .B(n16984), .ZN(
        n16986) );
  AOI21_X1 U20200 ( .B1(n9663), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(n16986), .ZN(n16987) );
  OAI211_X1 U20201 ( .C1(n17116), .C2(n17119), .A(n16988), .B(n16987), .ZN(
        n16989) );
  AOI211_X1 U20202 ( .C1(n17150), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n16990), .B(n16989), .ZN(n16991) );
  NAND3_X1 U20203 ( .A1(n16993), .A2(n16992), .A3(n16991), .ZN(n17305) );
  INV_X1 U20204 ( .A(n17305), .ZN(n16994) );
  OAI22_X1 U20205 ( .A1(n16996), .A2(n16995), .B1(n16994), .B2(n17251), .ZN(
        P3_U2681) );
  AOI21_X1 U20206 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17251), .A(n16997), .ZN(
        n17012) );
  AOI22_X1 U20207 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17010) );
  AOI22_X1 U20208 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17009) );
  OAI22_X1 U20209 ( .A1(n9746), .A2(n16999), .B1(n17015), .B2(n16998), .ZN(
        n17007) );
  OAI22_X1 U20210 ( .A1(n17116), .A2(n17236), .B1(n17053), .B2(n17000), .ZN(
        n17001) );
  AOI21_X1 U20211 ( .B1(n11202), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n17001), .ZN(n17005) );
  AOI22_X1 U20212 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17004) );
  AOI22_X1 U20213 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17003) );
  AOI22_X1 U20214 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9663), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17002) );
  NAND4_X1 U20215 ( .A1(n17005), .A2(n17004), .A3(n17003), .A4(n17002), .ZN(
        n17006) );
  AOI211_X1 U20216 ( .C1(n17150), .C2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n17007), .B(n17006), .ZN(n17008) );
  NAND3_X1 U20217 ( .A1(n17010), .A2(n17009), .A3(n17008), .ZN(n17312) );
  INV_X1 U20218 ( .A(n17312), .ZN(n17011) );
  OAI22_X1 U20219 ( .A1(n17013), .A2(n17012), .B1(n17011), .B2(n17251), .ZN(
        P3_U2682) );
  AOI22_X1 U20220 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9663), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17025) );
  AOI22_X1 U20221 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17014) );
  OAI21_X1 U20222 ( .B1(n17015), .B2(n17136), .A(n17014), .ZN(n17023) );
  OAI22_X1 U20223 ( .A1(n9746), .A2(n17016), .B1(n17116), .B2(n17240), .ZN(
        n17017) );
  AOI21_X1 U20224 ( .B1(n17149), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n17017), .ZN(n17021) );
  AOI22_X1 U20225 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17020) );
  AOI22_X1 U20226 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17019) );
  AOI22_X1 U20227 ( .A1(n11202), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17018) );
  NAND4_X1 U20228 ( .A1(n17021), .A2(n17020), .A3(n17019), .A4(n17018), .ZN(
        n17022) );
  AOI211_X1 U20229 ( .C1(n17167), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n17023), .B(n17022), .ZN(n17024) );
  OAI211_X1 U20230 ( .C1(n11187), .C2(n17026), .A(n17025), .B(n17024), .ZN(
        n17317) );
  INV_X1 U20231 ( .A(n17317), .ZN(n17029) );
  OAI21_X1 U20232 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17044), .A(n17027), .ZN(
        n17028) );
  AOI22_X1 U20233 ( .A1(n17257), .A2(n17029), .B1(n17028), .B2(n17251), .ZN(
        P3_U2683) );
  AOI22_X1 U20234 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17030) );
  OAI21_X1 U20235 ( .B1(n17133), .B2(n17031), .A(n17030), .ZN(n17042) );
  AOI22_X1 U20236 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17039) );
  OAI22_X1 U20237 ( .A1(n17116), .A2(n17244), .B1(n17053), .B2(n17032), .ZN(
        n17037) );
  AOI22_X1 U20238 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17035) );
  AOI22_X1 U20239 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17034) );
  AOI22_X1 U20240 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9663), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17033) );
  NAND3_X1 U20241 ( .A1(n17035), .A2(n17034), .A3(n17033), .ZN(n17036) );
  AOI211_X1 U20242 ( .C1(n11202), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n17037), .B(n17036), .ZN(n17038) );
  OAI211_X1 U20243 ( .C1(n17040), .C2(n17154), .A(n17039), .B(n17038), .ZN(
        n17041) );
  AOI211_X1 U20244 ( .C1(n17212), .C2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A(
        n17042), .B(n17041), .ZN(n17325) );
  NAND2_X1 U20245 ( .A1(n17251), .A2(n17043), .ZN(n17062) );
  NAND2_X1 U20246 ( .A1(n18266), .A2(n17044), .ZN(n17045) );
  OAI21_X1 U20247 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17062), .A(n17045), .ZN(
        n17046) );
  AOI21_X1 U20248 ( .B1(n17257), .B2(n17325), .A(n17046), .ZN(P3_U2684) );
  AOI22_X1 U20249 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17047) );
  OAI21_X1 U20250 ( .B1(n17188), .B2(n17048), .A(n17047), .ZN(n17060) );
  AOI22_X1 U20251 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17057) );
  AOI22_X1 U20252 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17050) );
  OAI21_X1 U20253 ( .B1(n17191), .B2(n17170), .A(n17050), .ZN(n17055) );
  AOI22_X1 U20254 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17167), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17052) );
  AOI22_X1 U20255 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17051) );
  OAI211_X1 U20256 ( .C1(n17053), .C2(n17179), .A(n17052), .B(n17051), .ZN(
        n17054) );
  AOI211_X1 U20257 ( .C1(n9663), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n17055), .B(n17054), .ZN(n17056) );
  OAI211_X1 U20258 ( .C1(n9746), .C2(n17058), .A(n17057), .B(n17056), .ZN(
        n17059) );
  AOI211_X1 U20259 ( .C1(n17185), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n17060), .B(n17059), .ZN(n17330) );
  NOR2_X1 U20260 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17061), .ZN(n17063) );
  OAI22_X1 U20261 ( .A1(n17330), .A2(n17251), .B1(n17063), .B2(n17062), .ZN(
        P3_U2685) );
  AOI22_X1 U20262 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17149), .ZN(n17064) );
  OAI21_X1 U20263 ( .B1(n17065), .B2(n17133), .A(n17064), .ZN(n17074) );
  AOI22_X1 U20264 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n11217), .ZN(n17072) );
  INV_X1 U20265 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17190) );
  OAI22_X1 U20266 ( .A1(n17200), .A2(n17053), .B1(n17191), .B2(n17190), .ZN(
        n17070) );
  AOI22_X1 U20267 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17184), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17068) );
  AOI22_X1 U20268 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n9649), .ZN(n17067) );
  AOI22_X1 U20269 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9663), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17066) );
  NAND3_X1 U20270 ( .A1(n17068), .A2(n17067), .A3(n17066), .ZN(n17069) );
  AOI211_X1 U20271 ( .C1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .C2(n17150), .A(
        n17070), .B(n17069), .ZN(n17071) );
  OAI211_X1 U20272 ( .C1(n17252), .C2(n17116), .A(n17072), .B(n17071), .ZN(
        n17073) );
  AOI211_X1 U20273 ( .C1(n17212), .C2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A(
        n17074), .B(n17073), .ZN(n17335) );
  INV_X1 U20274 ( .A(n17255), .ZN(n17256) );
  OAI211_X1 U20275 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n17076), .A(n17256), .B(
        n17075), .ZN(n17078) );
  NAND2_X1 U20276 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17079), .ZN(n17077) );
  OAI211_X1 U20277 ( .C1(n17335), .C2(n17251), .A(n17078), .B(n17077), .ZN(
        P3_U2686) );
  AOI21_X1 U20278 ( .B1(n18266), .B2(n17091), .A(n17079), .ZN(n17109) );
  AOI22_X1 U20279 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17089) );
  AOI22_X1 U20280 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17081) );
  AOI22_X1 U20281 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17080) );
  OAI211_X1 U20282 ( .C1(n17191), .C2(n17209), .A(n17081), .B(n17080), .ZN(
        n17087) );
  AOI22_X1 U20283 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17085) );
  AOI22_X1 U20284 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17084) );
  AOI22_X1 U20285 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9663), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17083) );
  NAND2_X1 U20286 ( .A1(n17213), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n17082) );
  NAND4_X1 U20287 ( .A1(n17085), .A2(n17084), .A3(n17083), .A4(n17082), .ZN(
        n17086) );
  AOI211_X1 U20288 ( .C1(n17049), .C2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n17087), .B(n17086), .ZN(n17088) );
  OAI211_X1 U20289 ( .C1(n17116), .C2(n17090), .A(n17089), .B(n17088), .ZN(
        n17336) );
  NOR2_X1 U20290 ( .A1(n17091), .A2(n17255), .ZN(n17092) );
  AOI22_X1 U20291 ( .A1(n17257), .A2(n17336), .B1(n17092), .B2(n17094), .ZN(
        n17093) );
  OAI21_X1 U20292 ( .B1(n17094), .B2(n17109), .A(n17093), .ZN(P3_U2687) );
  AOI22_X1 U20293 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17095) );
  OAI21_X1 U20294 ( .B1(n17133), .B2(n18580), .A(n17095), .ZN(n17107) );
  AOI22_X1 U20295 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17104) );
  OAI22_X1 U20296 ( .A1(n17116), .A2(n17097), .B1(n17199), .B2(n17096), .ZN(
        n17102) );
  AOI22_X1 U20297 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17100) );
  AOI22_X1 U20298 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17099) );
  AOI22_X1 U20299 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9663), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17098) );
  NAND3_X1 U20300 ( .A1(n17100), .A2(n17099), .A3(n17098), .ZN(n17101) );
  AOI211_X1 U20301 ( .C1(n11207), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n17102), .B(n17101), .ZN(n17103) );
  OAI211_X1 U20302 ( .C1(n17191), .C2(n17105), .A(n17104), .B(n17103), .ZN(
        n17106) );
  AOI211_X1 U20303 ( .C1(n17212), .C2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n17107), .B(n17106), .ZN(n17348) );
  NAND2_X1 U20304 ( .A1(n17260), .A2(n17108), .ZN(n17112) );
  NOR2_X1 U20305 ( .A1(n17113), .A2(n17112), .ZN(n17111) );
  NOR2_X1 U20306 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17111), .ZN(n17110) );
  OAI22_X1 U20307 ( .A1(n17348), .A2(n17251), .B1(n17110), .B2(n17109), .ZN(
        P3_U2688) );
  AOI21_X1 U20308 ( .B1(n17113), .B2(n17112), .A(n17111), .ZN(n17129) );
  AOI22_X1 U20309 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17128) );
  AOI22_X1 U20310 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17167), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17127) );
  OAI22_X1 U20311 ( .A1(n17116), .A2(n17115), .B1(n11186), .B2(n17114), .ZN(
        n17125) );
  AOI22_X1 U20312 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17122) );
  AOI22_X1 U20313 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17118) );
  AOI22_X1 U20314 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17117) );
  OAI211_X1 U20315 ( .C1(n17191), .C2(n17119), .A(n17118), .B(n17117), .ZN(
        n17120) );
  AOI21_X1 U20316 ( .B1(n17049), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n17120), .ZN(n17121) );
  OAI211_X1 U20317 ( .C1(n11187), .C2(n17123), .A(n17122), .B(n17121), .ZN(
        n17124) );
  AOI211_X1 U20318 ( .C1(n17213), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n17125), .B(n17124), .ZN(n17126) );
  NAND3_X1 U20319 ( .A1(n17128), .A2(n17127), .A3(n17126), .ZN(n17351) );
  MUX2_X1 U20320 ( .A(n17129), .B(n17351), .S(n17257), .Z(P3_U2689) );
  NAND2_X1 U20321 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17242), .ZN(n17232) );
  NOR2_X1 U20322 ( .A1(n17345), .A2(n17232), .ZN(n17233) );
  NAND2_X1 U20323 ( .A1(n17131), .A2(n17233), .ZN(n17164) );
  AOI22_X1 U20324 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17132) );
  OAI21_X1 U20325 ( .B1(n17133), .B2(n18565), .A(n17132), .ZN(n17145) );
  AOI22_X1 U20326 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17143) );
  OAI22_X1 U20327 ( .A1(n17116), .A2(n17136), .B1(n17135), .B2(n17134), .ZN(
        n17141) );
  AOI22_X1 U20328 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17167), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17139) );
  AOI22_X1 U20329 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17138) );
  AOI22_X1 U20330 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9663), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17137) );
  NAND3_X1 U20331 ( .A1(n17139), .A2(n17138), .A3(n17137), .ZN(n17140) );
  AOI211_X1 U20332 ( .C1(n17210), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n17141), .B(n17140), .ZN(n17142) );
  OAI211_X1 U20333 ( .C1(n17191), .C2(n17240), .A(n17143), .B(n17142), .ZN(
        n17144) );
  AOI211_X1 U20334 ( .C1(n11207), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n17145), .B(n17144), .ZN(n17360) );
  NAND3_X1 U20335 ( .A1(n17164), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n17251), 
        .ZN(n17146) );
  OAI221_X1 U20336 ( .B1(n17164), .B2(P3_EBX_REG_12__SCAN_IN), .C1(n17251), 
        .C2(n17360), .A(n17146), .ZN(P3_U2691) );
  OAI22_X1 U20337 ( .A1(n17116), .A2(n17148), .B1(n17188), .B2(n17147), .ZN(
        n17163) );
  AOI22_X1 U20338 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17161) );
  AOI22_X1 U20339 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17160) );
  AOI22_X1 U20340 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17151) );
  OAI21_X1 U20341 ( .B1(n17191), .B2(n17244), .A(n17151), .ZN(n17157) );
  AOI22_X1 U20342 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17153) );
  AOI22_X1 U20343 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17152) );
  OAI211_X1 U20344 ( .C1(n17155), .C2(n17154), .A(n17153), .B(n17152), .ZN(
        n17156) );
  AOI211_X1 U20345 ( .C1(n9663), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n17157), .B(n17156), .ZN(n17159) );
  NAND3_X1 U20346 ( .A1(n17161), .A2(n17160), .A3(n17159), .ZN(n17162) );
  AOI211_X1 U20347 ( .C1(n17185), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n17163), .B(n17162), .ZN(n17364) );
  INV_X1 U20348 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17227) );
  NOR2_X1 U20349 ( .A1(n17227), .A2(n17224), .ZN(n17204) );
  NAND2_X1 U20350 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17204), .ZN(n17203) );
  INV_X1 U20351 ( .A(n17203), .ZN(n17180) );
  AND2_X1 U20352 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17180), .ZN(n17182) );
  NOR2_X1 U20353 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17182), .ZN(n17166) );
  NAND2_X1 U20354 ( .A1(n17251), .A2(n17164), .ZN(n17165) );
  OAI22_X1 U20355 ( .A1(n17364), .A2(n17251), .B1(n17166), .B2(n17165), .ZN(
        P3_U2692) );
  AOI22_X1 U20356 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17178) );
  AOI22_X1 U20357 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17169) );
  AOI22_X1 U20358 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17168) );
  OAI211_X1 U20359 ( .C1(n11186), .C2(n17170), .A(n17169), .B(n17168), .ZN(
        n17176) );
  AOI22_X1 U20360 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17174) );
  AOI22_X1 U20361 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17173) );
  AOI22_X1 U20362 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17172) );
  NAND2_X1 U20363 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n17171) );
  NAND4_X1 U20364 ( .A1(n17174), .A2(n17173), .A3(n17172), .A4(n17171), .ZN(
        n17175) );
  AOI211_X1 U20365 ( .C1(n11202), .C2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n17176), .B(n17175), .ZN(n17177) );
  OAI211_X1 U20366 ( .C1(n17199), .C2(n17179), .A(n17178), .B(n17177), .ZN(
        n17367) );
  INV_X1 U20367 ( .A(n17367), .ZN(n17183) );
  OAI21_X1 U20368 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17180), .A(n17251), .ZN(
        n17181) );
  OAI22_X1 U20369 ( .A1(n17183), .A2(n17251), .B1(n17182), .B2(n17181), .ZN(
        P3_U2693) );
  AOI22_X1 U20370 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17186) );
  OAI21_X1 U20371 ( .B1(n17188), .B2(n17187), .A(n17186), .ZN(n17202) );
  AOI22_X1 U20372 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17189), .ZN(n17198) );
  OAI22_X1 U20373 ( .A1(n17252), .A2(n17191), .B1(n17190), .B2(n11186), .ZN(
        n17196) );
  AOI22_X1 U20374 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n11217), .ZN(n17194) );
  AOI22_X1 U20375 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n9649), .ZN(n17193) );
  AOI22_X1 U20376 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17049), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17192) );
  NAND3_X1 U20377 ( .A1(n17194), .A2(n17193), .A3(n17192), .ZN(n17195) );
  AOI211_X1 U20378 ( .C1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .C2(n17150), .A(
        n17196), .B(n17195), .ZN(n17197) );
  OAI211_X1 U20379 ( .C1(n17200), .C2(n17199), .A(n17198), .B(n17197), .ZN(
        n17201) );
  AOI211_X1 U20380 ( .C1(n17167), .C2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n17202), .B(n17201), .ZN(n17372) );
  OAI21_X1 U20381 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17204), .A(n17203), .ZN(
        n17205) );
  AOI22_X1 U20382 ( .A1(n17257), .A2(n17372), .B1(n17205), .B2(n17251), .ZN(
        P3_U2694) );
  NAND2_X1 U20383 ( .A1(n17251), .A2(n17224), .ZN(n17230) );
  INV_X1 U20384 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18478) );
  AOI22_X1 U20385 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17222) );
  AOI22_X1 U20386 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17208) );
  AOI22_X1 U20387 ( .A1(n9644), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17207) );
  OAI211_X1 U20388 ( .C1(n11186), .C2(n17209), .A(n17208), .B(n17207), .ZN(
        n17220) );
  AOI22_X1 U20389 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17210), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17218) );
  AOI22_X1 U20390 ( .A1(n17212), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11217), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17217) );
  AOI22_X1 U20391 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17213), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17216) );
  NAND2_X1 U20392 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n17215) );
  NAND4_X1 U20393 ( .A1(n17218), .A2(n17217), .A3(n17216), .A4(n17215), .ZN(
        n17219) );
  AOI211_X1 U20394 ( .C1(n11202), .C2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A(
        n17220), .B(n17219), .ZN(n17221) );
  OAI211_X1 U20395 ( .C1(n17223), .C2(n18478), .A(n17222), .B(n17221), .ZN(
        n17379) );
  NOR3_X1 U20396 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17345), .A3(n17224), .ZN(
        n17225) );
  AOI21_X1 U20397 ( .B1(n17257), .B2(n17379), .A(n17225), .ZN(n17226) );
  OAI21_X1 U20398 ( .B1(n17227), .B2(n17230), .A(n17226), .ZN(P3_U2695) );
  NOR2_X1 U20399 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17235), .ZN(n17228) );
  AOI22_X1 U20400 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17257), .B1(
        n17233), .B2(n17228), .ZN(n17229) );
  OAI21_X1 U20401 ( .B1(n17231), .B2(n17230), .A(n17229), .ZN(P3_U2696) );
  NAND2_X1 U20402 ( .A1(n17251), .A2(n17232), .ZN(n17237) );
  AOI22_X1 U20403 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17257), .B1(
        n17233), .B2(n17235), .ZN(n17234) );
  OAI21_X1 U20404 ( .B1(n17235), .B2(n17237), .A(n17234), .ZN(P3_U2697) );
  NOR2_X1 U20405 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17242), .ZN(n17238) );
  OAI22_X1 U20406 ( .A1(n17238), .A2(n17237), .B1(n17236), .B2(n17251), .ZN(
        P3_U2698) );
  NOR2_X1 U20407 ( .A1(n17239), .A2(n17255), .ZN(n17248) );
  AOI22_X1 U20408 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17251), .B1(
        P3_EBX_REG_3__SCAN_IN), .B2(n17248), .ZN(n17241) );
  OAI22_X1 U20409 ( .A1(n17242), .A2(n17241), .B1(n17240), .B2(n17251), .ZN(
        P3_U2699) );
  INV_X1 U20410 ( .A(n17248), .ZN(n17245) );
  NAND3_X1 U20411 ( .A1(n17245), .A2(P3_EBX_REG_3__SCAN_IN), .A3(n17251), .ZN(
        n17243) );
  OAI221_X1 U20412 ( .B1(n17245), .B2(P3_EBX_REG_3__SCAN_IN), .C1(n17251), 
        .C2(n17244), .A(n17243), .ZN(P3_U2700) );
  INV_X1 U20413 ( .A(n17246), .ZN(n17247) );
  AOI221_X1 U20414 ( .B1(n17247), .B2(n17260), .C1(n17345), .C2(n17260), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17249) );
  AOI211_X1 U20415 ( .C1(n17257), .C2(n17250), .A(n17249), .B(n17248), .ZN(
        P3_U2701) );
  OAI222_X1 U20416 ( .A1(n17255), .A2(n17254), .B1(n17253), .B2(n17260), .C1(
        n17252), .C2(n17251), .ZN(P3_U2702) );
  AOI22_X1 U20417 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17257), .B1(
        n17256), .B2(n17259), .ZN(n17258) );
  OAI21_X1 U20418 ( .B1(n17260), .B2(n17259), .A(n17258), .ZN(P3_U2703) );
  INV_X1 U20419 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17422) );
  INV_X1 U20420 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17426) );
  INV_X1 U20421 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17432) );
  INV_X1 U20422 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17531) );
  INV_X1 U20423 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17459) );
  NAND2_X1 U20424 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n17401) );
  INV_X1 U20425 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17464) );
  INV_X1 U20426 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17466) );
  NAND4_X1 U20427 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17261) );
  NOR4_X1 U20428 ( .A1(n17401), .A2(n17464), .A3(n17466), .A4(n17261), .ZN(
        n17384) );
  INV_X1 U20429 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17453) );
  NAND4_X1 U20430 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(P3_EAX_REG_13__SCAN_IN), .A4(P3_EAX_REG_12__SCAN_IN), .ZN(n17263)
         );
  NOR2_X1 U20431 ( .A1(n17453), .A2(n17263), .ZN(n17349) );
  INV_X1 U20432 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17440) );
  INV_X1 U20433 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17482) );
  NOR2_X1 U20434 ( .A1(n17440), .A2(n17482), .ZN(n17306) );
  NAND4_X1 U20435 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_19__SCAN_IN), .A4(n17306), .ZN(n17311) );
  NAND2_X1 U20436 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17300), .ZN(n17299) );
  NAND2_X1 U20437 ( .A1(n17268), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17267) );
  OAI22_X1 U20438 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17400), .B1(n17376), 
        .B2(n17268), .ZN(n17264) );
  AOI22_X1 U20439 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17337), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17264), .ZN(n17265) );
  OAI21_X1 U20440 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17267), .A(n17265), .ZN(
        P3_U2704) );
  NOR2_X2 U20441 ( .A1(n17266), .A2(n17407), .ZN(n17331) );
  AOI22_X1 U20442 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17331), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17337), .ZN(n17270) );
  OAI211_X1 U20443 ( .C1(n17268), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17407), .B(
        n17267), .ZN(n17269) );
  OAI211_X1 U20444 ( .C1(n17271), .C2(n17402), .A(n17270), .B(n17269), .ZN(
        P3_U2705) );
  AOI22_X1 U20445 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17331), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17337), .ZN(n17274) );
  OAI211_X1 U20446 ( .C1(n9719), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17407), .B(
        n17272), .ZN(n17273) );
  OAI211_X1 U20447 ( .C1(n17275), .C2(n17402), .A(n17274), .B(n17273), .ZN(
        P3_U2706) );
  INV_X1 U20448 ( .A(n17337), .ZN(n17289) );
  AOI22_X1 U20449 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17331), .B1(n17410), .B2(
        n17276), .ZN(n17279) );
  AOI211_X1 U20450 ( .C1(n17422), .C2(n17280), .A(n9719), .B(n17376), .ZN(
        n17277) );
  INV_X1 U20451 ( .A(n17277), .ZN(n17278) );
  OAI211_X1 U20452 ( .C1(n17289), .C2(n18248), .A(n17279), .B(n17278), .ZN(
        P3_U2707) );
  AOI22_X1 U20453 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17331), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17337), .ZN(n17282) );
  OAI211_X1 U20454 ( .C1(n17285), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17407), .B(
        n17280), .ZN(n17281) );
  OAI211_X1 U20455 ( .C1(n17283), .C2(n17402), .A(n17282), .B(n17281), .ZN(
        P3_U2708) );
  AOI22_X1 U20456 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17331), .B1(n17410), .B2(
        n17284), .ZN(n17288) );
  AOI211_X1 U20457 ( .C1(n17426), .C2(n9712), .A(n17285), .B(n17376), .ZN(
        n17286) );
  INV_X1 U20458 ( .A(n17286), .ZN(n17287) );
  OAI211_X1 U20459 ( .C1(n17289), .C2(n18239), .A(n17288), .B(n17287), .ZN(
        P3_U2709) );
  AOI22_X1 U20460 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17331), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17337), .ZN(n17292) );
  OAI211_X1 U20461 ( .C1(n17290), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17407), .B(
        n9712), .ZN(n17291) );
  OAI211_X1 U20462 ( .C1(n17293), .C2(n17402), .A(n17292), .B(n17291), .ZN(
        P3_U2710) );
  INV_X1 U20463 ( .A(n17331), .ZN(n17343) );
  AOI22_X1 U20464 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n17337), .B1(n17410), .B2(
        n17294), .ZN(n17298) );
  OAI211_X1 U20465 ( .C1(n17296), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17407), .B(
        n17295), .ZN(n17297) );
  OAI211_X1 U20466 ( .C1(n17343), .C2(n17510), .A(n17298), .B(n17297), .ZN(
        P3_U2711) );
  AOI22_X1 U20467 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17331), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17337), .ZN(n17302) );
  OAI211_X1 U20468 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17300), .A(n17407), .B(
        n17299), .ZN(n17301) );
  OAI211_X1 U20469 ( .C1(n17303), .C2(n17402), .A(n17302), .B(n17301), .ZN(
        P3_U2712) );
  NAND2_X1 U20470 ( .A1(n17338), .A2(n17432), .ZN(n17310) );
  AOI22_X1 U20471 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17337), .B1(n17410), .B2(
        n17305), .ZN(n17309) );
  NAND2_X1 U20472 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17326), .ZN(n17322) );
  INV_X1 U20473 ( .A(n17322), .ZN(n17318) );
  NAND2_X1 U20474 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17318), .ZN(n17316) );
  NAND2_X1 U20475 ( .A1(n17407), .A2(n17316), .ZN(n17313) );
  OAI21_X1 U20476 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17400), .A(n17313), .ZN(
        n17307) );
  AOI22_X1 U20477 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17331), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17307), .ZN(n17308) );
  OAI211_X1 U20478 ( .C1(n17311), .C2(n17310), .A(n17309), .B(n17308), .ZN(
        P3_U2713) );
  AOI22_X1 U20479 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n17337), .B1(n17410), .B2(
        n17312), .ZN(n17315) );
  INV_X1 U20480 ( .A(n17313), .ZN(n17319) );
  AOI22_X1 U20481 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17331), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(n17319), .ZN(n17314) );
  OAI211_X1 U20482 ( .C1(P3_EAX_REG_21__SCAN_IN), .C2(n17316), .A(n17315), .B(
        n17314), .ZN(P3_U2714) );
  AOI22_X1 U20483 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17337), .B1(n17410), .B2(
        n17317), .ZN(n17321) );
  INV_X1 U20484 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17436) );
  AOI22_X1 U20485 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17319), .B1(n17318), 
        .B2(n17436), .ZN(n17320) );
  OAI211_X1 U20486 ( .C1(n18249), .C2(n17343), .A(n17321), .B(n17320), .ZN(
        P3_U2715) );
  AOI22_X1 U20487 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17331), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17337), .ZN(n17324) );
  OAI211_X1 U20488 ( .C1(n17326), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17407), .B(
        n17322), .ZN(n17323) );
  OAI211_X1 U20489 ( .C1(n17325), .C2(n17402), .A(n17324), .B(n17323), .ZN(
        P3_U2716) );
  AOI22_X1 U20490 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17331), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17337), .ZN(n17329) );
  NAND2_X1 U20491 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17338), .ZN(n17332) );
  AOI211_X1 U20492 ( .C1(n17440), .C2(n17332), .A(n17326), .B(n17376), .ZN(
        n17327) );
  INV_X1 U20493 ( .A(n17327), .ZN(n17328) );
  OAI211_X1 U20494 ( .C1(n17330), .C2(n17402), .A(n17329), .B(n17328), .ZN(
        P3_U2717) );
  AOI22_X1 U20495 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17331), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17337), .ZN(n17334) );
  OAI211_X1 U20496 ( .C1(n17338), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17407), .B(
        n17332), .ZN(n17333) );
  OAI211_X1 U20497 ( .C1(n17335), .C2(n17402), .A(n17334), .B(n17333), .ZN(
        P3_U2718) );
  AOI22_X1 U20498 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n17337), .B1(n17410), .B2(
        n17336), .ZN(n17342) );
  INV_X1 U20499 ( .A(n17338), .ZN(n17339) );
  OAI211_X1 U20500 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17340), .A(n17407), .B(
        n17339), .ZN(n17341) );
  OAI211_X1 U20501 ( .C1(n17343), .C2(n18230), .A(n17342), .B(n17341), .ZN(
        P3_U2719) );
  INV_X1 U20502 ( .A(n17350), .ZN(n17344) );
  OAI33_X1 U20503 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(n17345), .A3(n17350), 
        .B1(n17531), .B2(n17376), .B3(n17344), .ZN(n17346) );
  AOI21_X1 U20504 ( .B1(BUF2_REG_15__SCAN_IN), .B2(n17411), .A(n17346), .ZN(
        n17347) );
  OAI21_X1 U20505 ( .B1(n17348), .B2(n17402), .A(n17347), .ZN(P3_U2720) );
  NAND2_X1 U20506 ( .A1(n18266), .A2(n17375), .ZN(n17355) );
  INV_X1 U20507 ( .A(n17355), .ZN(n17371) );
  NAND2_X1 U20508 ( .A1(n17349), .A2(n17371), .ZN(n17354) );
  INV_X1 U20509 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17526) );
  NAND2_X1 U20510 ( .A1(n17407), .A2(n17350), .ZN(n17353) );
  AOI22_X1 U20511 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17411), .B1(n17410), .B2(
        n17351), .ZN(n17352) );
  OAI221_X1 U20512 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17354), .C1(n17526), 
        .C2(n17353), .A(n17352), .ZN(P3_U2721) );
  INV_X1 U20513 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17457) );
  NOR2_X1 U20514 ( .A1(n17457), .A2(n17355), .ZN(n17374) );
  NAND2_X1 U20515 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17374), .ZN(n17368) );
  NOR2_X1 U20516 ( .A1(n17453), .A2(n17368), .ZN(n17366) );
  NAND2_X1 U20517 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17366), .ZN(n17359) );
  NAND2_X1 U20518 ( .A1(n17359), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n17358) );
  AOI22_X1 U20519 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17411), .B1(n17410), .B2(
        n17356), .ZN(n17357) );
  OAI221_X1 U20520 ( .B1(n17359), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n17358), 
        .C2(n17376), .A(n17357), .ZN(P3_U2722) );
  INV_X1 U20521 ( .A(n17359), .ZN(n17362) );
  AOI21_X1 U20522 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17407), .A(n17366), .ZN(
        n17361) );
  OAI222_X1 U20523 ( .A1(n17405), .A2(n17522), .B1(n17362), .B2(n17361), .C1(
        n17402), .C2(n17360), .ZN(P3_U2723) );
  INV_X1 U20524 ( .A(n17368), .ZN(n17363) );
  AOI21_X1 U20525 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17407), .A(n17363), .ZN(
        n17365) );
  OAI222_X1 U20526 ( .A1(n17405), .A2(n17517), .B1(n17366), .B2(n17365), .C1(
        n17402), .C2(n17364), .ZN(P3_U2724) );
  AOI22_X1 U20527 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17411), .B1(n17410), .B2(
        n17367), .ZN(n17370) );
  OAI211_X1 U20528 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n17374), .A(n17407), .B(
        n17368), .ZN(n17369) );
  NAND2_X1 U20529 ( .A1(n17370), .A2(n17369), .ZN(P3_U2725) );
  AOI21_X1 U20530 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17407), .A(n17371), .ZN(
        n17373) );
  OAI222_X1 U20531 ( .A1(n17405), .A2(n17512), .B1(n17374), .B2(n17373), .C1(
        n17402), .C2(n17372), .ZN(P3_U2726) );
  AOI211_X1 U20532 ( .C1(n17459), .C2(n17377), .A(n17376), .B(n17375), .ZN(
        n17378) );
  AOI21_X1 U20533 ( .B1(n17410), .B2(n17379), .A(n17378), .ZN(n17380) );
  OAI21_X1 U20534 ( .B1(n17510), .B2(n17405), .A(n17380), .ZN(P3_U2727) );
  INV_X1 U20535 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17462) );
  INV_X1 U20536 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17470) );
  NOR3_X1 U20537 ( .A1(n17401), .A2(n17470), .A3(n17400), .ZN(n17404) );
  NAND2_X1 U20538 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17404), .ZN(n17393) );
  NOR2_X1 U20539 ( .A1(n17466), .A2(n17393), .ZN(n17396) );
  NAND2_X1 U20540 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17396), .ZN(n17386) );
  NOR2_X1 U20541 ( .A1(n17462), .A2(n17386), .ZN(n17388) );
  AOI21_X1 U20542 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17407), .A(n17388), .ZN(
        n17385) );
  INV_X1 U20543 ( .A(n17400), .ZN(n17383) );
  AOI22_X1 U20544 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17411), .B1(n17410), .B2(
        n17381), .ZN(n17382) );
  OAI221_X1 U20545 ( .B1(n17385), .B2(n17384), .C1(n17385), .C2(n17383), .A(
        n17382), .ZN(P3_U2728) );
  INV_X1 U20546 ( .A(n17386), .ZN(n17391) );
  AOI21_X1 U20547 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17407), .A(n17391), .ZN(
        n17389) );
  OAI222_X1 U20548 ( .A1(n17405), .A2(n18258), .B1(n17389), .B2(n17388), .C1(
        n17402), .C2(n17387), .ZN(P3_U2729) );
  AOI21_X1 U20549 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17407), .A(n17396), .ZN(
        n17392) );
  OAI222_X1 U20550 ( .A1(n17405), .A2(n18253), .B1(n17392), .B2(n17391), .C1(
        n17402), .C2(n17390), .ZN(P3_U2730) );
  INV_X1 U20551 ( .A(n17393), .ZN(n17399) );
  AOI21_X1 U20552 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17407), .A(n17399), .ZN(
        n17395) );
  OAI222_X1 U20553 ( .A1(n18249), .A2(n17405), .B1(n17396), .B2(n17395), .C1(
        n17402), .C2(n17394), .ZN(P3_U2731) );
  AOI21_X1 U20554 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17407), .A(n17404), .ZN(
        n17398) );
  OAI222_X1 U20555 ( .A1(n18244), .A2(n17405), .B1(n17399), .B2(n17398), .C1(
        n17402), .C2(n17397), .ZN(P3_U2732) );
  NOR2_X1 U20556 ( .A1(n17401), .A2(n17400), .ZN(n17414) );
  AOI21_X1 U20557 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17407), .A(n17414), .ZN(
        n17403) );
  OAI222_X1 U20558 ( .A1(n18240), .A2(n17405), .B1(n17404), .B2(n17403), .C1(
        n17402), .C2(n11237), .ZN(P3_U2733) );
  NOR2_X1 U20559 ( .A1(n17406), .A2(n17476), .ZN(n17408) );
  OAI21_X1 U20560 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n17408), .A(n17407), .ZN(
        n17413) );
  AOI22_X1 U20561 ( .A1(n17411), .A2(BUF2_REG_1__SCAN_IN), .B1(n17410), .B2(
        n17409), .ZN(n17412) );
  OAI21_X1 U20562 ( .B1(n17414), .B2(n17413), .A(n17412), .ZN(P3_U2734) );
  NAND2_X1 U20563 ( .A1(n17416), .A2(n17415), .ZN(n17417) );
  AND2_X1 U20564 ( .A1(n17442), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20565 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17498) );
  NAND2_X1 U20566 ( .A1(n17446), .A2(n17418), .ZN(n17444) );
  AOI22_X1 U20567 ( .A1(n18903), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17472), .ZN(n17419) );
  OAI21_X1 U20568 ( .B1(n17498), .B2(n17444), .A(n17419), .ZN(P3_U2737) );
  INV_X1 U20569 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17496) );
  AOI22_X1 U20570 ( .A1(n18903), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17472), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17420) );
  OAI21_X1 U20571 ( .B1(n17496), .B2(n17444), .A(n17420), .ZN(P3_U2738) );
  AOI22_X1 U20572 ( .A1(n18903), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17472), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17421) );
  OAI21_X1 U20573 ( .B1(n17422), .B2(n17444), .A(n17421), .ZN(P3_U2739) );
  INV_X1 U20574 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17424) );
  AOI22_X1 U20575 ( .A1(n18903), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17442), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17423) );
  OAI21_X1 U20576 ( .B1(n17424), .B2(n17444), .A(n17423), .ZN(P3_U2740) );
  AOI22_X1 U20577 ( .A1(n18903), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17472), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17425) );
  OAI21_X1 U20578 ( .B1(n17426), .B2(n17444), .A(n17425), .ZN(P3_U2741) );
  INV_X1 U20579 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17428) );
  AOI22_X1 U20580 ( .A1(n18903), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17442), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17427) );
  OAI21_X1 U20581 ( .B1(n17428), .B2(n17444), .A(n17427), .ZN(P3_U2742) );
  AOI22_X1 U20582 ( .A1(n18903), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17442), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17429) );
  OAI21_X1 U20583 ( .B1(n9853), .B2(n17444), .A(n17429), .ZN(P3_U2743) );
  INV_X1 U20584 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17489) );
  CLKBUF_X1 U20585 ( .A(n18903), .Z(n17473) );
  AOI22_X1 U20586 ( .A1(n17473), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17472), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17430) );
  OAI21_X1 U20587 ( .B1(n17489), .B2(n17444), .A(n17430), .ZN(P3_U2744) );
  AOI22_X1 U20588 ( .A1(n17473), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17442), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17431) );
  OAI21_X1 U20589 ( .B1(n17432), .B2(n17444), .A(n17431), .ZN(P3_U2745) );
  INV_X1 U20590 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17434) );
  AOI22_X1 U20591 ( .A1(n17473), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17442), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17433) );
  OAI21_X1 U20592 ( .B1(n17434), .B2(n17444), .A(n17433), .ZN(P3_U2746) );
  AOI22_X1 U20593 ( .A1(n17473), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17442), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17435) );
  OAI21_X1 U20594 ( .B1(n17436), .B2(n17444), .A(n17435), .ZN(P3_U2747) );
  INV_X1 U20595 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17438) );
  AOI22_X1 U20596 ( .A1(n17473), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17442), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17437) );
  OAI21_X1 U20597 ( .B1(n17438), .B2(n17444), .A(n17437), .ZN(P3_U2748) );
  AOI22_X1 U20598 ( .A1(n17473), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17442), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17439) );
  OAI21_X1 U20599 ( .B1(n17440), .B2(n17444), .A(n17439), .ZN(P3_U2749) );
  AOI22_X1 U20600 ( .A1(n17473), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17442), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17441) );
  OAI21_X1 U20601 ( .B1(n17482), .B2(n17444), .A(n17441), .ZN(P3_U2750) );
  INV_X1 U20602 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17445) );
  AOI22_X1 U20603 ( .A1(n17473), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17442), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17443) );
  OAI21_X1 U20604 ( .B1(n17445), .B2(n17444), .A(n17443), .ZN(P3_U2751) );
  AOI22_X1 U20605 ( .A1(n17473), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17472), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17447) );
  OAI21_X1 U20606 ( .B1(n17531), .B2(n17475), .A(n17447), .ZN(P3_U2752) );
  AOI22_X1 U20607 ( .A1(n17473), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17472), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17448) );
  OAI21_X1 U20608 ( .B1(n17526), .B2(n17475), .A(n17448), .ZN(P3_U2753) );
  INV_X1 U20609 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17524) );
  AOI22_X1 U20610 ( .A1(n17473), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17472), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17449) );
  OAI21_X1 U20611 ( .B1(n17524), .B2(n17475), .A(n17449), .ZN(P3_U2754) );
  INV_X1 U20612 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17451) );
  AOI22_X1 U20613 ( .A1(n17473), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17472), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17450) );
  OAI21_X1 U20614 ( .B1(n17451), .B2(n17475), .A(n17450), .ZN(P3_U2755) );
  AOI22_X1 U20615 ( .A1(n17473), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17472), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17452) );
  OAI21_X1 U20616 ( .B1(n17453), .B2(n17475), .A(n17452), .ZN(P3_U2756) );
  INV_X1 U20617 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17455) );
  AOI22_X1 U20618 ( .A1(n17473), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17472), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17454) );
  OAI21_X1 U20619 ( .B1(n17455), .B2(n17475), .A(n17454), .ZN(P3_U2757) );
  AOI22_X1 U20620 ( .A1(n17473), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17472), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17456) );
  OAI21_X1 U20621 ( .B1(n17457), .B2(n17475), .A(n17456), .ZN(P3_U2758) );
  AOI22_X1 U20622 ( .A1(n17473), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17472), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17458) );
  OAI21_X1 U20623 ( .B1(n17459), .B2(n17475), .A(n17458), .ZN(P3_U2759) );
  INV_X1 U20624 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17508) );
  AOI22_X1 U20625 ( .A1(n17473), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17472), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17460) );
  OAI21_X1 U20626 ( .B1(n17508), .B2(n17475), .A(n17460), .ZN(P3_U2760) );
  AOI22_X1 U20627 ( .A1(n17473), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17472), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17461) );
  OAI21_X1 U20628 ( .B1(n17462), .B2(n17475), .A(n17461), .ZN(P3_U2761) );
  AOI22_X1 U20629 ( .A1(n17473), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17472), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17463) );
  OAI21_X1 U20630 ( .B1(n17464), .B2(n17475), .A(n17463), .ZN(P3_U2762) );
  AOI22_X1 U20631 ( .A1(n17473), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17472), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17465) );
  OAI21_X1 U20632 ( .B1(n17466), .B2(n17475), .A(n17465), .ZN(P3_U2763) );
  INV_X1 U20633 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17468) );
  AOI22_X1 U20634 ( .A1(n17473), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17472), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17467) );
  OAI21_X1 U20635 ( .B1(n17468), .B2(n17475), .A(n17467), .ZN(P3_U2764) );
  AOI22_X1 U20636 ( .A1(n17473), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17472), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17469) );
  OAI21_X1 U20637 ( .B1(n17470), .B2(n17475), .A(n17469), .ZN(P3_U2765) );
  INV_X1 U20638 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17501) );
  AOI22_X1 U20639 ( .A1(n17473), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17472), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17471) );
  OAI21_X1 U20640 ( .B1(n17501), .B2(n17475), .A(n17471), .ZN(P3_U2766) );
  AOI22_X1 U20641 ( .A1(n17473), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17472), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17474) );
  OAI21_X1 U20642 ( .B1(n17476), .B2(n17475), .A(n17474), .ZN(P3_U2767) );
  INV_X1 U20643 ( .A(n17479), .ZN(n17477) );
  OAI211_X1 U20644 ( .C1(n18907), .C2(n18906), .A(n17478), .B(n17477), .ZN(
        n17518) );
  NAND2_X1 U20645 ( .A1(n18906), .A2(n17478), .ZN(n18740) );
  AOI22_X1 U20646 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17515), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17527), .ZN(n17480) );
  OAI21_X1 U20647 ( .B1(n18230), .B2(n17521), .A(n17480), .ZN(P3_U2768) );
  AOI22_X1 U20648 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17528), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17527), .ZN(n17481) );
  OAI21_X1 U20649 ( .B1(n17482), .B2(n17530), .A(n17481), .ZN(P3_U2769) );
  AOI22_X1 U20650 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17515), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17527), .ZN(n17483) );
  OAI21_X1 U20651 ( .B1(n18240), .B2(n17521), .A(n17483), .ZN(P3_U2770) );
  AOI22_X1 U20652 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17515), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17527), .ZN(n17484) );
  OAI21_X1 U20653 ( .B1(n18244), .B2(n17521), .A(n17484), .ZN(P3_U2771) );
  AOI22_X1 U20654 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17519), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17527), .ZN(n17485) );
  OAI21_X1 U20655 ( .B1(n18249), .B2(n17521), .A(n17485), .ZN(P3_U2772) );
  AOI22_X1 U20656 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17515), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17527), .ZN(n17486) );
  OAI21_X1 U20657 ( .B1(n18253), .B2(n17521), .A(n17486), .ZN(P3_U2773) );
  AOI22_X1 U20658 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17519), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17527), .ZN(n17487) );
  OAI21_X1 U20659 ( .B1(n18258), .B2(n17521), .A(n17487), .ZN(P3_U2774) );
  AOI22_X1 U20660 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17528), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17527), .ZN(n17488) );
  OAI21_X1 U20661 ( .B1(n17489), .B2(n17530), .A(n17488), .ZN(P3_U2775) );
  AOI22_X1 U20662 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17519), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17527), .ZN(n17490) );
  OAI21_X1 U20663 ( .B1(n17510), .B2(n17521), .A(n17490), .ZN(P3_U2776) );
  AOI22_X1 U20664 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17515), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17527), .ZN(n17491) );
  OAI21_X1 U20665 ( .B1(n17512), .B2(n17521), .A(n17491), .ZN(P3_U2777) );
  AOI22_X1 U20666 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17519), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17527), .ZN(n17492) );
  OAI21_X1 U20667 ( .B1(n17514), .B2(n17521), .A(n17492), .ZN(P3_U2778) );
  AOI22_X1 U20668 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17515), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17527), .ZN(n17493) );
  OAI21_X1 U20669 ( .B1(n17517), .B2(n17521), .A(n17493), .ZN(P3_U2779) );
  AOI22_X1 U20670 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17519), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17527), .ZN(n17494) );
  OAI21_X1 U20671 ( .B1(n17522), .B2(n17521), .A(n17494), .ZN(P3_U2780) );
  AOI22_X1 U20672 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17528), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17527), .ZN(n17495) );
  OAI21_X1 U20673 ( .B1(n17496), .B2(n17530), .A(n17495), .ZN(P3_U2781) );
  AOI22_X1 U20674 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17528), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17527), .ZN(n17497) );
  OAI21_X1 U20675 ( .B1(n17498), .B2(n17530), .A(n17497), .ZN(P3_U2782) );
  AOI22_X1 U20676 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17519), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17527), .ZN(n17499) );
  OAI21_X1 U20677 ( .B1(n18230), .B2(n17521), .A(n17499), .ZN(P3_U2783) );
  AOI22_X1 U20678 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17528), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17527), .ZN(n17500) );
  OAI21_X1 U20679 ( .B1(n17501), .B2(n17530), .A(n17500), .ZN(P3_U2784) );
  AOI22_X1 U20680 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17519), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17527), .ZN(n17502) );
  OAI21_X1 U20681 ( .B1(n18240), .B2(n17521), .A(n17502), .ZN(P3_U2785) );
  AOI22_X1 U20682 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17519), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17518), .ZN(n17503) );
  OAI21_X1 U20683 ( .B1(n18244), .B2(n17521), .A(n17503), .ZN(P3_U2786) );
  AOI22_X1 U20684 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17515), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17518), .ZN(n17504) );
  OAI21_X1 U20685 ( .B1(n18249), .B2(n17521), .A(n17504), .ZN(P3_U2787) );
  AOI22_X1 U20686 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17519), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17518), .ZN(n17505) );
  OAI21_X1 U20687 ( .B1(n18253), .B2(n17521), .A(n17505), .ZN(P3_U2788) );
  AOI22_X1 U20688 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17519), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17518), .ZN(n17506) );
  OAI21_X1 U20689 ( .B1(n18258), .B2(n17521), .A(n17506), .ZN(P3_U2789) );
  AOI22_X1 U20690 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17528), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17518), .ZN(n17507) );
  OAI21_X1 U20691 ( .B1(n17508), .B2(n17530), .A(n17507), .ZN(P3_U2790) );
  AOI22_X1 U20692 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17515), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17518), .ZN(n17509) );
  OAI21_X1 U20693 ( .B1(n17510), .B2(n17521), .A(n17509), .ZN(P3_U2791) );
  AOI22_X1 U20694 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17515), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17518), .ZN(n17511) );
  OAI21_X1 U20695 ( .B1(n17512), .B2(n17521), .A(n17511), .ZN(P3_U2792) );
  AOI22_X1 U20696 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17519), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17518), .ZN(n17513) );
  OAI21_X1 U20697 ( .B1(n17514), .B2(n17521), .A(n17513), .ZN(P3_U2793) );
  AOI22_X1 U20698 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17515), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17518), .ZN(n17516) );
  OAI21_X1 U20699 ( .B1(n17517), .B2(n17521), .A(n17516), .ZN(P3_U2794) );
  AOI22_X1 U20700 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17519), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17518), .ZN(n17520) );
  OAI21_X1 U20701 ( .B1(n17522), .B2(n17521), .A(n17520), .ZN(P3_U2795) );
  AOI22_X1 U20702 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17528), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17527), .ZN(n17523) );
  OAI21_X1 U20703 ( .B1(n17524), .B2(n17530), .A(n17523), .ZN(P3_U2796) );
  AOI22_X1 U20704 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17528), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17527), .ZN(n17525) );
  OAI21_X1 U20705 ( .B1(n17526), .B2(n17530), .A(n17525), .ZN(P3_U2797) );
  AOI22_X1 U20706 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17528), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17527), .ZN(n17529) );
  OAI21_X1 U20707 ( .B1(n17531), .B2(n17530), .A(n17529), .ZN(P3_U2798) );
  NAND2_X1 U20708 ( .A1(n17562), .A2(n17534), .ZN(n17548) );
  OAI21_X1 U20709 ( .B1(n17532), .B2(n17896), .A(n17897), .ZN(n17533) );
  AOI21_X1 U20710 ( .B1(n17859), .B2(n17538), .A(n17533), .ZN(n17565) );
  OAI21_X1 U20711 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17642), .A(
        n17565), .ZN(n17550) );
  AOI22_X1 U20712 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17737), .B1(
        n17805), .B2(n17534), .ZN(n17536) );
  AOI211_X1 U20713 ( .C1(n17537), .C2(n17536), .A(n17535), .B(n17780), .ZN(
        n17544) );
  NOR2_X1 U20714 ( .A1(n17729), .A2(n17538), .ZN(n17556) );
  OAI211_X1 U20715 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17556), .B(n17539), .ZN(n17541) );
  OAI211_X1 U20716 ( .C1(n17746), .C2(n17542), .A(n17541), .B(n17540), .ZN(
        n17543) );
  AOI211_X1 U20717 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17550), .A(
        n17544), .B(n17543), .ZN(n17547) );
  NAND2_X1 U20718 ( .A1(n17901), .A2(n17809), .ZN(n17638) );
  AOI22_X1 U20719 ( .A1(n17888), .A2(n17911), .B1(n17761), .B2(n17545), .ZN(
        n17568) );
  NAND2_X1 U20720 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17568), .ZN(
        n17557) );
  NAND3_X1 U20721 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17638), .A3(
        n17557), .ZN(n17546) );
  OAI211_X1 U20722 ( .C1(n17549), .C2(n17548), .A(n17547), .B(n17546), .ZN(
        P3_U2802) );
  AOI22_X1 U20723 ( .A1(n17644), .A2(n17551), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n17550), .ZN(n17561) );
  NOR2_X1 U20724 ( .A1(n17553), .A2(n17552), .ZN(n17554) );
  XNOR2_X1 U20725 ( .A(n17805), .B(n17554), .ZN(n17914) );
  AOI22_X1 U20726 ( .A1(n17806), .A2(n17914), .B1(n17556), .B2(n17555), .ZN(
        n17560) );
  OAI221_X1 U20727 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17558), 
        .C1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n17562), .A(n17557), .ZN(
        n17559) );
  NAND2_X1 U20728 ( .A1(n9647), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17916) );
  NAND4_X1 U20729 ( .A1(n17561), .A2(n17560), .A3(n17559), .A4(n17916), .ZN(
        P3_U2803) );
  INV_X1 U20730 ( .A(n17562), .ZN(n17608) );
  NAND3_X1 U20731 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17929), .A3(
        n17925), .ZN(n17922) );
  AOI21_X1 U20732 ( .B1(n17563), .B2(n18257), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17564) );
  OAI22_X1 U20733 ( .A1(n17673), .A2(n17566), .B1(n17565), .B2(n17564), .ZN(
        n17570) );
  XNOR2_X1 U20734 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n17567), .ZN(
        n17919) );
  OAI22_X1 U20735 ( .A1(n17568), .A2(n17925), .B1(n17919), .B2(n17780), .ZN(
        n17569) );
  AOI211_X1 U20736 ( .C1(n9647), .C2(P3_REIP_REG_26__SCAN_IN), .A(n17570), .B(
        n17569), .ZN(n17571) );
  OAI21_X1 U20737 ( .B1(n17608), .B2(n17922), .A(n17571), .ZN(P3_U2804) );
  AOI21_X1 U20738 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n9774), .A(
        n17896), .ZN(n17572) );
  AOI211_X1 U20739 ( .C1(n18257), .C2(n17580), .A(n17857), .B(n17572), .ZN(
        n17604) );
  OAI21_X1 U20740 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17642), .A(
        n17604), .ZN(n17586) );
  AOI22_X1 U20741 ( .A1(n17644), .A2(n17573), .B1(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n17586), .ZN(n17584) );
  AOI21_X1 U20742 ( .B1(n17805), .B2(n17575), .A(n17574), .ZN(n17576) );
  XNOR2_X1 U20743 ( .A(n17576), .B(n17926), .ZN(n17938) );
  XNOR2_X1 U20744 ( .A(n17577), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17940) );
  XNOR2_X1 U20745 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17578), .ZN(
        n17936) );
  OAI22_X1 U20746 ( .A1(n17901), .A2(n17940), .B1(n17809), .B2(n17936), .ZN(
        n17579) );
  AOI21_X1 U20747 ( .B1(n17806), .B2(n17938), .A(n17579), .ZN(n17583) );
  NAND2_X1 U20748 ( .A1(n9647), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17934) );
  NOR2_X1 U20749 ( .A1(n17729), .A2(n17580), .ZN(n17588) );
  OAI211_X1 U20750 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17588), .B(n17581), .ZN(n17582) );
  NAND4_X1 U20751 ( .A1(n17584), .A2(n17583), .A3(n17934), .A4(n17582), .ZN(
        P3_U2805) );
  INV_X1 U20752 ( .A(n17585), .ZN(n17597) );
  NOR2_X1 U20753 ( .A1(n18217), .A2(n18821), .ZN(n17943) );
  AOI221_X1 U20754 ( .B1(n17588), .B2(n17587), .C1(n17586), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17943), .ZN(n17596) );
  NOR3_X1 U20755 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17941), .A3(
        n17589), .ZN(n17594) );
  AOI22_X1 U20756 ( .A1(n17888), .A2(n17945), .B1(n17761), .B2(n17947), .ZN(
        n17607) );
  AOI21_X1 U20757 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17591), .A(
        n17590), .ZN(n17955) );
  OAI22_X1 U20758 ( .A1(n17607), .A2(n17592), .B1(n17955), .B2(n17780), .ZN(
        n17593) );
  AOI21_X1 U20759 ( .B1(n17594), .B2(n17773), .A(n17593), .ZN(n17595) );
  OAI211_X1 U20760 ( .C1(n17746), .C2(n17597), .A(n17596), .B(n17595), .ZN(
        P3_U2806) );
  OAI21_X1 U20761 ( .B1(n17667), .B2(n17598), .A(n17610), .ZN(n17599) );
  OAI211_X1 U20762 ( .C1(n17805), .C2(n17974), .A(n17636), .B(n17599), .ZN(
        n17600) );
  XNOR2_X1 U20763 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n17600), .ZN(
        n17960) );
  AOI21_X1 U20764 ( .B1(n9774), .B2(n18257), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17603) );
  OAI21_X1 U20765 ( .B1(n17644), .B2(n17614), .A(n17601), .ZN(n17602) );
  NAND2_X1 U20766 ( .A1(n9647), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17961) );
  OAI211_X1 U20767 ( .C1(n17604), .C2(n17603), .A(n17602), .B(n17961), .ZN(
        n17605) );
  AOI21_X1 U20768 ( .B1(n17806), .B2(n17960), .A(n17605), .ZN(n17606) );
  OAI221_X1 U20769 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17608), 
        .C1(n17956), .C2(n17607), .A(n17606), .ZN(P3_U2807) );
  OAI22_X1 U20770 ( .A1(n17968), .A2(n17901), .B1(n17969), .B2(n17809), .ZN(
        n17683) );
  AOI21_X1 U20771 ( .B1(n17965), .B2(n17638), .A(n17683), .ZN(n17631) );
  AOI221_X1 U20772 ( .B1(n17684), .B2(n17610), .C1(n17965), .C2(n17610), .A(
        n17609), .ZN(n17611) );
  XNOR2_X1 U20773 ( .A(n17611), .B(n17974), .ZN(n17975) );
  NOR3_X1 U20774 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17965), .A3(
        n17696), .ZN(n17622) );
  AOI22_X1 U20775 ( .A1(n17859), .A2(n17615), .B1(n17725), .B2(n17612), .ZN(
        n17613) );
  NAND2_X1 U20776 ( .A1(n17613), .A2(n17897), .ZN(n17640) );
  AOI21_X1 U20777 ( .B1(n17614), .B2(n9951), .A(n17640), .ZN(n17624) );
  OR2_X1 U20778 ( .A1(n17615), .A2(n17729), .ZN(n17626) );
  AOI21_X1 U20779 ( .B1(n17625), .B2(n17620), .A(n17626), .ZN(n17617) );
  AOI22_X1 U20780 ( .A1(n17644), .A2(n17618), .B1(n17617), .B2(n17616), .ZN(
        n17619) );
  NAND2_X1 U20781 ( .A1(n9647), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17976) );
  OAI211_X1 U20782 ( .C1(n17624), .C2(n17620), .A(n17619), .B(n17976), .ZN(
        n17621) );
  AOI211_X1 U20783 ( .C1(n17975), .C2(n17806), .A(n17622), .B(n17621), .ZN(
        n17623) );
  OAI21_X1 U20784 ( .B1(n17631), .B2(n17974), .A(n17623), .ZN(P3_U2808) );
  NAND2_X1 U20785 ( .A1(n17981), .A2(n17630), .ZN(n17983) );
  INV_X1 U20786 ( .A(n17696), .ZN(n17668) );
  NAND2_X1 U20787 ( .A1(n17904), .A2(n17668), .ZN(n17659) );
  NAND2_X1 U20788 ( .A1(n9647), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n17987) );
  OAI221_X1 U20789 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17626), .C1(
        n17625), .C2(n17624), .A(n17987), .ZN(n17633) );
  AND3_X1 U20790 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17805), .A3(
        n17627), .ZN(n17648) );
  AOI22_X1 U20791 ( .A1(n17981), .A2(n17648), .B1(n17628), .B2(n17667), .ZN(
        n17629) );
  XNOR2_X1 U20792 ( .A(n17629), .B(n17630), .ZN(n17989) );
  OAI22_X1 U20793 ( .A1(n17631), .A2(n17630), .B1(n17989), .B2(n17780), .ZN(
        n17632) );
  AOI211_X1 U20794 ( .C1(n17644), .C2(n17634), .A(n17633), .B(n17632), .ZN(
        n17635) );
  OAI21_X1 U20795 ( .B1(n17983), .B2(n17659), .A(n17635), .ZN(P3_U2809) );
  OAI221_X1 U20796 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17665), 
        .C1(n18008), .C2(n17648), .A(n17636), .ZN(n17637) );
  XNOR2_X1 U20797 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17637), .ZN(
        n17997) );
  NAND2_X1 U20798 ( .A1(n17904), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17994) );
  AOI21_X1 U20799 ( .B1(n17638), .B2(n17994), .A(n17683), .ZN(n17658) );
  NAND2_X1 U20800 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17966), .ZN(
        n18002) );
  OAI22_X1 U20801 ( .A1(n17658), .A2(n17966), .B1(n17659), .B2(n18002), .ZN(
        n17639) );
  AOI21_X1 U20802 ( .B1(n17806), .B2(n17997), .A(n17639), .ZN(n17647) );
  NAND2_X1 U20803 ( .A1(n9647), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17999) );
  OAI221_X1 U20804 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17641), .C1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n18257), .A(n17640), .ZN(
        n17646) );
  OAI21_X1 U20805 ( .B1(n17644), .B2(n17614), .A(n17643), .ZN(n17645) );
  NAND4_X1 U20806 ( .A1(n17647), .A2(n17999), .A3(n17646), .A4(n17645), .ZN(
        P3_U2810) );
  AOI21_X1 U20807 ( .B1(n17667), .B2(n17665), .A(n17648), .ZN(n17649) );
  XNOR2_X1 U20808 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n17649), .ZN(
        n18004) );
  AOI21_X1 U20809 ( .B1(n17859), .B2(n17651), .A(n17857), .ZN(n17681) );
  OAI21_X1 U20810 ( .B1(n17650), .B2(n17896), .A(n17681), .ZN(n17662) );
  AOI22_X1 U20811 ( .A1(n9647), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17662), .ZN(n17654) );
  NOR2_X1 U20812 ( .A1(n17729), .A2(n17651), .ZN(n17664) );
  OAI211_X1 U20813 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17664), .B(n17652), .ZN(n17653) );
  OAI211_X1 U20814 ( .C1(n17746), .C2(n17655), .A(n17654), .B(n17653), .ZN(
        n17656) );
  AOI21_X1 U20815 ( .B1(n17806), .B2(n18004), .A(n17656), .ZN(n17657) );
  OAI221_X1 U20816 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17659), 
        .C1(n18008), .C2(n17658), .A(n17657), .ZN(P3_U2811) );
  AOI21_X1 U20817 ( .B1(n17668), .B2(n18012), .A(n17683), .ZN(n17677) );
  OAI22_X1 U20818 ( .A1(n18217), .A2(n18809), .B1(n17746), .B2(n17660), .ZN(
        n17661) );
  AOI221_X1 U20819 ( .B1(n17664), .B2(n17663), .C1(n17662), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17661), .ZN(n17670) );
  AOI21_X1 U20820 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17805), .A(
        n17665), .ZN(n17666) );
  XOR2_X1 U20821 ( .A(n17667), .B(n17666), .Z(n18023) );
  NOR2_X1 U20822 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18012), .ZN(
        n18022) );
  AOI22_X1 U20823 ( .A1(n17806), .A2(n18023), .B1(n17668), .B2(n18022), .ZN(
        n17669) );
  OAI211_X1 U20824 ( .C1(n17677), .C2(n17671), .A(n17670), .B(n17669), .ZN(
        P3_U2812) );
  AOI21_X1 U20825 ( .B1(n17672), .B2(n18257), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17682) );
  AOI22_X1 U20826 ( .A1(n9647), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n17674), 
        .B2(n17890), .ZN(n17680) );
  OAI21_X1 U20827 ( .B1(n17676), .B2(n18016), .A(n17675), .ZN(n18026) );
  NAND2_X1 U20828 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18016), .ZN(
        n18031) );
  OAI22_X1 U20829 ( .A1(n17677), .A2(n18016), .B1(n17696), .B2(n18031), .ZN(
        n17678) );
  AOI21_X1 U20830 ( .B1(n17806), .B2(n18026), .A(n17678), .ZN(n17679) );
  OAI211_X1 U20831 ( .C1(n17682), .C2(n17681), .A(n17680), .B(n17679), .ZN(
        P3_U2813) );
  INV_X1 U20832 ( .A(n17683), .ZN(n17695) );
  NOR2_X1 U20833 ( .A1(n17737), .A2(n17760), .ZN(n17781) );
  AOI22_X1 U20834 ( .A1(n17685), .A2(n17781), .B1(n17684), .B2(n17737), .ZN(
        n17686) );
  XNOR2_X1 U20835 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17686), .ZN(
        n18042) );
  AOI21_X1 U20836 ( .B1(n17859), .B2(n17688), .A(n17857), .ZN(n17714) );
  OAI21_X1 U20837 ( .B1(n17687), .B2(n17896), .A(n17714), .ZN(n17703) );
  AOI22_X1 U20838 ( .A1(n9647), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17703), .ZN(n17691) );
  NOR2_X1 U20839 ( .A1(n17729), .A2(n17688), .ZN(n17705) );
  OAI211_X1 U20840 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17705), .B(n17689), .ZN(n17690) );
  OAI211_X1 U20841 ( .C1(n17746), .C2(n17692), .A(n17691), .B(n17690), .ZN(
        n17693) );
  AOI21_X1 U20842 ( .B1(n17806), .B2(n18042), .A(n17693), .ZN(n17694) );
  OAI221_X1 U20843 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17696), 
        .C1(n18040), .C2(n17695), .A(n17694), .ZN(P3_U2814) );
  INV_X1 U20844 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18063) );
  NOR2_X1 U20845 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17698) );
  NOR2_X1 U20846 ( .A1(n17805), .A2(n17697), .ZN(n17782) );
  NAND2_X1 U20847 ( .A1(n17698), .A2(n17782), .ZN(n17764) );
  NOR2_X1 U20848 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17764), .ZN(
        n17743) );
  INV_X1 U20849 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17723) );
  NAND2_X1 U20850 ( .A1(n17743), .A2(n17723), .ZN(n17719) );
  OAI21_X1 U20851 ( .B1(n17736), .B2(n17716), .A(n17719), .ZN(n17699) );
  OAI221_X1 U20852 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18063), 
        .C1(n18084), .C2(n17805), .A(n17699), .ZN(n17700) );
  XNOR2_X1 U20853 ( .A(n18056), .B(n17700), .ZN(n18050) );
  OAI22_X1 U20854 ( .A1(n18217), .A2(n18803), .B1(n17746), .B2(n17701), .ZN(
        n17702) );
  AOI221_X1 U20855 ( .B1(n17705), .B2(n17704), .C1(n17703), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17702), .ZN(n17709) );
  INV_X1 U20856 ( .A(n17716), .ZN(n17706) );
  NOR2_X1 U20857 ( .A1(n18082), .A2(n18084), .ZN(n17724) );
  INV_X1 U20858 ( .A(n17724), .ZN(n18057) );
  NOR2_X1 U20859 ( .A1(n17762), .A2(n18057), .ZN(n18077) );
  NAND2_X1 U20860 ( .A1(n17706), .A2(n18077), .ZN(n17710) );
  AOI21_X1 U20861 ( .B1(n18056), .B2(n17710), .A(n17968), .ZN(n18053) );
  NOR2_X1 U20862 ( .A1(n17969), .A2(n17809), .ZN(n17707) );
  INV_X1 U20863 ( .A(n17760), .ZN(n18093) );
  NAND2_X1 U20864 ( .A1(n18093), .A2(n17724), .ZN(n18073) );
  OAI21_X1 U20865 ( .B1(n17716), .B2(n18073), .A(n18056), .ZN(n18048) );
  AOI22_X1 U20866 ( .A1(n17888), .A2(n18053), .B1(n17707), .B2(n18048), .ZN(
        n17708) );
  OAI211_X1 U20867 ( .C1(n17780), .C2(n18050), .A(n17709), .B(n17708), .ZN(
        P3_U2815) );
  NAND2_X1 U20868 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17724), .ZN(
        n17718) );
  INV_X1 U20869 ( .A(n17718), .ZN(n18058) );
  OAI221_X1 U20870 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18058), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n9804), .A(n17710), .ZN(
        n18070) );
  AOI21_X1 U20871 ( .B1(n17711), .B2(n18257), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17713) );
  OAI22_X1 U20872 ( .A1(n17714), .A2(n17713), .B1(n17673), .B2(n17712), .ZN(
        n17715) );
  AOI21_X1 U20873 ( .B1(n9647), .B2(P3_REIP_REG_14__SCAN_IN), .A(n17715), .ZN(
        n17722) );
  NOR2_X1 U20874 ( .A1(n17716), .A2(n18073), .ZN(n17717) );
  AOI221_X1 U20875 ( .B1(n17723), .B2(n18063), .C1(n18073), .C2(n18063), .A(
        n17717), .ZN(n18065) );
  INV_X1 U20876 ( .A(n17781), .ZN(n17765) );
  OAI22_X1 U20877 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17719), .B1(
        n17718), .B2(n17765), .ZN(n17720) );
  XNOR2_X1 U20878 ( .A(n18063), .B(n17720), .ZN(n18067) );
  AOI22_X1 U20879 ( .A1(n17761), .A2(n18065), .B1(n17806), .B2(n18067), .ZN(
        n17721) );
  OAI211_X1 U20880 ( .C1(n17901), .C2(n18070), .A(n17722), .B(n17721), .ZN(
        P3_U2816) );
  INV_X1 U20881 ( .A(n17773), .ZN(n17792) );
  NAND2_X1 U20882 ( .A1(n17724), .A2(n17723), .ZN(n18081) );
  AOI21_X1 U20883 ( .B1(n17859), .B2(n17728), .A(n17725), .ZN(n17726) );
  OAI21_X1 U20884 ( .B1(n17727), .B2(n17726), .A(n17897), .ZN(n17748) );
  NOR2_X1 U20885 ( .A1(n17729), .A2(n17728), .ZN(n17750) );
  OAI211_X1 U20886 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17750), .B(n17730), .ZN(n17732) );
  NAND2_X1 U20887 ( .A1(n9647), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17731) );
  OAI211_X1 U20888 ( .C1(n17746), .C2(n17733), .A(n17732), .B(n17731), .ZN(
        n17734) );
  AOI21_X1 U20889 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17748), .A(
        n17734), .ZN(n17742) );
  INV_X1 U20890 ( .A(n18073), .ZN(n17735) );
  OAI22_X1 U20891 ( .A1(n17735), .A2(n17809), .B1(n18077), .B2(n17901), .ZN(
        n17752) );
  INV_X1 U20892 ( .A(n17736), .ZN(n17739) );
  NOR2_X1 U20893 ( .A1(n18084), .A2(n17737), .ZN(n17738) );
  OAI22_X1 U20894 ( .A1(n17739), .A2(n18084), .B1(n17743), .B2(n17738), .ZN(
        n17740) );
  XNOR2_X1 U20895 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17740), .ZN(
        n18071) );
  AOI22_X1 U20896 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17752), .B1(
        n17806), .B2(n18071), .ZN(n17741) );
  OAI211_X1 U20897 ( .C1(n17792), .C2(n18081), .A(n17742), .B(n17741), .ZN(
        P3_U2817) );
  AOI21_X1 U20898 ( .B1(n17781), .B2(n18072), .A(n17743), .ZN(n17744) );
  XNOR2_X1 U20899 ( .A(n17744), .B(n18084), .ZN(n18088) );
  OAI22_X1 U20900 ( .A1(n18217), .A2(n18797), .B1(n17746), .B2(n17745), .ZN(
        n17747) );
  AOI221_X1 U20901 ( .B1(n17750), .B2(n17749), .C1(n17748), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17747), .ZN(n17754) );
  NOR2_X1 U20902 ( .A1(n17792), .A2(n18082), .ZN(n17751) );
  AOI22_X1 U20903 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17752), .B1(
        n17751), .B2(n18084), .ZN(n17753) );
  OAI211_X1 U20904 ( .C1(n18088), .C2(n17780), .A(n17754), .B(n17753), .ZN(
        P3_U2818) );
  OR2_X1 U20905 ( .A1(n18096), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18101) );
  NOR3_X1 U20906 ( .A1(n17821), .A2(n17827), .A3(n18263), .ZN(n17813) );
  NAND2_X1 U20907 ( .A1(n17755), .A2(n17813), .ZN(n17772) );
  NAND3_X1 U20908 ( .A1(n17891), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A3(
        n17772), .ZN(n17757) );
  NAND2_X1 U20909 ( .A1(n9647), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n17756) );
  OAI211_X1 U20910 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n17772), .A(
        n17757), .B(n17756), .ZN(n17758) );
  AOI21_X1 U20911 ( .B1(n17759), .B2(n17890), .A(n17758), .ZN(n17768) );
  AOI22_X1 U20912 ( .A1(n17888), .A2(n17762), .B1(n17761), .B2(n17760), .ZN(
        n17791) );
  OAI21_X1 U20913 ( .B1(n17763), .B2(n17792), .A(n17791), .ZN(n17776) );
  OAI21_X1 U20914 ( .B1(n17765), .B2(n18096), .A(n17764), .ZN(n17766) );
  XOR2_X1 U20915 ( .A(n17766), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(
        n18089) );
  AOI22_X1 U20916 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17776), .B1(
        n17806), .B2(n18089), .ZN(n17767) );
  OAI211_X1 U20917 ( .C1(n17792), .C2(n18101), .A(n17768), .B(n17767), .ZN(
        P3_U2819) );
  AOI22_X1 U20918 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17781), .B1(
        n17782), .B2(n9943), .ZN(n17769) );
  XOR2_X1 U20919 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n17769), .Z(
        n18110) );
  NAND3_X1 U20920 ( .A1(n17784), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        n17813), .ZN(n17785) );
  OAI21_X1 U20921 ( .B1(n17822), .B2(n17770), .A(n17785), .ZN(n17771) );
  AOI22_X1 U20922 ( .A1(n9647), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n17772), 
        .B2(n17771), .ZN(n17779) );
  AOI21_X1 U20923 ( .B1(n17773), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17774) );
  INV_X1 U20924 ( .A(n17774), .ZN(n17777) );
  AOI22_X1 U20925 ( .A1(n17777), .A2(n17776), .B1(n17775), .B2(n17890), .ZN(
        n17778) );
  OAI211_X1 U20926 ( .C1(n18110), .C2(n17780), .A(n17779), .B(n17778), .ZN(
        P3_U2820) );
  NOR2_X1 U20927 ( .A1(n17782), .A2(n17781), .ZN(n17783) );
  XNOR2_X1 U20928 ( .A(n17783), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18117) );
  AND2_X1 U20929 ( .A1(n17784), .A2(n17813), .ZN(n17786) );
  OAI211_X1 U20930 ( .C1(n17786), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n17891), .B(n17785), .ZN(n17787) );
  NAND2_X1 U20931 ( .A1(n9647), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n18118) );
  OAI211_X1 U20932 ( .C1(n17673), .C2(n17788), .A(n17787), .B(n18118), .ZN(
        n17789) );
  AOI21_X1 U20933 ( .B1(n17806), .B2(n18117), .A(n17789), .ZN(n17790) );
  OAI221_X1 U20934 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17792), .C1(
        n9943), .C2(n17791), .A(n17790), .ZN(P3_U2821) );
  INV_X1 U20935 ( .A(n17859), .ZN(n17793) );
  OAI21_X1 U20936 ( .B1(n17794), .B2(n17793), .A(n17897), .ZN(n17814) );
  NOR2_X1 U20937 ( .A1(n17795), .A2(n17812), .ZN(n17797) );
  OAI211_X1 U20938 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17797), .A(
        n18257), .B(n17796), .ZN(n17798) );
  NAND2_X1 U20939 ( .A1(n9647), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18127) );
  OAI211_X1 U20940 ( .C1(n17673), .C2(n17799), .A(n17798), .B(n18127), .ZN(
        n17800) );
  AOI21_X1 U20941 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17814), .A(
        n17800), .ZN(n17808) );
  AOI21_X1 U20942 ( .B1(n17802), .B2(n18130), .A(n17801), .ZN(n18132) );
  OAI21_X1 U20943 ( .B1(n17805), .B2(n17804), .A(n17803), .ZN(n18133) );
  AOI22_X1 U20944 ( .A1(n17888), .A2(n18132), .B1(n17806), .B2(n18133), .ZN(
        n17807) );
  OAI211_X1 U20945 ( .C1(n17809), .C2(n18138), .A(n17808), .B(n17807), .ZN(
        P3_U2822) );
  OAI21_X1 U20946 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17811), .A(
        n17810), .ZN(n18147) );
  NOR2_X1 U20947 ( .A1(n18217), .A2(n18787), .ZN(n18139) );
  AOI221_X1 U20948 ( .B1(n17814), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n17813), .C2(n17812), .A(n18139), .ZN(n17820) );
  NAND2_X1 U20949 ( .A1(n17816), .A2(n17815), .ZN(n17817) );
  XNOR2_X1 U20950 ( .A(n17817), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18143) );
  AOI22_X1 U20951 ( .A1(n17888), .A2(n18143), .B1(n17818), .B2(n17890), .ZN(
        n17819) );
  OAI211_X1 U20952 ( .C1(n9676), .C2(n18147), .A(n17820), .B(n17819), .ZN(
        P3_U2823) );
  NOR2_X1 U20953 ( .A1(n17821), .A2(n18263), .ZN(n17828) );
  NOR2_X1 U20954 ( .A1(n17822), .A2(n17828), .ZN(n17846) );
  OAI21_X1 U20955 ( .B1(n17825), .B2(n17824), .A(n17823), .ZN(n18155) );
  OAI22_X1 U20956 ( .A1(n9676), .A2(n18155), .B1(n18217), .B2(n18785), .ZN(
        n17826) );
  AOI221_X1 U20957 ( .B1(n17846), .B2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C1(
        n17828), .C2(n17827), .A(n17826), .ZN(n17832) );
  AOI21_X1 U20958 ( .B1(n18150), .B2(n17830), .A(n17829), .ZN(n18153) );
  NAND2_X1 U20959 ( .A1(n17888), .A2(n18153), .ZN(n17831) );
  OAI211_X1 U20960 ( .C1(n17673), .C2(n17833), .A(n17832), .B(n17831), .ZN(
        P3_U2824) );
  OAI21_X1 U20961 ( .B1(n17836), .B2(n17835), .A(n17834), .ZN(n17838) );
  XNOR2_X1 U20962 ( .A(n17838), .B(n17837), .ZN(n18164) );
  AOI21_X1 U20963 ( .B1(n17841), .B2(n17840), .A(n17839), .ZN(n18162) );
  AOI22_X1 U20964 ( .A1(n17888), .A2(n18162), .B1(n9647), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17848) );
  OAI21_X1 U20965 ( .B1(n17857), .B2(n17843), .A(n17842), .ZN(n17845) );
  AOI22_X1 U20966 ( .A1(n17846), .A2(n17845), .B1(n17844), .B2(n17890), .ZN(
        n17847) );
  OAI211_X1 U20967 ( .C1(n9676), .C2(n18164), .A(n17848), .B(n17847), .ZN(
        P3_U2825) );
  OAI21_X1 U20968 ( .B1(n17851), .B2(n17850), .A(n17849), .ZN(n18168) );
  INV_X1 U20969 ( .A(n17852), .ZN(n17854) );
  NOR2_X1 U20970 ( .A1(n17854), .A2(n17853), .ZN(n17855) );
  XNOR2_X1 U20971 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n17855), .ZN(
        n18174) );
  OAI22_X1 U20972 ( .A1(n17901), .A2(n18174), .B1(n18263), .B2(n17856), .ZN(
        n17863) );
  AOI21_X1 U20973 ( .B1(n17859), .B2(n17858), .A(n17857), .ZN(n17870) );
  OAI22_X1 U20974 ( .A1(n17673), .A2(n17861), .B1(n17860), .B2(n17870), .ZN(
        n17862) );
  AOI211_X1 U20975 ( .C1(n9647), .C2(P3_REIP_REG_4__SCAN_IN), .A(n17863), .B(
        n17862), .ZN(n17864) );
  OAI21_X1 U20976 ( .B1(n9676), .B2(n18168), .A(n17864), .ZN(P3_U2826) );
  OAI21_X1 U20977 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17866), .A(
        n17865), .ZN(n18179) );
  AOI21_X1 U20978 ( .B1(n17869), .B2(n17868), .A(n17867), .ZN(n18182) );
  AOI21_X1 U20979 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17897), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17871) );
  OAI22_X1 U20980 ( .A1(n17673), .A2(n17872), .B1(n17871), .B2(n17870), .ZN(
        n17873) );
  AOI21_X1 U20981 ( .B1(n17888), .B2(n18182), .A(n17873), .ZN(n17874) );
  NAND2_X1 U20982 ( .A1(n9647), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18178) );
  OAI211_X1 U20983 ( .C1(n9676), .C2(n18179), .A(n17874), .B(n18178), .ZN(
        P3_U2827) );
  AOI21_X1 U20984 ( .B1(n17877), .B2(n17876), .A(n17875), .ZN(n18197) );
  NOR2_X1 U20985 ( .A1(n18217), .A2(n18777), .ZN(n18185) );
  OAI21_X1 U20986 ( .B1(n17880), .B2(n17879), .A(n17878), .ZN(n18201) );
  OAI22_X1 U20987 ( .A1(n17673), .A2(n17881), .B1(n9676), .B2(n18201), .ZN(
        n17882) );
  AOI211_X1 U20988 ( .C1(n17888), .C2(n18197), .A(n18185), .B(n17882), .ZN(
        n17883) );
  OAI221_X1 U20989 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18263), .C1(
        n17884), .C2(n17897), .A(n17883), .ZN(P3_U2828) );
  OAI21_X1 U20990 ( .B1(n17886), .B2(n17894), .A(n17885), .ZN(n18211) );
  NAND2_X1 U20991 ( .A1(n18884), .A2(n17895), .ZN(n17887) );
  XNOR2_X1 U20992 ( .A(n17887), .B(n17886), .ZN(n18207) );
  AOI22_X1 U20993 ( .A1(n17888), .A2(n18207), .B1(n9647), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17893) );
  AOI22_X1 U20994 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17891), .B1(
        n17890), .B2(n17889), .ZN(n17892) );
  OAI211_X1 U20995 ( .C1(n9676), .C2(n18211), .A(n17893), .B(n17892), .ZN(
        P3_U2829) );
  AOI21_X1 U20996 ( .B1(n17895), .B2(n18884), .A(n17894), .ZN(n18215) );
  INV_X1 U20997 ( .A(n18215), .ZN(n18213) );
  NAND3_X1 U20998 ( .A1(n18865), .A2(n17897), .A3(n17896), .ZN(n17898) );
  AOI22_X1 U20999 ( .A1(n9647), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17898), .ZN(n17899) );
  OAI221_X1 U21000 ( .B1(n18215), .B2(n17901), .C1(n18213), .C2(n9676), .A(
        n17899), .ZN(P3_U2830) );
  NOR2_X1 U21001 ( .A1(n17902), .A2(n17957), .ZN(n17913) );
  NOR2_X1 U21002 ( .A1(n17903), .A2(n18092), .ZN(n17910) );
  NOR2_X1 U21003 ( .A1(n9640), .A2(n18219), .ZN(n18015) );
  NAND2_X1 U21004 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18032), .ZN(
        n18113) );
  NOR2_X1 U21005 ( .A1(n18021), .A2(n18113), .ZN(n18038) );
  NAND2_X1 U21006 ( .A1(n17904), .A2(n18038), .ZN(n17990) );
  OAI21_X1 U21007 ( .B1(n17905), .B2(n17990), .A(n9640), .ZN(n17971) );
  NAND2_X1 U21008 ( .A1(n17906), .A2(n17971), .ZN(n17946) );
  INV_X1 U21009 ( .A(n18015), .ZN(n18191) );
  OAI21_X1 U21010 ( .B1(n17927), .B2(n17946), .A(n18191), .ZN(n17931) );
  OAI211_X1 U21011 ( .C1(n17908), .C2(n18015), .A(n17931), .B(n17907), .ZN(
        n17909) );
  AOI211_X1 U21012 ( .C1(n18722), .C2(n17911), .A(n17910), .B(n17909), .ZN(
        n17921) );
  INV_X1 U21013 ( .A(n17921), .ZN(n17912) );
  MUX2_X1 U21014 ( .A(n17913), .B(n17912), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n17915) );
  AOI22_X1 U21015 ( .A1(n18196), .A2(n17915), .B1(n18134), .B2(n17914), .ZN(
        n17917) );
  OAI211_X1 U21016 ( .C1(n18203), .C2(n17918), .A(n17917), .B(n17916), .ZN(
        P3_U2835) );
  OAI222_X1 U21017 ( .A1(n17922), .A2(n17957), .B1(n17925), .B2(n17921), .C1(
        n17920), .C2(n17919), .ZN(n17923) );
  AOI22_X1 U21018 ( .A1(n9647), .A2(P3_REIP_REG_26__SCAN_IN), .B1(n18196), 
        .B2(n17923), .ZN(n17924) );
  OAI21_X1 U21019 ( .B1(n17925), .B2(n18203), .A(n17924), .ZN(P3_U2836) );
  AOI221_X1 U21020 ( .B1(n17927), .B2(n18723), .C1(n17950), .C2(n18723), .A(
        n17926), .ZN(n17932) );
  AOI21_X1 U21021 ( .B1(n17929), .B2(n17928), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17930) );
  AOI211_X1 U21022 ( .C1(n17932), .C2(n17931), .A(n17930), .B(n18218), .ZN(
        n17933) );
  AOI21_X1 U21023 ( .B1(n18186), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17933), .ZN(n17935) );
  OAI211_X1 U21024 ( .C1(n17936), .C2(n18137), .A(n17935), .B(n17934), .ZN(
        n17937) );
  AOI21_X1 U21025 ( .B1(n18134), .B2(n17938), .A(n17937), .ZN(n17939) );
  OAI21_X1 U21026 ( .B1(n18175), .B2(n17940), .A(n17939), .ZN(P3_U2837) );
  NOR2_X1 U21027 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17941), .ZN(
        n17944) );
  AOI21_X1 U21028 ( .B1(n17944), .B2(n17984), .A(n17943), .ZN(n17954) );
  INV_X1 U21029 ( .A(n17945), .ZN(n17949) );
  AOI22_X1 U21030 ( .A1(n18074), .A2(n17947), .B1(n18191), .B2(n17946), .ZN(
        n17948) );
  OAI211_X1 U21031 ( .C1(n17949), .C2(n18091), .A(n17948), .B(n18203), .ZN(
        n17952) );
  AOI211_X1 U21032 ( .C1(n18723), .C2(n17950), .A(n17956), .B(n17952), .ZN(
        n17951) );
  NOR2_X1 U21033 ( .A1(n9647), .A2(n17951), .ZN(n17959) );
  OAI211_X1 U21034 ( .C1(n18125), .C2(n17952), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17959), .ZN(n17953) );
  OAI211_X1 U21035 ( .C1(n17955), .C2(n18109), .A(n17954), .B(n17953), .ZN(
        P3_U2838) );
  OAI21_X1 U21036 ( .B1(n18186), .B2(n17957), .A(n17956), .ZN(n17958) );
  AOI22_X1 U21037 ( .A1(n18134), .A2(n17960), .B1(n17959), .B2(n17958), .ZN(
        n17962) );
  NAND2_X1 U21038 ( .A1(n17962), .A2(n17961), .ZN(P3_U2839) );
  AOI22_X1 U21039 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18196), .B1(
        n17963), .B2(n17984), .ZN(n17979) );
  AOI21_X1 U21040 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n18010), .A(
        n18188), .ZN(n17964) );
  AOI221_X1 U21041 ( .B1(n18009), .B2(n18219), .C1(n17994), .C2(n18219), .A(
        n17964), .ZN(n17992) );
  NAND2_X1 U21042 ( .A1(n18091), .A2(n18092), .ZN(n18095) );
  AOI22_X1 U21043 ( .A1(n18219), .A2(n17966), .B1(n17965), .B2(n18095), .ZN(
        n17967) );
  NAND2_X1 U21044 ( .A1(n17992), .A2(n17967), .ZN(n17980) );
  OAI22_X1 U21045 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18105), .B1(
        n17981), .B2(n18188), .ZN(n17973) );
  INV_X1 U21046 ( .A(n17968), .ZN(n17970) );
  NOR2_X1 U21047 ( .A1(n17969), .A2(n18092), .ZN(n18049) );
  AOI21_X1 U21048 ( .B1(n18722), .B2(n17970), .A(n18049), .ZN(n17993) );
  NAND2_X1 U21049 ( .A1(n17993), .A2(n17971), .ZN(n17972) );
  NOR4_X1 U21050 ( .A1(n17974), .A2(n17980), .A3(n17973), .A4(n17972), .ZN(
        n17978) );
  AOI22_X1 U21051 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18186), .B1(
        n18134), .B2(n17975), .ZN(n17977) );
  OAI211_X1 U21052 ( .C1(n17979), .C2(n17978), .A(n17977), .B(n17976), .ZN(
        P3_U2840) );
  NAND2_X1 U21053 ( .A1(n18196), .A2(n17993), .ZN(n18039) );
  AOI211_X1 U21054 ( .C1(n9640), .C2(n17990), .A(n18039), .B(n17980), .ZN(
        n17982) );
  AOI221_X1 U21055 ( .B1(n18202), .B2(n17982), .C1(n17981), .C2(n17982), .A(
        n9647), .ZN(n17986) );
  INV_X1 U21056 ( .A(n17983), .ZN(n17985) );
  NAND2_X1 U21057 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17984), .ZN(
        n18001) );
  INV_X1 U21058 ( .A(n18001), .ZN(n18003) );
  AOI22_X1 U21059 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17986), .B1(
        n17985), .B2(n18003), .ZN(n17988) );
  OAI211_X1 U21060 ( .C1(n17989), .C2(n18109), .A(n17988), .B(n17987), .ZN(
        P3_U2841) );
  NAND2_X1 U21061 ( .A1(n18008), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17996) );
  NAND2_X1 U21062 ( .A1(n9640), .A2(n17990), .ZN(n17991) );
  NAND4_X1 U21063 ( .A1(n17993), .A2(n17992), .A3(n18203), .A4(n17991), .ZN(
        n17995) );
  OAI221_X1 U21064 ( .B1(n17995), .B2(n17994), .C1(n17995), .C2(n18095), .A(
        n18217), .ZN(n18007) );
  OAI21_X1 U21065 ( .B1(n18202), .B2(n17996), .A(n18007), .ZN(n17998) );
  AOI22_X1 U21066 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17998), .B1(
        n18134), .B2(n17997), .ZN(n18000) );
  OAI211_X1 U21067 ( .C1(n18002), .C2(n18001), .A(n18000), .B(n17999), .ZN(
        P3_U2842) );
  AOI22_X1 U21068 ( .A1(n18134), .A2(n18004), .B1(n18003), .B2(n18008), .ZN(
        n18006) );
  NAND2_X1 U21069 ( .A1(n9647), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18005) );
  OAI211_X1 U21070 ( .C1(n18008), .C2(n18007), .A(n18006), .B(n18005), .ZN(
        P3_U2843) );
  NOR2_X1 U21071 ( .A1(n18701), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18189) );
  NOR3_X1 U21072 ( .A1(n18189), .A2(n18009), .A3(n18040), .ZN(n18014) );
  NOR2_X1 U21073 ( .A1(n18010), .A2(n18188), .ZN(n18011) );
  AOI211_X1 U21074 ( .C1(n18012), .C2(n18095), .A(n18011), .B(n18039), .ZN(
        n18013) );
  OAI21_X1 U21075 ( .B1(n18015), .B2(n18014), .A(n18013), .ZN(n18027) );
  OAI221_X1 U21076 ( .B1(n18027), .B2(n18016), .C1(n18027), .C2(n18191), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18025) );
  NAND2_X1 U21077 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18167) );
  INV_X1 U21078 ( .A(n18187), .ZN(n18017) );
  OAI22_X1 U21079 ( .A1(n18165), .A2(n18188), .B1(n18167), .B2(n18017), .ZN(
        n18121) );
  NAND2_X1 U21080 ( .A1(n18018), .A2(n18121), .ZN(n18141) );
  NOR2_X1 U21081 ( .A1(n18019), .A2(n18141), .ZN(n18045) );
  NOR2_X1 U21082 ( .A1(n18021), .A2(n18120), .ZN(n18041) );
  AOI22_X1 U21083 ( .A1(n18134), .A2(n18023), .B1(n18022), .B2(n18041), .ZN(
        n18024) );
  OAI221_X1 U21084 ( .B1(n9647), .B2(n18025), .C1(n18217), .C2(n18809), .A(
        n18024), .ZN(P3_U2844) );
  INV_X1 U21085 ( .A(n18041), .ZN(n18030) );
  AOI22_X1 U21086 ( .A1(n9647), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n18134), 
        .B2(n18026), .ZN(n18029) );
  NAND3_X1 U21087 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18217), .A3(
        n18027), .ZN(n18028) );
  OAI211_X1 U21088 ( .C1(n18031), .C2(n18030), .A(n18029), .B(n18028), .ZN(
        P3_U2845) );
  NOR2_X1 U21089 ( .A1(n9640), .A2(n18056), .ZN(n18037) );
  INV_X1 U21090 ( .A(n18032), .ZN(n18033) );
  AOI22_X1 U21091 ( .A1(n18723), .A2(n18034), .B1(n18219), .B2(n18033), .ZN(
        n18103) );
  AOI21_X1 U21092 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18058), .A(
        n18105), .ZN(n18035) );
  INV_X1 U21093 ( .A(n18035), .ZN(n18036) );
  OAI211_X1 U21094 ( .C1(n18038), .C2(n18037), .A(n18103), .B(n18036), .ZN(
        n18047) );
  OAI221_X1 U21095 ( .B1(n18039), .B2(n18125), .C1(n18039), .C2(n18047), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18044) );
  AOI22_X1 U21096 ( .A1(n18134), .A2(n18042), .B1(n18041), .B2(n18040), .ZN(
        n18043) );
  OAI221_X1 U21097 ( .B1(n9647), .B2(n18044), .C1(n18217), .C2(n18805), .A(
        n18043), .ZN(P3_U2846) );
  NAND2_X1 U21098 ( .A1(n18045), .A2(n18058), .ZN(n18061) );
  OAI21_X1 U21099 ( .B1(n18063), .B2(n18061), .A(n18056), .ZN(n18046) );
  AOI22_X1 U21100 ( .A1(n18049), .A2(n18048), .B1(n18047), .B2(n18046), .ZN(
        n18051) );
  OAI22_X1 U21101 ( .A1(n18051), .A2(n18218), .B1(n18109), .B2(n18050), .ZN(
        n18052) );
  AOI21_X1 U21102 ( .B1(n18214), .B2(n18053), .A(n18052), .ZN(n18055) );
  NAND2_X1 U21103 ( .A1(n9647), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18054) );
  OAI211_X1 U21104 ( .C1(n18203), .C2(n18056), .A(n18055), .B(n18054), .ZN(
        P3_U2847) );
  OAI21_X1 U21105 ( .B1(n18113), .B2(n18057), .A(n9640), .ZN(n18075) );
  OAI211_X1 U21106 ( .C1(n18059), .C2(n18058), .A(n18103), .B(n18075), .ZN(
        n18060) );
  OAI21_X1 U21107 ( .B1(n18063), .B2(n18060), .A(n18196), .ZN(n18062) );
  AOI222_X1 U21108 ( .A1(n18063), .A2(n18062), .B1(n18063), .B2(n18061), .C1(
        n18062), .C2(n18203), .ZN(n18064) );
  AOI21_X1 U21109 ( .B1(P3_REIP_REG_14__SCAN_IN), .B2(n9647), .A(n18064), .ZN(
        n18069) );
  INV_X1 U21110 ( .A(n18137), .ZN(n18066) );
  AOI22_X1 U21111 ( .A1(n18134), .A2(n18067), .B1(n18066), .B2(n18065), .ZN(
        n18068) );
  OAI211_X1 U21112 ( .C1(n18175), .C2(n18070), .A(n18069), .B(n18068), .ZN(
        P3_U2848) );
  AOI22_X1 U21113 ( .A1(n9647), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18134), 
        .B2(n18071), .ZN(n18080) );
  OAI21_X1 U21114 ( .B1(n18072), .B2(n18105), .A(n18103), .ZN(n18098) );
  AOI21_X1 U21115 ( .B1(n18074), .B2(n18073), .A(n18098), .ZN(n18076) );
  OAI211_X1 U21116 ( .C1(n18077), .C2(n18091), .A(n18076), .B(n18075), .ZN(
        n18085) );
  OAI21_X1 U21117 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18105), .A(
        n18196), .ZN(n18078) );
  OAI211_X1 U21118 ( .C1(n18085), .C2(n18078), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18217), .ZN(n18079) );
  OAI211_X1 U21119 ( .C1(n18120), .C2(n18081), .A(n18080), .B(n18079), .ZN(
        P3_U2849) );
  AOI22_X1 U21120 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18186), .B1(
        n9647), .B2(P3_REIP_REG_12__SCAN_IN), .ZN(n18087) );
  OAI22_X1 U21121 ( .A1(n18082), .A2(n18120), .B1(n18084), .B2(n18218), .ZN(
        n18083) );
  OAI21_X1 U21122 ( .B1(n18085), .B2(n18084), .A(n18083), .ZN(n18086) );
  OAI211_X1 U21123 ( .C1(n18088), .C2(n18109), .A(n18087), .B(n18086), .ZN(
        P3_U2850) );
  AOI22_X1 U21124 ( .A1(n9647), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18134), 
        .B2(n18089), .ZN(n18100) );
  OAI21_X1 U21125 ( .B1(n9943), .B2(n18113), .A(n9640), .ZN(n18090) );
  INV_X1 U21126 ( .A(n18090), .ZN(n18094) );
  OAI22_X1 U21127 ( .A1(n18093), .A2(n18092), .B1(n18091), .B2(n9804), .ZN(
        n18112) );
  AOI211_X1 U21128 ( .C1(n18096), .C2(n18095), .A(n18094), .B(n18112), .ZN(
        n18104) );
  OAI211_X1 U21129 ( .C1(n18701), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18196), .B(n18104), .ZN(n18097) );
  OAI211_X1 U21130 ( .C1(n18098), .C2(n18097), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18217), .ZN(n18099) );
  OAI211_X1 U21131 ( .C1(n18101), .C2(n18120), .A(n18100), .B(n18099), .ZN(
        P3_U2851) );
  NOR2_X1 U21132 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18120), .ZN(
        n18102) );
  AOI22_X1 U21133 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18102), .B1(
        n9647), .B2(P3_REIP_REG_10__SCAN_IN), .ZN(n18108) );
  NAND2_X1 U21134 ( .A1(n18196), .A2(n18103), .ZN(n18111) );
  OAI21_X1 U21135 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18105), .A(
        n18104), .ZN(n18106) );
  OAI211_X1 U21136 ( .C1(n18111), .C2(n18106), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n18217), .ZN(n18107) );
  OAI211_X1 U21137 ( .C1(n18110), .C2(n18109), .A(n18108), .B(n18107), .ZN(
        P3_U2852) );
  AOI211_X1 U21138 ( .C1(n9640), .C2(n18113), .A(n18112), .B(n18111), .ZN(
        n18115) );
  NOR3_X1 U21139 ( .A1(n9647), .A2(n18115), .A3(n9943), .ZN(n18116) );
  AOI21_X1 U21140 ( .B1(n18134), .B2(n18117), .A(n18116), .ZN(n18119) );
  OAI211_X1 U21141 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18120), .A(
        n18119), .B(n18118), .ZN(P3_U2853) );
  INV_X1 U21142 ( .A(n18121), .ZN(n18177) );
  INV_X1 U21143 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18184) );
  NOR3_X1 U21144 ( .A1(n18177), .A2(n18218), .A3(n18184), .ZN(n18172) );
  NAND3_X1 U21145 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n18172), .ZN(n18151) );
  NOR3_X1 U21146 ( .A1(n18142), .A2(n18150), .A3(n18151), .ZN(n18131) );
  OAI21_X1 U21147 ( .B1(n18189), .B2(n18122), .A(n18191), .ZN(n18123) );
  OAI21_X1 U21148 ( .B1(n18124), .B2(n18188), .A(n18123), .ZN(n18148) );
  AOI211_X1 U21149 ( .C1(n18125), .C2(n18150), .A(n18142), .B(n18148), .ZN(
        n18140) );
  INV_X1 U21150 ( .A(n18126), .ZN(n18204) );
  OAI21_X1 U21151 ( .B1(n18140), .B2(n18204), .A(n18203), .ZN(n18129) );
  INV_X1 U21152 ( .A(n18127), .ZN(n18128) );
  AOI221_X1 U21153 ( .B1(n18131), .B2(n18130), .C1(n18129), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18128), .ZN(n18136) );
  AOI22_X1 U21154 ( .A1(n18134), .A2(n18133), .B1(n18214), .B2(n18132), .ZN(
        n18135) );
  OAI211_X1 U21155 ( .C1(n18138), .C2(n18137), .A(n18136), .B(n18135), .ZN(
        P3_U2854) );
  AOI21_X1 U21156 ( .B1(n18186), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18139), .ZN(n18146) );
  AOI221_X1 U21157 ( .B1(n18150), .B2(n18142), .C1(n18141), .C2(n18142), .A(
        n18140), .ZN(n18144) );
  AOI22_X1 U21158 ( .A1(n18196), .A2(n18144), .B1(n18214), .B2(n18143), .ZN(
        n18145) );
  OAI211_X1 U21159 ( .C1(n18210), .C2(n18147), .A(n18146), .B(n18145), .ZN(
        P3_U2855) );
  AOI21_X1 U21160 ( .B1(n18196), .B2(n18148), .A(n18186), .ZN(n18157) );
  NAND2_X1 U21161 ( .A1(n9647), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n18149) );
  OAI221_X1 U21162 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18151), .C1(
        n18150), .C2(n18157), .A(n18149), .ZN(n18152) );
  AOI21_X1 U21163 ( .B1(n18214), .B2(n18153), .A(n18152), .ZN(n18154) );
  OAI21_X1 U21164 ( .B1(n18210), .B2(n18155), .A(n18154), .ZN(P3_U2856) );
  INV_X1 U21165 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18783) );
  NOR2_X1 U21166 ( .A1(n18217), .A2(n18783), .ZN(n18161) );
  INV_X1 U21167 ( .A(n18172), .ZN(n18156) );
  NOR2_X1 U21168 ( .A1(n18171), .A2(n18156), .ZN(n18159) );
  INV_X1 U21169 ( .A(n18157), .ZN(n18158) );
  MUX2_X1 U21170 ( .A(n18159), .B(n18158), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n18160) );
  AOI211_X1 U21171 ( .C1(n18214), .C2(n18162), .A(n18161), .B(n18160), .ZN(
        n18163) );
  OAI21_X1 U21172 ( .B1(n18210), .B2(n18164), .A(n18163), .ZN(P3_U2857) );
  NAND2_X1 U21173 ( .A1(n18723), .A2(n18165), .ZN(n18192) );
  NAND2_X1 U21174 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18192), .ZN(
        n18166) );
  AOI211_X1 U21175 ( .C1(n18167), .C2(n18191), .A(n18189), .B(n18166), .ZN(
        n18176) );
  OAI21_X1 U21176 ( .B1(n18176), .B2(n18204), .A(n18203), .ZN(n18170) );
  OAI22_X1 U21177 ( .A1(n18217), .A2(n18781), .B1(n18210), .B2(n18168), .ZN(
        n18169) );
  AOI221_X1 U21178 ( .B1(n18172), .B2(n18171), .C1(n18170), .C2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n18169), .ZN(n18173) );
  OAI21_X1 U21179 ( .B1(n18175), .B2(n18174), .A(n18173), .ZN(P3_U2858) );
  AOI211_X1 U21180 ( .C1(n18177), .C2(n18184), .A(n18176), .B(n18218), .ZN(
        n18181) );
  OAI21_X1 U21181 ( .B1(n18210), .B2(n18179), .A(n18178), .ZN(n18180) );
  AOI211_X1 U21182 ( .C1(n18182), .C2(n18214), .A(n18181), .B(n18180), .ZN(
        n18183) );
  OAI21_X1 U21183 ( .B1(n18184), .B2(n18203), .A(n18183), .ZN(P3_U2859) );
  AOI21_X1 U21184 ( .B1(n18186), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n18185), .ZN(n18200) );
  NAND2_X1 U21185 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18187), .ZN(
        n18195) );
  INV_X1 U21186 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18864) );
  NOR3_X1 U21187 ( .A1(n18188), .A2(n18884), .A3(n18864), .ZN(n18190) );
  AOI211_X1 U21188 ( .C1(n18864), .C2(n18191), .A(n18190), .B(n18189), .ZN(
        n18193) );
  OAI221_X1 U21189 ( .B1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n18195), .C1(
        n18194), .C2(n18193), .A(n18192), .ZN(n18198) );
  OAI221_X1 U21190 ( .B1(n18198), .B2(n18722), .C1(n18198), .C2(n18197), .A(
        n18196), .ZN(n18199) );
  OAI211_X1 U21191 ( .C1(n18201), .C2(n18210), .A(n18200), .B(n18199), .ZN(
        P3_U2860) );
  OR3_X1 U21192 ( .A1(n18218), .A2(n18202), .A3(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18221) );
  AOI21_X1 U21193 ( .B1(n18203), .B2(n18221), .A(n18864), .ZN(n18206) );
  AOI211_X1 U21194 ( .C1(n18703), .C2(n18884), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18204), .ZN(n18205) );
  AOI211_X1 U21195 ( .C1(n18214), .C2(n18207), .A(n18206), .B(n18205), .ZN(
        n18209) );
  NAND2_X1 U21196 ( .A1(n9647), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18208) );
  OAI211_X1 U21197 ( .C1(n18211), .C2(n18210), .A(n18209), .B(n18208), .ZN(
        P3_U2861) );
  AND2_X1 U21198 ( .A1(n9647), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18212) );
  AOI221_X1 U21199 ( .B1(n18216), .B2(n18215), .C1(n18214), .C2(n18213), .A(
        n18212), .ZN(n18222) );
  OAI211_X1 U21200 ( .C1(n18219), .C2(n18218), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n18217), .ZN(n18220) );
  NAND3_X1 U21201 ( .A1(n18222), .A2(n18221), .A3(n18220), .ZN(P3_U2862) );
  AOI211_X1 U21202 ( .C1(n18224), .C2(n18223), .A(n18749), .B(n18865), .ZN(
        n18742) );
  OAI21_X1 U21203 ( .B1(n18742), .B2(n18270), .A(n18229), .ZN(n18225) );
  OAI221_X1 U21204 ( .B1(n18707), .B2(n18900), .C1(n18707), .C2(n18229), .A(
        n18225), .ZN(P3_U2863) );
  NOR2_X1 U21205 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18717), .ZN(
        n18521) );
  NOR2_X1 U21206 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18714), .ZN(
        n18403) );
  NOR2_X1 U21207 ( .A1(n18521), .A2(n18403), .ZN(n18227) );
  OAI22_X1 U21208 ( .A1(n18228), .A2(n18717), .B1(n18227), .B2(n18226), .ZN(
        P3_U2866) );
  NOR2_X1 U21209 ( .A1(n18718), .A2(n18229), .ZN(P3_U2867) );
  NOR2_X1 U21210 ( .A1(n18714), .A2(n18717), .ZN(n18550) );
  INV_X1 U21211 ( .A(n18550), .ZN(n18231) );
  NOR2_X1 U21212 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18231), .ZN(
        n18627) );
  NAND2_X1 U21213 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18627), .ZN(
        n18663) );
  NAND2_X1 U21214 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18257), .ZN(n18631) );
  AND2_X1 U21215 ( .A1(n18257), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18624) );
  NAND2_X1 U21216 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18707), .ZN(
        n18376) );
  INV_X1 U21217 ( .A(n18376), .ZN(n18472) );
  NAND2_X1 U21218 ( .A1(n18550), .A2(n18472), .ZN(n18610) );
  INV_X1 U21219 ( .A(n18610), .ZN(n18617) );
  NOR2_X2 U21220 ( .A1(n18474), .A2(n18230), .ZN(n18623) );
  NOR2_X1 U21221 ( .A1(n18717), .A2(n18401), .ZN(n18626) );
  NAND2_X1 U21222 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18626), .ZN(
        n18309) );
  NAND2_X1 U21223 ( .A1(n18709), .A2(n18707), .ZN(n18710) );
  NAND2_X1 U21224 ( .A1(n18714), .A2(n18717), .ZN(n18310) );
  NOR2_X2 U21225 ( .A1(n18710), .A2(n18310), .ZN(n18325) );
  INV_X1 U21226 ( .A(n18325), .ZN(n18332) );
  NAND2_X1 U21227 ( .A1(n18309), .A2(n18332), .ZN(n18289) );
  AND2_X1 U21228 ( .A1(n18622), .A2(n18289), .ZN(n18264) );
  AOI22_X1 U21229 ( .A1(n18624), .A2(n18617), .B1(n18623), .B2(n18264), .ZN(
        n18236) );
  NOR2_X1 U21230 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18707), .ZN(
        n18447) );
  NOR2_X1 U21231 ( .A1(n18472), .A2(n18447), .ZN(n18523) );
  NOR2_X1 U21232 ( .A1(n18523), .A2(n18231), .ZN(n18586) );
  AOI21_X1 U21233 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18474), .ZN(n18583) );
  AOI22_X1 U21234 ( .A1(n18257), .A2(n18586), .B1(n18583), .B2(n18289), .ZN(
        n18267) );
  NAND2_X1 U21235 ( .A1(n18233), .A2(n18232), .ZN(n18265) );
  NOR2_X1 U21236 ( .A1(n18234), .A2(n18265), .ZN(n18628) );
  AOI22_X1 U21237 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18267), .B1(
        n18325), .B2(n18628), .ZN(n18235) );
  OAI211_X1 U21238 ( .C1(n18663), .C2(n18631), .A(n18236), .B(n18235), .ZN(
        P3_U2868) );
  NAND2_X1 U21239 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18257), .ZN(n18481) );
  NAND2_X1 U21240 ( .A1(n18257), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18637) );
  INV_X1 U21241 ( .A(n18637), .ZN(n18590) );
  AND2_X1 U21242 ( .A1(n18525), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18632) );
  AOI22_X1 U21243 ( .A1(n18617), .A2(n18590), .B1(n18264), .B2(n18632), .ZN(
        n18238) );
  NOR2_X2 U21244 ( .A1(n18906), .A2(n18265), .ZN(n18634) );
  AOI22_X1 U21245 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18267), .B1(
        n18325), .B2(n18634), .ZN(n18237) );
  OAI211_X1 U21246 ( .C1(n18663), .C2(n18481), .A(n18238), .B(n18237), .ZN(
        P3_U2869) );
  NAND2_X1 U21247 ( .A1(n18257), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18597) );
  INV_X1 U21248 ( .A(n18663), .ZN(n18673) );
  NOR2_X1 U21249 ( .A1(n18239), .A2(n18263), .ZN(n18594) );
  NOR2_X2 U21250 ( .A1(n18474), .A2(n18240), .ZN(n18638) );
  AOI22_X1 U21251 ( .A1(n18673), .A2(n18594), .B1(n18264), .B2(n18638), .ZN(
        n18243) );
  NOR2_X2 U21252 ( .A1(n18241), .A2(n18265), .ZN(n18640) );
  AOI22_X1 U21253 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18267), .B1(
        n18325), .B2(n18640), .ZN(n18242) );
  OAI211_X1 U21254 ( .C1(n18610), .C2(n18597), .A(n18243), .B(n18242), .ZN(
        P3_U2870) );
  NAND2_X1 U21255 ( .A1(n18257), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18534) );
  NAND2_X1 U21256 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18257), .ZN(n18649) );
  INV_X1 U21257 ( .A(n18649), .ZN(n18598) );
  NOR2_X2 U21258 ( .A1(n18474), .A2(n18244), .ZN(n18644) );
  AOI22_X1 U21259 ( .A1(n18673), .A2(n18598), .B1(n18264), .B2(n18644), .ZN(
        n18247) );
  NOR2_X2 U21260 ( .A1(n18245), .A2(n18265), .ZN(n18646) );
  AOI22_X1 U21261 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18267), .B1(
        n18325), .B2(n18646), .ZN(n18246) );
  OAI211_X1 U21262 ( .C1(n18610), .C2(n18534), .A(n18247), .B(n18246), .ZN(
        P3_U2871) );
  NAND2_X1 U21263 ( .A1(n18257), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18537) );
  NOR2_X1 U21264 ( .A1(n18248), .A2(n18263), .ZN(n18602) );
  NOR2_X2 U21265 ( .A1(n18474), .A2(n18249), .ZN(n18650) );
  AOI22_X1 U21266 ( .A1(n18673), .A2(n18602), .B1(n18264), .B2(n18650), .ZN(
        n18252) );
  NOR2_X2 U21267 ( .A1(n9677), .A2(n18265), .ZN(n18652) );
  AOI22_X1 U21268 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18267), .B1(
        n18325), .B2(n18652), .ZN(n18251) );
  OAI211_X1 U21269 ( .C1(n18610), .C2(n18537), .A(n18252), .B(n18251), .ZN(
        P3_U2872) );
  NAND2_X1 U21270 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n18257), .ZN(n18662) );
  NAND2_X1 U21271 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18257), .ZN(n18570) );
  INV_X1 U21272 ( .A(n18570), .ZN(n18658) );
  NOR2_X2 U21273 ( .A1(n18253), .A2(n18474), .ZN(n18656) );
  AOI22_X1 U21274 ( .A1(n18673), .A2(n18658), .B1(n18264), .B2(n18656), .ZN(
        n18256) );
  NOR2_X2 U21275 ( .A1(n18254), .A2(n18265), .ZN(n18659) );
  AOI22_X1 U21276 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18267), .B1(
        n18325), .B2(n18659), .ZN(n18255) );
  OAI211_X1 U21277 ( .C1(n18610), .C2(n18662), .A(n18256), .B(n18255), .ZN(
        P3_U2873) );
  NAND2_X1 U21278 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18257), .ZN(n18669) );
  NAND2_X1 U21279 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18257), .ZN(n18543) );
  INV_X1 U21280 ( .A(n18543), .ZN(n18665) );
  NOR2_X2 U21281 ( .A1(n18258), .A2(n18474), .ZN(n18664) );
  AOI22_X1 U21282 ( .A1(n18617), .A2(n18665), .B1(n18264), .B2(n18664), .ZN(
        n18261) );
  NOR2_X2 U21283 ( .A1(n18259), .A2(n18265), .ZN(n18666) );
  AOI22_X1 U21284 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18267), .B1(
        n18325), .B2(n18666), .ZN(n18260) );
  OAI211_X1 U21285 ( .C1(n18663), .C2(n18669), .A(n18261), .B(n18260), .ZN(
        P3_U2874) );
  NOR2_X1 U21286 ( .A1(n18263), .A2(n18262), .ZN(n18616) );
  INV_X1 U21287 ( .A(n18616), .ZN(n18680) );
  NAND2_X1 U21288 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18257), .ZN(n18621) );
  AND2_X1 U21289 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18525), .ZN(n18671) );
  AOI22_X1 U21290 ( .A1(n18617), .A2(n18672), .B1(n18264), .B2(n18671), .ZN(
        n18269) );
  NOR2_X2 U21291 ( .A1(n18266), .A2(n18265), .ZN(n18674) );
  AOI22_X1 U21292 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18267), .B1(
        n18325), .B2(n18674), .ZN(n18268) );
  OAI211_X1 U21293 ( .C1(n18663), .C2(n18680), .A(n18269), .B(n18268), .ZN(
        P3_U2875) );
  INV_X1 U21294 ( .A(n18309), .ZN(n18675) );
  NAND2_X1 U21295 ( .A1(n18709), .A2(n18622), .ZN(n18448) );
  NOR2_X1 U21296 ( .A1(n18310), .A2(n18448), .ZN(n18285) );
  AOI22_X1 U21297 ( .A1(n18675), .A2(n18624), .B1(n18623), .B2(n18285), .ZN(
        n18272) );
  INV_X1 U21298 ( .A(n18310), .ZN(n18312) );
  NOR2_X1 U21299 ( .A1(n18474), .A2(n18270), .ZN(n18625) );
  INV_X1 U21300 ( .A(n18625), .ZN(n18311) );
  NOR2_X1 U21301 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18311), .ZN(
        n18549) );
  AOI22_X1 U21302 ( .A1(n18257), .A2(n18626), .B1(n18312), .B2(n18549), .ZN(
        n18286) );
  NAND2_X1 U21303 ( .A1(n18447), .A2(n18312), .ZN(n18354) );
  INV_X1 U21304 ( .A(n18354), .ZN(n18347) );
  AOI22_X1 U21305 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18286), .B1(
        n18628), .B2(n18347), .ZN(n18271) );
  OAI211_X1 U21306 ( .C1(n18631), .C2(n18610), .A(n18272), .B(n18271), .ZN(
        P3_U2876) );
  AOI22_X1 U21307 ( .A1(n18617), .A2(n18633), .B1(n18632), .B2(n18285), .ZN(
        n18274) );
  AOI22_X1 U21308 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18286), .B1(
        n18634), .B2(n18347), .ZN(n18273) );
  OAI211_X1 U21309 ( .C1(n18309), .C2(n18637), .A(n18274), .B(n18273), .ZN(
        P3_U2877) );
  AOI22_X1 U21310 ( .A1(n18617), .A2(n18594), .B1(n18638), .B2(n18285), .ZN(
        n18276) );
  AOI22_X1 U21311 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18286), .B1(
        n18640), .B2(n18347), .ZN(n18275) );
  OAI211_X1 U21312 ( .C1(n18309), .C2(n18597), .A(n18276), .B(n18275), .ZN(
        P3_U2878) );
  AOI22_X1 U21313 ( .A1(n18617), .A2(n18598), .B1(n18644), .B2(n18285), .ZN(
        n18278) );
  AOI22_X1 U21314 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18286), .B1(
        n18646), .B2(n18347), .ZN(n18277) );
  OAI211_X1 U21315 ( .C1(n18309), .C2(n18534), .A(n18278), .B(n18277), .ZN(
        P3_U2879) );
  AOI22_X1 U21316 ( .A1(n18617), .A2(n18602), .B1(n18650), .B2(n18285), .ZN(
        n18280) );
  AOI22_X1 U21317 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18286), .B1(
        n18652), .B2(n18347), .ZN(n18279) );
  OAI211_X1 U21318 ( .C1(n18309), .C2(n18537), .A(n18280), .B(n18279), .ZN(
        P3_U2880) );
  INV_X1 U21319 ( .A(n18662), .ZN(n18606) );
  AOI22_X1 U21320 ( .A1(n18675), .A2(n18606), .B1(n18656), .B2(n18285), .ZN(
        n18282) );
  AOI22_X1 U21321 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18286), .B1(
        n18659), .B2(n18347), .ZN(n18281) );
  OAI211_X1 U21322 ( .C1(n18610), .C2(n18570), .A(n18282), .B(n18281), .ZN(
        P3_U2881) );
  INV_X1 U21323 ( .A(n18669), .ZN(n18571) );
  AOI22_X1 U21324 ( .A1(n18617), .A2(n18571), .B1(n18664), .B2(n18285), .ZN(
        n18284) );
  AOI22_X1 U21325 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18286), .B1(
        n18666), .B2(n18347), .ZN(n18283) );
  OAI211_X1 U21326 ( .C1(n18309), .C2(n18543), .A(n18284), .B(n18283), .ZN(
        P3_U2882) );
  AOI22_X1 U21327 ( .A1(n18675), .A2(n18672), .B1(n18671), .B2(n18285), .ZN(
        n18288) );
  AOI22_X1 U21328 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18286), .B1(
        n18674), .B2(n18347), .ZN(n18287) );
  OAI211_X1 U21329 ( .C1(n18610), .C2(n18680), .A(n18288), .B(n18287), .ZN(
        P3_U2883) );
  INV_X1 U21330 ( .A(n18628), .ZN(n18589) );
  NAND2_X1 U21331 ( .A1(n18472), .A2(n18312), .ZN(n18375) );
  INV_X1 U21332 ( .A(n18631), .ZN(n18581) );
  INV_X1 U21333 ( .A(n18375), .ZN(n18368) );
  NOR2_X1 U21334 ( .A1(n18347), .A2(n18368), .ZN(n18333) );
  NOR2_X1 U21335 ( .A1(n18750), .A2(n18333), .ZN(n18305) );
  AOI22_X1 U21336 ( .A1(n18581), .A2(n18675), .B1(n18623), .B2(n18305), .ZN(
        n18292) );
  INV_X1 U21337 ( .A(n18333), .ZN(n18290) );
  OAI221_X1 U21338 ( .B1(n18290), .B2(n18585), .C1(n18290), .C2(n18289), .A(
        n18583), .ZN(n18306) );
  AOI22_X1 U21339 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18306), .B1(
        n18325), .B2(n18624), .ZN(n18291) );
  OAI211_X1 U21340 ( .C1(n18589), .C2(n18375), .A(n18292), .B(n18291), .ZN(
        P3_U2884) );
  AOI22_X1 U21341 ( .A1(n18675), .A2(n18633), .B1(n18632), .B2(n18305), .ZN(
        n18294) );
  AOI22_X1 U21342 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18306), .B1(
        n18634), .B2(n18368), .ZN(n18293) );
  OAI211_X1 U21343 ( .C1(n18332), .C2(n18637), .A(n18294), .B(n18293), .ZN(
        P3_U2885) );
  AOI22_X1 U21344 ( .A1(n18675), .A2(n18594), .B1(n18638), .B2(n18305), .ZN(
        n18296) );
  AOI22_X1 U21345 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18306), .B1(
        n18640), .B2(n18368), .ZN(n18295) );
  OAI211_X1 U21346 ( .C1(n18332), .C2(n18597), .A(n18296), .B(n18295), .ZN(
        P3_U2886) );
  AOI22_X1 U21347 ( .A1(n18675), .A2(n18598), .B1(n18644), .B2(n18305), .ZN(
        n18298) );
  AOI22_X1 U21348 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18306), .B1(
        n18646), .B2(n18368), .ZN(n18297) );
  OAI211_X1 U21349 ( .C1(n18332), .C2(n18534), .A(n18298), .B(n18297), .ZN(
        P3_U2887) );
  AOI22_X1 U21350 ( .A1(n18675), .A2(n18602), .B1(n18650), .B2(n18305), .ZN(
        n18300) );
  AOI22_X1 U21351 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18306), .B1(
        n18652), .B2(n18368), .ZN(n18299) );
  OAI211_X1 U21352 ( .C1(n18332), .C2(n18537), .A(n18300), .B(n18299), .ZN(
        P3_U2888) );
  AOI22_X1 U21353 ( .A1(n18325), .A2(n18606), .B1(n18656), .B2(n18305), .ZN(
        n18302) );
  AOI22_X1 U21354 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18306), .B1(
        n18659), .B2(n18368), .ZN(n18301) );
  OAI211_X1 U21355 ( .C1(n18309), .C2(n18570), .A(n18302), .B(n18301), .ZN(
        P3_U2889) );
  AOI22_X1 U21356 ( .A1(n18675), .A2(n18571), .B1(n18664), .B2(n18305), .ZN(
        n18304) );
  AOI22_X1 U21357 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18306), .B1(
        n18666), .B2(n18368), .ZN(n18303) );
  OAI211_X1 U21358 ( .C1(n18332), .C2(n18543), .A(n18304), .B(n18303), .ZN(
        P3_U2890) );
  AOI22_X1 U21359 ( .A1(n18325), .A2(n18672), .B1(n18671), .B2(n18305), .ZN(
        n18308) );
  AOI22_X1 U21360 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18306), .B1(
        n18674), .B2(n18368), .ZN(n18307) );
  OAI211_X1 U21361 ( .C1(n18309), .C2(n18680), .A(n18308), .B(n18307), .ZN(
        P3_U2891) );
  NOR2_X1 U21362 ( .A1(n18709), .A2(n18310), .ZN(n18355) );
  AND2_X1 U21363 ( .A1(n18622), .A2(n18355), .ZN(n18328) );
  AOI22_X1 U21364 ( .A1(n18624), .A2(n18347), .B1(n18623), .B2(n18328), .ZN(
        n18314) );
  INV_X1 U21365 ( .A(n18585), .ZN(n18378) );
  AOI21_X1 U21366 ( .B1(n18709), .B2(n18378), .A(n18311), .ZN(n18402) );
  NAND2_X1 U21367 ( .A1(n18312), .A2(n18402), .ZN(n18329) );
  NAND2_X1 U21368 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18355), .ZN(
        n18400) );
  INV_X1 U21369 ( .A(n18400), .ZN(n18391) );
  AOI22_X1 U21370 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18329), .B1(
        n18628), .B2(n18391), .ZN(n18313) );
  OAI211_X1 U21371 ( .C1(n18631), .C2(n18332), .A(n18314), .B(n18313), .ZN(
        P3_U2892) );
  AOI22_X1 U21372 ( .A1(n18325), .A2(n18633), .B1(n18632), .B2(n18328), .ZN(
        n18316) );
  AOI22_X1 U21373 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18329), .B1(
        n18634), .B2(n18391), .ZN(n18315) );
  OAI211_X1 U21374 ( .C1(n18637), .C2(n18354), .A(n18316), .B(n18315), .ZN(
        P3_U2893) );
  AOI22_X1 U21375 ( .A1(n18325), .A2(n18594), .B1(n18638), .B2(n18328), .ZN(
        n18318) );
  AOI22_X1 U21376 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18329), .B1(
        n18640), .B2(n18391), .ZN(n18317) );
  OAI211_X1 U21377 ( .C1(n18597), .C2(n18354), .A(n18318), .B(n18317), .ZN(
        P3_U2894) );
  INV_X1 U21378 ( .A(n18534), .ZN(n18645) );
  AOI22_X1 U21379 ( .A1(n18645), .A2(n18347), .B1(n18644), .B2(n18328), .ZN(
        n18320) );
  AOI22_X1 U21380 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18329), .B1(
        n18646), .B2(n18391), .ZN(n18319) );
  OAI211_X1 U21381 ( .C1(n18332), .C2(n18649), .A(n18320), .B(n18319), .ZN(
        P3_U2895) );
  INV_X1 U21382 ( .A(n18602), .ZN(n18655) );
  INV_X1 U21383 ( .A(n18537), .ZN(n18651) );
  AOI22_X1 U21384 ( .A1(n18651), .A2(n18347), .B1(n18650), .B2(n18328), .ZN(
        n18322) );
  AOI22_X1 U21385 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18329), .B1(
        n18652), .B2(n18391), .ZN(n18321) );
  OAI211_X1 U21386 ( .C1(n18332), .C2(n18655), .A(n18322), .B(n18321), .ZN(
        P3_U2896) );
  AOI22_X1 U21387 ( .A1(n18325), .A2(n18658), .B1(n18656), .B2(n18328), .ZN(
        n18324) );
  AOI22_X1 U21388 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18329), .B1(
        n18659), .B2(n18391), .ZN(n18323) );
  OAI211_X1 U21389 ( .C1(n18662), .C2(n18354), .A(n18324), .B(n18323), .ZN(
        P3_U2897) );
  AOI22_X1 U21390 ( .A1(n18325), .A2(n18571), .B1(n18664), .B2(n18328), .ZN(
        n18327) );
  AOI22_X1 U21391 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18329), .B1(
        n18666), .B2(n18391), .ZN(n18326) );
  OAI211_X1 U21392 ( .C1(n18543), .C2(n18354), .A(n18327), .B(n18326), .ZN(
        P3_U2898) );
  AOI22_X1 U21393 ( .A1(n18672), .A2(n18347), .B1(n18671), .B2(n18328), .ZN(
        n18331) );
  AOI22_X1 U21394 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18329), .B1(
        n18674), .B2(n18391), .ZN(n18330) );
  OAI211_X1 U21395 ( .C1(n18332), .C2(n18680), .A(n18331), .B(n18330), .ZN(
        P3_U2899) );
  INV_X1 U21396 ( .A(n18710), .ZN(n18424) );
  NAND2_X1 U21397 ( .A1(n18424), .A2(n18403), .ZN(n18423) );
  INV_X1 U21398 ( .A(n18423), .ZN(n18416) );
  NOR2_X1 U21399 ( .A1(n18391), .A2(n18416), .ZN(n18379) );
  NOR2_X1 U21400 ( .A1(n18750), .A2(n18379), .ZN(n18350) );
  AOI22_X1 U21401 ( .A1(n18581), .A2(n18347), .B1(n18623), .B2(n18350), .ZN(
        n18336) );
  OAI21_X1 U21402 ( .B1(n18333), .B2(n18378), .A(n18379), .ZN(n18334) );
  OAI211_X1 U21403 ( .C1(n18416), .C2(n18854), .A(n18525), .B(n18334), .ZN(
        n18351) );
  AOI22_X1 U21404 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18351), .B1(
        n18624), .B2(n18368), .ZN(n18335) );
  OAI211_X1 U21405 ( .C1(n18589), .C2(n18423), .A(n18336), .B(n18335), .ZN(
        P3_U2900) );
  AOI22_X1 U21406 ( .A1(n18590), .A2(n18368), .B1(n18632), .B2(n18350), .ZN(
        n18338) );
  AOI22_X1 U21407 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18351), .B1(
        n18634), .B2(n18416), .ZN(n18337) );
  OAI211_X1 U21408 ( .C1(n18481), .C2(n18354), .A(n18338), .B(n18337), .ZN(
        P3_U2901) );
  INV_X1 U21409 ( .A(n18594), .ZN(n18643) );
  INV_X1 U21410 ( .A(n18597), .ZN(n18639) );
  AOI22_X1 U21411 ( .A1(n18639), .A2(n18368), .B1(n18638), .B2(n18350), .ZN(
        n18340) );
  AOI22_X1 U21412 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18351), .B1(
        n18640), .B2(n18416), .ZN(n18339) );
  OAI211_X1 U21413 ( .C1(n18643), .C2(n18354), .A(n18340), .B(n18339), .ZN(
        P3_U2902) );
  AOI22_X1 U21414 ( .A1(n18598), .A2(n18347), .B1(n18644), .B2(n18350), .ZN(
        n18342) );
  AOI22_X1 U21415 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18351), .B1(
        n18646), .B2(n18416), .ZN(n18341) );
  OAI211_X1 U21416 ( .C1(n18534), .C2(n18375), .A(n18342), .B(n18341), .ZN(
        P3_U2903) );
  AOI22_X1 U21417 ( .A1(n18651), .A2(n18368), .B1(n18650), .B2(n18350), .ZN(
        n18344) );
  AOI22_X1 U21418 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18351), .B1(
        n18652), .B2(n18416), .ZN(n18343) );
  OAI211_X1 U21419 ( .C1(n18655), .C2(n18354), .A(n18344), .B(n18343), .ZN(
        P3_U2904) );
  AOI22_X1 U21420 ( .A1(n18658), .A2(n18347), .B1(n18656), .B2(n18350), .ZN(
        n18346) );
  AOI22_X1 U21421 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18351), .B1(
        n18659), .B2(n18416), .ZN(n18345) );
  OAI211_X1 U21422 ( .C1(n18662), .C2(n18375), .A(n18346), .B(n18345), .ZN(
        P3_U2905) );
  AOI22_X1 U21423 ( .A1(n18571), .A2(n18347), .B1(n18664), .B2(n18350), .ZN(
        n18349) );
  AOI22_X1 U21424 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18351), .B1(
        n18666), .B2(n18416), .ZN(n18348) );
  OAI211_X1 U21425 ( .C1(n18543), .C2(n18375), .A(n18349), .B(n18348), .ZN(
        P3_U2906) );
  AOI22_X1 U21426 ( .A1(n18672), .A2(n18368), .B1(n18671), .B2(n18350), .ZN(
        n18353) );
  AOI22_X1 U21427 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18351), .B1(
        n18674), .B2(n18416), .ZN(n18352) );
  OAI211_X1 U21428 ( .C1(n18680), .C2(n18354), .A(n18353), .B(n18352), .ZN(
        P3_U2907) );
  NAND2_X1 U21429 ( .A1(n18403), .A2(n18447), .ZN(n18446) );
  INV_X1 U21430 ( .A(n18403), .ZN(n18377) );
  NOR2_X1 U21431 ( .A1(n18377), .A2(n18448), .ZN(n18371) );
  AOI22_X1 U21432 ( .A1(n18624), .A2(n18391), .B1(n18623), .B2(n18371), .ZN(
        n18357) );
  AOI22_X1 U21433 ( .A1(n18257), .A2(n18355), .B1(n18403), .B2(n18549), .ZN(
        n18372) );
  AOI22_X1 U21434 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18372), .B1(
        n18581), .B2(n18368), .ZN(n18356) );
  OAI211_X1 U21435 ( .C1(n18589), .C2(n18446), .A(n18357), .B(n18356), .ZN(
        P3_U2908) );
  INV_X1 U21436 ( .A(n18634), .ZN(n18593) );
  AOI22_X1 U21437 ( .A1(n18633), .A2(n18368), .B1(n18632), .B2(n18371), .ZN(
        n18359) );
  AOI22_X1 U21438 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18372), .B1(
        n18590), .B2(n18391), .ZN(n18358) );
  OAI211_X1 U21439 ( .C1(n18593), .C2(n18446), .A(n18359), .B(n18358), .ZN(
        P3_U2909) );
  AOI22_X1 U21440 ( .A1(n18639), .A2(n18391), .B1(n18638), .B2(n18371), .ZN(
        n18361) );
  INV_X1 U21441 ( .A(n18446), .ZN(n18429) );
  AOI22_X1 U21442 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18372), .B1(
        n18640), .B2(n18429), .ZN(n18360) );
  OAI211_X1 U21443 ( .C1(n18643), .C2(n18375), .A(n18361), .B(n18360), .ZN(
        P3_U2910) );
  AOI22_X1 U21444 ( .A1(n18598), .A2(n18368), .B1(n18644), .B2(n18371), .ZN(
        n18363) );
  AOI22_X1 U21445 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18372), .B1(
        n18646), .B2(n18429), .ZN(n18362) );
  OAI211_X1 U21446 ( .C1(n18534), .C2(n18400), .A(n18363), .B(n18362), .ZN(
        P3_U2911) );
  AOI22_X1 U21447 ( .A1(n18602), .A2(n18368), .B1(n18650), .B2(n18371), .ZN(
        n18365) );
  AOI22_X1 U21448 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18372), .B1(
        n18652), .B2(n18429), .ZN(n18364) );
  OAI211_X1 U21449 ( .C1(n18537), .C2(n18400), .A(n18365), .B(n18364), .ZN(
        P3_U2912) );
  AOI22_X1 U21450 ( .A1(n18606), .A2(n18391), .B1(n18656), .B2(n18371), .ZN(
        n18367) );
  AOI22_X1 U21451 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18372), .B1(
        n18659), .B2(n18429), .ZN(n18366) );
  OAI211_X1 U21452 ( .C1(n18570), .C2(n18375), .A(n18367), .B(n18366), .ZN(
        P3_U2913) );
  AOI22_X1 U21453 ( .A1(n18571), .A2(n18368), .B1(n18664), .B2(n18371), .ZN(
        n18370) );
  AOI22_X1 U21454 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18372), .B1(
        n18666), .B2(n18429), .ZN(n18369) );
  OAI211_X1 U21455 ( .C1(n18543), .C2(n18400), .A(n18370), .B(n18369), .ZN(
        P3_U2914) );
  AOI22_X1 U21456 ( .A1(n18672), .A2(n18391), .B1(n18671), .B2(n18371), .ZN(
        n18374) );
  AOI22_X1 U21457 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18372), .B1(
        n18674), .B2(n18429), .ZN(n18373) );
  OAI211_X1 U21458 ( .C1(n18680), .C2(n18375), .A(n18374), .B(n18373), .ZN(
        P3_U2915) );
  NOR2_X1 U21459 ( .A1(n18377), .A2(n18376), .ZN(n18461) );
  INV_X1 U21460 ( .A(n18461), .ZN(n18471) );
  NOR2_X1 U21461 ( .A1(n18429), .A2(n18464), .ZN(n18425) );
  NOR2_X1 U21462 ( .A1(n18750), .A2(n18425), .ZN(n18396) );
  AOI22_X1 U21463 ( .A1(n18624), .A2(n18416), .B1(n18623), .B2(n18396), .ZN(
        n18382) );
  OAI21_X1 U21464 ( .B1(n18379), .B2(n18378), .A(n18425), .ZN(n18380) );
  OAI211_X1 U21465 ( .C1(n18464), .C2(n18854), .A(n18525), .B(n18380), .ZN(
        n18397) );
  AOI22_X1 U21466 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18397), .B1(
        n18628), .B2(n18461), .ZN(n18381) );
  OAI211_X1 U21467 ( .C1(n18631), .C2(n18400), .A(n18382), .B(n18381), .ZN(
        P3_U2916) );
  AOI22_X1 U21468 ( .A1(n18633), .A2(n18391), .B1(n18632), .B2(n18396), .ZN(
        n18384) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18397), .B1(
        n18634), .B2(n18461), .ZN(n18383) );
  OAI211_X1 U21470 ( .C1(n18637), .C2(n18423), .A(n18384), .B(n18383), .ZN(
        P3_U2917) );
  AOI22_X1 U21471 ( .A1(n18639), .A2(n18416), .B1(n18638), .B2(n18396), .ZN(
        n18386) );
  AOI22_X1 U21472 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18397), .B1(
        n18640), .B2(n18464), .ZN(n18385) );
  OAI211_X1 U21473 ( .C1(n18643), .C2(n18400), .A(n18386), .B(n18385), .ZN(
        P3_U2918) );
  AOI22_X1 U21474 ( .A1(n18598), .A2(n18391), .B1(n18644), .B2(n18396), .ZN(
        n18388) );
  AOI22_X1 U21475 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18397), .B1(
        n18646), .B2(n18461), .ZN(n18387) );
  OAI211_X1 U21476 ( .C1(n18534), .C2(n18423), .A(n18388), .B(n18387), .ZN(
        P3_U2919) );
  AOI22_X1 U21477 ( .A1(n18651), .A2(n18416), .B1(n18650), .B2(n18396), .ZN(
        n18390) );
  AOI22_X1 U21478 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18397), .B1(
        n18652), .B2(n18461), .ZN(n18389) );
  OAI211_X1 U21479 ( .C1(n18655), .C2(n18400), .A(n18390), .B(n18389), .ZN(
        P3_U2920) );
  AOI22_X1 U21480 ( .A1(n18658), .A2(n18391), .B1(n18656), .B2(n18396), .ZN(
        n18393) );
  AOI22_X1 U21481 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18397), .B1(
        n18659), .B2(n18461), .ZN(n18392) );
  OAI211_X1 U21482 ( .C1(n18662), .C2(n18423), .A(n18393), .B(n18392), .ZN(
        P3_U2921) );
  AOI22_X1 U21483 ( .A1(n18664), .A2(n18396), .B1(n18665), .B2(n18416), .ZN(
        n18395) );
  AOI22_X1 U21484 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18397), .B1(
        n18666), .B2(n18464), .ZN(n18394) );
  OAI211_X1 U21485 ( .C1(n18669), .C2(n18400), .A(n18395), .B(n18394), .ZN(
        P3_U2922) );
  AOI22_X1 U21486 ( .A1(n18672), .A2(n18416), .B1(n18671), .B2(n18396), .ZN(
        n18399) );
  AOI22_X1 U21487 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18397), .B1(
        n18674), .B2(n18464), .ZN(n18398) );
  OAI211_X1 U21488 ( .C1(n18680), .C2(n18400), .A(n18399), .B(n18398), .ZN(
        P3_U2923) );
  NOR2_X1 U21489 ( .A1(n18401), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18449) );
  AND2_X1 U21490 ( .A1(n18622), .A2(n18449), .ZN(n18419) );
  AOI22_X1 U21491 ( .A1(n18624), .A2(n18429), .B1(n18623), .B2(n18419), .ZN(
        n18405) );
  NAND2_X1 U21492 ( .A1(n18403), .A2(n18402), .ZN(n18420) );
  NAND2_X1 U21493 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18449), .ZN(
        n18499) );
  INV_X1 U21494 ( .A(n18499), .ZN(n18490) );
  AOI22_X1 U21495 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18420), .B1(
        n18628), .B2(n18490), .ZN(n18404) );
  OAI211_X1 U21496 ( .C1(n18631), .C2(n18423), .A(n18405), .B(n18404), .ZN(
        P3_U2924) );
  AOI22_X1 U21497 ( .A1(n18633), .A2(n18416), .B1(n18632), .B2(n18419), .ZN(
        n18407) );
  AOI22_X1 U21498 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18420), .B1(
        n18634), .B2(n18490), .ZN(n18406) );
  OAI211_X1 U21499 ( .C1(n18637), .C2(n18446), .A(n18407), .B(n18406), .ZN(
        P3_U2925) );
  AOI22_X1 U21500 ( .A1(n18639), .A2(n18429), .B1(n18638), .B2(n18419), .ZN(
        n18409) );
  AOI22_X1 U21501 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18420), .B1(
        n18640), .B2(n18490), .ZN(n18408) );
  OAI211_X1 U21502 ( .C1(n18643), .C2(n18423), .A(n18409), .B(n18408), .ZN(
        P3_U2926) );
  AOI22_X1 U21503 ( .A1(n18645), .A2(n18429), .B1(n18644), .B2(n18419), .ZN(
        n18411) );
  AOI22_X1 U21504 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18420), .B1(
        n18646), .B2(n18490), .ZN(n18410) );
  OAI211_X1 U21505 ( .C1(n18649), .C2(n18423), .A(n18411), .B(n18410), .ZN(
        P3_U2927) );
  AOI22_X1 U21506 ( .A1(n18651), .A2(n18429), .B1(n18650), .B2(n18419), .ZN(
        n18413) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18420), .B1(
        n18652), .B2(n18490), .ZN(n18412) );
  OAI211_X1 U21508 ( .C1(n18655), .C2(n18423), .A(n18413), .B(n18412), .ZN(
        P3_U2928) );
  AOI22_X1 U21509 ( .A1(n18606), .A2(n18429), .B1(n18656), .B2(n18419), .ZN(
        n18415) );
  AOI22_X1 U21510 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18420), .B1(
        n18659), .B2(n18490), .ZN(n18414) );
  OAI211_X1 U21511 ( .C1(n18570), .C2(n18423), .A(n18415), .B(n18414), .ZN(
        P3_U2929) );
  AOI22_X1 U21512 ( .A1(n18571), .A2(n18416), .B1(n18664), .B2(n18419), .ZN(
        n18418) );
  AOI22_X1 U21513 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18420), .B1(
        n18666), .B2(n18490), .ZN(n18417) );
  OAI211_X1 U21514 ( .C1(n18543), .C2(n18446), .A(n18418), .B(n18417), .ZN(
        P3_U2930) );
  AOI22_X1 U21515 ( .A1(n18672), .A2(n18429), .B1(n18671), .B2(n18419), .ZN(
        n18422) );
  AOI22_X1 U21516 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18420), .B1(
        n18674), .B2(n18490), .ZN(n18421) );
  OAI211_X1 U21517 ( .C1(n18680), .C2(n18423), .A(n18422), .B(n18421), .ZN(
        P3_U2931) );
  NAND2_X1 U21518 ( .A1(n18424), .A2(n18521), .ZN(n18513) );
  NAND2_X1 U21519 ( .A1(n18499), .A2(n18513), .ZN(n18473) );
  INV_X1 U21520 ( .A(n18425), .ZN(n18426) );
  OAI221_X1 U21521 ( .B1(n18473), .B2(n18585), .C1(n18473), .C2(n18426), .A(
        n18583), .ZN(n18443) );
  AND2_X1 U21522 ( .A1(n18622), .A2(n18473), .ZN(n18442) );
  AOI22_X1 U21523 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18443), .B1(
        n18623), .B2(n18442), .ZN(n18428) );
  AOI22_X1 U21524 ( .A1(n18581), .A2(n18429), .B1(n18624), .B2(n18464), .ZN(
        n18427) );
  OAI211_X1 U21525 ( .C1(n18589), .C2(n18513), .A(n18428), .B(n18427), .ZN(
        P3_U2932) );
  AOI22_X1 U21526 ( .A1(n18633), .A2(n18429), .B1(n18632), .B2(n18442), .ZN(
        n18431) );
  AOI22_X1 U21527 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18443), .B1(
        n18590), .B2(n18464), .ZN(n18430) );
  OAI211_X1 U21528 ( .C1(n18593), .C2(n18513), .A(n18431), .B(n18430), .ZN(
        P3_U2933) );
  AOI22_X1 U21529 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18443), .B1(
        n18638), .B2(n18442), .ZN(n18433) );
  INV_X1 U21530 ( .A(n18513), .ZN(n18517) );
  AOI22_X1 U21531 ( .A1(n18639), .A2(n18464), .B1(n18640), .B2(n18517), .ZN(
        n18432) );
  OAI211_X1 U21532 ( .C1(n18643), .C2(n18446), .A(n18433), .B(n18432), .ZN(
        P3_U2934) );
  AOI22_X1 U21533 ( .A1(n18645), .A2(n18464), .B1(n18644), .B2(n18442), .ZN(
        n18435) );
  AOI22_X1 U21534 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18443), .B1(
        n18646), .B2(n18517), .ZN(n18434) );
  OAI211_X1 U21535 ( .C1(n18649), .C2(n18446), .A(n18435), .B(n18434), .ZN(
        P3_U2935) );
  AOI22_X1 U21536 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18443), .B1(
        n18650), .B2(n18442), .ZN(n18437) );
  AOI22_X1 U21537 ( .A1(n18651), .A2(n18464), .B1(n18652), .B2(n18517), .ZN(
        n18436) );
  OAI211_X1 U21538 ( .C1(n18655), .C2(n18446), .A(n18437), .B(n18436), .ZN(
        P3_U2936) );
  AOI22_X1 U21539 ( .A1(n18606), .A2(n18464), .B1(n18656), .B2(n18442), .ZN(
        n18439) );
  AOI22_X1 U21540 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18443), .B1(
        n18659), .B2(n18517), .ZN(n18438) );
  OAI211_X1 U21541 ( .C1(n18570), .C2(n18446), .A(n18439), .B(n18438), .ZN(
        P3_U2937) );
  AOI22_X1 U21542 ( .A1(n18664), .A2(n18442), .B1(n18665), .B2(n18461), .ZN(
        n18441) );
  AOI22_X1 U21543 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18443), .B1(
        n18666), .B2(n18517), .ZN(n18440) );
  OAI211_X1 U21544 ( .C1(n18669), .C2(n18446), .A(n18441), .B(n18440), .ZN(
        P3_U2938) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18443), .B1(
        n18671), .B2(n18442), .ZN(n18445) );
  AOI22_X1 U21546 ( .A1(n18674), .A2(n18517), .B1(n18672), .B2(n18464), .ZN(
        n18444) );
  OAI211_X1 U21547 ( .C1(n18680), .C2(n18446), .A(n18445), .B(n18444), .ZN(
        P3_U2939) );
  NAND2_X1 U21548 ( .A1(n18521), .A2(n18447), .ZN(n18548) );
  INV_X1 U21549 ( .A(n18521), .ZN(n18500) );
  NOR2_X1 U21550 ( .A1(n18500), .A2(n18448), .ZN(n18467) );
  AOI22_X1 U21551 ( .A1(n18581), .A2(n18464), .B1(n18623), .B2(n18467), .ZN(
        n18451) );
  AOI22_X1 U21552 ( .A1(n18257), .A2(n18449), .B1(n18521), .B2(n18549), .ZN(
        n18468) );
  AOI22_X1 U21553 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18468), .B1(
        n18624), .B2(n18490), .ZN(n18450) );
  OAI211_X1 U21554 ( .C1(n18589), .C2(n18548), .A(n18451), .B(n18450), .ZN(
        P3_U2940) );
  AOI22_X1 U21555 ( .A1(n18633), .A2(n18464), .B1(n18632), .B2(n18467), .ZN(
        n18453) );
  AOI22_X1 U21556 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18468), .B1(
        n18590), .B2(n18490), .ZN(n18452) );
  OAI211_X1 U21557 ( .C1(n18593), .C2(n18548), .A(n18453), .B(n18452), .ZN(
        P3_U2941) );
  INV_X1 U21558 ( .A(n18640), .ZN(n18456) );
  AOI22_X1 U21559 ( .A1(n18639), .A2(n18490), .B1(n18638), .B2(n18467), .ZN(
        n18455) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18468), .B1(
        n18594), .B2(n18461), .ZN(n18454) );
  OAI211_X1 U21561 ( .C1(n18456), .C2(n18548), .A(n18455), .B(n18454), .ZN(
        P3_U2942) );
  INV_X1 U21562 ( .A(n18646), .ZN(n18601) );
  AOI22_X1 U21563 ( .A1(n18645), .A2(n18490), .B1(n18644), .B2(n18467), .ZN(
        n18458) );
  AOI22_X1 U21564 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18468), .B1(
        n18598), .B2(n18461), .ZN(n18457) );
  OAI211_X1 U21565 ( .C1(n18601), .C2(n18548), .A(n18458), .B(n18457), .ZN(
        P3_U2943) );
  INV_X1 U21566 ( .A(n18652), .ZN(n18605) );
  AOI22_X1 U21567 ( .A1(n18651), .A2(n18490), .B1(n18650), .B2(n18467), .ZN(
        n18460) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18468), .B1(
        n18602), .B2(n18461), .ZN(n18459) );
  OAI211_X1 U21569 ( .C1(n18605), .C2(n18548), .A(n18460), .B(n18459), .ZN(
        P3_U2944) );
  INV_X1 U21570 ( .A(n18659), .ZN(n18609) );
  AOI22_X1 U21571 ( .A1(n18606), .A2(n18490), .B1(n18656), .B2(n18467), .ZN(
        n18463) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18468), .B1(
        n18658), .B2(n18461), .ZN(n18462) );
  OAI211_X1 U21573 ( .C1(n18609), .C2(n18548), .A(n18463), .B(n18462), .ZN(
        P3_U2945) );
  AOI22_X1 U21574 ( .A1(n18571), .A2(n18464), .B1(n18664), .B2(n18467), .ZN(
        n18466) );
  INV_X1 U21575 ( .A(n18548), .ZN(n18540) );
  AOI22_X1 U21576 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18468), .B1(
        n18666), .B2(n18540), .ZN(n18465) );
  OAI211_X1 U21577 ( .C1(n18543), .C2(n18499), .A(n18466), .B(n18465), .ZN(
        P3_U2946) );
  AOI22_X1 U21578 ( .A1(n18672), .A2(n18490), .B1(n18671), .B2(n18467), .ZN(
        n18470) );
  AOI22_X1 U21579 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18468), .B1(
        n18674), .B2(n18540), .ZN(n18469) );
  OAI211_X1 U21580 ( .C1(n18680), .C2(n18471), .A(n18470), .B(n18469), .ZN(
        P3_U2947) );
  NAND2_X1 U21581 ( .A1(n18521), .A2(n18472), .ZN(n18569) );
  INV_X1 U21582 ( .A(n18569), .ZN(n18576) );
  AOI211_X1 U21583 ( .C1(n18585), .C2(n18473), .A(n18540), .B(n18576), .ZN(
        n18475) );
  AOI211_X1 U21584 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(n18569), .A(n18475), 
        .B(n18474), .ZN(n18494) );
  AOI21_X1 U21585 ( .B1(n18548), .B2(n18569), .A(n18750), .ZN(n18495) );
  AOI22_X1 U21586 ( .A1(n18581), .A2(n18490), .B1(n18623), .B2(n18495), .ZN(
        n18477) );
  AOI22_X1 U21587 ( .A1(n18628), .A2(n18576), .B1(n18624), .B2(n18517), .ZN(
        n18476) );
  OAI211_X1 U21588 ( .C1(n18494), .C2(n18478), .A(n18477), .B(n18476), .ZN(
        P3_U2948) );
  AOI22_X1 U21589 ( .A1(n18590), .A2(n18517), .B1(n18632), .B2(n18495), .ZN(
        n18480) );
  INV_X1 U21590 ( .A(n18494), .ZN(n18496) );
  AOI22_X1 U21591 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18496), .B1(
        n18634), .B2(n18576), .ZN(n18479) );
  OAI211_X1 U21592 ( .C1(n18481), .C2(n18499), .A(n18480), .B(n18479), .ZN(
        P3_U2949) );
  AOI22_X1 U21593 ( .A1(n18639), .A2(n18517), .B1(n18638), .B2(n18495), .ZN(
        n18483) );
  AOI22_X1 U21594 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18496), .B1(
        n18640), .B2(n18576), .ZN(n18482) );
  OAI211_X1 U21595 ( .C1(n18643), .C2(n18499), .A(n18483), .B(n18482), .ZN(
        P3_U2950) );
  AOI22_X1 U21596 ( .A1(n18645), .A2(n18517), .B1(n18644), .B2(n18495), .ZN(
        n18485) );
  AOI22_X1 U21597 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18496), .B1(
        n18646), .B2(n18576), .ZN(n18484) );
  OAI211_X1 U21598 ( .C1(n18649), .C2(n18499), .A(n18485), .B(n18484), .ZN(
        P3_U2951) );
  AOI22_X1 U21599 ( .A1(n18602), .A2(n18490), .B1(n18650), .B2(n18495), .ZN(
        n18487) );
  AOI22_X1 U21600 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18496), .B1(
        n18652), .B2(n18576), .ZN(n18486) );
  OAI211_X1 U21601 ( .C1(n18537), .C2(n18513), .A(n18487), .B(n18486), .ZN(
        P3_U2952) );
  AOI22_X1 U21602 ( .A1(n18658), .A2(n18490), .B1(n18656), .B2(n18495), .ZN(
        n18489) );
  AOI22_X1 U21603 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18496), .B1(
        n18659), .B2(n18576), .ZN(n18488) );
  OAI211_X1 U21604 ( .C1(n18662), .C2(n18513), .A(n18489), .B(n18488), .ZN(
        P3_U2953) );
  AOI22_X1 U21605 ( .A1(n18571), .A2(n18490), .B1(n18664), .B2(n18495), .ZN(
        n18492) );
  AOI22_X1 U21606 ( .A1(n18666), .A2(n18576), .B1(n18665), .B2(n18517), .ZN(
        n18491) );
  OAI211_X1 U21607 ( .C1(n18494), .C2(n18493), .A(n18492), .B(n18491), .ZN(
        P3_U2954) );
  AOI22_X1 U21608 ( .A1(n18672), .A2(n18517), .B1(n18671), .B2(n18495), .ZN(
        n18498) );
  AOI22_X1 U21609 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18496), .B1(
        n18674), .B2(n18576), .ZN(n18497) );
  OAI211_X1 U21610 ( .C1(n18680), .C2(n18499), .A(n18498), .B(n18497), .ZN(
        P3_U2955) );
  NOR2_X1 U21611 ( .A1(n18709), .A2(n18500), .ZN(n18551) );
  AND2_X1 U21612 ( .A1(n18622), .A2(n18551), .ZN(n18516) );
  AOI22_X1 U21613 ( .A1(n18624), .A2(n18540), .B1(n18623), .B2(n18516), .ZN(
        n18502) );
  AOI22_X1 U21614 ( .A1(n18257), .A2(n18521), .B1(n18625), .B2(n18551), .ZN(
        n18518) );
  NAND2_X1 U21615 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18551), .ZN(
        n18613) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18518), .B1(
        n18628), .B2(n18615), .ZN(n18501) );
  OAI211_X1 U21617 ( .C1(n18631), .C2(n18513), .A(n18502), .B(n18501), .ZN(
        P3_U2956) );
  AOI22_X1 U21618 ( .A1(n18633), .A2(n18517), .B1(n18632), .B2(n18516), .ZN(
        n18504) );
  AOI22_X1 U21619 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18518), .B1(
        n18634), .B2(n18615), .ZN(n18503) );
  OAI211_X1 U21620 ( .C1(n18637), .C2(n18548), .A(n18504), .B(n18503), .ZN(
        P3_U2957) );
  AOI22_X1 U21621 ( .A1(n18594), .A2(n18517), .B1(n18638), .B2(n18516), .ZN(
        n18506) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18518), .B1(
        n18640), .B2(n18615), .ZN(n18505) );
  OAI211_X1 U21623 ( .C1(n18597), .C2(n18548), .A(n18506), .B(n18505), .ZN(
        P3_U2958) );
  AOI22_X1 U21624 ( .A1(n18598), .A2(n18517), .B1(n18644), .B2(n18516), .ZN(
        n18508) );
  AOI22_X1 U21625 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18518), .B1(
        n18646), .B2(n18615), .ZN(n18507) );
  OAI211_X1 U21626 ( .C1(n18534), .C2(n18548), .A(n18508), .B(n18507), .ZN(
        P3_U2959) );
  AOI22_X1 U21627 ( .A1(n18651), .A2(n18540), .B1(n18650), .B2(n18516), .ZN(
        n18510) );
  AOI22_X1 U21628 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18518), .B1(
        n18652), .B2(n18615), .ZN(n18509) );
  OAI211_X1 U21629 ( .C1(n18655), .C2(n18513), .A(n18510), .B(n18509), .ZN(
        P3_U2960) );
  AOI22_X1 U21630 ( .A1(n18606), .A2(n18540), .B1(n18656), .B2(n18516), .ZN(
        n18512) );
  AOI22_X1 U21631 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18518), .B1(
        n18659), .B2(n18615), .ZN(n18511) );
  OAI211_X1 U21632 ( .C1(n18570), .C2(n18513), .A(n18512), .B(n18511), .ZN(
        P3_U2961) );
  AOI22_X1 U21633 ( .A1(n18571), .A2(n18517), .B1(n18664), .B2(n18516), .ZN(
        n18515) );
  AOI22_X1 U21634 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18518), .B1(
        n18666), .B2(n18615), .ZN(n18514) );
  OAI211_X1 U21635 ( .C1(n18543), .C2(n18548), .A(n18515), .B(n18514), .ZN(
        P3_U2962) );
  AOI22_X1 U21636 ( .A1(n18616), .A2(n18517), .B1(n18671), .B2(n18516), .ZN(
        n18520) );
  AOI22_X1 U21637 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18518), .B1(
        n18674), .B2(n18615), .ZN(n18519) );
  OAI211_X1 U21638 ( .C1(n18621), .C2(n18548), .A(n18520), .B(n18519), .ZN(
        P3_U2963) );
  NAND2_X1 U21639 ( .A1(n18627), .A2(n18707), .ZN(n18679) );
  INV_X1 U21640 ( .A(n18679), .ZN(n18657) );
  NOR2_X1 U21641 ( .A1(n18615), .A2(n18657), .ZN(n18582) );
  NOR2_X1 U21642 ( .A1(n18750), .A2(n18582), .ZN(n18544) );
  AOI22_X1 U21643 ( .A1(n18624), .A2(n18576), .B1(n18623), .B2(n18544), .ZN(
        n18527) );
  NAND2_X1 U21644 ( .A1(n18585), .A2(n18521), .ZN(n18522) );
  OAI21_X1 U21645 ( .B1(n18523), .B2(n18522), .A(n18582), .ZN(n18524) );
  OAI211_X1 U21646 ( .C1(n18657), .C2(n18854), .A(n18525), .B(n18524), .ZN(
        n18545) );
  AOI22_X1 U21647 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18545), .B1(
        n18581), .B2(n18540), .ZN(n18526) );
  OAI211_X1 U21648 ( .C1(n18589), .C2(n18679), .A(n18527), .B(n18526), .ZN(
        P3_U2964) );
  AOI22_X1 U21649 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18545), .B1(
        n18632), .B2(n18544), .ZN(n18529) );
  AOI22_X1 U21650 ( .A1(n18633), .A2(n18540), .B1(n18634), .B2(n18657), .ZN(
        n18528) );
  OAI211_X1 U21651 ( .C1(n18637), .C2(n18569), .A(n18529), .B(n18528), .ZN(
        P3_U2965) );
  AOI22_X1 U21652 ( .A1(n18639), .A2(n18576), .B1(n18638), .B2(n18544), .ZN(
        n18531) );
  AOI22_X1 U21653 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18545), .B1(
        n18640), .B2(n18657), .ZN(n18530) );
  OAI211_X1 U21654 ( .C1(n18643), .C2(n18548), .A(n18531), .B(n18530), .ZN(
        P3_U2966) );
  AOI22_X1 U21655 ( .A1(n18598), .A2(n18540), .B1(n18644), .B2(n18544), .ZN(
        n18533) );
  AOI22_X1 U21656 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18545), .B1(
        n18646), .B2(n18657), .ZN(n18532) );
  OAI211_X1 U21657 ( .C1(n18534), .C2(n18569), .A(n18533), .B(n18532), .ZN(
        P3_U2967) );
  AOI22_X1 U21658 ( .A1(n18602), .A2(n18540), .B1(n18650), .B2(n18544), .ZN(
        n18536) );
  AOI22_X1 U21659 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18545), .B1(
        n18652), .B2(n18657), .ZN(n18535) );
  OAI211_X1 U21660 ( .C1(n18537), .C2(n18569), .A(n18536), .B(n18535), .ZN(
        P3_U2968) );
  AOI22_X1 U21661 ( .A1(n18658), .A2(n18540), .B1(n18656), .B2(n18544), .ZN(
        n18539) );
  AOI22_X1 U21662 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18545), .B1(
        n18659), .B2(n18657), .ZN(n18538) );
  OAI211_X1 U21663 ( .C1(n18662), .C2(n18569), .A(n18539), .B(n18538), .ZN(
        P3_U2969) );
  AOI22_X1 U21664 ( .A1(n18571), .A2(n18540), .B1(n18664), .B2(n18544), .ZN(
        n18542) );
  AOI22_X1 U21665 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18545), .B1(
        n18666), .B2(n18657), .ZN(n18541) );
  OAI211_X1 U21666 ( .C1(n18543), .C2(n18569), .A(n18542), .B(n18541), .ZN(
        P3_U2970) );
  AOI22_X1 U21667 ( .A1(n18672), .A2(n18576), .B1(n18671), .B2(n18544), .ZN(
        n18547) );
  AOI22_X1 U21668 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18545), .B1(
        n18674), .B2(n18657), .ZN(n18546) );
  OAI211_X1 U21669 ( .C1(n18680), .C2(n18548), .A(n18547), .B(n18546), .ZN(
        P3_U2971) );
  AOI22_X1 U21670 ( .A1(n18257), .A2(n18551), .B1(n18550), .B2(n18549), .ZN(
        n18566) );
  INV_X1 U21671 ( .A(n18566), .ZN(n18579) );
  AND2_X1 U21672 ( .A1(n18622), .A2(n18627), .ZN(n18575) );
  AOI22_X1 U21673 ( .A1(n18624), .A2(n18615), .B1(n18623), .B2(n18575), .ZN(
        n18553) );
  AOI22_X1 U21674 ( .A1(n18673), .A2(n18628), .B1(n18581), .B2(n18576), .ZN(
        n18552) );
  OAI211_X1 U21675 ( .C1(n18554), .C2(n18579), .A(n18553), .B(n18552), .ZN(
        P3_U2972) );
  AOI22_X1 U21676 ( .A1(n18590), .A2(n18615), .B1(n18632), .B2(n18575), .ZN(
        n18556) );
  AOI22_X1 U21677 ( .A1(n18673), .A2(n18634), .B1(n18633), .B2(n18576), .ZN(
        n18555) );
  OAI211_X1 U21678 ( .C1(n18557), .C2(n18579), .A(n18556), .B(n18555), .ZN(
        P3_U2973) );
  AOI22_X1 U21679 ( .A1(n18594), .A2(n18576), .B1(n18638), .B2(n18575), .ZN(
        n18559) );
  AOI22_X1 U21680 ( .A1(n18673), .A2(n18640), .B1(n18639), .B2(n18615), .ZN(
        n18558) );
  OAI211_X1 U21681 ( .C1(n18560), .C2(n18579), .A(n18559), .B(n18558), .ZN(
        P3_U2974) );
  AOI22_X1 U21682 ( .A1(n18645), .A2(n18615), .B1(n18644), .B2(n18575), .ZN(
        n18562) );
  AOI22_X1 U21683 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18566), .B1(
        n18673), .B2(n18646), .ZN(n18561) );
  OAI211_X1 U21684 ( .C1(n18649), .C2(n18569), .A(n18562), .B(n18561), .ZN(
        P3_U2975) );
  AOI22_X1 U21685 ( .A1(n18651), .A2(n18615), .B1(n18650), .B2(n18575), .ZN(
        n18564) );
  AOI22_X1 U21686 ( .A1(n18673), .A2(n18652), .B1(n18602), .B2(n18576), .ZN(
        n18563) );
  OAI211_X1 U21687 ( .C1(n18565), .C2(n18579), .A(n18564), .B(n18563), .ZN(
        P3_U2976) );
  AOI22_X1 U21688 ( .A1(n18606), .A2(n18615), .B1(n18656), .B2(n18575), .ZN(
        n18568) );
  AOI22_X1 U21689 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18566), .B1(
        n18673), .B2(n18659), .ZN(n18567) );
  OAI211_X1 U21690 ( .C1(n18570), .C2(n18569), .A(n18568), .B(n18567), .ZN(
        P3_U2977) );
  AOI22_X1 U21691 ( .A1(n18664), .A2(n18575), .B1(n18665), .B2(n18615), .ZN(
        n18573) );
  AOI22_X1 U21692 ( .A1(n18673), .A2(n18666), .B1(n18571), .B2(n18576), .ZN(
        n18572) );
  OAI211_X1 U21693 ( .C1(n18574), .C2(n18579), .A(n18573), .B(n18572), .ZN(
        P3_U2978) );
  AOI22_X1 U21694 ( .A1(n18672), .A2(n18615), .B1(n18671), .B2(n18575), .ZN(
        n18578) );
  AOI22_X1 U21695 ( .A1(n18673), .A2(n18674), .B1(n18616), .B2(n18576), .ZN(
        n18577) );
  OAI211_X1 U21696 ( .C1(n18580), .C2(n18579), .A(n18578), .B(n18577), .ZN(
        P3_U2979) );
  AND2_X1 U21697 ( .A1(n18622), .A2(n18586), .ZN(n18614) );
  AOI22_X1 U21698 ( .A1(n18581), .A2(n18615), .B1(n18623), .B2(n18614), .ZN(
        n18588) );
  INV_X1 U21699 ( .A(n18582), .ZN(n18584) );
  OAI221_X1 U21700 ( .B1(n18586), .B2(n18585), .C1(n18586), .C2(n18584), .A(
        n18583), .ZN(n18618) );
  AOI22_X1 U21701 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18618), .B1(
        n18624), .B2(n18657), .ZN(n18587) );
  OAI211_X1 U21702 ( .C1(n18589), .C2(n18610), .A(n18588), .B(n18587), .ZN(
        P3_U2980) );
  AOI22_X1 U21703 ( .A1(n18590), .A2(n18657), .B1(n18632), .B2(n18614), .ZN(
        n18592) );
  AOI22_X1 U21704 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18618), .B1(
        n18633), .B2(n18615), .ZN(n18591) );
  OAI211_X1 U21705 ( .C1(n18610), .C2(n18593), .A(n18592), .B(n18591), .ZN(
        P3_U2981) );
  AOI22_X1 U21706 ( .A1(n18594), .A2(n18615), .B1(n18638), .B2(n18614), .ZN(
        n18596) );
  AOI22_X1 U21707 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18618), .B1(
        n18617), .B2(n18640), .ZN(n18595) );
  OAI211_X1 U21708 ( .C1(n18597), .C2(n18679), .A(n18596), .B(n18595), .ZN(
        P3_U2982) );
  AOI22_X1 U21709 ( .A1(n18645), .A2(n18657), .B1(n18644), .B2(n18614), .ZN(
        n18600) );
  AOI22_X1 U21710 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18618), .B1(
        n18598), .B2(n18615), .ZN(n18599) );
  OAI211_X1 U21711 ( .C1(n18610), .C2(n18601), .A(n18600), .B(n18599), .ZN(
        P3_U2983) );
  AOI22_X1 U21712 ( .A1(n18651), .A2(n18657), .B1(n18650), .B2(n18614), .ZN(
        n18604) );
  AOI22_X1 U21713 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18618), .B1(
        n18602), .B2(n18615), .ZN(n18603) );
  OAI211_X1 U21714 ( .C1(n18610), .C2(n18605), .A(n18604), .B(n18603), .ZN(
        P3_U2984) );
  AOI22_X1 U21715 ( .A1(n18606), .A2(n18657), .B1(n18656), .B2(n18614), .ZN(
        n18608) );
  AOI22_X1 U21716 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18618), .B1(
        n18658), .B2(n18615), .ZN(n18607) );
  OAI211_X1 U21717 ( .C1(n18610), .C2(n18609), .A(n18608), .B(n18607), .ZN(
        P3_U2985) );
  AOI22_X1 U21718 ( .A1(n18664), .A2(n18614), .B1(n18665), .B2(n18657), .ZN(
        n18612) );
  AOI22_X1 U21719 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18618), .B1(
        n18617), .B2(n18666), .ZN(n18611) );
  OAI211_X1 U21720 ( .C1(n18669), .C2(n18613), .A(n18612), .B(n18611), .ZN(
        P3_U2986) );
  AOI22_X1 U21721 ( .A1(n18616), .A2(n18615), .B1(n18671), .B2(n18614), .ZN(
        n18620) );
  AOI22_X1 U21722 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18618), .B1(
        n18617), .B2(n18674), .ZN(n18619) );
  OAI211_X1 U21723 ( .C1(n18621), .C2(n18679), .A(n18620), .B(n18619), .ZN(
        P3_U2987) );
  AND2_X1 U21724 ( .A1(n18622), .A2(n18626), .ZN(n18670) );
  AOI22_X1 U21725 ( .A1(n18673), .A2(n18624), .B1(n18623), .B2(n18670), .ZN(
        n18630) );
  AOI22_X1 U21726 ( .A1(n18257), .A2(n18627), .B1(n18626), .B2(n18625), .ZN(
        n18676) );
  AOI22_X1 U21727 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18676), .B1(
        n18675), .B2(n18628), .ZN(n18629) );
  OAI211_X1 U21728 ( .C1(n18631), .C2(n18679), .A(n18630), .B(n18629), .ZN(
        P3_U2988) );
  AOI22_X1 U21729 ( .A1(n18633), .A2(n18657), .B1(n18632), .B2(n18670), .ZN(
        n18636) );
  AOI22_X1 U21730 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18676), .B1(
        n18675), .B2(n18634), .ZN(n18635) );
  OAI211_X1 U21731 ( .C1(n18663), .C2(n18637), .A(n18636), .B(n18635), .ZN(
        P3_U2989) );
  AOI22_X1 U21732 ( .A1(n18673), .A2(n18639), .B1(n18638), .B2(n18670), .ZN(
        n18642) );
  AOI22_X1 U21733 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18676), .B1(
        n18675), .B2(n18640), .ZN(n18641) );
  OAI211_X1 U21734 ( .C1(n18643), .C2(n18679), .A(n18642), .B(n18641), .ZN(
        P3_U2990) );
  AOI22_X1 U21735 ( .A1(n18673), .A2(n18645), .B1(n18644), .B2(n18670), .ZN(
        n18648) );
  AOI22_X1 U21736 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18676), .B1(
        n18675), .B2(n18646), .ZN(n18647) );
  OAI211_X1 U21737 ( .C1(n18649), .C2(n18679), .A(n18648), .B(n18647), .ZN(
        P3_U2991) );
  AOI22_X1 U21738 ( .A1(n18673), .A2(n18651), .B1(n18650), .B2(n18670), .ZN(
        n18654) );
  AOI22_X1 U21739 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18676), .B1(
        n18675), .B2(n18652), .ZN(n18653) );
  OAI211_X1 U21740 ( .C1(n18655), .C2(n18679), .A(n18654), .B(n18653), .ZN(
        P3_U2992) );
  AOI22_X1 U21741 ( .A1(n18658), .A2(n18657), .B1(n18656), .B2(n18670), .ZN(
        n18661) );
  AOI22_X1 U21742 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18676), .B1(
        n18675), .B2(n18659), .ZN(n18660) );
  OAI211_X1 U21743 ( .C1(n18663), .C2(n18662), .A(n18661), .B(n18660), .ZN(
        P3_U2993) );
  AOI22_X1 U21744 ( .A1(n18673), .A2(n18665), .B1(n18664), .B2(n18670), .ZN(
        n18668) );
  AOI22_X1 U21745 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18676), .B1(
        n18675), .B2(n18666), .ZN(n18667) );
  OAI211_X1 U21746 ( .C1(n18669), .C2(n18679), .A(n18668), .B(n18667), .ZN(
        P3_U2994) );
  AOI22_X1 U21747 ( .A1(n18673), .A2(n18672), .B1(n18671), .B2(n18670), .ZN(
        n18678) );
  AOI22_X1 U21748 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18676), .B1(
        n18675), .B2(n18674), .ZN(n18677) );
  OAI211_X1 U21749 ( .C1(n18680), .C2(n18679), .A(n18678), .B(n18677), .ZN(
        P3_U2995) );
  NAND2_X1 U21750 ( .A1(n18703), .A2(n18887), .ZN(n18704) );
  AOI22_X1 U21751 ( .A1(n18691), .A2(n18704), .B1(n18723), .B2(n18684), .ZN(
        n18855) );
  NOR2_X1 U21752 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18855), .ZN(
        n18688) );
  OAI21_X1 U21753 ( .B1(n18683), .B2(n18682), .A(n18681), .ZN(n18689) );
  OAI21_X1 U21754 ( .B1(n18691), .B2(n18703), .A(n18684), .ZN(n18685) );
  AOI21_X1 U21755 ( .B1(n18686), .B2(n18689), .A(n18685), .ZN(n18858) );
  NAND2_X1 U21756 ( .A1(n18734), .A2(n18858), .ZN(n18687) );
  AOI22_X1 U21757 ( .A1(n18734), .A2(n18688), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18687), .ZN(n18719) );
  INV_X1 U21758 ( .A(n18734), .ZN(n18712) );
  AOI21_X1 U21759 ( .B1(n18880), .B2(n18694), .A(n18689), .ZN(n18699) );
  NAND2_X1 U21760 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18690), .ZN(
        n18698) );
  AOI211_X1 U21761 ( .C1(n18880), .C2(n18872), .A(n18692), .B(n18691), .ZN(
        n18693) );
  INV_X1 U21762 ( .A(n18693), .ZN(n18697) );
  NOR2_X1 U21763 ( .A1(n18701), .A2(n18887), .ZN(n18695) );
  OAI211_X1 U21764 ( .C1(n18695), .C2(n18694), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n18872), .ZN(n18696) );
  OAI211_X1 U21765 ( .C1(n18699), .C2(n18698), .A(n18697), .B(n18696), .ZN(
        n18700) );
  AOI21_X1 U21766 ( .B1(n18723), .B2(n18866), .A(n18700), .ZN(n18869) );
  AOI22_X1 U21767 ( .A1(n18712), .A2(n18872), .B1(n18869), .B2(n18734), .ZN(
        n18716) );
  AND2_X1 U21768 ( .A1(n18702), .A2(n18701), .ZN(n18706) );
  AOI22_X1 U21769 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18703), .B1(
        n18706), .B2(n18887), .ZN(n18882) );
  INV_X1 U21770 ( .A(n18704), .ZN(n18705) );
  OAI22_X1 U21771 ( .A1(n18706), .A2(n18873), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18705), .ZN(n18878) );
  OR3_X1 U21772 ( .A1(n18882), .A2(n18709), .A3(n18707), .ZN(n18708) );
  AOI22_X1 U21773 ( .A1(n18882), .A2(n18709), .B1(n18878), .B2(n18708), .ZN(
        n18711) );
  OAI21_X1 U21774 ( .B1(n18712), .B2(n18711), .A(n18710), .ZN(n18713) );
  AOI222_X1 U21775 ( .A1(n18714), .A2(n18716), .B1(n18714), .B2(n18713), .C1(
        n18716), .C2(n18713), .ZN(n18715) );
  AOI211_X1 U21776 ( .C1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n18719), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n18715), .ZN(n18738) );
  INV_X1 U21777 ( .A(n18716), .ZN(n18721) );
  NAND2_X1 U21778 ( .A1(n18718), .A2(n18717), .ZN(n18720) );
  AOI21_X1 U21779 ( .B1(n18721), .B2(n18720), .A(n18719), .ZN(n18737) );
  NOR2_X1 U21780 ( .A1(n18723), .A2(n18722), .ZN(n18726) );
  OAI222_X1 U21781 ( .A1(n18729), .A2(n18728), .B1(n18727), .B2(n18726), .C1(
        n18725), .C2(n18724), .ZN(n18899) );
  AOI221_X1 U21782 ( .B1(P3_MORE_REG_SCAN_IN), .B2(n18731), .C1(
        P3_FLUSH_REG_SCAN_IN), .C2(n18731), .A(n18730), .ZN(n18732) );
  OAI211_X1 U21783 ( .C1(n18735), .C2(n18734), .A(n18733), .B(n18732), .ZN(
        n18736) );
  NOR4_X1 U21784 ( .A1(n18738), .A2(n18737), .A3(n18899), .A4(n18736), .ZN(
        n18748) );
  NOR2_X1 U21785 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18909) );
  AOI22_X1 U21786 ( .A1(n18881), .A2(n18909), .B1(n18766), .B2(n18903), .ZN(
        n18739) );
  INV_X1 U21787 ( .A(n18739), .ZN(n18744) );
  OAI211_X1 U21788 ( .C1(n18741), .C2(n18740), .A(n18901), .B(n18748), .ZN(
        n18853) );
  OAI21_X1 U21789 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18907), .A(n18853), 
        .ZN(n18751) );
  NOR2_X1 U21790 ( .A1(n18742), .A2(n18751), .ZN(n18743) );
  MUX2_X1 U21791 ( .A(n18744), .B(n18743), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18746) );
  OAI211_X1 U21792 ( .C1(n18748), .C2(n18747), .A(n18746), .B(n18745), .ZN(
        P3_U2996) );
  NAND2_X1 U21793 ( .A1(n18766), .A2(n18903), .ZN(n18754) );
  NAND4_X1 U21794 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n18766), .A4(n18749), .ZN(n18756) );
  OR3_X1 U21795 ( .A1(n18752), .A2(n18751), .A3(n18750), .ZN(n18753) );
  NAND4_X1 U21796 ( .A1(n18755), .A2(n18754), .A3(n18756), .A4(n18753), .ZN(
        P3_U2997) );
  INV_X1 U21797 ( .A(n18909), .ZN(n18758) );
  AND4_X1 U21798 ( .A1(n18758), .A2(n18757), .A3(n18756), .A4(n18852), .ZN(
        P3_U2998) );
  AND2_X1 U21799 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n9632), .ZN(P3_U2999) );
  AND2_X1 U21800 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n9631), .ZN(P3_U3000) );
  AND2_X1 U21801 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n9632), .ZN(P3_U3001) );
  AND2_X1 U21802 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n9631), .ZN(P3_U3002) );
  AND2_X1 U21803 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n9632), .ZN(P3_U3003) );
  AND2_X1 U21804 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n9631), .ZN(P3_U3004) );
  AND2_X1 U21805 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n9632), .ZN(P3_U3005) );
  AND2_X1 U21806 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n9631), .ZN(P3_U3006) );
  AND2_X1 U21807 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n9631), .ZN(P3_U3007) );
  AND2_X1 U21808 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n9632), .ZN(P3_U3008) );
  AND2_X1 U21809 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n9631), .ZN(P3_U3009) );
  AND2_X1 U21810 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n9632), .ZN(P3_U3010) );
  AND2_X1 U21811 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n9631), .ZN(P3_U3011) );
  AND2_X1 U21812 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n9632), .ZN(P3_U3012) );
  AND2_X1 U21813 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n9631), .ZN(P3_U3013) );
  AND2_X1 U21814 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n9632), .ZN(P3_U3014) );
  AND2_X1 U21815 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n9631), .ZN(P3_U3015) );
  AND2_X1 U21816 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n9632), .ZN(P3_U3016) );
  AND2_X1 U21817 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n9632), .ZN(P3_U3017) );
  AND2_X1 U21818 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n9631), .ZN(P3_U3018) );
  AND2_X1 U21819 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n9632), .ZN(P3_U3019) );
  AND2_X1 U21820 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n9631), .ZN(P3_U3020) );
  AND2_X1 U21821 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n9631), .ZN(P3_U3021)
         );
  AND2_X1 U21822 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n9632), .ZN(P3_U3022)
         );
  AND2_X1 U21823 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n9631), .ZN(P3_U3023)
         );
  AND2_X1 U21824 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n9632), .ZN(P3_U3024)
         );
  AND2_X1 U21825 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n9631), .ZN(P3_U3025)
         );
  AND2_X1 U21826 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n9632), .ZN(P3_U3026)
         );
  AND2_X1 U21827 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n9631), .ZN(P3_U3027)
         );
  AND2_X1 U21828 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n9632), .ZN(P3_U3028)
         );
  AOI21_X1 U21829 ( .B1(n18766), .B2(P3_STATE_REG_1__SCAN_IN), .A(n18771), 
        .ZN(n18772) );
  OAI21_X1 U21830 ( .B1(n18760), .B2(n21032), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18761) );
  INV_X1 U21831 ( .A(NA), .ZN(n20957) );
  NOR3_X1 U21832 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .A3(n20957), .ZN(n18773) );
  AOI21_X1 U21833 ( .B1(n18896), .B2(n18761), .A(n18773), .ZN(n18762) );
  OAI21_X1 U21834 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n18772), .A(n18762), 
        .ZN(P3_U3029) );
  AOI21_X1 U21835 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(HOLD), .A(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18763) );
  AOI21_X1 U21836 ( .B1(HOLD), .B2(P3_STATE_REG_2__SCAN_IN), .A(n18763), .ZN(
        n18764) );
  AOI22_X1 U21837 ( .A1(n18766), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n18764), .ZN(n18765) );
  NAND2_X1 U21838 ( .A1(n18765), .A2(n18904), .ZN(P3_U3030) );
  NOR2_X1 U21839 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(HOLD), .ZN(n18770)
         );
  NAND2_X1 U21840 ( .A1(n18766), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18767) );
  OAI22_X1 U21841 ( .A1(NA), .A2(n18767), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18768) );
  AOI21_X1 U21842 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(HOLD), .A(n18768), .ZN(
        n18769) );
  OAI33_X1 U21843 ( .A1(n18774), .A2(n18773), .A3(n18772), .B1(n18771), .B2(
        n18770), .B3(n18769), .ZN(P3_U3031) );
  NAND2_X1 U21844 ( .A1(n18830), .A2(n18774), .ZN(n18827) );
  CLKBUF_X1 U21845 ( .A(n18827), .Z(n18836) );
  OAI222_X1 U21846 ( .A1(n18776), .A2(n18833), .B1(n18775), .B2(n18830), .C1(
        n18777), .C2(n18836), .ZN(P3_U3032) );
  OAI222_X1 U21847 ( .A1(n18836), .A2(n18779), .B1(n18778), .B2(n18830), .C1(
        n18777), .C2(n18833), .ZN(P3_U3033) );
  OAI222_X1 U21848 ( .A1(n18827), .A2(n18781), .B1(n18780), .B2(n18830), .C1(
        n18779), .C2(n18833), .ZN(P3_U3034) );
  OAI222_X1 U21849 ( .A1(n18827), .A2(n18783), .B1(n18782), .B2(n18830), .C1(
        n18781), .C2(n18833), .ZN(P3_U3035) );
  OAI222_X1 U21850 ( .A1(n18827), .A2(n18785), .B1(n18784), .B2(n18830), .C1(
        n18783), .C2(n18833), .ZN(P3_U3036) );
  OAI222_X1 U21851 ( .A1(n18827), .A2(n18787), .B1(n18786), .B2(n18830), .C1(
        n18785), .C2(n18833), .ZN(P3_U3037) );
  INV_X1 U21852 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18790) );
  OAI222_X1 U21853 ( .A1(n18827), .A2(n18790), .B1(n18788), .B2(n18830), .C1(
        n18787), .C2(n18833), .ZN(P3_U3038) );
  INV_X1 U21854 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18791) );
  OAI222_X1 U21855 ( .A1(n18790), .A2(n18833), .B1(n18789), .B2(n18830), .C1(
        n18791), .C2(n18836), .ZN(P3_U3039) );
  OAI222_X1 U21856 ( .A1(n18836), .A2(n18793), .B1(n18792), .B2(n18830), .C1(
        n18791), .C2(n18833), .ZN(P3_U3040) );
  OAI222_X1 U21857 ( .A1(n18836), .A2(n18795), .B1(n18794), .B2(n18830), .C1(
        n18793), .C2(n18833), .ZN(P3_U3041) );
  OAI222_X1 U21858 ( .A1(n18836), .A2(n18797), .B1(n18796), .B2(n18830), .C1(
        n18795), .C2(n18833), .ZN(P3_U3042) );
  OAI222_X1 U21859 ( .A1(n18836), .A2(n18799), .B1(n18798), .B2(n18830), .C1(
        n18797), .C2(n18833), .ZN(P3_U3043) );
  OAI222_X1 U21860 ( .A1(n18836), .A2(n18802), .B1(n18800), .B2(n18830), .C1(
        n18799), .C2(n18833), .ZN(P3_U3044) );
  OAI222_X1 U21861 ( .A1(n18802), .A2(n18833), .B1(n18801), .B2(n18830), .C1(
        n18803), .C2(n18836), .ZN(P3_U3045) );
  OAI222_X1 U21862 ( .A1(n18836), .A2(n18805), .B1(n18804), .B2(n18830), .C1(
        n18803), .C2(n18840), .ZN(P3_U3046) );
  OAI222_X1 U21863 ( .A1(n18827), .A2(n18807), .B1(n18806), .B2(n18830), .C1(
        n18805), .C2(n18840), .ZN(P3_U3047) );
  OAI222_X1 U21864 ( .A1(n18827), .A2(n18809), .B1(n18808), .B2(n18830), .C1(
        n18807), .C2(n18840), .ZN(P3_U3048) );
  OAI222_X1 U21865 ( .A1(n18827), .A2(n18811), .B1(n18810), .B2(n18830), .C1(
        n18809), .C2(n18840), .ZN(P3_U3049) );
  OAI222_X1 U21866 ( .A1(n18827), .A2(n18814), .B1(n18812), .B2(n18830), .C1(
        n18811), .C2(n18840), .ZN(P3_U3050) );
  OAI222_X1 U21867 ( .A1(n18814), .A2(n18833), .B1(n18813), .B2(n18830), .C1(
        n18815), .C2(n18836), .ZN(P3_U3051) );
  OAI222_X1 U21868 ( .A1(n18827), .A2(n18817), .B1(n18816), .B2(n18830), .C1(
        n18815), .C2(n18840), .ZN(P3_U3052) );
  OAI222_X1 U21869 ( .A1(n18836), .A2(n18820), .B1(n18818), .B2(n18830), .C1(
        n18817), .C2(n18840), .ZN(P3_U3053) );
  OAI222_X1 U21870 ( .A1(n18820), .A2(n18833), .B1(n18819), .B2(n18830), .C1(
        n18821), .C2(n18836), .ZN(P3_U3054) );
  OAI222_X1 U21871 ( .A1(n18827), .A2(n18823), .B1(n18822), .B2(n18830), .C1(
        n18821), .C2(n18840), .ZN(P3_U3055) );
  OAI222_X1 U21872 ( .A1(n18836), .A2(n18825), .B1(n18824), .B2(n18830), .C1(
        n18823), .C2(n18833), .ZN(P3_U3056) );
  OAI222_X1 U21873 ( .A1(n18827), .A2(n18828), .B1(n18826), .B2(n18830), .C1(
        n18825), .C2(n18833), .ZN(P3_U3057) );
  INV_X1 U21874 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18832) );
  OAI222_X1 U21875 ( .A1(n18836), .A2(n18832), .B1(n18829), .B2(n18830), .C1(
        n18828), .C2(n18833), .ZN(P3_U3058) );
  INV_X1 U21876 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18834) );
  OAI222_X1 U21877 ( .A1(n18832), .A2(n18833), .B1(n18831), .B2(n18830), .C1(
        n18834), .C2(n18836), .ZN(P3_U3059) );
  OAI222_X1 U21878 ( .A1(n18836), .A2(n18839), .B1(n18835), .B2(n18830), .C1(
        n18834), .C2(n18833), .ZN(P3_U3060) );
  INV_X1 U21879 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18838) );
  OAI222_X1 U21880 ( .A1(n18840), .A2(n18839), .B1(n18838), .B2(n18830), .C1(
        n18837), .C2(n18836), .ZN(P3_U3061) );
  INV_X1 U21881 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18841) );
  AOI22_X1 U21882 ( .A1(n18830), .A2(n18842), .B1(n18841), .B2(n18896), .ZN(
        P3_U3274) );
  INV_X1 U21883 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18890) );
  INV_X1 U21884 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18843) );
  AOI22_X1 U21885 ( .A1(n18830), .A2(n18890), .B1(n18843), .B2(n18896), .ZN(
        P3_U3275) );
  INV_X1 U21886 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18844) );
  AOI22_X1 U21887 ( .A1(n18830), .A2(n18845), .B1(n18844), .B2(n18896), .ZN(
        P3_U3276) );
  INV_X1 U21888 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18893) );
  INV_X1 U21889 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18846) );
  AOI22_X1 U21890 ( .A1(n18830), .A2(n18893), .B1(n18846), .B2(n18896), .ZN(
        P3_U3277) );
  INV_X1 U21891 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18848) );
  AOI21_X1 U21892 ( .B1(n9632), .B2(n18848), .A(n18847), .ZN(P3_U3280) );
  OAI21_X1 U21893 ( .B1(n18851), .B2(n18850), .A(n18849), .ZN(P3_U3281) );
  OAI221_X1 U21894 ( .B1(n18854), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18854), 
        .C2(n18853), .A(n18852), .ZN(P3_U3282) );
  NOR3_X1 U21895 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18855), .A3(
        n18868), .ZN(n18856) );
  AOI21_X1 U21896 ( .B1(n18857), .B2(n18881), .A(n18856), .ZN(n18862) );
  INV_X1 U21897 ( .A(n18858), .ZN(n18859) );
  AOI21_X1 U21898 ( .B1(n18883), .B2(n18859), .A(n18888), .ZN(n18861) );
  OAI22_X1 U21899 ( .A1(n18888), .A2(n18862), .B1(n18861), .B2(n18860), .ZN(
        P3_U3285) );
  AOI22_X1 U21900 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n18864), .B2(n18863), .ZN(
        n18874) );
  NOR2_X1 U21901 ( .A1(n18865), .A2(n18884), .ZN(n18875) );
  OAI22_X1 U21902 ( .A1(n18869), .A2(n18868), .B1(n18867), .B2(n18866), .ZN(
        n18870) );
  AOI21_X1 U21903 ( .B1(n18874), .B2(n18875), .A(n18870), .ZN(n18871) );
  AOI22_X1 U21904 ( .A1(n18888), .A2(n18872), .B1(n18871), .B2(n18885), .ZN(
        P3_U3288) );
  INV_X1 U21905 ( .A(n18873), .ZN(n18877) );
  INV_X1 U21906 ( .A(n18874), .ZN(n18876) );
  AOI222_X1 U21907 ( .A1(n18878), .A2(n18883), .B1(n18881), .B2(n18877), .C1(
        n18876), .C2(n18875), .ZN(n18879) );
  AOI22_X1 U21908 ( .A1(n18888), .A2(n18880), .B1(n18879), .B2(n18885), .ZN(
        P3_U3289) );
  AOI222_X1 U21909 ( .A1(n18884), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18883), 
        .B2(n18882), .C1(n18887), .C2(n18881), .ZN(n18886) );
  AOI22_X1 U21910 ( .A1(n18888), .A2(n18887), .B1(n18886), .B2(n18885), .ZN(
        P3_U3290) );
  AOI211_X1 U21911 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_REIP_REG_1__SCAN_IN), .B(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18889) );
  AOI21_X1 U21912 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18889), .ZN(n18891) );
  AOI22_X1 U21913 ( .A1(n18895), .A2(n18891), .B1(n18890), .B2(n18892), .ZN(
        P3_U3292) );
  NOR2_X1 U21914 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n18894) );
  AOI22_X1 U21915 ( .A1(n18895), .A2(n18894), .B1(n18893), .B2(n18892), .ZN(
        P3_U3293) );
  INV_X1 U21916 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18897) );
  AOI22_X1 U21917 ( .A1(n18830), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18897), 
        .B2(n18896), .ZN(P3_U3294) );
  MUX2_X1 U21918 ( .A(P3_MORE_REG_SCAN_IN), .B(n18899), .S(n18898), .Z(
        P3_U3295) );
  OAI21_X1 U21919 ( .B1(n18901), .B2(n18900), .A(n18916), .ZN(n18902) );
  AOI21_X1 U21920 ( .B1(n18903), .B2(n18907), .A(n18902), .ZN(n18913) );
  AOI21_X1 U21921 ( .B1(n18906), .B2(n18905), .A(n18904), .ZN(n18908) );
  OAI211_X1 U21922 ( .C1(n18908), .C2(n18914), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18907), .ZN(n18910) );
  AOI21_X1 U21923 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18910), .A(n18909), 
        .ZN(n18912) );
  NAND2_X1 U21924 ( .A1(n18913), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18911) );
  OAI21_X1 U21925 ( .B1(n18913), .B2(n18912), .A(n18911), .ZN(P3_U3296) );
  MUX2_X1 U21926 ( .A(P3_M_IO_N_REG_SCAN_IN), .B(P3_MEMORYFETCH_REG_SCAN_IN), 
        .S(n18830), .Z(P3_U3297) );
  INV_X1 U21927 ( .A(n18914), .ZN(n18917) );
  OAI21_X1 U21928 ( .B1(P3_READREQUEST_REG_SCAN_IN), .B2(n18918), .A(n18916), 
        .ZN(n18915) );
  OAI21_X1 U21929 ( .B1(n18917), .B2(n18916), .A(n18915), .ZN(P3_U3298) );
  NOR2_X1 U21930 ( .A1(n18918), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18920)
         );
  OAI21_X1 U21931 ( .B1(n18921), .B2(n18920), .A(n18919), .ZN(P3_U3299) );
  INV_X1 U21932 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18922) );
  INV_X1 U21933 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19839) );
  NAND2_X1 U21934 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19839), .ZN(n19832) );
  OR2_X1 U21935 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n19828) );
  OAI21_X1 U21936 ( .B1(n19827), .B2(n19832), .A(n19828), .ZN(n19897) );
  OAI21_X1 U21937 ( .B1(n19827), .B2(n18922), .A(n9634), .ZN(P2_U2815) );
  INV_X1 U21938 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18924) );
  OAI22_X1 U21939 ( .A1(n19965), .A2(n18924), .B1(n9877), .B2(n18923), .ZN(
        P2_U2816) );
  NAND2_X1 U21940 ( .A1(n19971), .A2(n19833), .ZN(n19826) );
  AOI21_X1 U21941 ( .B1(n19827), .B2(n19826), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18925) );
  AOI21_X1 U21942 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n19974), .A(n18925), 
        .ZN(P2_U2817) );
  AOI21_X1 U21943 ( .B1(n19833), .B2(n21030), .A(n9634), .ZN(n19893) );
  INV_X1 U21944 ( .A(n19893), .ZN(n19895) );
  OAI21_X1 U21945 ( .B1(n19897), .B2(n19553), .A(n19895), .ZN(P2_U2818) );
  NOR4_X1 U21946 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18929) );
  NOR4_X1 U21947 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18928) );
  NOR4_X1 U21948 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18927) );
  NOR4_X1 U21949 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18926) );
  NAND4_X1 U21950 ( .A1(n18929), .A2(n18928), .A3(n18927), .A4(n18926), .ZN(
        n18935) );
  NOR4_X1 U21951 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n18933) );
  AOI211_X1 U21952 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n18932) );
  NOR4_X1 U21953 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n18931) );
  NOR4_X1 U21954 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n18930) );
  NAND4_X1 U21955 ( .A1(n18933), .A2(n18932), .A3(n18931), .A4(n18930), .ZN(
        n18934) );
  NOR2_X1 U21956 ( .A1(n18935), .A2(n18934), .ZN(n18943) );
  INV_X1 U21957 ( .A(n18943), .ZN(n18942) );
  NOR2_X1 U21958 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18942), .ZN(n18936) );
  INV_X1 U21959 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18937) );
  INV_X1 U21960 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19892) );
  AOI22_X1 U21961 ( .A1(n18936), .A2(n18937), .B1(n18942), .B2(n19892), .ZN(
        P2_U2820) );
  INV_X1 U21962 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19896) );
  INV_X1 U21963 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19894) );
  NAND3_X1 U21964 ( .A1(n18937), .A2(n19896), .A3(n19894), .ZN(n18941) );
  INV_X1 U21965 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19890) );
  AOI22_X1 U21966 ( .A1(n18936), .A2(n18941), .B1(n18942), .B2(n19890), .ZN(
        P2_U2821) );
  NAND2_X1 U21967 ( .A1(n18936), .A2(n19896), .ZN(n18940) );
  OAI21_X1 U21968 ( .B1(n10595), .B2(n18937), .A(n18943), .ZN(n18938) );
  OAI21_X1 U21969 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18943), .A(n18938), 
        .ZN(n18939) );
  OAI221_X1 U21970 ( .B1(n18940), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18940), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18939), .ZN(P2_U2822) );
  INV_X1 U21971 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19888) );
  OAI221_X1 U21972 ( .B1(n18943), .B2(n19888), .C1(n18942), .C2(n18941), .A(
        n18940), .ZN(P2_U2823) );
  NAND2_X1 U21973 ( .A1(n19049), .A2(n14079), .ZN(n19071) );
  AOI211_X1 U21974 ( .C1(n18951), .C2(n18945), .A(n18944), .B(n19071), .ZN(
        n18949) );
  AOI22_X1 U21975 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n18996), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n19054), .ZN(n18946) );
  OAI211_X1 U21976 ( .C1(n18947), .C2(n9646), .A(n18946), .B(n19033), .ZN(
        n18948) );
  AOI211_X1 U21977 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n19055), .A(n18949), .B(
        n18948), .ZN(n18953) );
  NOR2_X1 U21978 ( .A1(n19822), .A2(n14079), .ZN(n19067) );
  AOI22_X1 U21979 ( .A1(n18951), .A2(n19067), .B1(n19062), .B2(n18950), .ZN(
        n18952) );
  OAI211_X1 U21980 ( .C1(n18954), .C2(n19053), .A(n18953), .B(n18952), .ZN(
        P2_U2838) );
  NAND2_X1 U21981 ( .A1(n18963), .A2(n18955), .ZN(n18967) );
  INV_X1 U21982 ( .A(n18956), .ZN(n18965) );
  INV_X1 U21983 ( .A(n18957), .ZN(n18959) );
  AOI21_X1 U21984 ( .B1(n19055), .B2(P2_EBX_REG_15__SCAN_IN), .A(n19192), .ZN(
        n18958) );
  OAI21_X1 U21985 ( .B1(n18959), .B2(n19036), .A(n18958), .ZN(n18962) );
  OAI22_X1 U21986 ( .A1(n18960), .A2(n19006), .B1(n12839), .B2(n19035), .ZN(
        n18961) );
  AOI211_X1 U21987 ( .C1(n19067), .C2(n18963), .A(n18962), .B(n18961), .ZN(
        n18964) );
  OAI21_X1 U21988 ( .B1(n18965), .B2(n9646), .A(n18964), .ZN(n18966) );
  AOI21_X1 U21989 ( .B1(n18968), .B2(n18967), .A(n18966), .ZN(n18969) );
  OAI21_X1 U21990 ( .B1(n19087), .B2(n19053), .A(n18969), .ZN(P2_U2840) );
  NOR2_X1 U21991 ( .A1(n18993), .A2(n18970), .ZN(n18973) );
  XOR2_X1 U21992 ( .A(n18973), .B(n18972), .Z(n18980) );
  AOI22_X1 U21993 ( .A1(n18974), .A2(n19031), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n19055), .ZN(n18975) );
  OAI211_X1 U21994 ( .C1(n12810), .C2(n19035), .A(n18975), .B(n19033), .ZN(
        n18976) );
  AOI21_X1 U21995 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19068), .A(
        n18976), .ZN(n18979) );
  AOI22_X1 U21996 ( .A1(n18977), .A2(n19062), .B1(n19056), .B2(n19088), .ZN(
        n18978) );
  OAI211_X1 U21997 ( .C1(n19822), .C2(n18980), .A(n18979), .B(n18978), .ZN(
        P2_U2841) );
  OAI21_X1 U21998 ( .B1(n12807), .B2(n19035), .A(n19033), .ZN(n18984) );
  INV_X1 U21999 ( .A(n18981), .ZN(n18982) );
  OAI22_X1 U22000 ( .A1(n18982), .A2(n9646), .B1(n19017), .B2(n10474), .ZN(
        n18983) );
  AOI211_X1 U22001 ( .C1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n18996), .A(
        n18984), .B(n18983), .ZN(n18991) );
  NAND2_X1 U22002 ( .A1(n14079), .A2(n18985), .ZN(n18986) );
  XNOR2_X1 U22003 ( .A(n18987), .B(n18986), .ZN(n18989) );
  AOI22_X1 U22004 ( .A1(n18989), .A2(n19049), .B1(n19062), .B2(n18988), .ZN(
        n18990) );
  OAI211_X1 U22005 ( .C1(n19093), .C2(n19053), .A(n18991), .B(n18990), .ZN(
        P2_U2842) );
  NOR2_X1 U22006 ( .A1(n18993), .A2(n18992), .ZN(n18995) );
  XOR2_X1 U22007 ( .A(n18995), .B(n18994), .Z(n19003) );
  AOI22_X1 U22008 ( .A1(n19055), .A2(P2_EBX_REG_12__SCAN_IN), .B1(n18996), 
        .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18997) );
  OAI21_X1 U22009 ( .B1(n18998), .B2(n9646), .A(n18997), .ZN(n18999) );
  AOI211_X1 U22010 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19054), .A(n19192), 
        .B(n18999), .ZN(n19002) );
  AOI22_X1 U22011 ( .A1(n19094), .A2(n19056), .B1(n19062), .B2(n19000), .ZN(
        n19001) );
  OAI211_X1 U22012 ( .C1(n19822), .C2(n19003), .A(n19002), .B(n19001), .ZN(
        P2_U2843) );
  OAI222_X1 U22013 ( .A1(n19006), .A2(n16171), .B1(n19005), .B2(n19017), .C1(
        n19004), .C2(n9646), .ZN(n19007) );
  AOI211_X1 U22014 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n19054), .A(n19192), 
        .B(n19007), .ZN(n19014) );
  NAND2_X1 U22015 ( .A1(n14079), .A2(n19008), .ZN(n19009) );
  XNOR2_X1 U22016 ( .A(n19010), .B(n19009), .ZN(n19012) );
  AOI22_X1 U22017 ( .A1(n19012), .A2(n19049), .B1(n19062), .B2(n19011), .ZN(
        n19013) );
  OAI211_X1 U22018 ( .C1(n19099), .C2(n19053), .A(n19014), .B(n19013), .ZN(
        P2_U2844) );
  OAI21_X1 U22019 ( .B1(n12744), .B2(n19035), .A(n19033), .ZN(n19020) );
  INV_X1 U22020 ( .A(n19015), .ZN(n19018) );
  OAI22_X1 U22021 ( .A1(n19018), .A2(n9646), .B1(n19017), .B2(n19016), .ZN(
        n19019) );
  AOI211_X1 U22022 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n19068), .A(
        n19020), .B(n19019), .ZN(n19027) );
  NAND2_X1 U22023 ( .A1(n14079), .A2(n19021), .ZN(n19022) );
  XNOR2_X1 U22024 ( .A(n19023), .B(n19022), .ZN(n19025) );
  AOI22_X1 U22025 ( .A1(n19025), .A2(n19049), .B1(n19062), .B2(n19024), .ZN(
        n19026) );
  OAI211_X1 U22026 ( .C1(n19053), .C2(n19105), .A(n19027), .B(n19026), .ZN(
        P2_U2846) );
  NAND2_X1 U22027 ( .A1(n14079), .A2(n19028), .ZN(n19030) );
  XOR2_X1 U22028 ( .A(n19030), .B(n19029), .Z(n19041) );
  AOI22_X1 U22029 ( .A1(n19032), .A2(n19031), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19055), .ZN(n19034) );
  OAI211_X1 U22030 ( .C1(n19848), .C2(n19035), .A(n19034), .B(n19033), .ZN(
        n19039) );
  OAI22_X1 U22031 ( .A1(n19037), .A2(n19036), .B1(n19111), .B2(n19053), .ZN(
        n19038) );
  AOI211_X1 U22032 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19068), .A(
        n19039), .B(n19038), .ZN(n19040) );
  OAI21_X1 U22033 ( .B1(n19041), .B2(n19822), .A(n19040), .ZN(P2_U2848) );
  AOI22_X1 U22034 ( .A1(n19055), .A2(P2_EBX_REG_5__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n19068), .ZN(n19042) );
  OAI21_X1 U22035 ( .B1(n19043), .B2(n9646), .A(n19042), .ZN(n19044) );
  AOI211_X1 U22036 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19054), .A(n19192), .B(
        n19044), .ZN(n19052) );
  NAND2_X1 U22037 ( .A1(n14079), .A2(n19045), .ZN(n19046) );
  XNOR2_X1 U22038 ( .A(n19047), .B(n19046), .ZN(n19050) );
  AOI22_X1 U22039 ( .A1(n19050), .A2(n19049), .B1(n19062), .B2(n19048), .ZN(
        n19051) );
  OAI211_X1 U22040 ( .C1(n19053), .C2(n19118), .A(n19052), .B(n19051), .ZN(
        P2_U2850) );
  AOI22_X1 U22041 ( .A1(n19055), .A2(P2_EBX_REG_0__SCAN_IN), .B1(n19054), .B2(
        P2_REIP_REG_0__SCAN_IN), .ZN(n19059) );
  NAND2_X1 U22042 ( .A1(n19057), .A2(n19056), .ZN(n19058) );
  OAI211_X1 U22043 ( .C1(n19060), .C2(n9646), .A(n19059), .B(n19058), .ZN(
        n19061) );
  AOI21_X1 U22044 ( .B1(n19063), .B2(n19062), .A(n19061), .ZN(n19064) );
  OAI21_X1 U22045 ( .B1(n19933), .B2(n19065), .A(n19064), .ZN(n19066) );
  INV_X1 U22046 ( .A(n19066), .ZN(n19070) );
  OAI21_X1 U22047 ( .B1(n19068), .B2(n19067), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19069) );
  OAI211_X1 U22048 ( .C1(n19072), .C2(n19071), .A(n19070), .B(n19069), .ZN(
        P2_U2855) );
  AOI22_X1 U22049 ( .A1(n19073), .A2(n19131), .B1(n19078), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19075) );
  AOI22_X1 U22050 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19130), .B1(n19079), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19074) );
  NAND2_X1 U22051 ( .A1(n19075), .A2(n19074), .ZN(P2_U2888) );
  AOI22_X1 U22052 ( .A1(n19077), .A2(n19076), .B1(n19130), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19084) );
  AOI22_X1 U22053 ( .A1(n19079), .A2(BUF1_REG_16__SCAN_IN), .B1(n19078), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n19083) );
  AOI22_X1 U22054 ( .A1(n19081), .A2(n19085), .B1(n19131), .B2(n19080), .ZN(
        n19082) );
  NAND3_X1 U22055 ( .A1(n19084), .A2(n19083), .A3(n19082), .ZN(P2_U2903) );
  OAI222_X1 U22056 ( .A1(n19087), .A2(n19119), .B1(n13373), .B2(n19121), .C1(
        n19086), .C2(n19139), .ZN(P2_U2904) );
  INV_X1 U22057 ( .A(n19088), .ZN(n19091) );
  AOI22_X1 U22058 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19130), .B1(n19089), 
        .B2(n19107), .ZN(n19090) );
  OAI21_X1 U22059 ( .B1(n19119), .B2(n19091), .A(n19090), .ZN(P2_U2905) );
  INV_X1 U22060 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19145) );
  OAI222_X1 U22061 ( .A1(n19093), .A2(n19119), .B1(n19145), .B2(n19121), .C1(
        n19139), .C2(n19092), .ZN(P2_U2906) );
  INV_X1 U22062 ( .A(n19094), .ZN(n19097) );
  AOI22_X1 U22063 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19130), .B1(n19095), 
        .B2(n19107), .ZN(n19096) );
  OAI21_X1 U22064 ( .B1(n19119), .B2(n19097), .A(n19096), .ZN(P2_U2907) );
  INV_X1 U22065 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19149) );
  OAI222_X1 U22066 ( .A1(n19099), .A2(n19119), .B1(n19149), .B2(n19121), .C1(
        n19139), .C2(n19098), .ZN(P2_U2908) );
  INV_X1 U22067 ( .A(n19100), .ZN(n19103) );
  AOI22_X1 U22068 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19130), .B1(n19101), 
        .B2(n19107), .ZN(n19102) );
  OAI21_X1 U22069 ( .B1(n19119), .B2(n19103), .A(n19102), .ZN(P2_U2909) );
  INV_X1 U22070 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19153) );
  OAI222_X1 U22071 ( .A1(n19105), .A2(n19119), .B1(n19153), .B2(n19121), .C1(
        n19139), .C2(n19104), .ZN(P2_U2910) );
  INV_X1 U22072 ( .A(n19106), .ZN(n19110) );
  AOI22_X1 U22073 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19130), .B1(n19108), .B2(
        n19107), .ZN(n19109) );
  OAI21_X1 U22074 ( .B1(n19119), .B2(n19110), .A(n19109), .ZN(P2_U2911) );
  OAI222_X1 U22075 ( .A1(n19111), .A2(n19119), .B1(n19158), .B2(n19121), .C1(
        n19139), .C2(n19264), .ZN(P2_U2912) );
  INV_X1 U22076 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19160) );
  OAI222_X1 U22077 ( .A1(n19112), .A2(n19119), .B1(n19160), .B2(n19121), .C1(
        n19139), .C2(n19255), .ZN(P2_U2913) );
  INV_X1 U22078 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19162) );
  OAI22_X1 U22079 ( .A1(n19162), .A2(n19121), .B1(n19252), .B2(n19139), .ZN(
        n19113) );
  INV_X1 U22080 ( .A(n19113), .ZN(n19117) );
  OR3_X1 U22081 ( .A1(n19115), .A2(n19114), .A3(n19135), .ZN(n19116) );
  OAI211_X1 U22082 ( .C1(n19119), .C2(n19118), .A(n19117), .B(n19116), .ZN(
        P2_U2914) );
  INV_X1 U22083 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19120) );
  OAI22_X1 U22084 ( .A1(n19898), .A2(n19122), .B1(n19121), .B2(n19120), .ZN(
        n19123) );
  INV_X1 U22085 ( .A(n19123), .ZN(n19129) );
  AOI21_X1 U22086 ( .B1(n19126), .B2(n19125), .A(n19124), .ZN(n19127) );
  OR2_X1 U22087 ( .A1(n19127), .A2(n19135), .ZN(n19128) );
  OAI211_X1 U22088 ( .C1(n19243), .C2(n19139), .A(n19129), .B(n19128), .ZN(
        P2_U2916) );
  AOI22_X1 U22089 ( .A1(n19131), .A2(n19927), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19130), .ZN(n19138) );
  AOI21_X1 U22090 ( .B1(n19134), .B2(n19133), .A(n19132), .ZN(n19136) );
  OR2_X1 U22091 ( .A1(n19136), .A2(n19135), .ZN(n19137) );
  OAI211_X1 U22092 ( .C1(n19233), .C2(n19139), .A(n19138), .B(n19137), .ZN(
        P2_U2918) );
  AND2_X1 U22093 ( .A1(n19154), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U22094 ( .A1(n19968), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19170), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19141) );
  OAI21_X1 U22095 ( .B1(n13373), .B2(n19172), .A(n19141), .ZN(P2_U2936) );
  AOI22_X1 U22096 ( .A1(n19968), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19170), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19142) );
  OAI21_X1 U22097 ( .B1(n19143), .B2(n19172), .A(n19142), .ZN(P2_U2937) );
  AOI22_X1 U22098 ( .A1(n19968), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19170), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19144) );
  OAI21_X1 U22099 ( .B1(n19145), .B2(n19172), .A(n19144), .ZN(P2_U2938) );
  AOI22_X1 U22100 ( .A1(n19968), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19170), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19146) );
  OAI21_X1 U22101 ( .B1(n19147), .B2(n19172), .A(n19146), .ZN(P2_U2939) );
  AOI22_X1 U22102 ( .A1(n19968), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19154), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19148) );
  OAI21_X1 U22103 ( .B1(n19149), .B2(n19172), .A(n19148), .ZN(P2_U2940) );
  AOI22_X1 U22104 ( .A1(n19968), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19154), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19150) );
  OAI21_X1 U22105 ( .B1(n19151), .B2(n19172), .A(n19150), .ZN(P2_U2941) );
  AOI22_X1 U22106 ( .A1(n19968), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19154), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19152) );
  OAI21_X1 U22107 ( .B1(n19153), .B2(n19172), .A(n19152), .ZN(P2_U2942) );
  AOI22_X1 U22108 ( .A1(n19968), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19154), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19155) );
  OAI21_X1 U22109 ( .B1(n19156), .B2(n19172), .A(n19155), .ZN(P2_U2943) );
  AOI22_X1 U22110 ( .A1(n19968), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19170), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19157) );
  OAI21_X1 U22111 ( .B1(n19158), .B2(n19172), .A(n19157), .ZN(P2_U2944) );
  AOI22_X1 U22112 ( .A1(n19968), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19170), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19159) );
  OAI21_X1 U22113 ( .B1(n19160), .B2(n19172), .A(n19159), .ZN(P2_U2945) );
  AOI22_X1 U22114 ( .A1(n19968), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19170), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19161) );
  OAI21_X1 U22115 ( .B1(n19162), .B2(n19172), .A(n19161), .ZN(P2_U2946) );
  INV_X1 U22116 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19164) );
  AOI22_X1 U22117 ( .A1(n19968), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19170), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19163) );
  OAI21_X1 U22118 ( .B1(n19164), .B2(n19172), .A(n19163), .ZN(P2_U2947) );
  AOI22_X1 U22119 ( .A1(n19968), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19170), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19165) );
  OAI21_X1 U22120 ( .B1(n19120), .B2(n19172), .A(n19165), .ZN(P2_U2948) );
  AOI22_X1 U22121 ( .A1(n19968), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19170), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19166) );
  OAI21_X1 U22122 ( .B1(n19167), .B2(n19172), .A(n19166), .ZN(P2_U2949) );
  INV_X1 U22123 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19169) );
  AOI22_X1 U22124 ( .A1(n19968), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19170), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19168) );
  OAI21_X1 U22125 ( .B1(n19169), .B2(n19172), .A(n19168), .ZN(P2_U2950) );
  AOI22_X1 U22126 ( .A1(n19968), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19170), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19171) );
  OAI21_X1 U22127 ( .B1(n19173), .B2(n19172), .A(n19171), .ZN(P2_U2951) );
  AOI22_X1 U22128 ( .A1(n19187), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19174), .ZN(n19180) );
  INV_X1 U22129 ( .A(n19175), .ZN(n19177) );
  AOI222_X1 U22130 ( .A1(n19178), .A2(n11014), .B1(n19194), .B2(n19177), .C1(
        n19188), .C2(n19176), .ZN(n19179) );
  OAI211_X1 U22131 ( .C1(n19182), .C2(n19181), .A(n19180), .B(n19179), .ZN(
        P2_U3010) );
  AOI21_X1 U22132 ( .B1(n19185), .B2(n19184), .A(n19183), .ZN(n19186) );
  XNOR2_X1 U22133 ( .A(n19186), .B(n19191), .ZN(n19205) );
  AOI22_X1 U22134 ( .A1(n19205), .A2(n19188), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19187), .ZN(n19200) );
  AOI21_X1 U22135 ( .B1(n19191), .B2(n19190), .A(n19189), .ZN(n19203) );
  AND2_X1 U22136 ( .A1(n19192), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n19211) );
  AOI21_X1 U22137 ( .B1(n11014), .B2(n19203), .A(n19211), .ZN(n19198) );
  NAND2_X1 U22138 ( .A1(n19194), .A2(n19193), .ZN(n19197) );
  NAND2_X1 U22139 ( .A1(n19195), .A2(n14073), .ZN(n19196) );
  AND3_X1 U22140 ( .A1(n19198), .A2(n19197), .A3(n19196), .ZN(n19199) );
  NAND2_X1 U22141 ( .A1(n19200), .A2(n19199), .ZN(P2_U3013) );
  OAI21_X1 U22142 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n19201), .ZN(n19215) );
  AOI22_X1 U22143 ( .A1(n19204), .A2(n19203), .B1(n19202), .B2(n19927), .ZN(
        n19214) );
  INV_X1 U22144 ( .A(n19205), .ZN(n19208) );
  OAI22_X1 U22145 ( .A1(n19209), .A2(n19208), .B1(n19207), .B2(n19206), .ZN(
        n19210) );
  AOI211_X1 U22146 ( .C1(n19212), .C2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n19211), .B(n19210), .ZN(n19213) );
  OAI211_X1 U22147 ( .C1(n19216), .C2(n19215), .A(n19214), .B(n19213), .ZN(
        P2_U3045) );
  AOI22_X1 U22148 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19259), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19258), .ZN(n19726) );
  AOI22_X1 U22149 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19259), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19258), .ZN(n19766) );
  INV_X1 U22150 ( .A(n19250), .ZN(n19261) );
  AND2_X1 U22151 ( .A1(n19220), .A2(n19261), .ZN(n19755) );
  NOR2_X1 U22152 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19328) );
  NAND2_X1 U22153 ( .A1(n19328), .A2(n19929), .ZN(n19272) );
  NOR2_X1 U22154 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19272), .ZN(
        n19263) );
  AOI22_X1 U22155 ( .A1(n19798), .A2(n19714), .B1(n19755), .B2(n19263), .ZN(
        n19232) );
  OAI21_X1 U22156 ( .B1(n19798), .B2(n19294), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19221) );
  NAND2_X1 U22157 ( .A1(n19221), .A2(n19902), .ZN(n19230) );
  NOR2_X1 U22158 ( .A1(n19804), .A2(n19263), .ZN(n19229) );
  INV_X1 U22159 ( .A(n19229), .ZN(n19224) );
  INV_X1 U22160 ( .A(n19263), .ZN(n19222) );
  OAI211_X1 U22161 ( .C1(n10755), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19222), 
        .B(n19906), .ZN(n19223) );
  OAI211_X1 U22162 ( .C1(n19230), .C2(n19224), .A(n19761), .B(n19223), .ZN(
        n19266) );
  OAI21_X1 U22163 ( .B1(n19227), .B2(n19263), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19228) );
  AOI22_X1 U22164 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19266), .B1(
        n19226), .B2(n19265), .ZN(n19231) );
  OAI211_X1 U22165 ( .C1(n19726), .C2(n19291), .A(n19232), .B(n19231), .ZN(
        P2_U3048) );
  AOI22_X1 U22166 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19259), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19258), .ZN(n19771) );
  AOI22_X1 U22167 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19259), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19258), .ZN(n19674) );
  NOR2_X2 U22168 ( .A1(n13380), .A2(n19250), .ZN(n19767) );
  AOI22_X1 U22169 ( .A1(n19798), .A2(n19768), .B1(n19767), .B2(n19263), .ZN(
        n19236) );
  AOI22_X1 U22170 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19266), .B1(
        n19234), .B2(n19265), .ZN(n19235) );
  OAI211_X1 U22171 ( .C1(n19771), .C2(n19291), .A(n19236), .B(n19235), .ZN(
        P2_U3049) );
  AOI22_X1 U22172 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19259), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19258), .ZN(n19776) );
  AOI22_X1 U22173 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19258), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19259), .ZN(n19732) );
  INV_X1 U22174 ( .A(n19732), .ZN(n19773) );
  NOR2_X2 U22175 ( .A1(n19237), .A2(n19250), .ZN(n19772) );
  AOI22_X1 U22176 ( .A1(n19798), .A2(n19773), .B1(n19772), .B2(n19263), .ZN(
        n19241) );
  AOI22_X1 U22177 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19266), .B1(
        n19239), .B2(n19265), .ZN(n19240) );
  OAI211_X1 U22178 ( .C1(n19776), .C2(n19291), .A(n19241), .B(n19240), .ZN(
        P2_U3050) );
  AOI22_X1 U22179 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19259), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19258), .ZN(n19736) );
  AOI22_X1 U22180 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19259), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19258), .ZN(n19782) );
  AOI22_X1 U22181 ( .A1(n19798), .A2(n19733), .B1(n19777), .B2(n19263), .ZN(
        n19245) );
  NOR2_X2 U22182 ( .A1(n19243), .A2(n19618), .ZN(n19778) );
  AOI22_X1 U22183 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19266), .B1(
        n19778), .B2(n19265), .ZN(n19244) );
  OAI211_X1 U22184 ( .C1(n19736), .C2(n19291), .A(n19245), .B(n19244), .ZN(
        P2_U3051) );
  AOI22_X1 U22185 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19259), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19258), .ZN(n19788) );
  AOI22_X1 U22186 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19259), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19258), .ZN(n19740) );
  NOR2_X2 U22187 ( .A1(n10553), .A2(n19250), .ZN(n19783) );
  AOI22_X1 U22188 ( .A1(n19798), .A2(n19785), .B1(n19783), .B2(n19263), .ZN(
        n19248) );
  NOR2_X2 U22189 ( .A1(n19246), .A2(n19618), .ZN(n19784) );
  AOI22_X1 U22190 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19266), .B1(
        n19784), .B2(n19265), .ZN(n19247) );
  OAI211_X1 U22191 ( .C1(n19788), .C2(n19291), .A(n19248), .B(n19247), .ZN(
        P2_U3052) );
  AOI22_X2 U22192 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19259), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19258), .ZN(n19794) );
  AOI22_X1 U22193 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19259), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19258), .ZN(n19249) );
  NOR2_X2 U22194 ( .A1(n19251), .A2(n19250), .ZN(n19789) );
  AOI22_X1 U22195 ( .A1(n19798), .A2(n19791), .B1(n19789), .B2(n19263), .ZN(
        n19254) );
  NOR2_X2 U22196 ( .A1(n19252), .A2(n19618), .ZN(n19790) );
  AOI22_X1 U22197 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19266), .B1(
        n19790), .B2(n19265), .ZN(n19253) );
  OAI211_X1 U22198 ( .C1(n19794), .C2(n19291), .A(n19254), .B(n19253), .ZN(
        P2_U3053) );
  AOI22_X1 U22199 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19259), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19258), .ZN(n19702) );
  AOI22_X1 U22200 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19259), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19258), .ZN(n19802) );
  AND2_X1 U22201 ( .A1(n12904), .A2(n19261), .ZN(n19795) );
  AOI22_X1 U22202 ( .A1(n19798), .A2(n19699), .B1(n19795), .B2(n19263), .ZN(
        n19257) );
  NOR2_X2 U22203 ( .A1(n19255), .A2(n19618), .ZN(n19796) );
  AOI22_X1 U22204 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19266), .B1(
        n19796), .B2(n19265), .ZN(n19256) );
  OAI211_X1 U22205 ( .C1(n19702), .C2(n19291), .A(n19257), .B(n19256), .ZN(
        P2_U3054) );
  AOI22_X2 U22206 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19259), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19258), .ZN(n19813) );
  AOI22_X1 U22207 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19259), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19258), .ZN(n19260) );
  AND2_X1 U22208 ( .A1(n19262), .A2(n19261), .ZN(n19803) );
  AOI22_X1 U22209 ( .A1(n19798), .A2(n19807), .B1(n19803), .B2(n19263), .ZN(
        n19268) );
  NOR2_X2 U22210 ( .A1(n19264), .A2(n19618), .ZN(n19805) );
  AOI22_X1 U22211 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19266), .B1(
        n19805), .B2(n19265), .ZN(n19267) );
  OAI211_X1 U22212 ( .C1(n19813), .C2(n19291), .A(n19268), .B(n19267), .ZN(
        P2_U3055) );
  INV_X1 U22213 ( .A(n19269), .ZN(n19452) );
  NAND2_X1 U22214 ( .A1(n19929), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19518) );
  INV_X1 U22215 ( .A(n19328), .ZN(n19327) );
  NOR2_X1 U22216 ( .A1(n19518), .A2(n19327), .ZN(n19292) );
  OR2_X1 U22217 ( .A1(n19292), .A2(n19959), .ZN(n19270) );
  OR2_X1 U22218 ( .A1(n10741), .A2(n19270), .ZN(n19274) );
  INV_X1 U22219 ( .A(n19274), .ZN(n19271) );
  AOI211_X2 U22220 ( .C1(n19272), .C2(n19959), .A(n19452), .B(n19271), .ZN(
        n19293) );
  AOI22_X1 U22221 ( .A1(n19293), .A2(n19226), .B1(n19755), .B2(n19292), .ZN(
        n19278) );
  NAND2_X1 U22222 ( .A1(n19904), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19907) );
  OAI21_X1 U22223 ( .B1(n19907), .B2(n19520), .A(n19272), .ZN(n19275) );
  OR2_X1 U22224 ( .A1(n19292), .A2(n19931), .ZN(n19273) );
  NAND4_X1 U22225 ( .A1(n19275), .A2(n19761), .A3(n19274), .A4(n19273), .ZN(
        n19295) );
  NAND2_X1 U22226 ( .A1(n19276), .A2(n19454), .ZN(n19300) );
  INV_X1 U22227 ( .A(n19726), .ZN(n19763) );
  AOI22_X1 U22228 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19295), .B1(
        n19323), .B2(n19763), .ZN(n19277) );
  OAI211_X1 U22229 ( .C1(n19766), .C2(n19291), .A(n19278), .B(n19277), .ZN(
        P2_U3056) );
  AOI22_X1 U22230 ( .A1(n19293), .A2(n19234), .B1(n19767), .B2(n19292), .ZN(
        n19280) );
  INV_X1 U22231 ( .A(n19771), .ZN(n19671) );
  AOI22_X1 U22232 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19295), .B1(
        n19323), .B2(n19671), .ZN(n19279) );
  OAI211_X1 U22233 ( .C1(n19674), .C2(n19291), .A(n19280), .B(n19279), .ZN(
        P2_U3057) );
  AOI22_X1 U22234 ( .A1(n19293), .A2(n19239), .B1(n19772), .B2(n19292), .ZN(
        n19282) );
  INV_X1 U22235 ( .A(n19776), .ZN(n19729) );
  AOI22_X1 U22236 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19295), .B1(
        n19323), .B2(n19729), .ZN(n19281) );
  OAI211_X1 U22237 ( .C1(n19732), .C2(n19291), .A(n19282), .B(n19281), .ZN(
        P2_U3058) );
  AOI22_X1 U22238 ( .A1(n19293), .A2(n19778), .B1(n19777), .B2(n19292), .ZN(
        n19284) );
  INV_X1 U22239 ( .A(n19736), .ZN(n19779) );
  AOI22_X1 U22240 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19295), .B1(
        n19323), .B2(n19779), .ZN(n19283) );
  OAI211_X1 U22241 ( .C1(n19782), .C2(n19291), .A(n19284), .B(n19283), .ZN(
        P2_U3059) );
  AOI22_X1 U22242 ( .A1(n19293), .A2(n19784), .B1(n19783), .B2(n19292), .ZN(
        n19286) );
  INV_X1 U22243 ( .A(n19788), .ZN(n19737) );
  AOI22_X1 U22244 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19295), .B1(
        n19323), .B2(n19737), .ZN(n19285) );
  OAI211_X1 U22245 ( .C1(n19740), .C2(n19291), .A(n19286), .B(n19285), .ZN(
        P2_U3060) );
  AOI22_X1 U22246 ( .A1(n19293), .A2(n19790), .B1(n19789), .B2(n19292), .ZN(
        n19288) );
  AOI22_X1 U22247 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19295), .B1(
        n19294), .B2(n19791), .ZN(n19287) );
  OAI211_X1 U22248 ( .C1(n19794), .C2(n19300), .A(n19288), .B(n19287), .ZN(
        P2_U3061) );
  AOI22_X1 U22249 ( .A1(n19293), .A2(n19796), .B1(n19795), .B2(n19292), .ZN(
        n19290) );
  INV_X1 U22250 ( .A(n19702), .ZN(n19797) );
  AOI22_X1 U22251 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19295), .B1(
        n19323), .B2(n19797), .ZN(n19289) );
  OAI211_X1 U22252 ( .C1(n19802), .C2(n19291), .A(n19290), .B(n19289), .ZN(
        P2_U3062) );
  AOI22_X1 U22253 ( .A1(n19293), .A2(n19805), .B1(n19803), .B2(n19292), .ZN(
        n19297) );
  AOI22_X1 U22254 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19295), .B1(
        n19294), .B2(n19807), .ZN(n19296) );
  OAI211_X1 U22255 ( .C1(n19813), .C2(n19300), .A(n19297), .B(n19296), .ZN(
        P2_U3063) );
  NOR2_X1 U22256 ( .A1(n19929), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19549) );
  AND2_X1 U22257 ( .A1(n19549), .A2(n19328), .ZN(n19321) );
  OAI21_X1 U22258 ( .B1(n19303), .B2(n19321), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19299) );
  NOR2_X1 U22259 ( .A1(n19551), .A2(n19327), .ZN(n19301) );
  INV_X1 U22260 ( .A(n19301), .ZN(n19298) );
  NAND2_X1 U22261 ( .A1(n19299), .A2(n19298), .ZN(n19322) );
  AOI22_X1 U22262 ( .A1(n19322), .A2(n19226), .B1(n19755), .B2(n19321), .ZN(
        n19308) );
  AOI21_X1 U22263 ( .B1(n19346), .B2(n19300), .A(n19553), .ZN(n19302) );
  NOR2_X1 U22264 ( .A1(n19302), .A2(n19301), .ZN(n19305) );
  AOI21_X1 U22265 ( .B1(n19303), .B2(n19931), .A(n19321), .ZN(n19304) );
  MUX2_X1 U22266 ( .A(n19305), .B(n19304), .S(n19906), .Z(n19306) );
  AOI22_X1 U22267 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19714), .ZN(n19307) );
  OAI211_X1 U22268 ( .C1(n19726), .C2(n19346), .A(n19308), .B(n19307), .ZN(
        P2_U3064) );
  AOI22_X1 U22269 ( .A1(n19322), .A2(n19234), .B1(n19767), .B2(n19321), .ZN(
        n19310) );
  AOI22_X1 U22270 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19768), .ZN(n19309) );
  OAI211_X1 U22271 ( .C1(n19771), .C2(n19346), .A(n19310), .B(n19309), .ZN(
        P2_U3065) );
  AOI22_X1 U22272 ( .A1(n19322), .A2(n19239), .B1(n19772), .B2(n19321), .ZN(
        n19312) );
  AOI22_X1 U22273 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19773), .ZN(n19311) );
  OAI211_X1 U22274 ( .C1(n19776), .C2(n19346), .A(n19312), .B(n19311), .ZN(
        P2_U3066) );
  AOI22_X1 U22275 ( .A1(n19322), .A2(n19778), .B1(n19777), .B2(n19321), .ZN(
        n19314) );
  AOI22_X1 U22276 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19733), .ZN(n19313) );
  OAI211_X1 U22277 ( .C1(n19736), .C2(n19346), .A(n19314), .B(n19313), .ZN(
        P2_U3067) );
  AOI22_X1 U22278 ( .A1(n19322), .A2(n19784), .B1(n19783), .B2(n19321), .ZN(
        n19316) );
  AOI22_X1 U22279 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19785), .ZN(n19315) );
  OAI211_X1 U22280 ( .C1(n19788), .C2(n19346), .A(n19316), .B(n19315), .ZN(
        P2_U3068) );
  AOI22_X1 U22281 ( .A1(n19322), .A2(n19790), .B1(n19789), .B2(n19321), .ZN(
        n19318) );
  AOI22_X1 U22282 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19791), .ZN(n19317) );
  OAI211_X1 U22283 ( .C1(n19794), .C2(n19346), .A(n19318), .B(n19317), .ZN(
        P2_U3069) );
  AOI22_X1 U22284 ( .A1(n19322), .A2(n19796), .B1(n19795), .B2(n19321), .ZN(
        n19320) );
  AOI22_X1 U22285 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19699), .ZN(n19319) );
  OAI211_X1 U22286 ( .C1(n19702), .C2(n19346), .A(n19320), .B(n19319), .ZN(
        P2_U3070) );
  AOI22_X1 U22287 ( .A1(n19322), .A2(n19805), .B1(n19803), .B2(n19321), .ZN(
        n19326) );
  AOI22_X1 U22288 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19807), .ZN(n19325) );
  OAI211_X1 U22289 ( .C1(n19813), .C2(n19346), .A(n19326), .B(n19325), .ZN(
        P2_U3071) );
  NOR2_X1 U22290 ( .A1(n19581), .A2(n19327), .ZN(n19351) );
  AOI22_X1 U22291 ( .A1(n19763), .A2(n19384), .B1(n19351), .B2(n19755), .ZN(
        n19337) );
  OAI21_X1 U22292 ( .B1(n19907), .B2(n19589), .A(n19902), .ZN(n19335) );
  NAND2_X1 U22293 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19328), .ZN(
        n19334) );
  INV_X1 U22294 ( .A(n19334), .ZN(n19332) );
  INV_X1 U22295 ( .A(n19351), .ZN(n19329) );
  OAI211_X1 U22296 ( .C1(n19330), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19906), 
        .B(n19329), .ZN(n19331) );
  OAI211_X1 U22297 ( .C1(n19335), .C2(n19332), .A(n19761), .B(n19331), .ZN(
        n19354) );
  OAI21_X1 U22298 ( .B1(n10737), .B2(n19351), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19333) );
  OAI21_X1 U22299 ( .B1(n19335), .B2(n19334), .A(n19333), .ZN(n19353) );
  AOI22_X1 U22300 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19354), .B1(
        n19226), .B2(n19353), .ZN(n19336) );
  OAI211_X1 U22301 ( .C1(n19766), .C2(n19346), .A(n19337), .B(n19336), .ZN(
        P2_U3072) );
  AOI22_X1 U22302 ( .A1(n19671), .A2(n19384), .B1(n19351), .B2(n19767), .ZN(
        n19339) );
  AOI22_X1 U22303 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19354), .B1(
        n19234), .B2(n19353), .ZN(n19338) );
  OAI211_X1 U22304 ( .C1(n19674), .C2(n19346), .A(n19339), .B(n19338), .ZN(
        P2_U3073) );
  AOI22_X1 U22305 ( .A1(n19729), .A2(n19384), .B1(n19351), .B2(n19772), .ZN(
        n19341) );
  AOI22_X1 U22306 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19354), .B1(
        n19239), .B2(n19353), .ZN(n19340) );
  OAI211_X1 U22307 ( .C1(n19732), .C2(n19346), .A(n19341), .B(n19340), .ZN(
        P2_U3074) );
  AOI22_X1 U22308 ( .A1(n19779), .A2(n19384), .B1(n19351), .B2(n19777), .ZN(
        n19343) );
  AOI22_X1 U22309 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19354), .B1(
        n19778), .B2(n19353), .ZN(n19342) );
  OAI211_X1 U22310 ( .C1(n19782), .C2(n19346), .A(n19343), .B(n19342), .ZN(
        P2_U3075) );
  AOI22_X1 U22311 ( .A1(n19737), .A2(n19384), .B1(n19351), .B2(n19783), .ZN(
        n19345) );
  AOI22_X1 U22312 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19354), .B1(
        n19784), .B2(n19353), .ZN(n19344) );
  OAI211_X1 U22313 ( .C1(n19740), .C2(n19346), .A(n19345), .B(n19344), .ZN(
        P2_U3076) );
  INV_X1 U22314 ( .A(n19384), .ZN(n19362) );
  INV_X1 U22315 ( .A(n19346), .ZN(n19352) );
  AOI22_X1 U22316 ( .A1(n19352), .A2(n19791), .B1(n19351), .B2(n19789), .ZN(
        n19348) );
  AOI22_X1 U22317 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19354), .B1(
        n19790), .B2(n19353), .ZN(n19347) );
  OAI211_X1 U22318 ( .C1(n19794), .C2(n19362), .A(n19348), .B(n19347), .ZN(
        P2_U3077) );
  AOI22_X1 U22319 ( .A1(n19352), .A2(n19699), .B1(n19351), .B2(n19795), .ZN(
        n19350) );
  AOI22_X1 U22320 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19354), .B1(
        n19796), .B2(n19353), .ZN(n19349) );
  OAI211_X1 U22321 ( .C1(n19702), .C2(n19362), .A(n19350), .B(n19349), .ZN(
        P2_U3078) );
  AOI22_X1 U22322 ( .A1(n19352), .A2(n19807), .B1(n19351), .B2(n19803), .ZN(
        n19356) );
  AOI22_X1 U22323 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19354), .B1(
        n19805), .B2(n19353), .ZN(n19355) );
  OAI211_X1 U22324 ( .C1(n19813), .C2(n19362), .A(n19356), .B(n19355), .ZN(
        P2_U3079) );
  NOR2_X1 U22325 ( .A1(n19358), .A2(n19357), .ZN(n19614) );
  NAND2_X1 U22326 ( .A1(n19614), .A2(n19912), .ZN(n19361) );
  OR2_X1 U22327 ( .A1(n19361), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19360) );
  NAND3_X1 U22328 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19912), .A3(
        n19929), .ZN(n19393) );
  NOR2_X1 U22329 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19393), .ZN(
        n19382) );
  NOR3_X1 U22330 ( .A1(n19359), .A2(n19382), .A3(n19959), .ZN(n19363) );
  AOI21_X1 U22331 ( .B1(n19959), .B2(n19360), .A(n19363), .ZN(n19383) );
  AOI22_X1 U22332 ( .A1(n19383), .A2(n19226), .B1(n19755), .B2(n19382), .ZN(
        n19369) );
  INV_X1 U22333 ( .A(n19361), .ZN(n19367) );
  AOI21_X1 U22334 ( .B1(n19362), .B2(n19403), .A(n19553), .ZN(n19366) );
  INV_X1 U22335 ( .A(n19382), .ZN(n19364) );
  AOI211_X1 U22336 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19364), .A(n19618), 
        .B(n19363), .ZN(n19365) );
  AOI22_X1 U22337 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19385), .B1(
        n19384), .B2(n19714), .ZN(n19368) );
  OAI211_X1 U22338 ( .C1(n19726), .C2(n19403), .A(n19369), .B(n19368), .ZN(
        P2_U3080) );
  AOI22_X1 U22339 ( .A1(n19383), .A2(n19234), .B1(n19767), .B2(n19382), .ZN(
        n19371) );
  AOI22_X1 U22340 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19385), .B1(
        n19384), .B2(n19768), .ZN(n19370) );
  OAI211_X1 U22341 ( .C1(n19771), .C2(n19403), .A(n19371), .B(n19370), .ZN(
        P2_U3081) );
  AOI22_X1 U22342 ( .A1(n19383), .A2(n19239), .B1(n19772), .B2(n19382), .ZN(
        n19373) );
  AOI22_X1 U22343 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19385), .B1(
        n19384), .B2(n19773), .ZN(n19372) );
  OAI211_X1 U22344 ( .C1(n19776), .C2(n19403), .A(n19373), .B(n19372), .ZN(
        P2_U3082) );
  AOI22_X1 U22345 ( .A1(n19383), .A2(n19778), .B1(n19777), .B2(n19382), .ZN(
        n19375) );
  AOI22_X1 U22346 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19385), .B1(
        n19384), .B2(n19733), .ZN(n19374) );
  OAI211_X1 U22347 ( .C1(n19736), .C2(n19403), .A(n19375), .B(n19374), .ZN(
        P2_U3083) );
  AOI22_X1 U22348 ( .A1(n19383), .A2(n19784), .B1(n19783), .B2(n19382), .ZN(
        n19377) );
  AOI22_X1 U22349 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19385), .B1(
        n19384), .B2(n19785), .ZN(n19376) );
  OAI211_X1 U22350 ( .C1(n19788), .C2(n19403), .A(n19377), .B(n19376), .ZN(
        P2_U3084) );
  AOI22_X1 U22351 ( .A1(n19383), .A2(n19790), .B1(n19789), .B2(n19382), .ZN(
        n19379) );
  AOI22_X1 U22352 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19385), .B1(
        n19384), .B2(n19791), .ZN(n19378) );
  OAI211_X1 U22353 ( .C1(n19794), .C2(n19403), .A(n19379), .B(n19378), .ZN(
        P2_U3085) );
  AOI22_X1 U22354 ( .A1(n19383), .A2(n19796), .B1(n19795), .B2(n19382), .ZN(
        n19381) );
  AOI22_X1 U22355 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19385), .B1(
        n19384), .B2(n19699), .ZN(n19380) );
  OAI211_X1 U22356 ( .C1(n19702), .C2(n19403), .A(n19381), .B(n19380), .ZN(
        P2_U3086) );
  AOI22_X1 U22357 ( .A1(n19383), .A2(n19805), .B1(n19803), .B2(n19382), .ZN(
        n19387) );
  AOI22_X1 U22358 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19385), .B1(
        n19384), .B2(n19807), .ZN(n19386) );
  OAI211_X1 U22359 ( .C1(n19813), .C2(n19403), .A(n19387), .B(n19386), .ZN(
        P2_U3087) );
  NOR2_X1 U22360 ( .A1(n19939), .A2(n19393), .ZN(n19420) );
  AOI22_X1 U22361 ( .A1(n19763), .A2(n19440), .B1(n19420), .B2(n19755), .ZN(
        n19396) );
  OAI21_X1 U22362 ( .B1(n19907), .B2(n19651), .A(n19902), .ZN(n19394) );
  INV_X1 U22363 ( .A(n19393), .ZN(n19391) );
  OAI21_X1 U22364 ( .B1(n10742), .B2(n19959), .A(n19931), .ZN(n19389) );
  INV_X1 U22365 ( .A(n19420), .ZN(n19388) );
  AOI21_X1 U22366 ( .B1(n19389), .B2(n19388), .A(n19618), .ZN(n19390) );
  OAI21_X1 U22367 ( .B1(n19394), .B2(n19391), .A(n19390), .ZN(n19412) );
  OAI21_X1 U22368 ( .B1(n10742), .B2(n19420), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19392) );
  OAI21_X1 U22369 ( .B1(n19394), .B2(n19393), .A(n19392), .ZN(n19411) );
  AOI22_X1 U22370 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19412), .B1(
        n19226), .B2(n19411), .ZN(n19395) );
  OAI211_X1 U22371 ( .C1(n19766), .C2(n19403), .A(n19396), .B(n19395), .ZN(
        P2_U3088) );
  INV_X1 U22372 ( .A(n19403), .ZN(n19410) );
  AOI22_X1 U22373 ( .A1(n19410), .A2(n19768), .B1(n19767), .B2(n19420), .ZN(
        n19398) );
  AOI22_X1 U22374 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19412), .B1(
        n19234), .B2(n19411), .ZN(n19397) );
  OAI211_X1 U22375 ( .C1(n19771), .C2(n19437), .A(n19398), .B(n19397), .ZN(
        P2_U3089) );
  AOI22_X1 U22376 ( .A1(n19729), .A2(n19440), .B1(n19420), .B2(n19772), .ZN(
        n19400) );
  AOI22_X1 U22377 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19412), .B1(
        n19239), .B2(n19411), .ZN(n19399) );
  OAI211_X1 U22378 ( .C1(n19732), .C2(n19403), .A(n19400), .B(n19399), .ZN(
        P2_U3090) );
  AOI22_X1 U22379 ( .A1(n19779), .A2(n19440), .B1(n19420), .B2(n19777), .ZN(
        n19402) );
  AOI22_X1 U22380 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19412), .B1(
        n19778), .B2(n19411), .ZN(n19401) );
  OAI211_X1 U22381 ( .C1(n19782), .C2(n19403), .A(n19402), .B(n19401), .ZN(
        P2_U3091) );
  AOI22_X1 U22382 ( .A1(n19410), .A2(n19785), .B1(n19420), .B2(n19783), .ZN(
        n19405) );
  AOI22_X1 U22383 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19412), .B1(
        n19784), .B2(n19411), .ZN(n19404) );
  OAI211_X1 U22384 ( .C1(n19788), .C2(n19437), .A(n19405), .B(n19404), .ZN(
        P2_U3092) );
  AOI22_X1 U22385 ( .A1(n19410), .A2(n19791), .B1(n19420), .B2(n19789), .ZN(
        n19407) );
  AOI22_X1 U22386 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19412), .B1(
        n19790), .B2(n19411), .ZN(n19406) );
  OAI211_X1 U22387 ( .C1(n19794), .C2(n19437), .A(n19407), .B(n19406), .ZN(
        P2_U3093) );
  AOI22_X1 U22388 ( .A1(n19410), .A2(n19699), .B1(n19420), .B2(n19795), .ZN(
        n19409) );
  AOI22_X1 U22389 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19412), .B1(
        n19796), .B2(n19411), .ZN(n19408) );
  OAI211_X1 U22390 ( .C1(n19702), .C2(n19437), .A(n19409), .B(n19408), .ZN(
        P2_U3094) );
  AOI22_X1 U22391 ( .A1(n19410), .A2(n19807), .B1(n19420), .B2(n19803), .ZN(
        n19414) );
  AOI22_X1 U22392 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19412), .B1(
        n19805), .B2(n19411), .ZN(n19413) );
  OAI211_X1 U22393 ( .C1(n19813), .C2(n19437), .A(n19414), .B(n19413), .ZN(
        P2_U3095) );
  NAND2_X1 U22394 ( .A1(n19713), .A2(n19912), .ZN(n19453) );
  NOR2_X1 U22395 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19453), .ZN(
        n19438) );
  NOR2_X1 U22396 ( .A1(n19420), .A2(n19438), .ZN(n19416) );
  OR2_X1 U22397 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19416), .ZN(n19418) );
  NOR3_X1 U22398 ( .A1(n19417), .A2(n19438), .A3(n19959), .ZN(n19421) );
  AOI21_X1 U22399 ( .B1(n19959), .B2(n19418), .A(n19421), .ZN(n19439) );
  AOI22_X1 U22400 ( .A1(n19439), .A2(n19226), .B1(n19755), .B2(n19438), .ZN(
        n19424) );
  AOI21_X1 U22401 ( .B1(n19437), .B2(n19466), .A(n19553), .ZN(n19419) );
  AOI221_X1 U22402 ( .B1(n19931), .B2(n19420), .C1(n19931), .C2(n19419), .A(
        n19438), .ZN(n19422) );
  AOI22_X1 U22403 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19441), .B1(
        n19440), .B2(n19714), .ZN(n19423) );
  OAI211_X1 U22404 ( .C1(n19726), .C2(n19466), .A(n19424), .B(n19423), .ZN(
        P2_U3096) );
  AOI22_X1 U22405 ( .A1(n19439), .A2(n19234), .B1(n19767), .B2(n19438), .ZN(
        n19426) );
  AOI22_X1 U22406 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19441), .B1(
        n19440), .B2(n19768), .ZN(n19425) );
  OAI211_X1 U22407 ( .C1(n19771), .C2(n19466), .A(n19426), .B(n19425), .ZN(
        P2_U3097) );
  AOI22_X1 U22408 ( .A1(n19439), .A2(n19239), .B1(n19772), .B2(n19438), .ZN(
        n19428) );
  AOI22_X1 U22409 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19441), .B1(
        n19440), .B2(n19773), .ZN(n19427) );
  OAI211_X1 U22410 ( .C1(n19776), .C2(n19466), .A(n19428), .B(n19427), .ZN(
        P2_U3098) );
  AOI22_X1 U22411 ( .A1(n19439), .A2(n19778), .B1(n19777), .B2(n19438), .ZN(
        n19430) );
  AOI22_X1 U22412 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19441), .B1(
        n19440), .B2(n19733), .ZN(n19429) );
  OAI211_X1 U22413 ( .C1(n19736), .C2(n19466), .A(n19430), .B(n19429), .ZN(
        P2_U3099) );
  AOI22_X1 U22414 ( .A1(n19439), .A2(n19784), .B1(n19783), .B2(n19438), .ZN(
        n19432) );
  AOI22_X1 U22415 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19441), .B1(
        n19474), .B2(n19737), .ZN(n19431) );
  OAI211_X1 U22416 ( .C1(n19740), .C2(n19437), .A(n19432), .B(n19431), .ZN(
        P2_U3100) );
  AOI22_X1 U22417 ( .A1(n19439), .A2(n19790), .B1(n19789), .B2(n19438), .ZN(
        n19434) );
  AOI22_X1 U22418 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19441), .B1(
        n19440), .B2(n19791), .ZN(n19433) );
  OAI211_X1 U22419 ( .C1(n19794), .C2(n19466), .A(n19434), .B(n19433), .ZN(
        P2_U3101) );
  AOI22_X1 U22420 ( .A1(n19439), .A2(n19796), .B1(n19795), .B2(n19438), .ZN(
        n19436) );
  AOI22_X1 U22421 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19441), .B1(
        n19474), .B2(n19797), .ZN(n19435) );
  OAI211_X1 U22422 ( .C1(n19802), .C2(n19437), .A(n19436), .B(n19435), .ZN(
        P2_U3102) );
  AOI22_X1 U22423 ( .A1(n19439), .A2(n19805), .B1(n19803), .B2(n19438), .ZN(
        n19443) );
  AOI22_X1 U22424 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19441), .B1(
        n19440), .B2(n19807), .ZN(n19442) );
  OAI211_X1 U22425 ( .C1(n19813), .C2(n19466), .A(n19443), .B(n19442), .ZN(
        P2_U3103) );
  OAI21_X1 U22426 ( .B1(n19907), .B2(n19905), .A(n19453), .ZN(n19449) );
  NOR2_X1 U22427 ( .A1(n19939), .A2(n19453), .ZN(n19482) );
  INV_X1 U22428 ( .A(n19482), .ZN(n19444) );
  NAND2_X1 U22429 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19444), .ZN(n19445) );
  OR2_X1 U22430 ( .A1(n19446), .A2(n19445), .ZN(n19450) );
  OAI211_X1 U22431 ( .C1(n19931), .C2(n19482), .A(n19450), .B(n19761), .ZN(
        n19447) );
  INV_X1 U22432 ( .A(n19447), .ZN(n19448) );
  INV_X1 U22433 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n19457) );
  INV_X1 U22434 ( .A(n19450), .ZN(n19451) );
  AOI211_X2 U22435 ( .C1(n19453), .C2(n19959), .A(n19452), .B(n19451), .ZN(
        n19473) );
  AOI22_X1 U22436 ( .A1(n19473), .A2(n19226), .B1(n19755), .B2(n19482), .ZN(
        n19456) );
  NAND2_X1 U22437 ( .A1(n19756), .A2(n19454), .ZN(n19478) );
  AOI22_X1 U22438 ( .A1(n19474), .A2(n19714), .B1(n19512), .B2(n19763), .ZN(
        n19455) );
  OAI211_X1 U22439 ( .C1(n19472), .C2(n19457), .A(n19456), .B(n19455), .ZN(
        P2_U3104) );
  AOI22_X1 U22440 ( .A1(n19473), .A2(n19234), .B1(n19767), .B2(n19482), .ZN(
        n19459) );
  INV_X1 U22441 ( .A(n19472), .ZN(n19475) );
  AOI22_X1 U22442 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19475), .B1(
        n19512), .B2(n19671), .ZN(n19458) );
  OAI211_X1 U22443 ( .C1(n19674), .C2(n19466), .A(n19459), .B(n19458), .ZN(
        P2_U3105) );
  AOI22_X1 U22444 ( .A1(n19473), .A2(n19239), .B1(n19772), .B2(n19482), .ZN(
        n19461) );
  AOI22_X1 U22445 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19475), .B1(
        n19512), .B2(n19729), .ZN(n19460) );
  OAI211_X1 U22446 ( .C1(n19732), .C2(n19466), .A(n19461), .B(n19460), .ZN(
        P2_U3106) );
  AOI22_X1 U22447 ( .A1(n19473), .A2(n19778), .B1(n19777), .B2(n19482), .ZN(
        n19463) );
  AOI22_X1 U22448 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19475), .B1(
        n19512), .B2(n19779), .ZN(n19462) );
  OAI211_X1 U22449 ( .C1(n19782), .C2(n19466), .A(n19463), .B(n19462), .ZN(
        P2_U3107) );
  AOI22_X1 U22450 ( .A1(n19473), .A2(n19784), .B1(n19783), .B2(n19482), .ZN(
        n19465) );
  AOI22_X1 U22451 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19475), .B1(
        n19512), .B2(n19737), .ZN(n19464) );
  OAI211_X1 U22452 ( .C1(n19740), .C2(n19466), .A(n19465), .B(n19464), .ZN(
        P2_U3108) );
  AOI22_X1 U22453 ( .A1(n19473), .A2(n19790), .B1(n19789), .B2(n19482), .ZN(
        n19468) );
  AOI22_X1 U22454 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19475), .B1(
        n19474), .B2(n19791), .ZN(n19467) );
  OAI211_X1 U22455 ( .C1(n19794), .C2(n19478), .A(n19468), .B(n19467), .ZN(
        P2_U3109) );
  INV_X1 U22456 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n19471) );
  AOI22_X1 U22457 ( .A1(n19473), .A2(n19796), .B1(n19795), .B2(n19482), .ZN(
        n19470) );
  AOI22_X1 U22458 ( .A1(n19474), .A2(n19699), .B1(n19512), .B2(n19797), .ZN(
        n19469) );
  OAI211_X1 U22459 ( .C1(n19472), .C2(n19471), .A(n19470), .B(n19469), .ZN(
        P2_U3110) );
  AOI22_X1 U22460 ( .A1(n19473), .A2(n19805), .B1(n19803), .B2(n19482), .ZN(
        n19477) );
  AOI22_X1 U22461 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19475), .B1(
        n19474), .B2(n19807), .ZN(n19476) );
  OAI211_X1 U22462 ( .C1(n19813), .C2(n19478), .A(n19477), .B(n19476), .ZN(
        P2_U3111) );
  INV_X1 U22463 ( .A(n19712), .ZN(n19480) );
  NOR3_X1 U22464 ( .A1(n19544), .A2(n19906), .A3(n19512), .ZN(n19481) );
  AND2_X1 U22465 ( .A1(n19902), .A2(n19553), .ZN(n19901) );
  NOR2_X1 U22466 ( .A1(n19481), .A2(n19901), .ZN(n19487) );
  INV_X1 U22467 ( .A(n19487), .ZN(n19484) );
  NOR2_X1 U22468 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19912), .ZN(
        n19580) );
  NAND2_X1 U22469 ( .A1(n19580), .A2(n19929), .ZN(n19527) );
  NOR2_X1 U22470 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19527), .ZN(
        n19510) );
  NOR2_X1 U22471 ( .A1(n19510), .A2(n19482), .ZN(n19485) );
  AOI211_X1 U22472 ( .C1(n10749), .C2(n19931), .A(n19902), .B(n19510), .ZN(
        n19483) );
  INV_X1 U22473 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n19490) );
  AOI22_X1 U22474 ( .A1(n19544), .A2(n19763), .B1(n19755), .B2(n19510), .ZN(
        n19489) );
  OAI21_X1 U22475 ( .B1(n10749), .B2(n19510), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19486) );
  AOI22_X1 U22476 ( .A1(n19487), .A2(n19486), .B1(n19485), .B2(n19959), .ZN(
        n19513) );
  AOI22_X1 U22477 ( .A1(n19226), .A2(n19513), .B1(n19512), .B2(n19714), .ZN(
        n19488) );
  OAI211_X1 U22478 ( .C1(n19517), .C2(n19490), .A(n19489), .B(n19488), .ZN(
        P2_U3112) );
  INV_X1 U22479 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n19493) );
  AOI22_X1 U22480 ( .A1(n19544), .A2(n19671), .B1(n19767), .B2(n19510), .ZN(
        n19492) );
  AOI22_X1 U22481 ( .A1(n19234), .A2(n19513), .B1(n19512), .B2(n19768), .ZN(
        n19491) );
  OAI211_X1 U22482 ( .C1(n19517), .C2(n19493), .A(n19492), .B(n19491), .ZN(
        P2_U3113) );
  INV_X1 U22483 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n19496) );
  AOI22_X1 U22484 ( .A1(n19544), .A2(n19729), .B1(n19772), .B2(n19510), .ZN(
        n19495) );
  AOI22_X1 U22485 ( .A1(n19239), .A2(n19513), .B1(n19512), .B2(n19773), .ZN(
        n19494) );
  OAI211_X1 U22486 ( .C1(n19517), .C2(n19496), .A(n19495), .B(n19494), .ZN(
        P2_U3114) );
  INV_X1 U22487 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n19499) );
  AOI22_X1 U22488 ( .A1(n19544), .A2(n19779), .B1(n19777), .B2(n19510), .ZN(
        n19498) );
  AOI22_X1 U22489 ( .A1(n19778), .A2(n19513), .B1(n19512), .B2(n19733), .ZN(
        n19497) );
  OAI211_X1 U22490 ( .C1(n19517), .C2(n19499), .A(n19498), .B(n19497), .ZN(
        P2_U3115) );
  INV_X1 U22491 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n19502) );
  AOI22_X1 U22492 ( .A1(n19544), .A2(n19737), .B1(n19783), .B2(n19510), .ZN(
        n19501) );
  AOI22_X1 U22493 ( .A1(n19784), .A2(n19513), .B1(n19512), .B2(n19785), .ZN(
        n19500) );
  OAI211_X1 U22494 ( .C1(n19517), .C2(n19502), .A(n19501), .B(n19500), .ZN(
        P2_U3116) );
  INV_X1 U22495 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n19506) );
  INV_X1 U22496 ( .A(n19794), .ZN(n19503) );
  AOI22_X1 U22497 ( .A1(n19544), .A2(n19503), .B1(n19789), .B2(n19510), .ZN(
        n19505) );
  AOI22_X1 U22498 ( .A1(n19790), .A2(n19513), .B1(n19512), .B2(n19791), .ZN(
        n19504) );
  OAI211_X1 U22499 ( .C1(n19517), .C2(n19506), .A(n19505), .B(n19504), .ZN(
        P2_U3117) );
  AOI22_X1 U22500 ( .A1(n19544), .A2(n19797), .B1(n19795), .B2(n19510), .ZN(
        n19508) );
  AOI22_X1 U22501 ( .A1(n19796), .A2(n19513), .B1(n19512), .B2(n19699), .ZN(
        n19507) );
  OAI211_X1 U22502 ( .C1(n19517), .C2(n19509), .A(n19508), .B(n19507), .ZN(
        P2_U3118) );
  INV_X1 U22503 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n19516) );
  INV_X1 U22504 ( .A(n19813), .ZN(n19511) );
  AOI22_X1 U22505 ( .A1(n19544), .A2(n19511), .B1(n19803), .B2(n19510), .ZN(
        n19515) );
  AOI22_X1 U22506 ( .A1(n19805), .A2(n19513), .B1(n19512), .B2(n19807), .ZN(
        n19514) );
  OAI211_X1 U22507 ( .C1(n19517), .C2(n19516), .A(n19515), .B(n19514), .ZN(
        P2_U3119) );
  INV_X1 U22508 ( .A(n19544), .ZN(n19535) );
  INV_X1 U22509 ( .A(n19580), .ZN(n19586) );
  NOR2_X1 U22510 ( .A1(n19518), .A2(n19586), .ZN(n19555) );
  AOI22_X1 U22511 ( .A1(n19576), .A2(n19763), .B1(n19755), .B2(n19555), .ZN(
        n19530) );
  NAND2_X1 U22512 ( .A1(n19519), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19660) );
  OAI21_X1 U22513 ( .B1(n19660), .B2(n19520), .A(n19902), .ZN(n19528) );
  INV_X1 U22514 ( .A(n19527), .ZN(n19524) );
  INV_X1 U22515 ( .A(n19525), .ZN(n19522) );
  INV_X1 U22516 ( .A(n19555), .ZN(n19521) );
  OAI211_X1 U22517 ( .C1(n19522), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19906), 
        .B(n19521), .ZN(n19523) );
  OAI211_X1 U22518 ( .C1(n19528), .C2(n19524), .A(n19761), .B(n19523), .ZN(
        n19546) );
  OAI21_X1 U22519 ( .B1(n19525), .B2(n19555), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19526) );
  OAI21_X1 U22520 ( .B1(n19528), .B2(n19527), .A(n19526), .ZN(n19545) );
  AOI22_X1 U22521 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19546), .B1(
        n19226), .B2(n19545), .ZN(n19529) );
  OAI211_X1 U22522 ( .C1(n19766), .C2(n19535), .A(n19530), .B(n19529), .ZN(
        P2_U3120) );
  AOI22_X1 U22523 ( .A1(n19576), .A2(n19671), .B1(n19767), .B2(n19555), .ZN(
        n19532) );
  AOI22_X1 U22524 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19546), .B1(
        n19234), .B2(n19545), .ZN(n19531) );
  OAI211_X1 U22525 ( .C1(n19674), .C2(n19535), .A(n19532), .B(n19531), .ZN(
        P2_U3121) );
  AOI22_X1 U22526 ( .A1(n19576), .A2(n19729), .B1(n19772), .B2(n19555), .ZN(
        n19534) );
  AOI22_X1 U22527 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19546), .B1(
        n19239), .B2(n19545), .ZN(n19533) );
  OAI211_X1 U22528 ( .C1(n19732), .C2(n19535), .A(n19534), .B(n19533), .ZN(
        P2_U3122) );
  AOI22_X1 U22529 ( .A1(n19544), .A2(n19733), .B1(n19777), .B2(n19555), .ZN(
        n19537) );
  AOI22_X1 U22530 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19546), .B1(
        n19778), .B2(n19545), .ZN(n19536) );
  OAI211_X1 U22531 ( .C1(n19736), .C2(n19554), .A(n19537), .B(n19536), .ZN(
        P2_U3123) );
  AOI22_X1 U22532 ( .A1(n19544), .A2(n19785), .B1(n19783), .B2(n19555), .ZN(
        n19539) );
  AOI22_X1 U22533 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19546), .B1(
        n19784), .B2(n19545), .ZN(n19538) );
  OAI211_X1 U22534 ( .C1(n19788), .C2(n19554), .A(n19539), .B(n19538), .ZN(
        P2_U3124) );
  AOI22_X1 U22535 ( .A1(n19544), .A2(n19791), .B1(n19789), .B2(n19555), .ZN(
        n19541) );
  AOI22_X1 U22536 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19546), .B1(
        n19790), .B2(n19545), .ZN(n19540) );
  OAI211_X1 U22537 ( .C1(n19794), .C2(n19554), .A(n19541), .B(n19540), .ZN(
        P2_U3125) );
  AOI22_X1 U22538 ( .A1(n19544), .A2(n19699), .B1(n19795), .B2(n19555), .ZN(
        n19543) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19546), .B1(
        n19796), .B2(n19545), .ZN(n19542) );
  OAI211_X1 U22540 ( .C1(n19702), .C2(n19554), .A(n19543), .B(n19542), .ZN(
        P2_U3126) );
  AOI22_X1 U22541 ( .A1(n19544), .A2(n19807), .B1(n19803), .B2(n19555), .ZN(
        n19548) );
  AOI22_X1 U22542 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19546), .B1(
        n19805), .B2(n19545), .ZN(n19547) );
  OAI211_X1 U22543 ( .C1(n19813), .C2(n19554), .A(n19548), .B(n19547), .ZN(
        P2_U3127) );
  AND2_X1 U22544 ( .A1(n19549), .A2(n19580), .ZN(n19574) );
  OAI21_X1 U22545 ( .B1(n19552), .B2(n19574), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19550) );
  OAI21_X1 U22546 ( .B1(n19586), .B2(n19551), .A(n19550), .ZN(n19575) );
  AOI22_X1 U22547 ( .A1(n19575), .A2(n19226), .B1(n19755), .B2(n19574), .ZN(
        n19561) );
  INV_X1 U22548 ( .A(n19552), .ZN(n19558) );
  AOI21_X1 U22549 ( .B1(n19554), .B2(n19600), .A(n19553), .ZN(n19556) );
  NOR2_X1 U22550 ( .A1(n19556), .A2(n19555), .ZN(n19557) );
  AOI211_X1 U22551 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19558), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19557), .ZN(n19559) );
  OAI21_X1 U22552 ( .B1(n19559), .B2(n19574), .A(n19761), .ZN(n19577) );
  AOI22_X1 U22553 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19577), .B1(
        n19576), .B2(n19714), .ZN(n19560) );
  OAI211_X1 U22554 ( .C1(n19726), .C2(n19600), .A(n19561), .B(n19560), .ZN(
        P2_U3128) );
  AOI22_X1 U22555 ( .A1(n19575), .A2(n19234), .B1(n19767), .B2(n19574), .ZN(
        n19563) );
  AOI22_X1 U22556 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19577), .B1(
        n19576), .B2(n19768), .ZN(n19562) );
  OAI211_X1 U22557 ( .C1(n19771), .C2(n19600), .A(n19563), .B(n19562), .ZN(
        P2_U3129) );
  AOI22_X1 U22558 ( .A1(n19575), .A2(n19239), .B1(n19772), .B2(n19574), .ZN(
        n19565) );
  AOI22_X1 U22559 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19577), .B1(
        n19576), .B2(n19773), .ZN(n19564) );
  OAI211_X1 U22560 ( .C1(n19776), .C2(n19600), .A(n19565), .B(n19564), .ZN(
        P2_U3130) );
  AOI22_X1 U22561 ( .A1(n19575), .A2(n19778), .B1(n19777), .B2(n19574), .ZN(
        n19567) );
  AOI22_X1 U22562 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19577), .B1(
        n19576), .B2(n19733), .ZN(n19566) );
  OAI211_X1 U22563 ( .C1(n19736), .C2(n19600), .A(n19567), .B(n19566), .ZN(
        P2_U3131) );
  AOI22_X1 U22564 ( .A1(n19575), .A2(n19784), .B1(n19783), .B2(n19574), .ZN(
        n19569) );
  AOI22_X1 U22565 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19577), .B1(
        n19576), .B2(n19785), .ZN(n19568) );
  OAI211_X1 U22566 ( .C1(n19788), .C2(n19600), .A(n19569), .B(n19568), .ZN(
        P2_U3132) );
  AOI22_X1 U22567 ( .A1(n19575), .A2(n19790), .B1(n19789), .B2(n19574), .ZN(
        n19571) );
  AOI22_X1 U22568 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19577), .B1(
        n19576), .B2(n19791), .ZN(n19570) );
  OAI211_X1 U22569 ( .C1(n19794), .C2(n19600), .A(n19571), .B(n19570), .ZN(
        P2_U3133) );
  AOI22_X1 U22570 ( .A1(n19575), .A2(n19796), .B1(n19795), .B2(n19574), .ZN(
        n19573) );
  AOI22_X1 U22571 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19577), .B1(
        n19576), .B2(n19699), .ZN(n19572) );
  OAI211_X1 U22572 ( .C1(n19702), .C2(n19600), .A(n19573), .B(n19572), .ZN(
        P2_U3134) );
  AOI22_X1 U22573 ( .A1(n19575), .A2(n19805), .B1(n19803), .B2(n19574), .ZN(
        n19579) );
  AOI22_X1 U22574 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19577), .B1(
        n19576), .B2(n19807), .ZN(n19578) );
  OAI211_X1 U22575 ( .C1(n19813), .C2(n19600), .A(n19579), .B(n19578), .ZN(
        P2_U3135) );
  NAND2_X1 U22576 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19580), .ZN(
        n19583) );
  NOR2_X1 U22577 ( .A1(n19581), .A2(n19586), .ZN(n19605) );
  OAI21_X1 U22578 ( .B1(n19584), .B2(n19605), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19582) );
  OAI21_X1 U22579 ( .B1(n19583), .B2(n19906), .A(n19582), .ZN(n19606) );
  AOI22_X1 U22580 ( .A1(n19606), .A2(n19226), .B1(n19755), .B2(n19605), .ZN(
        n19591) );
  INV_X1 U22581 ( .A(n19584), .ZN(n19585) );
  AOI21_X1 U22582 ( .B1(n19585), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19588) );
  OAI22_X1 U22583 ( .A1(n19660), .A2(n19589), .B1(n19586), .B2(n19929), .ZN(
        n19587) );
  OAI211_X1 U22584 ( .C1(n19605), .C2(n19588), .A(n19587), .B(n19761), .ZN(
        n19608) );
  NOR2_X2 U22585 ( .A1(n19652), .A2(n19589), .ZN(n19647) );
  AOI22_X1 U22586 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19608), .B1(
        n19647), .B2(n19763), .ZN(n19590) );
  OAI211_X1 U22587 ( .C1(n19766), .C2(n19600), .A(n19591), .B(n19590), .ZN(
        P2_U3136) );
  AOI22_X1 U22588 ( .A1(n19606), .A2(n19234), .B1(n19767), .B2(n19605), .ZN(
        n19593) );
  AOI22_X1 U22589 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19608), .B1(
        n19647), .B2(n19671), .ZN(n19592) );
  OAI211_X1 U22590 ( .C1(n19674), .C2(n19600), .A(n19593), .B(n19592), .ZN(
        P2_U3137) );
  AOI22_X1 U22591 ( .A1(n19606), .A2(n19239), .B1(n19772), .B2(n19605), .ZN(
        n19595) );
  AOI22_X1 U22592 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19608), .B1(
        n19647), .B2(n19729), .ZN(n19594) );
  OAI211_X1 U22593 ( .C1(n19732), .C2(n19600), .A(n19595), .B(n19594), .ZN(
        P2_U3138) );
  AOI22_X1 U22594 ( .A1(n19606), .A2(n19778), .B1(n19777), .B2(n19605), .ZN(
        n19597) );
  AOI22_X1 U22595 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19608), .B1(
        n19647), .B2(n19779), .ZN(n19596) );
  OAI211_X1 U22596 ( .C1(n19782), .C2(n19600), .A(n19597), .B(n19596), .ZN(
        P2_U3139) );
  AOI22_X1 U22597 ( .A1(n19606), .A2(n19784), .B1(n19783), .B2(n19605), .ZN(
        n19599) );
  AOI22_X1 U22598 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19608), .B1(
        n19647), .B2(n19737), .ZN(n19598) );
  OAI211_X1 U22599 ( .C1(n19740), .C2(n19600), .A(n19599), .B(n19598), .ZN(
        P2_U3140) );
  INV_X1 U22600 ( .A(n19647), .ZN(n19611) );
  AOI22_X1 U22601 ( .A1(n19606), .A2(n19790), .B1(n19789), .B2(n19605), .ZN(
        n19602) );
  INV_X1 U22602 ( .A(n19600), .ZN(n19607) );
  AOI22_X1 U22603 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19608), .B1(
        n19607), .B2(n19791), .ZN(n19601) );
  OAI211_X1 U22604 ( .C1(n19794), .C2(n19611), .A(n19602), .B(n19601), .ZN(
        P2_U3141) );
  AOI22_X1 U22605 ( .A1(n19606), .A2(n19796), .B1(n19795), .B2(n19605), .ZN(
        n19604) );
  AOI22_X1 U22606 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19608), .B1(
        n19607), .B2(n19699), .ZN(n19603) );
  OAI211_X1 U22607 ( .C1(n19702), .C2(n19611), .A(n19604), .B(n19603), .ZN(
        P2_U3142) );
  AOI22_X1 U22608 ( .A1(n19606), .A2(n19805), .B1(n19803), .B2(n19605), .ZN(
        n19610) );
  AOI22_X1 U22609 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19608), .B1(
        n19607), .B2(n19807), .ZN(n19609) );
  OAI211_X1 U22610 ( .C1(n19813), .C2(n19611), .A(n19610), .B(n19609), .ZN(
        P2_U3143) );
  NAND3_X1 U22611 ( .A1(n19929), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19663) );
  NOR2_X1 U22612 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19663), .ZN(
        n19623) );
  INV_X1 U22613 ( .A(n19623), .ZN(n19644) );
  NAND2_X1 U22614 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19644), .ZN(n19612) );
  NOR2_X1 U22615 ( .A1(n19613), .A2(n19612), .ZN(n19619) );
  NAND2_X1 U22616 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19614), .ZN(
        n19620) );
  OAI21_X1 U22617 ( .B1(n19620), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19959), 
        .ZN(n19615) );
  INV_X1 U22618 ( .A(n19615), .ZN(n19616) );
  OR2_X1 U22619 ( .A1(n19619), .A2(n19616), .ZN(n19645) );
  INV_X1 U22620 ( .A(n19226), .ZN(n19658) );
  INV_X1 U22621 ( .A(n19755), .ZN(n19657) );
  OAI22_X1 U22622 ( .A1(n19645), .A2(n19658), .B1(n19657), .B2(n19644), .ZN(
        n19617) );
  INV_X1 U22623 ( .A(n19617), .ZN(n19625) );
  OAI21_X1 U22624 ( .B1(n19647), .B2(n19708), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19621) );
  AOI211_X1 U22625 ( .C1(n19621), .C2(n19620), .A(n19619), .B(n19618), .ZN(
        n19622) );
  AOI22_X1 U22626 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19648), .B1(
        n19647), .B2(n19714), .ZN(n19624) );
  OAI211_X1 U22627 ( .C1(n19726), .C2(n19690), .A(n19625), .B(n19624), .ZN(
        P2_U3144) );
  INV_X1 U22628 ( .A(n19234), .ZN(n19669) );
  INV_X1 U22629 ( .A(n19767), .ZN(n19668) );
  OAI22_X1 U22630 ( .A1(n19645), .A2(n19669), .B1(n19668), .B2(n19644), .ZN(
        n19626) );
  INV_X1 U22631 ( .A(n19626), .ZN(n19628) );
  AOI22_X1 U22632 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19648), .B1(
        n19647), .B2(n19768), .ZN(n19627) );
  OAI211_X1 U22633 ( .C1(n19771), .C2(n19690), .A(n19628), .B(n19627), .ZN(
        P2_U3145) );
  INV_X1 U22634 ( .A(n19239), .ZN(n19676) );
  INV_X1 U22635 ( .A(n19772), .ZN(n19675) );
  OAI22_X1 U22636 ( .A1(n19645), .A2(n19676), .B1(n19675), .B2(n19644), .ZN(
        n19629) );
  INV_X1 U22637 ( .A(n19629), .ZN(n19631) );
  AOI22_X1 U22638 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19648), .B1(
        n19647), .B2(n19773), .ZN(n19630) );
  OAI211_X1 U22639 ( .C1(n19776), .C2(n19690), .A(n19631), .B(n19630), .ZN(
        P2_U3146) );
  INV_X1 U22640 ( .A(n19778), .ZN(n19681) );
  INV_X1 U22641 ( .A(n19777), .ZN(n19680) );
  OAI22_X1 U22642 ( .A1(n19645), .A2(n19681), .B1(n19680), .B2(n19644), .ZN(
        n19632) );
  INV_X1 U22643 ( .A(n19632), .ZN(n19634) );
  AOI22_X1 U22644 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19648), .B1(
        n19647), .B2(n19733), .ZN(n19633) );
  OAI211_X1 U22645 ( .C1(n19736), .C2(n19690), .A(n19634), .B(n19633), .ZN(
        P2_U3147) );
  INV_X1 U22646 ( .A(n19784), .ZN(n19686) );
  INV_X1 U22647 ( .A(n19783), .ZN(n19685) );
  OAI22_X1 U22648 ( .A1(n19645), .A2(n19686), .B1(n19685), .B2(n19644), .ZN(
        n19635) );
  INV_X1 U22649 ( .A(n19635), .ZN(n19637) );
  AOI22_X1 U22650 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19648), .B1(
        n19647), .B2(n19785), .ZN(n19636) );
  OAI211_X1 U22651 ( .C1(n19788), .C2(n19690), .A(n19637), .B(n19636), .ZN(
        P2_U3148) );
  INV_X1 U22652 ( .A(n19790), .ZN(n19692) );
  INV_X1 U22653 ( .A(n19789), .ZN(n19691) );
  OAI22_X1 U22654 ( .A1(n19645), .A2(n19692), .B1(n19691), .B2(n19644), .ZN(
        n19638) );
  INV_X1 U22655 ( .A(n19638), .ZN(n19640) );
  AOI22_X1 U22656 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19648), .B1(
        n19647), .B2(n19791), .ZN(n19639) );
  OAI211_X1 U22657 ( .C1(n19794), .C2(n19690), .A(n19640), .B(n19639), .ZN(
        P2_U3149) );
  INV_X1 U22658 ( .A(n19796), .ZN(n19697) );
  INV_X1 U22659 ( .A(n19795), .ZN(n19696) );
  OAI22_X1 U22660 ( .A1(n19645), .A2(n19697), .B1(n19696), .B2(n19644), .ZN(
        n19641) );
  INV_X1 U22661 ( .A(n19641), .ZN(n19643) );
  AOI22_X1 U22662 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19648), .B1(
        n19647), .B2(n19699), .ZN(n19642) );
  OAI211_X1 U22663 ( .C1(n19702), .C2(n19690), .A(n19643), .B(n19642), .ZN(
        P2_U3150) );
  INV_X1 U22664 ( .A(n19805), .ZN(n19705) );
  INV_X1 U22665 ( .A(n19803), .ZN(n19704) );
  OAI22_X1 U22666 ( .A1(n19645), .A2(n19705), .B1(n19704), .B2(n19644), .ZN(
        n19646) );
  INV_X1 U22667 ( .A(n19646), .ZN(n19650) );
  AOI22_X1 U22668 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19648), .B1(
        n19647), .B2(n19807), .ZN(n19649) );
  OAI211_X1 U22669 ( .C1(n19813), .C2(n19690), .A(n19650), .B(n19649), .ZN(
        P2_U3151) );
  NOR2_X1 U22670 ( .A1(n19939), .A2(n19663), .ZN(n19716) );
  INV_X1 U22671 ( .A(n19716), .ZN(n19703) );
  NAND2_X1 U22672 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19703), .ZN(n19653) );
  NOR2_X1 U22673 ( .A1(n19654), .A2(n19653), .ZN(n19662) );
  INV_X1 U22674 ( .A(n19663), .ZN(n19655) );
  AOI21_X1 U22675 ( .B1(n19931), .B2(n19655), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19656) );
  OAI22_X1 U22676 ( .A1(n19706), .A2(n19658), .B1(n19657), .B2(n19703), .ZN(
        n19659) );
  INV_X1 U22677 ( .A(n19659), .ZN(n19667) );
  INV_X1 U22678 ( .A(n19660), .ZN(n19757) );
  NAND2_X1 U22679 ( .A1(n19757), .A2(n19661), .ZN(n19664) );
  AOI21_X1 U22680 ( .B1(n19664), .B2(n19663), .A(n19662), .ZN(n19665) );
  OAI211_X1 U22681 ( .C1(n19716), .C2(n19931), .A(n19665), .B(n19761), .ZN(
        n19709) );
  AOI22_X1 U22682 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n19714), .ZN(n19666) );
  OAI211_X1 U22683 ( .C1(n19726), .C2(n19745), .A(n19667), .B(n19666), .ZN(
        P2_U3152) );
  OAI22_X1 U22684 ( .A1(n19706), .A2(n19669), .B1(n19668), .B2(n19703), .ZN(
        n19670) );
  INV_X1 U22685 ( .A(n19670), .ZN(n19673) );
  AOI22_X1 U22686 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19709), .B1(
        n19747), .B2(n19671), .ZN(n19672) );
  OAI211_X1 U22687 ( .C1(n19674), .C2(n19690), .A(n19673), .B(n19672), .ZN(
        P2_U3153) );
  OAI22_X1 U22688 ( .A1(n19706), .A2(n19676), .B1(n19675), .B2(n19703), .ZN(
        n19677) );
  INV_X1 U22689 ( .A(n19677), .ZN(n19679) );
  AOI22_X1 U22690 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19709), .B1(
        n19747), .B2(n19729), .ZN(n19678) );
  OAI211_X1 U22691 ( .C1(n19732), .C2(n19690), .A(n19679), .B(n19678), .ZN(
        P2_U3154) );
  OAI22_X1 U22692 ( .A1(n19706), .A2(n19681), .B1(n19680), .B2(n19703), .ZN(
        n19682) );
  INV_X1 U22693 ( .A(n19682), .ZN(n19684) );
  AOI22_X1 U22694 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19709), .B1(
        n19747), .B2(n19779), .ZN(n19683) );
  OAI211_X1 U22695 ( .C1(n19782), .C2(n19690), .A(n19684), .B(n19683), .ZN(
        P2_U3155) );
  OAI22_X1 U22696 ( .A1(n19706), .A2(n19686), .B1(n19685), .B2(n19703), .ZN(
        n19687) );
  INV_X1 U22697 ( .A(n19687), .ZN(n19689) );
  AOI22_X1 U22698 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19709), .B1(
        n19747), .B2(n19737), .ZN(n19688) );
  OAI211_X1 U22699 ( .C1(n19740), .C2(n19690), .A(n19689), .B(n19688), .ZN(
        P2_U3156) );
  OAI22_X1 U22700 ( .A1(n19706), .A2(n19692), .B1(n19691), .B2(n19703), .ZN(
        n19693) );
  INV_X1 U22701 ( .A(n19693), .ZN(n19695) );
  AOI22_X1 U22702 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n19791), .ZN(n19694) );
  OAI211_X1 U22703 ( .C1(n19794), .C2(n19745), .A(n19695), .B(n19694), .ZN(
        P2_U3157) );
  OAI22_X1 U22704 ( .A1(n19706), .A2(n19697), .B1(n19696), .B2(n19703), .ZN(
        n19698) );
  INV_X1 U22705 ( .A(n19698), .ZN(n19701) );
  AOI22_X1 U22706 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n19699), .ZN(n19700) );
  OAI211_X1 U22707 ( .C1(n19702), .C2(n19745), .A(n19701), .B(n19700), .ZN(
        P2_U3158) );
  OAI22_X1 U22708 ( .A1(n19706), .A2(n19705), .B1(n19704), .B2(n19703), .ZN(
        n19707) );
  INV_X1 U22709 ( .A(n19707), .ZN(n19711) );
  AOI22_X1 U22710 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n19807), .ZN(n19710) );
  OAI211_X1 U22711 ( .C1(n19813), .C2(n19745), .A(n19711), .B(n19710), .ZN(
        P2_U3159) );
  NAND2_X1 U22712 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19713), .ZN(
        n19759) );
  NOR2_X1 U22713 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19759), .ZN(
        n19746) );
  AOI22_X1 U22714 ( .A1(n19747), .A2(n19714), .B1(n19755), .B2(n19746), .ZN(
        n19725) );
  NOR3_X1 U22715 ( .A1(n19808), .A2(n19747), .A3(n19906), .ZN(n19715) );
  NOR2_X1 U22716 ( .A1(n19715), .A2(n19901), .ZN(n19723) );
  NOR2_X1 U22717 ( .A1(n19746), .A2(n19716), .ZN(n19722) );
  INV_X1 U22718 ( .A(n19722), .ZN(n19720) );
  INV_X1 U22719 ( .A(n10750), .ZN(n19718) );
  INV_X1 U22720 ( .A(n19746), .ZN(n19717) );
  OAI211_X1 U22721 ( .C1(n19718), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19906), 
        .B(n19717), .ZN(n19719) );
  OAI211_X1 U22722 ( .C1(n19723), .C2(n19720), .A(n19761), .B(n19719), .ZN(
        n19749) );
  OAI21_X1 U22723 ( .B1(n10750), .B2(n19746), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19721) );
  AOI22_X1 U22724 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19749), .B1(
        n19226), .B2(n19748), .ZN(n19724) );
  OAI211_X1 U22725 ( .C1(n19726), .C2(n19801), .A(n19725), .B(n19724), .ZN(
        P2_U3160) );
  AOI22_X1 U22726 ( .A1(n19747), .A2(n19768), .B1(n19767), .B2(n19746), .ZN(
        n19728) );
  AOI22_X1 U22727 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19749), .B1(
        n19234), .B2(n19748), .ZN(n19727) );
  OAI211_X1 U22728 ( .C1(n19771), .C2(n19801), .A(n19728), .B(n19727), .ZN(
        P2_U3161) );
  AOI22_X1 U22729 ( .A1(n19808), .A2(n19729), .B1(n19772), .B2(n19746), .ZN(
        n19731) );
  AOI22_X1 U22730 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19749), .B1(
        n19239), .B2(n19748), .ZN(n19730) );
  OAI211_X1 U22731 ( .C1(n19732), .C2(n19745), .A(n19731), .B(n19730), .ZN(
        P2_U3162) );
  AOI22_X1 U22732 ( .A1(n19747), .A2(n19733), .B1(n19777), .B2(n19746), .ZN(
        n19735) );
  AOI22_X1 U22733 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19749), .B1(
        n19778), .B2(n19748), .ZN(n19734) );
  OAI211_X1 U22734 ( .C1(n19736), .C2(n19801), .A(n19735), .B(n19734), .ZN(
        P2_U3163) );
  AOI22_X1 U22735 ( .A1(n19808), .A2(n19737), .B1(n19783), .B2(n19746), .ZN(
        n19739) );
  AOI22_X1 U22736 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19749), .B1(
        n19784), .B2(n19748), .ZN(n19738) );
  OAI211_X1 U22737 ( .C1(n19740), .C2(n19745), .A(n19739), .B(n19738), .ZN(
        P2_U3164) );
  AOI22_X1 U22738 ( .A1(n19747), .A2(n19791), .B1(n19789), .B2(n19746), .ZN(
        n19742) );
  AOI22_X1 U22739 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19749), .B1(
        n19790), .B2(n19748), .ZN(n19741) );
  OAI211_X1 U22740 ( .C1(n19794), .C2(n19801), .A(n19742), .B(n19741), .ZN(
        P2_U3165) );
  AOI22_X1 U22741 ( .A1(n19808), .A2(n19797), .B1(n19795), .B2(n19746), .ZN(
        n19744) );
  AOI22_X1 U22742 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19749), .B1(
        n19796), .B2(n19748), .ZN(n19743) );
  OAI211_X1 U22743 ( .C1(n19802), .C2(n19745), .A(n19744), .B(n19743), .ZN(
        P2_U3166) );
  AOI22_X1 U22744 ( .A1(n19747), .A2(n19807), .B1(n19803), .B2(n19746), .ZN(
        n19751) );
  AOI22_X1 U22745 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19749), .B1(
        n19805), .B2(n19748), .ZN(n19750) );
  OAI211_X1 U22746 ( .C1(n19813), .C2(n19801), .A(n19751), .B(n19750), .ZN(
        P2_U3167) );
  NOR3_X1 U22747 ( .A1(n19752), .A2(n19804), .A3(n19959), .ZN(n19758) );
  INV_X1 U22748 ( .A(n19759), .ZN(n19753) );
  AOI21_X1 U22749 ( .B1(n19931), .B2(n19753), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19754) );
  NOR2_X1 U22750 ( .A1(n19758), .A2(n19754), .ZN(n19806) );
  AOI22_X1 U22751 ( .A1(n19806), .A2(n19226), .B1(n19804), .B2(n19755), .ZN(
        n19765) );
  NAND2_X1 U22752 ( .A1(n19757), .A2(n19756), .ZN(n19760) );
  AOI21_X1 U22753 ( .B1(n19760), .B2(n19759), .A(n19758), .ZN(n19762) );
  OAI211_X1 U22754 ( .C1(n19804), .C2(n19931), .A(n19762), .B(n19761), .ZN(
        n19809) );
  AOI22_X1 U22755 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19809), .B1(
        n19798), .B2(n19763), .ZN(n19764) );
  OAI211_X1 U22756 ( .C1(n19766), .C2(n19801), .A(n19765), .B(n19764), .ZN(
        P2_U3168) );
  AOI22_X1 U22757 ( .A1(n19806), .A2(n19234), .B1(n19804), .B2(n19767), .ZN(
        n19770) );
  AOI22_X1 U22758 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19809), .B1(
        n19808), .B2(n19768), .ZN(n19769) );
  OAI211_X1 U22759 ( .C1(n19771), .C2(n19812), .A(n19770), .B(n19769), .ZN(
        P2_U3169) );
  AOI22_X1 U22760 ( .A1(n19806), .A2(n19239), .B1(n19804), .B2(n19772), .ZN(
        n19775) );
  AOI22_X1 U22761 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19809), .B1(
        n19808), .B2(n19773), .ZN(n19774) );
  OAI211_X1 U22762 ( .C1(n19776), .C2(n19812), .A(n19775), .B(n19774), .ZN(
        P2_U3170) );
  AOI22_X1 U22763 ( .A1(n19806), .A2(n19778), .B1(n19804), .B2(n19777), .ZN(
        n19781) );
  AOI22_X1 U22764 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19809), .B1(
        n19798), .B2(n19779), .ZN(n19780) );
  OAI211_X1 U22765 ( .C1(n19782), .C2(n19801), .A(n19781), .B(n19780), .ZN(
        P2_U3171) );
  AOI22_X1 U22766 ( .A1(n19806), .A2(n19784), .B1(n19804), .B2(n19783), .ZN(
        n19787) );
  AOI22_X1 U22767 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19809), .B1(
        n19808), .B2(n19785), .ZN(n19786) );
  OAI211_X1 U22768 ( .C1(n19788), .C2(n19812), .A(n19787), .B(n19786), .ZN(
        P2_U3172) );
  AOI22_X1 U22769 ( .A1(n19806), .A2(n19790), .B1(n19804), .B2(n19789), .ZN(
        n19793) );
  AOI22_X1 U22770 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19809), .B1(
        n19808), .B2(n19791), .ZN(n19792) );
  OAI211_X1 U22771 ( .C1(n19794), .C2(n19812), .A(n19793), .B(n19792), .ZN(
        P2_U3173) );
  AOI22_X1 U22772 ( .A1(n19806), .A2(n19796), .B1(n19804), .B2(n19795), .ZN(
        n19800) );
  AOI22_X1 U22773 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19809), .B1(
        n19798), .B2(n19797), .ZN(n19799) );
  OAI211_X1 U22774 ( .C1(n19802), .C2(n19801), .A(n19800), .B(n19799), .ZN(
        P2_U3174) );
  AOI22_X1 U22775 ( .A1(n19806), .A2(n19805), .B1(n19804), .B2(n19803), .ZN(
        n19811) );
  AOI22_X1 U22776 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19809), .B1(
        n19808), .B2(n19807), .ZN(n19810) );
  OAI211_X1 U22777 ( .C1(n19813), .C2(n19812), .A(n19811), .B(n19810), .ZN(
        P2_U3175) );
  NOR2_X1 U22778 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n9877), .ZN(n19814) );
  OAI211_X1 U22779 ( .C1(n19815), .C2(n19814), .A(n19960), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19821) );
  NOR3_X1 U22780 ( .A1(n19960), .A2(n19816), .A3(n9877), .ZN(n19818) );
  OAI21_X1 U22781 ( .B1(n19819), .B2(n19818), .A(n19817), .ZN(n19820) );
  NAND3_X1 U22782 ( .A1(n19822), .A2(n19821), .A3(n19820), .ZN(P2_U3177) );
  AND2_X1 U22783 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n9635), .ZN(P2_U3179) );
  AND2_X1 U22784 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n9634), .ZN(P2_U3180) );
  AND2_X1 U22785 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n9635), .ZN(P2_U3181) );
  AND2_X1 U22786 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n9634), .ZN(P2_U3182) );
  AND2_X1 U22787 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n9635), .ZN(P2_U3183) );
  AND2_X1 U22788 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n9634), .ZN(P2_U3184) );
  AND2_X1 U22789 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n9635), .ZN(P2_U3185) );
  AND2_X1 U22790 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n9634), .ZN(P2_U3186) );
  AND2_X1 U22791 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n9634), .ZN(P2_U3187) );
  AND2_X1 U22792 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n9635), .ZN(P2_U3188) );
  AND2_X1 U22793 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n9634), .ZN(P2_U3189) );
  AND2_X1 U22794 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n9635), .ZN(P2_U3190) );
  AND2_X1 U22795 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n9634), .ZN(P2_U3191) );
  AND2_X1 U22796 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n9635), .ZN(P2_U3192) );
  AND2_X1 U22797 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n9634), .ZN(P2_U3193) );
  AND2_X1 U22798 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n9635), .ZN(P2_U3194) );
  AND2_X1 U22799 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n9634), .ZN(P2_U3195) );
  AND2_X1 U22800 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n9635), .ZN(P2_U3196) );
  AND2_X1 U22801 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n9635), .ZN(P2_U3197) );
  AND2_X1 U22802 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n9634), .ZN(P2_U3198) );
  AND2_X1 U22803 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n9635), .ZN(P2_U3199) );
  AND2_X1 U22804 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n9634), .ZN(P2_U3200) );
  AND2_X1 U22805 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n9634), .ZN(P2_U3201)
         );
  AND2_X1 U22806 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n9635), .ZN(P2_U3202)
         );
  AND2_X1 U22807 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n9634), .ZN(P2_U3203)
         );
  AND2_X1 U22808 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n9635), .ZN(P2_U3204)
         );
  AND2_X1 U22809 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n9634), .ZN(P2_U3205)
         );
  AND2_X1 U22810 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n9635), .ZN(P2_U3206)
         );
  AND2_X1 U22811 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n9634), .ZN(P2_U3207)
         );
  AND2_X1 U22812 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n9635), .ZN(P2_U3208)
         );
  NAND2_X1 U22813 ( .A1(n19960), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19836) );
  NAND3_X1 U22814 ( .A1(n19836), .A2(P2_STATE_REG_0__SCAN_IN), .A3(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19824) );
  OAI21_X1 U22815 ( .B1(n20957), .B2(n19828), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19838) );
  NAND2_X1 U22816 ( .A1(n19824), .A2(n19838), .ZN(n19825) );
  OAI221_X1 U22817 ( .B1(n19826), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .C1(
        n19826), .C2(n21032), .A(n19825), .ZN(P2_U3209) );
  NOR2_X1 U22818 ( .A1(HOLD), .A2(n19827), .ZN(n19837) );
  OAI211_X1 U22819 ( .C1(n19837), .C2(n19839), .A(
        P2_REQUESTPENDING_REG_SCAN_IN), .B(n19828), .ZN(n19829) );
  AND3_X1 U22820 ( .A1(n19830), .A2(n19836), .A3(n19829), .ZN(n19831) );
  OAI21_X1 U22821 ( .B1(n21032), .B2(n19832), .A(n19831), .ZN(P2_U3210) );
  OAI22_X1 U22822 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19833), .B1(NA), 
        .B2(n19836), .ZN(n19834) );
  OAI211_X1 U22823 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19834), .ZN(n19835) );
  OAI221_X1 U22824 ( .B1(n19838), .B2(n19837), .C1(n19838), .C2(n19836), .A(
        n19835), .ZN(P2_U3211) );
  OAI222_X1 U22825 ( .A1(n19886), .A2(n19841), .B1(n19840), .B2(n19974), .C1(
        n10595), .C2(n19884), .ZN(P2_U3212) );
  OAI222_X1 U22826 ( .A1(n19886), .A2(n12705), .B1(n19842), .B2(n19974), .C1(
        n19841), .C2(n19884), .ZN(P2_U3213) );
  OAI222_X1 U22827 ( .A1(n19886), .A2(n12677), .B1(n19843), .B2(n19974), .C1(
        n12705), .C2(n19884), .ZN(P2_U3214) );
  OAI222_X1 U22828 ( .A1(n19886), .A2(n12673), .B1(n19844), .B2(n19974), .C1(
        n12677), .C2(n19884), .ZN(P2_U3215) );
  OAI222_X1 U22829 ( .A1(n19886), .A2(n19846), .B1(n19845), .B2(n19974), .C1(
        n12673), .C2(n19884), .ZN(P2_U3216) );
  OAI222_X1 U22830 ( .A1(n19886), .A2(n19848), .B1(n19847), .B2(n19974), .C1(
        n19846), .C2(n19884), .ZN(P2_U3217) );
  INV_X1 U22831 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19850) );
  OAI222_X1 U22832 ( .A1(n19886), .A2(n19850), .B1(n19849), .B2(n19974), .C1(
        n19848), .C2(n19884), .ZN(P2_U3218) );
  OAI222_X1 U22833 ( .A1(n19886), .A2(n12744), .B1(n19851), .B2(n19974), .C1(
        n19850), .C2(n19884), .ZN(P2_U3219) );
  OAI222_X1 U22834 ( .A1(n19886), .A2(n12747), .B1(n19852), .B2(n19974), .C1(
        n12744), .C2(n19884), .ZN(P2_U3220) );
  INV_X1 U22835 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19854) );
  OAI222_X1 U22836 ( .A1(n19886), .A2(n19854), .B1(n19853), .B2(n19974), .C1(
        n12747), .C2(n19884), .ZN(P2_U3221) );
  OAI222_X1 U22837 ( .A1(n19886), .A2(n19856), .B1(n19855), .B2(n19974), .C1(
        n19854), .C2(n19884), .ZN(P2_U3222) );
  OAI222_X1 U22838 ( .A1(n19886), .A2(n12807), .B1(n19857), .B2(n19974), .C1(
        n19856), .C2(n19884), .ZN(P2_U3223) );
  OAI222_X1 U22839 ( .A1(n19886), .A2(n12810), .B1(n19858), .B2(n19974), .C1(
        n12807), .C2(n19884), .ZN(P2_U3224) );
  OAI222_X1 U22840 ( .A1(n19886), .A2(n12839), .B1(n19859), .B2(n19974), .C1(
        n12810), .C2(n19884), .ZN(P2_U3225) );
  OAI222_X1 U22841 ( .A1(n19886), .A2(n12843), .B1(n19860), .B2(n19974), .C1(
        n12839), .C2(n19884), .ZN(P2_U3226) );
  OAI222_X1 U22842 ( .A1(n19886), .A2(n19862), .B1(n19861), .B2(n19974), .C1(
        n12843), .C2(n19884), .ZN(P2_U3227) );
  OAI222_X1 U22843 ( .A1(n19886), .A2(n14914), .B1(n19863), .B2(n19974), .C1(
        n19862), .C2(n19884), .ZN(P2_U3228) );
  OAI222_X1 U22844 ( .A1(n19886), .A2(n19865), .B1(n19864), .B2(n19974), .C1(
        n14914), .C2(n19884), .ZN(P2_U3229) );
  OAI222_X1 U22845 ( .A1(n19886), .A2(n19867), .B1(n19866), .B2(n19974), .C1(
        n19865), .C2(n19884), .ZN(P2_U3230) );
  OAI222_X1 U22846 ( .A1(n19886), .A2(n19869), .B1(n19868), .B2(n19974), .C1(
        n19867), .C2(n19884), .ZN(P2_U3231) );
  OAI222_X1 U22847 ( .A1(n19886), .A2(n12856), .B1(n19870), .B2(n19974), .C1(
        n19869), .C2(n19884), .ZN(P2_U3232) );
  OAI222_X1 U22848 ( .A1(n19886), .A2(n19872), .B1(n19871), .B2(n19974), .C1(
        n12856), .C2(n19884), .ZN(P2_U3233) );
  OAI222_X1 U22849 ( .A1(n19886), .A2(n19874), .B1(n19873), .B2(n19974), .C1(
        n19872), .C2(n19884), .ZN(P2_U3234) );
  OAI222_X1 U22850 ( .A1(n19886), .A2(n19876), .B1(n19875), .B2(n19974), .C1(
        n19874), .C2(n19884), .ZN(P2_U3235) );
  OAI222_X1 U22851 ( .A1(n19886), .A2(n16073), .B1(n19877), .B2(n19974), .C1(
        n19876), .C2(n19884), .ZN(P2_U3236) );
  OAI222_X1 U22852 ( .A1(n19886), .A2(n19880), .B1(n19878), .B2(n19974), .C1(
        n16073), .C2(n19884), .ZN(P2_U3237) );
  OAI222_X1 U22853 ( .A1(n19884), .A2(n19880), .B1(n19879), .B2(n19974), .C1(
        n12870), .C2(n19886), .ZN(P2_U3238) );
  OAI222_X1 U22854 ( .A1(n19886), .A2(n19882), .B1(n19881), .B2(n19974), .C1(
        n12870), .C2(n19884), .ZN(P2_U3239) );
  OAI222_X1 U22855 ( .A1(n19886), .A2(n12876), .B1(n19883), .B2(n19974), .C1(
        n19882), .C2(n19884), .ZN(P2_U3240) );
  INV_X1 U22856 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19885) );
  OAI222_X1 U22857 ( .A1(n19886), .A2(n14833), .B1(n19885), .B2(n19974), .C1(
        n12876), .C2(n19884), .ZN(P2_U3241) );
  INV_X1 U22858 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19887) );
  AOI22_X1 U22859 ( .A1(n19974), .A2(n19888), .B1(n19887), .B2(n19971), .ZN(
        P2_U3585) );
  MUX2_X1 U22860 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n19974), .Z(P2_U3586) );
  INV_X1 U22861 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n19889) );
  AOI22_X1 U22862 ( .A1(n19974), .A2(n19890), .B1(n19889), .B2(n19971), .ZN(
        P2_U3587) );
  INV_X1 U22863 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19891) );
  AOI22_X1 U22864 ( .A1(n19974), .A2(n19892), .B1(n19891), .B2(n19971), .ZN(
        P2_U3588) );
  AOI21_X1 U22865 ( .B1(n9635), .B2(n19894), .A(n19893), .ZN(P2_U3591) );
  OAI21_X1 U22866 ( .B1(n19897), .B2(n19896), .A(n19895), .ZN(P2_U3592) );
  INV_X1 U22867 ( .A(n19898), .ZN(n19910) );
  AND2_X1 U22868 ( .A1(n19902), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19925) );
  NAND2_X1 U22869 ( .A1(n19899), .A2(n19925), .ZN(n19916) );
  OR2_X1 U22870 ( .A1(n19901), .A2(n19900), .ZN(n19924) );
  AOI21_X1 U22871 ( .B1(n19903), .B2(n19902), .A(n19924), .ZN(n19914) );
  AOI21_X1 U22872 ( .B1(n19916), .B2(n19914), .A(n19904), .ZN(n19909) );
  NOR3_X1 U22873 ( .A1(n19907), .A2(n19906), .A3(n19905), .ZN(n19908) );
  AOI211_X1 U22874 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19910), .A(n19909), 
        .B(n19908), .ZN(n19911) );
  AOI22_X1 U22875 ( .A1(n19940), .A2(n19912), .B1(n19911), .B2(n19937), .ZN(
        P2_U3602) );
  INV_X1 U22876 ( .A(n19913), .ZN(n19920) );
  INV_X1 U22877 ( .A(n19914), .ZN(n19919) );
  NOR2_X1 U22878 ( .A1(n19915), .A2(n19931), .ZN(n19918) );
  INV_X1 U22879 ( .A(n19916), .ZN(n19917) );
  AOI211_X1 U22880 ( .C1(n19920), .C2(n19919), .A(n19918), .B(n19917), .ZN(
        n19921) );
  AOI22_X1 U22881 ( .A1(n19940), .A2(n19922), .B1(n19921), .B2(n19937), .ZN(
        P2_U3603) );
  MUX2_X1 U22882 ( .A(n19925), .B(n19924), .S(n19923), .Z(n19926) );
  AOI21_X1 U22883 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19927), .A(n19926), 
        .ZN(n19928) );
  AOI22_X1 U22884 ( .A1(n19940), .A2(n19929), .B1(n19928), .B2(n19937), .ZN(
        P2_U3604) );
  INV_X1 U22885 ( .A(n19930), .ZN(n19932) );
  OAI22_X1 U22886 ( .A1(n19933), .A2(n19932), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19931), .ZN(n19934) );
  AOI21_X1 U22887 ( .B1(n19936), .B2(n19935), .A(n19934), .ZN(n19938) );
  AOI22_X1 U22888 ( .A1(n19940), .A2(n19939), .B1(n19938), .B2(n19937), .ZN(
        P2_U3605) );
  INV_X1 U22889 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19941) );
  AOI22_X1 U22890 ( .A1(n19974), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19941), 
        .B2(n19971), .ZN(P2_U3608) );
  INV_X1 U22891 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n19954) );
  INV_X1 U22892 ( .A(n19942), .ZN(n19953) );
  INV_X1 U22893 ( .A(n19943), .ZN(n19947) );
  INV_X1 U22894 ( .A(n19944), .ZN(n19945) );
  OAI22_X1 U22895 ( .A1(n19948), .A2(n19947), .B1(n19946), .B2(n19945), .ZN(
        n19949) );
  INV_X1 U22896 ( .A(n19949), .ZN(n19952) );
  NOR2_X1 U22897 ( .A1(n19953), .A2(n19950), .ZN(n19951) );
  AOI22_X1 U22898 ( .A1(n19954), .A2(n19953), .B1(n19952), .B2(n19951), .ZN(
        P2_U3609) );
  OAI21_X1 U22899 ( .B1(n19956), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19955), 
        .ZN(n19957) );
  NAND3_X1 U22900 ( .A1(n19958), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n19957), 
        .ZN(n19963) );
  OAI22_X1 U22901 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19961), .B1(n19960), 
        .B2(n19959), .ZN(n19962) );
  NAND2_X1 U22902 ( .A1(n19963), .A2(n19962), .ZN(n19970) );
  AOI21_X1 U22903 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19964), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19966) );
  AOI211_X1 U22904 ( .C1(n19968), .C2(n19967), .A(n19966), .B(n19965), .ZN(
        n19969) );
  MUX2_X1 U22905 ( .A(n19970), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n19969), 
        .Z(P2_U3610) );
  INV_X1 U22906 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n19972) );
  AOI22_X1 U22907 ( .A1(n19974), .A2(n19973), .B1(n19972), .B2(n19971), .ZN(
        P2_U3611) );
  AOI21_X1 U22908 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n11603), .A(n12453), 
        .ZN(n19981) );
  INV_X1 U22909 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20982) );
  NOR2_X1 U22910 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20778), .ZN(n20840) );
  INV_X1 U22911 ( .A(n20883), .ZN(n20885) );
  AOI21_X1 U22912 ( .B1(n19981), .B2(n20982), .A(n20885), .ZN(P1_U2802) );
  INV_X1 U22913 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n20984) );
  AOI21_X1 U22914 ( .B1(n19976), .B2(n19975), .A(n20984), .ZN(n19977) );
  AOI21_X1 U22915 ( .B1(n11773), .B2(n19978), .A(n19977), .ZN(n19979) );
  INV_X1 U22916 ( .A(n19979), .ZN(P1_U2803) );
  INV_X1 U22917 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n20991) );
  NOR2_X1 U22918 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19982) );
  NOR2_X1 U22919 ( .A1(n20885), .A2(n19982), .ZN(n19980) );
  AOI22_X1 U22920 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(n20885), .B1(n20991), 
        .B2(n19980), .ZN(P1_U2804) );
  NOR2_X1 U22921 ( .A1(n20885), .A2(n19981), .ZN(n20854) );
  OAI21_X1 U22922 ( .B1(BS16), .B2(n19982), .A(n20854), .ZN(n20852) );
  OAI21_X1 U22923 ( .B1(n20854), .B2(n20874), .A(n20852), .ZN(P1_U2805) );
  OAI21_X1 U22924 ( .B1(n19984), .B2(n19983), .A(n20172), .ZN(P1_U2806) );
  NOR4_X1 U22925 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19988) );
  NOR4_X1 U22926 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19987) );
  NOR4_X1 U22927 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19986) );
  NOR4_X1 U22928 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19985) );
  NAND4_X1 U22929 ( .A1(n19988), .A2(n19987), .A3(n19986), .A4(n19985), .ZN(
        n19994) );
  NOR4_X1 U22930 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19992) );
  AOI211_X1 U22931 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19991) );
  NOR4_X1 U22932 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19990) );
  NOR4_X1 U22933 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19989) );
  NAND4_X1 U22934 ( .A1(n19992), .A2(n19991), .A3(n19990), .A4(n19989), .ZN(
        n19993) );
  NOR2_X1 U22935 ( .A1(n19994), .A2(n19993), .ZN(n20867) );
  INV_X1 U22936 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20847) );
  NOR3_X1 U22937 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19996) );
  OAI21_X1 U22938 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19996), .A(n20867), .ZN(
        n19995) );
  OAI21_X1 U22939 ( .B1(n20867), .B2(n20847), .A(n19995), .ZN(P1_U2807) );
  INV_X1 U22940 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20853) );
  AOI21_X1 U22941 ( .B1(n13342), .B2(n20853), .A(n19996), .ZN(n19997) );
  INV_X1 U22942 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20844) );
  INV_X1 U22943 ( .A(n20867), .ZN(n20863) );
  AOI22_X1 U22944 ( .A1(n20867), .A2(n19997), .B1(n20844), .B2(n20863), .ZN(
        P1_U2808) );
  NAND2_X1 U22945 ( .A1(n20021), .A2(n19998), .ZN(n20020) );
  INV_X1 U22946 ( .A(n19999), .ZN(n20062) );
  NOR2_X1 U22947 ( .A1(n20000), .A2(n11886), .ZN(n20001) );
  AOI211_X1 U22948 ( .C1(n20002), .C2(n20027), .A(n20040), .B(n20001), .ZN(
        n20005) );
  INV_X1 U22949 ( .A(n20003), .ZN(n20061) );
  NAND2_X1 U22950 ( .A1(n20047), .A2(n20061), .ZN(n20004) );
  OAI211_X1 U22951 ( .C1(n20064), .C2(n20054), .A(n20005), .B(n20004), .ZN(
        n20006) );
  AOI21_X1 U22952 ( .B1(n20062), .B2(n20041), .A(n20006), .ZN(n20007) );
  OAI221_X1 U22953 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n20008), .C1(n20804), 
        .C2(n20020), .A(n20007), .ZN(P1_U2831) );
  OAI22_X1 U22954 ( .A1(n20054), .A2(n20010), .B1(n20009), .B2(n20053), .ZN(
        n20011) );
  INV_X1 U22955 ( .A(n20011), .ZN(n20012) );
  OAI21_X1 U22956 ( .B1(n20014), .B2(n20013), .A(n20012), .ZN(n20015) );
  AOI211_X1 U22957 ( .C1(n20048), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n20040), .B(n20015), .ZN(n20019) );
  AOI22_X1 U22958 ( .A1(n20017), .A2(n20041), .B1(n20016), .B2(n20802), .ZN(
        n20018) );
  OAI211_X1 U22959 ( .C1(n20802), .C2(n20020), .A(n20019), .B(n20018), .ZN(
        P1_U2832) );
  OAI21_X1 U22960 ( .B1(n20023), .B2(n20022), .A(n20021), .ZN(n20045) );
  NOR3_X1 U22961 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20051), .A3(n20023), .ZN(
        n20024) );
  AOI211_X1 U22962 ( .C1(n20047), .C2(n20065), .A(n20040), .B(n20024), .ZN(
        n20029) );
  INV_X1 U22963 ( .A(n20025), .ZN(n20026) );
  AOI22_X1 U22964 ( .A1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n20048), .B1(
        n20027), .B2(n20026), .ZN(n20028) );
  OAI211_X1 U22965 ( .C1(n20068), .C2(n20054), .A(n20029), .B(n20028), .ZN(
        n20030) );
  AOI21_X1 U22966 ( .B1(n20041), .B2(n20066), .A(n20030), .ZN(n20031) );
  OAI21_X1 U22967 ( .B1(n20045), .B2(n20800), .A(n20031), .ZN(P1_U2833) );
  INV_X1 U22968 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20798) );
  OAI22_X1 U22969 ( .A1(n20054), .A2(n20033), .B1(n20032), .B2(n20053), .ZN(
        n20034) );
  INV_X1 U22970 ( .A(n20034), .ZN(n20044) );
  AOI22_X1 U22971 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n20048), .B1(
        n20047), .B2(n20035), .ZN(n20038) );
  INV_X1 U22972 ( .A(n20051), .ZN(n20036) );
  NAND3_X1 U22973 ( .A1(n20036), .A2(n20798), .A3(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20037) );
  NAND2_X1 U22974 ( .A1(n20038), .A2(n20037), .ZN(n20039) );
  AOI211_X1 U22975 ( .C1(n20042), .C2(n20041), .A(n20040), .B(n20039), .ZN(
        n20043) );
  OAI211_X1 U22976 ( .C1(n20045), .C2(n20798), .A(n20044), .B(n20043), .ZN(
        P1_U2834) );
  INV_X1 U22977 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20796) );
  NAND2_X1 U22978 ( .A1(n20072), .A2(n20046), .ZN(n20058) );
  AOI22_X1 U22979 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20048), .B1(
        n20047), .B2(n20069), .ZN(n20050) );
  OAI211_X1 U22980 ( .C1(P1_REIP_REG_5__SCAN_IN), .C2(n20051), .A(n20050), .B(
        n20049), .ZN(n20056) );
  INV_X1 U22981 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20074) );
  OAI22_X1 U22982 ( .A1(n20054), .A2(n20074), .B1(n20053), .B2(n20052), .ZN(
        n20055) );
  NOR2_X1 U22983 ( .A1(n20056), .A2(n20055), .ZN(n20057) );
  AND2_X1 U22984 ( .A1(n20058), .A2(n20057), .ZN(n20059) );
  OAI21_X1 U22985 ( .B1(n20796), .B2(n20060), .A(n20059), .ZN(P1_U2835) );
  AOI22_X1 U22986 ( .A1(n20062), .A2(n20071), .B1(n20070), .B2(n20061), .ZN(
        n20063) );
  OAI21_X1 U22987 ( .B1(n20075), .B2(n20064), .A(n20063), .ZN(P1_U2863) );
  AOI22_X1 U22988 ( .A1(n20066), .A2(n20071), .B1(n20070), .B2(n20065), .ZN(
        n20067) );
  OAI21_X1 U22989 ( .B1(n20075), .B2(n20068), .A(n20067), .ZN(P1_U2865) );
  AOI22_X1 U22990 ( .A1(n20072), .A2(n20071), .B1(n20070), .B2(n20069), .ZN(
        n20073) );
  OAI21_X1 U22991 ( .B1(n20075), .B2(n20074), .A(n20073), .ZN(P1_U2867) );
  AOI22_X1 U22992 ( .A1(n20872), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20101), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20077) );
  OAI21_X1 U22993 ( .B1(n20078), .B2(n20104), .A(n20077), .ZN(P1_U2921) );
  AOI22_X1 U22994 ( .A1(n20872), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20101), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20079) );
  OAI21_X1 U22995 ( .B1(n14552), .B2(n20104), .A(n20079), .ZN(P1_U2922) );
  AOI22_X1 U22996 ( .A1(n20872), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20101), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20080) );
  OAI21_X1 U22997 ( .B1(n14556), .B2(n20104), .A(n20080), .ZN(P1_U2923) );
  AOI22_X1 U22998 ( .A1(n20872), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20101), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20081) );
  OAI21_X1 U22999 ( .B1(n20082), .B2(n20104), .A(n20081), .ZN(P1_U2924) );
  AOI22_X1 U23000 ( .A1(n20872), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20101), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20083) );
  OAI21_X1 U23001 ( .B1(n14563), .B2(n20104), .A(n20083), .ZN(P1_U2925) );
  AOI22_X1 U23002 ( .A1(n20872), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20101), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20084) );
  OAI21_X1 U23003 ( .B1(n14224), .B2(n20104), .A(n20084), .ZN(P1_U2926) );
  AOI22_X1 U23004 ( .A1(n20872), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20101), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20085) );
  OAI21_X1 U23005 ( .B1(n20086), .B2(n20104), .A(n20085), .ZN(P1_U2927) );
  AOI22_X1 U23006 ( .A1(n20872), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20101), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20087) );
  OAI21_X1 U23007 ( .B1(n20088), .B2(n20104), .A(n20087), .ZN(P1_U2928) );
  AOI22_X1 U23008 ( .A1(n20102), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20101), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20089) );
  OAI21_X1 U23009 ( .B1(n11779), .B2(n20104), .A(n20089), .ZN(P1_U2929) );
  AOI22_X1 U23010 ( .A1(n20102), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20101), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20090) );
  OAI21_X1 U23011 ( .B1(n11784), .B2(n20104), .A(n20090), .ZN(P1_U2930) );
  AOI22_X1 U23012 ( .A1(n20102), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20101), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20091) );
  OAI21_X1 U23013 ( .B1(n20092), .B2(n20104), .A(n20091), .ZN(P1_U2931) );
  AOI22_X1 U23014 ( .A1(n20102), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20101), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20093) );
  OAI21_X1 U23015 ( .B1(n20094), .B2(n20104), .A(n20093), .ZN(P1_U2932) );
  AOI22_X1 U23016 ( .A1(n20102), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20101), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20095) );
  OAI21_X1 U23017 ( .B1(n20096), .B2(n20104), .A(n20095), .ZN(P1_U2933) );
  AOI22_X1 U23018 ( .A1(n20102), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20101), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20097) );
  OAI21_X1 U23019 ( .B1(n20098), .B2(n20104), .A(n20097), .ZN(P1_U2934) );
  AOI22_X1 U23020 ( .A1(n20102), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20101), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20099) );
  OAI21_X1 U23021 ( .B1(n20100), .B2(n20104), .A(n20099), .ZN(P1_U2935) );
  AOI22_X1 U23022 ( .A1(n20102), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20101), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20103) );
  OAI21_X1 U23023 ( .B1(n20105), .B2(n20104), .A(n20103), .ZN(P1_U2936) );
  AOI22_X1 U23024 ( .A1(n20131), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20147), .ZN(n20106) );
  OAI21_X1 U23025 ( .B1(n20214), .B2(n20150), .A(n20106), .ZN(P1_U2937) );
  AOI22_X1 U23026 ( .A1(n20131), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20147), .ZN(n20107) );
  OAI21_X1 U23027 ( .B1(n20118), .B2(n20150), .A(n20107), .ZN(P1_U2938) );
  AOI22_X1 U23028 ( .A1(n20131), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20147), .ZN(n20108) );
  OAI21_X1 U23029 ( .B1(n20120), .B2(n20150), .A(n20108), .ZN(P1_U2939) );
  AOI22_X1 U23030 ( .A1(n20131), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20147), .ZN(n20109) );
  OAI21_X1 U23031 ( .B1(n20228), .B2(n20150), .A(n20109), .ZN(P1_U2940) );
  AOI22_X1 U23032 ( .A1(n20131), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20147), .ZN(n20110) );
  OAI21_X1 U23033 ( .B1(n20123), .B2(n20150), .A(n20110), .ZN(P1_U2941) );
  AOI22_X1 U23034 ( .A1(n20131), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20147), .ZN(n20111) );
  OAI21_X1 U23035 ( .B1(n20125), .B2(n20150), .A(n20111), .ZN(P1_U2942) );
  AOI22_X1 U23036 ( .A1(n20131), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20147), .ZN(n20112) );
  OAI21_X1 U23037 ( .B1(n20246), .B2(n20150), .A(n20112), .ZN(P1_U2943) );
  AOI22_X1 U23038 ( .A1(n20131), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20147), .ZN(n20113) );
  OAI21_X1 U23039 ( .B1(n20128), .B2(n20150), .A(n20113), .ZN(P1_U2944) );
  AOI22_X1 U23040 ( .A1(n20131), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20147), .ZN(n20114) );
  OAI21_X1 U23041 ( .B1(n20130), .B2(n20150), .A(n20114), .ZN(P1_U2945) );
  AOI22_X1 U23042 ( .A1(n20131), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20147), .ZN(n20115) );
  OAI21_X1 U23043 ( .B1(n20139), .B2(n20150), .A(n20115), .ZN(P1_U2949) );
  AOI22_X1 U23044 ( .A1(n20131), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20147), .ZN(n20116) );
  OAI21_X1 U23045 ( .B1(n20214), .B2(n20150), .A(n20116), .ZN(P1_U2952) );
  AOI22_X1 U23046 ( .A1(n20131), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20147), .ZN(n20117) );
  OAI21_X1 U23047 ( .B1(n20118), .B2(n20150), .A(n20117), .ZN(P1_U2953) );
  AOI22_X1 U23048 ( .A1(n9678), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20147), .ZN(n20119) );
  OAI21_X1 U23049 ( .B1(n20120), .B2(n20150), .A(n20119), .ZN(P1_U2954) );
  AOI22_X1 U23050 ( .A1(n9678), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20147), .ZN(n20121) );
  OAI21_X1 U23051 ( .B1(n20228), .B2(n20150), .A(n20121), .ZN(P1_U2955) );
  AOI22_X1 U23052 ( .A1(n9678), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20147), .ZN(n20122) );
  OAI21_X1 U23053 ( .B1(n20123), .B2(n20150), .A(n20122), .ZN(P1_U2956) );
  AOI22_X1 U23054 ( .A1(n20131), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20147), .ZN(n20124) );
  OAI21_X1 U23055 ( .B1(n20125), .B2(n20150), .A(n20124), .ZN(P1_U2957) );
  AOI22_X1 U23056 ( .A1(n9678), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20147), .ZN(n20126) );
  OAI21_X1 U23057 ( .B1(n20246), .B2(n20150), .A(n20126), .ZN(P1_U2958) );
  AOI22_X1 U23058 ( .A1(n9678), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20147), .ZN(n20127) );
  OAI21_X1 U23059 ( .B1(n20128), .B2(n20150), .A(n20127), .ZN(P1_U2959) );
  AOI22_X1 U23060 ( .A1(n9678), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20147), .ZN(n20129) );
  OAI21_X1 U23061 ( .B1(n20130), .B2(n20150), .A(n20129), .ZN(P1_U2960) );
  AOI22_X1 U23062 ( .A1(n20131), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20147), .ZN(n20134) );
  NAND2_X1 U23063 ( .A1(n20144), .A2(n20132), .ZN(n20133) );
  NAND2_X1 U23064 ( .A1(n20134), .A2(n20133), .ZN(P1_U2962) );
  AOI22_X1 U23065 ( .A1(n9678), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20147), .ZN(n20137) );
  NAND2_X1 U23066 ( .A1(n20144), .A2(n20135), .ZN(n20136) );
  NAND2_X1 U23067 ( .A1(n20137), .A2(n20136), .ZN(P1_U2963) );
  AOI22_X1 U23068 ( .A1(n9678), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20147), .ZN(n20138) );
  OAI21_X1 U23069 ( .B1(n20139), .B2(n20150), .A(n20138), .ZN(P1_U2964) );
  AOI22_X1 U23070 ( .A1(n9678), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20147), .ZN(n20142) );
  NAND2_X1 U23071 ( .A1(n20144), .A2(n20140), .ZN(n20141) );
  NAND2_X1 U23072 ( .A1(n20142), .A2(n20141), .ZN(P1_U2965) );
  AOI22_X1 U23073 ( .A1(n9678), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20147), .ZN(n20146) );
  NAND2_X1 U23074 ( .A1(n20144), .A2(n20143), .ZN(n20145) );
  NAND2_X1 U23075 ( .A1(n20146), .A2(n20145), .ZN(P1_U2966) );
  AOI22_X1 U23076 ( .A1(n9678), .A2(P1_EAX_REG_15__SCAN_IN), .B1(
        P1_LWORD_REG_15__SCAN_IN), .B2(n20147), .ZN(n20149) );
  OAI21_X1 U23077 ( .B1(n20151), .B2(n20150), .A(n20149), .ZN(P1_U2967) );
  AOI22_X1 U23078 ( .A1(n20152), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20190), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20159) );
  INV_X1 U23079 ( .A(n20153), .ZN(n20157) );
  AOI22_X1 U23080 ( .A1(n20157), .A2(n20156), .B1(n20155), .B2(n20154), .ZN(
        n20158) );
  OAI211_X1 U23081 ( .C1(n20161), .C2(n20160), .A(n20159), .B(n20158), .ZN(
        P1_U2995) );
  OAI21_X1 U23082 ( .B1(n20163), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n20162), .ZN(n20207) );
  NAND2_X1 U23083 ( .A1(n20165), .A2(n20164), .ZN(n20166) );
  AOI22_X1 U23084 ( .A1(n20168), .A2(n20167), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20166), .ZN(n20171) );
  INV_X1 U23085 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n20169) );
  OR2_X1 U23086 ( .A1(n20170), .A2(n20169), .ZN(n20197) );
  OAI211_X1 U23087 ( .C1(n20172), .C2(n20207), .A(n20171), .B(n20197), .ZN(
        P1_U2999) );
  AOI21_X1 U23088 ( .B1(n20203), .B2(n20174), .A(n20173), .ZN(n20178) );
  AOI22_X1 U23089 ( .A1(n20176), .A2(n20179), .B1(n20175), .B2(n20188), .ZN(
        n20177) );
  OAI211_X1 U23090 ( .C1(n20180), .C2(n20179), .A(n20178), .B(n20177), .ZN(
        P1_U3028) );
  NAND2_X1 U23091 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20182) );
  OAI21_X1 U23092 ( .B1(n20182), .B2(n20191), .A(n20181), .ZN(n20184) );
  AOI22_X1 U23093 ( .A1(n20185), .A2(n20184), .B1(n20203), .B2(n20183), .ZN(
        n20196) );
  INV_X1 U23094 ( .A(n20186), .ZN(n20189) );
  AOI22_X1 U23095 ( .A1(n20189), .A2(n20188), .B1(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20187), .ZN(n20195) );
  NAND2_X1 U23096 ( .A1(n20190), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n20194) );
  NAND3_X1 U23097 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20192), .A3(
        n20191), .ZN(n20193) );
  NAND4_X1 U23098 ( .A1(n20196), .A2(n20195), .A3(n20194), .A4(n20193), .ZN(
        P1_U3029) );
  INV_X1 U23099 ( .A(n20197), .ZN(n20202) );
  AOI21_X1 U23100 ( .B1(n20200), .B2(n20199), .A(n20198), .ZN(n20201) );
  AOI211_X1 U23101 ( .C1(n20204), .C2(n20203), .A(n20202), .B(n20201), .ZN(
        n20206) );
  OAI211_X1 U23102 ( .C1(n20208), .C2(n20207), .A(n20206), .B(n20205), .ZN(
        P1_U3031) );
  NOR2_X1 U23103 ( .A1(n20210), .A2(n20209), .ZN(P1_U3032) );
  INV_X1 U23104 ( .A(DATAI_24_), .ZN(n20933) );
  INV_X1 U23105 ( .A(n20722), .ZN(n20645) );
  NOR2_X2 U23106 ( .A1(n20235), .A2(n20212), .ZN(n20713) );
  INV_X1 U23107 ( .A(n20713), .ZN(n20583) );
  OAI22_X1 U23108 ( .A1(n20773), .A2(n20645), .B1(n20583), .B2(n20244), .ZN(
        n20213) );
  INV_X1 U23109 ( .A(n20213), .ZN(n20217) );
  INV_X1 U23110 ( .A(DATAI_16_), .ZN(n21026) );
  OAI22_X1 U23111 ( .A1(n20215), .A2(n20248), .B1(n21026), .B2(n20247), .ZN(
        n20642) );
  AOI22_X1 U23112 ( .A1(n20712), .A2(n20250), .B1(n20279), .B2(n20642), .ZN(
        n20216) );
  OAI211_X1 U23113 ( .C1(n20254), .C2(n20218), .A(n20217), .B(n20216), .ZN(
        P1_U3033) );
  INV_X1 U23114 ( .A(DATAI_25_), .ZN(n21033) );
  INV_X1 U23115 ( .A(n20728), .ZN(n20649) );
  NOR2_X2 U23116 ( .A1(n20235), .A2(n20220), .ZN(n20727) );
  INV_X1 U23117 ( .A(n20727), .ZN(n20595) );
  OAI22_X1 U23118 ( .A1(n20773), .A2(n20649), .B1(n20595), .B2(n20244), .ZN(
        n20221) );
  INV_X1 U23119 ( .A(n20221), .ZN(n20225) );
  NAND2_X1 U23120 ( .A1(n20261), .A2(n20222), .ZN(n20599) );
  INV_X1 U23121 ( .A(n20599), .ZN(n20726) );
  INV_X1 U23122 ( .A(DATAI_17_), .ZN(n20990) );
  OAI22_X1 U23123 ( .A1(n20990), .A2(n20247), .B1(n20223), .B2(n20248), .ZN(
        n20646) );
  AOI22_X1 U23124 ( .A1(n20726), .A2(n20250), .B1(n20279), .B2(n20646), .ZN(
        n20224) );
  OAI211_X1 U23125 ( .C1(n20254), .C2(n11673), .A(n20225), .B(n20224), .ZN(
        P1_U3034) );
  INV_X1 U23126 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n20232) );
  INV_X1 U23127 ( .A(DATAI_27_), .ZN(n20922) );
  INV_X1 U23128 ( .A(n20235), .ZN(n20243) );
  NAND2_X1 U23129 ( .A1(n20243), .A2(n20227), .ZN(n20605) );
  AOI22_X1 U23130 ( .A1(n20759), .A2(n20688), .B1(n20236), .B2(n20739), .ZN(
        n20231) );
  INV_X1 U23131 ( .A(DATAI_19_), .ZN(n20988) );
  OAI22_X1 U23132 ( .A1(n20229), .A2(n20248), .B1(n20988), .B2(n20247), .ZN(
        n20740) );
  AOI22_X1 U23133 ( .A1(n20738), .A2(n20250), .B1(n20279), .B2(n20740), .ZN(
        n20230) );
  OAI211_X1 U23134 ( .C1(n20254), .C2(n20232), .A(n20231), .B(n20230), .ZN(
        P1_U3036) );
  INV_X1 U23135 ( .A(DATAI_29_), .ZN(n20233) );
  NOR2_X2 U23136 ( .A1(n20235), .A2(n11606), .ZN(n20751) );
  AOI22_X1 U23137 ( .A1(n20759), .A2(n20694), .B1(n20236), .B2(n20751), .ZN(
        n20241) );
  NAND2_X1 U23138 ( .A1(n20261), .A2(n20237), .ZN(n20619) );
  INV_X1 U23139 ( .A(n20619), .ZN(n20750) );
  INV_X1 U23140 ( .A(DATAI_21_), .ZN(n20239) );
  AOI22_X1 U23141 ( .A1(n20750), .A2(n20250), .B1(n20279), .B2(n20752), .ZN(
        n20240) );
  OAI211_X1 U23142 ( .C1(n20254), .C2(n20242), .A(n20241), .B(n20240), .ZN(
        P1_U3038) );
  INV_X1 U23143 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20253) );
  INV_X1 U23144 ( .A(DATAI_30_), .ZN(n21027) );
  INV_X1 U23145 ( .A(n20698), .ZN(n20763) );
  OAI22_X1 U23146 ( .A1(n20773), .A2(n20763), .B1(n20244), .B2(n20620), .ZN(
        n20245) );
  INV_X1 U23147 ( .A(n20245), .ZN(n20252) );
  INV_X1 U23148 ( .A(DATAI_22_), .ZN(n20952) );
  OAI22_X1 U23149 ( .A1(n20249), .A2(n20248), .B1(n20952), .B2(n20247), .ZN(
        n20758) );
  AOI22_X1 U23150 ( .A1(n20756), .A2(n20250), .B1(n20279), .B2(n20758), .ZN(
        n20251) );
  OAI211_X1 U23151 ( .C1(n20254), .C2(n20253), .A(n20252), .B(n20251), .ZN(
        P1_U3039) );
  INV_X1 U23152 ( .A(n20642), .ZN(n20725) );
  INV_X1 U23153 ( .A(n20641), .ZN(n20255) );
  NOR2_X1 U23154 ( .A1(n20634), .A2(n20259), .ZN(n20278) );
  INV_X1 U23155 ( .A(n20318), .ZN(n20257) );
  INV_X1 U23156 ( .A(n20256), .ZN(n20636) );
  AOI21_X1 U23157 ( .B1(n20257), .B2(n20636), .A(n20278), .ZN(n20258) );
  OAI22_X1 U23158 ( .A1(n20258), .A2(n20719), .B1(n20259), .B2(n11773), .ZN(
        n20277) );
  AOI22_X1 U23159 ( .A1(n20713), .A2(n20278), .B1(n20277), .B2(n20712), .ZN(
        n20264) );
  OAI21_X1 U23160 ( .B1(n20326), .B2(n20260), .A(n20259), .ZN(n20262) );
  OAI21_X1 U23161 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n20590), .A(
        n20261), .ZN(n20321) );
  NAND2_X1 U23162 ( .A1(n20262), .A2(n20717), .ZN(n20280) );
  AOI22_X1 U23163 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20280), .B1(
        n20279), .B2(n20722), .ZN(n20263) );
  OAI211_X1 U23164 ( .C1(n20725), .C2(n20296), .A(n20264), .B(n20263), .ZN(
        P1_U3041) );
  INV_X1 U23165 ( .A(n20646), .ZN(n20731) );
  AOI22_X1 U23166 ( .A1(n20727), .A2(n20278), .B1(n20277), .B2(n20726), .ZN(
        n20266) );
  AOI22_X1 U23167 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20280), .B1(
        n20279), .B2(n20728), .ZN(n20265) );
  OAI211_X1 U23168 ( .C1(n20731), .C2(n20296), .A(n20266), .B(n20265), .ZN(
        P1_U3042) );
  INV_X1 U23169 ( .A(n20734), .ZN(n20687) );
  AOI22_X1 U23170 ( .A1(n20733), .A2(n20278), .B1(n20277), .B2(n20732), .ZN(
        n20268) );
  AOI22_X1 U23171 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20280), .B1(
        n20279), .B2(n20684), .ZN(n20267) );
  OAI211_X1 U23172 ( .C1(n20687), .C2(n20296), .A(n20268), .B(n20267), .ZN(
        P1_U3043) );
  INV_X1 U23173 ( .A(n20740), .ZN(n20691) );
  AOI22_X1 U23174 ( .A1(n20739), .A2(n20278), .B1(n20277), .B2(n20738), .ZN(
        n20270) );
  AOI22_X1 U23175 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20280), .B1(
        n20279), .B2(n20688), .ZN(n20269) );
  OAI211_X1 U23176 ( .C1(n20691), .C2(n20296), .A(n20270), .B(n20269), .ZN(
        P1_U3044) );
  INV_X1 U23177 ( .A(n20654), .ZN(n20749) );
  AOI22_X1 U23178 ( .A1(n20278), .A2(n20745), .B1(n20277), .B2(n20744), .ZN(
        n20272) );
  AOI22_X1 U23179 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20280), .B1(
        n20279), .B2(n20746), .ZN(n20271) );
  OAI211_X1 U23180 ( .C1(n20749), .C2(n20296), .A(n20272), .B(n20271), .ZN(
        P1_U3045) );
  INV_X1 U23181 ( .A(n20752), .ZN(n20697) );
  AOI22_X1 U23182 ( .A1(n20751), .A2(n20278), .B1(n20277), .B2(n20750), .ZN(
        n20274) );
  AOI22_X1 U23183 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20280), .B1(
        n20279), .B2(n20694), .ZN(n20273) );
  OAI211_X1 U23184 ( .C1(n20697), .C2(n20296), .A(n20274), .B(n20273), .ZN(
        P1_U3046) );
  INV_X1 U23185 ( .A(n20758), .ZN(n20701) );
  AOI22_X1 U23186 ( .A1(n20757), .A2(n20278), .B1(n20756), .B2(n20277), .ZN(
        n20276) );
  AOI22_X1 U23187 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20280), .B1(
        n20279), .B2(n20698), .ZN(n20275) );
  OAI211_X1 U23188 ( .C1(n20701), .C2(n20296), .A(n20276), .B(n20275), .ZN(
        P1_U3047) );
  INV_X1 U23189 ( .A(n20664), .ZN(n20774) );
  AOI22_X1 U23190 ( .A1(n20278), .A2(n20767), .B1(n20277), .B2(n20764), .ZN(
        n20282) );
  AOI22_X1 U23191 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20280), .B1(
        n20279), .B2(n20768), .ZN(n20281) );
  OAI211_X1 U23192 ( .C1(n20774), .C2(n20296), .A(n20282), .B(n20281), .ZN(
        P1_U3048) );
  NAND2_X1 U23193 ( .A1(n20296), .A2(n20721), .ZN(n20284) );
  OAI21_X1 U23194 ( .B1(n20342), .B2(n20284), .A(n20577), .ZN(n20286) );
  NOR2_X1 U23195 ( .A1(n20318), .A2(n20455), .ZN(n20288) );
  INV_X1 U23196 ( .A(n20712), .ZN(n20594) );
  NAND3_X1 U23197 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20546), .A3(
        n12312), .ZN(n20322) );
  NOR2_X1 U23198 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20322), .ZN(
        n20307) );
  INV_X1 U23199 ( .A(n20307), .ZN(n20292) );
  OAI22_X1 U23200 ( .A1(n20296), .A2(n20645), .B1(n20583), .B2(n20292), .ZN(
        n20285) );
  INV_X1 U23201 ( .A(n20285), .ZN(n20291) );
  INV_X1 U23202 ( .A(n20286), .ZN(n20289) );
  NOR2_X1 U23203 ( .A1(n10297), .A2(n11773), .ZN(n20402) );
  AOI211_X1 U23204 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20292), .A(n20402), 
        .B(n20458), .ZN(n20287) );
  AOI22_X1 U23205 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20309), .B1(
        n20342), .B2(n20642), .ZN(n20290) );
  OAI211_X1 U23206 ( .C1(n20312), .C2(n20594), .A(n20291), .B(n20290), .ZN(
        P1_U3049) );
  OAI22_X1 U23207 ( .A1(n20296), .A2(n20649), .B1(n20595), .B2(n20292), .ZN(
        n20293) );
  INV_X1 U23208 ( .A(n20293), .ZN(n20295) );
  AOI22_X1 U23209 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20309), .B1(
        n20342), .B2(n20646), .ZN(n20294) );
  OAI211_X1 U23210 ( .C1(n20312), .C2(n20599), .A(n20295), .B(n20294), .ZN(
        P1_U3050) );
  INV_X1 U23211 ( .A(n20732), .ZN(n20604) );
  AOI22_X1 U23212 ( .A1(n20342), .A2(n20734), .B1(n20733), .B2(n20307), .ZN(
        n20298) );
  AOI22_X1 U23213 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20309), .B1(
        n20308), .B2(n20684), .ZN(n20297) );
  OAI211_X1 U23214 ( .C1(n20312), .C2(n20604), .A(n20298), .B(n20297), .ZN(
        P1_U3051) );
  INV_X1 U23215 ( .A(n20738), .ZN(n20609) );
  AOI22_X1 U23216 ( .A1(n20342), .A2(n20740), .B1(n20739), .B2(n20307), .ZN(
        n20300) );
  AOI22_X1 U23217 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20309), .B1(
        n20308), .B2(n20688), .ZN(n20299) );
  OAI211_X1 U23218 ( .C1(n20312), .C2(n20609), .A(n20300), .B(n20299), .ZN(
        P1_U3052) );
  AOI22_X1 U23219 ( .A1(n20342), .A2(n20654), .B1(n20745), .B2(n20307), .ZN(
        n20302) );
  AOI22_X1 U23220 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20309), .B1(
        n20308), .B2(n20746), .ZN(n20301) );
  OAI211_X1 U23221 ( .C1(n20312), .C2(n20614), .A(n20302), .B(n20301), .ZN(
        P1_U3053) );
  AOI22_X1 U23222 ( .A1(n20342), .A2(n20752), .B1(n20751), .B2(n20307), .ZN(
        n20304) );
  AOI22_X1 U23223 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20309), .B1(
        n20308), .B2(n20694), .ZN(n20303) );
  OAI211_X1 U23224 ( .C1(n20312), .C2(n20619), .A(n20304), .B(n20303), .ZN(
        P1_U3054) );
  INV_X1 U23225 ( .A(n20756), .ZN(n20624) );
  AOI22_X1 U23226 ( .A1(n20342), .A2(n20758), .B1(n20757), .B2(n20307), .ZN(
        n20306) );
  AOI22_X1 U23227 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20309), .B1(
        n20308), .B2(n20698), .ZN(n20305) );
  OAI211_X1 U23228 ( .C1(n20312), .C2(n20624), .A(n20306), .B(n20305), .ZN(
        P1_U3055) );
  AOI22_X1 U23229 ( .A1(n20342), .A2(n20664), .B1(n20767), .B2(n20307), .ZN(
        n20311) );
  AOI22_X1 U23230 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20309), .B1(
        n20308), .B2(n20768), .ZN(n20310) );
  OAI211_X1 U23231 ( .C1(n20312), .C2(n20632), .A(n20311), .B(n20310), .ZN(
        P1_U3056) );
  INV_X1 U23232 ( .A(n20322), .ZN(n20319) );
  INV_X1 U23233 ( .A(n20715), .ZN(n20313) );
  AOI21_X1 U23234 ( .B1(n20314), .B2(n20313), .A(n20719), .ZN(n20320) );
  AND2_X1 U23235 ( .A1(n20315), .A2(n9664), .ZN(n20709) );
  INV_X1 U23236 ( .A(n20709), .ZN(n20317) );
  NOR2_X1 U23237 ( .A1(n20547), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20341) );
  INV_X1 U23238 ( .A(n20341), .ZN(n20316) );
  OAI21_X1 U23239 ( .B1(n20318), .B2(n20317), .A(n20316), .ZN(n20324) );
  AOI22_X1 U23240 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20319), .B1(n20320), 
        .B2(n20324), .ZN(n20346) );
  AOI22_X1 U23241 ( .A1(n20342), .A2(n20722), .B1(n20713), .B2(n20341), .ZN(
        n20328) );
  INV_X1 U23242 ( .A(n20320), .ZN(n20325) );
  AOI21_X1 U23243 ( .B1(n20719), .B2(n20322), .A(n20321), .ZN(n20323) );
  OAI21_X1 U23244 ( .B1(n20325), .B2(n20324), .A(n20323), .ZN(n20343) );
  AOI22_X1 U23245 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20343), .B1(
        n20371), .B2(n20642), .ZN(n20327) );
  OAI211_X1 U23246 ( .C1(n20346), .C2(n20594), .A(n20328), .B(n20327), .ZN(
        P1_U3057) );
  AOI22_X1 U23247 ( .A1(n20371), .A2(n20646), .B1(n20727), .B2(n20341), .ZN(
        n20330) );
  AOI22_X1 U23248 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20343), .B1(
        n20342), .B2(n20728), .ZN(n20329) );
  OAI211_X1 U23249 ( .C1(n20346), .C2(n20599), .A(n20330), .B(n20329), .ZN(
        P1_U3058) );
  AOI22_X1 U23250 ( .A1(n20342), .A2(n20684), .B1(n20733), .B2(n20341), .ZN(
        n20332) );
  AOI22_X1 U23251 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20343), .B1(
        n20371), .B2(n20734), .ZN(n20331) );
  OAI211_X1 U23252 ( .C1(n20346), .C2(n20604), .A(n20332), .B(n20331), .ZN(
        P1_U3059) );
  AOI22_X1 U23253 ( .A1(n20342), .A2(n20688), .B1(n20739), .B2(n20341), .ZN(
        n20334) );
  AOI22_X1 U23254 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20343), .B1(
        n20371), .B2(n20740), .ZN(n20333) );
  OAI211_X1 U23255 ( .C1(n20346), .C2(n20609), .A(n20334), .B(n20333), .ZN(
        P1_U3060) );
  AOI22_X1 U23256 ( .A1(n20342), .A2(n20746), .B1(n20745), .B2(n20341), .ZN(
        n20336) );
  AOI22_X1 U23257 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20343), .B1(
        n20371), .B2(n20654), .ZN(n20335) );
  OAI211_X1 U23258 ( .C1(n20346), .C2(n20614), .A(n20336), .B(n20335), .ZN(
        P1_U3061) );
  AOI22_X1 U23259 ( .A1(n20371), .A2(n20752), .B1(n20751), .B2(n20341), .ZN(
        n20338) );
  AOI22_X1 U23260 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20343), .B1(
        n20342), .B2(n20694), .ZN(n20337) );
  OAI211_X1 U23261 ( .C1(n20346), .C2(n20619), .A(n20338), .B(n20337), .ZN(
        P1_U3062) );
  AOI22_X1 U23262 ( .A1(n20371), .A2(n20758), .B1(n20757), .B2(n20341), .ZN(
        n20340) );
  AOI22_X1 U23263 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20343), .B1(
        n20342), .B2(n20698), .ZN(n20339) );
  OAI211_X1 U23264 ( .C1(n20346), .C2(n20624), .A(n20340), .B(n20339), .ZN(
        P1_U3063) );
  AOI22_X1 U23265 ( .A1(n20342), .A2(n20768), .B1(n20767), .B2(n20341), .ZN(
        n20345) );
  AOI22_X1 U23266 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20343), .B1(
        n20371), .B2(n20664), .ZN(n20344) );
  OAI211_X1 U23267 ( .C1(n20346), .C2(n20632), .A(n20345), .B(n20344), .ZN(
        P1_U3064) );
  INV_X1 U23268 ( .A(n20453), .ZN(n20575) );
  NAND3_X1 U23269 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20546), .A3(
        n20582), .ZN(n20375) );
  NOR2_X1 U23270 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20375), .ZN(
        n20370) );
  NOR2_X1 U23271 ( .A1(n10245), .A2(n20347), .ZN(n20428) );
  NAND3_X1 U23272 ( .A1(n20428), .A2(n20455), .A3(n20721), .ZN(n20348) );
  OAI21_X1 U23273 ( .B1(n20672), .B2(n20349), .A(n20348), .ZN(n20369) );
  AOI22_X1 U23274 ( .A1(n20713), .A2(n20370), .B1(n20712), .B2(n20369), .ZN(
        n20356) );
  INV_X1 U23275 ( .A(n20371), .ZN(n20350) );
  AOI21_X1 U23276 ( .B1(n20350), .B2(n20398), .A(n20874), .ZN(n20351) );
  AOI21_X1 U23277 ( .B1(n20428), .B2(n20455), .A(n20351), .ZN(n20352) );
  NOR2_X1 U23278 ( .A1(n20352), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20354) );
  AOI22_X1 U23279 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20372), .B1(
        n20371), .B2(n20722), .ZN(n20355) );
  OAI211_X1 U23280 ( .C1(n20725), .C2(n20398), .A(n20356), .B(n20355), .ZN(
        P1_U3065) );
  AOI22_X1 U23281 ( .A1(n20727), .A2(n20370), .B1(n20726), .B2(n20369), .ZN(
        n20358) );
  AOI22_X1 U23282 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20372), .B1(
        n20371), .B2(n20728), .ZN(n20357) );
  OAI211_X1 U23283 ( .C1(n20731), .C2(n20398), .A(n20358), .B(n20357), .ZN(
        P1_U3066) );
  AOI22_X1 U23284 ( .A1(n20733), .A2(n20370), .B1(n20732), .B2(n20369), .ZN(
        n20360) );
  AOI22_X1 U23285 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20372), .B1(
        n20371), .B2(n20684), .ZN(n20359) );
  OAI211_X1 U23286 ( .C1(n20687), .C2(n20398), .A(n20360), .B(n20359), .ZN(
        P1_U3067) );
  AOI22_X1 U23287 ( .A1(n20739), .A2(n20370), .B1(n20738), .B2(n20369), .ZN(
        n20362) );
  AOI22_X1 U23288 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20372), .B1(
        n20371), .B2(n20688), .ZN(n20361) );
  OAI211_X1 U23289 ( .C1(n20691), .C2(n20398), .A(n20362), .B(n20361), .ZN(
        P1_U3068) );
  AOI22_X1 U23290 ( .A1(n20745), .A2(n20370), .B1(n20744), .B2(n20369), .ZN(
        n20364) );
  AOI22_X1 U23291 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20372), .B1(
        n20371), .B2(n20746), .ZN(n20363) );
  OAI211_X1 U23292 ( .C1(n20749), .C2(n20398), .A(n20364), .B(n20363), .ZN(
        P1_U3069) );
  AOI22_X1 U23293 ( .A1(n20751), .A2(n20370), .B1(n20750), .B2(n20369), .ZN(
        n20366) );
  AOI22_X1 U23294 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20372), .B1(
        n20371), .B2(n20694), .ZN(n20365) );
  OAI211_X1 U23295 ( .C1(n20697), .C2(n20398), .A(n20366), .B(n20365), .ZN(
        P1_U3070) );
  AOI22_X1 U23296 ( .A1(n20757), .A2(n20370), .B1(n20756), .B2(n20369), .ZN(
        n20368) );
  AOI22_X1 U23297 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20372), .B1(
        n20371), .B2(n20698), .ZN(n20367) );
  OAI211_X1 U23298 ( .C1(n20701), .C2(n20398), .A(n20368), .B(n20367), .ZN(
        P1_U3071) );
  AOI22_X1 U23299 ( .A1(n20767), .A2(n20370), .B1(n20764), .B2(n20369), .ZN(
        n20374) );
  AOI22_X1 U23300 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20372), .B1(
        n20371), .B2(n20768), .ZN(n20373) );
  OAI211_X1 U23301 ( .C1(n20774), .C2(n20398), .A(n20374), .B(n20373), .ZN(
        P1_U3072) );
  NOR2_X1 U23302 ( .A1(n20634), .A2(n20375), .ZN(n20394) );
  AOI21_X1 U23303 ( .B1(n20428), .B2(n20636), .A(n20394), .ZN(n20376) );
  OAI22_X1 U23304 ( .A1(n20376), .A2(n20719), .B1(n20375), .B2(n11773), .ZN(
        n20393) );
  AOI22_X1 U23305 ( .A1(n20713), .A2(n20394), .B1(n20393), .B2(n20712), .ZN(
        n20380) );
  INV_X1 U23306 ( .A(n20375), .ZN(n20378) );
  OAI21_X1 U23307 ( .B1(n20426), .B2(n20874), .A(n20376), .ZN(n20377) );
  OAI221_X1 U23308 ( .B1(n20721), .B2(n20378), .C1(n20719), .C2(n20377), .A(
        n20717), .ZN(n20395) );
  AOI22_X1 U23309 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20395), .B1(
        n20421), .B2(n20642), .ZN(n20379) );
  OAI211_X1 U23310 ( .C1(n20645), .C2(n20398), .A(n20380), .B(n20379), .ZN(
        P1_U3073) );
  AOI22_X1 U23311 ( .A1(n20727), .A2(n20394), .B1(n20393), .B2(n20726), .ZN(
        n20382) );
  AOI22_X1 U23312 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20395), .B1(
        n20421), .B2(n20646), .ZN(n20381) );
  OAI211_X1 U23313 ( .C1(n20649), .C2(n20398), .A(n20382), .B(n20381), .ZN(
        P1_U3074) );
  INV_X1 U23314 ( .A(n20684), .ZN(n20737) );
  AOI22_X1 U23315 ( .A1(n20733), .A2(n20394), .B1(n20393), .B2(n20732), .ZN(
        n20384) );
  AOI22_X1 U23316 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20395), .B1(
        n20421), .B2(n20734), .ZN(n20383) );
  OAI211_X1 U23317 ( .C1(n20737), .C2(n20398), .A(n20384), .B(n20383), .ZN(
        P1_U3075) );
  INV_X1 U23318 ( .A(n20688), .ZN(n20743) );
  AOI22_X1 U23319 ( .A1(n20739), .A2(n20394), .B1(n20738), .B2(n20393), .ZN(
        n20386) );
  AOI22_X1 U23320 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20395), .B1(
        n20421), .B2(n20740), .ZN(n20385) );
  OAI211_X1 U23321 ( .C1(n20743), .C2(n20398), .A(n20386), .B(n20385), .ZN(
        P1_U3076) );
  INV_X1 U23322 ( .A(n20746), .ZN(n20657) );
  AOI22_X1 U23323 ( .A1(n20745), .A2(n20394), .B1(n20393), .B2(n20744), .ZN(
        n20388) );
  AOI22_X1 U23324 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20395), .B1(
        n20421), .B2(n20654), .ZN(n20387) );
  OAI211_X1 U23325 ( .C1(n20657), .C2(n20398), .A(n20388), .B(n20387), .ZN(
        P1_U3077) );
  INV_X1 U23326 ( .A(n20694), .ZN(n20755) );
  AOI22_X1 U23327 ( .A1(n20751), .A2(n20394), .B1(n20393), .B2(n20750), .ZN(
        n20390) );
  AOI22_X1 U23328 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20395), .B1(
        n20421), .B2(n20752), .ZN(n20389) );
  OAI211_X1 U23329 ( .C1(n20755), .C2(n20398), .A(n20390), .B(n20389), .ZN(
        P1_U3078) );
  AOI22_X1 U23330 ( .A1(n20757), .A2(n20394), .B1(n20756), .B2(n20393), .ZN(
        n20392) );
  AOI22_X1 U23331 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20395), .B1(
        n20421), .B2(n20758), .ZN(n20391) );
  OAI211_X1 U23332 ( .C1(n20763), .C2(n20398), .A(n20392), .B(n20391), .ZN(
        P1_U3079) );
  INV_X1 U23333 ( .A(n20768), .ZN(n20669) );
  AOI22_X1 U23334 ( .A1(n20767), .A2(n20394), .B1(n20393), .B2(n20764), .ZN(
        n20397) );
  AOI22_X1 U23335 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20395), .B1(
        n20421), .B2(n20664), .ZN(n20396) );
  OAI211_X1 U23336 ( .C1(n20669), .C2(n20398), .A(n20397), .B(n20396), .ZN(
        P1_U3080) );
  INV_X1 U23337 ( .A(n20421), .ZN(n20399) );
  NAND2_X1 U23338 ( .A1(n20399), .A2(n20721), .ZN(n20400) );
  OAI21_X1 U23339 ( .B1(n20400), .B2(n20449), .A(n20577), .ZN(n20404) );
  AND2_X1 U23340 ( .A1(n20428), .A2(n20674), .ZN(n20401) );
  INV_X1 U23341 ( .A(n20672), .ZN(n20581) );
  INV_X1 U23342 ( .A(n20431), .ZN(n20429) );
  NOR2_X1 U23343 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20429), .ZN(
        n20420) );
  AOI22_X1 U23344 ( .A1(n20421), .A2(n20722), .B1(n20713), .B2(n20420), .ZN(
        n20407) );
  INV_X1 U23345 ( .A(n20401), .ZN(n20403) );
  AOI21_X1 U23346 ( .B1(n20404), .B2(n20403), .A(n20402), .ZN(n20405) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20422), .B1(
        n20449), .B2(n20642), .ZN(n20406) );
  OAI211_X1 U23348 ( .C1(n20425), .C2(n20594), .A(n20407), .B(n20406), .ZN(
        P1_U3081) );
  AOI22_X1 U23349 ( .A1(n20421), .A2(n20728), .B1(n20420), .B2(n20727), .ZN(
        n20409) );
  AOI22_X1 U23350 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20422), .B1(
        n20449), .B2(n20646), .ZN(n20408) );
  OAI211_X1 U23351 ( .C1(n20425), .C2(n20599), .A(n20409), .B(n20408), .ZN(
        P1_U3082) );
  AOI22_X1 U23352 ( .A1(n20421), .A2(n20684), .B1(n20733), .B2(n20420), .ZN(
        n20411) );
  AOI22_X1 U23353 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20422), .B1(
        n20449), .B2(n20734), .ZN(n20410) );
  OAI211_X1 U23354 ( .C1(n20425), .C2(n20604), .A(n20411), .B(n20410), .ZN(
        P1_U3083) );
  AOI22_X1 U23355 ( .A1(n20449), .A2(n20740), .B1(n20420), .B2(n20739), .ZN(
        n20413) );
  AOI22_X1 U23356 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20422), .B1(
        n20421), .B2(n20688), .ZN(n20412) );
  OAI211_X1 U23357 ( .C1(n20425), .C2(n20609), .A(n20413), .B(n20412), .ZN(
        P1_U3084) );
  AOI22_X1 U23358 ( .A1(n20421), .A2(n20746), .B1(n20745), .B2(n20420), .ZN(
        n20415) );
  AOI22_X1 U23359 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20422), .B1(
        n20449), .B2(n20654), .ZN(n20414) );
  OAI211_X1 U23360 ( .C1(n20425), .C2(n20614), .A(n20415), .B(n20414), .ZN(
        P1_U3085) );
  AOI22_X1 U23361 ( .A1(n20449), .A2(n20752), .B1(n20420), .B2(n20751), .ZN(
        n20417) );
  AOI22_X1 U23362 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20422), .B1(
        n20421), .B2(n20694), .ZN(n20416) );
  OAI211_X1 U23363 ( .C1(n20425), .C2(n20619), .A(n20417), .B(n20416), .ZN(
        P1_U3086) );
  AOI22_X1 U23364 ( .A1(n20449), .A2(n20758), .B1(n20420), .B2(n20757), .ZN(
        n20419) );
  AOI22_X1 U23365 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20422), .B1(
        n20421), .B2(n20698), .ZN(n20418) );
  OAI211_X1 U23366 ( .C1(n20425), .C2(n20624), .A(n20419), .B(n20418), .ZN(
        P1_U3087) );
  AOI22_X1 U23367 ( .A1(n20449), .A2(n20664), .B1(n20767), .B2(n20420), .ZN(
        n20424) );
  AOI22_X1 U23368 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20422), .B1(
        n20421), .B2(n20768), .ZN(n20423) );
  OAI211_X1 U23369 ( .C1(n20425), .C2(n20632), .A(n20424), .B(n20423), .ZN(
        P1_U3088) );
  INV_X1 U23370 ( .A(n20427), .ZN(n20448) );
  AOI21_X1 U23371 ( .B1(n20428), .B2(n20709), .A(n20448), .ZN(n20430) );
  OAI22_X1 U23372 ( .A1(n20430), .A2(n20719), .B1(n20429), .B2(n11773), .ZN(
        n20447) );
  AOI22_X1 U23373 ( .A1(n20713), .A2(n20448), .B1(n20712), .B2(n20447), .ZN(
        n20434) );
  OAI21_X1 U23374 ( .B1(n20432), .B2(n20431), .A(n20717), .ZN(n20450) );
  AOI22_X1 U23375 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20450), .B1(
        n20449), .B2(n20722), .ZN(n20433) );
  OAI211_X1 U23376 ( .C1(n20725), .C2(n20459), .A(n20434), .B(n20433), .ZN(
        P1_U3089) );
  AOI22_X1 U23377 ( .A1(n20727), .A2(n20448), .B1(n20726), .B2(n20447), .ZN(
        n20436) );
  AOI22_X1 U23378 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20450), .B1(
        n20449), .B2(n20728), .ZN(n20435) );
  OAI211_X1 U23379 ( .C1(n20731), .C2(n20459), .A(n20436), .B(n20435), .ZN(
        P1_U3090) );
  AOI22_X1 U23380 ( .A1(n20733), .A2(n20448), .B1(n20732), .B2(n20447), .ZN(
        n20438) );
  AOI22_X1 U23381 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20450), .B1(
        n20449), .B2(n20684), .ZN(n20437) );
  OAI211_X1 U23382 ( .C1(n20687), .C2(n20459), .A(n20438), .B(n20437), .ZN(
        P1_U3091) );
  AOI22_X1 U23383 ( .A1(n20739), .A2(n20448), .B1(n20738), .B2(n20447), .ZN(
        n20440) );
  AOI22_X1 U23384 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20450), .B1(
        n20449), .B2(n20688), .ZN(n20439) );
  OAI211_X1 U23385 ( .C1(n20691), .C2(n20459), .A(n20440), .B(n20439), .ZN(
        P1_U3092) );
  AOI22_X1 U23386 ( .A1(n20745), .A2(n20448), .B1(n20744), .B2(n20447), .ZN(
        n20442) );
  AOI22_X1 U23387 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20450), .B1(
        n20449), .B2(n20746), .ZN(n20441) );
  OAI211_X1 U23388 ( .C1(n20749), .C2(n20459), .A(n20442), .B(n20441), .ZN(
        P1_U3093) );
  AOI22_X1 U23389 ( .A1(n20751), .A2(n20448), .B1(n20750), .B2(n20447), .ZN(
        n20444) );
  AOI22_X1 U23390 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20450), .B1(
        n20449), .B2(n20694), .ZN(n20443) );
  OAI211_X1 U23391 ( .C1(n20697), .C2(n20459), .A(n20444), .B(n20443), .ZN(
        P1_U3094) );
  AOI22_X1 U23392 ( .A1(n20757), .A2(n20448), .B1(n20756), .B2(n20447), .ZN(
        n20446) );
  AOI22_X1 U23393 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20450), .B1(
        n20449), .B2(n20698), .ZN(n20445) );
  OAI211_X1 U23394 ( .C1(n20701), .C2(n20459), .A(n20446), .B(n20445), .ZN(
        P1_U3095) );
  AOI22_X1 U23395 ( .A1(n20767), .A2(n20448), .B1(n20764), .B2(n20447), .ZN(
        n20452) );
  AOI22_X1 U23396 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20450), .B1(
        n20449), .B2(n20768), .ZN(n20451) );
  OAI211_X1 U23397 ( .C1(n20774), .C2(n20459), .A(n20452), .B(n20451), .ZN(
        P1_U3096) );
  NAND3_X1 U23398 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12312), .A3(
        n20582), .ZN(n20484) );
  NOR2_X1 U23399 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20484), .ZN(
        n20479) );
  AND2_X1 U23400 ( .A1(n20454), .A2(n10245), .ZN(n20548) );
  AOI21_X1 U23401 ( .B1(n20548), .B2(n20455), .A(n20479), .ZN(n20461) );
  AND2_X1 U23402 ( .A1(n20456), .A2(n20512), .ZN(n20580) );
  INV_X1 U23403 ( .A(n20580), .ZN(n20586) );
  OAI22_X1 U23404 ( .A1(n20461), .A2(n20719), .B1(n20586), .B2(n20457), .ZN(
        n20478) );
  AOI22_X1 U23405 ( .A1(n20713), .A2(n20479), .B1(n20478), .B2(n20712), .ZN(
        n20465) );
  INV_X1 U23406 ( .A(n20458), .ZN(n20516) );
  INV_X1 U23407 ( .A(n20507), .ZN(n20460) );
  OAI21_X1 U23408 ( .B1(n20460), .B2(n20480), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20462) );
  NAND2_X1 U23409 ( .A1(n20462), .A2(n20461), .ZN(n20463) );
  AOI22_X1 U23410 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20481), .B1(
        n20480), .B2(n20722), .ZN(n20464) );
  OAI211_X1 U23411 ( .C1(n20725), .C2(n20507), .A(n20465), .B(n20464), .ZN(
        P1_U3097) );
  AOI22_X1 U23412 ( .A1(n20727), .A2(n20479), .B1(n20478), .B2(n20726), .ZN(
        n20467) );
  AOI22_X1 U23413 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20481), .B1(
        n20480), .B2(n20728), .ZN(n20466) );
  OAI211_X1 U23414 ( .C1(n20731), .C2(n20507), .A(n20467), .B(n20466), .ZN(
        P1_U3098) );
  AOI22_X1 U23415 ( .A1(n20733), .A2(n20479), .B1(n20478), .B2(n20732), .ZN(
        n20469) );
  AOI22_X1 U23416 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20481), .B1(
        n20480), .B2(n20684), .ZN(n20468) );
  OAI211_X1 U23417 ( .C1(n20687), .C2(n20507), .A(n20469), .B(n20468), .ZN(
        P1_U3099) );
  AOI22_X1 U23418 ( .A1(n20739), .A2(n20479), .B1(n20478), .B2(n20738), .ZN(
        n20471) );
  AOI22_X1 U23419 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20481), .B1(
        n20480), .B2(n20688), .ZN(n20470) );
  OAI211_X1 U23420 ( .C1(n20691), .C2(n20507), .A(n20471), .B(n20470), .ZN(
        P1_U3100) );
  AOI22_X1 U23421 ( .A1(n20479), .A2(n20745), .B1(n20478), .B2(n20744), .ZN(
        n20473) );
  AOI22_X1 U23422 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20481), .B1(
        n20480), .B2(n20746), .ZN(n20472) );
  OAI211_X1 U23423 ( .C1(n20749), .C2(n20507), .A(n20473), .B(n20472), .ZN(
        P1_U3101) );
  AOI22_X1 U23424 ( .A1(n20751), .A2(n20479), .B1(n20478), .B2(n20750), .ZN(
        n20475) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20481), .B1(
        n20480), .B2(n20694), .ZN(n20474) );
  OAI211_X1 U23426 ( .C1(n20697), .C2(n20507), .A(n20475), .B(n20474), .ZN(
        P1_U3102) );
  AOI22_X1 U23427 ( .A1(n20757), .A2(n20479), .B1(n20756), .B2(n20478), .ZN(
        n20477) );
  AOI22_X1 U23428 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20481), .B1(
        n20480), .B2(n20698), .ZN(n20476) );
  OAI211_X1 U23429 ( .C1(n20701), .C2(n20507), .A(n20477), .B(n20476), .ZN(
        P1_U3103) );
  AOI22_X1 U23430 ( .A1(n20479), .A2(n20767), .B1(n20478), .B2(n20764), .ZN(
        n20483) );
  AOI22_X1 U23431 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20481), .B1(
        n20480), .B2(n20768), .ZN(n20482) );
  OAI211_X1 U23432 ( .C1(n20774), .C2(n20507), .A(n20483), .B(n20482), .ZN(
        P1_U3104) );
  NOR2_X1 U23433 ( .A1(n20634), .A2(n20484), .ZN(n20503) );
  AOI21_X1 U23434 ( .B1(n20548), .B2(n20636), .A(n20503), .ZN(n20485) );
  OAI22_X1 U23435 ( .A1(n20485), .A2(n20719), .B1(n20484), .B2(n11773), .ZN(
        n20502) );
  AOI22_X1 U23436 ( .A1(n20713), .A2(n20503), .B1(n20502), .B2(n20712), .ZN(
        n20489) );
  INV_X1 U23437 ( .A(n20484), .ZN(n20487) );
  OAI21_X1 U23438 ( .B1(n20554), .B2(n20874), .A(n20485), .ZN(n20486) );
  OAI221_X1 U23439 ( .B1(n20721), .B2(n20487), .C1(n20719), .C2(n20486), .A(
        n20717), .ZN(n20504) );
  AOI22_X1 U23440 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20504), .B1(
        n20541), .B2(n20642), .ZN(n20488) );
  OAI211_X1 U23441 ( .C1(n20645), .C2(n20507), .A(n20489), .B(n20488), .ZN(
        P1_U3105) );
  AOI22_X1 U23442 ( .A1(n20727), .A2(n20503), .B1(n20502), .B2(n20726), .ZN(
        n20491) );
  AOI22_X1 U23443 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20504), .B1(
        n20541), .B2(n20646), .ZN(n20490) );
  OAI211_X1 U23444 ( .C1(n20649), .C2(n20507), .A(n20491), .B(n20490), .ZN(
        P1_U3106) );
  AOI22_X1 U23445 ( .A1(n20733), .A2(n20503), .B1(n20502), .B2(n20732), .ZN(
        n20493) );
  AOI22_X1 U23446 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20504), .B1(
        n20541), .B2(n20734), .ZN(n20492) );
  OAI211_X1 U23447 ( .C1(n20737), .C2(n20507), .A(n20493), .B(n20492), .ZN(
        P1_U3107) );
  AOI22_X1 U23448 ( .A1(n20739), .A2(n20503), .B1(n20502), .B2(n20738), .ZN(
        n20495) );
  AOI22_X1 U23449 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20504), .B1(
        n20541), .B2(n20740), .ZN(n20494) );
  OAI211_X1 U23450 ( .C1(n20743), .C2(n20507), .A(n20495), .B(n20494), .ZN(
        P1_U3108) );
  AOI22_X1 U23451 ( .A1(n20503), .A2(n20745), .B1(n20502), .B2(n20744), .ZN(
        n20497) );
  AOI22_X1 U23452 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20504), .B1(
        n20541), .B2(n20654), .ZN(n20496) );
  OAI211_X1 U23453 ( .C1(n20657), .C2(n20507), .A(n20497), .B(n20496), .ZN(
        P1_U3109) );
  AOI22_X1 U23454 ( .A1(n20751), .A2(n20503), .B1(n20502), .B2(n20750), .ZN(
        n20499) );
  AOI22_X1 U23455 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20504), .B1(
        n20541), .B2(n20752), .ZN(n20498) );
  OAI211_X1 U23456 ( .C1(n20755), .C2(n20507), .A(n20499), .B(n20498), .ZN(
        P1_U3110) );
  AOI22_X1 U23457 ( .A1(n20757), .A2(n20503), .B1(n20756), .B2(n20502), .ZN(
        n20501) );
  AOI22_X1 U23458 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20504), .B1(
        n20541), .B2(n20758), .ZN(n20500) );
  OAI211_X1 U23459 ( .C1(n20763), .C2(n20507), .A(n20501), .B(n20500), .ZN(
        P1_U3111) );
  AOI22_X1 U23460 ( .A1(n20503), .A2(n20767), .B1(n20502), .B2(n20764), .ZN(
        n20506) );
  AOI22_X1 U23461 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20504), .B1(
        n20541), .B2(n20664), .ZN(n20505) );
  OAI211_X1 U23462 ( .C1(n20669), .C2(n20507), .A(n20506), .B(n20505), .ZN(
        P1_U3112) );
  INV_X1 U23463 ( .A(n20541), .ZN(n20510) );
  NAND3_X1 U23464 ( .A1(n20510), .A2(n20721), .A3(n20574), .ZN(n20511) );
  NAND2_X1 U23465 ( .A1(n20511), .A2(n20577), .ZN(n20519) );
  AND2_X1 U23466 ( .A1(n20548), .A2(n20674), .ZN(n20515) );
  OR2_X1 U23467 ( .A1(n20512), .A2(n20546), .ZN(n20673) );
  INV_X1 U23468 ( .A(n20673), .ZN(n20513) );
  NAND3_X1 U23469 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n12312), .ZN(n20550) );
  NOR2_X1 U23470 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20550), .ZN(
        n20532) );
  AOI22_X1 U23471 ( .A1(n20541), .A2(n20722), .B1(n20713), .B2(n20532), .ZN(
        n20522) );
  INV_X1 U23472 ( .A(n20515), .ZN(n20518) );
  NAND2_X1 U23473 ( .A1(n20673), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20677) );
  OAI211_X1 U23474 ( .C1(n20590), .C2(n20532), .A(n20677), .B(n20516), .ZN(
        n20517) );
  AOI21_X1 U23475 ( .B1(n20519), .B2(n20518), .A(n20517), .ZN(n20520) );
  INV_X1 U23476 ( .A(n20574), .ZN(n20533) );
  AOI22_X1 U23477 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20542), .B1(
        n20533), .B2(n20642), .ZN(n20521) );
  OAI211_X1 U23478 ( .C1(n20545), .C2(n20594), .A(n20522), .B(n20521), .ZN(
        P1_U3113) );
  AOI22_X1 U23479 ( .A1(n20541), .A2(n20728), .B1(n20727), .B2(n20532), .ZN(
        n20524) );
  AOI22_X1 U23480 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20542), .B1(
        n20533), .B2(n20646), .ZN(n20523) );
  OAI211_X1 U23481 ( .C1(n20545), .C2(n20599), .A(n20524), .B(n20523), .ZN(
        P1_U3114) );
  AOI22_X1 U23482 ( .A1(n20541), .A2(n20684), .B1(n20733), .B2(n20532), .ZN(
        n20526) );
  AOI22_X1 U23483 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20542), .B1(
        n20533), .B2(n20734), .ZN(n20525) );
  OAI211_X1 U23484 ( .C1(n20545), .C2(n20604), .A(n20526), .B(n20525), .ZN(
        P1_U3115) );
  INV_X1 U23485 ( .A(n20532), .ZN(n20539) );
  OAI22_X1 U23486 ( .A1(n20574), .A2(n20691), .B1(n20605), .B2(n20539), .ZN(
        n20527) );
  INV_X1 U23487 ( .A(n20527), .ZN(n20529) );
  AOI22_X1 U23488 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20542), .B1(
        n20541), .B2(n20688), .ZN(n20528) );
  OAI211_X1 U23489 ( .C1(n20545), .C2(n20609), .A(n20529), .B(n20528), .ZN(
        P1_U3116) );
  AOI22_X1 U23490 ( .A1(n20541), .A2(n20746), .B1(n20745), .B2(n20532), .ZN(
        n20531) );
  AOI22_X1 U23491 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20542), .B1(
        n20533), .B2(n20654), .ZN(n20530) );
  OAI211_X1 U23492 ( .C1(n20545), .C2(n20614), .A(n20531), .B(n20530), .ZN(
        P1_U3117) );
  AOI22_X1 U23493 ( .A1(n20541), .A2(n20694), .B1(n20751), .B2(n20532), .ZN(
        n20535) );
  AOI22_X1 U23494 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20542), .B1(
        n20533), .B2(n20752), .ZN(n20534) );
  OAI211_X1 U23495 ( .C1(n20545), .C2(n20619), .A(n20535), .B(n20534), .ZN(
        P1_U3118) );
  OAI22_X1 U23496 ( .A1(n20574), .A2(n20701), .B1(n20620), .B2(n20539), .ZN(
        n20536) );
  INV_X1 U23497 ( .A(n20536), .ZN(n20538) );
  AOI22_X1 U23498 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20542), .B1(
        n20541), .B2(n20698), .ZN(n20537) );
  OAI211_X1 U23499 ( .C1(n20545), .C2(n20624), .A(n20538), .B(n20537), .ZN(
        P1_U3119) );
  INV_X1 U23500 ( .A(n20767), .ZN(n20626) );
  OAI22_X1 U23501 ( .A1(n20574), .A2(n20774), .B1(n20626), .B2(n20539), .ZN(
        n20540) );
  INV_X1 U23502 ( .A(n20540), .ZN(n20544) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20542), .B1(
        n20541), .B2(n20768), .ZN(n20543) );
  OAI211_X1 U23504 ( .C1(n20545), .C2(n20632), .A(n20544), .B(n20543), .ZN(
        P1_U3120) );
  NOR2_X1 U23505 ( .A1(n20547), .A2(n20546), .ZN(n20570) );
  AOI21_X1 U23506 ( .B1(n20548), .B2(n20709), .A(n20570), .ZN(n20549) );
  OAI22_X1 U23507 ( .A1(n20549), .A2(n20719), .B1(n20550), .B2(n11773), .ZN(
        n20569) );
  AOI22_X1 U23508 ( .A1(n20713), .A2(n20570), .B1(n20569), .B2(n20712), .ZN(
        n20556) );
  OAI21_X1 U23509 ( .B1(n20554), .B2(n20551), .A(n20550), .ZN(n20552) );
  NAND2_X1 U23510 ( .A1(n20552), .A2(n20717), .ZN(n20571) );
  AOI22_X1 U23511 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20571), .B1(
        n20628), .B2(n20642), .ZN(n20555) );
  OAI211_X1 U23512 ( .C1(n20645), .C2(n20574), .A(n20556), .B(n20555), .ZN(
        P1_U3121) );
  AOI22_X1 U23513 ( .A1(n20727), .A2(n20570), .B1(n20569), .B2(n20726), .ZN(
        n20558) );
  AOI22_X1 U23514 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20571), .B1(
        n20628), .B2(n20646), .ZN(n20557) );
  OAI211_X1 U23515 ( .C1(n20649), .C2(n20574), .A(n20558), .B(n20557), .ZN(
        P1_U3122) );
  AOI22_X1 U23516 ( .A1(n20733), .A2(n20570), .B1(n20569), .B2(n20732), .ZN(
        n20560) );
  AOI22_X1 U23517 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20571), .B1(
        n20628), .B2(n20734), .ZN(n20559) );
  OAI211_X1 U23518 ( .C1(n20737), .C2(n20574), .A(n20560), .B(n20559), .ZN(
        P1_U3123) );
  AOI22_X1 U23519 ( .A1(n20739), .A2(n20570), .B1(n20738), .B2(n20569), .ZN(
        n20562) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20571), .B1(
        n20628), .B2(n20740), .ZN(n20561) );
  OAI211_X1 U23521 ( .C1(n20743), .C2(n20574), .A(n20562), .B(n20561), .ZN(
        P1_U3124) );
  AOI22_X1 U23522 ( .A1(n20745), .A2(n20570), .B1(n20569), .B2(n20744), .ZN(
        n20564) );
  AOI22_X1 U23523 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20571), .B1(
        n20628), .B2(n20654), .ZN(n20563) );
  OAI211_X1 U23524 ( .C1(n20657), .C2(n20574), .A(n20564), .B(n20563), .ZN(
        P1_U3125) );
  AOI22_X1 U23525 ( .A1(n20751), .A2(n20570), .B1(n20569), .B2(n20750), .ZN(
        n20566) );
  AOI22_X1 U23526 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20571), .B1(
        n20628), .B2(n20752), .ZN(n20565) );
  OAI211_X1 U23527 ( .C1(n20755), .C2(n20574), .A(n20566), .B(n20565), .ZN(
        P1_U3126) );
  AOI22_X1 U23528 ( .A1(n20757), .A2(n20570), .B1(n20756), .B2(n20569), .ZN(
        n20568) );
  AOI22_X1 U23529 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20571), .B1(
        n20628), .B2(n20758), .ZN(n20567) );
  OAI211_X1 U23530 ( .C1(n20763), .C2(n20574), .A(n20568), .B(n20567), .ZN(
        P1_U3127) );
  AOI22_X1 U23531 ( .A1(n20767), .A2(n20570), .B1(n20569), .B2(n20764), .ZN(
        n20573) );
  AOI22_X1 U23532 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20571), .B1(
        n20628), .B2(n20664), .ZN(n20572) );
  OAI211_X1 U23533 ( .C1(n20669), .C2(n20574), .A(n20573), .B(n20572), .ZN(
        P1_U3128) );
  INV_X1 U23534 ( .A(n20628), .ZN(n20576) );
  NAND3_X1 U23535 ( .A1(n20576), .A2(n20721), .A3(n20668), .ZN(n20578) );
  NAND2_X1 U23536 ( .A1(n20578), .A2(n20577), .ZN(n20588) );
  OR2_X1 U23537 ( .A1(n10245), .A2(n20579), .ZN(n20635) );
  NOR2_X1 U23538 ( .A1(n20635), .A2(n20674), .ZN(n20585) );
  NAND3_X1 U23539 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20582), .ZN(n20638) );
  NOR2_X1 U23540 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20638), .ZN(
        n20591) );
  INV_X1 U23541 ( .A(n20591), .ZN(n20625) );
  OAI22_X1 U23542 ( .A1(n20668), .A2(n20725), .B1(n20583), .B2(n20625), .ZN(
        n20584) );
  INV_X1 U23543 ( .A(n20584), .ZN(n20593) );
  INV_X1 U23544 ( .A(n20585), .ZN(n20587) );
  AOI22_X1 U23545 ( .A1(n20588), .A2(n20587), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20586), .ZN(n20589) );
  AOI22_X1 U23546 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20629), .B1(
        n20628), .B2(n20722), .ZN(n20592) );
  OAI211_X1 U23547 ( .C1(n20633), .C2(n20594), .A(n20593), .B(n20592), .ZN(
        P1_U3129) );
  OAI22_X1 U23548 ( .A1(n20668), .A2(n20731), .B1(n20595), .B2(n20625), .ZN(
        n20596) );
  INV_X1 U23549 ( .A(n20596), .ZN(n20598) );
  AOI22_X1 U23550 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20629), .B1(
        n20628), .B2(n20728), .ZN(n20597) );
  OAI211_X1 U23551 ( .C1(n20633), .C2(n20599), .A(n20598), .B(n20597), .ZN(
        P1_U3130) );
  INV_X1 U23552 ( .A(n20733), .ZN(n20600) );
  OAI22_X1 U23553 ( .A1(n20668), .A2(n20687), .B1(n20600), .B2(n20625), .ZN(
        n20601) );
  INV_X1 U23554 ( .A(n20601), .ZN(n20603) );
  AOI22_X1 U23555 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20629), .B1(
        n20628), .B2(n20684), .ZN(n20602) );
  OAI211_X1 U23556 ( .C1(n20633), .C2(n20604), .A(n20603), .B(n20602), .ZN(
        P1_U3131) );
  OAI22_X1 U23557 ( .A1(n20668), .A2(n20691), .B1(n20605), .B2(n20625), .ZN(
        n20606) );
  INV_X1 U23558 ( .A(n20606), .ZN(n20608) );
  AOI22_X1 U23559 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20629), .B1(
        n20628), .B2(n20688), .ZN(n20607) );
  OAI211_X1 U23560 ( .C1(n20633), .C2(n20609), .A(n20608), .B(n20607), .ZN(
        P1_U3132) );
  INV_X1 U23561 ( .A(n20745), .ZN(n20610) );
  OAI22_X1 U23562 ( .A1(n20668), .A2(n20749), .B1(n20610), .B2(n20625), .ZN(
        n20611) );
  INV_X1 U23563 ( .A(n20611), .ZN(n20613) );
  AOI22_X1 U23564 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20629), .B1(
        n20628), .B2(n20746), .ZN(n20612) );
  OAI211_X1 U23565 ( .C1(n20633), .C2(n20614), .A(n20613), .B(n20612), .ZN(
        P1_U3133) );
  INV_X1 U23566 ( .A(n20751), .ZN(n20615) );
  OAI22_X1 U23567 ( .A1(n20668), .A2(n20697), .B1(n20615), .B2(n20625), .ZN(
        n20616) );
  INV_X1 U23568 ( .A(n20616), .ZN(n20618) );
  AOI22_X1 U23569 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20629), .B1(
        n20628), .B2(n20694), .ZN(n20617) );
  OAI211_X1 U23570 ( .C1(n20633), .C2(n20619), .A(n20618), .B(n20617), .ZN(
        P1_U3134) );
  OAI22_X1 U23571 ( .A1(n20668), .A2(n20701), .B1(n20620), .B2(n20625), .ZN(
        n20621) );
  INV_X1 U23572 ( .A(n20621), .ZN(n20623) );
  AOI22_X1 U23573 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20629), .B1(
        n20628), .B2(n20698), .ZN(n20622) );
  OAI211_X1 U23574 ( .C1(n20633), .C2(n20624), .A(n20623), .B(n20622), .ZN(
        P1_U3135) );
  OAI22_X1 U23575 ( .A1(n20668), .A2(n20774), .B1(n20626), .B2(n20625), .ZN(
        n20627) );
  INV_X1 U23576 ( .A(n20627), .ZN(n20631) );
  AOI22_X1 U23577 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20629), .B1(
        n20628), .B2(n20768), .ZN(n20630) );
  OAI211_X1 U23578 ( .C1(n20633), .C2(n20632), .A(n20631), .B(n20630), .ZN(
        P1_U3136) );
  NOR2_X1 U23579 ( .A1(n20634), .A2(n20638), .ZN(n20663) );
  INV_X1 U23580 ( .A(n20635), .ZN(n20710) );
  AOI21_X1 U23581 ( .B1(n20710), .B2(n20636), .A(n20663), .ZN(n20637) );
  OAI22_X1 U23582 ( .A1(n20637), .A2(n20719), .B1(n20638), .B2(n11773), .ZN(
        n20662) );
  AOI22_X1 U23583 ( .A1(n20713), .A2(n20663), .B1(n20712), .B2(n20662), .ZN(
        n20644) );
  INV_X1 U23584 ( .A(n20638), .ZN(n20640) );
  OAI21_X1 U23585 ( .B1(n20640), .B2(n20639), .A(n20717), .ZN(n20665) );
  NOR2_X2 U23586 ( .A1(n20716), .A2(n20641), .ZN(n20704) );
  AOI22_X1 U23587 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20665), .B1(
        n20704), .B2(n20642), .ZN(n20643) );
  OAI211_X1 U23588 ( .C1(n20645), .C2(n20668), .A(n20644), .B(n20643), .ZN(
        P1_U3137) );
  AOI22_X1 U23589 ( .A1(n20727), .A2(n20663), .B1(n20726), .B2(n20662), .ZN(
        n20648) );
  AOI22_X1 U23590 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20665), .B1(
        n20704), .B2(n20646), .ZN(n20647) );
  OAI211_X1 U23591 ( .C1(n20649), .C2(n20668), .A(n20648), .B(n20647), .ZN(
        P1_U3138) );
  AOI22_X1 U23592 ( .A1(n20733), .A2(n20663), .B1(n20732), .B2(n20662), .ZN(
        n20651) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20665), .B1(
        n20704), .B2(n20734), .ZN(n20650) );
  OAI211_X1 U23594 ( .C1(n20737), .C2(n20668), .A(n20651), .B(n20650), .ZN(
        P1_U3139) );
  AOI22_X1 U23595 ( .A1(n20739), .A2(n20663), .B1(n20738), .B2(n20662), .ZN(
        n20653) );
  AOI22_X1 U23596 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20665), .B1(
        n20704), .B2(n20740), .ZN(n20652) );
  OAI211_X1 U23597 ( .C1(n20743), .C2(n20668), .A(n20653), .B(n20652), .ZN(
        P1_U3140) );
  AOI22_X1 U23598 ( .A1(n20745), .A2(n20663), .B1(n20744), .B2(n20662), .ZN(
        n20656) );
  AOI22_X1 U23599 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20665), .B1(
        n20704), .B2(n20654), .ZN(n20655) );
  OAI211_X1 U23600 ( .C1(n20657), .C2(n20668), .A(n20656), .B(n20655), .ZN(
        P1_U3141) );
  AOI22_X1 U23601 ( .A1(n20751), .A2(n20663), .B1(n20750), .B2(n20662), .ZN(
        n20659) );
  AOI22_X1 U23602 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20665), .B1(
        n20704), .B2(n20752), .ZN(n20658) );
  OAI211_X1 U23603 ( .C1(n20755), .C2(n20668), .A(n20659), .B(n20658), .ZN(
        P1_U3142) );
  AOI22_X1 U23604 ( .A1(n20757), .A2(n20663), .B1(n20756), .B2(n20662), .ZN(
        n20661) );
  AOI22_X1 U23605 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20665), .B1(
        n20704), .B2(n20758), .ZN(n20660) );
  OAI211_X1 U23606 ( .C1(n20763), .C2(n20668), .A(n20661), .B(n20660), .ZN(
        P1_U3143) );
  AOI22_X1 U23607 ( .A1(n20767), .A2(n20663), .B1(n20764), .B2(n20662), .ZN(
        n20667) );
  AOI22_X1 U23608 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20665), .B1(
        n20704), .B2(n20664), .ZN(n20666) );
  OAI211_X1 U23609 ( .C1(n20669), .C2(n20668), .A(n20667), .B(n20666), .ZN(
        P1_U3144) );
  NOR2_X1 U23610 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20711), .ZN(
        n20703) );
  NAND3_X1 U23611 ( .A1(n20710), .A2(n20674), .A3(n20721), .ZN(n20671) );
  OAI21_X1 U23612 ( .B1(n20673), .B2(n20672), .A(n20671), .ZN(n20702) );
  AOI22_X1 U23613 ( .A1(n20713), .A2(n20703), .B1(n20712), .B2(n20702), .ZN(
        n20681) );
  OAI21_X1 U23614 ( .B1(n20704), .B2(n20769), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20676) );
  NAND2_X1 U23615 ( .A1(n20710), .A2(n20674), .ZN(n20675) );
  AOI21_X1 U23616 ( .B1(n20676), .B2(n20675), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20679) );
  AOI22_X1 U23617 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20705), .B1(
        n20704), .B2(n20722), .ZN(n20680) );
  OAI211_X1 U23618 ( .C1(n20725), .C2(n20762), .A(n20681), .B(n20680), .ZN(
        P1_U3145) );
  AOI22_X1 U23619 ( .A1(n20727), .A2(n20703), .B1(n20726), .B2(n20702), .ZN(
        n20683) );
  AOI22_X1 U23620 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20705), .B1(
        n20704), .B2(n20728), .ZN(n20682) );
  OAI211_X1 U23621 ( .C1(n20731), .C2(n20762), .A(n20683), .B(n20682), .ZN(
        P1_U3146) );
  AOI22_X1 U23622 ( .A1(n20733), .A2(n20703), .B1(n20732), .B2(n20702), .ZN(
        n20686) );
  AOI22_X1 U23623 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20705), .B1(
        n20704), .B2(n20684), .ZN(n20685) );
  OAI211_X1 U23624 ( .C1(n20687), .C2(n20762), .A(n20686), .B(n20685), .ZN(
        P1_U3147) );
  AOI22_X1 U23625 ( .A1(n20739), .A2(n20703), .B1(n20738), .B2(n20702), .ZN(
        n20690) );
  AOI22_X1 U23626 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20705), .B1(
        n20704), .B2(n20688), .ZN(n20689) );
  OAI211_X1 U23627 ( .C1(n20691), .C2(n20762), .A(n20690), .B(n20689), .ZN(
        P1_U3148) );
  AOI22_X1 U23628 ( .A1(n20745), .A2(n20703), .B1(n20744), .B2(n20702), .ZN(
        n20693) );
  AOI22_X1 U23629 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20705), .B1(
        n20704), .B2(n20746), .ZN(n20692) );
  OAI211_X1 U23630 ( .C1(n20749), .C2(n20762), .A(n20693), .B(n20692), .ZN(
        P1_U3149) );
  AOI22_X1 U23631 ( .A1(n20751), .A2(n20703), .B1(n20750), .B2(n20702), .ZN(
        n20696) );
  AOI22_X1 U23632 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20705), .B1(
        n20704), .B2(n20694), .ZN(n20695) );
  OAI211_X1 U23633 ( .C1(n20697), .C2(n20762), .A(n20696), .B(n20695), .ZN(
        P1_U3150) );
  AOI22_X1 U23634 ( .A1(n20757), .A2(n20703), .B1(n20756), .B2(n20702), .ZN(
        n20700) );
  AOI22_X1 U23635 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20705), .B1(
        n20704), .B2(n20698), .ZN(n20699) );
  OAI211_X1 U23636 ( .C1(n20701), .C2(n20762), .A(n20700), .B(n20699), .ZN(
        P1_U3151) );
  AOI22_X1 U23637 ( .A1(n20767), .A2(n20703), .B1(n20764), .B2(n20702), .ZN(
        n20707) );
  AOI22_X1 U23638 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20705), .B1(
        n20704), .B2(n20768), .ZN(n20706) );
  OAI211_X1 U23639 ( .C1(n20774), .C2(n20762), .A(n20707), .B(n20706), .ZN(
        P1_U3152) );
  INV_X1 U23640 ( .A(n20708), .ZN(n20766) );
  AOI21_X1 U23641 ( .B1(n20710), .B2(n20709), .A(n20766), .ZN(n20714) );
  OAI22_X1 U23642 ( .A1(n20714), .A2(n20719), .B1(n20711), .B2(n11773), .ZN(
        n20765) );
  AOI22_X1 U23643 ( .A1(n20713), .A2(n20766), .B1(n20765), .B2(n20712), .ZN(
        n20724) );
  OAI21_X1 U23644 ( .B1(n20716), .B2(n20715), .A(n20714), .ZN(n20718) );
  OAI221_X1 U23645 ( .B1(n20721), .B2(n20720), .C1(n20719), .C2(n20718), .A(
        n20717), .ZN(n20770) );
  AOI22_X1 U23646 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20770), .B1(
        n20769), .B2(n20722), .ZN(n20723) );
  OAI211_X1 U23647 ( .C1(n20725), .C2(n20773), .A(n20724), .B(n20723), .ZN(
        P1_U3153) );
  AOI22_X1 U23648 ( .A1(n20727), .A2(n20766), .B1(n20765), .B2(n20726), .ZN(
        n20730) );
  AOI22_X1 U23649 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20770), .B1(
        n20769), .B2(n20728), .ZN(n20729) );
  OAI211_X1 U23650 ( .C1(n20731), .C2(n20773), .A(n20730), .B(n20729), .ZN(
        P1_U3154) );
  AOI22_X1 U23651 ( .A1(n20733), .A2(n20766), .B1(n20765), .B2(n20732), .ZN(
        n20736) );
  AOI22_X1 U23652 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20770), .B1(
        n20759), .B2(n20734), .ZN(n20735) );
  OAI211_X1 U23653 ( .C1(n20737), .C2(n20762), .A(n20736), .B(n20735), .ZN(
        P1_U3155) );
  AOI22_X1 U23654 ( .A1(n20739), .A2(n20766), .B1(n20738), .B2(n20765), .ZN(
        n20742) );
  AOI22_X1 U23655 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20770), .B1(
        n20759), .B2(n20740), .ZN(n20741) );
  OAI211_X1 U23656 ( .C1(n20743), .C2(n20762), .A(n20742), .B(n20741), .ZN(
        P1_U3156) );
  AOI22_X1 U23657 ( .A1(n20745), .A2(n20766), .B1(n20765), .B2(n20744), .ZN(
        n20748) );
  AOI22_X1 U23658 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20770), .B1(
        n20769), .B2(n20746), .ZN(n20747) );
  OAI211_X1 U23659 ( .C1(n20749), .C2(n20773), .A(n20748), .B(n20747), .ZN(
        P1_U3157) );
  AOI22_X1 U23660 ( .A1(n20751), .A2(n20766), .B1(n20765), .B2(n20750), .ZN(
        n20754) );
  AOI22_X1 U23661 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20770), .B1(
        n20759), .B2(n20752), .ZN(n20753) );
  OAI211_X1 U23662 ( .C1(n20755), .C2(n20762), .A(n20754), .B(n20753), .ZN(
        P1_U3158) );
  AOI22_X1 U23663 ( .A1(n20757), .A2(n20766), .B1(n20756), .B2(n20765), .ZN(
        n20761) );
  AOI22_X1 U23664 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20770), .B1(
        n20759), .B2(n20758), .ZN(n20760) );
  OAI211_X1 U23665 ( .C1(n20763), .C2(n20762), .A(n20761), .B(n20760), .ZN(
        P1_U3159) );
  AOI22_X1 U23666 ( .A1(n20767), .A2(n20766), .B1(n20765), .B2(n20764), .ZN(
        n20772) );
  AOI22_X1 U23667 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20770), .B1(
        n20769), .B2(n20768), .ZN(n20771) );
  OAI211_X1 U23668 ( .C1(n20774), .C2(n20773), .A(n20772), .B(n20771), .ZN(
        P1_U3160) );
  OAI221_X1 U23669 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20777), .C1(n11773), 
        .C2(n20776), .A(n20775), .ZN(P1_U3163) );
  AND2_X1 U23670 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20850), .ZN(
        P1_U3164) );
  AND2_X1 U23671 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20850), .ZN(
        P1_U3165) );
  AND2_X1 U23672 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20850), .ZN(
        P1_U3166) );
  AND2_X1 U23673 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20850), .ZN(
        P1_U3167) );
  AND2_X1 U23674 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20850), .ZN(
        P1_U3168) );
  AND2_X1 U23675 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20850), .ZN(
        P1_U3169) );
  AND2_X1 U23676 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20850), .ZN(
        P1_U3170) );
  AND2_X1 U23677 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20850), .ZN(
        P1_U3171) );
  AND2_X1 U23678 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20850), .ZN(
        P1_U3172) );
  AND2_X1 U23679 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20850), .ZN(
        P1_U3173) );
  AND2_X1 U23680 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20850), .ZN(
        P1_U3174) );
  AND2_X1 U23681 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20850), .ZN(
        P1_U3175) );
  AND2_X1 U23682 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20850), .ZN(
        P1_U3176) );
  AND2_X1 U23683 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20850), .ZN(
        P1_U3177) );
  AND2_X1 U23684 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20850), .ZN(
        P1_U3178) );
  AND2_X1 U23685 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20850), .ZN(
        P1_U3179) );
  AND2_X1 U23686 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20850), .ZN(
        P1_U3180) );
  AND2_X1 U23687 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20850), .ZN(
        P1_U3181) );
  AND2_X1 U23688 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20850), .ZN(
        P1_U3182) );
  AND2_X1 U23689 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20850), .ZN(
        P1_U3183) );
  AND2_X1 U23690 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20850), .ZN(
        P1_U3184) );
  AND2_X1 U23691 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20850), .ZN(
        P1_U3185) );
  AND2_X1 U23692 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20850), .ZN(P1_U3186) );
  AND2_X1 U23693 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20850), .ZN(P1_U3187) );
  AND2_X1 U23694 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20850), .ZN(P1_U3188) );
  AND2_X1 U23695 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20850), .ZN(P1_U3189) );
  AND2_X1 U23696 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20850), .ZN(P1_U3190) );
  AND2_X1 U23697 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20850), .ZN(P1_U3191) );
  AND2_X1 U23698 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20850), .ZN(P1_U3192) );
  AND2_X1 U23699 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20850), .ZN(P1_U3193) );
  OAI21_X1 U23700 ( .B1(n20778), .B2(n20871), .A(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20784) );
  INV_X1 U23701 ( .A(n20784), .ZN(n20782) );
  NOR2_X1 U23702 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20779) );
  OAI22_X1 U23703 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20957), .B1(n20779), 
        .B2(n21032), .ZN(n20780) );
  NOR2_X1 U23704 ( .A1(n20967), .A2(n20780), .ZN(n20781) );
  OAI22_X1 U23705 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20782), .B1(n20885), 
        .B2(n20781), .ZN(P1_U3194) );
  OAI211_X1 U23706 ( .C1(NA), .C2(n20871), .A(P1_STATE_REG_1__SCAN_IN), .B(
        n11603), .ZN(n20783) );
  OAI211_X1 U23707 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20967), .A(
        P1_STATE_REG_0__SCAN_IN), .B(n20783), .ZN(n20788) );
  OAI211_X1 U23708 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20957), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20784), .ZN(n20787) );
  NOR2_X1 U23709 ( .A1(NA), .A2(n20871), .ZN(n20785) );
  NAND4_X1 U23710 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .A3(P1_REQUESTPENDING_REG_SCAN_IN), .A4(n20785), .ZN(n20786) );
  OAI211_X1 U23711 ( .C1(n21032), .C2(n20788), .A(n20787), .B(n20786), .ZN(
        P1_U3196) );
  NAND2_X1 U23712 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20885), .ZN(n20842) );
  INV_X1 U23713 ( .A(n20842), .ZN(n20818) );
  INV_X1 U23714 ( .A(n20818), .ZN(n20836) );
  NOR2_X1 U23715 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20883), .ZN(n20815) );
  AOI22_X1 U23716 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(n20883), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20815), .ZN(n20789) );
  OAI21_X1 U23717 ( .B1(n13342), .B2(n20836), .A(n20789), .ZN(P1_U3197) );
  AOI22_X1 U23718 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20883), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20818), .ZN(n20790) );
  OAI21_X1 U23719 ( .B1(n20792), .B2(n20838), .A(n20790), .ZN(P1_U3198) );
  OAI222_X1 U23720 ( .A1(n20836), .A2(n20792), .B1(n20791), .B2(n20840), .C1(
        n20793), .C2(n20838), .ZN(P1_U3199) );
  INV_X1 U23721 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20794) );
  OAI222_X1 U23722 ( .A1(n20838), .A2(n20796), .B1(n20794), .B2(n20840), .C1(
        n20793), .C2(n20836), .ZN(P1_U3200) );
  INV_X1 U23723 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20795) );
  OAI222_X1 U23724 ( .A1(n20842), .A2(n20796), .B1(n20795), .B2(n20840), .C1(
        n20798), .C2(n20838), .ZN(P1_U3201) );
  INV_X1 U23725 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20797) );
  OAI222_X1 U23726 ( .A1(n20842), .A2(n20798), .B1(n20797), .B2(n20840), .C1(
        n20800), .C2(n20838), .ZN(P1_U3202) );
  INV_X1 U23727 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20799) );
  OAI222_X1 U23728 ( .A1(n20836), .A2(n20800), .B1(n20799), .B2(n20840), .C1(
        n20802), .C2(n20838), .ZN(P1_U3203) );
  INV_X1 U23729 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20801) );
  OAI222_X1 U23730 ( .A1(n20836), .A2(n20802), .B1(n20801), .B2(n20840), .C1(
        n20804), .C2(n20838), .ZN(P1_U3204) );
  INV_X1 U23731 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20803) );
  OAI222_X1 U23732 ( .A1(n20842), .A2(n20804), .B1(n20803), .B2(n20840), .C1(
        n20806), .C2(n20838), .ZN(P1_U3205) );
  AOI22_X1 U23733 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n20883), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n20815), .ZN(n20805) );
  OAI21_X1 U23734 ( .B1(n20806), .B2(n20836), .A(n20805), .ZN(P1_U3206) );
  AOI22_X1 U23735 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20883), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n20818), .ZN(n20807) );
  OAI21_X1 U23736 ( .B1(n20809), .B2(n20838), .A(n20807), .ZN(P1_U3207) );
  INV_X1 U23737 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20808) );
  OAI222_X1 U23738 ( .A1(n20842), .A2(n20809), .B1(n20808), .B2(n20885), .C1(
        n20811), .C2(n20838), .ZN(P1_U3208) );
  AOI22_X1 U23739 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20883), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20815), .ZN(n20810) );
  OAI21_X1 U23740 ( .B1(n20811), .B2(n20836), .A(n20810), .ZN(P1_U3209) );
  AOI22_X1 U23741 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20883), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20818), .ZN(n20812) );
  OAI21_X1 U23742 ( .B1(n20814), .B2(n20838), .A(n20812), .ZN(P1_U3210) );
  INV_X1 U23743 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20813) );
  OAI222_X1 U23744 ( .A1(n20842), .A2(n20814), .B1(n20813), .B2(n20840), .C1(
        n20817), .C2(n20838), .ZN(P1_U3211) );
  AOI22_X1 U23745 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20883), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20815), .ZN(n20816) );
  OAI21_X1 U23746 ( .B1(n20817), .B2(n20836), .A(n20816), .ZN(P1_U3212) );
  AOI22_X1 U23747 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20883), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20818), .ZN(n20819) );
  OAI21_X1 U23748 ( .B1(n20821), .B2(n20838), .A(n20819), .ZN(P1_U3213) );
  INV_X1 U23749 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20820) );
  OAI222_X1 U23750 ( .A1(n20842), .A2(n20821), .B1(n20820), .B2(n20885), .C1(
        n20823), .C2(n20838), .ZN(P1_U3214) );
  INV_X1 U23751 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n20822) );
  OAI222_X1 U23752 ( .A1(n20842), .A2(n20823), .B1(n20822), .B2(n20840), .C1(
        n20824), .C2(n20838), .ZN(P1_U3215) );
  INV_X1 U23753 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20825) );
  OAI222_X1 U23754 ( .A1(n20838), .A2(n20985), .B1(n20825), .B2(n20885), .C1(
        n20824), .C2(n20836), .ZN(P1_U3216) );
  INV_X1 U23755 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20826) );
  OAI222_X1 U23756 ( .A1(n20842), .A2(n20985), .B1(n20826), .B2(n20885), .C1(
        n21023), .C2(n20838), .ZN(P1_U3217) );
  INV_X1 U23757 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20827) );
  INV_X1 U23758 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20829) );
  OAI222_X1 U23759 ( .A1(n20842), .A2(n21023), .B1(n20827), .B2(n20885), .C1(
        n20829), .C2(n20838), .ZN(P1_U3218) );
  INV_X1 U23760 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20828) );
  OAI222_X1 U23761 ( .A1(n20842), .A2(n20829), .B1(n20828), .B2(n20885), .C1(
        n21010), .C2(n20838), .ZN(P1_U3219) );
  INV_X1 U23762 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20830) );
  OAI222_X1 U23763 ( .A1(n20838), .A2(n21011), .B1(n20830), .B2(n20885), .C1(
        n21010), .C2(n20836), .ZN(P1_U3220) );
  INV_X1 U23764 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20831) );
  OAI222_X1 U23765 ( .A1(n20838), .A2(n21013), .B1(n20831), .B2(n20885), .C1(
        n21011), .C2(n20836), .ZN(P1_U3221) );
  INV_X1 U23766 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20832) );
  OAI222_X1 U23767 ( .A1(n20838), .A2(n20948), .B1(n20832), .B2(n20885), .C1(
        n21013), .C2(n20836), .ZN(P1_U3222) );
  INV_X1 U23768 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20833) );
  OAI222_X1 U23769 ( .A1(n20836), .A2(n20948), .B1(n20833), .B2(n20885), .C1(
        n20835), .C2(n20838), .ZN(P1_U3223) );
  INV_X1 U23770 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20834) );
  OAI222_X1 U23771 ( .A1(n20836), .A2(n20835), .B1(n20834), .B2(n20885), .C1(
        n20963), .C2(n20838), .ZN(P1_U3224) );
  INV_X1 U23772 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n20837) );
  OAI222_X1 U23773 ( .A1(n20842), .A2(n20963), .B1(n20837), .B2(n20885), .C1(
        n21017), .C2(n20838), .ZN(P1_U3225) );
  INV_X1 U23774 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20841) );
  OAI222_X1 U23775 ( .A1(n20842), .A2(n21017), .B1(n20841), .B2(n20840), .C1(
        n20839), .C2(n20838), .ZN(P1_U3226) );
  INV_X1 U23776 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20843) );
  AOI22_X1 U23777 ( .A1(n20885), .A2(n20844), .B1(n20843), .B2(n20883), .ZN(
        P1_U3458) );
  INV_X1 U23778 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20864) );
  INV_X1 U23779 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20845) );
  AOI22_X1 U23780 ( .A1(n20885), .A2(n20864), .B1(n20845), .B2(n20883), .ZN(
        P1_U3459) );
  INV_X1 U23781 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20846) );
  AOI22_X1 U23782 ( .A1(n20885), .A2(n20847), .B1(n20846), .B2(n20883), .ZN(
        P1_U3460) );
  INV_X1 U23783 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21016) );
  INV_X1 U23784 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20848) );
  AOI22_X1 U23785 ( .A1(n20885), .A2(n21016), .B1(n20848), .B2(n20883), .ZN(
        P1_U3461) );
  INV_X1 U23786 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20851) );
  INV_X1 U23787 ( .A(n20852), .ZN(n20849) );
  AOI21_X1 U23788 ( .B1(n20851), .B2(n20850), .A(n20849), .ZN(P1_U3464) );
  OAI21_X1 U23789 ( .B1(n20854), .B2(n20853), .A(n20852), .ZN(P1_U3465) );
  AOI22_X1 U23790 ( .A1(n20858), .A2(n20857), .B1(n20856), .B2(n20855), .ZN(
        n20859) );
  INV_X1 U23791 ( .A(n20859), .ZN(n20861) );
  MUX2_X1 U23792 ( .A(n20861), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n20860), .Z(P1_U3469) );
  AOI21_X1 U23793 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20862) );
  AOI22_X1 U23794 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20862), .B2(n13342), .ZN(n20865) );
  AOI22_X1 U23795 ( .A1(n20867), .A2(n20865), .B1(n20864), .B2(n20863), .ZN(
        P1_U3481) );
  OAI21_X1 U23796 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20867), .ZN(n20866) );
  OAI21_X1 U23797 ( .B1(n20867), .B2(n21016), .A(n20866), .ZN(P1_U3482) );
  INV_X1 U23798 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20868) );
  AOI22_X1 U23799 ( .A1(n20885), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20868), 
        .B2(n20883), .ZN(P1_U3483) );
  AOI211_X1 U23800 ( .C1(n20872), .C2(n20871), .A(n20870), .B(n20869), .ZN(
        n20882) );
  OAI21_X1 U23801 ( .B1(n20875), .B2(n20874), .A(n20873), .ZN(n20876) );
  NAND3_X1 U23802 ( .A1(n20877), .A2(n20876), .A3(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n20878) );
  NAND2_X1 U23803 ( .A1(n20878), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20881) );
  NOR2_X1 U23804 ( .A1(n20882), .A2(n20879), .ZN(n20880) );
  AOI22_X1 U23805 ( .A1(n20967), .A2(n20882), .B1(n20881), .B2(n20880), .ZN(
        P1_U3485) );
  INV_X1 U23806 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n20884) );
  AOI22_X1 U23807 ( .A1(n20885), .A2(n20884), .B1(n21002), .B2(n20883), .ZN(
        P1_U3486) );
  INV_X1 U23808 ( .A(DATAI_6_), .ZN(n21081) );
  AOI22_X1 U23809 ( .A1(P1_READREQUEST_REG_SCAN_IN), .A2(keyinput_f38), .B1(
        DATAI_31_), .B2(keyinput_f1), .ZN(n20886) );
  OAI221_X1 U23810 ( .B1(P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_f38), .C1(
        DATAI_31_), .C2(keyinput_f1), .A(n20886), .ZN(n20945) );
  AOI22_X1 U23811 ( .A1(READY1), .A2(keyinput_f36), .B1(
        P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_f44), .ZN(n20887) );
  OAI221_X1 U23812 ( .B1(READY1), .B2(keyinput_f36), .C1(
        P1_STATEBS16_REG_SCAN_IN), .C2(keyinput_f44), .A(n20887), .ZN(n20944)
         );
  AOI22_X1 U23813 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_f0), .B1(
        n21026), .B2(keyinput_f16), .ZN(n20888) );
  OAI221_X1 U23814 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_f0), .C1(
        n21026), .C2(keyinput_f16), .A(n20888), .ZN(n20898) );
  OAI22_X1 U23815 ( .A1(DATAI_7_), .A2(keyinput_f25), .B1(
        P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_f51), .ZN(n20889) );
  AOI221_X1 U23816 ( .B1(DATAI_7_), .B2(keyinput_f25), .C1(keyinput_f51), .C2(
        P1_BYTEENABLE_REG_3__SCAN_IN), .A(n20889), .ZN(n20896) );
  OAI22_X1 U23817 ( .A1(DATAI_26_), .A2(keyinput_f6), .B1(keyinput_f39), .B2(
        P1_ADS_N_REG_SCAN_IN), .ZN(n20890) );
  AOI221_X1 U23818 ( .B1(DATAI_26_), .B2(keyinput_f6), .C1(
        P1_ADS_N_REG_SCAN_IN), .C2(keyinput_f39), .A(n20890), .ZN(n20895) );
  OAI22_X1 U23819 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(keyinput_f63), .B1(
        keyinput_f13), .B2(DATAI_19_), .ZN(n20891) );
  AOI221_X1 U23820 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(keyinput_f63), .C1(
        DATAI_19_), .C2(keyinput_f13), .A(n20891), .ZN(n20894) );
  OAI22_X1 U23821 ( .A1(DATAI_8_), .A2(keyinput_f24), .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_f46), .ZN(n20892) );
  AOI221_X1 U23822 ( .B1(DATAI_8_), .B2(keyinput_f24), .C1(keyinput_f46), .C2(
        P1_FLUSH_REG_SCAN_IN), .A(n20892), .ZN(n20893) );
  NAND4_X1 U23823 ( .A1(n20896), .A2(n20895), .A3(n20894), .A4(n20893), .ZN(
        n20897) );
  AOI211_X1 U23824 ( .C1(keyinput_f18), .C2(DATAI_14_), .A(n20898), .B(n20897), 
        .ZN(n20899) );
  OAI21_X1 U23825 ( .B1(keyinput_f18), .B2(DATAI_14_), .A(n20899), .ZN(n20943)
         );
  AOI22_X1 U23826 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(keyinput_f55), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(keyinput_f60), .ZN(n20900) );
  OAI221_X1 U23827 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(keyinput_f55), .C1(
        P1_REIP_REG_23__SCAN_IN), .C2(keyinput_f60), .A(n20900), .ZN(n20907)
         );
  AOI22_X1 U23828 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(keyinput_f40), .B1(
        DATAI_20_), .B2(keyinput_f12), .ZN(n20901) );
  OAI221_X1 U23829 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_f40), .C1(
        DATAI_20_), .C2(keyinput_f12), .A(n20901), .ZN(n20906) );
  AOI22_X1 U23830 ( .A1(DATAI_5_), .A2(keyinput_f27), .B1(DATAI_23_), .B2(
        keyinput_f9), .ZN(n20902) );
  OAI221_X1 U23831 ( .B1(DATAI_5_), .B2(keyinput_f27), .C1(DATAI_23_), .C2(
        keyinput_f9), .A(n20902), .ZN(n20905) );
  AOI22_X1 U23832 ( .A1(keyinput_f49), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        DATAI_2_), .B2(keyinput_f30), .ZN(n20903) );
  OAI221_X1 U23833 ( .B1(keyinput_f49), .B2(P1_BYTEENABLE_REG_1__SCAN_IN), 
        .C1(DATAI_2_), .C2(keyinput_f30), .A(n20903), .ZN(n20904) );
  NOR4_X1 U23834 ( .A1(n20907), .A2(n20906), .A3(n20905), .A4(n20904), .ZN(
        n20941) );
  AOI22_X1 U23835 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(keyinput_f57), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(keyinput_f53), .ZN(n20908) );
  OAI221_X1 U23836 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_f57), .C1(
        P1_REIP_REG_30__SCAN_IN), .C2(keyinput_f53), .A(n20908), .ZN(n20915)
         );
  AOI22_X1 U23837 ( .A1(DATAI_28_), .A2(keyinput_f4), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(keyinput_f58), .ZN(n20909) );
  OAI221_X1 U23838 ( .B1(DATAI_28_), .B2(keyinput_f4), .C1(
        P1_REIP_REG_25__SCAN_IN), .C2(keyinput_f58), .A(n20909), .ZN(n20914)
         );
  AOI22_X1 U23839 ( .A1(DATAI_17_), .A2(keyinput_f15), .B1(DATAI_10_), .B2(
        keyinput_f22), .ZN(n20910) );
  OAI221_X1 U23840 ( .B1(DATAI_17_), .B2(keyinput_f15), .C1(DATAI_10_), .C2(
        keyinput_f22), .A(n20910), .ZN(n20913) );
  AOI22_X1 U23841 ( .A1(DATAI_0_), .A2(keyinput_f32), .B1(DATAI_29_), .B2(
        keyinput_f3), .ZN(n20911) );
  OAI221_X1 U23842 ( .B1(DATAI_0_), .B2(keyinput_f32), .C1(DATAI_29_), .C2(
        keyinput_f3), .A(n20911), .ZN(n20912) );
  NOR4_X1 U23843 ( .A1(n20915), .A2(n20914), .A3(n20913), .A4(n20912), .ZN(
        n20940) );
  AOI22_X1 U23844 ( .A1(n14549), .A2(keyinput_f17), .B1(keyinput_f33), .B2(
        n21032), .ZN(n20916) );
  OAI221_X1 U23845 ( .B1(n14549), .B2(keyinput_f17), .C1(n21032), .C2(
        keyinput_f33), .A(n20916), .ZN(n20927) );
  INV_X1 U23846 ( .A(keyinput_f47), .ZN(n20918) );
  AOI22_X1 U23847 ( .A1(n20919), .A2(keyinput_f45), .B1(P1_W_R_N_REG_SCAN_IN), 
        .B2(n20918), .ZN(n20917) );
  OAI221_X1 U23848 ( .B1(n20919), .B2(keyinput_f45), .C1(n20918), .C2(
        P1_W_R_N_REG_SCAN_IN), .A(n20917), .ZN(n20926) );
  AOI22_X1 U23849 ( .A1(n21023), .A2(keyinput_f61), .B1(keyinput_f35), .B2(
        n21030), .ZN(n20920) );
  OAI221_X1 U23850 ( .B1(n21023), .B2(keyinput_f61), .C1(n21030), .C2(
        keyinput_f35), .A(n20920), .ZN(n20925) );
  AOI22_X1 U23851 ( .A1(n20923), .A2(keyinput_f28), .B1(n20922), .B2(
        keyinput_f5), .ZN(n20921) );
  OAI221_X1 U23852 ( .B1(n20923), .B2(keyinput_f28), .C1(n20922), .C2(
        keyinput_f5), .A(n20921), .ZN(n20924) );
  NOR4_X1 U23853 ( .A1(n20927), .A2(n20926), .A3(n20925), .A4(n20924), .ZN(
        n20939) );
  AOI22_X1 U23854 ( .A1(DATAI_25_), .A2(keyinput_f7), .B1(DATAI_30_), .B2(
        keyinput_f2), .ZN(n20928) );
  OAI221_X1 U23855 ( .B1(DATAI_25_), .B2(keyinput_f7), .C1(DATAI_30_), .C2(
        keyinput_f2), .A(n20928), .ZN(n20937) );
  AOI22_X1 U23856 ( .A1(DATAI_21_), .A2(keyinput_f11), .B1(
        P1_REIP_REG_31__SCAN_IN), .B2(keyinput_f52), .ZN(n20929) );
  OAI221_X1 U23857 ( .B1(DATAI_21_), .B2(keyinput_f11), .C1(
        P1_REIP_REG_31__SCAN_IN), .C2(keyinput_f52), .A(n20929), .ZN(n20936)
         );
  INV_X1 U23858 ( .A(DATAI_3_), .ZN(n20987) );
  AOI22_X1 U23859 ( .A1(n20987), .A2(keyinput_f29), .B1(keyinput_f42), .B2(
        n20991), .ZN(n20930) );
  OAI221_X1 U23860 ( .B1(n20987), .B2(keyinput_f29), .C1(n20991), .C2(
        keyinput_f42), .A(n20930), .ZN(n20935) );
  INV_X1 U23861 ( .A(keyinput_f50), .ZN(n20932) );
  AOI22_X1 U23862 ( .A1(n20933), .A2(keyinput_f8), .B1(
        P1_BYTEENABLE_REG_2__SCAN_IN), .B2(n20932), .ZN(n20931) );
  OAI221_X1 U23863 ( .B1(n20933), .B2(keyinput_f8), .C1(n20932), .C2(
        P1_BYTEENABLE_REG_2__SCAN_IN), .A(n20931), .ZN(n20934) );
  NOR4_X1 U23864 ( .A1(n20937), .A2(n20936), .A3(n20935), .A4(n20934), .ZN(
        n20938) );
  NAND4_X1 U23865 ( .A1(n20941), .A2(n20940), .A3(n20939), .A4(n20938), .ZN(
        n20942) );
  NOR4_X1 U23866 ( .A1(n20945), .A2(n20944), .A3(n20943), .A4(n20942), .ZN(
        n20979) );
  AOI22_X1 U23867 ( .A1(n20948), .A2(keyinput_f56), .B1(keyinput_f21), .B2(
        n20947), .ZN(n20946) );
  OAI221_X1 U23868 ( .B1(n20948), .B2(keyinput_f56), .C1(n20947), .C2(
        keyinput_f21), .A(n20946), .ZN(n20976) );
  AOI22_X1 U23869 ( .A1(n20950), .A2(keyinput_f31), .B1(n21010), .B2(
        keyinput_f59), .ZN(n20949) );
  OAI221_X1 U23870 ( .B1(n20950), .B2(keyinput_f31), .C1(n21010), .C2(
        keyinput_f59), .A(n20949), .ZN(n20975) );
  OAI22_X1 U23871 ( .A1(n20953), .A2(keyinput_f19), .B1(n20952), .B2(
        keyinput_f10), .ZN(n20951) );
  AOI221_X1 U23872 ( .B1(n20953), .B2(keyinput_f19), .C1(keyinput_f10), .C2(
        n20952), .A(n20951), .ZN(n20956) );
  XOR2_X1 U23873 ( .A(keyinput_f41), .B(P1_M_IO_N_REG_SCAN_IN), .Z(n20954) );
  AOI21_X1 U23874 ( .B1(keyinput_f34), .B2(n20957), .A(n20954), .ZN(n20955) );
  OAI211_X1 U23875 ( .C1(keyinput_f34), .C2(n20957), .A(n20956), .B(n20955), 
        .ZN(n20974) );
  INV_X1 U23876 ( .A(DATAI_12_), .ZN(n20960) );
  OAI22_X1 U23877 ( .A1(n20960), .A2(keyinput_f20), .B1(n20959), .B2(
        keyinput_f14), .ZN(n20958) );
  AOI221_X1 U23878 ( .B1(n20960), .B2(keyinput_f20), .C1(keyinput_f14), .C2(
        n20959), .A(n20958), .ZN(n20972) );
  INV_X1 U23879 ( .A(READY2), .ZN(n20962) );
  OAI22_X1 U23880 ( .A1(n20963), .A2(keyinput_f54), .B1(n20962), .B2(
        keyinput_f37), .ZN(n20961) );
  AOI221_X1 U23881 ( .B1(n20963), .B2(keyinput_f54), .C1(keyinput_f37), .C2(
        n20962), .A(n20961), .ZN(n20971) );
  INV_X1 U23882 ( .A(keyinput_f48), .ZN(n20965) );
  OAI22_X1 U23883 ( .A1(n20985), .A2(keyinput_f62), .B1(n20965), .B2(
        P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20964) );
  AOI221_X1 U23884 ( .B1(n20985), .B2(keyinput_f62), .C1(
        P1_BYTEENABLE_REG_0__SCAN_IN), .C2(n20965), .A(n20964), .ZN(n20970) );
  OAI22_X1 U23885 ( .A1(n20968), .A2(keyinput_f23), .B1(n20967), .B2(
        keyinput_f43), .ZN(n20966) );
  AOI221_X1 U23886 ( .B1(n20968), .B2(keyinput_f23), .C1(keyinput_f43), .C2(
        n20967), .A(n20966), .ZN(n20969) );
  NAND4_X1 U23887 ( .A1(n20972), .A2(n20971), .A3(n20970), .A4(n20969), .ZN(
        n20973) );
  NOR4_X1 U23888 ( .A1(n20976), .A2(n20975), .A3(n20974), .A4(n20973), .ZN(
        n20978) );
  NOR2_X1 U23889 ( .A1(n21081), .A2(keyinput_f26), .ZN(n20977) );
  AOI221_X1 U23890 ( .B1(n20979), .B2(n20978), .C1(keyinput_f26), .C2(n21081), 
        .A(n20977), .ZN(n21080) );
  AOI22_X1 U23891 ( .A1(n20982), .A2(keyinput_g39), .B1(n20981), .B2(
        keyinput_g4), .ZN(n20980) );
  OAI221_X1 U23892 ( .B1(n20982), .B2(keyinput_g39), .C1(n20981), .C2(
        keyinput_g4), .A(n20980), .ZN(n20995) );
  AOI22_X1 U23893 ( .A1(n20985), .A2(keyinput_g62), .B1(keyinput_g40), .B2(
        n20984), .ZN(n20983) );
  OAI221_X1 U23894 ( .B1(n20985), .B2(keyinput_g62), .C1(n20984), .C2(
        keyinput_g40), .A(n20983), .ZN(n20994) );
  AOI22_X1 U23895 ( .A1(n20988), .A2(keyinput_g13), .B1(n20987), .B2(
        keyinput_g29), .ZN(n20986) );
  OAI221_X1 U23896 ( .B1(n20988), .B2(keyinput_g13), .C1(n20987), .C2(
        keyinput_g29), .A(n20986), .ZN(n20993) );
  AOI22_X1 U23897 ( .A1(n20991), .A2(keyinput_g42), .B1(n20990), .B2(
        keyinput_g15), .ZN(n20989) );
  OAI221_X1 U23898 ( .B1(n20991), .B2(keyinput_g42), .C1(n20990), .C2(
        keyinput_g15), .A(n20989), .ZN(n20992) );
  NOR4_X1 U23899 ( .A1(n20995), .A2(n20994), .A3(n20993), .A4(n20992), .ZN(
        n21041) );
  AOI22_X1 U23900 ( .A1(READY2), .A2(keyinput_g37), .B1(DATAI_29_), .B2(
        keyinput_g3), .ZN(n20996) );
  OAI221_X1 U23901 ( .B1(READY2), .B2(keyinput_g37), .C1(DATAI_29_), .C2(
        keyinput_g3), .A(n20996), .ZN(n21006) );
  AOI22_X1 U23902 ( .A1(DATAI_7_), .A2(keyinput_g25), .B1(
        P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_g44), .ZN(n20997) );
  OAI221_X1 U23903 ( .B1(DATAI_7_), .B2(keyinput_g25), .C1(
        P1_STATEBS16_REG_SCAN_IN), .C2(keyinput_g44), .A(n20997), .ZN(n21005)
         );
  INV_X1 U23904 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n20999) );
  AOI22_X1 U23905 ( .A1(n21000), .A2(keyinput_g1), .B1(keyinput_g38), .B2(
        n20999), .ZN(n20998) );
  OAI221_X1 U23906 ( .B1(n21000), .B2(keyinput_g1), .C1(n20999), .C2(
        keyinput_g38), .A(n20998), .ZN(n21004) );
  AOI22_X1 U23907 ( .A1(P1_BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_g49), .B1(
        n21002), .B2(keyinput_g41), .ZN(n21001) );
  OAI221_X1 U23908 ( .B1(P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_g49), 
        .C1(n21002), .C2(keyinput_g41), .A(n21001), .ZN(n21003) );
  NOR4_X1 U23909 ( .A1(n21006), .A2(n21005), .A3(n21004), .A4(n21003), .ZN(
        n21040) );
  INV_X1 U23910 ( .A(READY1), .ZN(n21008) );
  AOI22_X1 U23911 ( .A1(n14549), .A2(keyinput_g17), .B1(n21008), .B2(
        keyinput_g36), .ZN(n21007) );
  OAI221_X1 U23912 ( .B1(n14549), .B2(keyinput_g17), .C1(n21008), .C2(
        keyinput_g36), .A(n21007), .ZN(n21021) );
  AOI22_X1 U23913 ( .A1(n21011), .A2(keyinput_g58), .B1(n21010), .B2(
        keyinput_g59), .ZN(n21009) );
  OAI221_X1 U23914 ( .B1(n21011), .B2(keyinput_g58), .C1(n21010), .C2(
        keyinput_g59), .A(n21009), .ZN(n21020) );
  AOI22_X1 U23915 ( .A1(n21014), .A2(keyinput_g6), .B1(n21013), .B2(
        keyinput_g57), .ZN(n21012) );
  OAI221_X1 U23916 ( .B1(n21014), .B2(keyinput_g6), .C1(n21013), .C2(
        keyinput_g57), .A(n21012), .ZN(n21019) );
  AOI22_X1 U23917 ( .A1(n21017), .A2(keyinput_g53), .B1(keyinput_g48), .B2(
        n21016), .ZN(n21015) );
  OAI221_X1 U23918 ( .B1(n21017), .B2(keyinput_g53), .C1(n21016), .C2(
        keyinput_g48), .A(n21015), .ZN(n21018) );
  NOR4_X1 U23919 ( .A1(n21021), .A2(n21020), .A3(n21019), .A4(n21018), .ZN(
        n21039) );
  AOI22_X1 U23920 ( .A1(n21024), .A2(keyinput_g18), .B1(n21023), .B2(
        keyinput_g61), .ZN(n21022) );
  OAI221_X1 U23921 ( .B1(n21024), .B2(keyinput_g18), .C1(n21023), .C2(
        keyinput_g61), .A(n21022), .ZN(n21037) );
  AOI22_X1 U23922 ( .A1(n21027), .A2(keyinput_g2), .B1(keyinput_g16), .B2(
        n21026), .ZN(n21025) );
  OAI221_X1 U23923 ( .B1(n21027), .B2(keyinput_g2), .C1(n21026), .C2(
        keyinput_g16), .A(n21025), .ZN(n21036) );
  INV_X1 U23924 ( .A(DATAI_2_), .ZN(n21029) );
  AOI22_X1 U23925 ( .A1(n21030), .A2(keyinput_g35), .B1(n21029), .B2(
        keyinput_g30), .ZN(n21028) );
  OAI221_X1 U23926 ( .B1(n21030), .B2(keyinput_g35), .C1(n21029), .C2(
        keyinput_g30), .A(n21028), .ZN(n21035) );
  AOI22_X1 U23927 ( .A1(n21033), .A2(keyinput_g7), .B1(keyinput_g33), .B2(
        n21032), .ZN(n21031) );
  OAI221_X1 U23928 ( .B1(n21033), .B2(keyinput_g7), .C1(n21032), .C2(
        keyinput_g33), .A(n21031), .ZN(n21034) );
  NOR4_X1 U23929 ( .A1(n21037), .A2(n21036), .A3(n21035), .A4(n21034), .ZN(
        n21038) );
  NAND4_X1 U23930 ( .A1(n21041), .A2(n21040), .A3(n21039), .A4(n21038), .ZN(
        n21078) );
  AOI22_X1 U23931 ( .A1(DATAI_10_), .A2(keyinput_g22), .B1(
        P1_REIP_REG_27__SCAN_IN), .B2(keyinput_g56), .ZN(n21042) );
  OAI221_X1 U23932 ( .B1(DATAI_10_), .B2(keyinput_g22), .C1(
        P1_REIP_REG_27__SCAN_IN), .C2(keyinput_g56), .A(n21042), .ZN(n21049)
         );
  AOI22_X1 U23933 ( .A1(DATAI_0_), .A2(keyinput_g32), .B1(DATAI_18_), .B2(
        keyinput_g14), .ZN(n21043) );
  OAI221_X1 U23934 ( .B1(DATAI_0_), .B2(keyinput_g32), .C1(DATAI_18_), .C2(
        keyinput_g14), .A(n21043), .ZN(n21048) );
  AOI22_X1 U23935 ( .A1(DATAI_20_), .A2(keyinput_g12), .B1(DATAI_5_), .B2(
        keyinput_g27), .ZN(n21044) );
  OAI221_X1 U23936 ( .B1(DATAI_20_), .B2(keyinput_g12), .C1(DATAI_5_), .C2(
        keyinput_g27), .A(n21044), .ZN(n21047) );
  AOI22_X1 U23937 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(keyinput_g55), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(keyinput_g63), .ZN(n21045) );
  OAI221_X1 U23938 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(keyinput_g55), .C1(
        P1_REIP_REG_20__SCAN_IN), .C2(keyinput_g63), .A(n21045), .ZN(n21046)
         );
  NOR4_X1 U23939 ( .A1(n21049), .A2(n21048), .A3(n21047), .A4(n21046), .ZN(
        n21076) );
  XOR2_X1 U23940 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(keyinput_g51), .Z(
        n21056) );
  AOI22_X1 U23941 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_g0), .B1(
        DATAI_9_), .B2(keyinput_g23), .ZN(n21050) );
  OAI221_X1 U23942 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_g0), .C1(
        DATAI_9_), .C2(keyinput_g23), .A(n21050), .ZN(n21055) );
  AOI22_X1 U23943 ( .A1(NA), .A2(keyinput_g34), .B1(P1_FLUSH_REG_SCAN_IN), 
        .B2(keyinput_g46), .ZN(n21051) );
  OAI221_X1 U23944 ( .B1(NA), .B2(keyinput_g34), .C1(P1_FLUSH_REG_SCAN_IN), 
        .C2(keyinput_g46), .A(n21051), .ZN(n21054) );
  AOI22_X1 U23945 ( .A1(DATAI_13_), .A2(keyinput_g19), .B1(
        P1_REIP_REG_31__SCAN_IN), .B2(keyinput_g52), .ZN(n21052) );
  OAI221_X1 U23946 ( .B1(DATAI_13_), .B2(keyinput_g19), .C1(
        P1_REIP_REG_31__SCAN_IN), .C2(keyinput_g52), .A(n21052), .ZN(n21053)
         );
  NOR4_X1 U23947 ( .A1(n21056), .A2(n21055), .A3(n21054), .A4(n21053), .ZN(
        n21075) );
  AOI22_X1 U23948 ( .A1(P1_W_R_N_REG_SCAN_IN), .A2(keyinput_g47), .B1(
        DATAI_27_), .B2(keyinput_g5), .ZN(n21057) );
  OAI221_X1 U23949 ( .B1(P1_W_R_N_REG_SCAN_IN), .B2(keyinput_g47), .C1(
        DATAI_27_), .C2(keyinput_g5), .A(n21057), .ZN(n21064) );
  AOI22_X1 U23950 ( .A1(DATAI_8_), .A2(keyinput_g24), .B1(DATAI_12_), .B2(
        keyinput_g20), .ZN(n21058) );
  OAI221_X1 U23951 ( .B1(DATAI_8_), .B2(keyinput_g24), .C1(DATAI_12_), .C2(
        keyinput_g20), .A(n21058), .ZN(n21063) );
  AOI22_X1 U23952 ( .A1(P1_BYTEENABLE_REG_2__SCAN_IN), .A2(keyinput_g50), .B1(
        DATAI_1_), .B2(keyinput_g31), .ZN(n21059) );
  OAI221_X1 U23953 ( .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_g50), 
        .C1(DATAI_1_), .C2(keyinput_g31), .A(n21059), .ZN(n21062) );
  AOI22_X1 U23954 ( .A1(P1_REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_g43), 
        .B1(P1_MORE_REG_SCAN_IN), .B2(keyinput_g45), .ZN(n21060) );
  OAI221_X1 U23955 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_g43), 
        .C1(P1_MORE_REG_SCAN_IN), .C2(keyinput_g45), .A(n21060), .ZN(n21061)
         );
  NOR4_X1 U23956 ( .A1(n21064), .A2(n21063), .A3(n21062), .A4(n21061), .ZN(
        n21074) );
  AOI22_X1 U23957 ( .A1(DATAI_21_), .A2(keyinput_g11), .B1(DATAI_22_), .B2(
        keyinput_g10), .ZN(n21065) );
  OAI221_X1 U23958 ( .B1(DATAI_21_), .B2(keyinput_g11), .C1(DATAI_22_), .C2(
        keyinput_g10), .A(n21065), .ZN(n21072) );
  AOI22_X1 U23959 ( .A1(DATAI_24_), .A2(keyinput_g8), .B1(DATAI_11_), .B2(
        keyinput_g21), .ZN(n21066) );
  OAI221_X1 U23960 ( .B1(DATAI_24_), .B2(keyinput_g8), .C1(DATAI_11_), .C2(
        keyinput_g21), .A(n21066), .ZN(n21071) );
  AOI22_X1 U23961 ( .A1(DATAI_23_), .A2(keyinput_g9), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(keyinput_g60), .ZN(n21067) );
  OAI221_X1 U23962 ( .B1(DATAI_23_), .B2(keyinput_g9), .C1(
        P1_REIP_REG_23__SCAN_IN), .C2(keyinput_g60), .A(n21067), .ZN(n21070)
         );
  AOI22_X1 U23963 ( .A1(DATAI_4_), .A2(keyinput_g28), .B1(
        P1_REIP_REG_29__SCAN_IN), .B2(keyinput_g54), .ZN(n21068) );
  OAI221_X1 U23964 ( .B1(DATAI_4_), .B2(keyinput_g28), .C1(
        P1_REIP_REG_29__SCAN_IN), .C2(keyinput_g54), .A(n21068), .ZN(n21069)
         );
  NOR4_X1 U23965 ( .A1(n21072), .A2(n21071), .A3(n21070), .A4(n21069), .ZN(
        n21073) );
  NAND4_X1 U23966 ( .A1(n21076), .A2(n21075), .A3(n21074), .A4(n21073), .ZN(
        n21077) );
  OAI22_X1 U23967 ( .A1(keyinput_g26), .A2(n21081), .B1(n21078), .B2(n21077), 
        .ZN(n21079) );
  AOI211_X1 U23968 ( .C1(keyinput_g26), .C2(n21081), .A(n21080), .B(n21079), 
        .ZN(n21083) );
  AOI22_X1 U23969 ( .A1(n16499), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n16501), .ZN(n21082) );
  XNOR2_X1 U23970 ( .A(n21083), .B(n21082), .ZN(U355) );
  INV_X1 U11111 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10510) );
  INV_X2 U11088 ( .A(n10770), .ZN(n19251) );
  AND2_X2 U11576 ( .A1(n9650), .A2(n10510), .ZN(n10727) );
  AND2_X2 U11131 ( .A1(n14181), .A2(n10639), .ZN(n13047) );
  CLKBUF_X1 U11158 ( .A(n12442), .Z(n9638) );
  INV_X1 U11206 ( .A(n11576), .ZN(n11622) );
  CLKBUF_X1 U11219 ( .A(n10558), .Z(n10573) );
  INV_X2 U11367 ( .A(n17155), .ZN(n17049) );
  NAND2_X1 U11454 ( .A1(n10523), .A2(n10522), .ZN(n10556) );
  AND2_X2 U12326 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10183) );
  CLKBUF_X1 U12423 ( .A(n10556), .Z(n19262) );
  CLKBUF_X1 U12424 ( .A(n19154), .Z(n19170) );
  CLKBUF_X1 U12813 ( .A(n18840), .Z(n18833) );
  CLKBUF_X1 U13245 ( .A(n16481), .Z(n16495) );
endmodule

