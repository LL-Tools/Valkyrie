

module b14_C_AntiSAT_k_256_1 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2218, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083;

  AND2_X1 U2460 ( .A1(n3176), .A2(n2959), .ZN(n2918) );
  CLKBUF_X1 U2461 ( .A(n2541), .Z(n2222) );
  CLKBUF_X1 U2462 ( .A(n3742), .Z(n2218) );
  NOR2_X1 U2463 ( .A1(n2979), .A2(n2976), .ZN(n3742) );
  NAND2_X2 U2464 ( .A1(n5047), .A2(n2819), .ZN(n2904) );
  INV_X1 U2465 ( .A(n2918), .ZN(n2906) );
  INV_X1 U2466 ( .A(IR_REG_31__SCAN_IN), .ZN(n2964) );
  INV_X1 U2467 ( .A(n5070), .ZN(n5047) );
  AOI21_X2 U2469 ( .B1(n3730), .B2(n3726), .A(n3727), .ZN(n3648) );
  OAI21_X2 U2470 ( .B1(n3689), .B2(n3692), .A(n3690), .ZN(n3670) );
  NOR2_X1 U2471 ( .A1(n4216), .A2(n4193), .ZN(n4196) );
  NAND4_X1 U2472 ( .A1(n2605), .A2(n2604), .A3(n2603), .A4(n2602), .ZN(n3928)
         );
  NAND2_X1 U2473 ( .A1(n2559), .A2(n2558), .ZN(n3931) );
  CLKBUF_X3 U2474 ( .A(n2583), .Z(n2221) );
  BUF_X2 U2475 ( .A(n2540), .Z(n3137) );
  NAND2_X1 U2476 ( .A1(n2934), .A2(n2484), .ZN(n3112) );
  XNOR2_X1 U2477 ( .A(n2488), .B(n2487), .ZN(n2504) );
  AND3_X1 U2478 ( .A1(n2462), .A2(n2433), .A3(n2225), .ZN(n2477) );
  OR2_X1 U2479 ( .A1(n2950), .A2(n2946), .ZN(n2986) );
  AND2_X1 U2480 ( .A1(n2309), .A2(n2236), .ZN(n4750) );
  OR2_X1 U2481 ( .A1(n3467), .A2(n3846), .ZN(n3469) );
  NAND2_X1 U2482 ( .A1(n4216), .A2(n4193), .ZN(n4194) );
  NAND2_X1 U2483 ( .A1(n2446), .A2(n2641), .ZN(n3926) );
  AND4_X1 U2484 ( .A1(n2623), .A2(n2622), .A3(n2621), .A4(n2620), .ZN(n2627)
         );
  AND4_X1 U2485 ( .A1(n2545), .A2(n2544), .A3(n2543), .A4(n2542), .ZN(n3162)
         );
  AND4_X1 U2486 ( .A1(n2576), .A2(n2575), .A3(n2574), .A4(n2573), .ZN(n2580)
         );
  AND3_X1 U2487 ( .A1(n2557), .A2(n2556), .A3(n2555), .ZN(n2558) );
  CLKBUF_X3 U2488 ( .A(n2222), .Z(n2971) );
  INV_X2 U2489 ( .A(n2904), .ZN(n2915) );
  AND2_X2 U2490 ( .A1(n2471), .A2(n3118), .ZN(n2583) );
  INV_X2 U2491 ( .A(n2819), .ZN(n2920) );
  INV_X1 U2492 ( .A(n2472), .ZN(n3118) );
  AND2_X2 U2493 ( .A1(n3112), .A2(n3176), .ZN(n2819) );
  INV_X2 U2494 ( .A(n4791), .ZN(U4043) );
  AOI21_X1 U2495 ( .B1(n2967), .B2(n2242), .A(n2347), .ZN(n2346) );
  XNOR2_X1 U2496 ( .A(n2468), .B(n3614), .ZN(n2471) );
  AND2_X1 U2497 ( .A1(n2506), .A2(n2505), .ZN(n5039) );
  NAND2_X1 U2498 ( .A1(n2504), .A2(n3905), .ZN(n3176) );
  XNOR2_X1 U2499 ( .A(n2481), .B(n2480), .ZN(n2932) );
  XNOR2_X1 U2500 ( .A(n2502), .B(IR_REG_22__SCAN_IN), .ZN(n3913) );
  NAND2_X1 U2501 ( .A1(n2479), .A2(IR_REG_31__SCAN_IN), .ZN(n2481) );
  NAND2_X1 U2502 ( .A1(n2501), .A2(IR_REG_31__SCAN_IN), .ZN(n2488) );
  OR2_X1 U2503 ( .A1(n2477), .A2(n2964), .ZN(n2478) );
  NAND2_X1 U2504 ( .A1(n2462), .A2(n2461), .ZN(n2485) );
  INV_X1 U2505 ( .A(n2756), .ZN(n2462) );
  AND3_X1 U2506 ( .A1(n2458), .A2(n2281), .A3(n2563), .ZN(n2307) );
  NOR2_X1 U2507 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2514)
         );
  NOR2_X1 U2508 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2464)
         );
  OAI22_X1 U2509 ( .A1(n3162), .A2(n2905), .B1(n2920), .B2(n3301), .ZN(n2546)
         );
  OAI22_X1 U2510 ( .A1(n2627), .A2(n2905), .B1(n2920), .B2(n3340), .ZN(n2626)
         );
  BUF_X4 U2511 ( .A(n2591), .Z(n2905) );
  BUF_X4 U2512 ( .A(n2583), .Z(n2220) );
  INV_X1 U2514 ( .A(IR_REG_19__SCAN_IN), .ZN(n2498) );
  AOI21_X1 U2515 ( .B1(n2422), .B2(n2425), .A(n4099), .ZN(n2421) );
  INV_X1 U2516 ( .A(n4096), .ZN(n2425) );
  NOR2_X1 U2517 ( .A1(n2371), .A2(n3886), .ZN(n2368) );
  INV_X1 U2518 ( .A(n3479), .ZN(n3086) );
  NAND2_X1 U2519 ( .A1(n2963), .A2(n2493), .ZN(n2967) );
  NAND2_X1 U2520 ( .A1(n2435), .A2(n2466), .ZN(n2434) );
  INV_X1 U2521 ( .A(IR_REG_21__SCAN_IN), .ZN(n2466) );
  INV_X1 U2522 ( .A(n2465), .ZN(n2435) );
  NOR2_X1 U2523 ( .A1(n2588), .A2(n2306), .ZN(n2402) );
  NAND2_X1 U2524 ( .A1(n2460), .A2(n2459), .ZN(n2306) );
  NOR2_X1 U2525 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2378)
         );
  AND2_X1 U2526 ( .A1(n2898), .A2(REG3_REG_27__SCAN_IN), .ZN(n2908) );
  OR3_X1 U2527 ( .A1(n2850), .A2(n2849), .A3(n3717), .ZN(n2866) );
  AOI21_X1 U2528 ( .B1(n2485), .B2(IR_REG_31__SCAN_IN), .A(n2329), .ZN(n2328)
         );
  NAND2_X1 U2529 ( .A1(n2330), .A2(n2498), .ZN(n2329) );
  NAND2_X1 U2530 ( .A1(n2332), .A2(IR_REG_31__SCAN_IN), .ZN(n2330) );
  NAND2_X1 U2531 ( .A1(n2409), .A2(n2406), .ZN(n3099) );
  AOI21_X1 U2532 ( .B1(n2408), .B2(n2239), .A(n2407), .ZN(n2406) );
  NOR2_X1 U2533 ( .A1(n3036), .A2(n4031), .ZN(n2407) );
  NAND2_X1 U2534 ( .A1(n3851), .A2(n3033), .ZN(n3034) );
  INV_X1 U2535 ( .A(n3105), .ZN(n3088) );
  INV_X1 U2536 ( .A(IR_REG_28__SCAN_IN), .ZN(n2493) );
  INV_X1 U2537 ( .A(n2495), .ZN(n2494) );
  OR2_X1 U2538 ( .A1(n4935), .A2(n2299), .ZN(n2298) );
  NAND2_X1 U2539 ( .A1(n2300), .A2(n4381), .ZN(n2299) );
  NAND2_X1 U2540 ( .A1(n2297), .A2(n2300), .ZN(n2296) );
  INV_X1 U2541 ( .A(n2231), .ZN(n2297) );
  NAND2_X1 U2542 ( .A1(n3419), .A2(n2316), .ZN(n2315) );
  INV_X1 U2543 ( .A(n3487), .ZN(n2316) );
  INV_X1 U2544 ( .A(n3886), .ZN(n2369) );
  AND2_X1 U2545 ( .A1(n3879), .A2(n3062), .ZN(n2371) );
  OR2_X1 U2546 ( .A1(n2372), .A2(n3881), .ZN(n2370) );
  AND2_X1 U2547 ( .A1(n3749), .A2(n2373), .ZN(n2372) );
  INV_X1 U2548 ( .A(n3750), .ZN(n2373) );
  INV_X1 U2549 ( .A(n3737), .ZN(n2327) );
  NOR2_X1 U2550 ( .A1(n4852), .A2(n2280), .ZN(n2279) );
  INV_X1 U2551 ( .A(n4026), .ZN(n4029) );
  AOI21_X1 U2552 ( .B1(n2421), .B2(n2419), .A(n2246), .ZN(n2418) );
  INV_X1 U2553 ( .A(n2422), .ZN(n2419) );
  INV_X1 U2554 ( .A(n2421), .ZN(n2420) );
  NOR2_X1 U2555 ( .A1(n3865), .A2(n2437), .ZN(n2436) );
  INV_X1 U2556 ( .A(n3014), .ZN(n2437) );
  NOR2_X1 U2557 ( .A1(n3794), .A2(n2349), .ZN(n2348) );
  INV_X1 U2558 ( .A(n3770), .ZN(n2349) );
  OR2_X1 U2559 ( .A1(n3764), .A2(n2358), .ZN(n2357) );
  INV_X1 U2560 ( .A(n2357), .ZN(n2356) );
  AND2_X1 U2561 ( .A1(n3761), .A2(n3762), .ZN(n2360) );
  NAND2_X1 U2562 ( .A1(n2990), .A2(n3190), .ZN(n3752) );
  NAND2_X1 U2563 ( .A1(n2987), .A2(n3178), .ZN(n3755) );
  AND2_X1 U2564 ( .A1(n3913), .A2(n3905), .ZN(n3132) );
  AND2_X1 U2565 ( .A1(n3012), .A2(n2241), .ZN(n2439) );
  NOR2_X1 U2566 ( .A1(n3455), .A2(n3425), .ZN(n2387) );
  NOR2_X1 U2567 ( .A1(n3496), .A2(n3639), .ZN(n3477) );
  AND2_X1 U2568 ( .A1(n3041), .A2(n2991), .ZN(n2440) );
  NAND2_X1 U2569 ( .A1(n2477), .A2(n2467), .ZN(n2495) );
  INV_X1 U2570 ( .A(IR_REG_26__SCAN_IN), .ZN(n2467) );
  OAI21_X1 U2571 ( .B1(n2243), .B2(n3666), .A(n2327), .ZN(n2324) );
  INV_X1 U2572 ( .A(n2761), .ZN(n2308) );
  AND2_X1 U2573 ( .A1(n2961), .A2(n2960), .ZN(n3911) );
  NOR2_X1 U2574 ( .A1(n2932), .A2(n4709), .ZN(n2484) );
  NOR2_X1 U2575 ( .A1(n3936), .A2(n4720), .ZN(n3937) );
  NAND2_X1 U2576 ( .A1(n4725), .A2(n3969), .ZN(n2263) );
  NOR2_X1 U2577 ( .A1(n2266), .A2(n2390), .ZN(n2265) );
  INV_X1 U2578 ( .A(n2277), .ZN(n2271) );
  NOR2_X1 U2579 ( .A1(n5029), .A2(n2278), .ZN(n2277) );
  AND2_X1 U2580 ( .A1(n2276), .A2(n2275), .ZN(n2274) );
  OR2_X1 U2581 ( .A1(n5029), .A2(n3975), .ZN(n2276) );
  NAND2_X1 U2582 ( .A1(n2278), .A2(n2279), .ZN(n2275) );
  INV_X1 U2583 ( .A(n2279), .ZN(n2273) );
  XNOR2_X1 U2584 ( .A(n3948), .B(n4895), .ZN(n4890) );
  NAND2_X1 U2585 ( .A1(n4881), .A2(n2260), .ZN(n3982) );
  NAND2_X1 U2586 ( .A1(n3964), .A2(REG2_REG_11__SCAN_IN), .ZN(n2260) );
  AOI21_X1 U2587 ( .B1(n4902), .B2(n3984), .A(n2391), .ZN(n3985) );
  AND2_X1 U2588 ( .A1(n4900), .A2(REG2_REG_13__SCAN_IN), .ZN(n2391) );
  NAND2_X1 U2589 ( .A1(n2259), .A2(n2258), .ZN(n2257) );
  INV_X1 U2590 ( .A(n4922), .ZN(n2258) );
  INV_X1 U2591 ( .A(n2401), .ZN(n2399) );
  AND2_X1 U2592 ( .A1(n4009), .A2(n2910), .ZN(n4018) );
  INV_X1 U2593 ( .A(n3621), .ZN(n4038) );
  OR2_X1 U2594 ( .A1(n3816), .A2(n3817), .ZN(n4026) );
  NAND2_X1 U2595 ( .A1(n2414), .A2(n2412), .ZN(n2411) );
  INV_X1 U2596 ( .A(n3031), .ZN(n2412) );
  AND2_X1 U2597 ( .A1(n2885), .A2(n2884), .ZN(n2898) );
  NOR2_X1 U2598 ( .A1(n2866), .A2(n4503), .ZN(n2885) );
  OAI22_X1 U2599 ( .A1(n4077), .A2(n3029), .B1(n3694), .B2(n4110), .ZN(n4062)
         );
  AND2_X1 U2600 ( .A1(n2431), .A2(n3024), .ZN(n2430) );
  INV_X1 U2601 ( .A(n4181), .ZN(n2431) );
  NAND2_X1 U2602 ( .A1(n4204), .A2(n3023), .ZN(n2432) );
  AND2_X1 U2603 ( .A1(n2438), .A2(n2436), .ZN(n3562) );
  NOR2_X1 U2604 ( .A1(n3791), .A2(n2345), .ZN(n2344) );
  INV_X1 U2605 ( .A(n3790), .ZN(n2345) );
  AND2_X1 U2606 ( .A1(n3796), .A2(n3777), .ZN(n3865) );
  NAND2_X1 U2607 ( .A1(n3470), .A2(n3790), .ZN(n3454) );
  NAND2_X1 U2608 ( .A1(n3112), .A2(n3129), .ZN(n3170) );
  NAND2_X1 U2609 ( .A1(n3267), .A2(n3861), .ZN(n2361) );
  AND2_X1 U2610 ( .A1(n3762), .A2(n3766), .ZN(n3844) );
  NAND2_X1 U2611 ( .A1(n3292), .A2(n3756), .ZN(n3267) );
  AND2_X1 U2612 ( .A1(n3761), .A2(n3758), .ZN(n3861) );
  INV_X1 U2613 ( .A(n3041), .ZN(n3843) );
  NAND2_X1 U2614 ( .A1(n3859), .A2(n3164), .ZN(n3163) );
  NAND2_X1 U2615 ( .A1(n3755), .A2(n3752), .ZN(n3859) );
  AND2_X1 U2616 ( .A1(n3069), .A2(n3068), .ZN(n4213) );
  NAND2_X1 U2617 ( .A1(n3088), .A2(n3821), .ZN(n4230) );
  AND2_X1 U2618 ( .A1(n2230), .A2(n3106), .ZN(n2384) );
  NAND2_X1 U2619 ( .A1(n3594), .A2(n4731), .ZN(n4215) );
  NAND2_X1 U2620 ( .A1(n2935), .A2(n2934), .ZN(n3123) );
  NAND2_X1 U2621 ( .A1(n2444), .A2(IR_REG_31__SCAN_IN), .ZN(n2468) );
  NAND2_X1 U2622 ( .A1(n2444), .A2(n2346), .ZN(n2472) );
  NOR2_X1 U2623 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .ZN(n2347)
         );
  INV_X1 U2624 ( .A(IR_REG_23__SCAN_IN), .ZN(n2941) );
  INV_X1 U2625 ( .A(IR_REG_24__SCAN_IN), .ZN(n2480) );
  NAND4_X1 U2626 ( .A1(n2464), .A2(n2463), .A3(n2498), .A4(n2771), .ZN(n2465)
         );
  NAND2_X1 U2627 ( .A1(n2404), .A2(n2459), .ZN(n2727) );
  NOR2_X1 U2628 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2381)
         );
  NOR2_X1 U2629 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2379)
         );
  NOR2_X1 U2630 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2380)
         );
  AND2_X1 U2631 ( .A1(n2660), .A2(n2659), .ZN(n2685) );
  INV_X1 U2632 ( .A(IR_REG_1__SCAN_IN), .ZN(n2395) );
  OAI21_X1 U2633 ( .B1(n2525), .B2(n4716), .A(n2383), .ZN(n3294) );
  NAND2_X1 U2634 ( .A1(n2525), .A2(DATAI_2_), .ZN(n2383) );
  INV_X1 U2635 ( .A(n4189), .ZN(n4734) );
  INV_X1 U2636 ( .A(n4714), .ZN(n4774) );
  XNOR2_X1 U2637 ( .A(n3937), .B(n4718), .ZN(n4803) );
  NAND2_X1 U2638 ( .A1(n4830), .A2(n3974), .ZN(n4842) );
  NAND2_X1 U2639 ( .A1(n4882), .A2(n4883), .ZN(n4881) );
  XNOR2_X1 U2640 ( .A(n3982), .B(n4895), .ZN(n4892) );
  NAND2_X1 U2641 ( .A1(n4892), .A2(REG2_REG_12__SCAN_IN), .ZN(n4891) );
  OR2_X1 U2642 ( .A1(n4935), .A2(REG1_REG_16__SCAN_IN), .ZN(n2301) );
  INV_X1 U2643 ( .A(n4824), .ZN(n4955) );
  AND3_X1 U2644 ( .A1(n2298), .A2(n2296), .A3(n2255), .ZN(n4956) );
  NAND2_X1 U2645 ( .A1(n4950), .A2(n4951), .ZN(n2287) );
  NAND2_X1 U2646 ( .A1(n4941), .A2(n2401), .ZN(n4950) );
  AOI21_X1 U2647 ( .B1(n4941), .B2(n2253), .A(n4949), .ZN(n2286) );
  NAND2_X1 U2648 ( .A1(n2501), .A2(n2500), .ZN(n3998) );
  OAI21_X1 U2649 ( .B1(n2485), .B2(n2332), .A(IR_REG_31__SCAN_IN), .ZN(n2499)
         );
  XNOR2_X1 U2650 ( .A(n3099), .B(n3098), .ZN(n4016) );
  OR2_X1 U2651 ( .A1(n3170), .A2(n3081), .ZN(n4171) );
  INV_X1 U2652 ( .A(n4762), .ZN(n4223) );
  NOR2_X1 U2653 ( .A1(n2485), .A2(IR_REG_15__SCAN_IN), .ZN(n2790) );
  NAND2_X1 U2654 ( .A1(n5032), .A2(n5079), .ZN(n2294) );
  NAND2_X1 U2655 ( .A1(n2294), .A2(REG1_REG_6__SCAN_IN), .ZN(n2293) );
  AND2_X1 U2656 ( .A1(n2426), .A2(n2423), .ZN(n2422) );
  NAND2_X1 U2657 ( .A1(n2424), .A2(n4096), .ZN(n2423) );
  INV_X1 U2658 ( .A(n3837), .ZN(n2424) );
  INV_X1 U2659 ( .A(IR_REG_14__SCAN_IN), .ZN(n2460) );
  XNOR2_X1 U2660 ( .A(n2609), .B(n2906), .ZN(n2628) );
  AOI22_X1 U2661 ( .A1(n2312), .A2(n2317), .B1(n2311), .B2(n3420), .ZN(n2310)
         );
  INV_X1 U2662 ( .A(n2315), .ZN(n2311) );
  NAND2_X1 U2663 ( .A1(n2750), .A2(n2319), .ZN(n2317) );
  OR2_X1 U2664 ( .A1(n2747), .A2(n2318), .ZN(n2312) );
  OR2_X1 U2665 ( .A1(n2314), .A2(n2747), .ZN(n2313) );
  NAND2_X1 U2666 ( .A1(n2750), .A2(n2315), .ZN(n2314) );
  NAND2_X1 U2667 ( .A1(n2292), .A2(n2290), .ZN(n3942) );
  NAND2_X1 U2668 ( .A1(n2291), .A2(n2294), .ZN(n2290) );
  OR2_X1 U2669 ( .A1(n4826), .A2(n2293), .ZN(n2292) );
  NAND2_X1 U2670 ( .A1(n2234), .A2(n4834), .ZN(n2291) );
  NAND2_X1 U2671 ( .A1(n3988), .A2(REG2_REG_15__SCAN_IN), .ZN(n2256) );
  NAND2_X1 U2672 ( .A1(n3991), .A2(REG2_REG_18__SCAN_IN), .ZN(n2400) );
  INV_X1 U2673 ( .A(n3037), .ZN(n2410) );
  NOR2_X1 U2674 ( .A1(n2414), .A2(n3037), .ZN(n2408) );
  AND2_X1 U2675 ( .A1(n3884), .A2(n2367), .ZN(n2366) );
  NAND2_X1 U2676 ( .A1(n2370), .A2(n2368), .ZN(n2367) );
  NAND2_X1 U2677 ( .A1(n2365), .A2(n2370), .ZN(n4144) );
  NAND2_X1 U2678 ( .A1(n2375), .A2(n2371), .ZN(n2365) );
  INV_X1 U2679 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2648) );
  NOR2_X1 U2680 ( .A1(n3033), .A2(n3671), .ZN(n2385) );
  AND2_X1 U2681 ( .A1(n3087), .A2(n4152), .ZN(n2389) );
  AND2_X1 U2682 ( .A1(n4169), .A2(n4168), .ZN(n3087) );
  NAND2_X1 U2683 ( .A1(n2486), .A2(n2771), .ZN(n2334) );
  INV_X1 U2684 ( .A(IR_REG_17__SCAN_IN), .ZN(n2486) );
  NOR2_X1 U2685 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2723)
         );
  NOR2_X1 U2686 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2382)
         );
  NOR2_X1 U2687 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2655)
         );
  AND2_X1 U2688 ( .A1(n2666), .A2(REG3_REG_10__SCAN_IN), .ZN(n2679) );
  XNOR2_X1 U2689 ( .A(n2567), .B(n2906), .ZN(n2569) );
  INV_X1 U2690 ( .A(n4051), .ZN(n3036) );
  AND2_X1 U2691 ( .A1(n3819), .A2(DATAI_21_), .ZN(n3660) );
  XNOR2_X1 U2692 ( .A(n2592), .B(n2918), .ZN(n2595) );
  OAI22_X1 U2693 ( .A1(n2996), .A2(n2591), .B1(n2920), .B2(n3258), .ZN(n2592)
         );
  NOR2_X1 U2694 ( .A1(n3332), .A2(n2336), .ZN(n2335) );
  INV_X1 U2695 ( .A(n2338), .ZN(n2336) );
  NAND2_X1 U2696 ( .A1(n3221), .A2(n3222), .ZN(n2338) );
  NAND2_X1 U2697 ( .A1(n3220), .A2(n2339), .ZN(n2337) );
  OR2_X1 U2698 ( .A1(n3221), .A2(n3222), .ZN(n2339) );
  AND2_X1 U2699 ( .A1(n2796), .A2(n2795), .ZN(n2797) );
  AND3_X1 U2700 ( .A1(n3140), .A2(n3139), .A3(n3138), .ZN(n3900) );
  OR2_X1 U2701 ( .A1(n4782), .A2(n4781), .ZN(n2289) );
  AND2_X1 U2702 ( .A1(n2289), .A2(n2288), .ZN(n3935) );
  NAND2_X1 U2703 ( .A1(n4784), .A2(REG1_REG_2__SCAN_IN), .ZN(n2288) );
  OR2_X1 U2704 ( .A1(n4826), .A2(n4827), .ZN(n2295) );
  XNOR2_X1 U2705 ( .A(n3942), .B(n4852), .ZN(n4847) );
  NAND2_X1 U2706 ( .A1(n4878), .A2(n3947), .ZN(n3948) );
  NAND2_X1 U2707 ( .A1(n4906), .A2(n3950), .ZN(n3951) );
  OR2_X1 U2708 ( .A1(n4912), .A2(n3986), .ZN(n2259) );
  INV_X1 U2709 ( .A(n5018), .ZN(n3988) );
  NAND2_X1 U2710 ( .A1(n4926), .A2(n3953), .ZN(n3954) );
  AND2_X1 U2711 ( .A1(n3819), .A2(n3133), .ZN(n3962) );
  OR2_X1 U2712 ( .A1(n3990), .A2(REG2_REG_17__SCAN_IN), .ZN(n2401) );
  NAND2_X1 U2713 ( .A1(n2333), .A2(n2463), .ZN(n2332) );
  INV_X1 U2714 ( .A(n2334), .ZN(n2333) );
  INV_X1 U2715 ( .A(n2400), .ZN(n2397) );
  AOI21_X1 U2716 ( .B1(n3100), .B2(n3066), .A(n3818), .ZN(n3067) );
  OAI21_X1 U2717 ( .B1(n4045), .B2(n2342), .A(n2340), .ZN(n3100) );
  AOI21_X1 U2718 ( .B1(n2341), .B2(n3809), .A(n3817), .ZN(n2340) );
  NAND2_X1 U2719 ( .A1(n2343), .A2(n2341), .ZN(n4028) );
  NAND2_X1 U2720 ( .A1(n2417), .A2(n2416), .ZN(n4077) );
  AOI21_X1 U2721 ( .B1(n2418), .B2(n2420), .A(n2245), .ZN(n2416) );
  AND2_X1 U2722 ( .A1(n4122), .A2(n4132), .ZN(n4124) );
  NAND2_X1 U2723 ( .A1(n3027), .A2(n3837), .ZN(n4141) );
  NAND2_X1 U2724 ( .A1(n2374), .A2(n3749), .ZN(n4159) );
  NAND2_X1 U2725 ( .A1(n2375), .A2(n3879), .ZN(n2374) );
  NOR2_X1 U2726 ( .A1(n2827), .A2(n2469), .ZN(n2829) );
  NAND2_X1 U2727 ( .A1(n2801), .A2(REG3_REG_18__SCAN_IN), .ZN(n2827) );
  INV_X1 U2728 ( .A(n2430), .ZN(n2429) );
  AOI21_X1 U2729 ( .B1(n2430), .B2(n2428), .A(n2244), .ZN(n2427) );
  INV_X1 U2730 ( .A(n3023), .ZN(n2428) );
  AND2_X1 U2731 ( .A1(n2454), .A2(n3858), .ZN(n4205) );
  NAND2_X1 U2732 ( .A1(n2751), .A2(REG3_REG_15__SCAN_IN), .ZN(n2763) );
  AND2_X1 U2733 ( .A1(n3876), .A2(n3878), .ZN(n3864) );
  AND4_X1 U2734 ( .A1(n2770), .A2(n2769), .A3(n2768), .A4(n2767), .ZN(n3567)
         );
  NOR2_X1 U2735 ( .A1(n2717), .A2(n3424), .ZN(n2738) );
  NAND2_X1 U2736 ( .A1(n2679), .A2(REG3_REG_11__SCAN_IN), .ZN(n2702) );
  OR2_X1 U2737 ( .A1(n2702), .A2(n2701), .ZN(n2717) );
  AND2_X1 U2738 ( .A1(n3453), .A2(n3790), .ZN(n3846) );
  NAND2_X1 U2739 ( .A1(n3049), .A2(n3793), .ZN(n3470) );
  INV_X1 U2740 ( .A(n4211), .ZN(n4188) );
  AND4_X1 U2741 ( .A1(n2684), .A2(n2683), .A3(n2682), .A4(n2681), .ZN(n3505)
         );
  NAND2_X1 U2742 ( .A1(n2350), .A2(n3770), .ZN(n3400) );
  INV_X1 U2743 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4628) );
  AND2_X1 U2744 ( .A1(n3044), .A2(n3771), .ZN(n3845) );
  NOR2_X1 U2745 ( .A1(n2600), .A2(n4415), .ZN(n2618) );
  INV_X1 U2746 ( .A(REG3_REG_6__SCAN_IN), .ZN(n4415) );
  NAND2_X1 U2747 ( .A1(n2355), .A2(n2353), .ZN(n3357) );
  INV_X1 U2748 ( .A(n2354), .ZN(n2353) );
  OAI21_X1 U2749 ( .B1(n2360), .B2(n2357), .A(n3781), .ZN(n2354) );
  INV_X1 U2750 ( .A(n4208), .ZN(n4185) );
  OAI211_X1 U2751 ( .C1(n3267), .C2(n2352), .A(n2351), .B(n3766), .ZN(n3257)
         );
  INV_X1 U2752 ( .A(n2360), .ZN(n2352) );
  NAND2_X1 U2753 ( .A1(n2359), .A2(n2360), .ZN(n2351) );
  INV_X1 U2754 ( .A(n3861), .ZN(n2359) );
  INV_X1 U2755 ( .A(n3320), .ZN(n3315) );
  NAND2_X1 U2756 ( .A1(n3843), .A2(n2362), .ZN(n3292) );
  OAI21_X1 U2757 ( .B1(n3859), .B2(n3203), .A(n3755), .ZN(n3293) );
  INV_X1 U2758 ( .A(n4213), .ZN(n4183) );
  NAND2_X1 U2759 ( .A1(n3994), .A2(n3132), .ZN(n4208) );
  NAND2_X1 U2760 ( .A1(n4711), .A2(n5039), .ZN(n4207) );
  NOR2_X1 U2761 ( .A1(n4230), .A2(n4232), .ZN(n4229) );
  INV_X1 U2762 ( .A(n4207), .ZN(n4231) );
  NAND2_X1 U2763 ( .A1(n4089), .A2(n2385), .ZN(n4054) );
  NAND2_X1 U2764 ( .A1(n4089), .A2(n4069), .ZN(n4071) );
  AND2_X1 U2765 ( .A1(n4113), .A2(n4087), .ZN(n4089) );
  NAND2_X1 U2766 ( .A1(n3819), .A2(DATAI_24_), .ZN(n4087) );
  AND2_X1 U2767 ( .A1(n4196), .A2(n2388), .ZN(n4113) );
  AND2_X1 U2768 ( .A1(n2229), .A2(n4115), .ZN(n2388) );
  NAND2_X1 U2769 ( .A1(n4196), .A2(n2229), .ZN(n4126) );
  NAND2_X1 U2770 ( .A1(n4196), .A2(n2389), .ZN(n4151) );
  INV_X1 U2771 ( .A(n3660), .ZN(n4152) );
  NAND2_X1 U2772 ( .A1(n3819), .A2(DATAI_20_), .ZN(n4168) );
  INV_X1 U2773 ( .A(n3646), .ZN(n4169) );
  OR2_X1 U2774 ( .A1(n4215), .A2(n3682), .ZN(n4216) );
  AND2_X1 U2775 ( .A1(n3478), .A2(n2228), .ZN(n3594) );
  NAND2_X1 U2776 ( .A1(n2438), .A2(n3014), .ZN(n3526) );
  NAND2_X1 U2777 ( .A1(n3478), .A2(n2387), .ZN(n3539) );
  AND2_X1 U2778 ( .A1(n3477), .A2(n3086), .ZN(n3478) );
  NAND2_X1 U2779 ( .A1(n3478), .A2(n3461), .ZN(n3538) );
  OR2_X1 U2780 ( .A1(n3441), .A2(n3405), .ZN(n3496) );
  NOR2_X1 U2781 ( .A1(n3367), .A2(n3345), .ZN(n3440) );
  OR2_X1 U2782 ( .A1(n3365), .A2(n3364), .ZN(n3367) );
  OR2_X1 U2783 ( .A1(n3314), .A2(n3254), .ZN(n3365) );
  INV_X1 U2784 ( .A(n3258), .ZN(n3254) );
  NOR2_X1 U2785 ( .A1(n3300), .A2(n3274), .ZN(n3316) );
  NOR2_X1 U2786 ( .A1(n3178), .A2(n3179), .ZN(n3302) );
  NAND2_X1 U2787 ( .A1(n3302), .A2(n3301), .ZN(n3300) );
  INV_X1 U2788 ( .A(n3294), .ZN(n3301) );
  NAND2_X1 U2789 ( .A1(n3163), .A2(n2991), .ZN(n3291) );
  NAND2_X1 U2790 ( .A1(n2495), .A2(IR_REG_31__SCAN_IN), .ZN(n3073) );
  NOR2_X1 U2791 ( .A1(n2223), .A2(IR_REG_16__SCAN_IN), .ZN(n2377) );
  AND2_X1 U2792 ( .A1(n2642), .A2(n2625), .ZN(n4835) );
  INV_X1 U2793 ( .A(IR_REG_4__SCAN_IN), .ZN(n2458) );
  OR2_X1 U2794 ( .A1(n2908), .A2(n2899), .ZN(n3621) );
  NAND2_X1 U2795 ( .A1(n2320), .A2(n2324), .ZN(n3618) );
  OAI21_X1 U2796 ( .B1(n3423), .B2(n3420), .A(n3419), .ZN(n3489) );
  AND2_X1 U2797 ( .A1(n3625), .A2(n3626), .ZN(n2862) );
  AND4_X1 U2798 ( .A1(n2805), .A2(n2804), .A3(n2803), .A4(n2802), .ZN(n4209)
         );
  OAI21_X1 U2799 ( .B1(n3670), .B2(n2323), .A(n2321), .ZN(n2950) );
  INV_X1 U2800 ( .A(n2324), .ZN(n2323) );
  AND2_X1 U2801 ( .A1(n3617), .A2(n2322), .ZN(n2321) );
  NAND2_X1 U2802 ( .A1(n2326), .A2(n2324), .ZN(n2322) );
  INV_X1 U2803 ( .A(n3178), .ZN(n3190) );
  AND4_X1 U2804 ( .A1(n2847), .A2(n2846), .A3(n2845), .A4(n2844), .ZN(n4142)
         );
  INV_X1 U2805 ( .A(n3021), .ZN(n4731) );
  OAI21_X1 U2806 ( .B1(n4748), .B2(n2782), .A(n2781), .ZN(n3681) );
  NAND2_X1 U2807 ( .A1(n2778), .A2(n2780), .ZN(n2781) );
  INV_X1 U2808 ( .A(n2779), .ZN(n2780) );
  AND4_X1 U2809 ( .A1(n2880), .A2(n2879), .A3(n2878), .A4(n2877), .ZN(n4083)
         );
  INV_X1 U2810 ( .A(n3926), .ZN(n3341) );
  NAND2_X1 U2811 ( .A1(n2337), .A2(n2338), .ZN(n3331) );
  INV_X1 U2812 ( .A(n4743), .ZN(n3741) );
  AND4_X1 U2813 ( .A1(n2744), .A2(n2743), .A3(n2742), .A4(n2741), .ZN(n4745)
         );
  INV_X1 U2814 ( .A(n3705), .ZN(n4743) );
  INV_X1 U2815 ( .A(n3900), .ZN(n4004) );
  NAND4_X1 U2816 ( .A1(n2871), .A2(n2870), .A3(n2869), .A4(n2868), .ZN(n4110)
         );
  INV_X1 U2817 ( .A(n4158), .ZN(n3707) );
  INV_X1 U2818 ( .A(n3567), .ZN(n4747) );
  INV_X1 U2819 ( .A(n4745), .ZN(n3923) );
  NAND4_X1 U2820 ( .A1(n2721), .A2(n2720), .A3(n2719), .A4(n2718), .ZN(n3523)
         );
  INV_X1 U2821 ( .A(n3505), .ZN(n3640) );
  INV_X1 U2822 ( .A(n2627), .ZN(n3927) );
  INV_X1 U2823 ( .A(n2580), .ZN(n3930) );
  CLKBUF_X1 U2824 ( .A(n2988), .Z(n2990) );
  NAND2_X1 U2825 ( .A1(n2540), .A2(REG2_REG_0__SCAN_IN), .ZN(n2524) );
  OR2_X1 U2826 ( .A1(n3112), .A2(n5010), .ZN(n4791) );
  XNOR2_X1 U2827 ( .A(n3935), .B(n4729), .ZN(n4721) );
  AND2_X1 U2828 ( .A1(n4803), .A2(REG1_REG_4__SCAN_IN), .ZN(n4809) );
  NAND2_X1 U2829 ( .A1(n4805), .A2(REG2_REG_4__SCAN_IN), .ZN(n4804) );
  NAND2_X1 U2830 ( .A1(n2267), .A2(n2264), .ZN(n4805) );
  OAI21_X1 U2831 ( .B1(n2262), .B2(n2261), .A(n3971), .ZN(n4819) );
  NAND2_X1 U2832 ( .A1(n3938), .A2(n2304), .ZN(n2302) );
  INV_X1 U2833 ( .A(n4814), .ZN(n2304) );
  NOR2_X1 U2834 ( .A1(n4809), .A2(n3938), .ZN(n4815) );
  AND2_X1 U2835 ( .A1(n2295), .A2(n2234), .ZN(n4838) );
  OAI211_X1 U2836 ( .C1(n4842), .C2(n2272), .A(REG2_REG_8__SCAN_IN), .B(n2269), 
        .ZN(n4848) );
  NAND2_X1 U2837 ( .A1(n2274), .A2(n2273), .ZN(n2272) );
  AND2_X1 U2838 ( .A1(n2271), .A2(n2274), .ZN(n2270) );
  OAI211_X1 U2839 ( .C1(n4842), .C2(n2273), .A(n2274), .B(n2268), .ZN(n4849)
         );
  NAND2_X1 U2840 ( .A1(n4842), .A2(n2277), .ZN(n2268) );
  NAND2_X1 U2841 ( .A1(n4871), .A2(n3981), .ZN(n4882) );
  NAND2_X1 U2842 ( .A1(n4891), .A2(n3983), .ZN(n4902) );
  NOR2_X1 U2843 ( .A1(n4913), .A2(n3533), .ZN(n4912) );
  INV_X1 U2844 ( .A(n2257), .ZN(n4921) );
  INV_X1 U2845 ( .A(n2259), .ZN(n4923) );
  INV_X1 U2846 ( .A(n4952), .ZN(n2284) );
  OR2_X1 U2847 ( .A1(n4768), .A2(n4787), .ZN(n4824) );
  NAND2_X1 U2848 ( .A1(n2398), .A2(n2396), .ZN(n3993) );
  OR2_X1 U2849 ( .A1(n2253), .A2(n2397), .ZN(n2396) );
  OAI21_X1 U2850 ( .B1(n3032), .B2(n2413), .A(n2239), .ZN(n4027) );
  OR2_X1 U2851 ( .A1(n2898), .A2(n2886), .ZN(n4057) );
  NAND2_X1 U2852 ( .A1(n2432), .A2(n2430), .ZN(n4180) );
  NAND2_X1 U2853 ( .A1(n2432), .A2(n3024), .ZN(n4178) );
  NAND2_X1 U2854 ( .A1(n3478), .A2(n2227), .ZN(n4290) );
  NAND2_X1 U2855 ( .A1(n2361), .A2(n3761), .ZN(n3317) );
  INV_X1 U2856 ( .A(n3179), .ZN(n5040) );
  INV_X1 U2857 ( .A(n5010), .ZN(n3129) );
  AND2_X1 U2858 ( .A1(n2442), .A2(n2492), .ZN(n2441) );
  AND2_X1 U2859 ( .A1(n2493), .A2(n2443), .ZN(n2442) );
  INV_X1 U2860 ( .A(IR_REG_29__SCAN_IN), .ZN(n2443) );
  INV_X1 U2861 ( .A(IR_REG_30__SCAN_IN), .ZN(n3614) );
  INV_X1 U2862 ( .A(n3994), .ZN(n4789) );
  NAND2_X1 U2863 ( .A1(n3131), .A2(STATE_REG_SCAN_IN), .ZN(n5010) );
  OAI21_X1 U2864 ( .B1(n2485), .B2(n2465), .A(IR_REG_31__SCAN_IN), .ZN(n2489)
         );
  INV_X1 U2865 ( .A(n3998), .ZN(n4712) );
  NOR2_X1 U2866 ( .A1(n2727), .A2(n2405), .ZN(n2745) );
  NOR2_X1 U2867 ( .A1(n2661), .A2(n2685), .ZN(n4856) );
  OR2_X1 U2868 ( .A1(n2514), .A2(n2964), .ZN(n2282) );
  NAND2_X1 U2869 ( .A1(n2515), .A2(n2392), .ZN(n4714) );
  AND2_X1 U2870 ( .A1(n2394), .A2(n2393), .ZN(n2392) );
  INV_X1 U2871 ( .A(IR_REG_0__SCAN_IN), .ZN(n5038) );
  NAND2_X1 U2872 ( .A1(n2296), .A2(n2298), .ZN(n4946) );
  AOI21_X1 U2873 ( .B1(n2287), .B2(n2286), .A(n2283), .ZN(n4959) );
  NAND2_X1 U2874 ( .A1(n2285), .A2(n2284), .ZN(n2283) );
  AOI211_X1 U2875 ( .C1(n4023), .C2(n4223), .A(n4022), .B(n4021), .ZN(n4024)
         );
  OR2_X1 U2876 ( .A1(n4010), .A2(n4288), .ZN(n3095) );
  OR2_X1 U2877 ( .A1(n4017), .A2(n4288), .ZN(n3107) );
  AND2_X1 U2878 ( .A1(n3090), .A2(n3089), .ZN(n3091) );
  OR2_X1 U2879 ( .A1(n4017), .A2(n4706), .ZN(n3110) );
  AND2_X1 U2880 ( .A1(n3919), .A2(n3671), .ZN(n3030) );
  MUX2_X2 U2881 ( .A(n2497), .B(n2496), .S(n3073), .Z(n2525) );
  AND2_X2 U2882 ( .A1(n3112), .A2(n2491), .ZN(n2513) );
  INV_X1 U2883 ( .A(n4843), .ZN(n2278) );
  INV_X1 U2884 ( .A(n4718), .ZN(n2390) );
  NAND2_X1 U2885 ( .A1(n2941), .A2(n2480), .ZN(n2223) );
  NAND3_X1 U2886 ( .A1(n2462), .A2(n2433), .A3(n2461), .ZN(n2224) );
  AND2_X1 U2887 ( .A1(n2377), .A2(n2376), .ZN(n2225) );
  AND2_X1 U2888 ( .A1(n2343), .A2(n3893), .ZN(n2226) );
  AND2_X1 U2889 ( .A1(n2387), .A2(n3015), .ZN(n2227) );
  AND2_X1 U2890 ( .A1(n2227), .A2(n4742), .ZN(n2228) );
  INV_X1 U2891 ( .A(n3030), .ZN(n2415) );
  AND2_X1 U2892 ( .A1(n2389), .A2(n3718), .ZN(n2229) );
  AND2_X1 U2893 ( .A1(n2385), .A2(n4031), .ZN(n2230) );
  NOR2_X1 U2894 ( .A1(n2471), .A2(n2472), .ZN(n2541) );
  AND4_X1 U2895 ( .A1(n2587), .A2(n2586), .A3(n2585), .A4(n2584), .ZN(n2996)
         );
  AND2_X1 U2896 ( .A1(n3121), .A2(n2472), .ZN(n2540) );
  OR2_X1 U2897 ( .A1(n5015), .A2(n3954), .ZN(n2231) );
  AND2_X1 U2898 ( .A1(n2539), .A2(n2538), .ZN(n2232) );
  INV_X1 U2899 ( .A(n3420), .ZN(n2319) );
  AND2_X1 U2900 ( .A1(n2734), .A2(n2735), .ZN(n3420) );
  OR2_X1 U2901 ( .A1(n2485), .A2(n2434), .ZN(n2233) );
  OR2_X1 U2902 ( .A1(n3941), .A2(n3940), .ZN(n2234) );
  AND2_X1 U2903 ( .A1(n2564), .A2(n2577), .ZN(n3967) );
  INV_X1 U2904 ( .A(n3967), .ZN(n4729) );
  AND2_X1 U2905 ( .A1(n2257), .A2(n2256), .ZN(n2235) );
  INV_X1 U2906 ( .A(IR_REG_15__SCAN_IN), .ZN(n2771) );
  INV_X1 U2907 ( .A(IR_REG_16__SCAN_IN), .ZN(n2461) );
  INV_X1 U2908 ( .A(n2342), .ZN(n2341) );
  NAND2_X1 U2909 ( .A1(n4029), .A2(n3893), .ZN(n2342) );
  AND2_X1 U2910 ( .A1(n2310), .A2(n2308), .ZN(n2236) );
  AND2_X1 U2911 ( .A1(n4774), .A2(REG1_REG_1__SCAN_IN), .ZN(n2237) );
  AND2_X1 U2912 ( .A1(n2301), .A2(n2231), .ZN(n2238) );
  INV_X1 U2913 ( .A(IR_REG_3__SCAN_IN), .ZN(n2563) );
  INV_X1 U2914 ( .A(IR_REG_2__SCAN_IN), .ZN(n2281) );
  NAND2_X1 U2915 ( .A1(n3013), .A2(n2439), .ZN(n2438) );
  AND2_X1 U2916 ( .A1(n2411), .A2(n3035), .ZN(n2239) );
  INV_X1 U2917 ( .A(IR_REG_7__SCAN_IN), .ZN(n2459) );
  AND2_X1 U2918 ( .A1(n4196), .A2(n3087), .ZN(n4150) );
  NAND2_X1 U2919 ( .A1(n2307), .A2(n2514), .ZN(n2588) );
  AND2_X1 U2920 ( .A1(n4089), .A2(n2230), .ZN(n2240) );
  AND2_X1 U2921 ( .A1(n3603), .A2(n3059), .ZN(n3879) );
  NAND2_X1 U2922 ( .A1(n3469), .A2(n3010), .ZN(n3459) );
  INV_X1 U2923 ( .A(IR_REG_25__SCAN_IN), .ZN(n2376) );
  INV_X1 U2924 ( .A(n5029), .ZN(n4852) );
  OR2_X1 U2925 ( .A1(n3523), .A2(n3425), .ZN(n2241) );
  INV_X1 U2926 ( .A(n4716), .ZN(n4784) );
  XNOR2_X1 U2927 ( .A(n2282), .B(n2281), .ZN(n4716) );
  AND2_X1 U2928 ( .A1(IR_REG_29__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2242)
         );
  NOR2_X1 U2929 ( .A1(n2897), .A2(n2896), .ZN(n2243) );
  INV_X1 U2930 ( .A(n2414), .ZN(n2413) );
  AND2_X1 U2931 ( .A1(n2415), .A2(n3034), .ZN(n2414) );
  AND2_X1 U2932 ( .A1(n4209), .A2(n3025), .ZN(n2244) );
  NOR2_X1 U2933 ( .A1(n3720), .A2(n4115), .ZN(n2245) );
  NOR2_X1 U2934 ( .A1(n4135), .A2(n3630), .ZN(n2246) );
  AND2_X1 U2935 ( .A1(n3679), .A2(n2797), .ZN(n2247) );
  INV_X1 U2936 ( .A(n2326), .ZN(n2325) );
  NAND2_X1 U2937 ( .A1(n2327), .A2(n3667), .ZN(n2326) );
  NAND2_X1 U2938 ( .A1(n3925), .A2(n3405), .ZN(n2248) );
  NOR2_X1 U2939 ( .A1(n4814), .A2(n2305), .ZN(n2249) );
  AND2_X1 U2940 ( .A1(n2436), .A2(n3016), .ZN(n2250) );
  AND2_X1 U2941 ( .A1(n2370), .A2(n2369), .ZN(n2251) );
  AND2_X1 U2942 ( .A1(n2239), .A2(n2410), .ZN(n2252) );
  XNOR2_X1 U2943 ( .A(n2478), .B(IR_REG_26__SCAN_IN), .ZN(n2934) );
  NAND2_X1 U2944 ( .A1(n2337), .A2(n2335), .ZN(n3329) );
  AND2_X1 U2945 ( .A1(n2494), .A2(n2492), .ZN(n2963) );
  AND2_X1 U2946 ( .A1(n3819), .A2(DATAI_22_), .ZN(n4134) );
  INV_X1 U2947 ( .A(n4115), .ZN(n3630) );
  INV_X1 U2948 ( .A(n2331), .ZN(n2806) );
  NOR2_X1 U2949 ( .A1(n2485), .A2(n2334), .ZN(n2331) );
  INV_X1 U2950 ( .A(n4945), .ZN(n2300) );
  NOR2_X1 U2951 ( .A1(n2399), .A2(n4951), .ZN(n2253) );
  INV_X1 U2952 ( .A(n4031), .ZN(n4036) );
  INV_X1 U2953 ( .A(n3671), .ZN(n4069) );
  AND2_X1 U2954 ( .A1(n3819), .A2(DATAI_25_), .ZN(n3671) );
  INV_X1 U2955 ( .A(n3766), .ZN(n2358) );
  AND2_X1 U2956 ( .A1(n4942), .A2(n2400), .ZN(n2254) );
  OR2_X1 U2957 ( .A1(n3990), .A2(REG1_REG_17__SCAN_IN), .ZN(n2255) );
  INV_X1 U2958 ( .A(n3106), .ZN(n2386) );
  INV_X1 U2959 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2305) );
  NAND2_X1 U2960 ( .A1(n4953), .A2(ADDR_REG_18__SCAN_IN), .ZN(n2285) );
  NAND2_X1 U2961 ( .A1(n2265), .A2(n4725), .ZN(n2264) );
  NAND2_X1 U2962 ( .A1(n2263), .A2(n2390), .ZN(n2267) );
  OAI21_X1 U2963 ( .B1(n4725), .B2(n2390), .A(REG2_REG_4__SCAN_IN), .ZN(n2261)
         );
  AOI21_X1 U2964 ( .B1(n2263), .B2(n2390), .A(n2265), .ZN(n2262) );
  NAND2_X1 U2965 ( .A1(n4725), .A2(n3969), .ZN(n3970) );
  INV_X1 U2966 ( .A(n3969), .ZN(n2266) );
  NAND2_X1 U2967 ( .A1(n4842), .A2(n2270), .ZN(n2269) );
  NAND2_X1 U2968 ( .A1(n4842), .A2(n4843), .ZN(n4841) );
  NAND2_X1 U2969 ( .A1(n4841), .A2(n3975), .ZN(n3976) );
  INV_X1 U2970 ( .A(n3975), .ZN(n2280) );
  INV_X1 U2971 ( .A(n2289), .ZN(n4780) );
  NOR2_X1 U2972 ( .A1(n4770), .A2(n2237), .ZN(n4782) );
  INV_X1 U2973 ( .A(n2295), .ZN(n4825) );
  INV_X1 U2974 ( .A(n2301), .ZN(n4936) );
  NAND2_X1 U2975 ( .A1(n4803), .A2(n2249), .ZN(n2303) );
  NAND2_X1 U2976 ( .A1(n2303), .A2(n2302), .ZN(n4813) );
  NAND2_X1 U2977 ( .A1(n3423), .A2(n2313), .ZN(n2309) );
  NAND2_X1 U2978 ( .A1(n2309), .A2(n2310), .ZN(n2762) );
  INV_X1 U2979 ( .A(n2750), .ZN(n2318) );
  NAND2_X1 U2980 ( .A1(n3670), .A2(n2325), .ZN(n2320) );
  AOI21_X1 U2981 ( .B1(n3670), .B2(n3667), .A(n3666), .ZN(n3739) );
  INV_X1 U2982 ( .A(n2328), .ZN(n2501) );
  NAND2_X1 U2983 ( .A1(n2716), .A2(n2715), .ZN(n3423) );
  NAND2_X1 U2984 ( .A1(n3714), .A2(n3715), .ZN(n3713) );
  AND2_X2 U2985 ( .A1(n3713), .A2(n2862), .ZN(n3628) );
  NOR2_X2 U2986 ( .A1(n4750), .A2(n4749), .ZN(n4748) );
  OAI21_X1 U2987 ( .B1(n3374), .B2(n3376), .A(n3375), .ZN(n2716) );
  OAI22_X2 U2988 ( .A1(n3648), .A2(n3649), .B1(n2825), .B2(n2824), .ZN(n3703)
         );
  NAND2_X1 U2989 ( .A1(n2700), .A2(n2699), .ZN(n3374) );
  NAND2_X1 U2990 ( .A1(n3280), .A2(n2636), .ZN(n3220) );
  NOR2_X2 U2991 ( .A1(n3628), .A2(n2452), .ZN(n3689) );
  NAND2_X1 U2992 ( .A1(n3279), .A2(n2633), .ZN(n3280) );
  NAND2_X1 U2993 ( .A1(n2534), .A2(n2533), .ZN(n3188) );
  NAND2_X1 U2994 ( .A1(n2232), .A2(n3156), .ZN(n3155) );
  AOI21_X1 U2995 ( .B1(n3656), .B2(n3657), .A(n2843), .ZN(n3714) );
  OAI21_X1 U2996 ( .B1(n3681), .B2(n2247), .A(n2799), .ZN(n2800) );
  NAND2_X1 U2997 ( .A1(n2395), .A2(n2964), .ZN(n2394) );
  XNOR2_X1 U2998 ( .A(n3960), .B(n3959), .ZN(n4002) );
  NAND2_X1 U2999 ( .A1(n4954), .A2(n2447), .ZN(n3960) );
  XNOR2_X1 U3000 ( .A(n3941), .B(n3940), .ZN(n4826) );
  NAND2_X1 U3001 ( .A1(n2517), .A2(n2516), .ZN(n2518) );
  NAND2_X1 U3002 ( .A1(n4045), .A2(n3897), .ZN(n2343) );
  XNOR2_X1 U3003 ( .A(n3100), .B(n3855), .ZN(n3103) );
  NAND2_X1 U3004 ( .A1(n3470), .A2(n2344), .ZN(n3053) );
  NAND2_X1 U3005 ( .A1(n2350), .A2(n2348), .ZN(n3048) );
  NAND2_X1 U3006 ( .A1(n3433), .A2(n3773), .ZN(n2350) );
  NAND3_X1 U3007 ( .A1(n3861), .A2(n3267), .A3(n2356), .ZN(n2355) );
  INV_X1 U3008 ( .A(n3752), .ZN(n2363) );
  OAI21_X1 U3009 ( .B1(n3203), .B2(n2363), .A(n3755), .ZN(n2362) );
  INV_X1 U3010 ( .A(n3601), .ZN(n2375) );
  NAND2_X1 U3011 ( .A1(n2364), .A2(n2366), .ZN(n4080) );
  NAND2_X1 U3012 ( .A1(n3601), .A2(n2251), .ZN(n2364) );
  NAND3_X1 U3013 ( .A1(n2462), .A2(n2433), .A3(n2377), .ZN(n2482) );
  NAND4_X1 U3014 ( .A1(n2381), .A2(n2380), .A3(n2379), .A4(n2378), .ZN(n2405)
         );
  NAND2_X1 U3015 ( .A1(n2382), .A2(n2655), .ZN(n2725) );
  NAND2_X1 U3016 ( .A1(n4089), .A2(n2384), .ZN(n3105) );
  NAND3_X1 U3017 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .A3(
        IR_REG_31__SCAN_IN), .ZN(n2393) );
  NAND2_X1 U3018 ( .A1(n4940), .A2(n2254), .ZN(n2398) );
  NAND2_X1 U3019 ( .A1(n4940), .A2(n4942), .ZN(n4941) );
  INV_X1 U3020 ( .A(n2405), .ZN(n2403) );
  NAND2_X1 U3021 ( .A1(n2403), .A2(n2402), .ZN(n2756) );
  INV_X1 U3022 ( .A(n2588), .ZN(n2404) );
  NAND2_X1 U3023 ( .A1(n3032), .A2(n2252), .ZN(n2409) );
  AOI21_X1 U3024 ( .B1(n3032), .B2(n3031), .A(n3030), .ZN(n4043) );
  NAND2_X1 U3025 ( .A1(n3027), .A2(n2418), .ZN(n2417) );
  NOR2_X1 U3026 ( .A1(n4095), .A2(n4098), .ZN(n2426) );
  OAI21_X1 U3027 ( .B1(n4204), .B2(n2429), .A(n2427), .ZN(n3600) );
  NOR2_X2 U3028 ( .A1(n2434), .A2(IR_REG_22__SCAN_IN), .ZN(n2433) );
  NAND2_X1 U3029 ( .A1(n2438), .A2(n2250), .ZN(n3018) );
  NAND2_X1 U3030 ( .A1(n3013), .A2(n3012), .ZN(n3541) );
  NAND2_X1 U3031 ( .A1(n3163), .A2(n2440), .ZN(n3289) );
  NAND2_X1 U3032 ( .A1(n2494), .A2(n2441), .ZN(n2444) );
  XNOR2_X1 U3033 ( .A(n2518), .B(n2918), .ZN(n2535) );
  AOI22_X1 U3034 ( .A1(n3099), .A2(n3855), .B1(n2386), .B2(n4033), .ZN(n3038)
         );
  NAND2_X1 U3035 ( .A1(n3175), .A2(n4171), .ZN(n4173) );
  AND2_X2 U3036 ( .A1(n3093), .A2(n3174), .ZN(n5073) );
  AND2_X2 U3037 ( .A1(n3093), .A2(n3092), .ZN(n5081) );
  NAND2_X1 U3038 ( .A1(n3231), .A2(n2615), .ZN(n2445) );
  AND2_X1 U3039 ( .A1(n2640), .A2(n2639), .ZN(n2446) );
  OR2_X1 U3040 ( .A1(n5013), .A2(n3956), .ZN(n2447) );
  AND2_X1 U3041 ( .A1(n2785), .A2(REG0_REG_8__SCAN_IN), .ZN(n2448) );
  AND2_X1 U3042 ( .A1(n2220), .A2(REG1_REG_8__SCAN_IN), .ZN(n2449) );
  AND3_X1 U3043 ( .A1(n2523), .A2(n2522), .A3(n2521), .ZN(n2450) );
  AND2_X1 U3044 ( .A1(n3047), .A2(n3401), .ZN(n2451) );
  OR2_X1 U3045 ( .A1(n2455), .A2(n2875), .ZN(n2452) );
  AND3_X1 U3046 ( .A1(n2949), .A2(n2951), .A3(n4752), .ZN(n2453) );
  NAND2_X1 U3047 ( .A1(n2798), .A2(n3678), .ZN(n2799) );
  INV_X1 U3048 ( .A(n3851), .ZN(n4065) );
  NAND2_X1 U3049 ( .A1(n4734), .A2(n4217), .ZN(n2454) );
  NOR2_X1 U3050 ( .A1(n2865), .A2(n2864), .ZN(n2455) );
  AND2_X1 U3051 ( .A1(n2984), .A2(n2983), .ZN(n2456) );
  NAND2_X1 U3052 ( .A1(n3819), .A2(DATAI_26_), .ZN(n4055) );
  INV_X1 U3053 ( .A(n4055), .ZN(n3033) );
  AOI21_X1 U3054 ( .B1(n4080), .B2(n3887), .A(n3834), .ZN(n4063) );
  NOR2_X1 U3055 ( .A1(n3396), .A2(n2451), .ZN(n2457) );
  INV_X1 U3056 ( .A(n3964), .ZN(n5026) );
  INV_X1 U3057 ( .A(IR_REG_18__SCAN_IN), .ZN(n2463) );
  NAND2_X1 U3058 ( .A1(n3931), .A2(n2961), .ZN(n2566) );
  NAND2_X1 U3059 ( .A1(n2597), .A2(n2596), .ZN(n2615) );
  XNOR2_X1 U3060 ( .A(n2546), .B(n2918), .ZN(n2552) );
  INV_X1 U3061 ( .A(n3864), .ZN(n3019) );
  INV_X1 U3062 ( .A(n3924), .ZN(n3472) );
  INV_X1 U3063 ( .A(IR_REG_27__SCAN_IN), .ZN(n2492) );
  NAND2_X1 U3064 ( .A1(n2550), .A2(n2549), .ZN(n2553) );
  AND2_X1 U3065 ( .A1(REG3_REG_17__SCAN_IN), .A2(n2783), .ZN(n2801) );
  INV_X1 U3066 ( .A(n5033), .ZN(n3940) );
  NAND2_X1 U3067 ( .A1(n4869), .A2(n3946), .ZN(n4879) );
  NAND2_X1 U3068 ( .A1(n4065), .A2(n4055), .ZN(n3035) );
  AND2_X1 U3069 ( .A1(n4104), .A2(n3064), .ZN(n4098) );
  AND2_X1 U3070 ( .A1(n3602), .A2(n3603), .ZN(n4181) );
  NOR2_X1 U3071 ( .A1(n2649), .A2(n2648), .ZN(n2666) );
  OR2_X1 U3072 ( .A1(n3812), .A2(n3818), .ZN(n3855) );
  NOR2_X1 U3073 ( .A1(n2763), .A2(n4730), .ZN(n2783) );
  AOI21_X1 U3074 ( .B1(n2989), .B2(n2961), .A(n2526), .ZN(n2532) );
  INV_X1 U3075 ( .A(n4135), .ZN(n3720) );
  INV_X1 U3076 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3424) );
  INV_X1 U3077 ( .A(n3855), .ZN(n3098) );
  INV_X1 U3078 ( .A(n4098), .ZN(n4132) );
  AND4_X1 U3079 ( .A1(n2476), .A2(n2475), .A3(n2474), .A4(n2473), .ZN(n4158)
         );
  OR2_X1 U3080 ( .A1(n2637), .A2(n4628), .ZN(n2649) );
  AND2_X1 U3081 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2581) );
  INV_X1 U3082 ( .A(n3123), .ZN(n2940) );
  INV_X1 U3083 ( .A(n4217), .ZN(n3682) );
  INV_X1 U3084 ( .A(n3455), .ZN(n3461) );
  AND2_X1 U3085 ( .A1(n3046), .A2(n3772), .ZN(n3842) );
  NAND2_X1 U3086 ( .A1(n2952), .A2(n4752), .ZN(n2946) );
  INV_X1 U3087 ( .A(n4758), .ZN(n3723) );
  INV_X1 U3088 ( .A(n3699), .ZN(n4752) );
  AND2_X1 U3089 ( .A1(n2738), .A2(REG3_REG_14__SCAN_IN), .ZN(n2751) );
  NAND4_X1 U3090 ( .A1(n2891), .A2(n2890), .A3(n2889), .A4(n2888), .ZN(n3851)
         );
  NAND4_X1 U3091 ( .A1(n2855), .A2(n2854), .A3(n2853), .A4(n2852), .ZN(n4135)
         );
  AND4_X1 U3092 ( .A1(n2789), .A2(n2788), .A3(n2787), .A4(n2786), .ZN(n4189)
         );
  NAND2_X1 U3093 ( .A1(n4907), .A2(n4908), .ZN(n4906) );
  XNOR2_X1 U3094 ( .A(n3954), .B(n5015), .ZN(n4935) );
  AND2_X1 U3095 ( .A1(n4789), .A2(n3132), .ZN(n4211) );
  AND2_X1 U3096 ( .A1(n4173), .A2(n3252), .ZN(n4167) );
  INV_X1 U3097 ( .A(n4221), .ZN(n4991) );
  INV_X1 U3098 ( .A(n4171), .ZN(n4987) );
  AOI21_X1 U3099 ( .B1(n2940), .B2(n3127), .A(n2939), .ZN(n3092) );
  NAND2_X1 U3100 ( .A1(n3819), .A2(DATAI_23_), .ZN(n4115) );
  OR2_X1 U3101 ( .A1(n3349), .A2(n3845), .ZN(n5062) );
  NAND2_X1 U3102 ( .A1(n3527), .A2(n5065), .ZN(n4285) );
  AND3_X1 U3103 ( .A1(n3085), .A2(n3084), .A3(n3083), .ZN(n3093) );
  INV_X1 U3104 ( .A(n2932), .ZN(n3125) );
  AND2_X1 U3105 ( .A1(n2689), .A2(n2708), .ZN(n3964) );
  NAND2_X1 U3106 ( .A1(n2945), .A2(n2944), .ZN(n3699) );
  AND2_X1 U3107 ( .A1(n2962), .A2(n3150), .ZN(n4758) );
  NAND4_X1 U3108 ( .A1(n2903), .A2(n2902), .A3(n2901), .A4(n2900), .ZN(n4051)
         );
  NAND4_X1 U3109 ( .A1(n2818), .A2(n2817), .A3(n2816), .A4(n2815), .ZN(n4186)
         );
  INV_X1 U3110 ( .A(n4785), .ZN(n4960) );
  OR2_X1 U3111 ( .A1(n4199), .A2(n5047), .ZN(n4221) );
  OR2_X1 U3112 ( .A1(n4124), .A2(n4123), .ZN(n4257) );
  AND2_X1 U3113 ( .A1(n3509), .A2(n3508), .ZN(n4967) );
  INV_X1 U3114 ( .A(n4167), .ZN(n4225) );
  AND2_X1 U3115 ( .A1(n3095), .A2(n3094), .ZN(n3096) );
  NAND2_X1 U3116 ( .A1(n5081), .A2(n5070), .ZN(n4288) );
  NAND2_X1 U3117 ( .A1(n5073), .A2(n5070), .ZN(n4706) );
  INV_X1 U3118 ( .A(n5073), .ZN(n5071) );
  INV_X1 U3119 ( .A(n5007), .ZN(n5009) );
  NAND2_X1 U3120 ( .A1(n3124), .A2(n3123), .ZN(n5007) );
  OR2_X1 U3121 ( .A1(n2792), .A2(n2331), .ZN(n5014) );
  INV_X1 U3122 ( .A(n4835), .ZN(n5032) );
  AND2_X4 U3123 ( .A1(n2471), .A2(n2472), .ZN(n2785) );
  NAND2_X1 U3124 ( .A1(n2785), .A2(REG0_REG_21__SCAN_IN), .ZN(n2476) );
  NAND2_X1 U3125 ( .A1(n2221), .A2(REG1_REG_21__SCAN_IN), .ZN(n2475) );
  NAND2_X1 U3126 ( .A1(n2581), .A2(REG3_REG_5__SCAN_IN), .ZN(n2600) );
  NAND2_X1 U3127 ( .A1(n2618), .A2(REG3_REG_7__SCAN_IN), .ZN(n2637) );
  INV_X1 U3128 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2701) );
  INV_X1 U3129 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4730) );
  NAND2_X1 U3130 ( .A1(REG3_REG_19__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .ZN(
        n2469) );
  NAND2_X1 U3131 ( .A1(n2829), .A2(REG3_REG_21__SCAN_IN), .ZN(n2850) );
  OR2_X1 U3132 ( .A1(n2829), .A2(REG3_REG_21__SCAN_IN), .ZN(n2470) );
  AND2_X1 U3133 ( .A1(n2850), .A2(n2470), .ZN(n4153) );
  NAND2_X1 U3134 ( .A1(n2971), .A2(n4153), .ZN(n2474) );
  INV_X1 U3135 ( .A(n2471), .ZN(n3121) );
  NAND2_X1 U3136 ( .A1(n3137), .A2(REG2_REG_21__SCAN_IN), .ZN(n2473) );
  NAND2_X1 U3137 ( .A1(n2224), .A2(IR_REG_31__SCAN_IN), .ZN(n2942) );
  NAND2_X1 U3138 ( .A1(n2942), .A2(n2941), .ZN(n2479) );
  NAND2_X1 U3139 ( .A1(n2482), .A2(IR_REG_31__SCAN_IN), .ZN(n2483) );
  XNOR2_X1 U3140 ( .A(n2483), .B(n2376), .ZN(n4709) );
  INV_X1 U3141 ( .A(IR_REG_20__SCAN_IN), .ZN(n2487) );
  MUX2_X1 U3142 ( .A(IR_REG_31__SCAN_IN), .B(n2489), .S(IR_REG_21__SCAN_IN), 
        .Z(n2490) );
  AND2_X1 U3143 ( .A1(n2233), .A2(n2490), .ZN(n3905) );
  INV_X1 U3144 ( .A(n3176), .ZN(n2491) );
  NAND2_X1 U3145 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2497) );
  NAND2_X1 U3146 ( .A1(n2493), .A2(n2492), .ZN(n2496) );
  OAI22_X1 U3147 ( .A1(n4158), .A2(n2905), .B1(n2920), .B2(n4152), .ZN(n2503)
         );
  OR2_X1 U31480 ( .A1(n2499), .A2(n2498), .ZN(n2500) );
  NAND2_X1 U31490 ( .A1(n2233), .A2(IR_REG_31__SCAN_IN), .ZN(n2502) );
  NAND2_X1 U3150 ( .A1(n3998), .A2(n3913), .ZN(n2959) );
  XNOR2_X1 U3151 ( .A(n2503), .B(n2906), .ZN(n3656) );
  INV_X1 U3152 ( .A(n3913), .ZN(n2506) );
  INV_X1 U3153 ( .A(n3905), .ZN(n2505) );
  AND2_X2 U3154 ( .A1(n2504), .A2(n5039), .ZN(n5070) );
  OR2_X1 U3155 ( .A1(n4158), .A2(n2904), .ZN(n2508) );
  NAND2_X1 U3156 ( .A1(n3660), .A2(n2513), .ZN(n2507) );
  NAND2_X1 U3157 ( .A1(n2508), .A2(n2507), .ZN(n3657) );
  NAND2_X1 U3158 ( .A1(n2785), .A2(REG0_REG_1__SCAN_IN), .ZN(n2512) );
  NAND2_X1 U3159 ( .A1(n2583), .A2(REG1_REG_1__SCAN_IN), .ZN(n2511) );
  NAND2_X1 U3160 ( .A1(n2540), .A2(REG2_REG_1__SCAN_IN), .ZN(n2510) );
  NAND2_X1 U3161 ( .A1(n2222), .A2(REG3_REG_1__SCAN_IN), .ZN(n2509) );
  NAND4_X1 U3162 ( .A1(n2512), .A2(n2511), .A3(n2510), .A4(n2509), .ZN(n2988)
         );
  INV_X1 U3163 ( .A(n2513), .ZN(n2591) );
  NAND2_X1 U3164 ( .A1(n2988), .A2(n2513), .ZN(n2517) );
  INV_X1 U3165 ( .A(n2514), .ZN(n2515) );
  MUX2_X1 U3166 ( .A(n4774), .B(DATAI_1_), .S(n2525), .Z(n3178) );
  NAND2_X1 U3167 ( .A1(n3178), .A2(n2819), .ZN(n2516) );
  INV_X1 U3168 ( .A(n2988), .ZN(n2987) );
  OR2_X1 U3169 ( .A1(n2987), .A2(n2904), .ZN(n2520) );
  INV_X2 U3170 ( .A(n2591), .ZN(n2961) );
  NAND2_X1 U3171 ( .A1(n3178), .A2(n2961), .ZN(n2519) );
  NAND2_X1 U3172 ( .A1(n2520), .A2(n2519), .ZN(n2536) );
  XNOR2_X1 U3173 ( .A(n2535), .B(n2536), .ZN(n3187) );
  NAND2_X1 U3174 ( .A1(n2221), .A2(REG1_REG_0__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U3175 ( .A1(n2222), .A2(REG3_REG_0__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U3176 ( .A1(n2785), .A2(REG0_REG_0__SCAN_IN), .ZN(n2521) );
  NAND2_X2 U3177 ( .A1(n2524), .A2(n2450), .ZN(n2989) );
  MUX2_X1 U3178 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2525), .Z(n3179) );
  AND2_X1 U3179 ( .A1(n3179), .A2(n2819), .ZN(n2526) );
  INV_X1 U3180 ( .A(n3112), .ZN(n2527) );
  NAND2_X1 U3181 ( .A1(n2527), .A2(REG1_REG_0__SCAN_IN), .ZN(n2528) );
  NAND2_X1 U3182 ( .A1(n2532), .A2(n2528), .ZN(n3149) );
  NAND2_X1 U3183 ( .A1(n2989), .A2(n2915), .ZN(n2531) );
  NOR2_X1 U3184 ( .A1(n3112), .A2(n5038), .ZN(n2529) );
  AOI21_X1 U3185 ( .B1(n3179), .B2(n2961), .A(n2529), .ZN(n2530) );
  NAND2_X1 U3186 ( .A1(n2531), .A2(n2530), .ZN(n3148) );
  NAND2_X1 U3187 ( .A1(n3149), .A2(n3148), .ZN(n2534) );
  NAND2_X1 U3188 ( .A1(n2532), .A2(n2918), .ZN(n2533) );
  NAND2_X1 U3189 ( .A1(n3187), .A2(n3188), .ZN(n2539) );
  INV_X1 U3190 ( .A(n2535), .ZN(n2537) );
  NAND2_X1 U3191 ( .A1(n2537), .A2(n2536), .ZN(n2538) );
  NAND2_X1 U3192 ( .A1(n2540), .A2(REG2_REG_2__SCAN_IN), .ZN(n2545) );
  NAND2_X1 U3193 ( .A1(n2220), .A2(REG1_REG_2__SCAN_IN), .ZN(n2544) );
  NAND2_X1 U3194 ( .A1(n2222), .A2(REG3_REG_2__SCAN_IN), .ZN(n2543) );
  NAND2_X1 U3195 ( .A1(n2785), .A2(REG0_REG_2__SCAN_IN), .ZN(n2542) );
  INV_X1 U3196 ( .A(n2552), .ZN(n2550) );
  OR2_X1 U3197 ( .A1(n3162), .A2(n2904), .ZN(n2548) );
  NAND2_X1 U3198 ( .A1(n3294), .A2(n2961), .ZN(n2547) );
  AND2_X1 U3199 ( .A1(n2548), .A2(n2547), .ZN(n2551) );
  INV_X1 U3200 ( .A(n2551), .ZN(n2549) );
  NAND2_X1 U3201 ( .A1(n2552), .A2(n2551), .ZN(n2554) );
  AND2_X1 U3202 ( .A1(n2553), .A2(n2554), .ZN(n3156) );
  NAND2_X1 U3203 ( .A1(n3155), .A2(n2554), .ZN(n3196) );
  NAND2_X1 U3204 ( .A1(n2220), .A2(REG1_REG_3__SCAN_IN), .ZN(n2559) );
  NAND2_X1 U3205 ( .A1(n2785), .A2(REG0_REG_3__SCAN_IN), .ZN(n2557) );
  NAND2_X1 U3206 ( .A1(n2540), .A2(REG2_REG_3__SCAN_IN), .ZN(n2556) );
  INV_X1 U3207 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4981) );
  NAND2_X1 U3208 ( .A1(n2222), .A2(n4981), .ZN(n2555) );
  NOR3_X1 U3209 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .A3(
        IR_REG_2__SCAN_IN), .ZN(n2562) );
  INV_X1 U32100 ( .A(n2562), .ZN(n2560) );
  NAND2_X1 U32110 ( .A1(IR_REG_31__SCAN_IN), .A2(n2560), .ZN(n2561) );
  MUX2_X1 U32120 ( .A(n2561), .B(IR_REG_31__SCAN_IN), .S(n2563), .Z(n2564) );
  NAND2_X1 U32130 ( .A1(n2563), .A2(n2562), .ZN(n2577) );
  MUX2_X1 U32140 ( .A(n3967), .B(DATAI_3_), .S(n2525), .Z(n3274) );
  NAND2_X1 U32150 ( .A1(n3274), .A2(n2819), .ZN(n2565) );
  NAND2_X1 U32160 ( .A1(n2566), .A2(n2565), .ZN(n2567) );
  AND2_X1 U32170 ( .A1(n3274), .A2(n2961), .ZN(n2568) );
  AOI21_X1 U32180 ( .B1(n3931), .B2(n2915), .A(n2568), .ZN(n2570) );
  XNOR2_X1 U32190 ( .A(n2569), .B(n2570), .ZN(n3197) );
  NAND2_X1 U32200 ( .A1(n3196), .A2(n3197), .ZN(n3195) );
  INV_X1 U32210 ( .A(n2569), .ZN(n2571) );
  NAND2_X1 U32220 ( .A1(n2571), .A2(n2570), .ZN(n3242) );
  NAND2_X1 U32230 ( .A1(n2785), .A2(REG0_REG_4__SCAN_IN), .ZN(n2576) );
  NAND2_X1 U32240 ( .A1(n2221), .A2(REG1_REG_4__SCAN_IN), .ZN(n2575) );
  NOR2_X1 U32250 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2572) );
  NOR2_X1 U32260 ( .A1(n2581), .A2(n2572), .ZN(n3326) );
  NAND2_X1 U32270 ( .A1(n2222), .A2(n3326), .ZN(n2574) );
  NAND2_X1 U32280 ( .A1(n2540), .A2(REG2_REG_4__SCAN_IN), .ZN(n2573) );
  NAND2_X1 U32290 ( .A1(n2577), .A2(IR_REG_31__SCAN_IN), .ZN(n2578) );
  XNOR2_X1 U32300 ( .A(n2578), .B(IR_REG_4__SCAN_IN), .ZN(n4718) );
  MUX2_X1 U32310 ( .A(n4718), .B(DATAI_4_), .S(n2525), .Z(n3320) );
  OAI22_X1 U32320 ( .A1(n2580), .A2(n2905), .B1(n2920), .B2(n3315), .ZN(n2579)
         );
  XNOR2_X1 U32330 ( .A(n2579), .B(n2918), .ZN(n2612) );
  OAI22_X1 U32340 ( .A1(n2580), .A2(n2904), .B1(n2905), .B2(n3315), .ZN(n2613)
         );
  XNOR2_X1 U32350 ( .A(n2612), .B(n2613), .ZN(n3241) );
  AND2_X1 U32360 ( .A1(n3242), .A2(n3241), .ZN(n3230) );
  OAI21_X1 U32370 ( .B1(n2581), .B2(REG3_REG_5__SCAN_IN), .A(n2600), .ZN(n3255) );
  INV_X1 U32380 ( .A(n3255), .ZN(n2582) );
  NAND2_X1 U32390 ( .A1(n2222), .A2(n2582), .ZN(n2587) );
  NAND2_X1 U32400 ( .A1(n2221), .A2(REG1_REG_5__SCAN_IN), .ZN(n2586) );
  NAND2_X1 U32410 ( .A1(n2540), .A2(REG2_REG_5__SCAN_IN), .ZN(n2585) );
  NAND2_X1 U32420 ( .A1(n2785), .A2(REG0_REG_5__SCAN_IN), .ZN(n2584) );
  NAND2_X1 U32430 ( .A1(n2588), .A2(IR_REG_31__SCAN_IN), .ZN(n2589) );
  XNOR2_X1 U32440 ( .A(n2589), .B(IR_REG_5__SCAN_IN), .ZN(n5035) );
  INV_X1 U32450 ( .A(n5035), .ZN(n4823) );
  INV_X1 U32460 ( .A(DATAI_5_), .ZN(n2590) );
  MUX2_X1 U32470 ( .A(n4823), .B(n2590), .S(n2525), .Z(n3258) );
  OR2_X1 U32480 ( .A1(n2996), .A2(n2904), .ZN(n2594) );
  NAND2_X1 U32490 ( .A1(n3254), .A2(n2961), .ZN(n2593) );
  NAND2_X1 U32500 ( .A1(n2594), .A2(n2593), .ZN(n2596) );
  XNOR2_X1 U32510 ( .A(n2595), .B(n2596), .ZN(n3229) );
  INV_X1 U32520 ( .A(n3229), .ZN(n2598) );
  INV_X1 U32530 ( .A(n2595), .ZN(n2597) );
  NAND2_X1 U32540 ( .A1(n2598), .A2(n2615), .ZN(n2616) );
  AND2_X1 U32550 ( .A1(n3230), .A2(n2616), .ZN(n2599) );
  NAND2_X1 U32560 ( .A1(n3195), .A2(n2599), .ZN(n3210) );
  AND2_X1 U32570 ( .A1(n2600), .A2(n4415), .ZN(n2601) );
  NOR2_X1 U32580 ( .A1(n2618), .A2(n2601), .ZN(n4974) );
  NAND2_X1 U32590 ( .A1(n2971), .A2(n4974), .ZN(n2605) );
  NAND2_X1 U32600 ( .A1(n2221), .A2(REG1_REG_6__SCAN_IN), .ZN(n2604) );
  NAND2_X1 U32610 ( .A1(n3137), .A2(REG2_REG_6__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U32620 ( .A1(n2785), .A2(REG0_REG_6__SCAN_IN), .ZN(n2602) );
  NAND2_X1 U32630 ( .A1(n3928), .A2(n2961), .ZN(n2608) );
  OR2_X1 U32640 ( .A1(n2588), .A2(IR_REG_5__SCAN_IN), .ZN(n2657) );
  NAND2_X1 U32650 ( .A1(n2657), .A2(IR_REG_31__SCAN_IN), .ZN(n2606) );
  XNOR2_X1 U32660 ( .A(n2606), .B(IR_REG_6__SCAN_IN), .ZN(n5033) );
  MUX2_X1 U32670 ( .A(n5033), .B(DATAI_6_), .S(n2525), .Z(n3364) );
  NAND2_X1 U32680 ( .A1(n3364), .A2(n2819), .ZN(n2607) );
  NAND2_X1 U32690 ( .A1(n2608), .A2(n2607), .ZN(n2609) );
  NAND2_X1 U32700 ( .A1(n3928), .A2(n2915), .ZN(n2611) );
  NAND2_X1 U32710 ( .A1(n3364), .A2(n2961), .ZN(n2610) );
  NAND2_X1 U32720 ( .A1(n2611), .A2(n2610), .ZN(n2629) );
  NAND2_X1 U32730 ( .A1(n2628), .A2(n2629), .ZN(n3211) );
  INV_X1 U32740 ( .A(n2612), .ZN(n2614) );
  NAND2_X1 U32750 ( .A1(n2614), .A2(n2613), .ZN(n3231) );
  NAND2_X1 U32760 ( .A1(n2445), .A2(n2616), .ZN(n3209) );
  AND2_X1 U32770 ( .A1(n3211), .A2(n3209), .ZN(n2617) );
  NAND2_X1 U32780 ( .A1(n3210), .A2(n2617), .ZN(n3279) );
  NAND2_X1 U32790 ( .A1(n2785), .A2(REG0_REG_7__SCAN_IN), .ZN(n2623) );
  NAND2_X1 U32800 ( .A1(n2221), .A2(REG1_REG_7__SCAN_IN), .ZN(n2622) );
  OR2_X1 U32810 ( .A1(n2618), .A2(REG3_REG_7__SCAN_IN), .ZN(n2619) );
  AND2_X1 U32820 ( .A1(n2637), .A2(n2619), .ZN(n3284) );
  NAND2_X1 U32830 ( .A1(n2971), .A2(n3284), .ZN(n2621) );
  NAND2_X1 U32840 ( .A1(n2540), .A2(REG2_REG_7__SCAN_IN), .ZN(n2620) );
  OAI21_X1 U32850 ( .B1(n2657), .B2(IR_REG_6__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2624) );
  NAND2_X1 U32860 ( .A1(n2624), .A2(n2459), .ZN(n2642) );
  OR2_X1 U32870 ( .A1(n2624), .A2(n2459), .ZN(n2625) );
  MUX2_X1 U32880 ( .A(n4835), .B(DATAI_7_), .S(n2525), .Z(n3345) );
  INV_X1 U32890 ( .A(n3345), .ZN(n3340) );
  XNOR2_X1 U32900 ( .A(n2626), .B(n2906), .ZN(n2635) );
  OAI22_X1 U32910 ( .A1(n2627), .A2(n2904), .B1(n2905), .B2(n3340), .ZN(n2634)
         );
  XNOR2_X1 U32920 ( .A(n2635), .B(n2634), .ZN(n3283) );
  INV_X1 U32930 ( .A(n3283), .ZN(n2632) );
  INV_X1 U32940 ( .A(n2628), .ZN(n2631) );
  INV_X1 U32950 ( .A(n2629), .ZN(n2630) );
  NAND2_X1 U32960 ( .A1(n2631), .A2(n2630), .ZN(n3278) );
  AND2_X1 U32970 ( .A1(n2632), .A2(n3278), .ZN(n2633) );
  NAND2_X1 U32980 ( .A1(n2635), .A2(n2634), .ZN(n2636) );
  NAND2_X1 U32990 ( .A1(n2637), .A2(n4628), .ZN(n2638) );
  AND2_X1 U33000 ( .A1(n2649), .A2(n2638), .ZN(n4968) );
  NAND2_X1 U33010 ( .A1(n2971), .A2(n4968), .ZN(n2640) );
  NOR2_X1 U33020 ( .A1(n2448), .A2(n2449), .ZN(n2639) );
  NAND2_X1 U33030 ( .A1(n3137), .A2(REG2_REG_8__SCAN_IN), .ZN(n2641) );
  OR2_X1 U33040 ( .A1(n3341), .A2(n2904), .ZN(n2646) );
  NAND2_X1 U33050 ( .A1(n2642), .A2(IR_REG_31__SCAN_IN), .ZN(n2643) );
  XNOR2_X1 U33060 ( .A(n2643), .B(IR_REG_8__SCAN_IN), .ZN(n5029) );
  INV_X1 U33070 ( .A(DATAI_8_), .ZN(n2644) );
  MUX2_X1 U33080 ( .A(n4852), .B(n2644), .S(n2525), .Z(n3434) );
  INV_X1 U33090 ( .A(n3434), .ZN(n3444) );
  NAND2_X1 U33100 ( .A1(n3444), .A2(n2513), .ZN(n2645) );
  NAND2_X1 U33110 ( .A1(n2646), .A2(n2645), .ZN(n3222) );
  OAI22_X1 U33120 ( .A1(n3341), .A2(n2905), .B1(n2920), .B2(n3434), .ZN(n2647)
         );
  XNOR2_X1 U33130 ( .A(n2647), .B(n2906), .ZN(n3221) );
  AND2_X1 U33140 ( .A1(n2649), .A2(n2648), .ZN(n2650) );
  OR2_X1 U33150 ( .A1(n2650), .A2(n2666), .ZN(n3408) );
  INV_X1 U33160 ( .A(n3408), .ZN(n3336) );
  NAND2_X1 U33170 ( .A1(n2971), .A2(n3336), .ZN(n2654) );
  NAND2_X1 U33180 ( .A1(n2221), .A2(REG1_REG_9__SCAN_IN), .ZN(n2653) );
  NAND2_X1 U33190 ( .A1(n3137), .A2(REG2_REG_9__SCAN_IN), .ZN(n2652) );
  NAND2_X1 U33200 ( .A1(n2785), .A2(REG0_REG_9__SCAN_IN), .ZN(n2651) );
  NAND4_X1 U33210 ( .A1(n2654), .A2(n2653), .A3(n2652), .A4(n2651), .ZN(n3925)
         );
  NAND2_X1 U33220 ( .A1(n3925), .A2(n2961), .ZN(n2663) );
  NAND2_X1 U33230 ( .A1(n2655), .A2(n2459), .ZN(n2656) );
  NOR2_X1 U33240 ( .A1(n2657), .A2(n2656), .ZN(n2660) );
  NOR2_X1 U33250 ( .A1(n2660), .A2(n2964), .ZN(n2658) );
  MUX2_X1 U33260 ( .A(n2964), .B(n2658), .S(IR_REG_9__SCAN_IN), .Z(n2661) );
  INV_X1 U33270 ( .A(IR_REG_9__SCAN_IN), .ZN(n2659) );
  MUX2_X1 U33280 ( .A(n4856), .B(DATAI_9_), .S(n2525), .Z(n3405) );
  NAND2_X1 U33290 ( .A1(n3405), .A2(n2819), .ZN(n2662) );
  NAND2_X1 U33300 ( .A1(n2663), .A2(n2662), .ZN(n2664) );
  XNOR2_X1 U33310 ( .A(n2664), .B(n2918), .ZN(n2678) );
  AND2_X1 U33320 ( .A1(n3405), .A2(n2961), .ZN(n2665) );
  AOI21_X1 U33330 ( .B1(n3925), .B2(n2915), .A(n2665), .ZN(n2677) );
  XNOR2_X1 U33340 ( .A(n2678), .B(n2677), .ZN(n3332) );
  NOR2_X1 U33350 ( .A1(n2666), .A2(REG3_REG_10__SCAN_IN), .ZN(n2667) );
  OR2_X1 U33360 ( .A1(n2679), .A2(n2667), .ZN(n3641) );
  INV_X1 U33370 ( .A(n3641), .ZN(n4961) );
  NAND2_X1 U33380 ( .A1(n2971), .A2(n4961), .ZN(n2671) );
  NAND2_X1 U33390 ( .A1(n2221), .A2(REG1_REG_10__SCAN_IN), .ZN(n2670) );
  NAND2_X1 U33400 ( .A1(n3137), .A2(REG2_REG_10__SCAN_IN), .ZN(n2669) );
  NAND2_X1 U33410 ( .A1(n2785), .A2(REG0_REG_10__SCAN_IN), .ZN(n2668) );
  NAND4_X1 U33420 ( .A1(n2671), .A2(n2670), .A3(n2669), .A4(n2668), .ZN(n3924)
         );
  NAND2_X1 U33430 ( .A1(n3924), .A2(n2513), .ZN(n2674) );
  OR2_X1 U33440 ( .A1(n2685), .A2(n2964), .ZN(n2672) );
  XNOR2_X1 U33450 ( .A(n2672), .B(IR_REG_10__SCAN_IN), .ZN(n3979) );
  MUX2_X1 U33460 ( .A(n3979), .B(DATAI_10_), .S(n2525), .Z(n3639) );
  NAND2_X1 U33470 ( .A1(n3639), .A2(n2819), .ZN(n2673) );
  NAND2_X1 U33480 ( .A1(n2674), .A2(n2673), .ZN(n2675) );
  XNOR2_X1 U33490 ( .A(n2675), .B(n2906), .ZN(n2694) );
  AND2_X1 U33500 ( .A1(n3639), .A2(n2961), .ZN(n2676) );
  AOI21_X1 U33510 ( .B1(n3924), .B2(n2915), .A(n2676), .ZN(n2692) );
  XNOR2_X1 U33520 ( .A(n2694), .B(n2692), .ZN(n3637) );
  NAND2_X1 U3353 ( .A1(n2678), .A2(n2677), .ZN(n3635) );
  AND2_X1 U33540 ( .A1(n3637), .A2(n3635), .ZN(n3384) );
  NAND2_X1 U3355 ( .A1(n2785), .A2(REG0_REG_11__SCAN_IN), .ZN(n2684) );
  NAND2_X1 U3356 ( .A1(n2220), .A2(REG1_REG_11__SCAN_IN), .ZN(n2683) );
  OR2_X1 U3357 ( .A1(n2679), .A2(REG3_REG_11__SCAN_IN), .ZN(n2680) );
  AND2_X1 U3358 ( .A1(n2702), .A2(n2680), .ZN(n3390) );
  NAND2_X1 U3359 ( .A1(n2971), .A2(n3390), .ZN(n2682) );
  NAND2_X1 U3360 ( .A1(n3137), .A2(REG2_REG_11__SCAN_IN), .ZN(n2681) );
  INV_X1 U3361 ( .A(IR_REG_10__SCAN_IN), .ZN(n2722) );
  AOI21_X1 U3362 ( .B1(n2685), .B2(n2722), .A(n2964), .ZN(n2686) );
  NAND2_X1 U3363 ( .A1(n2686), .A2(IR_REG_11__SCAN_IN), .ZN(n2689) );
  INV_X1 U3364 ( .A(n2686), .ZN(n2688) );
  INV_X1 U3365 ( .A(IR_REG_11__SCAN_IN), .ZN(n2687) );
  NAND2_X1 U3366 ( .A1(n2688), .A2(n2687), .ZN(n2708) );
  MUX2_X1 U3367 ( .A(n3964), .B(DATAI_11_), .S(n2525), .Z(n3479) );
  OAI22_X1 U3368 ( .A1(n3505), .A2(n2905), .B1(n2920), .B2(n3086), .ZN(n2690)
         );
  XNOR2_X1 U3369 ( .A(n2690), .B(n2906), .ZN(n2696) );
  OAI22_X1 U3370 ( .A1(n3505), .A2(n2904), .B1(n2905), .B2(n3086), .ZN(n2695)
         );
  OR2_X1 U3371 ( .A1(n2696), .A2(n2695), .ZN(n3387) );
  AND2_X1 U3372 ( .A1(n3384), .A2(n3387), .ZN(n2691) );
  NAND2_X1 U3373 ( .A1(n3329), .A2(n2691), .ZN(n2700) );
  INV_X1 U3374 ( .A(n3387), .ZN(n2698) );
  INV_X1 U3375 ( .A(n2692), .ZN(n2693) );
  NAND2_X1 U3376 ( .A1(n2694), .A2(n2693), .ZN(n3385) );
  NAND2_X1 U3377 ( .A1(n2696), .A2(n2695), .ZN(n3386) );
  AND2_X1 U3378 ( .A1(n3385), .A2(n3386), .ZN(n2697) );
  OR2_X1 U3379 ( .A1(n2698), .A2(n2697), .ZN(n2699) );
  NAND2_X1 U3380 ( .A1(n2785), .A2(REG0_REG_12__SCAN_IN), .ZN(n2707) );
  NAND2_X1 U3381 ( .A1(n2220), .A2(REG1_REG_12__SCAN_IN), .ZN(n2706) );
  NAND2_X1 U3382 ( .A1(n2702), .A2(n2701), .ZN(n2703) );
  AND2_X1 U3383 ( .A1(n2717), .A2(n2703), .ZN(n3463) );
  NAND2_X1 U3384 ( .A1(n2971), .A2(n3463), .ZN(n2705) );
  NAND2_X1 U3385 ( .A1(n3137), .A2(REG2_REG_12__SCAN_IN), .ZN(n2704) );
  NAND4_X1 U3386 ( .A1(n2707), .A2(n2706), .A3(n2705), .A4(n2704), .ZN(n3553)
         );
  NAND2_X1 U3387 ( .A1(n3553), .A2(n2513), .ZN(n2711) );
  NAND2_X1 U3388 ( .A1(n2708), .A2(IR_REG_31__SCAN_IN), .ZN(n2709) );
  XNOR2_X1 U3389 ( .A(n2709), .B(IR_REG_12__SCAN_IN), .ZN(n5023) );
  MUX2_X1 U3390 ( .A(n5023), .B(DATAI_12_), .S(n2525), .Z(n3455) );
  NAND2_X1 U3391 ( .A1(n3455), .A2(n2819), .ZN(n2710) );
  NAND2_X1 U3392 ( .A1(n2711), .A2(n2710), .ZN(n2712) );
  XNOR2_X1 U3393 ( .A(n2712), .B(n2906), .ZN(n3376) );
  NAND2_X1 U3394 ( .A1(n3553), .A2(n2915), .ZN(n2714) );
  NAND2_X1 U3395 ( .A1(n3455), .A2(n2961), .ZN(n2713) );
  NAND2_X1 U3396 ( .A1(n2714), .A2(n2713), .ZN(n3375) );
  NAND2_X1 U3397 ( .A1(n3374), .A2(n3376), .ZN(n2715) );
  NAND2_X1 U3398 ( .A1(n2785), .A2(REG0_REG_13__SCAN_IN), .ZN(n2721) );
  NAND2_X1 U3399 ( .A1(n2221), .A2(REG1_REG_13__SCAN_IN), .ZN(n2720) );
  AOI21_X1 U3400 ( .B1(n2717), .B2(n3424), .A(n2738), .ZN(n3580) );
  NAND2_X1 U3401 ( .A1(n2971), .A2(n3580), .ZN(n2719) );
  NAND2_X1 U3402 ( .A1(n3137), .A2(REG2_REG_13__SCAN_IN), .ZN(n2718) );
  NAND2_X1 U3403 ( .A1(n3523), .A2(n2961), .ZN(n2730) );
  NAND2_X1 U3404 ( .A1(n2723), .A2(n2722), .ZN(n2724) );
  OR2_X1 U3405 ( .A1(n2725), .A2(n2724), .ZN(n2726) );
  OAI21_X1 U3406 ( .B1(n2727), .B2(n2726), .A(IR_REG_31__SCAN_IN), .ZN(n2728)
         );
  XNOR2_X1 U3407 ( .A(n2728), .B(IR_REG_13__SCAN_IN), .ZN(n4900) );
  MUX2_X1 U3408 ( .A(n4900), .B(DATAI_13_), .S(n3819), .Z(n3425) );
  NAND2_X1 U3409 ( .A1(n3425), .A2(n2819), .ZN(n2729) );
  NAND2_X1 U3410 ( .A1(n2730), .A2(n2729), .ZN(n2731) );
  XNOR2_X1 U3411 ( .A(n2731), .B(n2906), .ZN(n2734) );
  NAND2_X1 U3412 ( .A1(n3523), .A2(n2915), .ZN(n2733) );
  NAND2_X1 U3413 ( .A1(n3425), .A2(n2961), .ZN(n2732) );
  NAND2_X1 U3414 ( .A1(n2733), .A2(n2732), .ZN(n2735) );
  INV_X1 U3415 ( .A(n2734), .ZN(n2737) );
  INV_X1 U3416 ( .A(n2735), .ZN(n2736) );
  NAND2_X1 U3417 ( .A1(n2737), .A2(n2736), .ZN(n3419) );
  NAND2_X1 U3418 ( .A1(n2785), .A2(REG0_REG_14__SCAN_IN), .ZN(n2744) );
  NAND2_X1 U3419 ( .A1(n2220), .A2(REG1_REG_14__SCAN_IN), .ZN(n2743) );
  INV_X1 U3420 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2740) );
  INV_X1 U3421 ( .A(n2738), .ZN(n2739) );
  AOI21_X1 U3422 ( .B1(n2740), .B2(n2739), .A(n2751), .ZN(n3490) );
  NAND2_X1 U3423 ( .A1(n2971), .A2(n3490), .ZN(n2742) );
  NAND2_X1 U3424 ( .A1(n3137), .A2(REG2_REG_14__SCAN_IN), .ZN(n2741) );
  OR2_X1 U3425 ( .A1(n2745), .A2(n2964), .ZN(n2746) );
  XNOR2_X1 U3426 ( .A(n2746), .B(IR_REG_14__SCAN_IN), .ZN(n5019) );
  MUX2_X1 U3427 ( .A(n5019), .B(DATAI_14_), .S(n3819), .Z(n3531) );
  INV_X1 U3428 ( .A(n3531), .ZN(n3015) );
  OAI22_X1 U3429 ( .A1(n4745), .A2(n2904), .B1(n2905), .B2(n3015), .ZN(n3486)
         );
  AND2_X1 U3430 ( .A1(n3419), .A2(n3486), .ZN(n2747) );
  INV_X1 U3431 ( .A(n3486), .ZN(n2749) );
  OAI22_X1 U3432 ( .A1(n4745), .A2(n2905), .B1(n2920), .B2(n3015), .ZN(n2748)
         );
  XNOR2_X1 U3433 ( .A(n2748), .B(n2918), .ZN(n3487) );
  OR2_X1 U3434 ( .A1(n2749), .A2(n3487), .ZN(n2750) );
  OAI21_X1 U3435 ( .B1(REG3_REG_15__SCAN_IN), .B2(n2751), .A(n2763), .ZN(n4757) );
  INV_X1 U3436 ( .A(n4757), .ZN(n3574) );
  NAND2_X1 U3437 ( .A1(n2971), .A2(n3574), .ZN(n2755) );
  NAND2_X1 U3438 ( .A1(n2220), .A2(REG1_REG_15__SCAN_IN), .ZN(n2754) );
  NAND2_X1 U3439 ( .A1(n3137), .A2(REG2_REG_15__SCAN_IN), .ZN(n2753) );
  NAND2_X1 U3440 ( .A1(n2785), .A2(REG0_REG_15__SCAN_IN), .ZN(n2752) );
  NAND4_X1 U3441 ( .A1(n2755), .A2(n2754), .A3(n2753), .A4(n2752), .ZN(n3922)
         );
  NAND2_X1 U3442 ( .A1(n3922), .A2(n2961), .ZN(n2758) );
  NAND2_X1 U3443 ( .A1(n2756), .A2(IR_REG_31__SCAN_IN), .ZN(n2772) );
  XNOR2_X1 U3444 ( .A(n2772), .B(n2771), .ZN(n5018) );
  MUX2_X1 U3445 ( .A(n3988), .B(DATAI_15_), .S(n3819), .Z(n3571) );
  NAND2_X1 U3446 ( .A1(n3571), .A2(n2819), .ZN(n2757) );
  NAND2_X1 U3447 ( .A1(n2758), .A2(n2757), .ZN(n2759) );
  XNOR2_X1 U3448 ( .A(n2759), .B(n2906), .ZN(n2761) );
  AND2_X1 U3449 ( .A1(n3571), .A2(n2961), .ZN(n2760) );
  AOI21_X1 U3450 ( .B1(n3922), .B2(n2915), .A(n2760), .ZN(n4749) );
  NAND2_X1 U3451 ( .A1(n2762), .A2(n2761), .ZN(n4735) );
  INV_X1 U3452 ( .A(n2763), .ZN(n2765) );
  INV_X1 U3453 ( .A(n2783), .ZN(n2764) );
  OAI21_X1 U3454 ( .B1(REG3_REG_16__SCAN_IN), .B2(n2765), .A(n2764), .ZN(n4741) );
  INV_X1 U3455 ( .A(n4741), .ZN(n2766) );
  NAND2_X1 U3456 ( .A1(n2971), .A2(n2766), .ZN(n2770) );
  NAND2_X1 U3457 ( .A1(n2221), .A2(REG1_REG_16__SCAN_IN), .ZN(n2769) );
  NAND2_X1 U34580 ( .A1(n3137), .A2(REG2_REG_16__SCAN_IN), .ZN(n2768) );
  NAND2_X1 U34590 ( .A1(n2785), .A2(REG0_REG_16__SCAN_IN), .ZN(n2767) );
  NAND2_X1 U3460 ( .A1(n2772), .A2(n2771), .ZN(n2773) );
  NAND2_X1 U3461 ( .A1(n2773), .A2(IR_REG_31__SCAN_IN), .ZN(n2774) );
  XNOR2_X1 U3462 ( .A(n2774), .B(IR_REG_16__SCAN_IN), .ZN(n5015) );
  MUX2_X1 U3463 ( .A(n5015), .B(DATAI_16_), .S(n2525), .Z(n3021) );
  OAI22_X1 U3464 ( .A1(n3567), .A2(n2905), .B1(n2920), .B2(n4731), .ZN(n2775)
         );
  XNOR2_X1 U3465 ( .A(n2775), .B(n2918), .ZN(n2778) );
  OR2_X1 U3466 ( .A1(n3567), .A2(n2904), .ZN(n2777) );
  NAND2_X1 U34670 ( .A1(n3021), .A2(n2513), .ZN(n2776) );
  NAND2_X1 U3468 ( .A1(n2777), .A2(n2776), .ZN(n2779) );
  XNOR2_X1 U34690 ( .A(n2778), .B(n2779), .ZN(n4736) );
  NAND2_X1 U3470 ( .A1(n4735), .A2(n4736), .ZN(n2782) );
  NOR2_X1 U34710 ( .A1(REG3_REG_17__SCAN_IN), .A2(n2783), .ZN(n2784) );
  NOR2_X1 U3472 ( .A1(n2801), .A2(n2784), .ZN(n4219) );
  NAND2_X1 U34730 ( .A1(n2971), .A2(n4219), .ZN(n2789) );
  NAND2_X1 U3474 ( .A1(n2220), .A2(REG1_REG_17__SCAN_IN), .ZN(n2788) );
  NAND2_X1 U34750 ( .A1(n3137), .A2(REG2_REG_17__SCAN_IN), .ZN(n2787) );
  NAND2_X1 U3476 ( .A1(n2785), .A2(REG0_REG_17__SCAN_IN), .ZN(n2786) );
  NOR2_X1 U34770 ( .A1(n2790), .A2(n2964), .ZN(n2791) );
  MUX2_X1 U3478 ( .A(n2964), .B(n2791), .S(IR_REG_17__SCAN_IN), .Z(n2792) );
  INV_X1 U34790 ( .A(DATAI_17_), .ZN(n2793) );
  MUX2_X1 U3480 ( .A(n5014), .B(n2793), .S(n2525), .Z(n4217) );
  OAI22_X1 U34810 ( .A1(n4189), .A2(n2905), .B1(n2920), .B2(n4217), .ZN(n2794)
         );
  XNOR2_X1 U3482 ( .A(n2794), .B(n2918), .ZN(n3679) );
  OR2_X1 U34830 ( .A1(n4189), .A2(n2904), .ZN(n2796) );
  NAND2_X1 U3484 ( .A1(n3682), .A2(n2513), .ZN(n2795) );
  INV_X1 U34850 ( .A(n3679), .ZN(n2798) );
  INV_X1 U3486 ( .A(n2797), .ZN(n3678) );
  INV_X1 U34870 ( .A(n2800), .ZN(n3730) );
  NAND2_X1 U3488 ( .A1(n2785), .A2(REG0_REG_18__SCAN_IN), .ZN(n2805) );
  NAND2_X1 U34890 ( .A1(n2220), .A2(REG1_REG_18__SCAN_IN), .ZN(n2804) );
  OAI21_X1 U3490 ( .B1(n2801), .B2(REG3_REG_18__SCAN_IN), .A(n2827), .ZN(n3733) );
  INV_X1 U34910 ( .A(n3733), .ZN(n4197) );
  NAND2_X1 U3492 ( .A1(n2971), .A2(n4197), .ZN(n2803) );
  NAND2_X1 U34930 ( .A1(n3137), .A2(REG2_REG_18__SCAN_IN), .ZN(n2802) );
  NAND2_X1 U3494 ( .A1(n2806), .A2(IR_REG_31__SCAN_IN), .ZN(n2807) );
  XNOR2_X1 U34950 ( .A(n2807), .B(IR_REG_18__SCAN_IN), .ZN(n3991) );
  MUX2_X1 U3496 ( .A(n3991), .B(DATAI_18_), .S(n3819), .Z(n4193) );
  INV_X1 U34970 ( .A(n4193), .ZN(n3025) );
  OAI22_X1 U3498 ( .A1(n4209), .A2(n2905), .B1(n2920), .B2(n3025), .ZN(n2808)
         );
  XNOR2_X1 U34990 ( .A(n2808), .B(n2918), .ZN(n2814) );
  INV_X1 U3500 ( .A(n2814), .ZN(n2811) );
  OR2_X1 U35010 ( .A1(n4209), .A2(n2904), .ZN(n2810) );
  NAND2_X1 U3502 ( .A1(n4193), .A2(n2513), .ZN(n2809) );
  NAND2_X1 U35030 ( .A1(n2810), .A2(n2809), .ZN(n2812) );
  NAND2_X1 U3504 ( .A1(n2811), .A2(n2812), .ZN(n3726) );
  INV_X1 U35050 ( .A(n2812), .ZN(n2813) );
  AND2_X1 U35060 ( .A1(n2814), .A2(n2813), .ZN(n3727) );
  NAND2_X1 U35070 ( .A1(n2785), .A2(REG0_REG_19__SCAN_IN), .ZN(n2818) );
  NAND2_X1 U35080 ( .A1(n2221), .A2(REG1_REG_19__SCAN_IN), .ZN(n2817) );
  XNOR2_X1 U35090 ( .A(n2827), .B(REG3_REG_19__SCAN_IN), .ZN(n3653) );
  NAND2_X1 U35100 ( .A1(n2971), .A2(n3653), .ZN(n2816) );
  NAND2_X1 U35110 ( .A1(n3137), .A2(REG2_REG_19__SCAN_IN), .ZN(n2815) );
  MUX2_X1 U35120 ( .A(n4712), .B(DATAI_19_), .S(n3819), .Z(n3646) );
  AOI22_X1 U35130 ( .A1(n4186), .A2(n2915), .B1(n2961), .B2(n3646), .ZN(n2823)
         );
  NAND2_X1 U35140 ( .A1(n4186), .A2(n2513), .ZN(n2821) );
  NAND2_X1 U35150 ( .A1(n3646), .A2(n2819), .ZN(n2820) );
  NAND2_X1 U35160 ( .A1(n2821), .A2(n2820), .ZN(n2822) );
  XNOR2_X1 U35170 ( .A(n2822), .B(n2906), .ZN(n2825) );
  XOR2_X1 U35180 ( .A(n2823), .B(n2825), .Z(n3649) );
  INV_X1 U35190 ( .A(n2823), .ZN(n2824) );
  NAND2_X1 U35200 ( .A1(n2785), .A2(REG0_REG_20__SCAN_IN), .ZN(n2835) );
  NAND2_X1 U35210 ( .A1(n2220), .A2(REG1_REG_20__SCAN_IN), .ZN(n2834) );
  INV_X1 U35220 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4616) );
  INV_X1 U35230 ( .A(REG3_REG_20__SCAN_IN), .ZN(n2826) );
  OAI21_X1 U35240 ( .B1(n2827), .B2(n4616), .A(n2826), .ZN(n2828) );
  INV_X1 U35250 ( .A(n2828), .ZN(n2830) );
  OR2_X1 U35260 ( .A1(n2830), .A2(n2829), .ZN(n4172) );
  INV_X1 U35270 ( .A(n4172), .ZN(n2831) );
  NAND2_X1 U35280 ( .A1(n2971), .A2(n2831), .ZN(n2833) );
  NAND2_X1 U35290 ( .A1(n3137), .A2(REG2_REG_20__SCAN_IN), .ZN(n2832) );
  NAND4_X1 U35300 ( .A1(n2835), .A2(n2834), .A3(n2833), .A4(n2832), .ZN(n4148)
         );
  NAND2_X1 U35310 ( .A1(n4148), .A2(n2513), .ZN(n2837) );
  OR2_X1 U35320 ( .A1(n4168), .A2(n2920), .ZN(n2836) );
  NAND2_X1 U35330 ( .A1(n2837), .A2(n2836), .ZN(n2838) );
  XNOR2_X1 U35340 ( .A(n2838), .B(n2918), .ZN(n2841) );
  NOR2_X1 U35350 ( .A1(n4168), .A2(n2905), .ZN(n2839) );
  AOI21_X1 U35360 ( .B1(n4148), .B2(n2915), .A(n2839), .ZN(n2840) );
  OR2_X1 U35370 ( .A1(n2841), .A2(n2840), .ZN(n3702) );
  NAND2_X1 U35380 ( .A1(n2841), .A2(n2840), .ZN(n3701) );
  OAI21_X1 U35390 ( .B1(n3656), .B2(n3657), .A(n3701), .ZN(n2842) );
  AOI21_X1 U35400 ( .B1(n3703), .B2(n3702), .A(n2842), .ZN(n2843) );
  NAND2_X1 U35410 ( .A1(n2785), .A2(REG0_REG_22__SCAN_IN), .ZN(n2847) );
  NAND2_X1 U35420 ( .A1(n2221), .A2(REG1_REG_22__SCAN_IN), .ZN(n2846) );
  XNOR2_X1 U35430 ( .A(n2850), .B(REG3_REG_22__SCAN_IN), .ZN(n4127) );
  NAND2_X1 U35440 ( .A1(n2971), .A2(n4127), .ZN(n2845) );
  NAND2_X1 U35450 ( .A1(n3137), .A2(REG2_REG_22__SCAN_IN), .ZN(n2844) );
  INV_X1 U35460 ( .A(n4134), .ZN(n3718) );
  OAI22_X1 U35470 ( .A1(n4142), .A2(n2904), .B1(n2905), .B2(n3718), .ZN(n2859)
         );
  OAI22_X1 U35480 ( .A1(n4142), .A2(n2905), .B1(n2920), .B2(n3718), .ZN(n2848)
         );
  XNOR2_X1 U35490 ( .A(n2848), .B(n2906), .ZN(n2858) );
  XOR2_X1 U35500 ( .A(n2859), .B(n2858), .Z(n3715) );
  NAND2_X1 U35510 ( .A1(n2785), .A2(REG0_REG_23__SCAN_IN), .ZN(n2855) );
  NAND2_X1 U35520 ( .A1(n2220), .A2(REG1_REG_23__SCAN_IN), .ZN(n2854) );
  INV_X1 U35530 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3717) );
  INV_X1 U35540 ( .A(REG3_REG_23__SCAN_IN), .ZN(n2849) );
  OAI21_X1 U35550 ( .B1(n2850), .B2(n3717), .A(n2849), .ZN(n2851) );
  AND2_X1 U35560 ( .A1(n2851), .A2(n2866), .ZN(n3629) );
  NAND2_X1 U35570 ( .A1(n2971), .A2(n3629), .ZN(n2853) );
  NAND2_X1 U35580 ( .A1(n3137), .A2(REG2_REG_23__SCAN_IN), .ZN(n2852) );
  OAI22_X1 U35590 ( .A1(n3720), .A2(n2905), .B1(n2920), .B2(n4115), .ZN(n2856)
         );
  XNOR2_X1 U35600 ( .A(n2856), .B(n2906), .ZN(n2863) );
  NOR2_X1 U35610 ( .A1(n4115), .A2(n2905), .ZN(n2857) );
  AOI21_X1 U35620 ( .B1(n4135), .B2(n2915), .A(n2857), .ZN(n2864) );
  XNOR2_X1 U35630 ( .A(n2863), .B(n2864), .ZN(n3625) );
  INV_X1 U35640 ( .A(n2858), .ZN(n2861) );
  INV_X1 U35650 ( .A(n2859), .ZN(n2860) );
  NAND2_X1 U35660 ( .A1(n2861), .A2(n2860), .ZN(n3626) );
  INV_X1 U35670 ( .A(n2863), .ZN(n2865) );
  NAND2_X1 U35680 ( .A1(n2785), .A2(REG0_REG_24__SCAN_IN), .ZN(n2871) );
  NAND2_X1 U35690 ( .A1(n2221), .A2(REG1_REG_24__SCAN_IN), .ZN(n2870) );
  INV_X1 U35700 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4503) );
  AND2_X1 U35710 ( .A1(n2866), .A2(n4503), .ZN(n2867) );
  NOR2_X1 U35720 ( .A1(n2885), .A2(n2867), .ZN(n4090) );
  NAND2_X1 U35730 ( .A1(n2971), .A2(n4090), .ZN(n2869) );
  NAND2_X1 U35740 ( .A1(n3137), .A2(REG2_REG_24__SCAN_IN), .ZN(n2868) );
  NOR2_X1 U35750 ( .A1(n4087), .A2(n2905), .ZN(n2872) );
  AOI21_X1 U35760 ( .B1(n4110), .B2(n2915), .A(n2872), .ZN(n2874) );
  INV_X1 U35770 ( .A(n4110), .ZN(n3028) );
  OAI22_X1 U35780 ( .A1(n3028), .A2(n2905), .B1(n2920), .B2(n4087), .ZN(n2873)
         );
  XOR2_X1 U35790 ( .A(n2906), .B(n2873), .Z(n3692) );
  INV_X1 U35800 ( .A(n2874), .ZN(n2875) );
  OAI21_X2 U35810 ( .B1(n3628), .B2(n2455), .A(n2875), .ZN(n3690) );
  NAND2_X1 U3582 ( .A1(n2785), .A2(REG0_REG_25__SCAN_IN), .ZN(n2880) );
  NAND2_X1 U3583 ( .A1(n2221), .A2(REG1_REG_25__SCAN_IN), .ZN(n2879) );
  INV_X1 U3584 ( .A(REG3_REG_25__SCAN_IN), .ZN(n2876) );
  XNOR2_X1 U3585 ( .A(n2885), .B(n2876), .ZN(n4072) );
  NAND2_X1 U3586 ( .A1(n2971), .A2(n4072), .ZN(n2878) );
  NAND2_X1 U3587 ( .A1(n3137), .A2(REG2_REG_25__SCAN_IN), .ZN(n2877) );
  OAI22_X1 U3588 ( .A1(n4083), .A2(n2905), .B1(n2920), .B2(n4069), .ZN(n2881)
         );
  XNOR2_X1 U3589 ( .A(n2881), .B(n2906), .ZN(n2883) );
  OAI22_X1 U3590 ( .A1(n4083), .A2(n2904), .B1(n2905), .B2(n4069), .ZN(n2882)
         );
  OR2_X1 U3591 ( .A1(n2883), .A2(n2882), .ZN(n3667) );
  AND2_X1 U3592 ( .A1(n2883), .A2(n2882), .ZN(n3666) );
  NAND2_X1 U3593 ( .A1(n2785), .A2(REG0_REG_26__SCAN_IN), .ZN(n2891) );
  NAND2_X1 U3594 ( .A1(n2220), .A2(REG1_REG_26__SCAN_IN), .ZN(n2890) );
  AND2_X1 U3595 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2884) );
  AOI21_X1 U3596 ( .B1(n2885), .B2(REG3_REG_25__SCAN_IN), .A(
        REG3_REG_26__SCAN_IN), .ZN(n2886) );
  INV_X1 U3597 ( .A(n4057), .ZN(n2887) );
  NAND2_X1 U3598 ( .A1(n2971), .A2(n2887), .ZN(n2889) );
  NAND2_X1 U3599 ( .A1(n3137), .A2(REG2_REG_26__SCAN_IN), .ZN(n2888) );
  NAND2_X1 U3600 ( .A1(n3851), .A2(n2513), .ZN(n2893) );
  OR2_X1 U3601 ( .A1(n4055), .A2(n2920), .ZN(n2892) );
  NAND2_X1 U3602 ( .A1(n2893), .A2(n2892), .ZN(n2894) );
  XNOR2_X1 U3603 ( .A(n2894), .B(n2918), .ZN(n2897) );
  NOR2_X1 U3604 ( .A1(n4055), .A2(n2905), .ZN(n2895) );
  AOI21_X1 U3605 ( .B1(n3851), .B2(n2915), .A(n2895), .ZN(n2896) );
  AND2_X1 U3606 ( .A1(n2897), .A2(n2896), .ZN(n3737) );
  NAND2_X1 U3607 ( .A1(n2785), .A2(REG0_REG_27__SCAN_IN), .ZN(n2903) );
  NAND2_X1 U3608 ( .A1(n2220), .A2(REG1_REG_27__SCAN_IN), .ZN(n2902) );
  NOR2_X1 U3609 ( .A1(n2898), .A2(REG3_REG_27__SCAN_IN), .ZN(n2899) );
  NAND2_X1 U3610 ( .A1(n2971), .A2(n4038), .ZN(n2901) );
  NAND2_X1 U3611 ( .A1(n3137), .A2(REG2_REG_27__SCAN_IN), .ZN(n2900) );
  NAND2_X1 U3612 ( .A1(n3819), .A2(DATAI_27_), .ZN(n4031) );
  OAI22_X1 U3613 ( .A1(n3036), .A2(n2904), .B1(n4031), .B2(n2905), .ZN(n2947)
         );
  OAI22_X1 U3614 ( .A1(n3036), .A2(n2905), .B1(n4031), .B2(n2920), .ZN(n2907)
         );
  XNOR2_X1 U3615 ( .A(n2907), .B(n2906), .ZN(n2948) );
  XOR2_X1 U3616 ( .A(n2947), .B(n2948), .Z(n3617) );
  NAND2_X1 U3617 ( .A1(n2785), .A2(REG0_REG_28__SCAN_IN), .ZN(n2914) );
  NAND2_X1 U3618 ( .A1(n2221), .A2(REG1_REG_28__SCAN_IN), .ZN(n2913) );
  NAND2_X1 U3619 ( .A1(n2908), .A2(REG3_REG_28__SCAN_IN), .ZN(n4009) );
  INV_X1 U3620 ( .A(n2908), .ZN(n2909) );
  INV_X1 U3621 ( .A(REG3_REG_28__SCAN_IN), .ZN(n4504) );
  NAND2_X1 U3622 ( .A1(n2909), .A2(n4504), .ZN(n2910) );
  NAND2_X1 U3623 ( .A1(n2971), .A2(n4018), .ZN(n2912) );
  NAND2_X1 U3624 ( .A1(n3137), .A2(REG2_REG_28__SCAN_IN), .ZN(n2911) );
  NAND4_X1 U3625 ( .A1(n2914), .A2(n2913), .A3(n2912), .A4(n2911), .ZN(n4033)
         );
  NAND2_X1 U3626 ( .A1(n4033), .A2(n2915), .ZN(n2917) );
  NAND2_X1 U3627 ( .A1(n3819), .A2(DATAI_28_), .ZN(n3106) );
  NAND2_X1 U3628 ( .A1(n2386), .A2(n2513), .ZN(n2916) );
  NAND2_X1 U3629 ( .A1(n2917), .A2(n2916), .ZN(n2919) );
  XNOR2_X1 U3630 ( .A(n2919), .B(n2918), .ZN(n2923) );
  NOR2_X1 U3631 ( .A1(n3106), .A2(n2920), .ZN(n2921) );
  AOI21_X1 U3632 ( .B1(n4033), .B2(n2961), .A(n2921), .ZN(n2922) );
  XNOR2_X1 U3633 ( .A(n2923), .B(n2922), .ZN(n2952) );
  NOR4_X1 U3634 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2927) );
  NOR4_X1 U3635 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2926) );
  NOR4_X1 U3636 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2925) );
  NOR4_X1 U3637 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2924) );
  NAND4_X1 U3638 ( .A1(n2927), .A2(n2926), .A3(n2925), .A4(n2924), .ZN(n2937)
         );
  NOR2_X1 U3639 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_13__SCAN_IN), .ZN(n2931)
         );
  NOR4_X1 U3640 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2930) );
  NOR4_X1 U3641 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_22__SCAN_IN), .ZN(n2929) );
  NOR4_X1 U3642 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2928) );
  NAND4_X1 U3643 ( .A1(n2931), .A2(n2930), .A3(n2929), .A4(n2928), .ZN(n2936)
         );
  NAND2_X1 U3644 ( .A1(n2932), .A2(n4709), .ZN(n2933) );
  MUX2_X1 U3645 ( .A(n2932), .B(n2933), .S(B_REG_SCAN_IN), .Z(n2935) );
  OAI21_X1 U3646 ( .B1(n2937), .B2(n2936), .A(n2940), .ZN(n3083) );
  INV_X1 U3647 ( .A(n2934), .ZN(n2938) );
  NAND2_X1 U3648 ( .A1(n2938), .A2(n4709), .ZN(n3128) );
  AND2_X1 U3649 ( .A1(n3083), .A2(n3128), .ZN(n3173) );
  INV_X1 U3650 ( .A(D_REG_0__SCAN_IN), .ZN(n3127) );
  NOR2_X1 U3651 ( .A1(n2934), .A2(n3125), .ZN(n2939) );
  INV_X1 U3652 ( .A(D_REG_1__SCAN_IN), .ZN(n3169) );
  NAND2_X1 U3653 ( .A1(n2940), .A2(n3169), .ZN(n3080) );
  NAND3_X1 U3654 ( .A1(n3173), .A2(n3092), .A3(n3080), .ZN(n2979) );
  INV_X1 U3655 ( .A(n2979), .ZN(n2945) );
  XNOR2_X1 U3656 ( .A(n2942), .B(n2941), .ZN(n3131) );
  INV_X1 U3657 ( .A(n2504), .ZN(n4711) );
  AOI21_X1 U3658 ( .B1(n4712), .B2(n5039), .A(n3132), .ZN(n2943) );
  NAND2_X1 U3659 ( .A1(n4207), .A2(n2943), .ZN(n2954) );
  NOR2_X1 U3660 ( .A1(n3170), .A2(n2954), .ZN(n2944) );
  INV_X1 U3661 ( .A(n2952), .ZN(n2949) );
  NAND2_X1 U3662 ( .A1(n2948), .A2(n2947), .ZN(n2951) );
  NAND2_X1 U3663 ( .A1(n2950), .A2(n2453), .ZN(n2985) );
  INV_X1 U3664 ( .A(n2951), .ZN(n2953) );
  NAND3_X1 U3665 ( .A1(n2953), .A2(n4752), .A3(n2952), .ZN(n2984) );
  NAND2_X1 U3666 ( .A1(n2954), .A2(n4207), .ZN(n2955) );
  NAND2_X1 U3667 ( .A1(n2979), .A2(n2955), .ZN(n2957) );
  NAND2_X1 U3668 ( .A1(n2504), .A2(n3998), .ZN(n2956) );
  NAND2_X1 U3669 ( .A1(n2956), .A2(n3132), .ZN(n3172) );
  NAND2_X1 U3670 ( .A1(n2957), .A2(n3172), .ZN(n3151) );
  NAND2_X1 U3671 ( .A1(n3112), .A2(n3131), .ZN(n2958) );
  OAI21_X1 U3672 ( .B1(n3151), .B2(n2958), .A(STATE_REG_SCAN_IN), .ZN(n2962)
         );
  NOR2_X1 U3673 ( .A1(n5010), .A2(n2959), .ZN(n2960) );
  NAND2_X1 U3674 ( .A1(n2979), .A2(n3911), .ZN(n3150) );
  NOR2_X1 U3675 ( .A1(n2963), .A2(n2964), .ZN(n2965) );
  MUX2_X1 U3676 ( .A(n2964), .B(n2965), .S(IR_REG_28__SCAN_IN), .Z(n2966) );
  INV_X1 U3677 ( .A(n2966), .ZN(n2968) );
  NAND2_X1 U3678 ( .A1(n2968), .A2(n2967), .ZN(n3994) );
  NAND2_X1 U3679 ( .A1(n4789), .A2(n3911), .ZN(n2969) );
  NOR2_X2 U3680 ( .A1(n2979), .A2(n2969), .ZN(n3740) );
  INV_X1 U3681 ( .A(n3740), .ZN(n4744) );
  OAI22_X1 U3682 ( .A1(n4744), .A2(n3036), .B1(STATE_REG_SCAN_IN), .B2(n4504), 
        .ZN(n2982) );
  NAND2_X1 U3683 ( .A1(n2785), .A2(REG0_REG_29__SCAN_IN), .ZN(n2975) );
  NAND2_X1 U3684 ( .A1(n2220), .A2(REG1_REG_29__SCAN_IN), .ZN(n2974) );
  INV_X1 U3685 ( .A(n4009), .ZN(n2970) );
  NAND2_X1 U3686 ( .A1(n2971), .A2(n2970), .ZN(n2973) );
  NAND2_X1 U3687 ( .A1(n3137), .A2(REG2_REG_29__SCAN_IN), .ZN(n2972) );
  NAND4_X1 U3688 ( .A1(n2975), .A2(n2974), .A3(n2973), .A4(n2972), .ZN(n3918)
         );
  INV_X1 U3689 ( .A(n3918), .ZN(n2980) );
  NAND2_X1 U3690 ( .A1(n3994), .A2(n3911), .ZN(n2976) );
  INV_X1 U3691 ( .A(n2218), .ZN(n3719) );
  INV_X1 U3692 ( .A(n3170), .ZN(n3124) );
  NAND2_X1 U3693 ( .A1(n3124), .A2(n4231), .ZN(n2978) );
  NOR2_X1 U3694 ( .A1(n3998), .A2(n3913), .ZN(n2977) );
  NAND2_X1 U3695 ( .A1(n2504), .A2(n2977), .ZN(n5065) );
  OR2_X1 U3696 ( .A1(n5065), .A2(n3905), .ZN(n3081) );
  OAI21_X1 U3697 ( .B1(n2979), .B2(n2978), .A(n4171), .ZN(n3705) );
  OAI22_X1 U3698 ( .A1(n2980), .A2(n3719), .B1(n4743), .B2(n3106), .ZN(n2981)
         );
  AOI211_X1 U3699 ( .C1(n4018), .C2(n3723), .A(n2982), .B(n2981), .ZN(n2983)
         );
  NAND3_X1 U3700 ( .A1(n2986), .A2(n2985), .A3(n2456), .ZN(U3217) );
  AND2_X1 U3701 ( .A1(n2989), .A2(n3179), .ZN(n3164) );
  NAND2_X1 U3702 ( .A1(n2990), .A2(n3178), .ZN(n2991) );
  INV_X1 U3703 ( .A(n3162), .ZN(n3932) );
  NAND2_X1 U3704 ( .A1(n3932), .A2(n3301), .ZN(n3759) );
  NAND2_X1 U3705 ( .A1(n3162), .A2(n3294), .ZN(n3756) );
  NAND2_X1 U3706 ( .A1(n3759), .A2(n3756), .ZN(n3041) );
  NAND2_X1 U3707 ( .A1(n3162), .A2(n3301), .ZN(n2992) );
  NAND2_X1 U3708 ( .A1(n3289), .A2(n2992), .ZN(n3266) );
  NAND2_X1 U3709 ( .A1(n3931), .A2(n3274), .ZN(n2993) );
  NAND2_X1 U3710 ( .A1(n3266), .A2(n2993), .ZN(n2995) );
  INV_X1 U3711 ( .A(n3931), .ZN(n3296) );
  INV_X1 U3712 ( .A(n3274), .ZN(n3042) );
  NAND2_X1 U3713 ( .A1(n3296), .A2(n3042), .ZN(n2994) );
  NAND2_X1 U3714 ( .A1(n2995), .A2(n2994), .ZN(n3248) );
  NAND2_X1 U3715 ( .A1(n2580), .A2(n3320), .ZN(n3762) );
  NAND2_X1 U3716 ( .A1(n3930), .A2(n3315), .ZN(n3766) );
  AND2_X1 U3717 ( .A1(n2996), .A2(n3258), .ZN(n2999) );
  OR2_X1 U3718 ( .A1(n3844), .A2(n2999), .ZN(n3001) );
  NAND2_X1 U3719 ( .A1(n3930), .A2(n3320), .ZN(n3249) );
  INV_X1 U3720 ( .A(n2996), .ZN(n3929) );
  NAND2_X1 U3721 ( .A1(n3929), .A2(n3254), .ZN(n2997) );
  AND2_X1 U3722 ( .A1(n3249), .A2(n2997), .ZN(n2998) );
  OR2_X1 U3723 ( .A1(n2999), .A2(n2998), .ZN(n3000) );
  OAI21_X1 U3724 ( .B1(n3248), .B2(n3001), .A(n3000), .ZN(n3356) );
  AND2_X1 U3725 ( .A1(n3928), .A2(n3364), .ZN(n3002) );
  OAI22_X1 U3726 ( .A1(n3356), .A2(n3002), .B1(n3364), .B2(n3928), .ZN(n3349)
         );
  INV_X1 U3727 ( .A(n3349), .ZN(n3008) );
  NAND2_X1 U3728 ( .A1(n2627), .A2(n3345), .ZN(n3044) );
  NAND2_X1 U3729 ( .A1(n3927), .A2(n3340), .ZN(n3771) );
  AND2_X1 U3730 ( .A1(n3341), .A2(n3434), .ZN(n3005) );
  OR2_X1 U3731 ( .A1(n3845), .A2(n3005), .ZN(n3396) );
  INV_X1 U3732 ( .A(n3925), .ZN(n3047) );
  INV_X1 U3733 ( .A(n3405), .ZN(n3401) );
  NAND2_X1 U3734 ( .A1(n3927), .A2(n3345), .ZN(n3431) );
  NAND2_X1 U3735 ( .A1(n3926), .A2(n3444), .ZN(n3003) );
  AND2_X1 U3736 ( .A1(n3431), .A2(n3003), .ZN(n3004) );
  OR2_X1 U3737 ( .A1(n3005), .A2(n3004), .ZN(n3397) );
  AND2_X1 U3738 ( .A1(n2248), .A2(n3397), .ZN(n3006) );
  NOR2_X1 U3739 ( .A1(n2451), .A2(n3006), .ZN(n3007) );
  AOI21_X1 U3740 ( .B1(n3008), .B2(n2457), .A(n3007), .ZN(n3501) );
  NOR2_X1 U3741 ( .A1(n3924), .A2(n3639), .ZN(n3009) );
  INV_X1 U3742 ( .A(n3639), .ZN(n3498) );
  OAI22_X1 U3743 ( .A1(n3501), .A2(n3009), .B1(n3472), .B2(n3498), .ZN(n3467)
         );
  NAND2_X1 U3744 ( .A1(n3505), .A2(n3479), .ZN(n3453) );
  NAND2_X1 U3745 ( .A1(n3640), .A2(n3086), .ZN(n3790) );
  NAND2_X1 U3746 ( .A1(n3505), .A2(n3086), .ZN(n3010) );
  NAND2_X1 U3747 ( .A1(n3553), .A2(n3455), .ZN(n3011) );
  NAND2_X1 U3748 ( .A1(n3459), .A2(n3011), .ZN(n3013) );
  INV_X1 U3749 ( .A(n3553), .ZN(n3051) );
  NAND2_X1 U3750 ( .A1(n3051), .A2(n3461), .ZN(n3012) );
  NAND2_X1 U3751 ( .A1(n3523), .A2(n3425), .ZN(n3014) );
  NAND2_X1 U3752 ( .A1(n4745), .A2(n3531), .ZN(n3796) );
  NAND2_X1 U3753 ( .A1(n3923), .A2(n3015), .ZN(n3777) );
  NAND2_X1 U3754 ( .A1(n3922), .A2(n3571), .ZN(n3016) );
  NOR2_X1 U3755 ( .A1(n3923), .A2(n3531), .ZN(n3561) );
  INV_X1 U3756 ( .A(n3922), .ZN(n4732) );
  INV_X1 U3757 ( .A(n3571), .ZN(n4742) );
  AOI22_X1 U3758 ( .A1(n3561), .A2(n3016), .B1(n4732), .B2(n4742), .ZN(n3017)
         );
  NAND2_X1 U3759 ( .A1(n3018), .A2(n3017), .ZN(n3589) );
  INV_X1 U3760 ( .A(n3589), .ZN(n3020) );
  NAND2_X1 U3761 ( .A1(n3567), .A2(n3021), .ZN(n3876) );
  NAND2_X1 U3762 ( .A1(n4747), .A2(n4731), .ZN(n3878) );
  NAND2_X1 U3763 ( .A1(n3020), .A2(n3019), .ZN(n3587) );
  NAND2_X1 U3764 ( .A1(n4747), .A2(n3021), .ZN(n3022) );
  NAND2_X1 U3765 ( .A1(n3587), .A2(n3022), .ZN(n4204) );
  NAND2_X1 U3766 ( .A1(n4189), .A2(n4217), .ZN(n3023) );
  NAND2_X1 U3767 ( .A1(n4734), .A2(n3682), .ZN(n3024) );
  NAND2_X1 U3768 ( .A1(n4209), .A2(n4193), .ZN(n3602) );
  INV_X1 U3769 ( .A(n4209), .ZN(n3921) );
  NAND2_X1 U3770 ( .A1(n3921), .A2(n3025), .ZN(n3603) );
  NOR2_X1 U3771 ( .A1(n4186), .A2(n3646), .ZN(n4163) );
  INV_X1 U3772 ( .A(n4168), .ZN(n3706) );
  NAND2_X1 U3773 ( .A1(n4148), .A2(n3706), .ZN(n3836) );
  NAND2_X1 U3774 ( .A1(n4186), .A2(n3646), .ZN(n4164) );
  AND2_X1 U3775 ( .A1(n3836), .A2(n4164), .ZN(n3026) );
  OAI21_X1 U3776 ( .B1(n3600), .B2(n4163), .A(n3026), .ZN(n3027) );
  INV_X1 U3777 ( .A(n4148), .ZN(n3606) );
  NAND2_X1 U3778 ( .A1(n3606), .A2(n4168), .ZN(n3837) );
  NAND2_X1 U3779 ( .A1(n3707), .A2(n3660), .ZN(n4096) );
  NAND2_X1 U3780 ( .A1(n4142), .A2(n4134), .ZN(n4104) );
  INV_X1 U3781 ( .A(n4142), .ZN(n3920) );
  NAND2_X1 U3782 ( .A1(n3920), .A2(n3718), .ZN(n3064) );
  NOR2_X1 U3783 ( .A1(n3707), .A2(n3660), .ZN(n4095) );
  AND2_X1 U3784 ( .A1(n3920), .A2(n4134), .ZN(n4099) );
  NOR2_X1 U3785 ( .A1(n3028), .A2(n4087), .ZN(n3029) );
  INV_X1 U3786 ( .A(n4087), .ZN(n3694) );
  INV_X1 U3787 ( .A(n4062), .ZN(n3032) );
  NAND2_X1 U3788 ( .A1(n4083), .A2(n4069), .ZN(n3031) );
  INV_X1 U3789 ( .A(n4083), .ZN(n3919) );
  NOR2_X1 U3790 ( .A1(n4051), .A2(n4036), .ZN(n3037) );
  AND2_X1 U3791 ( .A1(n4033), .A2(n3106), .ZN(n3812) );
  NOR2_X1 U3792 ( .A1(n4033), .A2(n3106), .ZN(n3818) );
  NAND2_X1 U3793 ( .A1(n3819), .A2(DATAI_29_), .ZN(n3821) );
  XNOR2_X1 U3794 ( .A(n3918), .B(n3821), .ZN(n3866) );
  XNOR2_X1 U3795 ( .A(n3038), .B(n3866), .ZN(n4008) );
  XNOR2_X1 U3796 ( .A(n3176), .B(n3913), .ZN(n3039) );
  NAND2_X1 U3797 ( .A1(n3039), .A2(n3998), .ZN(n3527) );
  INV_X1 U3798 ( .A(n2989), .ZN(n3040) );
  NAND2_X1 U3799 ( .A1(n3040), .A2(n3179), .ZN(n3203) );
  NAND2_X1 U3800 ( .A1(n3296), .A2(n3274), .ZN(n3761) );
  NAND2_X1 U3801 ( .A1(n3931), .A2(n3042), .ZN(n3758) );
  AND2_X1 U3802 ( .A1(n3929), .A2(n3258), .ZN(n3764) );
  NAND2_X1 U3803 ( .A1(n2996), .A2(n3254), .ZN(n3781) );
  INV_X1 U3804 ( .A(n3364), .ZN(n3358) );
  NAND2_X1 U3805 ( .A1(n3928), .A2(n3358), .ZN(n3779) );
  NAND2_X1 U3806 ( .A1(n3357), .A2(n3779), .ZN(n3043) );
  INV_X1 U3807 ( .A(n3928), .ZN(n3259) );
  NAND2_X1 U3808 ( .A1(n3259), .A2(n3364), .ZN(n3768) );
  NAND2_X1 U3809 ( .A1(n3043), .A2(n3768), .ZN(n3339) );
  INV_X1 U3810 ( .A(n3044), .ZN(n3045) );
  OAI21_X1 U3811 ( .B1(n3339), .B2(n3045), .A(n3771), .ZN(n3433) );
  NAND2_X1 U3812 ( .A1(n3341), .A2(n3444), .ZN(n3773) );
  NAND2_X1 U3813 ( .A1(n3926), .A2(n3434), .ZN(n3770) );
  AND2_X1 U3814 ( .A1(n3925), .A2(n3401), .ZN(n3794) );
  INV_X1 U3815 ( .A(n3794), .ZN(n3046) );
  NAND2_X1 U3816 ( .A1(n3047), .A2(n3405), .ZN(n3772) );
  NAND2_X1 U3817 ( .A1(n3048), .A2(n3772), .ZN(n3503) );
  NAND2_X1 U3818 ( .A1(n3924), .A2(n3498), .ZN(n3789) );
  NAND2_X1 U3819 ( .A1(n3503), .A2(n3789), .ZN(n3049) );
  NAND2_X1 U3820 ( .A1(n3472), .A2(n3639), .ZN(n3793) );
  NAND2_X1 U3821 ( .A1(n3553), .A2(n3461), .ZN(n3546) );
  INV_X1 U3822 ( .A(n3425), .ZN(n3551) );
  NAND2_X1 U3823 ( .A1(n3523), .A2(n3551), .ZN(n3542) );
  NAND2_X1 U3824 ( .A1(n3546), .A2(n3542), .ZN(n3791) );
  INV_X1 U3825 ( .A(n3791), .ZN(n3050) );
  NAND2_X1 U3826 ( .A1(n3051), .A2(n3455), .ZN(n3545) );
  NAND2_X1 U3827 ( .A1(n3453), .A2(n3545), .ZN(n3052) );
  NOR2_X1 U3828 ( .A1(n3523), .A2(n3551), .ZN(n3543) );
  AOI21_X1 U3829 ( .B1(n3052), .B2(n3050), .A(n3543), .ZN(n3798) );
  NAND2_X1 U3830 ( .A1(n3053), .A2(n3798), .ZN(n3875) );
  NAND2_X1 U3831 ( .A1(n3875), .A2(n3865), .ZN(n3564) );
  NAND2_X1 U3832 ( .A1(n4732), .A2(n3571), .ZN(n3795) );
  NAND2_X1 U3833 ( .A1(n3922), .A2(n4742), .ZN(n3778) );
  NAND2_X1 U3834 ( .A1(n3795), .A2(n3778), .ZN(n3565) );
  INV_X1 U3835 ( .A(n3796), .ZN(n3054) );
  NOR2_X1 U3836 ( .A1(n3565), .A2(n3054), .ZN(n3055) );
  NAND2_X1 U3837 ( .A1(n3564), .A2(n3055), .ZN(n3056) );
  NAND2_X1 U3838 ( .A1(n3056), .A2(n3778), .ZN(n3590) );
  NAND2_X1 U3839 ( .A1(n3590), .A2(n3864), .ZN(n3057) );
  NAND2_X1 U3840 ( .A1(n3057), .A2(n3878), .ZN(n4206) );
  INV_X1 U3841 ( .A(n4206), .ZN(n3058) );
  NAND2_X1 U3842 ( .A1(n3058), .A2(n2454), .ZN(n3601) );
  NAND2_X1 U3843 ( .A1(n4186), .A2(n4169), .ZN(n3059) );
  NAND2_X1 U3844 ( .A1(n4189), .A2(n3682), .ZN(n3858) );
  NAND2_X1 U3845 ( .A1(n3602), .A2(n3858), .ZN(n3061) );
  NOR2_X1 U3846 ( .A1(n4186), .A2(n4169), .ZN(n3060) );
  AOI21_X1 U3847 ( .B1(n3061), .B2(n3879), .A(n3060), .ZN(n3749) );
  NOR2_X1 U3848 ( .A1(n4148), .A2(n4168), .ZN(n3750) );
  AND2_X1 U3849 ( .A1(n4148), .A2(n4168), .ZN(n3881) );
  INV_X1 U3850 ( .A(n3881), .ZN(n3062) );
  NAND2_X1 U3851 ( .A1(n4158), .A2(n3660), .ZN(n3854) );
  NAND2_X1 U3852 ( .A1(n4104), .A2(n3854), .ZN(n3886) );
  NOR2_X1 U3853 ( .A1(n4158), .A2(n3660), .ZN(n4101) );
  NAND2_X1 U3854 ( .A1(n4135), .A2(n4115), .ZN(n3063) );
  NAND2_X1 U3855 ( .A1(n3064), .A2(n3063), .ZN(n3807) );
  AOI21_X1 U3856 ( .B1(n4101), .B2(n4104), .A(n3807), .ZN(n3884) );
  NOR2_X1 U3857 ( .A1(n4110), .A2(n4087), .ZN(n3835) );
  NOR2_X1 U3858 ( .A1(n4135), .A2(n4115), .ZN(n4078) );
  NOR2_X1 U3859 ( .A1(n3835), .A2(n4078), .ZN(n3887) );
  AND2_X1 U3860 ( .A1(n4110), .A2(n4087), .ZN(n3834) );
  OR2_X1 U3861 ( .A1(n4083), .A2(n3671), .ZN(n3833) );
  NAND2_X1 U3862 ( .A1(n4063), .A2(n3833), .ZN(n4045) );
  NAND2_X1 U3863 ( .A1(n4083), .A2(n3671), .ZN(n4044) );
  NAND2_X1 U3864 ( .A1(n4065), .A2(n3033), .ZN(n3065) );
  NAND2_X1 U3865 ( .A1(n4044), .A2(n3065), .ZN(n3809) );
  INV_X1 U3866 ( .A(n3809), .ZN(n3897) );
  NAND2_X1 U3867 ( .A1(n3851), .A2(n4055), .ZN(n3893) );
  INV_X1 U3868 ( .A(n3893), .ZN(n3815) );
  AND2_X1 U3869 ( .A1(n4051), .A2(n4031), .ZN(n3816) );
  NOR2_X1 U3870 ( .A1(n4051), .A2(n4031), .ZN(n3817) );
  INV_X1 U3871 ( .A(n3812), .ZN(n3066) );
  XOR2_X1 U3872 ( .A(n3866), .B(n3067), .Z(n3079) );
  NAND2_X1 U3873 ( .A1(n4711), .A2(n3905), .ZN(n3069) );
  NAND2_X1 U3874 ( .A1(n4712), .A2(n3913), .ZN(n3068) );
  NAND2_X1 U3875 ( .A1(n4033), .A2(n4211), .ZN(n3077) );
  NAND2_X1 U3876 ( .A1(n2221), .A2(REG1_REG_30__SCAN_IN), .ZN(n3072) );
  NAND2_X1 U3877 ( .A1(n3137), .A2(REG2_REG_30__SCAN_IN), .ZN(n3071) );
  NAND2_X1 U3878 ( .A1(n2785), .A2(REG0_REG_30__SCAN_IN), .ZN(n3070) );
  NAND3_X1 U3879 ( .A1(n3072), .A2(n3071), .A3(n3070), .ZN(n3825) );
  XNOR2_X1 U3880 ( .A(n3073), .B(IR_REG_27__SCAN_IN), .ZN(n4787) );
  AND2_X1 U3881 ( .A1(n4787), .A2(B_REG_SCAN_IN), .ZN(n3074) );
  NOR2_X1 U3882 ( .A1(n4208), .A2(n3074), .ZN(n4003) );
  NOR2_X1 U3883 ( .A1(n3821), .A2(n4207), .ZN(n3075) );
  AOI21_X1 U3884 ( .B1(n3825), .B2(n4003), .A(n3075), .ZN(n3076) );
  AND2_X1 U3885 ( .A1(n3077), .A2(n3076), .ZN(n3078) );
  OAI21_X1 U3886 ( .B1(n3079), .B2(n4213), .A(n3078), .ZN(n4012) );
  AOI21_X1 U3887 ( .B1(n4008), .B2(n4285), .A(n4012), .ZN(n3097) );
  NAND2_X1 U3888 ( .A1(n3080), .A2(n3128), .ZN(n3085) );
  NAND2_X1 U3889 ( .A1(n3081), .A2(n3172), .ZN(n3082) );
  NOR2_X1 U3890 ( .A1(n3170), .A2(n3082), .ZN(n3084) );
  INV_X1 U3891 ( .A(n3092), .ZN(n3174) );
  NAND2_X1 U3892 ( .A1(n3316), .A2(n3315), .ZN(n3314) );
  NAND2_X1 U3893 ( .A1(n3440), .A2(n3434), .ZN(n3441) );
  OAI21_X1 U3894 ( .B1(n3088), .B2(n3821), .A(n4230), .ZN(n4010) );
  OR2_X1 U3895 ( .A1(n4010), .A2(n4706), .ZN(n3090) );
  NAND2_X1 U3896 ( .A1(n5071), .A2(REG0_REG_29__SCAN_IN), .ZN(n3089) );
  OAI21_X1 U3897 ( .B1(n3097), .B2(n5071), .A(n3091), .ZN(U3515) );
  NAND2_X1 U3898 ( .A1(n3451), .A2(REG1_REG_29__SCAN_IN), .ZN(n3094) );
  OAI21_X1 U3899 ( .B1(n3097), .B2(n3451), .A(n3096), .ZN(U3547) );
  INV_X1 U3900 ( .A(REG1_REG_28__SCAN_IN), .ZN(n3104) );
  AOI22_X1 U3901 ( .A1(n3918), .A2(n4185), .B1(n4231), .B2(n2386), .ZN(n3102)
         );
  NAND2_X1 U3902 ( .A1(n4051), .A2(n4211), .ZN(n3101) );
  OAI211_X1 U3903 ( .C1(n3103), .C2(n4213), .A(n3102), .B(n3101), .ZN(n4023)
         );
  AOI21_X1 U3904 ( .B1(n4016), .B2(n4285), .A(n4023), .ZN(n3109) );
  MUX2_X1 U3905 ( .A(n3104), .B(n3109), .S(n5081), .Z(n3108) );
  OAI21_X1 U3906 ( .B1(n2240), .B2(n3106), .A(n3105), .ZN(n4017) );
  NAND2_X1 U3907 ( .A1(n3108), .A2(n3107), .ZN(U3546) );
  INV_X1 U3908 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4549) );
  MUX2_X1 U3909 ( .A(n4549), .B(n3109), .S(n5073), .Z(n3111) );
  NAND2_X1 U3910 ( .A1(n3111), .A2(n3110), .ZN(U3514) );
  INV_X2 U3911 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3912 ( .A(DATAI_21_), .ZN(n3114) );
  NAND2_X1 U3913 ( .A1(n3905), .A2(STATE_REG_SCAN_IN), .ZN(n3113) );
  OAI21_X1 U3914 ( .B1(STATE_REG_SCAN_IN), .B2(n3114), .A(n3113), .ZN(U3331)
         );
  INV_X1 U3915 ( .A(DATAI_22_), .ZN(n4618) );
  NAND2_X1 U3916 ( .A1(n3913), .A2(STATE_REG_SCAN_IN), .ZN(n3115) );
  OAI21_X1 U3917 ( .B1(STATE_REG_SCAN_IN), .B2(n4618), .A(n3115), .ZN(U3330)
         );
  INV_X1 U3918 ( .A(DATAI_24_), .ZN(n3116) );
  MUX2_X1 U3919 ( .A(n3116), .B(n2932), .S(STATE_REG_SCAN_IN), .Z(n3117) );
  INV_X1 U3920 ( .A(n3117), .ZN(U3328) );
  INV_X1 U3921 ( .A(DATAI_29_), .ZN(n3120) );
  NAND2_X1 U3922 ( .A1(n3118), .A2(STATE_REG_SCAN_IN), .ZN(n3119) );
  OAI21_X1 U3923 ( .B1(STATE_REG_SCAN_IN), .B2(n3120), .A(n3119), .ZN(U3323)
         );
  INV_X1 U3924 ( .A(DATAI_30_), .ZN(n4362) );
  NAND2_X1 U3925 ( .A1(n3121), .A2(STATE_REG_SCAN_IN), .ZN(n3122) );
  OAI21_X1 U3926 ( .B1(STATE_REG_SCAN_IN), .B2(n4362), .A(n3122), .ZN(U3322)
         );
  NOR3_X1 U3927 ( .A1(n2934), .A2(n3125), .A3(n5010), .ZN(n3126) );
  AOI21_X1 U3928 ( .B1(n5007), .B2(n3127), .A(n3126), .ZN(U3458) );
  INV_X1 U3929 ( .A(n3128), .ZN(n3130) );
  AOI22_X1 U3930 ( .A1(n5007), .A2(n3169), .B1(n3130), .B2(n3129), .ZN(U3459)
         );
  OR2_X1 U3931 ( .A1(n3131), .A2(U3149), .ZN(n3916) );
  NAND2_X1 U3932 ( .A1(n3170), .A2(n3916), .ZN(n3961) );
  INV_X1 U3933 ( .A(n3961), .ZN(n3134) );
  NAND2_X1 U3934 ( .A1(n3132), .A2(n3131), .ZN(n3133) );
  NOR2_X2 U3935 ( .A1(n3134), .A2(n3962), .ZN(n4953) );
  NOR2_X1 U3936 ( .A1(n4953), .A2(U4043), .ZN(U3148) );
  INV_X1 U3937 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4630) );
  NAND2_X1 U3938 ( .A1(n3825), .A2(U4043), .ZN(n3135) );
  OAI21_X1 U3939 ( .B1(U4043), .B2(n4630), .A(n3135), .ZN(U3580) );
  INV_X1 U3940 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n4413) );
  NAND2_X1 U3941 ( .A1(n4135), .A2(U4043), .ZN(n3136) );
  OAI21_X1 U3942 ( .B1(U4043), .B2(n4413), .A(n3136), .ZN(U3573) );
  INV_X1 U3943 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n4416) );
  NAND2_X1 U3944 ( .A1(n2220), .A2(REG1_REG_31__SCAN_IN), .ZN(n3140) );
  NAND2_X1 U3945 ( .A1(n3137), .A2(REG2_REG_31__SCAN_IN), .ZN(n3139) );
  NAND2_X1 U3946 ( .A1(n2785), .A2(REG0_REG_31__SCAN_IN), .ZN(n3138) );
  NAND2_X1 U3947 ( .A1(n4004), .A2(U4043), .ZN(n3141) );
  OAI21_X1 U3948 ( .B1(U4043), .B2(n4416), .A(n3141), .ZN(U3581) );
  INV_X1 U3949 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n4608) );
  NAND2_X1 U3950 ( .A1(n2990), .A2(U4043), .ZN(n3142) );
  OAI21_X1 U3951 ( .B1(U4043), .B2(n4608), .A(n3142), .ZN(U3551) );
  INV_X1 U3952 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n4407) );
  NAND2_X1 U3953 ( .A1(n3553), .A2(U4043), .ZN(n3143) );
  OAI21_X1 U3954 ( .B1(U4043), .B2(n4407), .A(n3143), .ZN(U3562) );
  INV_X1 U3955 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n4603) );
  NAND2_X1 U3956 ( .A1(n3523), .A2(U4043), .ZN(n3144) );
  OAI21_X1 U3957 ( .B1(U4043), .B2(n4603), .A(n3144), .ZN(U3563) );
  INV_X1 U3958 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n4522) );
  NAND2_X1 U3959 ( .A1(n3707), .A2(U4043), .ZN(n3145) );
  OAI21_X1 U3960 ( .B1(U4043), .B2(n4522), .A(n3145), .ZN(U3571) );
  INV_X1 U3961 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n4625) );
  NAND2_X1 U3962 ( .A1(n3640), .A2(U4043), .ZN(n3146) );
  OAI21_X1 U3963 ( .B1(U4043), .B2(n4625), .A(n3146), .ZN(U3561) );
  INV_X1 U3964 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n4627) );
  NAND2_X1 U3965 ( .A1(n3851), .A2(U4043), .ZN(n3147) );
  OAI21_X1 U3966 ( .B1(U4043), .B2(n4627), .A(n3147), .ZN(U3576) );
  XNOR2_X1 U3967 ( .A(n3149), .B(n3148), .ZN(n4790) );
  INV_X1 U3968 ( .A(n3150), .ZN(n3152) );
  NOR3_X1 U3969 ( .A1(n3152), .A2(n3151), .A3(n3170), .ZN(n3161) );
  INV_X1 U3970 ( .A(n3161), .ZN(n3192) );
  OAI22_X1 U3971 ( .A1(n2987), .A2(n3719), .B1(n4743), .B2(n5040), .ZN(n3153)
         );
  AOI21_X1 U3972 ( .B1(n3192), .B2(REG3_REG_0__SCAN_IN), .A(n3153), .ZN(n3154)
         );
  OAI21_X1 U3973 ( .B1(n4790), .B2(n3699), .A(n3154), .ZN(U3229) );
  INV_X1 U3974 ( .A(REG3_REG_2__SCAN_IN), .ZN(n4533) );
  OAI21_X1 U3975 ( .B1(n2232), .B2(n3156), .A(n3155), .ZN(n3157) );
  NAND2_X1 U3976 ( .A1(n3157), .A2(n4752), .ZN(n3160) );
  OAI22_X1 U3977 ( .A1(n3296), .A2(n3719), .B1(n4744), .B2(n2987), .ZN(n3158)
         );
  AOI21_X1 U3978 ( .B1(n3294), .B2(n3741), .A(n3158), .ZN(n3159) );
  OAI211_X1 U3979 ( .C1(n3161), .C2(n4533), .A(n3160), .B(n3159), .ZN(U3234)
         );
  INV_X1 U3980 ( .A(n3203), .ZN(n3754) );
  XNOR2_X1 U3981 ( .A(n3859), .B(n3754), .ZN(n3168) );
  OAI22_X1 U3982 ( .A1(n3162), .A2(n4208), .B1(n4207), .B2(n3190), .ZN(n3166)
         );
  OAI21_X1 U3983 ( .B1(n3859), .B2(n3164), .A(n3163), .ZN(n5048) );
  NOR2_X1 U3984 ( .A1(n5048), .A2(n3527), .ZN(n3165) );
  AOI211_X1 U3985 ( .C1(n4211), .C2(n2989), .A(n3166), .B(n3165), .ZN(n3167)
         );
  OAI21_X1 U3986 ( .B1(n4213), .B2(n3168), .A(n3167), .ZN(n5050) );
  INV_X1 U3987 ( .A(n5050), .ZN(n3186) );
  OAI21_X1 U3988 ( .B1(n3170), .B2(n3169), .A(n5007), .ZN(n3171) );
  NAND4_X1 U3989 ( .A1(n3174), .A2(n3173), .A3(n3172), .A4(n3171), .ZN(n3175)
         );
  INV_X2 U3990 ( .A(n4173), .ZN(n4762) );
  INV_X1 U3991 ( .A(n5048), .ZN(n3184) );
  OR2_X1 U3992 ( .A1(n3176), .A2(n3998), .ZN(n3251) );
  INV_X1 U3993 ( .A(n3251), .ZN(n3177) );
  NAND2_X1 U3994 ( .A1(n4173), .A2(n3177), .ZN(n3485) );
  INV_X1 U3995 ( .A(n3485), .ZN(n4992) );
  NAND2_X1 U3996 ( .A1(n4173), .A2(n3998), .ZN(n4199) );
  INV_X1 U3997 ( .A(n3302), .ZN(n3181) );
  NAND2_X1 U3998 ( .A1(n3179), .A2(n3178), .ZN(n3180) );
  NAND2_X1 U3999 ( .A1(n3181), .A2(n3180), .ZN(n5046) );
  AOI22_X1 U4000 ( .A1(n4762), .A2(REG2_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(n4987), .ZN(n3182) );
  OAI21_X1 U4001 ( .B1(n4221), .B2(n5046), .A(n3182), .ZN(n3183) );
  AOI21_X1 U4002 ( .B1(n3184), .B2(n4992), .A(n3183), .ZN(n3185) );
  OAI21_X1 U4003 ( .B1(n3186), .B2(n4762), .A(n3185), .ZN(U3289) );
  XNOR2_X1 U4004 ( .A(n3188), .B(n3187), .ZN(n3194) );
  AOI22_X1 U4005 ( .A1(n3932), .A2(n2218), .B1(n3740), .B2(n2989), .ZN(n3189)
         );
  OAI21_X1 U4006 ( .B1(n4743), .B2(n3190), .A(n3189), .ZN(n3191) );
  AOI21_X1 U4007 ( .B1(REG3_REG_1__SCAN_IN), .B2(n3192), .A(n3191), .ZN(n3193)
         );
  OAI21_X1 U4008 ( .B1(n3194), .B2(n3699), .A(n3193), .ZN(U3219) );
  OAI21_X1 U4009 ( .B1(n3197), .B2(n3196), .A(n3195), .ZN(n3201) );
  AOI22_X1 U4010 ( .A1(n3932), .A2(n3740), .B1(n3274), .B2(n3741), .ZN(n3199)
         );
  NOR2_X1 U4011 ( .A1(STATE_REG_SCAN_IN), .A2(n4981), .ZN(n4724) );
  AOI21_X1 U4012 ( .B1(n3930), .B2(n2218), .A(n4724), .ZN(n3198) );
  OAI211_X1 U4013 ( .C1(REG3_REG_3__SCAN_IN), .C2(n4758), .A(n3199), .B(n3198), 
        .ZN(n3200) );
  AOI21_X1 U4014 ( .B1(n3201), .B2(n4752), .A(n3200), .ZN(n3202) );
  INV_X1 U4015 ( .A(n3202), .ZN(U3215) );
  NAND2_X1 U4016 ( .A1(n2989), .A2(n5040), .ZN(n3753) );
  AND2_X1 U4017 ( .A1(n3203), .A2(n3753), .ZN(n5042) );
  AND2_X1 U4018 ( .A1(n3527), .A2(n4213), .ZN(n3204) );
  OAI22_X1 U4019 ( .A1(n5042), .A2(n3204), .B1(n2987), .B2(n4208), .ZN(n5044)
         );
  AOI21_X1 U4020 ( .B1(n5039), .B2(n3998), .A(n4231), .ZN(n3205) );
  NOR2_X1 U4021 ( .A1(n5040), .A2(n3205), .ZN(n3206) );
  OAI21_X1 U4022 ( .B1(n5044), .B2(n3206), .A(n4223), .ZN(n3208) );
  AOI22_X1 U4023 ( .A1(n4762), .A2(REG2_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(n4987), .ZN(n3207) );
  OAI211_X1 U4024 ( .C1(n5042), .C2(n3485), .A(n3208), .B(n3207), .ZN(U3290)
         );
  NAND2_X1 U4025 ( .A1(n3210), .A2(n3209), .ZN(n3213) );
  NAND2_X1 U4026 ( .A1(n3211), .A2(n3278), .ZN(n3212) );
  XNOR2_X1 U4027 ( .A(n3213), .B(n3212), .ZN(n3218) );
  INV_X1 U4028 ( .A(n4974), .ZN(n3216) );
  AOI22_X1 U4029 ( .A1(n3929), .A2(n3740), .B1(n3364), .B2(n3705), .ZN(n3215)
         );
  NOR2_X1 U4030 ( .A1(STATE_REG_SCAN_IN), .A2(n4415), .ZN(n4828) );
  AOI21_X1 U4031 ( .B1(n3927), .B2(n2218), .A(n4828), .ZN(n3214) );
  OAI211_X1 U4032 ( .C1(n4758), .C2(n3216), .A(n3215), .B(n3214), .ZN(n3217)
         );
  AOI21_X1 U4033 ( .B1(n3218), .B2(n4752), .A(n3217), .ZN(n3219) );
  INV_X1 U4034 ( .A(n3219), .ZN(U3236) );
  XOR2_X1 U4035 ( .A(n3222), .B(n3221), .Z(n3223) );
  XNOR2_X1 U4036 ( .A(n3220), .B(n3223), .ZN(n3228) );
  NOR2_X1 U4037 ( .A1(STATE_REG_SCAN_IN), .A2(n4628), .ZN(n4854) );
  AOI21_X1 U4038 ( .B1(n2218), .B2(n3925), .A(n4854), .ZN(n3225) );
  NAND2_X1 U4039 ( .A1(n3705), .A2(n3444), .ZN(n3224) );
  OAI211_X1 U4040 ( .C1(n4744), .C2(n2627), .A(n3225), .B(n3224), .ZN(n3226)
         );
  AOI21_X1 U4041 ( .B1(n3723), .B2(n4968), .A(n3226), .ZN(n3227) );
  OAI21_X1 U4042 ( .B1(n3228), .B2(n3699), .A(n3227), .ZN(U3218) );
  NAND2_X1 U40430 ( .A1(n3195), .A2(n3230), .ZN(n3240) );
  NAND2_X1 U4044 ( .A1(n3240), .A2(n3231), .ZN(n3232) );
  XOR2_X1 U4045 ( .A(n3229), .B(n3232), .Z(n3236) );
  AOI22_X1 U4046 ( .A1(n3930), .A2(n3740), .B1(n3254), .B2(n3705), .ZN(n3234)
         );
  AND2_X1 U4047 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n4816) );
  AOI21_X1 U4048 ( .B1(n2218), .B2(n3928), .A(n4816), .ZN(n3233) );
  OAI211_X1 U4049 ( .C1(n4758), .C2(n3255), .A(n3234), .B(n3233), .ZN(n3235)
         );
  AOI21_X1 U4050 ( .B1(n3236), .B2(n4752), .A(n3235), .ZN(n3237) );
  INV_X1 U4051 ( .A(n3237), .ZN(U3224) );
  AOI22_X1 U4052 ( .A1(n3740), .A2(n3931), .B1(n3741), .B2(n3320), .ZN(n3239)
         );
  INV_X1 U4053 ( .A(REG3_REG_4__SCAN_IN), .ZN(n4553) );
  NOR2_X1 U4054 ( .A1(STATE_REG_SCAN_IN), .A2(n4553), .ZN(n4811) );
  INV_X1 U4055 ( .A(n4811), .ZN(n3238) );
  OAI211_X1 U4056 ( .C1(n2996), .C2(n3719), .A(n3239), .B(n3238), .ZN(n3246)
         );
  INV_X1 U4057 ( .A(n3240), .ZN(n3244) );
  AOI21_X1 U4058 ( .B1(n3195), .B2(n3242), .A(n3241), .ZN(n3243) );
  NOR3_X1 U4059 ( .A1(n3244), .A2(n3243), .A3(n3699), .ZN(n3245) );
  AOI211_X1 U4060 ( .C1(n3326), .C2(n3723), .A(n3246), .B(n3245), .ZN(n3247)
         );
  INV_X1 U4061 ( .A(n3247), .ZN(U3227) );
  XNOR2_X1 U4062 ( .A(n2996), .B(n3254), .ZN(n3853) );
  OR2_X1 U4063 ( .A1(n3248), .A2(n3844), .ZN(n3319) );
  NAND2_X1 U4064 ( .A1(n3319), .A2(n3249), .ZN(n3250) );
  XOR2_X1 U4065 ( .A(n3853), .B(n3250), .Z(n3309) );
  INV_X1 U4066 ( .A(n3309), .ZN(n3265) );
  NAND2_X1 U4067 ( .A1(n3527), .A2(n3251), .ZN(n3252) );
  INV_X1 U4068 ( .A(n3365), .ZN(n3253) );
  AOI21_X1 U4069 ( .B1(n3254), .B2(n3314), .A(n3253), .ZN(n3311) );
  INV_X1 U4070 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3966) );
  OAI22_X1 U4071 ( .A1(n3255), .A2(n4171), .B1(n3966), .B2(n4173), .ZN(n3256)
         );
  AOI21_X1 U4072 ( .B1(n3311), .B2(n4991), .A(n3256), .ZN(n3264) );
  XOR2_X1 U4073 ( .A(n3853), .B(n3257), .Z(n3262) );
  OAI22_X1 U4074 ( .A1(n3259), .A2(n4208), .B1(n4207), .B2(n3258), .ZN(n3260)
         );
  AOI21_X1 U4075 ( .B1(n4211), .B2(n3930), .A(n3260), .ZN(n3261) );
  OAI21_X1 U4076 ( .B1(n3262), .B2(n4213), .A(n3261), .ZN(n3308) );
  NAND2_X1 U4077 ( .A1(n3308), .A2(n4223), .ZN(n3263) );
  OAI211_X1 U4078 ( .C1(n3265), .C2(n4225), .A(n3264), .B(n3263), .ZN(U3285)
         );
  INV_X1 U4079 ( .A(n5065), .ZN(n5055) );
  XNOR2_X1 U4080 ( .A(n3266), .B(n3861), .ZN(n3269) );
  INV_X1 U4081 ( .A(n3269), .ZN(n4983) );
  XNOR2_X1 U4082 ( .A(n3267), .B(n3861), .ZN(n3272) );
  AOI22_X1 U4083 ( .A1(n3932), .A2(n4211), .B1(n4231), .B2(n3274), .ZN(n3268)
         );
  OAI21_X1 U4084 ( .B1(n2580), .B2(n4208), .A(n3268), .ZN(n3271) );
  NOR2_X1 U4085 ( .A1(n3269), .A2(n3527), .ZN(n3270) );
  AOI211_X1 U4086 ( .C1(n3272), .C2(n4183), .A(n3271), .B(n3270), .ZN(n4986)
         );
  INV_X1 U4087 ( .A(n4986), .ZN(n3273) );
  AOI21_X1 U4088 ( .B1(n5055), .B2(n4983), .A(n3273), .ZN(n3277) );
  AOI21_X1 U4089 ( .B1(n3274), .B2(n3300), .A(n3316), .ZN(n4982) );
  INV_X1 U4090 ( .A(n4706), .ZN(n3447) );
  AOI22_X1 U4091 ( .A1(n4982), .A2(n3447), .B1(REG0_REG_3__SCAN_IN), .B2(n5071), .ZN(n3275) );
  OAI21_X1 U4092 ( .B1(n3277), .B2(n5071), .A(n3275), .ZN(U3473) );
  INV_X1 U4093 ( .A(n4288), .ZN(n3449) );
  AOI22_X1 U4094 ( .A1(n4982), .A2(n3449), .B1(REG1_REG_3__SCAN_IN), .B2(n3451), .ZN(n3276) );
  OAI21_X1 U4095 ( .B1(n3277), .B2(n3451), .A(n3276), .ZN(U3521) );
  NAND2_X1 U4096 ( .A1(n3279), .A2(n3278), .ZN(n3282) );
  INV_X1 U4097 ( .A(n3280), .ZN(n3281) );
  AOI211_X1 U4098 ( .C1(n3283), .C2(n3282), .A(n3699), .B(n3281), .ZN(n3288)
         );
  INV_X1 U4099 ( .A(n3284), .ZN(n3348) );
  AOI22_X1 U4100 ( .A1(n3926), .A2(n2218), .B1(n3345), .B2(n3705), .ZN(n3286)
         );
  INV_X1 U4101 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4371) );
  NOR2_X1 U4102 ( .A1(STATE_REG_SCAN_IN), .A2(n4371), .ZN(n4840) );
  AOI21_X1 U4103 ( .B1(n3740), .B2(n3928), .A(n4840), .ZN(n3285) );
  OAI211_X1 U4104 ( .C1(n4758), .C2(n3348), .A(n3286), .B(n3285), .ZN(n3287)
         );
  OR2_X1 U4105 ( .A1(n3288), .A2(n3287), .ZN(U3210) );
  INV_X1 U4106 ( .A(n3289), .ZN(n3290) );
  AOI21_X1 U4107 ( .B1(n3843), .B2(n3291), .A(n3290), .ZN(n4988) );
  OAI21_X1 U4108 ( .B1(n3843), .B2(n3293), .A(n3292), .ZN(n3299) );
  AOI22_X1 U4109 ( .A1(n2990), .A2(n4211), .B1(n4231), .B2(n3294), .ZN(n3295)
         );
  OAI21_X1 U4110 ( .B1(n3296), .B2(n4208), .A(n3295), .ZN(n3298) );
  NOR2_X1 U4111 ( .A1(n4988), .A2(n3527), .ZN(n3297) );
  AOI211_X1 U4112 ( .C1(n4183), .C2(n3299), .A(n3298), .B(n3297), .ZN(n4996)
         );
  OAI21_X1 U4113 ( .B1(n4988), .B2(n5065), .A(n4996), .ZN(n3306) );
  OAI21_X1 U4114 ( .B1(n3302), .B2(n3301), .A(n3300), .ZN(n4989) );
  INV_X1 U4115 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4493) );
  OAI22_X1 U4116 ( .A1(n4288), .A2(n4989), .B1(n5081), .B2(n4493), .ZN(n3303)
         );
  AOI21_X1 U4117 ( .B1(n3306), .B2(n5081), .A(n3303), .ZN(n3304) );
  INV_X1 U4118 ( .A(n3304), .ZN(U3520) );
  INV_X1 U4119 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4632) );
  OAI22_X1 U4120 ( .A1(n4706), .A2(n4989), .B1(n5073), .B2(n4632), .ZN(n3305)
         );
  AOI21_X1 U4121 ( .B1(n3306), .B2(n5073), .A(n3305), .ZN(n3307) );
  INV_X1 U4122 ( .A(n3307), .ZN(U3471) );
  AOI21_X1 U4123 ( .B1(n3309), .B2(n4285), .A(n3308), .ZN(n3313) );
  AOI22_X1 U4124 ( .A1(n3311), .A2(n3447), .B1(REG0_REG_5__SCAN_IN), .B2(n5071), .ZN(n3310) );
  OAI21_X1 U4125 ( .B1(n3313), .B2(n5071), .A(n3310), .ZN(U3477) );
  AOI22_X1 U4126 ( .A1(n3311), .A2(n3449), .B1(REG1_REG_5__SCAN_IN), .B2(n3451), .ZN(n3312) );
  OAI21_X1 U4127 ( .B1(n3313), .B2(n3451), .A(n3312), .ZN(U3523) );
  OAI211_X1 U4128 ( .C1(n3316), .C2(n3315), .A(n3314), .B(n5070), .ZN(n5052)
         );
  NOR2_X1 U4129 ( .A1(n5052), .A2(n4712), .ZN(n3325) );
  XOR2_X1 U4130 ( .A(n3844), .B(n3317), .Z(n3324) );
  NAND2_X1 U4131 ( .A1(n3248), .A2(n3844), .ZN(n3318) );
  AND2_X1 U4132 ( .A1(n3319), .A2(n3318), .ZN(n5056) );
  INV_X1 U4133 ( .A(n3527), .ZN(n3502) );
  AOI22_X1 U4134 ( .A1(n3931), .A2(n4211), .B1(n4231), .B2(n3320), .ZN(n3321)
         );
  OAI21_X1 U4135 ( .B1(n2996), .B2(n4208), .A(n3321), .ZN(n3322) );
  AOI21_X1 U4136 ( .B1(n5056), .B2(n3502), .A(n3322), .ZN(n3323) );
  OAI21_X1 U4137 ( .B1(n4213), .B2(n3324), .A(n3323), .ZN(n5053) );
  AOI211_X1 U4138 ( .C1(n4987), .C2(n3326), .A(n3325), .B(n5053), .ZN(n3328)
         );
  AOI22_X1 U4139 ( .A1(n5056), .A2(n4992), .B1(REG2_REG_4__SCAN_IN), .B2(n4762), .ZN(n3327) );
  OAI21_X1 U4140 ( .B1(n3328), .B2(n4762), .A(n3327), .ZN(U3286) );
  INV_X1 U4141 ( .A(n3329), .ZN(n3330) );
  AOI21_X1 U4142 ( .B1(n3332), .B2(n3331), .A(n3330), .ZN(n3338) );
  AND2_X1 U4143 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4867) );
  AOI21_X1 U4144 ( .B1(n2218), .B2(n3924), .A(n4867), .ZN(n3334) );
  NAND2_X1 U4145 ( .A1(n3705), .A2(n3405), .ZN(n3333) );
  OAI211_X1 U4146 ( .C1(n4744), .C2(n3341), .A(n3334), .B(n3333), .ZN(n3335)
         );
  AOI21_X1 U4147 ( .B1(n3723), .B2(n3336), .A(n3335), .ZN(n3337) );
  OAI21_X1 U4148 ( .B1(n3338), .B2(n3699), .A(n3337), .ZN(U3228) );
  XOR2_X1 U4149 ( .A(n3845), .B(n3339), .Z(n3344) );
  OAI22_X1 U4150 ( .A1(n3341), .A2(n4208), .B1(n4207), .B2(n3340), .ZN(n3342)
         );
  AOI21_X1 U4151 ( .B1(n4211), .B2(n3928), .A(n3342), .ZN(n3343) );
  OAI21_X1 U4152 ( .B1(n3344), .B2(n4213), .A(n3343), .ZN(n5060) );
  INV_X1 U4153 ( .A(n5060), .ZN(n3355) );
  INV_X1 U4154 ( .A(n4199), .ZN(n3353) );
  NAND2_X1 U4155 ( .A1(n3367), .A2(n3345), .ZN(n3346) );
  NAND2_X1 U4156 ( .A1(n3346), .A2(n5070), .ZN(n3347) );
  NOR2_X1 U4157 ( .A1(n3440), .A2(n3347), .ZN(n5061) );
  INV_X1 U4158 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3965) );
  OAI22_X1 U4159 ( .A1(n4173), .A2(n3965), .B1(n3348), .B2(n4171), .ZN(n3352)
         );
  INV_X1 U4160 ( .A(n5062), .ZN(n3350) );
  AND2_X1 U4161 ( .A1(n3349), .A2(n3845), .ZN(n5059) );
  NOR3_X1 U4162 ( .A1(n3350), .A2(n5059), .A3(n4225), .ZN(n3351) );
  AOI211_X1 U4163 ( .C1(n3353), .C2(n5061), .A(n3352), .B(n3351), .ZN(n3354)
         );
  OAI21_X1 U4164 ( .B1(n4762), .B2(n3355), .A(n3354), .ZN(U3283) );
  AND2_X1 U4165 ( .A1(n3779), .A2(n3768), .ZN(n3863) );
  XNOR2_X1 U4166 ( .A(n3356), .B(n3863), .ZN(n4977) );
  INV_X1 U4167 ( .A(n4977), .ZN(n3363) );
  XOR2_X1 U4168 ( .A(n3863), .B(n3357), .Z(n3361) );
  OAI22_X1 U4169 ( .A1(n2996), .A2(n4188), .B1(n4207), .B2(n3358), .ZN(n3359)
         );
  AOI21_X1 U4170 ( .B1(n4185), .B2(n3927), .A(n3359), .ZN(n3360) );
  OAI21_X1 U4171 ( .B1(n3361), .B2(n4213), .A(n3360), .ZN(n3362) );
  AOI21_X1 U4172 ( .B1(n3502), .B2(n4977), .A(n3362), .ZN(n4980) );
  OAI21_X1 U4173 ( .B1(n5065), .B2(n3363), .A(n4980), .ZN(n3372) );
  NAND2_X1 U4174 ( .A1(n3365), .A2(n3364), .ZN(n3366) );
  NAND2_X1 U4175 ( .A1(n3367), .A2(n3366), .ZN(n4975) );
  INV_X1 U4176 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3368) );
  OAI22_X1 U4177 ( .A1(n4975), .A2(n4706), .B1(n5073), .B2(n3368), .ZN(n3369)
         );
  AOI21_X1 U4178 ( .B1(n3372), .B2(n5073), .A(n3369), .ZN(n3370) );
  INV_X1 U4179 ( .A(n3370), .ZN(U3479) );
  INV_X1 U4180 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4827) );
  OAI22_X1 U4181 ( .A1(n4975), .A2(n4288), .B1(n5081), .B2(n4827), .ZN(n3371)
         );
  AOI21_X1 U4182 ( .B1(n3372), .B2(n5081), .A(n3371), .ZN(n3373) );
  INV_X1 U4183 ( .A(n3373), .ZN(U3524) );
  XNOR2_X1 U4184 ( .A(n3376), .B(n3375), .ZN(n3377) );
  XNOR2_X1 U4185 ( .A(n3374), .B(n3377), .ZN(n3382) );
  INV_X1 U4186 ( .A(n3463), .ZN(n3380) );
  NOR2_X1 U4187 ( .A1(STATE_REG_SCAN_IN), .A2(n2701), .ZN(n4897) );
  AOI21_X1 U4188 ( .B1(n3640), .B2(n3740), .A(n4897), .ZN(n3379) );
  AOI22_X1 U4189 ( .A1(n2218), .A2(n3523), .B1(n3741), .B2(n3455), .ZN(n3378)
         );
  OAI211_X1 U4190 ( .C1(n4758), .C2(n3380), .A(n3379), .B(n3378), .ZN(n3381)
         );
  AOI21_X1 U4191 ( .B1(n3382), .B2(n4752), .A(n3381), .ZN(n3383) );
  INV_X1 U4192 ( .A(n3383), .ZN(U3221) );
  NAND2_X1 U4193 ( .A1(n3329), .A2(n3384), .ZN(n3636) );
  NAND2_X1 U4194 ( .A1(n3636), .A2(n3385), .ZN(n3389) );
  NAND2_X1 U4195 ( .A1(n3387), .A2(n3386), .ZN(n3388) );
  XNOR2_X1 U4196 ( .A(n3389), .B(n3388), .ZN(n3394) );
  INV_X1 U4197 ( .A(n3390), .ZN(n3480) );
  AND2_X1 U4198 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4887) );
  AOI21_X1 U4199 ( .B1(n3740), .B2(n3924), .A(n4887), .ZN(n3392) );
  AOI22_X1 U4200 ( .A1(n2218), .A2(n3553), .B1(n3741), .B2(n3479), .ZN(n3391)
         );
  OAI211_X1 U4201 ( .C1(n4758), .C2(n3480), .A(n3392), .B(n3391), .ZN(n3393)
         );
  AOI21_X1 U4202 ( .B1(n3394), .B2(n4752), .A(n3393), .ZN(n3395) );
  INV_X1 U4203 ( .A(n3395), .ZN(U3233) );
  OR2_X1 U4204 ( .A1(n3349), .A2(n3396), .ZN(n3398) );
  NAND2_X1 U4205 ( .A1(n3398), .A2(n3397), .ZN(n3399) );
  XNOR2_X1 U4206 ( .A(n3399), .B(n3842), .ZN(n3414) );
  INV_X1 U4207 ( .A(n3414), .ZN(n3412) );
  XNOR2_X1 U4208 ( .A(n3400), .B(n3842), .ZN(n3404) );
  OAI22_X1 U4209 ( .A1(n3472), .A2(n4208), .B1(n4207), .B2(n3401), .ZN(n3402)
         );
  AOI21_X1 U4210 ( .B1(n4211), .B2(n3926), .A(n3402), .ZN(n3403) );
  OAI21_X1 U4211 ( .B1(n3404), .B2(n4213), .A(n3403), .ZN(n3413) );
  NAND2_X1 U4212 ( .A1(n3413), .A2(n4223), .ZN(n3411) );
  NAND2_X1 U4213 ( .A1(n3441), .A2(n3405), .ZN(n3406) );
  AND2_X1 U4214 ( .A1(n3496), .A2(n3406), .ZN(n3416) );
  INV_X1 U4215 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3407) );
  OAI22_X1 U4216 ( .A1(n3408), .A2(n4171), .B1(n3407), .B2(n4173), .ZN(n3409)
         );
  AOI21_X1 U4217 ( .B1(n3416), .B2(n4991), .A(n3409), .ZN(n3410) );
  OAI211_X1 U4218 ( .C1(n3412), .C2(n4225), .A(n3411), .B(n3410), .ZN(U3281)
         );
  AOI21_X1 U4219 ( .B1(n3414), .B2(n4285), .A(n3413), .ZN(n3418) );
  INV_X1 U4220 ( .A(n5081), .ZN(n3451) );
  AOI22_X1 U4221 ( .A1(n3416), .A2(n3449), .B1(REG1_REG_9__SCAN_IN), .B2(n3451), .ZN(n3415) );
  OAI21_X1 U4222 ( .B1(n3418), .B2(n3451), .A(n3415), .ZN(U3527) );
  AOI22_X1 U4223 ( .A1(n3416), .A2(n3447), .B1(REG0_REG_9__SCAN_IN), .B2(n5071), .ZN(n3417) );
  OAI21_X1 U4224 ( .B1(n3418), .B2(n5071), .A(n3417), .ZN(U3485) );
  INV_X1 U4225 ( .A(n3419), .ZN(n3421) );
  NOR2_X1 U4226 ( .A1(n3421), .A2(n3420), .ZN(n3422) );
  XNOR2_X1 U4227 ( .A(n3423), .B(n3422), .ZN(n3430) );
  NOR2_X1 U4228 ( .A1(STATE_REG_SCAN_IN), .A2(n3424), .ZN(n4905) );
  AOI21_X1 U4229 ( .B1(n3740), .B2(n3553), .A(n4905), .ZN(n3427) );
  NAND2_X1 U4230 ( .A1(n3705), .A2(n3425), .ZN(n3426) );
  OAI211_X1 U4231 ( .C1(n3719), .C2(n4745), .A(n3427), .B(n3426), .ZN(n3428)
         );
  AOI21_X1 U4232 ( .B1(n3723), .B2(n3580), .A(n3428), .ZN(n3429) );
  OAI21_X1 U4233 ( .B1(n3430), .B2(n3699), .A(n3429), .ZN(U3231) );
  NAND2_X1 U4234 ( .A1(n5062), .A2(n3431), .ZN(n3432) );
  AND2_X1 U4235 ( .A1(n3773), .A2(n3770), .ZN(n3840) );
  XNOR2_X1 U4236 ( .A(n3432), .B(n3840), .ZN(n4970) );
  XNOR2_X1 U4237 ( .A(n3433), .B(n3840), .ZN(n3437) );
  OAI22_X1 U4238 ( .A1(n2627), .A2(n4188), .B1(n4207), .B2(n3434), .ZN(n3435)
         );
  AOI21_X1 U4239 ( .B1(n4185), .B2(n3925), .A(n3435), .ZN(n3436) );
  OAI21_X1 U4240 ( .B1(n3437), .B2(n4213), .A(n3436), .ZN(n3438) );
  AOI21_X1 U4241 ( .B1(n3502), .B2(n4970), .A(n3438), .ZN(n4973) );
  INV_X1 U4242 ( .A(n4973), .ZN(n3439) );
  AOI21_X1 U4243 ( .B1(n5055), .B2(n4970), .A(n3439), .ZN(n3452) );
  INV_X1 U4244 ( .A(n3440), .ZN(n3443) );
  INV_X1 U4245 ( .A(n3441), .ZN(n3442) );
  AOI21_X1 U4246 ( .B1(n3444), .B2(n3443), .A(n3442), .ZN(n4969) );
  INV_X1 U4247 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3445) );
  NOR2_X1 U4248 ( .A1(n5073), .A2(n3445), .ZN(n3446) );
  AOI21_X1 U4249 ( .B1(n4969), .B2(n3447), .A(n3446), .ZN(n3448) );
  OAI21_X1 U4250 ( .B1(n3452), .B2(n5071), .A(n3448), .ZN(U3483) );
  AOI22_X1 U4251 ( .A1(n4969), .A2(n3449), .B1(n3451), .B2(REG1_REG_8__SCAN_IN), .ZN(n3450) );
  OAI21_X1 U4252 ( .B1(n3452), .B2(n3451), .A(n3450), .ZN(U3526) );
  NAND2_X1 U4253 ( .A1(n3454), .A2(n3453), .ZN(n3548) );
  AND2_X1 U4254 ( .A1(n3545), .A2(n3546), .ZN(n3841) );
  XNOR2_X1 U4255 ( .A(n3548), .B(n3841), .ZN(n3458) );
  AOI22_X1 U4256 ( .A1(n3523), .A2(n4185), .B1(n4231), .B2(n3455), .ZN(n3456)
         );
  OAI21_X1 U4257 ( .B1(n3505), .B2(n4188), .A(n3456), .ZN(n3457) );
  AOI21_X1 U4258 ( .B1(n3458), .B2(n4183), .A(n3457), .ZN(n3517) );
  INV_X1 U4259 ( .A(n3841), .ZN(n3460) );
  XNOR2_X1 U4260 ( .A(n3459), .B(n3460), .ZN(n3516) );
  OR2_X1 U4261 ( .A1(n3478), .A2(n3461), .ZN(n3462) );
  NAND2_X1 U4262 ( .A1(n3538), .A2(n3462), .ZN(n3522) );
  AOI22_X1 U4263 ( .A1(n4762), .A2(REG2_REG_12__SCAN_IN), .B1(n3463), .B2(
        n4987), .ZN(n3464) );
  OAI21_X1 U4264 ( .B1(n3522), .B2(n4221), .A(n3464), .ZN(n3465) );
  AOI21_X1 U4265 ( .B1(n3516), .B2(n4167), .A(n3465), .ZN(n3466) );
  OAI21_X1 U4266 ( .B1(n4762), .B2(n3517), .A(n3466), .ZN(U3278) );
  NAND2_X1 U4267 ( .A1(n3467), .A2(n3846), .ZN(n3468) );
  NAND2_X1 U4268 ( .A1(n3469), .A2(n3468), .ZN(n3474) );
  INV_X1 U4269 ( .A(n3474), .ZN(n5066) );
  XOR2_X1 U4270 ( .A(n3846), .B(n3470), .Z(n3476) );
  AOI22_X1 U4271 ( .A1(n3553), .A2(n4185), .B1(n4231), .B2(n3479), .ZN(n3471)
         );
  OAI21_X1 U4272 ( .B1(n3472), .B2(n4188), .A(n3471), .ZN(n3473) );
  AOI21_X1 U4273 ( .B1(n3474), .B2(n3502), .A(n3473), .ZN(n3475) );
  OAI21_X1 U4274 ( .B1(n4213), .B2(n3476), .A(n3475), .ZN(n5067) );
  NAND2_X1 U4275 ( .A1(n5067), .A2(n4223), .ZN(n3484) );
  INV_X1 U4276 ( .A(n3477), .ZN(n3497) );
  AOI21_X1 U4277 ( .B1(n3479), .B2(n3497), .A(n3478), .ZN(n5069) );
  INV_X1 U4278 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3481) );
  OAI22_X1 U4279 ( .A1(n4173), .A2(n3481), .B1(n3480), .B2(n4171), .ZN(n3482)
         );
  AOI21_X1 U4280 ( .B1(n5069), .B2(n4991), .A(n3482), .ZN(n3483) );
  OAI211_X1 U4281 ( .C1(n5066), .C2(n3485), .A(n3484), .B(n3483), .ZN(U3279)
         );
  XNOR2_X1 U4282 ( .A(n3487), .B(n3486), .ZN(n3488) );
  XNOR2_X1 U4283 ( .A(n3489), .B(n3488), .ZN(n3494) );
  INV_X1 U4284 ( .A(n3490), .ZN(n3532) );
  AND2_X1 U4285 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4915) );
  AOI21_X1 U4286 ( .B1(n2218), .B2(n3922), .A(n4915), .ZN(n3492) );
  AOI22_X1 U4287 ( .A1(n3740), .A2(n3523), .B1(n3741), .B2(n3531), .ZN(n3491)
         );
  OAI211_X1 U4288 ( .C1(n4758), .C2(n3532), .A(n3492), .B(n3491), .ZN(n3493)
         );
  AOI21_X1 U4289 ( .B1(n3494), .B2(n4752), .A(n3493), .ZN(n3495) );
  INV_X1 U4290 ( .A(n3495), .ZN(U3212) );
  INV_X1 U4291 ( .A(n3496), .ZN(n3499) );
  OAI21_X1 U4292 ( .B1(n3499), .B2(n3498), .A(n3497), .ZN(n4962) );
  AND2_X1 U4293 ( .A1(n3793), .A2(n3789), .ZN(n3860) );
  INV_X1 U4294 ( .A(n3860), .ZN(n3500) );
  XNOR2_X1 U4295 ( .A(n3501), .B(n3500), .ZN(n4964) );
  NAND2_X1 U4296 ( .A1(n4964), .A2(n3502), .ZN(n3509) );
  XNOR2_X1 U4297 ( .A(n3503), .B(n3860), .ZN(n3507) );
  AOI22_X1 U4298 ( .A1(n3925), .A2(n4211), .B1(n4231), .B2(n3639), .ZN(n3504)
         );
  OAI21_X1 U4299 ( .B1(n3505), .B2(n4208), .A(n3504), .ZN(n3506) );
  AOI21_X1 U4300 ( .B1(n3507), .B2(n4183), .A(n3506), .ZN(n3508) );
  NAND2_X1 U4301 ( .A1(n4964), .A2(n5055), .ZN(n3510) );
  AND2_X1 U4302 ( .A1(n4967), .A2(n3510), .ZN(n3513) );
  INV_X1 U4303 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3511) );
  MUX2_X1 U4304 ( .A(n3513), .B(n3511), .S(n5071), .Z(n3512) );
  OAI21_X1 U4305 ( .B1(n4962), .B2(n4706), .A(n3512), .ZN(U3487) );
  INV_X1 U4306 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3514) );
  MUX2_X1 U4307 ( .A(n3514), .B(n3513), .S(n5081), .Z(n3515) );
  OAI21_X1 U4308 ( .B1(n4962), .B2(n4288), .A(n3515), .ZN(U3528) );
  NAND2_X1 U4309 ( .A1(n3516), .A2(n4285), .ZN(n3518) );
  AND2_X1 U4310 ( .A1(n3518), .A2(n3517), .ZN(n3520) );
  INV_X1 U4311 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4605) );
  MUX2_X1 U4312 ( .A(n3520), .B(n4605), .S(n3451), .Z(n3519) );
  OAI21_X1 U4313 ( .B1(n3522), .B2(n4288), .A(n3519), .ZN(U3530) );
  INV_X1 U4314 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4337) );
  MUX2_X1 U4315 ( .A(n4337), .B(n3520), .S(n5073), .Z(n3521) );
  OAI21_X1 U4316 ( .B1(n3522), .B2(n4706), .A(n3521), .ZN(U3491) );
  OAI21_X1 U4317 ( .B1(n3865), .B2(n3875), .A(n3564), .ZN(n3530) );
  INV_X1 U4318 ( .A(n3523), .ZN(n3525) );
  AOI22_X1 U4319 ( .A1(n3922), .A2(n4185), .B1(n4231), .B2(n3531), .ZN(n3524)
         );
  OAI21_X1 U4320 ( .B1(n3525), .B2(n4188), .A(n3524), .ZN(n3529) );
  AOI21_X1 U4321 ( .B1(n3865), .B2(n3526), .A(n3562), .ZN(n4293) );
  NOR2_X1 U4322 ( .A1(n4293), .A2(n3527), .ZN(n3528) );
  AOI211_X1 U4323 ( .C1(n4183), .C2(n3530), .A(n3529), .B(n3528), .ZN(n4292)
         );
  INV_X1 U4324 ( .A(n4293), .ZN(n3536) );
  NAND2_X1 U4325 ( .A1(n3539), .A2(n3531), .ZN(n4289) );
  AND3_X1 U4326 ( .A1(n4290), .A2(n4991), .A3(n4289), .ZN(n3535) );
  INV_X1 U4327 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3533) );
  OAI22_X1 U4328 ( .A1(n4173), .A2(n3533), .B1(n3532), .B2(n4171), .ZN(n3534)
         );
  AOI211_X1 U4329 ( .C1(n3536), .C2(n4992), .A(n3535), .B(n3534), .ZN(n3537)
         );
  OAI21_X1 U4330 ( .B1(n4292), .B2(n4762), .A(n3537), .ZN(U3276) );
  INV_X1 U4331 ( .A(n3538), .ZN(n3540) );
  OAI21_X1 U4332 ( .B1(n3540), .B2(n3551), .A(n3539), .ZN(n3583) );
  INV_X1 U4333 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3556) );
  INV_X1 U4334 ( .A(n3542), .ZN(n3544) );
  OR2_X1 U4335 ( .A1(n3544), .A2(n3543), .ZN(n3549) );
  XNOR2_X1 U4336 ( .A(n3541), .B(n3549), .ZN(n3585) );
  INV_X1 U4337 ( .A(n3545), .ZN(n3547) );
  OAI21_X1 U4338 ( .B1(n3548), .B2(n3547), .A(n3546), .ZN(n3550) );
  INV_X1 U4339 ( .A(n3549), .ZN(n3839) );
  XNOR2_X1 U4340 ( .A(n3550), .B(n3839), .ZN(n3555) );
  OAI22_X1 U4341 ( .A1(n4745), .A2(n4208), .B1(n4207), .B2(n3551), .ZN(n3552)
         );
  AOI21_X1 U4342 ( .B1(n4211), .B2(n3553), .A(n3552), .ZN(n3554) );
  OAI21_X1 U4343 ( .B1(n3555), .B2(n4213), .A(n3554), .ZN(n3579) );
  AOI21_X1 U4344 ( .B1(n4285), .B2(n3585), .A(n3579), .ZN(n3558) );
  MUX2_X1 U4345 ( .A(n3556), .B(n3558), .S(n5073), .Z(n3557) );
  OAI21_X1 U4346 ( .B1(n3583), .B2(n4706), .A(n3557), .ZN(U3493) );
  INV_X1 U4347 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3559) );
  MUX2_X1 U4348 ( .A(n3559), .B(n3558), .S(n5081), .Z(n3560) );
  OAI21_X1 U4349 ( .B1(n4288), .B2(n3583), .A(n3560), .ZN(U3531) );
  NOR2_X1 U4350 ( .A1(n3562), .A2(n3561), .ZN(n3563) );
  INV_X1 U4351 ( .A(n3565), .ZN(n3856) );
  XNOR2_X1 U4352 ( .A(n3563), .B(n3856), .ZN(n4286) );
  INV_X1 U4353 ( .A(n4286), .ZN(n3578) );
  NAND2_X1 U4354 ( .A1(n3564), .A2(n3796), .ZN(n3566) );
  XNOR2_X1 U4355 ( .A(n3566), .B(n3565), .ZN(n3570) );
  OAI22_X1 U4356 ( .A1(n3567), .A2(n4208), .B1(n4742), .B2(n4207), .ZN(n3568)
         );
  AOI21_X1 U4357 ( .B1(n4211), .B2(n3923), .A(n3568), .ZN(n3569) );
  OAI21_X1 U4358 ( .B1(n3570), .B2(n4213), .A(n3569), .ZN(n4284) );
  INV_X1 U4359 ( .A(n3594), .ZN(n3573) );
  NAND2_X1 U4360 ( .A1(n4290), .A2(n3571), .ZN(n3572) );
  NAND2_X1 U4361 ( .A1(n3573), .A2(n3572), .ZN(n4707) );
  AOI22_X1 U4362 ( .A1(n4762), .A2(REG2_REG_15__SCAN_IN), .B1(n3574), .B2(
        n4987), .ZN(n3575) );
  OAI21_X1 U4363 ( .B1(n4707), .B2(n4221), .A(n3575), .ZN(n3576) );
  AOI21_X1 U4364 ( .B1(n4284), .B2(n4223), .A(n3576), .ZN(n3577) );
  OAI21_X1 U4365 ( .B1(n3578), .B2(n4225), .A(n3577), .ZN(U3275) );
  NAND2_X1 U4366 ( .A1(n3579), .A2(n4223), .ZN(n3582) );
  AOI22_X1 U4367 ( .A1(n4762), .A2(REG2_REG_13__SCAN_IN), .B1(n3580), .B2(
        n4987), .ZN(n3581) );
  OAI211_X1 U4368 ( .C1(n3583), .C2(n4221), .A(n3582), .B(n3581), .ZN(n3584)
         );
  AOI21_X1 U4369 ( .B1(n4167), .B2(n3585), .A(n3584), .ZN(n3586) );
  INV_X1 U4370 ( .A(n3586), .ZN(U3277) );
  INV_X1 U4371 ( .A(n3587), .ZN(n3588) );
  AOI21_X1 U4372 ( .B1(n3864), .B2(n3589), .A(n3588), .ZN(n4282) );
  INV_X1 U4373 ( .A(n4282), .ZN(n3599) );
  XNOR2_X1 U4374 ( .A(n3590), .B(n3864), .ZN(n3593) );
  OAI22_X1 U4375 ( .A1(n4189), .A2(n4208), .B1(n4207), .B2(n4731), .ZN(n3591)
         );
  AOI21_X1 U4376 ( .B1(n4211), .B2(n3922), .A(n3591), .ZN(n3592) );
  OAI21_X1 U4377 ( .B1(n3593), .B2(n4213), .A(n3592), .ZN(n4281) );
  OAI21_X1 U4378 ( .B1(n3594), .B2(n4731), .A(n4215), .ZN(n4702) );
  NOR2_X1 U4379 ( .A1(n4702), .A2(n4221), .ZN(n3597) );
  INV_X1 U4380 ( .A(REG2_REG_16__SCAN_IN), .ZN(n3595) );
  OAI22_X1 U4381 ( .A1(n4173), .A2(n3595), .B1(n4741), .B2(n4171), .ZN(n3596)
         );
  AOI211_X1 U4382 ( .C1(n4281), .C2(n4223), .A(n3597), .B(n3596), .ZN(n3598)
         );
  OAI21_X1 U4383 ( .B1(n3599), .B2(n4225), .A(n3598), .ZN(U3274) );
  XNOR2_X1 U4384 ( .A(n4186), .B(n4169), .ZN(n3852) );
  XOR2_X1 U4385 ( .A(n3852), .B(n3600), .Z(n4272) );
  NAND2_X1 U4386 ( .A1(n3601), .A2(n3858), .ZN(n4182) );
  INV_X1 U4387 ( .A(n3602), .ZN(n3604) );
  OAI21_X1 U4388 ( .B1(n4182), .B2(n3604), .A(n3603), .ZN(n3605) );
  XOR2_X1 U4389 ( .A(n3852), .B(n3605), .Z(n3609) );
  OAI22_X1 U4390 ( .A1(n3606), .A2(n4208), .B1(n4207), .B2(n4169), .ZN(n3607)
         );
  AOI21_X1 U4391 ( .B1(n4211), .B2(n3921), .A(n3607), .ZN(n3608) );
  OAI21_X1 U4392 ( .B1(n3609), .B2(n4213), .A(n3608), .ZN(n4269) );
  XNOR2_X1 U4393 ( .A(n4196), .B(n3646), .ZN(n4270) );
  INV_X1 U4394 ( .A(n4270), .ZN(n3611) );
  AOI22_X1 U4395 ( .A1(n4762), .A2(REG2_REG_19__SCAN_IN), .B1(n3653), .B2(
        n4987), .ZN(n3610) );
  OAI21_X1 U4396 ( .B1(n3611), .B2(n4221), .A(n3610), .ZN(n3612) );
  AOI21_X1 U4397 ( .B1(n4269), .B2(n4223), .A(n3612), .ZN(n3613) );
  OAI21_X1 U4398 ( .B1(n4272), .B2(n4225), .A(n3613), .ZN(U3271) );
  NAND3_X1 U4399 ( .A1(n3614), .A2(STATE_REG_SCAN_IN), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n3616) );
  INV_X1 U4400 ( .A(DATAI_31_), .ZN(n3615) );
  OAI22_X1 U4401 ( .A1(n2444), .A2(n3616), .B1(STATE_REG_SCAN_IN), .B2(n3615), 
        .ZN(U3321) );
  XNOR2_X1 U4402 ( .A(n3618), .B(n3617), .ZN(n3624) );
  AOI22_X1 U4403 ( .A1(n2218), .A2(n4033), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3620) );
  AOI22_X1 U4404 ( .A1(n3740), .A2(n3851), .B1(n3741), .B2(n4036), .ZN(n3619)
         );
  OAI211_X1 U4405 ( .C1(n4758), .C2(n3621), .A(n3620), .B(n3619), .ZN(n3622)
         );
  INV_X1 U4406 ( .A(n3622), .ZN(n3623) );
  OAI21_X1 U4407 ( .B1(n3624), .B2(n3699), .A(n3623), .ZN(U3211) );
  AOI21_X1 U4408 ( .B1(n3713), .B2(n3626), .A(n3625), .ZN(n3627) );
  NOR3_X1 U4409 ( .A1(n3628), .A2(n3627), .A3(n3699), .ZN(n3634) );
  INV_X1 U4410 ( .A(n3629), .ZN(n4117) );
  AOI22_X1 U4411 ( .A1(n3920), .A2(n3740), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3632) );
  AOI22_X1 U4412 ( .A1(n2218), .A2(n4110), .B1(n3741), .B2(n3630), .ZN(n3631)
         );
  OAI211_X1 U4413 ( .C1(n4758), .C2(n4117), .A(n3632), .B(n3631), .ZN(n3633)
         );
  OR2_X1 U4414 ( .A1(n3634), .A2(n3633), .ZN(U3213) );
  AND2_X1 U4415 ( .A1(n3329), .A2(n3635), .ZN(n3638) );
  OAI211_X1 U4416 ( .C1(n3638), .C2(n3637), .A(n4752), .B(n3636), .ZN(n3645)
         );
  INV_X1 U4417 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4606) );
  NOR2_X1 U4418 ( .A1(STATE_REG_SCAN_IN), .A2(n4606), .ZN(n4876) );
  AOI21_X1 U4419 ( .B1(n3740), .B2(n3925), .A(n4876), .ZN(n3644) );
  AOI22_X1 U4420 ( .A1(n3640), .A2(n2218), .B1(n3639), .B2(n3705), .ZN(n3643)
         );
  OR2_X1 U4421 ( .A1(n4758), .A2(n3641), .ZN(n3642) );
  NAND4_X1 U4422 ( .A1(n3645), .A2(n3644), .A3(n3643), .A4(n3642), .ZN(U3214)
         );
  AOI22_X1 U4423 ( .A1(n2218), .A2(n4148), .B1(n3741), .B2(n3646), .ZN(n3647)
         );
  NAND2_X1 U4424 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3997) );
  OAI211_X1 U4425 ( .C1(n4209), .C2(n4744), .A(n3647), .B(n3997), .ZN(n3652)
         );
  XOR2_X1 U4426 ( .A(n3649), .B(n3648), .Z(n3650) );
  NOR2_X1 U4427 ( .A1(n3650), .A2(n3699), .ZN(n3651) );
  AOI211_X1 U4428 ( .C1(n3653), .C2(n3723), .A(n3652), .B(n3651), .ZN(n3654)
         );
  INV_X1 U4429 ( .A(n3654), .ZN(U3216) );
  INV_X1 U4430 ( .A(n3701), .ZN(n3655) );
  OAI21_X1 U4431 ( .B1(n3703), .B2(n3655), .A(n3702), .ZN(n3659) );
  XOR2_X1 U4432 ( .A(n3657), .B(n3656), .Z(n3658) );
  XNOR2_X1 U4433 ( .A(n3659), .B(n3658), .ZN(n3665) );
  AOI22_X1 U4434 ( .A1(n3740), .A2(n4148), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3662) );
  NAND2_X1 U4435 ( .A1(n3741), .A2(n3660), .ZN(n3661) );
  OAI211_X1 U4436 ( .C1(n4142), .C2(n3719), .A(n3662), .B(n3661), .ZN(n3663)
         );
  AOI21_X1 U4437 ( .B1(n3723), .B2(n4153), .A(n3663), .ZN(n3664) );
  OAI21_X1 U4438 ( .B1(n3665), .B2(n3699), .A(n3664), .ZN(U3220) );
  INV_X1 U4439 ( .A(n3666), .ZN(n3668) );
  NAND2_X1 U4440 ( .A1(n3668), .A2(n3667), .ZN(n3669) );
  XNOR2_X1 U4441 ( .A(n3670), .B(n3669), .ZN(n3676) );
  INV_X1 U4442 ( .A(n4072), .ZN(n3674) );
  AOI22_X1 U4443 ( .A1(n3740), .A2(n4110), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3673) );
  AOI22_X1 U4444 ( .A1(n2218), .A2(n3851), .B1(n3741), .B2(n3671), .ZN(n3672)
         );
  OAI211_X1 U4445 ( .C1(n4758), .C2(n3674), .A(n3673), .B(n3672), .ZN(n3675)
         );
  AOI21_X1 U4446 ( .B1(n3676), .B2(n4752), .A(n3675), .ZN(n3677) );
  INV_X1 U4447 ( .A(n3677), .ZN(U3222) );
  XNOR2_X1 U4448 ( .A(n3679), .B(n3678), .ZN(n3680) );
  XNOR2_X1 U4449 ( .A(n3681), .B(n3680), .ZN(n3687) );
  INV_X1 U4450 ( .A(n4219), .ZN(n3685) );
  AOI22_X1 U4451 ( .A1(n3921), .A2(n2218), .B1(n3682), .B2(n3705), .ZN(n3684)
         );
  AND2_X1 U4452 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4944) );
  AOI21_X1 U4453 ( .B1(n4747), .B2(n3740), .A(n4944), .ZN(n3683) );
  OAI211_X1 U4454 ( .C1(n4758), .C2(n3685), .A(n3684), .B(n3683), .ZN(n3686)
         );
  AOI21_X1 U4455 ( .B1(n3687), .B2(n4752), .A(n3686), .ZN(n3688) );
  INV_X1 U4456 ( .A(n3688), .ZN(U3225) );
  INV_X1 U4457 ( .A(n3689), .ZN(n3691) );
  NAND2_X1 U4458 ( .A1(n3691), .A2(n3690), .ZN(n3693) );
  XNOR2_X1 U4459 ( .A(n3693), .B(n3692), .ZN(n3700) );
  AOI22_X1 U4460 ( .A1(n3740), .A2(n4135), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3696) );
  NAND2_X1 U4461 ( .A1(n3705), .A2(n3694), .ZN(n3695) );
  OAI211_X1 U4462 ( .C1(n4083), .C2(n3719), .A(n3696), .B(n3695), .ZN(n3697)
         );
  AOI21_X1 U4463 ( .B1(n3723), .B2(n4090), .A(n3697), .ZN(n3698) );
  OAI21_X1 U4464 ( .B1(n3700), .B2(n3699), .A(n3698), .ZN(U3226) );
  NAND2_X1 U4465 ( .A1(n3702), .A2(n3701), .ZN(n3704) );
  XOR2_X1 U4466 ( .A(n3704), .B(n3703), .Z(n3711) );
  AOI22_X1 U4467 ( .A1(n3740), .A2(n4186), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n3709) );
  AOI22_X1 U4468 ( .A1(n3707), .A2(n2218), .B1(n3706), .B2(n3705), .ZN(n3708)
         );
  OAI211_X1 U4469 ( .C1(n4758), .C2(n4172), .A(n3709), .B(n3708), .ZN(n3710)
         );
  AOI21_X1 U4470 ( .B1(n3711), .B2(n4752), .A(n3710), .ZN(n3712) );
  INV_X1 U4471 ( .A(n3712), .ZN(U3230) );
  OAI21_X1 U4472 ( .B1(n3715), .B2(n3714), .A(n3713), .ZN(n3716) );
  NAND2_X1 U4473 ( .A1(n3716), .A2(n4752), .ZN(n3725) );
  OAI22_X1 U4474 ( .A1(n4744), .A2(n4158), .B1(STATE_REG_SCAN_IN), .B2(n3717), 
        .ZN(n3722) );
  OAI22_X1 U4475 ( .A1(n3720), .A2(n3719), .B1(n4743), .B2(n3718), .ZN(n3721)
         );
  AOI211_X1 U4476 ( .C1(n4127), .C2(n3723), .A(n3722), .B(n3721), .ZN(n3724)
         );
  NAND2_X1 U4477 ( .A1(n3725), .A2(n3724), .ZN(U3232) );
  INV_X1 U4478 ( .A(n3726), .ZN(n3728) );
  NOR2_X1 U4479 ( .A1(n3728), .A2(n3727), .ZN(n3729) );
  XNOR2_X1 U4480 ( .A(n3730), .B(n3729), .ZN(n3735) );
  INV_X1 U4481 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4515) );
  NOR2_X1 U4482 ( .A1(STATE_REG_SCAN_IN), .A2(n4515), .ZN(n4952) );
  AOI21_X1 U4483 ( .B1(n4734), .B2(n3740), .A(n4952), .ZN(n3732) );
  AOI22_X1 U4484 ( .A1(n2218), .A2(n4186), .B1(n3741), .B2(n4193), .ZN(n3731)
         );
  OAI211_X1 U4485 ( .C1(n4758), .C2(n3733), .A(n3732), .B(n3731), .ZN(n3734)
         );
  AOI21_X1 U4486 ( .B1(n3735), .B2(n4752), .A(n3734), .ZN(n3736) );
  INV_X1 U4487 ( .A(n3736), .ZN(U3235) );
  NOR2_X1 U4488 ( .A1(n2243), .A2(n3737), .ZN(n3738) );
  XNOR2_X1 U4489 ( .A(n3739), .B(n3738), .ZN(n3746) );
  AOI22_X1 U4490 ( .A1(n3919), .A2(n3740), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3744) );
  AOI22_X1 U4491 ( .A1(n2218), .A2(n4051), .B1(n3741), .B2(n3033), .ZN(n3743)
         );
  OAI211_X1 U4492 ( .C1(n4758), .C2(n4057), .A(n3744), .B(n3743), .ZN(n3745)
         );
  AOI21_X1 U4493 ( .B1(n3746), .B2(n4752), .A(n3745), .ZN(n3747) );
  INV_X1 U4494 ( .A(n3747), .ZN(U3237) );
  INV_X1 U4495 ( .A(n3833), .ZN(n3748) );
  NOR2_X1 U4496 ( .A1(n3748), .A2(n3834), .ZN(n3892) );
  INV_X1 U4497 ( .A(n3749), .ZN(n3751) );
  NOR2_X1 U4498 ( .A1(n3751), .A2(n3750), .ZN(n3883) );
  OAI211_X1 U4499 ( .C1(n3754), .C2(n3905), .A(n3753), .B(n3752), .ZN(n3757)
         );
  NAND3_X1 U4500 ( .A1(n3757), .A2(n3756), .A3(n3755), .ZN(n3760) );
  NAND3_X1 U4501 ( .A1(n3760), .A2(n3759), .A3(n3758), .ZN(n3763) );
  NAND3_X1 U4502 ( .A1(n3763), .A2(n3762), .A3(n3761), .ZN(n3767) );
  INV_X1 U4503 ( .A(n3764), .ZN(n3765) );
  NAND4_X1 U4504 ( .A1(n3767), .A2(n3766), .A3(n3765), .A4(n3779), .ZN(n3769)
         );
  NAND3_X1 U4505 ( .A1(n3769), .A2(n3845), .A3(n3768), .ZN(n3776) );
  AND2_X1 U4506 ( .A1(n3771), .A2(n3770), .ZN(n3780) );
  INV_X1 U4507 ( .A(n3772), .ZN(n3775) );
  INV_X1 U4508 ( .A(n3773), .ZN(n3774) );
  AOI211_X1 U4509 ( .C1(n3776), .C2(n3780), .A(n3775), .B(n3774), .ZN(n3788)
         );
  NAND2_X1 U4510 ( .A1(n3778), .A2(n3777), .ZN(n3787) );
  INV_X1 U4511 ( .A(n3779), .ZN(n3783) );
  INV_X1 U4512 ( .A(n3780), .ZN(n3782) );
  NOR3_X1 U4513 ( .A1(n3783), .A2(n3782), .A3(n3781), .ZN(n3785) );
  INV_X1 U4514 ( .A(n3793), .ZN(n3784) );
  NAND2_X1 U4515 ( .A1(n3787), .A2(n3795), .ZN(n3873) );
  OAI21_X1 U4516 ( .B1(n3785), .B2(n3784), .A(n3873), .ZN(n3786) );
  OAI21_X1 U4517 ( .B1(n3788), .B2(n3787), .A(n3786), .ZN(n3801) );
  NAND2_X1 U4518 ( .A1(n3790), .A2(n3789), .ZN(n3792) );
  AOI211_X1 U4519 ( .C1(n3794), .C2(n3793), .A(n3792), .B(n3791), .ZN(n3800)
         );
  NAND2_X1 U4520 ( .A1(n3796), .A2(n3795), .ZN(n3874) );
  INV_X1 U4521 ( .A(n3874), .ZN(n3797) );
  NAND2_X1 U4522 ( .A1(n3798), .A2(n3797), .ZN(n3799) );
  AOI22_X1 U4523 ( .A1(n3801), .A2(n3800), .B1(n3873), .B2(n3799), .ZN(n3803)
         );
  INV_X1 U4524 ( .A(n3878), .ZN(n3802) );
  OAI21_X1 U4525 ( .B1(n3803), .B2(n3802), .A(n3876), .ZN(n3804) );
  NAND3_X1 U4526 ( .A1(n3804), .A2(n3879), .A3(n2454), .ZN(n3805) );
  AOI211_X1 U4527 ( .C1(n3883), .C2(n3805), .A(n4101), .B(n3881), .ZN(n3806)
         );
  NOR2_X1 U4528 ( .A1(n3806), .A2(n3886), .ZN(n3808) );
  OAI21_X1 U4529 ( .B1(n3808), .B2(n3807), .A(n3887), .ZN(n3810) );
  AOI21_X1 U4530 ( .B1(n3892), .B2(n3810), .A(n3809), .ZN(n3814) );
  AND2_X1 U4531 ( .A1(n3918), .A2(n3821), .ZN(n3811) );
  NOR2_X1 U4532 ( .A1(n3812), .A2(n3811), .ZN(n3894) );
  INV_X1 U4533 ( .A(n3894), .ZN(n3813) );
  NOR4_X1 U4534 ( .A1(n3816), .A2(n3815), .A3(n3814), .A4(n3813), .ZN(n3823)
         );
  OR2_X1 U4535 ( .A1(n3818), .A2(n3817), .ZN(n3890) );
  AND2_X1 U4536 ( .A1(n2525), .A2(DATAI_30_), .ZN(n4232) );
  INV_X1 U4537 ( .A(n4232), .ZN(n3824) );
  NAND2_X1 U4538 ( .A1(n3819), .A2(DATAI_31_), .ZN(n4005) );
  NAND2_X1 U4539 ( .A1(n4004), .A2(n4005), .ZN(n3828) );
  OAI21_X1 U4540 ( .B1(n3825), .B2(n3824), .A(n3828), .ZN(n3830) );
  INV_X1 U4541 ( .A(n3830), .ZN(n3820) );
  OAI21_X1 U4542 ( .B1(n3918), .B2(n3821), .A(n3820), .ZN(n3889) );
  AOI21_X1 U4543 ( .B1(n3890), .B2(n3894), .A(n3889), .ZN(n3896) );
  INV_X1 U4544 ( .A(n3896), .ZN(n3822) );
  NOR2_X1 U4545 ( .A1(n3823), .A2(n3822), .ZN(n3829) );
  NOR2_X1 U4546 ( .A1(n4004), .A2(n4005), .ZN(n3902) );
  INV_X1 U4547 ( .A(n3902), .ZN(n3827) );
  AND2_X1 U4548 ( .A1(n3825), .A2(n3824), .ZN(n3903) );
  INV_X1 U4549 ( .A(n3903), .ZN(n3826) );
  NAND2_X1 U4550 ( .A1(n3827), .A2(n3826), .ZN(n3831) );
  OAI21_X1 U4551 ( .B1(n3829), .B2(n3831), .A(n3828), .ZN(n3909) );
  NOR2_X1 U4552 ( .A1(n3831), .A2(n3830), .ZN(n3832) );
  NAND2_X1 U4553 ( .A1(n4029), .A2(n3832), .ZN(n3850) );
  NAND2_X1 U4554 ( .A1(n3833), .A2(n4044), .ZN(n4064) );
  INV_X1 U4555 ( .A(n4064), .ZN(n3838) );
  NOR2_X1 U4556 ( .A1(n3835), .A2(n3834), .ZN(n4082) );
  NAND2_X1 U4557 ( .A1(n3837), .A2(n3836), .ZN(n4165) );
  NAND4_X1 U4558 ( .A1(n3839), .A2(n3838), .A3(n4082), .A4(n4165), .ZN(n3849)
         );
  NAND4_X1 U4559 ( .A1(n3842), .A2(n4181), .A3(n3841), .A4(n3840), .ZN(n3848)
         );
  NAND4_X1 U4560 ( .A1(n3846), .A2(n3845), .A3(n3844), .A4(n3843), .ZN(n3847)
         );
  NOR4_X1 U4561 ( .A1(n3850), .A2(n3849), .A3(n3848), .A4(n3847), .ZN(n3872)
         );
  XNOR2_X1 U4562 ( .A(n3851), .B(n4055), .ZN(n4046) );
  XNOR2_X1 U4563 ( .A(n4135), .B(n4115), .ZN(n4105) );
  NOR4_X1 U4564 ( .A1(n4046), .A2(n3853), .A3(n4105), .A4(n3852), .ZN(n3871)
         );
  INV_X1 U4565 ( .A(n3854), .ZN(n4102) );
  OR2_X1 U4566 ( .A1(n4101), .A2(n4102), .ZN(n4143) );
  INV_X1 U4567 ( .A(n4143), .ZN(n3857) );
  NAND4_X1 U4568 ( .A1(n3857), .A2(n3098), .A3(n3856), .A4(n5042), .ZN(n3869)
         );
  INV_X1 U4569 ( .A(n3859), .ZN(n3862) );
  NAND4_X1 U4570 ( .A1(n4205), .A2(n3862), .A3(n3861), .A4(n3860), .ZN(n3868)
         );
  NAND4_X1 U4571 ( .A1(n3865), .A2(n4098), .A3(n3864), .A4(n3863), .ZN(n3867)
         );
  NOR4_X1 U4572 ( .A1(n3869), .A2(n3868), .A3(n3867), .A4(n3866), .ZN(n3870)
         );
  AND3_X1 U4573 ( .A1(n3872), .A2(n3871), .A3(n3870), .ZN(n3907) );
  INV_X1 U4574 ( .A(n4005), .ZN(n3904) );
  OAI21_X1 U4575 ( .B1(n3875), .B2(n3874), .A(n3873), .ZN(n3877) );
  NAND2_X1 U4576 ( .A1(n3877), .A2(n3876), .ZN(n3880) );
  NAND4_X1 U4577 ( .A1(n3880), .A2(n3879), .A3(n3878), .A4(n2454), .ZN(n3882)
         );
  AOI21_X1 U4578 ( .B1(n3883), .B2(n3882), .A(n3881), .ZN(n3885) );
  OAI21_X1 U4579 ( .B1(n3886), .B2(n3885), .A(n3884), .ZN(n3888) );
  NAND2_X1 U4580 ( .A1(n3888), .A2(n3887), .ZN(n3891) );
  AOI211_X1 U4581 ( .C1(n3892), .C2(n3891), .A(n3890), .B(n3889), .ZN(n3898)
         );
  NAND3_X1 U4582 ( .A1(n4029), .A2(n3894), .A3(n3893), .ZN(n3895) );
  AOI22_X1 U4583 ( .A1(n3898), .A2(n3897), .B1(n3896), .B2(n3895), .ZN(n3899)
         );
  AOI21_X1 U4584 ( .B1(n4232), .B2(n3900), .A(n3899), .ZN(n3901) );
  AOI211_X1 U4585 ( .C1(n3904), .C2(n3903), .A(n3902), .B(n3901), .ZN(n3906)
         );
  MUX2_X1 U4586 ( .A(n3907), .B(n3906), .S(n3905), .Z(n3908) );
  MUX2_X1 U4587 ( .A(n3909), .B(n3908), .S(n4711), .Z(n3910) );
  XNOR2_X1 U4588 ( .A(n3910), .B(n4712), .ZN(n3917) );
  NAND2_X1 U4589 ( .A1(n4789), .A2(n4787), .ZN(n4796) );
  INV_X1 U4590 ( .A(n3911), .ZN(n3912) );
  NOR2_X1 U4591 ( .A1(n4796), .A2(n3912), .ZN(n3915) );
  OAI21_X1 U4592 ( .B1(n3916), .B2(n3913), .A(B_REG_SCAN_IN), .ZN(n3914) );
  OAI22_X1 U4593 ( .A1(n3917), .A2(n3916), .B1(n3915), .B2(n3914), .ZN(U3239)
         );
  MUX2_X1 U4594 ( .A(n3918), .B(DATAO_REG_29__SCAN_IN), .S(n4791), .Z(U3579)
         );
  MUX2_X1 U4595 ( .A(n4033), .B(DATAO_REG_28__SCAN_IN), .S(n4791), .Z(U3578)
         );
  MUX2_X1 U4596 ( .A(n4051), .B(DATAO_REG_27__SCAN_IN), .S(n4791), .Z(U3577)
         );
  MUX2_X1 U4597 ( .A(DATAO_REG_25__SCAN_IN), .B(n3919), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4598 ( .A(n4110), .B(DATAO_REG_24__SCAN_IN), .S(n4791), .Z(U3574)
         );
  MUX2_X1 U4599 ( .A(DATAO_REG_22__SCAN_IN), .B(n3920), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4600 ( .A(n4148), .B(DATAO_REG_20__SCAN_IN), .S(n4791), .Z(U3570)
         );
  MUX2_X1 U4601 ( .A(n4186), .B(DATAO_REG_19__SCAN_IN), .S(n4791), .Z(U3569)
         );
  MUX2_X1 U4602 ( .A(DATAO_REG_18__SCAN_IN), .B(n3921), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4603 ( .A(DATAO_REG_17__SCAN_IN), .B(n4734), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4604 ( .A(DATAO_REG_16__SCAN_IN), .B(n4747), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4605 ( .A(n3922), .B(DATAO_REG_15__SCAN_IN), .S(n4791), .Z(U3565)
         );
  MUX2_X1 U4606 ( .A(DATAO_REG_14__SCAN_IN), .B(n3923), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4607 ( .A(n3924), .B(DATAO_REG_10__SCAN_IN), .S(n4791), .Z(U3560)
         );
  MUX2_X1 U4608 ( .A(n3925), .B(DATAO_REG_9__SCAN_IN), .S(n4791), .Z(U3559) );
  MUX2_X1 U4609 ( .A(DATAO_REG_8__SCAN_IN), .B(n3926), .S(U4043), .Z(U3558) );
  MUX2_X1 U4610 ( .A(DATAO_REG_7__SCAN_IN), .B(n3927), .S(U4043), .Z(U3557) );
  MUX2_X1 U4611 ( .A(n3928), .B(DATAO_REG_6__SCAN_IN), .S(n4791), .Z(U3556) );
  MUX2_X1 U4612 ( .A(DATAO_REG_5__SCAN_IN), .B(n3929), .S(U4043), .Z(U3555) );
  MUX2_X1 U4613 ( .A(DATAO_REG_4__SCAN_IN), .B(n3930), .S(U4043), .Z(U3554) );
  MUX2_X1 U4614 ( .A(n3931), .B(DATAO_REG_3__SCAN_IN), .S(n4791), .Z(U3553) );
  MUX2_X1 U4615 ( .A(DATAO_REG_2__SCAN_IN), .B(n3932), .S(U4043), .Z(U3552) );
  MUX2_X1 U4616 ( .A(n2989), .B(DATAO_REG_0__SCAN_IN), .S(n4791), .Z(U3550) );
  INV_X1 U4617 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3956) );
  INV_X1 U4618 ( .A(n3991), .ZN(n5013) );
  AOI22_X1 U4619 ( .A1(n3991), .A2(REG1_REG_18__SCAN_IN), .B1(n3956), .B2(
        n5013), .ZN(n4957) );
  INV_X1 U4620 ( .A(n5014), .ZN(n3990) );
  INV_X1 U4621 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4382) );
  AOI22_X1 U4622 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3988), .B1(n5018), .B2(
        n4382), .ZN(n4928) );
  INV_X1 U4623 ( .A(REG1_REG_11__SCAN_IN), .ZN(n5082) );
  AOI22_X1 U4624 ( .A1(n3964), .A2(REG1_REG_11__SCAN_IN), .B1(n5082), .B2(
        n5026), .ZN(n4880) );
  NAND2_X1 U4625 ( .A1(n4856), .A2(REG1_REG_9__SCAN_IN), .ZN(n3944) );
  INV_X1 U4626 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3933) );
  MUX2_X1 U4627 ( .A(n3933), .B(REG1_REG_9__SCAN_IN), .S(n4856), .Z(n3934) );
  INV_X1 U4628 ( .A(n3934), .ZN(n4858) );
  INV_X1 U4629 ( .A(REG1_REG_0__SCAN_IN), .ZN(n5074) );
  INV_X1 U4630 ( .A(REG1_REG_1__SCAN_IN), .ZN(n5076) );
  AOI22_X1 U4631 ( .A1(REG1_REG_1__SCAN_IN), .A2(n4714), .B1(n4774), .B2(n5076), .ZN(n4772) );
  NOR3_X1 U4632 ( .A1(n5038), .A2(n5074), .A3(n4772), .ZN(n4770) );
  AOI22_X1 U4633 ( .A1(n4784), .A2(n4493), .B1(REG1_REG_2__SCAN_IN), .B2(n4716), .ZN(n4781) );
  NOR2_X1 U4634 ( .A1(n3935), .A2(n4729), .ZN(n3936) );
  INV_X1 U4635 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4722) );
  NOR2_X1 U4636 ( .A1(n4722), .A2(n4721), .ZN(n4720) );
  NOR2_X1 U4637 ( .A1(n3937), .A2(n2390), .ZN(n3938) );
  NAND2_X1 U4638 ( .A1(n5035), .A2(REG1_REG_5__SCAN_IN), .ZN(n3939) );
  OAI21_X1 U4639 ( .B1(n5035), .B2(REG1_REG_5__SCAN_IN), .A(n3939), .ZN(n4814)
         );
  AOI21_X1 U4640 ( .B1(REG1_REG_5__SCAN_IN), .B2(n5035), .A(n4813), .ZN(n3941)
         );
  NAND2_X1 U4641 ( .A1(REG1_REG_7__SCAN_IN), .A2(n4835), .ZN(n4834) );
  INV_X1 U4642 ( .A(REG1_REG_7__SCAN_IN), .ZN(n5079) );
  NAND2_X1 U4643 ( .A1(n5029), .A2(n3942), .ZN(n3943) );
  NAND2_X1 U4644 ( .A1(REG1_REG_8__SCAN_IN), .A2(n4847), .ZN(n4846) );
  NAND2_X1 U4645 ( .A1(n3943), .A2(n4846), .ZN(n4859) );
  NAND2_X1 U4646 ( .A1(n4858), .A2(n4859), .ZN(n4857) );
  NAND2_X1 U4647 ( .A1(n3944), .A2(n4857), .ZN(n3945) );
  INV_X1 U4648 ( .A(n3979), .ZN(n5028) );
  XNOR2_X1 U4649 ( .A(n3945), .B(n5028), .ZN(n4870) );
  NAND2_X1 U4650 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4870), .ZN(n4869) );
  NAND2_X1 U4651 ( .A1(n3979), .A2(n3945), .ZN(n3946) );
  NAND2_X1 U4652 ( .A1(n4880), .A2(n4879), .ZN(n4878) );
  NAND2_X1 U4653 ( .A1(n3964), .A2(REG1_REG_11__SCAN_IN), .ZN(n3947) );
  NAND2_X1 U4654 ( .A1(n5023), .A2(n3948), .ZN(n3949) );
  INV_X1 U4655 ( .A(n5023), .ZN(n4895) );
  NAND2_X1 U4656 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4890), .ZN(n4889) );
  NAND2_X1 U4657 ( .A1(n3949), .A2(n4889), .ZN(n4907) );
  INV_X1 U4658 ( .A(n4900), .ZN(n5022) );
  AOI22_X1 U4659 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4900), .B1(n5022), .B2(
        n3559), .ZN(n4908) );
  NAND2_X1 U4660 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4900), .ZN(n3950) );
  NAND2_X1 U4661 ( .A1(n5019), .A2(n3951), .ZN(n3952) );
  INV_X1 U4662 ( .A(n5019), .ZN(n4920) );
  XNOR2_X1 U4663 ( .A(n3951), .B(n4920), .ZN(n4917) );
  NAND2_X1 U4664 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4917), .ZN(n4916) );
  NAND2_X1 U4665 ( .A1(n3952), .A2(n4916), .ZN(n4927) );
  NAND2_X1 U4666 ( .A1(n4928), .A2(n4927), .ZN(n4926) );
  OR2_X1 U4667 ( .A1(n5018), .A2(n4382), .ZN(n3953) );
  INV_X1 U4668 ( .A(n5015), .ZN(n4939) );
  INV_X1 U4669 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4670 ( .A1(n3990), .A2(n3955), .B1(REG1_REG_17__SCAN_IN), .B2(
        n5014), .ZN(n4945) );
  NAND2_X1 U4671 ( .A1(n4957), .A2(n4956), .ZN(n4954) );
  INV_X1 U4672 ( .A(REG1_REG_19__SCAN_IN), .ZN(n3957) );
  MUX2_X1 U4673 ( .A(REG1_REG_19__SCAN_IN), .B(n3957), .S(n3998), .Z(n3958) );
  INV_X1 U4674 ( .A(n3958), .ZN(n3959) );
  NAND2_X1 U4675 ( .A1(n3962), .A2(n3961), .ZN(n4768) );
  INV_X1 U4676 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4677 ( .A1(n3991), .A2(n3963), .B1(REG2_REG_18__SCAN_IN), .B2(
        n5013), .ZN(n4951) );
  INV_X1 U4678 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4639) );
  AOI22_X1 U4679 ( .A1(n3990), .A2(REG2_REG_17__SCAN_IN), .B1(n4639), .B2(
        n5014), .ZN(n4942) );
  AOI22_X1 U4680 ( .A1(n3964), .A2(REG2_REG_11__SCAN_IN), .B1(n3481), .B2(
        n5026), .ZN(n4883) );
  NAND2_X1 U4681 ( .A1(n4856), .A2(REG2_REG_9__SCAN_IN), .ZN(n3978) );
  MUX2_X1 U4682 ( .A(REG2_REG_9__SCAN_IN), .B(n3407), .S(n4856), .Z(n4861) );
  NAND2_X1 U4683 ( .A1(REG2_REG_7__SCAN_IN), .A2(n4835), .ZN(n3975) );
  AOI22_X1 U4684 ( .A1(REG2_REG_7__SCAN_IN), .A2(n4835), .B1(n5032), .B2(n3965), .ZN(n4843) );
  NAND2_X1 U4685 ( .A1(n5035), .A2(REG2_REG_5__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4686 ( .A1(n5035), .A2(REG2_REG_5__SCAN_IN), .B1(n3966), .B2(n4823), .ZN(n4820) );
  INV_X1 U4687 ( .A(REG2_REG_2__SCAN_IN), .ZN(n4641) );
  AOI22_X1 U4688 ( .A1(n4784), .A2(REG2_REG_2__SCAN_IN), .B1(n4641), .B2(n4716), .ZN(n4799) );
  INV_X1 U4689 ( .A(REG2_REG_1__SCAN_IN), .ZN(n4384) );
  AOI22_X1 U4690 ( .A1(REG2_REG_1__SCAN_IN), .A2(n4774), .B1(n4714), .B2(n4384), .ZN(n4776) );
  INV_X1 U4691 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4763) );
  NOR2_X1 U4692 ( .A1(n5038), .A2(n4763), .ZN(n4786) );
  NAND2_X1 U4693 ( .A1(n4776), .A2(n4786), .ZN(n4775) );
  OAI21_X1 U4694 ( .B1(n4714), .B2(n4384), .A(n4775), .ZN(n4798) );
  NAND2_X1 U4695 ( .A1(n4799), .A2(n4798), .ZN(n4797) );
  OAI21_X1 U4696 ( .B1(n4641), .B2(n4716), .A(n4797), .ZN(n3968) );
  NAND2_X1 U4697 ( .A1(n3967), .A2(n3968), .ZN(n3969) );
  XNOR2_X1 U4698 ( .A(n4729), .B(n3968), .ZN(n4726) );
  NAND2_X1 U4699 ( .A1(REG2_REG_3__SCAN_IN), .A2(n4726), .ZN(n4725) );
  NAND2_X1 U4700 ( .A1(n4718), .A2(n3970), .ZN(n3971) );
  NAND2_X1 U4701 ( .A1(n4820), .A2(n4819), .ZN(n4818) );
  NAND2_X1 U4702 ( .A1(n3972), .A2(n4818), .ZN(n3973) );
  NAND2_X1 U4703 ( .A1(n5033), .A2(n3973), .ZN(n3974) );
  XNOR2_X1 U4704 ( .A(n3973), .B(n3940), .ZN(n4831) );
  NAND2_X1 U4705 ( .A1(REG2_REG_6__SCAN_IN), .A2(n4831), .ZN(n4830) );
  NAND2_X1 U4706 ( .A1(n5029), .A2(n3976), .ZN(n3977) );
  NAND2_X1 U4707 ( .A1(n3977), .A2(n4848), .ZN(n4862) );
  NAND2_X1 U4708 ( .A1(n4861), .A2(n4862), .ZN(n4860) );
  NAND2_X1 U4709 ( .A1(n3978), .A2(n4860), .ZN(n3980) );
  NAND2_X1 U4710 ( .A1(n3979), .A2(n3980), .ZN(n3981) );
  XNOR2_X1 U4711 ( .A(n3980), .B(n5028), .ZN(n4872) );
  NAND2_X1 U4712 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4872), .ZN(n4871) );
  NAND2_X1 U4713 ( .A1(n5023), .A2(n3982), .ZN(n3983) );
  INV_X1 U4714 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4899) );
  NAND2_X1 U4715 ( .A1(n4899), .A2(n5022), .ZN(n3984) );
  NOR2_X1 U4716 ( .A1(n3985), .A2(n4920), .ZN(n3986) );
  XOR2_X1 U4717 ( .A(n3985), .B(n5019), .Z(n4913) );
  NAND2_X1 U4718 ( .A1(REG2_REG_15__SCAN_IN), .A2(n3988), .ZN(n3987) );
  OAI21_X1 U4719 ( .B1(REG2_REG_15__SCAN_IN), .B2(n3988), .A(n3987), .ZN(n4922) );
  NAND2_X1 U4720 ( .A1(n2235), .A2(n4939), .ZN(n3989) );
  XNOR2_X1 U4721 ( .A(n2235), .B(n5015), .ZN(n4932) );
  NAND2_X1 U4722 ( .A1(n4932), .A2(n3595), .ZN(n4931) );
  NAND2_X1 U4723 ( .A1(n3989), .A2(n4931), .ZN(n4940) );
  XNOR2_X1 U4724 ( .A(n3998), .B(REG2_REG_19__SCAN_IN), .ZN(n3992) );
  XNOR2_X1 U4725 ( .A(n3993), .B(n3992), .ZN(n4000) );
  NOR2_X2 U4726 ( .A1(n4796), .A2(n4768), .ZN(n4911) );
  INV_X1 U4727 ( .A(n4768), .ZN(n3995) );
  AND2_X1 U4728 ( .A1(n3995), .A2(n3994), .ZN(n4785) );
  NAND2_X1 U4729 ( .A1(n4953), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3996) );
  OAI211_X1 U4730 ( .C1(n4960), .C2(n3998), .A(n3997), .B(n3996), .ZN(n3999)
         );
  AOI21_X1 U4731 ( .B1(n4000), .B2(n4911), .A(n3999), .ZN(n4001) );
  OAI21_X1 U4732 ( .B1(n4002), .B2(n4824), .A(n4001), .ZN(U3259) );
  XNOR2_X1 U4733 ( .A(n4229), .B(n4005), .ZN(n4297) );
  NAND2_X1 U4734 ( .A1(n4004), .A2(n4003), .ZN(n4234) );
  OAI21_X1 U4735 ( .B1(n4005), .B2(n4207), .A(n4234), .ZN(n4294) );
  NAND2_X1 U4736 ( .A1(n4294), .A2(n4223), .ZN(n4007) );
  NAND2_X1 U4737 ( .A1(n4762), .A2(REG2_REG_31__SCAN_IN), .ZN(n4006) );
  OAI211_X1 U4738 ( .C1(n4297), .C2(n4221), .A(n4007), .B(n4006), .ZN(U3260)
         );
  INV_X1 U4739 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4015) );
  NAND2_X1 U4740 ( .A1(n4008), .A2(n4167), .ZN(n4014) );
  OAI22_X1 U4741 ( .A1(n4010), .A2(n4221), .B1(n4009), .B2(n4171), .ZN(n4011)
         );
  OAI21_X1 U4742 ( .B1(n4012), .B2(n4011), .A(n4173), .ZN(n4013) );
  OAI211_X1 U4743 ( .C1(n4173), .C2(n4015), .A(n4014), .B(n4013), .ZN(U3354)
         );
  INV_X1 U4744 ( .A(n4016), .ZN(n4025) );
  NOR2_X1 U4745 ( .A1(n4017), .A2(n4221), .ZN(n4022) );
  INV_X1 U4746 ( .A(REG2_REG_28__SCAN_IN), .ZN(n4020) );
  INV_X1 U4747 ( .A(n4018), .ZN(n4019) );
  OAI22_X1 U4748 ( .A1(n4173), .A2(n4020), .B1(n4019), .B2(n4171), .ZN(n4021)
         );
  OAI21_X1 U4749 ( .B1(n4025), .B2(n4225), .A(n4024), .ZN(U3262) );
  XNOR2_X1 U4750 ( .A(n4027), .B(n4026), .ZN(n4238) );
  INV_X1 U4751 ( .A(n4238), .ZN(n4042) );
  OAI21_X1 U4752 ( .B1(n2226), .B2(n4029), .A(n4028), .ZN(n4030) );
  NAND2_X1 U4753 ( .A1(n4030), .A2(n4183), .ZN(n4035) );
  NOR2_X1 U4754 ( .A1(n4031), .A2(n4207), .ZN(n4032) );
  AOI21_X1 U4755 ( .B1(n4033), .B2(n4185), .A(n4032), .ZN(n4034) );
  OAI211_X1 U4756 ( .C1(n4065), .C2(n4188), .A(n4035), .B(n4034), .ZN(n4237)
         );
  AND2_X1 U4757 ( .A1(n4054), .A2(n4036), .ZN(n4037) );
  OR2_X1 U4758 ( .A1(n4037), .A2(n2240), .ZN(n4304) );
  AOI22_X1 U4759 ( .A1(n4762), .A2(REG2_REG_27__SCAN_IN), .B1(n4038), .B2(
        n4987), .ZN(n4039) );
  OAI21_X1 U4760 ( .B1(n4304), .B2(n4221), .A(n4039), .ZN(n4040) );
  AOI21_X1 U4761 ( .B1(n4237), .B2(n4223), .A(n4040), .ZN(n4041) );
  OAI21_X1 U4762 ( .B1(n4042), .B2(n4225), .A(n4041), .ZN(U3263) );
  XNOR2_X1 U4763 ( .A(n4043), .B(n4046), .ZN(n4242) );
  INV_X1 U4764 ( .A(n4242), .ZN(n4061) );
  NAND2_X1 U4765 ( .A1(n4045), .A2(n4044), .ZN(n4048) );
  INV_X1 U4766 ( .A(n4046), .ZN(n4047) );
  XNOR2_X1 U4767 ( .A(n4048), .B(n4047), .ZN(n4049) );
  NAND2_X1 U4768 ( .A1(n4049), .A2(n4183), .ZN(n4053) );
  NOR2_X1 U4769 ( .A1(n4055), .A2(n4207), .ZN(n4050) );
  AOI21_X1 U4770 ( .B1(n4051), .B2(n4185), .A(n4050), .ZN(n4052) );
  OAI211_X1 U4771 ( .C1(n4083), .C2(n4188), .A(n4053), .B(n4052), .ZN(n4241)
         );
  INV_X1 U4772 ( .A(n4071), .ZN(n4056) );
  OAI21_X1 U4773 ( .B1(n4056), .B2(n4055), .A(n4054), .ZN(n4307) );
  NOR2_X1 U4774 ( .A1(n4307), .A2(n4221), .ZN(n4059) );
  INV_X1 U4775 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4550) );
  OAI22_X1 U4776 ( .A1(n4173), .A2(n4550), .B1(n4057), .B2(n4171), .ZN(n4058)
         );
  AOI211_X1 U4777 ( .C1(n4241), .C2(n4223), .A(n4059), .B(n4058), .ZN(n4060)
         );
  OAI21_X1 U4778 ( .B1(n4061), .B2(n4225), .A(n4060), .ZN(U3264) );
  XNOR2_X1 U4779 ( .A(n4062), .B(n4064), .ZN(n4245) );
  INV_X1 U4780 ( .A(n4245), .ZN(n4076) );
  XNOR2_X1 U4781 ( .A(n4063), .B(n4064), .ZN(n4068) );
  OAI22_X1 U4782 ( .A1(n4065), .A2(n4208), .B1(n4207), .B2(n4069), .ZN(n4066)
         );
  AOI21_X1 U4783 ( .B1(n4211), .B2(n4110), .A(n4066), .ZN(n4067) );
  OAI21_X1 U4784 ( .B1(n4068), .B2(n4213), .A(n4067), .ZN(n4244) );
  OR2_X1 U4785 ( .A1(n4089), .A2(n4069), .ZN(n4070) );
  NAND2_X1 U4786 ( .A1(n4071), .A2(n4070), .ZN(n4311) );
  AOI22_X1 U4787 ( .A1(n4762), .A2(REG2_REG_25__SCAN_IN), .B1(n4072), .B2(
        n4987), .ZN(n4073) );
  OAI21_X1 U4788 ( .B1(n4311), .B2(n4221), .A(n4073), .ZN(n4074) );
  AOI21_X1 U4789 ( .B1(n4244), .B2(n4223), .A(n4074), .ZN(n4075) );
  OAI21_X1 U4790 ( .B1(n4076), .B2(n4225), .A(n4075), .ZN(U3265) );
  XNOR2_X1 U4791 ( .A(n4077), .B(n4082), .ZN(n4249) );
  INV_X1 U4792 ( .A(n4249), .ZN(n4094) );
  INV_X1 U4793 ( .A(n4078), .ZN(n4079) );
  NAND2_X1 U4794 ( .A1(n4080), .A2(n4079), .ZN(n4081) );
  XOR2_X1 U4795 ( .A(n4082), .B(n4081), .Z(n4086) );
  OAI22_X1 U4796 ( .A1(n4083), .A2(n4208), .B1(n4207), .B2(n4087), .ZN(n4084)
         );
  AOI21_X1 U4797 ( .B1(n4211), .B2(n4135), .A(n4084), .ZN(n4085) );
  OAI21_X1 U4798 ( .B1(n4086), .B2(n4213), .A(n4085), .ZN(n4248) );
  NOR2_X1 U4799 ( .A1(n4113), .A2(n4087), .ZN(n4088) );
  OR2_X1 U4800 ( .A1(n4089), .A2(n4088), .ZN(n4315) );
  AOI22_X1 U4801 ( .A1(n4762), .A2(REG2_REG_24__SCAN_IN), .B1(n4090), .B2(
        n4987), .ZN(n4091) );
  OAI21_X1 U4802 ( .B1(n4315), .B2(n4221), .A(n4091), .ZN(n4092) );
  AOI21_X1 U4803 ( .B1(n4248), .B2(n4223), .A(n4092), .ZN(n4093) );
  OAI21_X1 U4804 ( .B1(n4094), .B2(n4225), .A(n4093), .ZN(U3266) );
  OR2_X1 U4805 ( .A1(n4141), .A2(n4095), .ZN(n4097) );
  NAND2_X1 U4806 ( .A1(n4097), .A2(n4096), .ZN(n4122) );
  NOR2_X1 U4807 ( .A1(n4124), .A2(n4099), .ZN(n4100) );
  XNOR2_X1 U4808 ( .A(n4100), .B(n4105), .ZN(n4253) );
  INV_X1 U4809 ( .A(n4253), .ZN(n4121) );
  INV_X1 U4810 ( .A(n4101), .ZN(n4103) );
  AOI21_X1 U4811 ( .B1(n4144), .B2(n4103), .A(n4102), .ZN(n4133) );
  OAI21_X1 U4812 ( .B1(n4133), .B2(n4132), .A(n4104), .ZN(n4107) );
  INV_X1 U4813 ( .A(n4105), .ZN(n4106) );
  XNOR2_X1 U4814 ( .A(n4107), .B(n4106), .ZN(n4108) );
  NAND2_X1 U4815 ( .A1(n4108), .A2(n4183), .ZN(n4112) );
  NOR2_X1 U4816 ( .A1(n4115), .A2(n4207), .ZN(n4109) );
  AOI21_X1 U4817 ( .B1(n4110), .B2(n4185), .A(n4109), .ZN(n4111) );
  OAI211_X1 U4818 ( .C1(n4142), .C2(n4188), .A(n4112), .B(n4111), .ZN(n4252)
         );
  INV_X1 U4819 ( .A(n4126), .ZN(n4116) );
  INV_X1 U4820 ( .A(n4113), .ZN(n4114) );
  OAI21_X1 U4821 ( .B1(n4116), .B2(n4115), .A(n4114), .ZN(n4319) );
  NOR2_X1 U4822 ( .A1(n4319), .A2(n4221), .ZN(n4119) );
  OAI22_X1 U4823 ( .A1(n4173), .A2(n4643), .B1(n4117), .B2(n4171), .ZN(n4118)
         );
  AOI211_X1 U4824 ( .C1(n4252), .C2(n4223), .A(n4119), .B(n4118), .ZN(n4120)
         );
  OAI21_X1 U4825 ( .B1(n4121), .B2(n4225), .A(n4120), .ZN(U3267) );
  NOR2_X1 U4826 ( .A1(n4122), .A2(n4132), .ZN(n4123) );
  NAND2_X1 U4827 ( .A1(n4151), .A2(n4134), .ZN(n4125) );
  NAND2_X1 U4828 ( .A1(n4126), .A2(n4125), .ZN(n4323) );
  INV_X1 U4829 ( .A(n4323), .ZN(n4131) );
  INV_X1 U4830 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4129) );
  INV_X1 U4831 ( .A(n4127), .ZN(n4128) );
  OAI22_X1 U4832 ( .A1(n4173), .A2(n4129), .B1(n4128), .B2(n4171), .ZN(n4130)
         );
  AOI21_X1 U4833 ( .B1(n4131), .B2(n4991), .A(n4130), .ZN(n4140) );
  XNOR2_X1 U4834 ( .A(n4133), .B(n4132), .ZN(n4138) );
  AOI22_X1 U4835 ( .A1(n4135), .A2(n4185), .B1(n4231), .B2(n4134), .ZN(n4136)
         );
  OAI21_X1 U4836 ( .B1(n4158), .B2(n4188), .A(n4136), .ZN(n4137) );
  AOI21_X1 U4837 ( .B1(n4138), .B2(n4183), .A(n4137), .ZN(n4256) );
  OR2_X1 U4838 ( .A1(n4256), .A2(n4762), .ZN(n4139) );
  OAI211_X1 U4839 ( .C1(n4257), .C2(n4225), .A(n4140), .B(n4139), .ZN(U3268)
         );
  XNOR2_X1 U4840 ( .A(n4141), .B(n4143), .ZN(n4261) );
  INV_X1 U4841 ( .A(n4261), .ZN(n4157) );
  OAI22_X1 U4842 ( .A1(n4142), .A2(n4208), .B1(n4207), .B2(n4152), .ZN(n4147)
         );
  XNOR2_X1 U4843 ( .A(n4144), .B(n4143), .ZN(n4145) );
  NOR2_X1 U4844 ( .A1(n4145), .A2(n4213), .ZN(n4146) );
  AOI211_X1 U4845 ( .C1(n4211), .C2(n4148), .A(n4147), .B(n4146), .ZN(n4149)
         );
  INV_X1 U4846 ( .A(n4149), .ZN(n4260) );
  OAI21_X1 U4847 ( .B1(n4150), .B2(n4152), .A(n4151), .ZN(n4327) );
  AOI22_X1 U4848 ( .A1(n4762), .A2(REG2_REG_21__SCAN_IN), .B1(n4153), .B2(
        n4987), .ZN(n4154) );
  OAI21_X1 U4849 ( .B1(n4327), .B2(n4221), .A(n4154), .ZN(n4155) );
  AOI21_X1 U4850 ( .B1(n4260), .B2(n4223), .A(n4155), .ZN(n4156) );
  OAI21_X1 U4851 ( .B1(n4157), .B2(n4225), .A(n4156), .ZN(U3269) );
  OAI22_X1 U4852 ( .A1(n4158), .A2(n4208), .B1(n4207), .B2(n4168), .ZN(n4162)
         );
  XOR2_X1 U4853 ( .A(n4165), .B(n4159), .Z(n4160) );
  NOR2_X1 U4854 ( .A1(n4160), .A2(n4213), .ZN(n4161) );
  AOI211_X1 U4855 ( .C1(n4211), .C2(n4186), .A(n4162), .B(n4161), .ZN(n4264)
         );
  AOI21_X1 U4856 ( .B1(n3600), .B2(n4164), .A(n4163), .ZN(n4166) );
  XNOR2_X1 U4857 ( .A(n4166), .B(n4165), .ZN(n4266) );
  NAND2_X1 U4858 ( .A1(n4266), .A2(n4167), .ZN(n4177) );
  AOI21_X1 U4859 ( .B1(n4196), .B2(n4169), .A(n4168), .ZN(n4170) );
  OR2_X1 U4860 ( .A1(n4150), .A2(n4170), .ZN(n4331) );
  INV_X1 U4861 ( .A(n4331), .ZN(n4175) );
  INV_X1 U4862 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4509) );
  OAI22_X1 U4863 ( .A1(n4173), .A2(n4509), .B1(n4172), .B2(n4171), .ZN(n4174)
         );
  AOI21_X1 U4864 ( .B1(n4175), .B2(n4991), .A(n4174), .ZN(n4176) );
  OAI211_X1 U4865 ( .C1(n4762), .C2(n4264), .A(n4177), .B(n4176), .ZN(U3270)
         );
  NAND2_X1 U4866 ( .A1(n4178), .A2(n4181), .ZN(n4179) );
  NAND2_X1 U4867 ( .A1(n4180), .A2(n4179), .ZN(n4273) );
  INV_X1 U4868 ( .A(n4273), .ZN(n4203) );
  XNOR2_X1 U4869 ( .A(n4182), .B(n4181), .ZN(n4184) );
  NAND2_X1 U4870 ( .A1(n4184), .A2(n4183), .ZN(n4192) );
  AOI22_X1 U4871 ( .A1(n4186), .A2(n4185), .B1(n4231), .B2(n4193), .ZN(n4187)
         );
  OAI21_X1 U4872 ( .B1(n4189), .B2(n4188), .A(n4187), .ZN(n4190) );
  INV_X1 U4873 ( .A(n4190), .ZN(n4191) );
  NAND2_X1 U4874 ( .A1(n4192), .A2(n4191), .ZN(n4275) );
  NAND2_X1 U4875 ( .A1(n4194), .A2(n5070), .ZN(n4195) );
  NOR2_X1 U4876 ( .A1(n4196), .A2(n4195), .ZN(n4274) );
  INV_X1 U4877 ( .A(n4274), .ZN(n4200) );
  AOI22_X1 U4878 ( .A1(n4762), .A2(REG2_REG_18__SCAN_IN), .B1(n4197), .B2(
        n4987), .ZN(n4198) );
  OAI21_X1 U4879 ( .B1(n4200), .B2(n4199), .A(n4198), .ZN(n4201) );
  AOI21_X1 U4880 ( .B1(n4275), .B2(n4223), .A(n4201), .ZN(n4202) );
  OAI21_X1 U4881 ( .B1(n4203), .B2(n4225), .A(n4202), .ZN(U3272) );
  XNOR2_X1 U4882 ( .A(n4204), .B(n4205), .ZN(n4279) );
  INV_X1 U4883 ( .A(n4279), .ZN(n4226) );
  XNOR2_X1 U4884 ( .A(n4206), .B(n4205), .ZN(n4214) );
  OAI22_X1 U4885 ( .A1(n4209), .A2(n4208), .B1(n4207), .B2(n4217), .ZN(n4210)
         );
  AOI21_X1 U4886 ( .B1(n4211), .B2(n4747), .A(n4210), .ZN(n4212) );
  OAI21_X1 U4887 ( .B1(n4214), .B2(n4213), .A(n4212), .ZN(n4278) );
  INV_X1 U4888 ( .A(n4215), .ZN(n4218) );
  AOI22_X1 U4889 ( .A1(n4762), .A2(REG2_REG_17__SCAN_IN), .B1(n4219), .B2(
        n4987), .ZN(n4220) );
  OAI21_X1 U4890 ( .B1(n4698), .B2(n4221), .A(n4220), .ZN(n4222) );
  AOI21_X1 U4891 ( .B1(n4278), .B2(n4223), .A(n4222), .ZN(n4224) );
  OAI21_X1 U4892 ( .B1(n4226), .B2(n4225), .A(n4224), .ZN(U3273) );
  NAND2_X1 U4893 ( .A1(n4294), .A2(n5081), .ZN(n4228) );
  NAND2_X1 U4894 ( .A1(n3451), .A2(REG1_REG_31__SCAN_IN), .ZN(n4227) );
  OAI211_X1 U4895 ( .C1(n4297), .C2(n4288), .A(n4228), .B(n4227), .ZN(U3549)
         );
  AOI21_X1 U4896 ( .B1(n4232), .B2(n4230), .A(n4229), .ZN(n4759) );
  INV_X1 U4897 ( .A(n4759), .ZN(n4300) );
  INV_X1 U4898 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4235) );
  NAND2_X1 U4899 ( .A1(n4232), .A2(n4231), .ZN(n4233) );
  AND2_X1 U4900 ( .A1(n4234), .A2(n4233), .ZN(n4761) );
  MUX2_X1 U4901 ( .A(n4235), .B(n4761), .S(n5081), .Z(n4236) );
  OAI21_X1 U4902 ( .B1(n4300), .B2(n4288), .A(n4236), .ZN(U3548) );
  INV_X1 U4903 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4239) );
  AOI21_X1 U4904 ( .B1(n4238), .B2(n4285), .A(n4237), .ZN(n4301) );
  MUX2_X1 U4905 ( .A(n4239), .B(n4301), .S(n5081), .Z(n4240) );
  OAI21_X1 U4906 ( .B1(n4288), .B2(n4304), .A(n4240), .ZN(U3545) );
  INV_X1 U4907 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4547) );
  AOI21_X1 U4908 ( .B1(n4242), .B2(n4285), .A(n4241), .ZN(n4305) );
  MUX2_X1 U4909 ( .A(n4547), .B(n4305), .S(n5081), .Z(n4243) );
  OAI21_X1 U4910 ( .B1(n4288), .B2(n4307), .A(n4243), .ZN(U3544) );
  INV_X1 U4911 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4246) );
  AOI21_X1 U4912 ( .B1(n4245), .B2(n4285), .A(n4244), .ZN(n4308) );
  MUX2_X1 U4913 ( .A(n4246), .B(n4308), .S(n5081), .Z(n4247) );
  OAI21_X1 U4914 ( .B1(n4288), .B2(n4311), .A(n4247), .ZN(U3543) );
  INV_X1 U4915 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4250) );
  AOI21_X1 U4916 ( .B1(n4249), .B2(n4285), .A(n4248), .ZN(n4312) );
  MUX2_X1 U4917 ( .A(n4250), .B(n4312), .S(n5081), .Z(n4251) );
  OAI21_X1 U4918 ( .B1(n4288), .B2(n4315), .A(n4251), .ZN(U3542) );
  INV_X1 U4919 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4254) );
  AOI21_X1 U4920 ( .B1(n4253), .B2(n4285), .A(n4252), .ZN(n4316) );
  MUX2_X1 U4921 ( .A(n4254), .B(n4316), .S(n5081), .Z(n4255) );
  OAI21_X1 U4922 ( .B1(n4288), .B2(n4319), .A(n4255), .ZN(U3541) );
  INV_X1 U4923 ( .A(n4285), .ZN(n5058) );
  OAI21_X1 U4924 ( .B1(n4257), .B2(n5058), .A(n4256), .ZN(n4320) );
  MUX2_X1 U4925 ( .A(n4320), .B(REG1_REG_22__SCAN_IN), .S(n3451), .Z(n4258) );
  INV_X1 U4926 ( .A(n4258), .ZN(n4259) );
  OAI21_X1 U4927 ( .B1(n4288), .B2(n4323), .A(n4259), .ZN(U3540) );
  INV_X1 U4928 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4262) );
  AOI21_X1 U4929 ( .B1(n4285), .B2(n4261), .A(n4260), .ZN(n4324) );
  MUX2_X1 U4930 ( .A(n4262), .B(n4324), .S(n5081), .Z(n4263) );
  OAI21_X1 U4931 ( .B1(n4288), .B2(n4327), .A(n4263), .ZN(U3539) );
  INV_X1 U4932 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4267) );
  INV_X1 U4933 ( .A(n4264), .ZN(n4265) );
  AOI21_X1 U4934 ( .B1(n4266), .B2(n4285), .A(n4265), .ZN(n4328) );
  MUX2_X1 U4935 ( .A(n4267), .B(n4328), .S(n5081), .Z(n4268) );
  OAI21_X1 U4936 ( .B1(n4288), .B2(n4331), .A(n4268), .ZN(U3538) );
  AOI21_X1 U4937 ( .B1(n5070), .B2(n4270), .A(n4269), .ZN(n4271) );
  OAI21_X1 U4938 ( .B1(n4272), .B2(n5058), .A(n4271), .ZN(n4332) );
  MUX2_X1 U4939 ( .A(REG1_REG_19__SCAN_IN), .B(n4332), .S(n5081), .Z(U3537) );
  NAND2_X1 U4940 ( .A1(n4273), .A2(n4285), .ZN(n4277) );
  NOR2_X1 U4941 ( .A1(n4275), .A2(n4274), .ZN(n4276) );
  NAND2_X1 U4942 ( .A1(n4277), .A2(n4276), .ZN(n4694) );
  MUX2_X1 U4943 ( .A(n4694), .B(REG1_REG_18__SCAN_IN), .S(n3451), .Z(U3536) );
  AOI21_X1 U4944 ( .B1(n4279), .B2(n4285), .A(n4278), .ZN(n4695) );
  MUX2_X1 U4945 ( .A(n3955), .B(n4695), .S(n5081), .Z(n4280) );
  OAI21_X1 U4946 ( .B1(n4288), .B2(n4698), .A(n4280), .ZN(U3535) );
  INV_X1 U4947 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4381) );
  AOI21_X1 U4948 ( .B1(n4282), .B2(n4285), .A(n4281), .ZN(n4699) );
  MUX2_X1 U4949 ( .A(n4381), .B(n4699), .S(n5081), .Z(n4283) );
  OAI21_X1 U4950 ( .B1(n4288), .B2(n4702), .A(n4283), .ZN(U3534) );
  AOI21_X1 U4951 ( .B1(n4286), .B2(n4285), .A(n4284), .ZN(n4703) );
  MUX2_X1 U4952 ( .A(n4382), .B(n4703), .S(n5081), .Z(n4287) );
  OAI21_X1 U4953 ( .B1(n4288), .B2(n4707), .A(n4287), .ZN(U3533) );
  NAND3_X1 U4954 ( .A1(n4290), .A2(n5070), .A3(n4289), .ZN(n4291) );
  OAI211_X1 U4955 ( .C1(n4293), .C2(n5065), .A(n4292), .B(n4291), .ZN(n4708)
         );
  MUX2_X1 U4956 ( .A(REG1_REG_14__SCAN_IN), .B(n4708), .S(n5081), .Z(U3532) );
  NAND2_X1 U4957 ( .A1(n4294), .A2(n5073), .ZN(n4296) );
  NAND2_X1 U4958 ( .A1(n5071), .A2(REG0_REG_31__SCAN_IN), .ZN(n4295) );
  OAI211_X1 U4959 ( .C1(n4297), .C2(n4706), .A(n4296), .B(n4295), .ZN(U3517)
         );
  INV_X1 U4960 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4298) );
  MUX2_X1 U4961 ( .A(n4298), .B(n4761), .S(n5073), .Z(n4299) );
  OAI21_X1 U4962 ( .B1(n4300), .B2(n4706), .A(n4299), .ZN(U3516) );
  INV_X1 U4963 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4302) );
  MUX2_X1 U4964 ( .A(n4302), .B(n4301), .S(n5073), .Z(n4303) );
  OAI21_X1 U4965 ( .B1(n4304), .B2(n4706), .A(n4303), .ZN(U3513) );
  INV_X1 U4966 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4490) );
  MUX2_X1 U4967 ( .A(n4490), .B(n4305), .S(n5073), .Z(n4306) );
  OAI21_X1 U4968 ( .B1(n4307), .B2(n4706), .A(n4306), .ZN(U3512) );
  INV_X1 U4969 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4309) );
  MUX2_X1 U4970 ( .A(n4309), .B(n4308), .S(n5073), .Z(n4310) );
  OAI21_X1 U4971 ( .B1(n4311), .B2(n4706), .A(n4310), .ZN(U3511) );
  INV_X1 U4972 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4313) );
  MUX2_X1 U4973 ( .A(n4313), .B(n4312), .S(n5073), .Z(n4314) );
  OAI21_X1 U4974 ( .B1(n4315), .B2(n4706), .A(n4314), .ZN(U3510) );
  INV_X1 U4975 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4317) );
  MUX2_X1 U4976 ( .A(n4317), .B(n4316), .S(n5073), .Z(n4318) );
  OAI21_X1 U4977 ( .B1(n4319), .B2(n4706), .A(n4318), .ZN(U3509) );
  MUX2_X1 U4978 ( .A(REG0_REG_22__SCAN_IN), .B(n4320), .S(n5073), .Z(n4321) );
  INV_X1 U4979 ( .A(n4321), .ZN(n4322) );
  OAI21_X1 U4980 ( .B1(n4323), .B2(n4706), .A(n4322), .ZN(U3508) );
  INV_X1 U4981 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4325) );
  MUX2_X1 U4982 ( .A(n4325), .B(n4324), .S(n5073), .Z(n4326) );
  OAI21_X1 U4983 ( .B1(n4327), .B2(n4706), .A(n4326), .ZN(U3507) );
  INV_X1 U4984 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4329) );
  MUX2_X1 U4985 ( .A(n4329), .B(n4328), .S(n5073), .Z(n4330) );
  OAI21_X1 U4986 ( .B1(n4331), .B2(n4706), .A(n4330), .ZN(U3506) );
  MUX2_X1 U4987 ( .A(REG0_REG_19__SCAN_IN), .B(n4332), .S(n5073), .Z(n4693) );
  INV_X1 U4988 ( .A(D_REG_19__SCAN_IN), .ZN(n5002) );
  INV_X1 U4989 ( .A(D_REG_22__SCAN_IN), .ZN(n5001) );
  AOI22_X1 U4990 ( .A1(n5002), .A2(keyinput139), .B1(keyinput151), .B2(n5001), 
        .ZN(n4333) );
  OAI221_X1 U4991 ( .B1(n5002), .B2(keyinput139), .C1(n5001), .C2(keyinput151), 
        .A(n4333), .ZN(n4341) );
  INV_X1 U4992 ( .A(D_REG_28__SCAN_IN), .ZN(n4999) );
  INV_X1 U4993 ( .A(D_REG_27__SCAN_IN), .ZN(n5000) );
  AOI22_X1 U4994 ( .A1(n4999), .A2(keyinput206), .B1(keyinput225), .B2(n5000), 
        .ZN(n4334) );
  OAI221_X1 U4995 ( .B1(n4999), .B2(keyinput206), .C1(n5000), .C2(keyinput225), 
        .A(n4334), .ZN(n4340) );
  INV_X1 U4996 ( .A(D_REG_31__SCAN_IN), .ZN(n4997) );
  AOI22_X1 U4997 ( .A1(n4997), .A2(keyinput215), .B1(keyinput194), .B2(n4632), 
        .ZN(n4335) );
  OAI221_X1 U4998 ( .B1(n4997), .B2(keyinput215), .C1(n4632), .C2(keyinput194), 
        .A(n4335), .ZN(n4339) );
  INV_X1 U4999 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4516) );
  AOI22_X1 U5000 ( .A1(n4337), .A2(keyinput138), .B1(n4516), .B2(keyinput185), 
        .ZN(n4336) );
  OAI221_X1 U5001 ( .B1(n4337), .B2(keyinput138), .C1(n4516), .C2(keyinput185), 
        .A(n4336), .ZN(n4338) );
  OR4_X1 U5002 ( .A1(n4341), .A2(n4340), .A3(n4339), .A4(n4338), .ZN(n4488) );
  AOI22_X1 U5003 ( .A1(REG1_REG_18__SCAN_IN), .A2(keyinput243), .B1(
        REG1_REG_27__SCAN_IN), .B2(keyinput147), .ZN(n4342) );
  OAI221_X1 U5004 ( .B1(REG1_REG_18__SCAN_IN), .B2(keyinput243), .C1(
        REG1_REG_27__SCAN_IN), .C2(keyinput147), .A(n4342), .ZN(n4349) );
  AOI22_X1 U5005 ( .A1(REG2_REG_0__SCAN_IN), .A2(keyinput214), .B1(
        REG2_REG_8__SCAN_IN), .B2(keyinput129), .ZN(n4343) );
  OAI221_X1 U5006 ( .B1(REG2_REG_0__SCAN_IN), .B2(keyinput214), .C1(
        REG2_REG_8__SCAN_IN), .C2(keyinput129), .A(n4343), .ZN(n4348) );
  AOI22_X1 U5007 ( .A1(REG2_REG_13__SCAN_IN), .A2(keyinput208), .B1(
        REG2_REG_7__SCAN_IN), .B2(keyinput182), .ZN(n4344) );
  OAI221_X1 U5008 ( .B1(REG2_REG_13__SCAN_IN), .B2(keyinput208), .C1(
        REG2_REG_7__SCAN_IN), .C2(keyinput182), .A(n4344), .ZN(n4347) );
  AOI22_X1 U5009 ( .A1(REG2_REG_24__SCAN_IN), .A2(keyinput218), .B1(
        REG2_REG_25__SCAN_IN), .B2(keyinput132), .ZN(n4345) );
  OAI221_X1 U5010 ( .B1(REG2_REG_24__SCAN_IN), .B2(keyinput218), .C1(
        REG2_REG_25__SCAN_IN), .C2(keyinput132), .A(n4345), .ZN(n4346) );
  NOR4_X1 U5011 ( .A1(n4349), .A2(n4348), .A3(n4347), .A4(n4346), .ZN(n4379)
         );
  AOI22_X1 U5012 ( .A1(REG2_REG_27__SCAN_IN), .A2(keyinput199), .B1(
        REG2_REG_28__SCAN_IN), .B2(keyinput190), .ZN(n4350) );
  OAI221_X1 U5013 ( .B1(REG2_REG_27__SCAN_IN), .B2(keyinput199), .C1(
        REG2_REG_28__SCAN_IN), .C2(keyinput190), .A(n4350), .ZN(n4357) );
  AOI22_X1 U5014 ( .A1(ADDR_REG_16__SCAN_IN), .A2(keyinput233), .B1(
        REG2_REG_29__SCAN_IN), .B2(keyinput158), .ZN(n4351) );
  OAI221_X1 U5015 ( .B1(ADDR_REG_16__SCAN_IN), .B2(keyinput233), .C1(
        REG2_REG_29__SCAN_IN), .C2(keyinput158), .A(n4351), .ZN(n4356) );
  AOI22_X1 U5016 ( .A1(DATAO_REG_11__SCAN_IN), .A2(keyinput232), .B1(
        DATAO_REG_7__SCAN_IN), .B2(keyinput159), .ZN(n4352) );
  OAI221_X1 U5017 ( .B1(DATAO_REG_11__SCAN_IN), .B2(keyinput232), .C1(
        DATAO_REG_7__SCAN_IN), .C2(keyinput159), .A(n4352), .ZN(n4355) );
  AOI22_X1 U5018 ( .A1(DATAO_REG_18__SCAN_IN), .A2(keyinput211), .B1(
        DATAO_REG_13__SCAN_IN), .B2(keyinput235), .ZN(n4353) );
  OAI221_X1 U5019 ( .B1(DATAO_REG_18__SCAN_IN), .B2(keyinput211), .C1(
        DATAO_REG_13__SCAN_IN), .C2(keyinput235), .A(n4353), .ZN(n4354) );
  NOR4_X1 U5020 ( .A1(n4357), .A2(n4356), .A3(n4355), .A4(n4354), .ZN(n4378)
         );
  AOI22_X1 U5021 ( .A1(DATAO_REG_30__SCAN_IN), .A2(keyinput143), .B1(
        DATAO_REG_29__SCAN_IN), .B2(keyinput195), .ZN(n4358) );
  OAI221_X1 U5022 ( .B1(DATAO_REG_30__SCAN_IN), .B2(keyinput143), .C1(
        DATAO_REG_29__SCAN_IN), .C2(keyinput195), .A(n4358), .ZN(n4366) );
  AOI22_X1 U5023 ( .A1(REG3_REG_2__SCAN_IN), .A2(keyinput240), .B1(
        B_REG_SCAN_IN), .B2(keyinput168), .ZN(n4359) );
  OAI221_X1 U5024 ( .B1(REG3_REG_2__SCAN_IN), .B2(keyinput240), .C1(
        B_REG_SCAN_IN), .C2(keyinput168), .A(n4359), .ZN(n4365) );
  AOI22_X1 U5025 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput207), .B1(
        REG3_REG_25__SCAN_IN), .B2(keyinput197), .ZN(n4360) );
  OAI221_X1 U5026 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput207), .C1(
        REG3_REG_25__SCAN_IN), .C2(keyinput197), .A(n4360), .ZN(n4364) );
  INV_X1 U5027 ( .A(DATAI_25_), .ZN(n4527) );
  AOI22_X1 U5028 ( .A1(n4362), .A2(keyinput248), .B1(n4527), .B2(keyinput221), 
        .ZN(n4361) );
  OAI221_X1 U5029 ( .B1(n4362), .B2(keyinput248), .C1(n4527), .C2(keyinput221), 
        .A(n4361), .ZN(n4363) );
  NOR4_X1 U5030 ( .A1(n4366), .A2(n4365), .A3(n4364), .A4(n4363), .ZN(n4377)
         );
  INV_X1 U5031 ( .A(DATAI_18_), .ZN(n5012) );
  AOI22_X1 U5032 ( .A1(n5012), .A2(keyinput216), .B1(n4618), .B2(keyinput191), 
        .ZN(n4367) );
  OAI221_X1 U5033 ( .B1(n5012), .B2(keyinput216), .C1(n4618), .C2(keyinput191), 
        .A(n4367), .ZN(n4375) );
  INV_X1 U5034 ( .A(DATAI_10_), .ZN(n5027) );
  INV_X1 U5035 ( .A(DATAI_9_), .ZN(n4614) );
  AOI22_X1 U5036 ( .A1(n5027), .A2(keyinput201), .B1(n4614), .B2(keyinput210), 
        .ZN(n4368) );
  OAI221_X1 U5037 ( .B1(n5027), .B2(keyinput201), .C1(n4614), .C2(keyinput210), 
        .A(n4368), .ZN(n4374) );
  INV_X1 U5038 ( .A(DATAI_2_), .ZN(n4715) );
  INV_X1 U5039 ( .A(DATAI_0_), .ZN(n5037) );
  AOI22_X1 U5040 ( .A1(n4715), .A2(keyinput135), .B1(keyinput136), .B2(n5037), 
        .ZN(n4369) );
  OAI221_X1 U5041 ( .B1(n4715), .B2(keyinput135), .C1(n5037), .C2(keyinput136), 
        .A(n4369), .ZN(n4373) );
  AOI22_X1 U5042 ( .A1(n4371), .A2(keyinput145), .B1(n4628), .B2(keyinput167), 
        .ZN(n4370) );
  OAI221_X1 U5043 ( .B1(n4371), .B2(keyinput145), .C1(n4628), .C2(keyinput167), 
        .A(n4370), .ZN(n4372) );
  NOR4_X1 U5044 ( .A1(n4375), .A2(n4374), .A3(n4373), .A4(n4372), .ZN(n4376)
         );
  NAND4_X1 U5045 ( .A1(n4379), .A2(n4378), .A3(n4377), .A4(n4376), .ZN(n4487)
         );
  AOI22_X1 U5046 ( .A1(n4382), .A2(keyinput172), .B1(n4381), .B2(keyinput130), 
        .ZN(n4380) );
  OAI221_X1 U5047 ( .B1(n4382), .B2(keyinput172), .C1(n4381), .C2(keyinput130), 
        .A(n4380), .ZN(n4390) );
  AOI22_X1 U5048 ( .A1(n4547), .A2(keyinput161), .B1(keyinput134), .B2(n4384), 
        .ZN(n4383) );
  OAI221_X1 U5049 ( .B1(n4547), .B2(keyinput161), .C1(n4384), .C2(keyinput134), 
        .A(n4383), .ZN(n4389) );
  INV_X1 U5050 ( .A(REG2_REG_3__SCAN_IN), .ZN(n4500) );
  AOI22_X1 U5051 ( .A1(n4641), .A2(keyinput252), .B1(keyinput186), .B2(n4500), 
        .ZN(n4385) );
  OAI221_X1 U5052 ( .B1(n4641), .B2(keyinput252), .C1(n4500), .C2(keyinput186), 
        .A(n4385), .ZN(n4388) );
  INV_X1 U5053 ( .A(REG2_REG_6__SCAN_IN), .ZN(n4538) );
  AOI22_X1 U5054 ( .A1(n4538), .A2(keyinput245), .B1(keyinput219), .B2(n3481), 
        .ZN(n4386) );
  OAI221_X1 U5055 ( .B1(n4538), .B2(keyinput245), .C1(n3481), .C2(keyinput219), 
        .A(n4386), .ZN(n4387) );
  NOR4_X1 U5056 ( .A1(n4390), .A2(n4389), .A3(n4388), .A4(n4387), .ZN(n4428)
         );
  AOI22_X1 U5057 ( .A1(n3595), .A2(keyinput163), .B1(keyinput155), .B2(n4639), 
        .ZN(n4391) );
  OAI221_X1 U5058 ( .B1(n3595), .B2(keyinput163), .C1(n4639), .C2(keyinput155), 
        .A(n4391), .ZN(n4400) );
  INV_X1 U5059 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4393) );
  AOI22_X1 U5060 ( .A1(n4393), .A2(keyinput156), .B1(n4509), .B2(keyinput171), 
        .ZN(n4392) );
  OAI221_X1 U5061 ( .B1(n4393), .B2(keyinput156), .C1(n4509), .C2(keyinput171), 
        .A(n4392), .ZN(n4399) );
  INV_X1 U5062 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4643) );
  AOI22_X1 U5063 ( .A1(n4129), .A2(keyinput152), .B1(n4643), .B2(keyinput242), 
        .ZN(n4394) );
  OAI221_X1 U5064 ( .B1(n4129), .B2(keyinput152), .C1(n4643), .C2(keyinput242), 
        .A(n4394), .ZN(n4398) );
  INV_X1 U5065 ( .A(ADDR_REG_17__SCAN_IN), .ZN(n4540) );
  INV_X1 U5066 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4396) );
  AOI22_X1 U5067 ( .A1(n4540), .A2(keyinput183), .B1(keyinput249), .B2(n4396), 
        .ZN(n4395) );
  OAI221_X1 U5068 ( .B1(n4540), .B2(keyinput183), .C1(n4396), .C2(keyinput249), 
        .A(n4395), .ZN(n4397) );
  NOR4_X1 U5069 ( .A1(n4400), .A2(n4399), .A3(n4398), .A4(n4397), .ZN(n4427)
         );
  INV_X1 U5070 ( .A(ADDR_REG_9__SCAN_IN), .ZN(n4402) );
  INV_X1 U5071 ( .A(ADDR_REG_12__SCAN_IN), .ZN(n4541) );
  AOI22_X1 U5072 ( .A1(n4402), .A2(keyinput166), .B1(keyinput162), .B2(n4541), 
        .ZN(n4401) );
  OAI221_X1 U5073 ( .B1(n4402), .B2(keyinput166), .C1(n4541), .C2(keyinput162), 
        .A(n4401), .ZN(n4411) );
  INV_X1 U5074 ( .A(ADDR_REG_7__SCAN_IN), .ZN(n4537) );
  INV_X1 U5075 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n4404) );
  AOI22_X1 U5076 ( .A1(n4537), .A2(keyinput247), .B1(keyinput203), .B2(n4404), 
        .ZN(n4403) );
  OAI221_X1 U5077 ( .B1(n4537), .B2(keyinput247), .C1(n4404), .C2(keyinput203), 
        .A(n4403), .ZN(n4410) );
  INV_X1 U5078 ( .A(ADDR_REG_2__SCAN_IN), .ZN(n4535) );
  AOI22_X1 U5079 ( .A1(n4535), .A2(keyinput184), .B1(keyinput253), .B2(n4608), 
        .ZN(n4405) );
  OAI221_X1 U5080 ( .B1(n4535), .B2(keyinput184), .C1(n4608), .C2(keyinput253), 
        .A(n4405), .ZN(n4409) );
  AOI22_X1 U5081 ( .A1(n4407), .A2(keyinput205), .B1(keyinput181), .B2(n4522), 
        .ZN(n4406) );
  OAI221_X1 U5082 ( .B1(n4407), .B2(keyinput205), .C1(n4522), .C2(keyinput181), 
        .A(n4406), .ZN(n4408) );
  NOR4_X1 U5083 ( .A1(n4411), .A2(n4410), .A3(n4409), .A4(n4408), .ZN(n4426)
         );
  AOI22_X1 U5084 ( .A1(n4413), .A2(keyinput229), .B1(keyinput131), .B2(n4627), 
        .ZN(n4412) );
  OAI221_X1 U5085 ( .B1(n4413), .B2(keyinput229), .C1(n4627), .C2(keyinput131), 
        .A(n4412), .ZN(n4424) );
  AOI22_X1 U5086 ( .A1(n4416), .A2(keyinput226), .B1(n4415), .B2(keyinput176), 
        .ZN(n4414) );
  OAI221_X1 U5087 ( .B1(n4416), .B2(keyinput226), .C1(n4415), .C2(keyinput176), 
        .A(n4414), .ZN(n4423) );
  INV_X1 U5088 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4418) );
  AOI22_X1 U5089 ( .A1(n4515), .A2(keyinput157), .B1(n4418), .B2(keyinput193), 
        .ZN(n4417) );
  OAI221_X1 U5090 ( .B1(n4515), .B2(keyinput157), .C1(n4418), .C2(keyinput193), 
        .A(n4417), .ZN(n4422) );
  INV_X1 U5091 ( .A(ADDR_REG_19__SCAN_IN), .ZN(n4420) );
  AOI22_X1 U5092 ( .A1(n4420), .A2(keyinput223), .B1(n4550), .B2(keyinput202), 
        .ZN(n4419) );
  OAI221_X1 U5093 ( .B1(n4420), .B2(keyinput223), .C1(n4550), .C2(keyinput202), 
        .A(n4419), .ZN(n4421) );
  NOR4_X1 U5094 ( .A1(n4424), .A2(n4423), .A3(n4422), .A4(n4421), .ZN(n4425)
         );
  NAND4_X1 U5095 ( .A1(n4428), .A2(n4427), .A3(n4426), .A4(n4425), .ZN(n4486)
         );
  INV_X1 U5096 ( .A(D_REG_11__SCAN_IN), .ZN(n5004) );
  INV_X1 U5097 ( .A(D_REG_12__SCAN_IN), .ZN(n5003) );
  AOI22_X1 U5098 ( .A1(n5004), .A2(keyinput170), .B1(n5003), .B2(keyinput140), 
        .ZN(n4429) );
  OAI221_X1 U5099 ( .B1(n5004), .B2(keyinput170), .C1(n5003), .C2(keyinput140), 
        .A(n4429), .ZN(n4442) );
  INV_X1 U5100 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4601) );
  AOI22_X1 U5101 ( .A1(n4601), .A2(keyinput222), .B1(n4503), .B2(keyinput142), 
        .ZN(n4430) );
  OAI221_X1 U5102 ( .B1(n4601), .B2(keyinput222), .C1(n4503), .C2(keyinput142), 
        .A(n4430), .ZN(n4441) );
  XNOR2_X1 U5103 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput255), .ZN(n4434) );
  XNOR2_X1 U5104 ( .A(IR_REG_17__SCAN_IN), .B(keyinput187), .ZN(n4433) );
  XNOR2_X1 U5105 ( .A(IR_REG_9__SCAN_IN), .B(keyinput173), .ZN(n4432) );
  XNOR2_X1 U5106 ( .A(IR_REG_23__SCAN_IN), .B(keyinput133), .ZN(n4431) );
  NAND4_X1 U5107 ( .A1(n4434), .A2(n4433), .A3(n4432), .A4(n4431), .ZN(n4440)
         );
  XNOR2_X1 U5108 ( .A(IR_REG_21__SCAN_IN), .B(keyinput244), .ZN(n4438) );
  XNOR2_X1 U5109 ( .A(IR_REG_27__SCAN_IN), .B(keyinput227), .ZN(n4437) );
  XNOR2_X1 U5110 ( .A(IR_REG_26__SCAN_IN), .B(keyinput213), .ZN(n4436) );
  XNOR2_X1 U5111 ( .A(IR_REG_28__SCAN_IN), .B(keyinput204), .ZN(n4435) );
  NAND4_X1 U5112 ( .A1(n4438), .A2(n4437), .A3(n4436), .A4(n4435), .ZN(n4439)
         );
  OR4_X1 U5113 ( .A1(n4442), .A2(n4441), .A3(n4440), .A4(n4439), .ZN(n4484) );
  AOI22_X1 U5114 ( .A1(DATAI_23_), .A2(keyinput146), .B1(DATAI_28_), .B2(
        keyinput189), .ZN(n4443) );
  OAI221_X1 U5115 ( .B1(DATAI_23_), .B2(keyinput146), .C1(DATAI_28_), .C2(
        keyinput189), .A(n4443), .ZN(n4450) );
  AOI22_X1 U5116 ( .A1(DATAI_15_), .A2(keyinput198), .B1(DATAI_17_), .B2(
        keyinput141), .ZN(n4444) );
  OAI221_X1 U5117 ( .B1(DATAI_15_), .B2(keyinput198), .C1(DATAI_17_), .C2(
        keyinput141), .A(n4444), .ZN(n4449) );
  AOI22_X1 U5118 ( .A1(DATAI_1_), .A2(keyinput150), .B1(REG3_REG_28__SCAN_IN), 
        .B2(keyinput149), .ZN(n4445) );
  OAI221_X1 U5119 ( .B1(DATAI_1_), .B2(keyinput150), .C1(REG3_REG_28__SCAN_IN), 
        .C2(keyinput149), .A(n4445), .ZN(n4448) );
  AOI22_X1 U5120 ( .A1(REG3_REG_10__SCAN_IN), .A2(keyinput148), .B1(
        REG3_REG_12__SCAN_IN), .B2(keyinput174), .ZN(n4446) );
  OAI221_X1 U5121 ( .B1(REG3_REG_10__SCAN_IN), .B2(keyinput148), .C1(
        REG3_REG_12__SCAN_IN), .C2(keyinput174), .A(n4446), .ZN(n4447) );
  NOR4_X1 U5122 ( .A1(n4450), .A2(n4449), .A3(n4448), .A4(n4447), .ZN(n4478)
         );
  AOI22_X1 U5123 ( .A1(REG3_REG_20__SCAN_IN), .A2(keyinput169), .B1(
        IR_REG_0__SCAN_IN), .B2(keyinput196), .ZN(n4451) );
  OAI221_X1 U5124 ( .B1(REG3_REG_20__SCAN_IN), .B2(keyinput169), .C1(
        IR_REG_0__SCAN_IN), .C2(keyinput196), .A(n4451), .ZN(n4458) );
  AOI22_X1 U5125 ( .A1(IR_REG_6__SCAN_IN), .A2(keyinput238), .B1(
        IR_REG_14__SCAN_IN), .B2(keyinput179), .ZN(n4452) );
  OAI221_X1 U5126 ( .B1(IR_REG_6__SCAN_IN), .B2(keyinput238), .C1(
        IR_REG_14__SCAN_IN), .C2(keyinput179), .A(n4452), .ZN(n4457) );
  AOI22_X1 U5127 ( .A1(D_REG_2__SCAN_IN), .A2(keyinput217), .B1(
        D_REG_5__SCAN_IN), .B2(keyinput137), .ZN(n4453) );
  OAI221_X1 U5128 ( .B1(D_REG_2__SCAN_IN), .B2(keyinput217), .C1(
        D_REG_5__SCAN_IN), .C2(keyinput137), .A(n4453), .ZN(n4456) );
  AOI22_X1 U5129 ( .A1(D_REG_10__SCAN_IN), .A2(keyinput234), .B1(
        D_REG_7__SCAN_IN), .B2(keyinput239), .ZN(n4454) );
  OAI221_X1 U5130 ( .B1(D_REG_10__SCAN_IN), .B2(keyinput234), .C1(
        D_REG_7__SCAN_IN), .C2(keyinput239), .A(n4454), .ZN(n4455) );
  NOR4_X1 U5131 ( .A1(n4458), .A2(n4457), .A3(n4456), .A4(n4455), .ZN(n4477)
         );
  AOI22_X1 U5132 ( .A1(D_REG_13__SCAN_IN), .A2(keyinput178), .B1(
        D_REG_14__SCAN_IN), .B2(keyinput164), .ZN(n4459) );
  OAI221_X1 U5133 ( .B1(D_REG_13__SCAN_IN), .B2(keyinput178), .C1(
        D_REG_14__SCAN_IN), .C2(keyinput164), .A(n4459), .ZN(n4466) );
  AOI22_X1 U5134 ( .A1(REG0_REG_0__SCAN_IN), .A2(keyinput128), .B1(
        D_REG_29__SCAN_IN), .B2(keyinput231), .ZN(n4460) );
  OAI221_X1 U5135 ( .B1(REG0_REG_0__SCAN_IN), .B2(keyinput128), .C1(
        D_REG_29__SCAN_IN), .C2(keyinput231), .A(n4460), .ZN(n4465) );
  AOI22_X1 U5136 ( .A1(REG0_REG_1__SCAN_IN), .A2(keyinput200), .B1(
        REG0_REG_8__SCAN_IN), .B2(keyinput228), .ZN(n4461) );
  OAI221_X1 U5137 ( .B1(REG0_REG_1__SCAN_IN), .B2(keyinput200), .C1(
        REG0_REG_8__SCAN_IN), .C2(keyinput228), .A(n4461), .ZN(n4464) );
  AOI22_X1 U5138 ( .A1(REG0_REG_11__SCAN_IN), .A2(keyinput180), .B1(
        REG0_REG_10__SCAN_IN), .B2(keyinput165), .ZN(n4462) );
  OAI221_X1 U5139 ( .B1(REG0_REG_11__SCAN_IN), .B2(keyinput180), .C1(
        REG0_REG_10__SCAN_IN), .C2(keyinput165), .A(n4462), .ZN(n4463) );
  NOR4_X1 U5140 ( .A1(n4466), .A2(n4465), .A3(n4464), .A4(n4463), .ZN(n4476)
         );
  AOI22_X1 U5141 ( .A1(REG0_REG_13__SCAN_IN), .A2(keyinput192), .B1(
        REG0_REG_16__SCAN_IN), .B2(keyinput220), .ZN(n4467) );
  OAI221_X1 U5142 ( .B1(REG0_REG_13__SCAN_IN), .B2(keyinput192), .C1(
        REG0_REG_16__SCAN_IN), .C2(keyinput220), .A(n4467), .ZN(n4474) );
  AOI22_X1 U5143 ( .A1(REG1_REG_0__SCAN_IN), .A2(keyinput177), .B1(
        REG0_REG_25__SCAN_IN), .B2(keyinput154), .ZN(n4468) );
  OAI221_X1 U5144 ( .B1(REG1_REG_0__SCAN_IN), .B2(keyinput177), .C1(
        REG0_REG_25__SCAN_IN), .C2(keyinput154), .A(n4468), .ZN(n4473) );
  AOI22_X1 U5145 ( .A1(REG1_REG_7__SCAN_IN), .A2(keyinput188), .B1(
        REG0_REG_28__SCAN_IN), .B2(keyinput246), .ZN(n4469) );
  OAI221_X1 U5146 ( .B1(REG1_REG_7__SCAN_IN), .B2(keyinput188), .C1(
        REG0_REG_28__SCAN_IN), .C2(keyinput246), .A(n4469), .ZN(n4472) );
  AOI22_X1 U5147 ( .A1(REG1_REG_10__SCAN_IN), .A2(keyinput175), .B1(
        REG1_REG_8__SCAN_IN), .B2(keyinput209), .ZN(n4470) );
  OAI221_X1 U5148 ( .B1(REG1_REG_10__SCAN_IN), .B2(keyinput175), .C1(
        REG1_REG_8__SCAN_IN), .C2(keyinput209), .A(n4470), .ZN(n4471) );
  NOR4_X1 U5149 ( .A1(n4474), .A2(n4473), .A3(n4472), .A4(n4471), .ZN(n4475)
         );
  NAND4_X1 U5150 ( .A1(n4478), .A2(n4477), .A3(n4476), .A4(n4475), .ZN(n4483)
         );
  INV_X1 U5151 ( .A(D_REG_4__SCAN_IN), .ZN(n5006) );
  AOI22_X1 U5152 ( .A1(n3169), .A2(keyinput230), .B1(keyinput160), .B2(n5006), 
        .ZN(n4479) );
  OAI221_X1 U5153 ( .B1(n3169), .B2(keyinput230), .C1(n5006), .C2(keyinput160), 
        .A(n4479), .ZN(n4482) );
  AOI22_X1 U5154 ( .A1(n2459), .A2(keyinput250), .B1(keyinput241), .B2(n2771), 
        .ZN(n4480) );
  OAI221_X1 U5155 ( .B1(n2459), .B2(keyinput250), .C1(n2771), .C2(keyinput241), 
        .A(n4480), .ZN(n4481) );
  OR4_X1 U5156 ( .A1(n4484), .A2(n4483), .A3(n4482), .A4(n4481), .ZN(n4485) );
  NOR4_X1 U5157 ( .A1(n4488), .A2(n4487), .A3(n4486), .A4(n4485), .ZN(n4563)
         );
  AOI22_X1 U5158 ( .A1(n4325), .A2(keyinput254), .B1(n4490), .B2(keyinput236), 
        .ZN(n4489) );
  OAI221_X1 U5159 ( .B1(n4325), .B2(keyinput254), .C1(n4490), .C2(keyinput236), 
        .A(n4489), .ZN(n4498) );
  AOI22_X1 U5160 ( .A1(n4302), .A2(keyinput251), .B1(keyinput237), .B2(n5076), 
        .ZN(n4491) );
  OAI221_X1 U5161 ( .B1(n4302), .B2(keyinput251), .C1(n5076), .C2(keyinput237), 
        .A(n4491), .ZN(n4497) );
  AOI22_X1 U5162 ( .A1(n4493), .A2(keyinput212), .B1(keyinput224), .B2(n2305), 
        .ZN(n4492) );
  OAI221_X1 U5163 ( .B1(n4493), .B2(keyinput212), .C1(n2305), .C2(keyinput224), 
        .A(n4492), .ZN(n4496) );
  AOI22_X1 U5164 ( .A1(n5082), .A2(keyinput153), .B1(n4605), .B2(keyinput144), 
        .ZN(n4494) );
  OAI221_X1 U5165 ( .B1(n5082), .B2(keyinput153), .C1(n4605), .C2(keyinput144), 
        .A(n4494), .ZN(n4495) );
  NOR4_X1 U5166 ( .A1(n4498), .A2(n4497), .A3(n4496), .A4(n4495), .ZN(n4562)
         );
  INV_X1 U5167 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4501) );
  AOI22_X1 U5168 ( .A1(n4501), .A2(keyinput4), .B1(keyinput58), .B2(n4500), 
        .ZN(n4499) );
  OAI221_X1 U5169 ( .B1(n4501), .B2(keyinput4), .C1(n4500), .C2(keyinput58), 
        .A(n4499), .ZN(n4513) );
  AOI22_X1 U5170 ( .A1(n4504), .A2(keyinput21), .B1(keyinput14), .B2(n4503), 
        .ZN(n4502) );
  OAI221_X1 U5171 ( .B1(n4504), .B2(keyinput21), .C1(n4503), .C2(keyinput14), 
        .A(n4502), .ZN(n4512) );
  INV_X1 U5172 ( .A(B_REG_SCAN_IN), .ZN(n4507) );
  INV_X1 U5173 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4506) );
  AOI22_X1 U5174 ( .A1(n4507), .A2(keyinput40), .B1(keyinput90), .B2(n4506), 
        .ZN(n4505) );
  OAI221_X1 U5175 ( .B1(n4507), .B2(keyinput40), .C1(n4506), .C2(keyinput90), 
        .A(n4505), .ZN(n4511) );
  AOI22_X1 U5176 ( .A1(n4129), .A2(keyinput24), .B1(keyinput43), .B2(n4509), 
        .ZN(n4508) );
  OAI221_X1 U5177 ( .B1(n4129), .B2(keyinput24), .C1(n4509), .C2(keyinput43), 
        .A(n4508), .ZN(n4510) );
  NOR4_X1 U5178 ( .A1(n4513), .A2(n4512), .A3(n4511), .A4(n4510), .ZN(n4531)
         );
  AOI22_X1 U5179 ( .A1(n4516), .A2(keyinput57), .B1(n4515), .B2(keyinput29), 
        .ZN(n4514) );
  OAI221_X1 U5180 ( .B1(n4516), .B2(keyinput57), .C1(n4515), .C2(keyinput29), 
        .A(n4514), .ZN(n4517) );
  INV_X1 U5181 ( .A(n4517), .ZN(n4520) );
  XNOR2_X1 U5182 ( .A(keyinput17), .B(REG3_REG_7__SCAN_IN), .ZN(n4519) );
  XNOR2_X1 U5183 ( .A(IR_REG_23__SCAN_IN), .B(keyinput5), .ZN(n4518) );
  NAND3_X1 U5184 ( .A1(n4520), .A2(n4519), .A3(n4518), .ZN(n4525) );
  INV_X1 U5185 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4523) );
  AOI22_X1 U5186 ( .A1(n4523), .A2(keyinput81), .B1(keyinput53), .B2(n4522), 
        .ZN(n4521) );
  OAI221_X1 U5187 ( .B1(n4523), .B2(keyinput81), .C1(n4522), .C2(keyinput53), 
        .A(n4521), .ZN(n4524) );
  NOR2_X1 U5188 ( .A1(n4525), .A2(n4524), .ZN(n4530) );
  AOI22_X1 U5189 ( .A1(n4527), .A2(keyinput93), .B1(keyinput73), .B2(n5027), 
        .ZN(n4526) );
  OAI221_X1 U5190 ( .B1(n4527), .B2(keyinput93), .C1(n5027), .C2(keyinput73), 
        .A(n4526), .ZN(n4528) );
  INV_X1 U5191 ( .A(n4528), .ZN(n4529) );
  NAND3_X1 U5192 ( .A1(n4531), .A2(n4530), .A3(n4529), .ZN(n4561) );
  AOI22_X1 U5193 ( .A1(n3595), .A2(keyinput35), .B1(keyinput112), .B2(n4533), 
        .ZN(n4532) );
  OAI221_X1 U5194 ( .B1(n3595), .B2(keyinput35), .C1(n4533), .C2(keyinput112), 
        .A(n4532), .ZN(n4545) );
  AOI22_X1 U5195 ( .A1(n4535), .A2(keyinput56), .B1(n5038), .B2(keyinput68), 
        .ZN(n4534) );
  OAI221_X1 U5196 ( .B1(n4535), .B2(keyinput56), .C1(n5038), .C2(keyinput68), 
        .A(n4534), .ZN(n4544) );
  AOI22_X1 U5197 ( .A1(n4538), .A2(keyinput117), .B1(keyinput119), .B2(n4537), 
        .ZN(n4536) );
  OAI221_X1 U5198 ( .B1(n4538), .B2(keyinput117), .C1(n4537), .C2(keyinput119), 
        .A(n4536), .ZN(n4543) );
  AOI22_X1 U5199 ( .A1(n4541), .A2(keyinput34), .B1(n4540), .B2(keyinput55), 
        .ZN(n4539) );
  OAI221_X1 U5200 ( .B1(n4541), .B2(keyinput34), .C1(n4540), .C2(keyinput55), 
        .A(n4539), .ZN(n4542) );
  NOR4_X1 U5201 ( .A1(n4545), .A2(n4544), .A3(n4543), .A4(n4542), .ZN(n4559)
         );
  AOI22_X1 U5202 ( .A1(n4309), .A2(keyinput26), .B1(n4547), .B2(keyinput33), 
        .ZN(n4546) );
  OAI221_X1 U5203 ( .B1(n4309), .B2(keyinput26), .C1(n4547), .C2(keyinput33), 
        .A(n4546), .ZN(n4557) );
  AOI22_X1 U5204 ( .A1(n4550), .A2(keyinput74), .B1(n4549), .B2(keyinput118), 
        .ZN(n4548) );
  OAI221_X1 U5205 ( .B1(n4550), .B2(keyinput74), .C1(n4549), .C2(keyinput118), 
        .A(n4548), .ZN(n4556) );
  INV_X1 U5206 ( .A(REG0_REG_0__SCAN_IN), .ZN(n5045) );
  AOI22_X1 U5207 ( .A1(n2459), .A2(keyinput122), .B1(keyinput0), .B2(n5045), 
        .ZN(n4551) );
  OAI221_X1 U5208 ( .B1(n2459), .B2(keyinput122), .C1(n5045), .C2(keyinput0), 
        .A(n4551), .ZN(n4555) );
  INV_X1 U5209 ( .A(D_REG_29__SCAN_IN), .ZN(n4998) );
  AOI22_X1 U5210 ( .A1(n4553), .A2(keyinput127), .B1(n4998), .B2(keyinput103), 
        .ZN(n4552) );
  OAI221_X1 U5211 ( .B1(n4553), .B2(keyinput127), .C1(n4998), .C2(keyinput103), 
        .A(n4552), .ZN(n4554) );
  NOR4_X1 U5212 ( .A1(n4557), .A2(n4556), .A3(n4555), .A4(n4554), .ZN(n4558)
         );
  NAND2_X1 U5213 ( .A1(n4559), .A2(n4558), .ZN(n4560) );
  AOI211_X1 U5214 ( .C1(n4563), .C2(n4562), .A(n4561), .B(n4560), .ZN(n4691)
         );
  OAI22_X1 U5215 ( .A1(REG1_REG_27__SCAN_IN), .A2(keyinput19), .B1(DATAI_30_), 
        .B2(keyinput120), .ZN(n4564) );
  AOI221_X1 U5216 ( .B1(REG1_REG_27__SCAN_IN), .B2(keyinput19), .C1(
        keyinput120), .C2(DATAI_30_), .A(n4564), .ZN(n4571) );
  OAI22_X1 U5217 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput65), .B1(
        REG3_REG_20__SCAN_IN), .B2(keyinput41), .ZN(n4565) );
  AOI221_X1 U5218 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput65), .C1(keyinput41), .C2(REG3_REG_20__SCAN_IN), .A(n4565), .ZN(n4570) );
  OAI22_X1 U5219 ( .A1(REG1_REG_0__SCAN_IN), .A2(keyinput49), .B1(
        REG1_REG_4__SCAN_IN), .B2(keyinput96), .ZN(n4566) );
  AOI221_X1 U5220 ( .B1(REG1_REG_0__SCAN_IN), .B2(keyinput49), .C1(keyinput96), 
        .C2(REG1_REG_4__SCAN_IN), .A(n4566), .ZN(n4569) );
  OAI22_X1 U5221 ( .A1(DATAI_28_), .A2(keyinput61), .B1(REG0_REG_16__SCAN_IN), 
        .B2(keyinput92), .ZN(n4567) );
  AOI221_X1 U5222 ( .B1(DATAI_28_), .B2(keyinput61), .C1(keyinput92), .C2(
        REG0_REG_16__SCAN_IN), .A(n4567), .ZN(n4568) );
  NAND4_X1 U5223 ( .A1(n4571), .A2(n4570), .A3(n4569), .A4(n4568), .ZN(n4599)
         );
  OAI22_X1 U5224 ( .A1(REG2_REG_28__SCAN_IN), .A2(keyinput62), .B1(
        REG2_REG_27__SCAN_IN), .B2(keyinput71), .ZN(n4572) );
  AOI221_X1 U5225 ( .B1(REG2_REG_28__SCAN_IN), .B2(keyinput62), .C1(keyinput71), .C2(REG2_REG_27__SCAN_IN), .A(n4572), .ZN(n4579) );
  OAI22_X1 U5226 ( .A1(REG3_REG_25__SCAN_IN), .A2(keyinput69), .B1(
        ADDR_REG_19__SCAN_IN), .B2(keyinput95), .ZN(n4573) );
  AOI221_X1 U5227 ( .B1(REG3_REG_25__SCAN_IN), .B2(keyinput69), .C1(keyinput95), .C2(ADDR_REG_19__SCAN_IN), .A(n4573), .ZN(n4578) );
  OAI22_X1 U5228 ( .A1(REG2_REG_29__SCAN_IN), .A2(keyinput30), .B1(keyinput31), 
        .B2(DATAO_REG_7__SCAN_IN), .ZN(n4574) );
  AOI221_X1 U5229 ( .B1(REG2_REG_29__SCAN_IN), .B2(keyinput30), .C1(
        DATAO_REG_7__SCAN_IN), .C2(keyinput31), .A(n4574), .ZN(n4577) );
  OAI22_X1 U5230 ( .A1(REG2_REG_19__SCAN_IN), .A2(keyinput28), .B1(keyinput115), .B2(REG1_REG_18__SCAN_IN), .ZN(n4575) );
  AOI221_X1 U5231 ( .B1(REG2_REG_19__SCAN_IN), .B2(keyinput28), .C1(
        REG1_REG_18__SCAN_IN), .C2(keyinput115), .A(n4575), .ZN(n4576) );
  NAND4_X1 U5232 ( .A1(n4579), .A2(n4578), .A3(n4577), .A4(n4576), .ZN(n4598)
         );
  OAI22_X1 U5233 ( .A1(D_REG_7__SCAN_IN), .A2(keyinput111), .B1(
        D_REG_5__SCAN_IN), .B2(keyinput9), .ZN(n4580) );
  AOI221_X1 U5234 ( .B1(D_REG_7__SCAN_IN), .B2(keyinput111), .C1(keyinput9), 
        .C2(D_REG_5__SCAN_IN), .A(n4580), .ZN(n4587) );
  OAI22_X1 U5235 ( .A1(D_REG_14__SCAN_IN), .A2(keyinput36), .B1(
        D_REG_13__SCAN_IN), .B2(keyinput50), .ZN(n4581) );
  AOI221_X1 U5236 ( .B1(D_REG_14__SCAN_IN), .B2(keyinput36), .C1(keyinput50), 
        .C2(D_REG_13__SCAN_IN), .A(n4581), .ZN(n4586) );
  OAI22_X1 U5237 ( .A1(REG0_REG_10__SCAN_IN), .A2(keyinput37), .B1(
        REG0_REG_11__SCAN_IN), .B2(keyinput52), .ZN(n4582) );
  AOI221_X1 U5238 ( .B1(REG0_REG_10__SCAN_IN), .B2(keyinput37), .C1(keyinput52), .C2(REG0_REG_11__SCAN_IN), .A(n4582), .ZN(n4585) );
  OAI22_X1 U5239 ( .A1(DATAI_23_), .A2(keyinput18), .B1(REG0_REG_8__SCAN_IN), 
        .B2(keyinput100), .ZN(n4583) );
  AOI221_X1 U5240 ( .B1(DATAI_23_), .B2(keyinput18), .C1(keyinput100), .C2(
        REG0_REG_8__SCAN_IN), .A(n4583), .ZN(n4584) );
  NAND4_X1 U5241 ( .A1(n4587), .A2(n4586), .A3(n4585), .A4(n4584), .ZN(n4597)
         );
  OAI22_X1 U5242 ( .A1(REG1_REG_15__SCAN_IN), .A2(keyinput44), .B1(keyinput105), .B2(ADDR_REG_16__SCAN_IN), .ZN(n4588) );
  AOI221_X1 U5243 ( .B1(REG1_REG_15__SCAN_IN), .B2(keyinput44), .C1(
        ADDR_REG_16__SCAN_IN), .C2(keyinput105), .A(n4588), .ZN(n4595) );
  OAI22_X1 U5244 ( .A1(REG2_REG_8__SCAN_IN), .A2(keyinput1), .B1(
        ADDR_REG_9__SCAN_IN), .B2(keyinput38), .ZN(n4589) );
  AOI221_X1 U5245 ( .B1(REG2_REG_8__SCAN_IN), .B2(keyinput1), .C1(keyinput38), 
        .C2(ADDR_REG_9__SCAN_IN), .A(n4589), .ZN(n4594) );
  OAI22_X1 U5246 ( .A1(REG2_REG_7__SCAN_IN), .A2(keyinput54), .B1(
        REG2_REG_11__SCAN_IN), .B2(keyinput91), .ZN(n4590) );
  AOI221_X1 U5247 ( .B1(REG2_REG_7__SCAN_IN), .B2(keyinput54), .C1(keyinput91), 
        .C2(REG2_REG_11__SCAN_IN), .A(n4590), .ZN(n4593) );
  OAI22_X1 U5248 ( .A1(REG1_REG_2__SCAN_IN), .A2(keyinput84), .B1(
        REG2_REG_1__SCAN_IN), .B2(keyinput6), .ZN(n4591) );
  AOI221_X1 U5249 ( .B1(REG1_REG_2__SCAN_IN), .B2(keyinput84), .C1(keyinput6), 
        .C2(REG2_REG_1__SCAN_IN), .A(n4591), .ZN(n4592) );
  NAND4_X1 U5250 ( .A1(n4595), .A2(n4594), .A3(n4593), .A4(n4592), .ZN(n4596)
         );
  NOR4_X1 U5251 ( .A1(n4599), .A2(n4598), .A3(n4597), .A4(n4596), .ZN(n4690)
         );
  INV_X1 U5252 ( .A(D_REG_10__SCAN_IN), .ZN(n5005) );
  AOI22_X1 U5253 ( .A1(n4601), .A2(keyinput94), .B1(n5005), .B2(keyinput106), 
        .ZN(n4600) );
  OAI221_X1 U5254 ( .B1(n4601), .B2(keyinput94), .C1(n5005), .C2(keyinput106), 
        .A(n4600), .ZN(n4612) );
  AOI22_X1 U5255 ( .A1(n4603), .A2(keyinput107), .B1(n5003), .B2(keyinput12), 
        .ZN(n4602) );
  OAI221_X1 U5256 ( .B1(n4603), .B2(keyinput107), .C1(n5003), .C2(keyinput12), 
        .A(n4602), .ZN(n4611) );
  AOI22_X1 U5257 ( .A1(n4606), .A2(keyinput20), .B1(keyinput16), .B2(n4605), 
        .ZN(n4604) );
  OAI221_X1 U5258 ( .B1(n4606), .B2(keyinput20), .C1(n4605), .C2(keyinput16), 
        .A(n4604), .ZN(n4610) );
  AOI22_X1 U5259 ( .A1(n2771), .A2(keyinput113), .B1(keyinput125), .B2(n4608), 
        .ZN(n4607) );
  OAI221_X1 U5260 ( .B1(n2771), .B2(keyinput113), .C1(n4608), .C2(keyinput125), 
        .A(n4607), .ZN(n4609) );
  NOR4_X1 U5261 ( .A1(n4612), .A2(n4611), .A3(n4610), .A4(n4609), .ZN(n4651)
         );
  AOI22_X1 U5262 ( .A1(n4763), .A2(keyinput86), .B1(n4614), .B2(keyinput82), 
        .ZN(n4613) );
  OAI221_X1 U5263 ( .B1(n4763), .B2(keyinput86), .C1(n4614), .C2(keyinput82), 
        .A(n4613), .ZN(n4623) );
  AOI22_X1 U5264 ( .A1(n4616), .A2(keyinput79), .B1(keyinput46), .B2(n2701), 
        .ZN(n4615) );
  OAI221_X1 U5265 ( .B1(n4616), .B2(keyinput79), .C1(n2701), .C2(keyinput46), 
        .A(n4615), .ZN(n4622) );
  AOI22_X1 U5266 ( .A1(n5004), .A2(keyinput42), .B1(keyinput63), .B2(n4618), 
        .ZN(n4617) );
  OAI221_X1 U5267 ( .B1(n5004), .B2(keyinput42), .C1(n4618), .C2(keyinput63), 
        .A(n4617), .ZN(n4621) );
  INV_X1 U5268 ( .A(D_REG_2__SCAN_IN), .ZN(n5008) );
  AOI22_X1 U5269 ( .A1(n5000), .A2(keyinput97), .B1(keyinput89), .B2(n5008), 
        .ZN(n4619) );
  OAI221_X1 U5270 ( .B1(n5000), .B2(keyinput97), .C1(n5008), .C2(keyinput89), 
        .A(n4619), .ZN(n4620) );
  NOR4_X1 U5271 ( .A1(n4623), .A2(n4622), .A3(n4621), .A4(n4620), .ZN(n4650)
         );
  INV_X1 U5272 ( .A(REG0_REG_1__SCAN_IN), .ZN(n5051) );
  AOI22_X1 U5273 ( .A1(n5051), .A2(keyinput72), .B1(keyinput104), .B2(n4625), 
        .ZN(n4624) );
  OAI221_X1 U5274 ( .B1(n5051), .B2(keyinput72), .C1(n4625), .C2(keyinput104), 
        .A(n4624), .ZN(n4636) );
  AOI22_X1 U5275 ( .A1(n4628), .A2(keyinput39), .B1(keyinput3), .B2(n4627), 
        .ZN(n4626) );
  OAI221_X1 U5276 ( .B1(n4628), .B2(keyinput39), .C1(n4627), .C2(keyinput3), 
        .A(n4626), .ZN(n4635) );
  AOI22_X1 U5277 ( .A1(n5001), .A2(keyinput23), .B1(keyinput15), .B2(n4630), 
        .ZN(n4629) );
  OAI221_X1 U5278 ( .B1(n5001), .B2(keyinput23), .C1(n4630), .C2(keyinput15), 
        .A(n4629), .ZN(n4634) );
  INV_X1 U5279 ( .A(DATAI_15_), .ZN(n5017) );
  AOI22_X1 U5280 ( .A1(n5017), .A2(keyinput70), .B1(n4632), .B2(keyinput66), 
        .ZN(n4631) );
  OAI221_X1 U5281 ( .B1(n5017), .B2(keyinput70), .C1(n4632), .C2(keyinput66), 
        .A(n4631), .ZN(n4633) );
  NOR4_X1 U5282 ( .A1(n4636), .A2(n4635), .A3(n4634), .A4(n4633), .ZN(n4649)
         );
  AOI22_X1 U5283 ( .A1(n5082), .A2(keyinput25), .B1(n5079), .B2(keyinput60), 
        .ZN(n4637) );
  OAI221_X1 U5284 ( .B1(n5082), .B2(keyinput25), .C1(n5079), .C2(keyinput60), 
        .A(n4637), .ZN(n4647) );
  AOI22_X1 U5285 ( .A1(n5076), .A2(keyinput109), .B1(keyinput27), .B2(n4639), 
        .ZN(n4638) );
  OAI221_X1 U5286 ( .B1(n5076), .B2(keyinput109), .C1(n4639), .C2(keyinput27), 
        .A(n4638), .ZN(n4646) );
  AOI22_X1 U5287 ( .A1(n4899), .A2(keyinput80), .B1(n4641), .B2(keyinput124), 
        .ZN(n4640) );
  OAI221_X1 U5288 ( .B1(n4899), .B2(keyinput80), .C1(n4641), .C2(keyinput124), 
        .A(n4640), .ZN(n4645) );
  AOI22_X1 U5289 ( .A1(n4325), .A2(keyinput126), .B1(n4643), .B2(keyinput114), 
        .ZN(n4642) );
  OAI221_X1 U5290 ( .B1(n4325), .B2(keyinput126), .C1(n4643), .C2(keyinput114), 
        .A(n4642), .ZN(n4644) );
  NOR4_X1 U5291 ( .A1(n4647), .A2(n4646), .A3(n4645), .A4(n4644), .ZN(n4648)
         );
  AND4_X1 U5292 ( .A1(n4651), .A2(n4650), .A3(n4649), .A4(n4648), .ZN(n4689)
         );
  OAI22_X1 U5293 ( .A1(IR_REG_9__SCAN_IN), .A2(keyinput45), .B1(keyinput77), 
        .B2(DATAO_REG_12__SCAN_IN), .ZN(n4652) );
  AOI221_X1 U5294 ( .B1(IR_REG_9__SCAN_IN), .B2(keyinput45), .C1(
        DATAO_REG_12__SCAN_IN), .C2(keyinput77), .A(n4652), .ZN(n4659) );
  OAI22_X1 U5295 ( .A1(IR_REG_26__SCAN_IN), .A2(keyinput85), .B1(keyinput101), 
        .B2(DATAO_REG_23__SCAN_IN), .ZN(n4653) );
  AOI221_X1 U5296 ( .B1(IR_REG_26__SCAN_IN), .B2(keyinput85), .C1(
        DATAO_REG_23__SCAN_IN), .C2(keyinput101), .A(n4653), .ZN(n4658) );
  OAI22_X1 U5297 ( .A1(IR_REG_28__SCAN_IN), .A2(keyinput76), .B1(keyinput88), 
        .B2(DATAI_18_), .ZN(n4654) );
  AOI221_X1 U5298 ( .B1(IR_REG_28__SCAN_IN), .B2(keyinput76), .C1(DATAI_18_), 
        .C2(keyinput88), .A(n4654), .ZN(n4657) );
  OAI22_X1 U5299 ( .A1(IR_REG_21__SCAN_IN), .A2(keyinput116), .B1(keyinput13), 
        .B2(DATAI_17_), .ZN(n4655) );
  AOI221_X1 U5300 ( .B1(IR_REG_21__SCAN_IN), .B2(keyinput116), .C1(DATAI_17_), 
        .C2(keyinput13), .A(n4655), .ZN(n4656) );
  NAND4_X1 U5301 ( .A1(n4659), .A2(n4658), .A3(n4657), .A4(n4656), .ZN(n4687)
         );
  OAI22_X1 U5302 ( .A1(REG0_REG_26__SCAN_IN), .A2(keyinput108), .B1(keyinput83), .B2(DATAO_REG_18__SCAN_IN), .ZN(n4660) );
  AOI221_X1 U5303 ( .B1(REG0_REG_26__SCAN_IN), .B2(keyinput108), .C1(
        DATAO_REG_18__SCAN_IN), .C2(keyinput83), .A(n4660), .ZN(n4667) );
  OAI22_X1 U5304 ( .A1(REG1_REG_10__SCAN_IN), .A2(keyinput47), .B1(keyinput64), 
        .B2(REG0_REG_13__SCAN_IN), .ZN(n4661) );
  AOI221_X1 U5305 ( .B1(REG1_REG_10__SCAN_IN), .B2(keyinput47), .C1(
        REG0_REG_13__SCAN_IN), .C2(keyinput64), .A(n4661), .ZN(n4666) );
  OAI22_X1 U5306 ( .A1(DATAI_0_), .A2(keyinput8), .B1(ADDR_REG_13__SCAN_IN), 
        .B2(keyinput121), .ZN(n4662) );
  AOI221_X1 U5307 ( .B1(DATAI_0_), .B2(keyinput8), .C1(keyinput121), .C2(
        ADDR_REG_13__SCAN_IN), .A(n4662), .ZN(n4665) );
  OAI22_X1 U5308 ( .A1(REG0_REG_27__SCAN_IN), .A2(keyinput123), .B1(
        DATAO_REG_29__SCAN_IN), .B2(keyinput67), .ZN(n4663) );
  AOI221_X1 U5309 ( .B1(REG0_REG_27__SCAN_IN), .B2(keyinput123), .C1(
        keyinput67), .C2(DATAO_REG_29__SCAN_IN), .A(n4663), .ZN(n4664) );
  NAND4_X1 U5310 ( .A1(n4667), .A2(n4666), .A3(n4665), .A4(n4664), .ZN(n4686)
         );
  OAI22_X1 U5311 ( .A1(IR_REG_14__SCAN_IN), .A2(keyinput51), .B1(keyinput11), 
        .B2(D_REG_19__SCAN_IN), .ZN(n4668) );
  AOI221_X1 U5312 ( .B1(IR_REG_14__SCAN_IN), .B2(keyinput51), .C1(
        D_REG_19__SCAN_IN), .C2(keyinput11), .A(n4668), .ZN(n4675) );
  OAI22_X1 U5313 ( .A1(D_REG_28__SCAN_IN), .A2(keyinput78), .B1(DATAI_2_), 
        .B2(keyinput7), .ZN(n4669) );
  AOI221_X1 U5314 ( .B1(D_REG_28__SCAN_IN), .B2(keyinput78), .C1(keyinput7), 
        .C2(DATAI_2_), .A(n4669), .ZN(n4674) );
  OAI22_X1 U5315 ( .A1(D_REG_31__SCAN_IN), .A2(keyinput87), .B1(
        IR_REG_27__SCAN_IN), .B2(keyinput99), .ZN(n4670) );
  AOI221_X1 U5316 ( .B1(D_REG_31__SCAN_IN), .B2(keyinput87), .C1(keyinput99), 
        .C2(IR_REG_27__SCAN_IN), .A(n4670), .ZN(n4673) );
  OAI22_X1 U5317 ( .A1(IR_REG_17__SCAN_IN), .A2(keyinput59), .B1(
        ADDR_REG_3__SCAN_IN), .B2(keyinput75), .ZN(n4671) );
  AOI221_X1 U5318 ( .B1(IR_REG_17__SCAN_IN), .B2(keyinput59), .C1(keyinput75), 
        .C2(ADDR_REG_3__SCAN_IN), .A(n4671), .ZN(n4672) );
  NAND4_X1 U5319 ( .A1(n4675), .A2(n4674), .A3(n4673), .A4(n4672), .ZN(n4685)
         );
  OAI22_X1 U5320 ( .A1(IR_REG_6__SCAN_IN), .A2(keyinput110), .B1(keyinput98), 
        .B2(DATAO_REG_31__SCAN_IN), .ZN(n4676) );
  AOI221_X1 U5321 ( .B1(IR_REG_6__SCAN_IN), .B2(keyinput110), .C1(
        DATAO_REG_31__SCAN_IN), .C2(keyinput98), .A(n4676), .ZN(n4683) );
  OAI22_X1 U5322 ( .A1(D_REG_4__SCAN_IN), .A2(keyinput32), .B1(
        REG3_REG_6__SCAN_IN), .B2(keyinput48), .ZN(n4677) );
  AOI221_X1 U5323 ( .B1(D_REG_4__SCAN_IN), .B2(keyinput32), .C1(keyinput48), 
        .C2(REG3_REG_6__SCAN_IN), .A(n4677), .ZN(n4682) );
  OAI22_X1 U5324 ( .A1(REG1_REG_16__SCAN_IN), .A2(keyinput2), .B1(keyinput10), 
        .B2(REG0_REG_12__SCAN_IN), .ZN(n4678) );
  AOI221_X1 U5325 ( .B1(REG1_REG_16__SCAN_IN), .B2(keyinput2), .C1(
        REG0_REG_12__SCAN_IN), .C2(keyinput10), .A(n4678), .ZN(n4681) );
  OAI22_X1 U5326 ( .A1(D_REG_1__SCAN_IN), .A2(keyinput102), .B1(DATAI_1_), 
        .B2(keyinput22), .ZN(n4679) );
  AOI221_X1 U5327 ( .B1(D_REG_1__SCAN_IN), .B2(keyinput102), .C1(keyinput22), 
        .C2(DATAI_1_), .A(n4679), .ZN(n4680) );
  NAND4_X1 U5328 ( .A1(n4683), .A2(n4682), .A3(n4681), .A4(n4680), .ZN(n4684)
         );
  NOR4_X1 U5329 ( .A1(n4687), .A2(n4686), .A3(n4685), .A4(n4684), .ZN(n4688)
         );
  NAND4_X1 U5330 ( .A1(n4691), .A2(n4690), .A3(n4689), .A4(n4688), .ZN(n4692)
         );
  XNOR2_X1 U5331 ( .A(n4693), .B(n4692), .ZN(U3505) );
  MUX2_X1 U5332 ( .A(n4694), .B(REG0_REG_18__SCAN_IN), .S(n5071), .Z(U3503) );
  INV_X1 U5333 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4696) );
  MUX2_X1 U5334 ( .A(n4696), .B(n4695), .S(n5073), .Z(n4697) );
  OAI21_X1 U5335 ( .B1(n4698), .B2(n4706), .A(n4697), .ZN(U3501) );
  INV_X1 U5336 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4700) );
  MUX2_X1 U5337 ( .A(n4700), .B(n4699), .S(n5073), .Z(n4701) );
  OAI21_X1 U5338 ( .B1(n4702), .B2(n4706), .A(n4701), .ZN(U3499) );
  INV_X1 U5339 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4704) );
  MUX2_X1 U5340 ( .A(n4704), .B(n4703), .S(n5073), .Z(n4705) );
  OAI21_X1 U5341 ( .B1(n4707), .B2(n4706), .A(n4705), .ZN(U3497) );
  MUX2_X1 U5342 ( .A(REG0_REG_14__SCAN_IN), .B(n4708), .S(n5073), .Z(U3495) );
  MUX2_X1 U5343 ( .A(DATAI_28_), .B(n4789), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U5344 ( .A(n4787), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U5345 ( .A(n2934), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  INV_X1 U5346 ( .A(n4709), .ZN(n4710) );
  MUX2_X1 U5347 ( .A(n4710), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U5348 ( .A(DATAI_20_), .B(n4711), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5349 ( .A(n4712), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5350 ( .A(DATAI_9_), .B(n4856), .S(STATE_REG_SCAN_IN), .Z(U3343) );
  INV_X1 U5351 ( .A(DATAI_1_), .ZN(n4713) );
  AOI22_X1 U5352 ( .A1(STATE_REG_SCAN_IN), .A2(n4714), .B1(n4713), .B2(U3149), 
        .ZN(U3351) );
  AOI22_X1 U5353 ( .A1(STATE_REG_SCAN_IN), .A2(n4716), .B1(n4715), .B2(U3149), 
        .ZN(U3350) );
  INV_X1 U5354 ( .A(DATAI_3_), .ZN(n4717) );
  AOI22_X1 U5355 ( .A1(STATE_REG_SCAN_IN), .A2(n4729), .B1(n4717), .B2(U3149), 
        .ZN(U3349) );
  OAI22_X1 U5356 ( .A1(U3149), .A2(n4718), .B1(DATAI_4_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4719) );
  INV_X1 U5357 ( .A(n4719), .ZN(U3348) );
  AOI211_X1 U5358 ( .C1(n4722), .C2(n4721), .A(n4720), .B(n4824), .ZN(n4723)
         );
  AOI211_X1 U5359 ( .C1(n4953), .C2(ADDR_REG_3__SCAN_IN), .A(n4724), .B(n4723), 
        .ZN(n4728) );
  OAI211_X1 U5360 ( .C1(REG2_REG_3__SCAN_IN), .C2(n4726), .A(n4911), .B(n4725), 
        .ZN(n4727) );
  OAI211_X1 U5361 ( .C1(n4960), .C2(n4729), .A(n4728), .B(n4727), .ZN(U3243)
         );
  NOR2_X1 U5362 ( .A1(STATE_REG_SCAN_IN), .A2(n4730), .ZN(n4934) );
  OAI22_X1 U5363 ( .A1(n4732), .A2(n4744), .B1(n4743), .B2(n4731), .ZN(n4733)
         );
  AOI211_X1 U5364 ( .C1(n2218), .C2(n4734), .A(n4934), .B(n4733), .ZN(n4740)
         );
  INV_X1 U5365 ( .A(n4735), .ZN(n4753) );
  NOR2_X1 U5366 ( .A1(n4748), .A2(n4753), .ZN(n4737) );
  XNOR2_X1 U5367 ( .A(n4737), .B(n4736), .ZN(n4738) );
  NAND2_X1 U5368 ( .A1(n4738), .A2(n4752), .ZN(n4739) );
  OAI211_X1 U5369 ( .C1(n4758), .C2(n4741), .A(n4740), .B(n4739), .ZN(U3223)
         );
  AND2_X1 U5370 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4925) );
  OAI22_X1 U5371 ( .A1(n4745), .A2(n4744), .B1(n4743), .B2(n4742), .ZN(n4746)
         );
  AOI211_X1 U5372 ( .C1(n2218), .C2(n4747), .A(n4925), .B(n4746), .ZN(n4756)
         );
  INV_X1 U5373 ( .A(n4748), .ZN(n4754) );
  OAI21_X1 U5374 ( .B1(n4750), .B2(n4753), .A(n4749), .ZN(n4751) );
  OAI211_X1 U5375 ( .C1(n4754), .C2(n4753), .A(n4752), .B(n4751), .ZN(n4755)
         );
  OAI211_X1 U5376 ( .C1(n4758), .C2(n4757), .A(n4756), .B(n4755), .ZN(U3238)
         );
  AOI22_X1 U5377 ( .A1(n4759), .A2(n4991), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4762), .ZN(n4760) );
  OAI21_X1 U5378 ( .B1(n4762), .B2(n4761), .A(n4760), .ZN(U3261) );
  NAND2_X1 U5379 ( .A1(n4787), .A2(n4763), .ZN(n4764) );
  NAND2_X1 U5380 ( .A1(n4789), .A2(n4764), .ZN(n4792) );
  INV_X1 U5381 ( .A(n4792), .ZN(n4765) );
  OAI21_X1 U5382 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4787), .A(n4765), .ZN(n4766)
         );
  XNOR2_X1 U5383 ( .A(n4766), .B(n5038), .ZN(n4769) );
  AOI22_X1 U5384 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4953), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4767) );
  OAI21_X1 U5385 ( .B1(n4769), .B2(n4768), .A(n4767), .ZN(U3240) );
  AOI22_X1 U5386 ( .A1(ADDR_REG_1__SCAN_IN), .A2(n4953), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4779) );
  NAND2_X1 U5387 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4771) );
  AOI211_X1 U5388 ( .C1(n4772), .C2(n4771), .A(n4770), .B(n4824), .ZN(n4773)
         );
  AOI21_X1 U5389 ( .B1(n4785), .B2(n4774), .A(n4773), .ZN(n4778) );
  OAI211_X1 U5390 ( .C1(n4776), .C2(n4786), .A(n4911), .B(n4775), .ZN(n4777)
         );
  NAND3_X1 U5391 ( .A1(n4779), .A2(n4778), .A3(n4777), .ZN(U3241) );
  AOI22_X1 U5392 ( .A1(n4953), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4802) );
  AOI211_X1 U5393 ( .C1(n4782), .C2(n4781), .A(n4780), .B(n4824), .ZN(n4783)
         );
  AOI21_X1 U5394 ( .B1(n4785), .B2(n4784), .A(n4783), .ZN(n4801) );
  INV_X1 U5395 ( .A(n4786), .ZN(n4795) );
  INV_X1 U5396 ( .A(n4787), .ZN(n4788) );
  NAND3_X1 U5397 ( .A1(n4790), .A2(n4789), .A3(n4788), .ZN(n4794) );
  AOI21_X1 U5398 ( .B1(n4792), .B2(n5038), .A(n4791), .ZN(n4793) );
  OAI211_X1 U5399 ( .C1(n4796), .C2(n4795), .A(n4794), .B(n4793), .ZN(n4806)
         );
  OAI211_X1 U5400 ( .C1(n4799), .C2(n4798), .A(n4911), .B(n4797), .ZN(n4800)
         );
  NAND4_X1 U5401 ( .A1(n4802), .A2(n4801), .A3(n4806), .A4(n4800), .ZN(U3242)
         );
  OAI21_X1 U5402 ( .B1(REG1_REG_4__SCAN_IN), .B2(n4803), .A(n4955), .ZN(n4808)
         );
  OAI211_X1 U5403 ( .C1(REG2_REG_4__SCAN_IN), .C2(n4805), .A(n4911), .B(n4804), 
        .ZN(n4807) );
  OAI211_X1 U5404 ( .C1(n4809), .C2(n4808), .A(n4807), .B(n4806), .ZN(n4810)
         );
  AOI211_X1 U5405 ( .C1(n4953), .C2(ADDR_REG_4__SCAN_IN), .A(n4811), .B(n4810), 
        .ZN(n4812) );
  OAI21_X1 U5406 ( .B1(n2390), .B2(n4960), .A(n4812), .ZN(U3244) );
  AOI211_X1 U5407 ( .C1(n4815), .C2(n4814), .A(n4813), .B(n4824), .ZN(n4817)
         );
  AOI211_X1 U5408 ( .C1(n4953), .C2(ADDR_REG_5__SCAN_IN), .A(n4817), .B(n4816), 
        .ZN(n4822) );
  OAI211_X1 U5409 ( .C1(n4820), .C2(n4819), .A(n4911), .B(n4818), .ZN(n4821)
         );
  OAI211_X1 U5410 ( .C1(n4960), .C2(n4823), .A(n4822), .B(n4821), .ZN(U3245)
         );
  AOI211_X1 U5411 ( .C1(n4827), .C2(n4826), .A(n4825), .B(n4824), .ZN(n4829)
         );
  AOI211_X1 U5412 ( .C1(n4953), .C2(ADDR_REG_6__SCAN_IN), .A(n4829), .B(n4828), 
        .ZN(n4833) );
  OAI211_X1 U5413 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4831), .A(n4911), .B(n4830), 
        .ZN(n4832) );
  OAI211_X1 U5414 ( .C1(n4960), .C2(n3940), .A(n4833), .B(n4832), .ZN(U3246)
         );
  OAI21_X1 U5415 ( .B1(REG1_REG_7__SCAN_IN), .B2(n4835), .A(n4834), .ZN(n4837)
         );
  OAI21_X1 U5416 ( .B1(n4838), .B2(n4837), .A(n4955), .ZN(n4836) );
  AOI21_X1 U5417 ( .B1(n4838), .B2(n4837), .A(n4836), .ZN(n4839) );
  AOI211_X1 U5418 ( .C1(n4953), .C2(ADDR_REG_7__SCAN_IN), .A(n4840), .B(n4839), 
        .ZN(n4845) );
  OAI211_X1 U5419 ( .C1(n4843), .C2(n4842), .A(n4911), .B(n4841), .ZN(n4844)
         );
  OAI211_X1 U5420 ( .C1(n4960), .C2(n5032), .A(n4845), .B(n4844), .ZN(U3247)
         );
  OAI211_X1 U5421 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4847), .A(n4955), .B(n4846), 
        .ZN(n4851) );
  OAI211_X1 U5422 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4849), .A(n4911), .B(n4848), 
        .ZN(n4850) );
  OAI211_X1 U5423 ( .C1(n4960), .C2(n4852), .A(n4851), .B(n4850), .ZN(n4853)
         );
  AOI211_X1 U5424 ( .C1(n4953), .C2(ADDR_REG_8__SCAN_IN), .A(n4854), .B(n4853), 
        .ZN(n4855) );
  INV_X1 U5425 ( .A(n4855), .ZN(U3248) );
  INV_X1 U5426 ( .A(n4856), .ZN(n4865) );
  OAI211_X1 U5427 ( .C1(n4859), .C2(n4858), .A(n4955), .B(n4857), .ZN(n4864)
         );
  OAI211_X1 U5428 ( .C1(n4862), .C2(n4861), .A(n4911), .B(n4860), .ZN(n4863)
         );
  OAI211_X1 U5429 ( .C1(n4960), .C2(n4865), .A(n4864), .B(n4863), .ZN(n4866)
         );
  AOI211_X1 U5430 ( .C1(n4953), .C2(ADDR_REG_9__SCAN_IN), .A(n4867), .B(n4866), 
        .ZN(n4868) );
  INV_X1 U5431 ( .A(n4868), .ZN(U3249) );
  OAI211_X1 U5432 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4870), .A(n4955), .B(n4869), .ZN(n4874) );
  OAI211_X1 U5433 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4872), .A(n4911), .B(n4871), .ZN(n4873) );
  OAI211_X1 U5434 ( .C1(n4960), .C2(n5028), .A(n4874), .B(n4873), .ZN(n4875)
         );
  AOI211_X1 U5435 ( .C1(n4953), .C2(ADDR_REG_10__SCAN_IN), .A(n4876), .B(n4875), .ZN(n4877) );
  INV_X1 U5436 ( .A(n4877), .ZN(U3250) );
  OAI211_X1 U5437 ( .C1(n4880), .C2(n4879), .A(n4955), .B(n4878), .ZN(n4885)
         );
  OAI211_X1 U5438 ( .C1(n4883), .C2(n4882), .A(n4911), .B(n4881), .ZN(n4884)
         );
  OAI211_X1 U5439 ( .C1(n4960), .C2(n5026), .A(n4885), .B(n4884), .ZN(n4886)
         );
  AOI211_X1 U5440 ( .C1(n4953), .C2(ADDR_REG_11__SCAN_IN), .A(n4887), .B(n4886), .ZN(n4888) );
  INV_X1 U5441 ( .A(n4888), .ZN(U3251) );
  OAI211_X1 U5442 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4890), .A(n4955), .B(n4889), .ZN(n4894) );
  OAI211_X1 U5443 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4892), .A(n4911), .B(n4891), .ZN(n4893) );
  OAI211_X1 U5444 ( .C1(n4960), .C2(n4895), .A(n4894), .B(n4893), .ZN(n4896)
         );
  AOI211_X1 U5445 ( .C1(n4953), .C2(ADDR_REG_12__SCAN_IN), .A(n4897), .B(n4896), .ZN(n4898) );
  INV_X1 U5446 ( .A(n4898), .ZN(U3252) );
  AOI22_X1 U5447 ( .A1(REG2_REG_13__SCAN_IN), .A2(n4900), .B1(n5022), .B2(
        n4899), .ZN(n4903) );
  OAI21_X1 U5448 ( .B1(n4903), .B2(n4902), .A(n4911), .ZN(n4901) );
  AOI21_X1 U5449 ( .B1(n4903), .B2(n4902), .A(n4901), .ZN(n4904) );
  AOI211_X1 U5450 ( .C1(ADDR_REG_13__SCAN_IN), .C2(n4953), .A(n4905), .B(n4904), .ZN(n4910) );
  OAI211_X1 U5451 ( .C1(n4908), .C2(n4907), .A(n4955), .B(n4906), .ZN(n4909)
         );
  OAI211_X1 U5452 ( .C1(n4960), .C2(n5022), .A(n4910), .B(n4909), .ZN(U3253)
         );
  INV_X1 U5453 ( .A(n4911), .ZN(n4949) );
  AOI211_X1 U5454 ( .C1(n3533), .C2(n4913), .A(n4912), .B(n4949), .ZN(n4914)
         );
  AOI211_X1 U5455 ( .C1(n4953), .C2(ADDR_REG_14__SCAN_IN), .A(n4915), .B(n4914), .ZN(n4919) );
  OAI211_X1 U5456 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4917), .A(n4955), .B(n4916), .ZN(n4918) );
  OAI211_X1 U5457 ( .C1(n4960), .C2(n4920), .A(n4919), .B(n4918), .ZN(U3254)
         );
  AOI211_X1 U5458 ( .C1(n4923), .C2(n4922), .A(n4921), .B(n4949), .ZN(n4924)
         );
  AOI211_X1 U5459 ( .C1(n4953), .C2(ADDR_REG_15__SCAN_IN), .A(n4925), .B(n4924), .ZN(n4930) );
  OAI211_X1 U5460 ( .C1(n4928), .C2(n4927), .A(n4955), .B(n4926), .ZN(n4929)
         );
  OAI211_X1 U5461 ( .C1(n4960), .C2(n5018), .A(n4930), .B(n4929), .ZN(U3255)
         );
  AOI221_X1 U5462 ( .B1(n4932), .B2(n4931), .C1(n3595), .C2(n4931), .A(n4949), 
        .ZN(n4933) );
  AOI211_X1 U5463 ( .C1(ADDR_REG_16__SCAN_IN), .C2(n4953), .A(n4934), .B(n4933), .ZN(n4938) );
  OAI221_X1 U5464 ( .B1(n4936), .B2(REG1_REG_16__SCAN_IN), .C1(n4936), .C2(
        n4935), .A(n4955), .ZN(n4937) );
  OAI211_X1 U5465 ( .C1(n4960), .C2(n4939), .A(n4938), .B(n4937), .ZN(U3256)
         );
  AOI221_X1 U5466 ( .B1(n4942), .B2(n4941), .C1(n4940), .C2(n4941), .A(n4949), 
        .ZN(n4943) );
  AOI211_X1 U5467 ( .C1(ADDR_REG_17__SCAN_IN), .C2(n4953), .A(n4944), .B(n4943), .ZN(n4948) );
  OAI221_X1 U5468 ( .B1(n4946), .B2(n2238), .C1(n4946), .C2(n4945), .A(n4955), 
        .ZN(n4947) );
  OAI211_X1 U5469 ( .C1(n4960), .C2(n5014), .A(n4948), .B(n4947), .ZN(U3257)
         );
  OAI211_X1 U5470 ( .C1(n4957), .C2(n4956), .A(n4955), .B(n4954), .ZN(n4958)
         );
  OAI211_X1 U5471 ( .C1(n4960), .C2(n5013), .A(n4959), .B(n4958), .ZN(U3258)
         );
  AOI22_X1 U5472 ( .A1(n4961), .A2(n4987), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4762), .ZN(n4966) );
  INV_X1 U5473 ( .A(n4962), .ZN(n4963) );
  AOI22_X1 U5474 ( .A1(n4964), .A2(n4992), .B1(n4991), .B2(n4963), .ZN(n4965)
         );
  OAI211_X1 U5475 ( .C1(n4762), .C2(n4967), .A(n4966), .B(n4965), .ZN(U3280)
         );
  AOI22_X1 U5476 ( .A1(n4968), .A2(n4987), .B1(REG2_REG_8__SCAN_IN), .B2(n4762), .ZN(n4972) );
  AOI22_X1 U5477 ( .A1(n4970), .A2(n4992), .B1(n4991), .B2(n4969), .ZN(n4971)
         );
  OAI211_X1 U5478 ( .C1(n4762), .C2(n4973), .A(n4972), .B(n4971), .ZN(U3282)
         );
  AOI22_X1 U5479 ( .A1(n4974), .A2(n4987), .B1(REG2_REG_6__SCAN_IN), .B2(n4762), .ZN(n4979) );
  INV_X1 U5480 ( .A(n4975), .ZN(n4976) );
  AOI22_X1 U5481 ( .A1(n4977), .A2(n4992), .B1(n4991), .B2(n4976), .ZN(n4978)
         );
  OAI211_X1 U5482 ( .C1(n4762), .C2(n4980), .A(n4979), .B(n4978), .ZN(U3284)
         );
  AOI22_X1 U5483 ( .A1(n4762), .A2(REG2_REG_3__SCAN_IN), .B1(n4987), .B2(n4981), .ZN(n4985) );
  AOI22_X1 U5484 ( .A1(n4983), .A2(n4992), .B1(n4991), .B2(n4982), .ZN(n4984)
         );
  OAI211_X1 U5485 ( .C1(n4762), .C2(n4986), .A(n4985), .B(n4984), .ZN(U3287)
         );
  AOI22_X1 U5486 ( .A1(REG3_REG_2__SCAN_IN), .A2(n4987), .B1(
        REG2_REG_2__SCAN_IN), .B2(n4762), .ZN(n4995) );
  INV_X1 U5487 ( .A(n4988), .ZN(n4993) );
  INV_X1 U5488 ( .A(n4989), .ZN(n4990) );
  AOI22_X1 U5489 ( .A1(n4993), .A2(n4992), .B1(n4991), .B2(n4990), .ZN(n4994)
         );
  OAI211_X1 U5490 ( .C1(n4762), .C2(n4996), .A(n4995), .B(n4994), .ZN(U3288)
         );
  NOR2_X1 U5491 ( .A1(n5009), .A2(n4997), .ZN(U3291) );
  AND2_X1 U5492 ( .A1(D_REG_30__SCAN_IN), .A2(n5007), .ZN(U3292) );
  NOR2_X1 U5493 ( .A1(n5009), .A2(n4998), .ZN(U3293) );
  NOR2_X1 U5494 ( .A1(n5009), .A2(n4999), .ZN(U3294) );
  NOR2_X1 U5495 ( .A1(n5009), .A2(n5000), .ZN(U3295) );
  AND2_X1 U5496 ( .A1(D_REG_26__SCAN_IN), .A2(n5007), .ZN(U3296) );
  AND2_X1 U5497 ( .A1(D_REG_25__SCAN_IN), .A2(n5007), .ZN(U3297) );
  AND2_X1 U5498 ( .A1(D_REG_24__SCAN_IN), .A2(n5007), .ZN(U3298) );
  AND2_X1 U5499 ( .A1(D_REG_23__SCAN_IN), .A2(n5007), .ZN(U3299) );
  NOR2_X1 U5500 ( .A1(n5009), .A2(n5001), .ZN(U3300) );
  AND2_X1 U5501 ( .A1(D_REG_21__SCAN_IN), .A2(n5007), .ZN(U3301) );
  AND2_X1 U5502 ( .A1(D_REG_20__SCAN_IN), .A2(n5007), .ZN(U3302) );
  NOR2_X1 U5503 ( .A1(n5009), .A2(n5002), .ZN(U3303) );
  AND2_X1 U5504 ( .A1(D_REG_18__SCAN_IN), .A2(n5007), .ZN(U3304) );
  AND2_X1 U5505 ( .A1(D_REG_17__SCAN_IN), .A2(n5007), .ZN(U3305) );
  AND2_X1 U5506 ( .A1(D_REG_16__SCAN_IN), .A2(n5007), .ZN(U3306) );
  AND2_X1 U5507 ( .A1(D_REG_15__SCAN_IN), .A2(n5007), .ZN(U3307) );
  AND2_X1 U5508 ( .A1(n5007), .A2(D_REG_14__SCAN_IN), .ZN(U3308) );
  AND2_X1 U5509 ( .A1(n5007), .A2(D_REG_13__SCAN_IN), .ZN(U3309) );
  NOR2_X1 U5510 ( .A1(n5009), .A2(n5003), .ZN(U3310) );
  NOR2_X1 U5511 ( .A1(n5009), .A2(n5004), .ZN(U3311) );
  NOR2_X1 U5512 ( .A1(n5009), .A2(n5005), .ZN(U3312) );
  AND2_X1 U5513 ( .A1(D_REG_9__SCAN_IN), .A2(n5007), .ZN(U3313) );
  AND2_X1 U5514 ( .A1(D_REG_8__SCAN_IN), .A2(n5007), .ZN(U3314) );
  AND2_X1 U5515 ( .A1(n5007), .A2(D_REG_7__SCAN_IN), .ZN(U3315) );
  AND2_X1 U5516 ( .A1(D_REG_6__SCAN_IN), .A2(n5007), .ZN(U3316) );
  AND2_X1 U5517 ( .A1(n5007), .A2(D_REG_5__SCAN_IN), .ZN(U3317) );
  NOR2_X1 U5518 ( .A1(n5009), .A2(n5006), .ZN(U3318) );
  AND2_X1 U5519 ( .A1(D_REG_3__SCAN_IN), .A2(n5007), .ZN(U3319) );
  NOR2_X1 U5520 ( .A1(n5009), .A2(n5008), .ZN(U3320) );
  OAI21_X1 U5521 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n5010), .ZN(
        n5011) );
  INV_X1 U5522 ( .A(n5011), .ZN(U3329) );
  AOI22_X1 U5523 ( .A1(STATE_REG_SCAN_IN), .A2(n5013), .B1(n5012), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5524 ( .A1(STATE_REG_SCAN_IN), .A2(n5014), .B1(n2793), .B2(U3149), 
        .ZN(U3335) );
  OAI22_X1 U5525 ( .A1(U3149), .A2(n5015), .B1(DATAI_16_), .B2(
        STATE_REG_SCAN_IN), .ZN(n5016) );
  INV_X1 U5526 ( .A(n5016), .ZN(U3336) );
  AOI22_X1 U5527 ( .A1(STATE_REG_SCAN_IN), .A2(n5018), .B1(n5017), .B2(U3149), 
        .ZN(U3337) );
  OAI22_X1 U5528 ( .A1(U3149), .A2(n5019), .B1(DATAI_14_), .B2(
        STATE_REG_SCAN_IN), .ZN(n5020) );
  INV_X1 U5529 ( .A(n5020), .ZN(U3338) );
  INV_X1 U5530 ( .A(DATAI_13_), .ZN(n5021) );
  AOI22_X1 U5531 ( .A1(STATE_REG_SCAN_IN), .A2(n5022), .B1(n5021), .B2(U3149), 
        .ZN(U3339) );
  OAI22_X1 U5532 ( .A1(U3149), .A2(n5023), .B1(DATAI_12_), .B2(
        STATE_REG_SCAN_IN), .ZN(n5024) );
  INV_X1 U5533 ( .A(n5024), .ZN(U3340) );
  INV_X1 U5534 ( .A(DATAI_11_), .ZN(n5025) );
  AOI22_X1 U5535 ( .A1(STATE_REG_SCAN_IN), .A2(n5026), .B1(n5025), .B2(U3149), 
        .ZN(U3341) );
  AOI22_X1 U5536 ( .A1(STATE_REG_SCAN_IN), .A2(n5028), .B1(n5027), .B2(U3149), 
        .ZN(U3342) );
  OAI22_X1 U5537 ( .A1(U3149), .A2(n5029), .B1(DATAI_8_), .B2(
        STATE_REG_SCAN_IN), .ZN(n5030) );
  INV_X1 U5538 ( .A(n5030), .ZN(U3344) );
  INV_X1 U5539 ( .A(DATAI_7_), .ZN(n5031) );
  AOI22_X1 U5540 ( .A1(STATE_REG_SCAN_IN), .A2(n5032), .B1(n5031), .B2(U3149), 
        .ZN(U3345) );
  OAI22_X1 U5541 ( .A1(U3149), .A2(n5033), .B1(DATAI_6_), .B2(
        STATE_REG_SCAN_IN), .ZN(n5034) );
  INV_X1 U5542 ( .A(n5034), .ZN(U3346) );
  OAI22_X1 U5543 ( .A1(U3149), .A2(n5035), .B1(DATAI_5_), .B2(
        STATE_REG_SCAN_IN), .ZN(n5036) );
  INV_X1 U5544 ( .A(n5036), .ZN(U3347) );
  AOI22_X1 U5545 ( .A1(STATE_REG_SCAN_IN), .A2(n5038), .B1(n5037), .B2(U3149), 
        .ZN(U3352) );
  INV_X1 U5546 ( .A(n5039), .ZN(n5041) );
  OAI22_X1 U5547 ( .A1(n5042), .A2(n5065), .B1(n5041), .B2(n5040), .ZN(n5043)
         );
  NOR2_X1 U5548 ( .A1(n5044), .A2(n5043), .ZN(n5075) );
  AOI22_X1 U5549 ( .A1(n5073), .A2(n5075), .B1(n5045), .B2(n5071), .ZN(U3467)
         );
  OAI22_X1 U5550 ( .A1(n5048), .A2(n5065), .B1(n5047), .B2(n5046), .ZN(n5049)
         );
  NOR2_X1 U5551 ( .A1(n5050), .A2(n5049), .ZN(n5077) );
  AOI22_X1 U5552 ( .A1(n5073), .A2(n5077), .B1(n5051), .B2(n5071), .ZN(U3469)
         );
  INV_X1 U5553 ( .A(n5052), .ZN(n5054) );
  AOI211_X1 U5554 ( .C1(n5056), .C2(n5055), .A(n5054), .B(n5053), .ZN(n5078)
         );
  INV_X1 U5555 ( .A(REG0_REG_4__SCAN_IN), .ZN(n5057) );
  AOI22_X1 U5556 ( .A1(n5073), .A2(n5078), .B1(n5057), .B2(n5071), .ZN(U3475)
         );
  NOR2_X1 U5557 ( .A1(n5059), .A2(n5058), .ZN(n5063) );
  AOI211_X1 U5558 ( .C1(n5063), .C2(n5062), .A(n5061), .B(n5060), .ZN(n5080)
         );
  INV_X1 U5559 ( .A(REG0_REG_7__SCAN_IN), .ZN(n5064) );
  AOI22_X1 U5560 ( .A1(n5073), .A2(n5080), .B1(n5064), .B2(n5071), .ZN(U3481)
         );
  NOR2_X1 U5561 ( .A1(n5066), .A2(n5065), .ZN(n5068) );
  AOI211_X1 U5562 ( .C1(n5070), .C2(n5069), .A(n5068), .B(n5067), .ZN(n5083)
         );
  INV_X1 U5563 ( .A(REG0_REG_11__SCAN_IN), .ZN(n5072) );
  AOI22_X1 U5564 ( .A1(n5073), .A2(n5083), .B1(n5072), .B2(n5071), .ZN(U3489)
         );
  AOI22_X1 U5565 ( .A1(n5081), .A2(n5075), .B1(n5074), .B2(n3451), .ZN(U3518)
         );
  AOI22_X1 U5566 ( .A1(n5081), .A2(n5077), .B1(n5076), .B2(n3451), .ZN(U3519)
         );
  AOI22_X1 U5567 ( .A1(n5081), .A2(n5078), .B1(n2305), .B2(n3451), .ZN(U3522)
         );
  AOI22_X1 U5568 ( .A1(n5081), .A2(n5080), .B1(n5079), .B2(n3451), .ZN(U3525)
         );
  AOI22_X1 U5569 ( .A1(n5081), .A2(n5083), .B1(n5082), .B2(n3451), .ZN(U3529)
         );
  CLKBUF_X1 U2468 ( .A(n2525), .Z(n3819) );
  OAI21_X1 U2513 ( .B1(n4218), .B2(n4217), .A(n4216), .ZN(n4698) );
endmodule

