

module b14_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, 
        DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, 
        DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, 
        DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, 
        DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, 
        DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257;

  NAND2_X1 U2517 ( .A1(n2876), .A2(n2929), .ZN(n2880) );
  NAND2_X1 U2518 ( .A1(n2874), .A2(n4625), .ZN(n2929) );
  OR2_X1 U2519 ( .A1(n2902), .A2(n2765), .ZN(n2845) );
  NOR2_X1 U2520 ( .A1(n2903), .A2(IR_REG_19__SCAN_IN), .ZN(n2902) );
  OAI21_X1 U2521 ( .B1(n2752), .B2(IR_REG_16__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2844) );
  CLKBUF_X2 U2522 ( .A(n2483), .Z(n4188) );
  NOR2_X1 U2524 ( .A1(n2675), .A2(IR_REG_9__SCAN_IN), .ZN(n2674) );
  INV_X1 U2525 ( .A(n4016), .ZN(n3968) );
  INV_X1 U2526 ( .A(n2937), .ZN(n4010) );
  NAND2_X2 U2527 ( .A1(n2609), .A2(n2555), .ZN(n4258) );
  OR2_X1 U2528 ( .A1(n3534), .A2(n3536), .ZN(n3558) );
  INV_X1 U2529 ( .A(n2950), .ZN(n4833) );
  NAND2_X1 U2530 ( .A1(n2552), .A2(IR_REG_31__SCAN_IN), .ZN(n2779) );
  NAND2_X1 U2531 ( .A1(n2770), .A2(n4623), .ZN(n2876) );
  CLKBUF_X3 U2532 ( .A(n2983), .Z(n2483) );
  NAND2_X2 U2533 ( .A1(n4423), .A2(n4433), .ZN(n4401) );
  NAND2_X2 U2534 ( .A1(n2790), .A2(n2791), .ZN(n2482) );
  NAND2_X2 U2535 ( .A1(n2790), .A2(n2791), .ZN(n2977) );
  NOR2_X1 U2536 ( .A1(n4620), .A2(n4621), .ZN(n2939) );
  NAND2_X1 U2537 ( .A1(n4620), .A2(n4621), .ZN(n3785) );
  AND2_X1 U2538 ( .A1(n2869), .A2(n4620), .ZN(n2981) );
  AND2_X1 U2539 ( .A1(n4371), .A2(n2537), .ZN(n2536) );
  AND2_X1 U2540 ( .A1(n4383), .A2(n4382), .ZN(n4385) );
  AOI21_X1 U2541 ( .B1(n4401), .B2(n3851), .A(n4209), .ZN(n4383) );
  AND2_X1 U2542 ( .A1(n3991), .A2(n3990), .ZN(n4078) );
  NAND2_X1 U2543 ( .A1(n2650), .A2(n4113), .ZN(n4067) );
  OAI21_X1 U2544 ( .B1(n5056), .B2(n5055), .A(n3927), .ZN(n5074) );
  AOI22_X1 U2545 ( .A1(n5037), .A2(n5038), .B1(n3920), .B2(n3919), .ZN(n5056)
         );
  OR2_X2 U2546 ( .A1(n4488), .A2(n4475), .ZN(n4473) );
  OAI21_X1 U2547 ( .B1(n3897), .B2(n2662), .A(n2659), .ZN(n2664) );
  OAI21_X1 U2548 ( .B1(n3556), .B2(n2584), .A(n2582), .ZN(n3643) );
  NAND2_X1 U2549 ( .A1(n3487), .A2(n4058), .ZN(n4104) );
  AND2_X1 U2550 ( .A1(n5142), .A2(n2545), .ZN(n5140) );
  OR2_X2 U2551 ( .A1(n3656), .A2(n5022), .ZN(n3676) );
  AOI21_X1 U2552 ( .B1(n3467), .B2(n3466), .A(n2678), .ZN(n4133) );
  INV_X2 U2553 ( .A(n4652), .ZN(n4656) );
  NAND2_X4 U2554 ( .A1(n5219), .A2(n3469), .ZN(n2937) );
  NAND4_X1 U2555 ( .A1(n2993), .A2(n2992), .A3(n2991), .A4(n2990), .ZN(n4331)
         );
  NAND4_X2 U2556 ( .A1(n2987), .A2(n2986), .A3(n2985), .A4(n2984), .ZN(n4332)
         );
  NAND2_X2 U2557 ( .A1(n2929), .A2(n2930), .ZN(n4016) );
  NAND4_X2 U2558 ( .A1(n2873), .A2(n2872), .A3(n2871), .A4(n2870), .ZN(n2951)
         );
  NAND2_X2 U2559 ( .A1(n2874), .A2(n2906), .ZN(n5219) );
  CLKBUF_X1 U2560 ( .A(n2981), .Z(n2484) );
  CLKBUF_X1 U2561 ( .A(n2790), .Z(n4805) );
  CLKBUF_X1 U2562 ( .A(n2791), .Z(n4657) );
  NAND2_X1 U2563 ( .A1(n2865), .A2(IR_REG_31__SCAN_IN), .ZN(n2864) );
  NAND2_X1 U2564 ( .A1(n2776), .A2(IR_REG_31__SCAN_IN), .ZN(n2777) );
  INV_X1 U2565 ( .A(n2767), .ZN(n2782) );
  AND2_X1 U2566 ( .A1(n2716), .A2(n2553), .ZN(n2551) );
  AND2_X1 U2567 ( .A1(n2674), .A2(n2673), .ZN(n2672) );
  NOR2_X1 U2568 ( .A1(n2764), .A2(IR_REG_25__SCAN_IN), .ZN(n2676) );
  AND2_X1 U2569 ( .A1(n2684), .A2(n2741), .ZN(n2553) );
  NOR2_X1 U2570 ( .A1(n2759), .A2(n2842), .ZN(n2760) );
  AND2_X1 U2571 ( .A1(n2781), .A2(n2762), .ZN(n2768) );
  NAND4_X1 U2572 ( .A1(n2758), .A2(n3179), .A3(n3374), .A4(n3377), .ZN(n2759)
         );
  AND2_X1 U2573 ( .A1(n3382), .A2(n3188), .ZN(n2763) );
  AND3_X1 U2574 ( .A1(n3348), .A2(n3352), .A3(n3351), .ZN(n2684) );
  INV_X1 U2575 ( .A(IR_REG_12__SCAN_IN), .ZN(n3170) );
  INV_X1 U2576 ( .A(IR_REG_11__SCAN_IN), .ZN(n3166) );
  INV_X1 U2577 ( .A(IR_REG_16__SCAN_IN), .ZN(n3179) );
  INV_X1 U2578 ( .A(IR_REG_17__SCAN_IN), .ZN(n3376) );
  INV_X1 U2579 ( .A(IR_REG_6__SCAN_IN), .ZN(n3352) );
  INV_X1 U2580 ( .A(IR_REG_19__SCAN_IN), .ZN(n3377) );
  INV_X1 U2581 ( .A(IR_REG_21__SCAN_IN), .ZN(n2781) );
  INV_X1 U2582 ( .A(IR_REG_23__SCAN_IN), .ZN(n3382) );
  INV_X1 U2583 ( .A(IR_REG_24__SCAN_IN), .ZN(n3188) );
  INV_X1 U2584 ( .A(IR_REG_7__SCAN_IN), .ZN(n3348) );
  INV_X2 U2585 ( .A(IR_REG_20__SCAN_IN), .ZN(n3374) );
  NAND2_X2 U2586 ( .A1(n2943), .A2(n2682), .ZN(n2978) );
  NOR2_X2 U2587 ( .A1(n2951), .A2(n4833), .ZN(n4260) );
  NOR2_X1 U2588 ( .A1(n2869), .A2(n4620), .ZN(n2983) );
  XNOR2_X2 U2589 ( .A(n2777), .B(n3391), .ZN(n2790) );
  BUF_X4 U2590 ( .A(n2981), .Z(n2485) );
  NAND2_X1 U2591 ( .A1(n2876), .A2(n2929), .ZN(n2486) );
  INV_X2 U2592 ( .A(n3785), .ZN(n2487) );
  NOR2_X1 U2593 ( .A1(n4122), .A2(n2649), .ZN(n2648) );
  INV_X1 U2594 ( .A(n4113), .ZN(n2649) );
  AND2_X1 U2595 ( .A1(n3541), .A2(n4149), .ZN(n3542) );
  NAND2_X1 U2596 ( .A1(n2551), .A2(n2672), .ZN(n2757) );
  INV_X1 U2597 ( .A(n2648), .ZN(n2647) );
  NOR2_X1 U2598 ( .A1(n2514), .A2(n2490), .ZN(n2645) );
  NAND2_X1 U2599 ( .A1(n3898), .A2(n3900), .ZN(n3901) );
  NOR2_X1 U2600 ( .A1(n4410), .A2(n4452), .ZN(n2566) );
  AOI21_X1 U2601 ( .B1(n3727), .B2(n2572), .A(n2570), .ZN(n2569) );
  OAI21_X1 U2602 ( .B1(n2571), .B2(n2579), .A(n2489), .ZN(n2570) );
  NOR2_X1 U2603 ( .A1(n3068), .A2(n2564), .ZN(n2563) );
  INV_X1 U2604 ( .A(n3543), .ZN(n2564) );
  OAI211_X1 U2605 ( .C1(n2966), .C2(n2965), .A(STATE_REG_SCAN_IN), .B(n2964), 
        .ZN(n4568) );
  OAI21_X1 U2606 ( .B1(n5108), .B2(n2656), .A(n2653), .ZN(n5182) );
  NAND2_X1 U2607 ( .A1(n2488), .A2(n2657), .ZN(n2656) );
  AOI21_X1 U2608 ( .B1(n2488), .B2(n2513), .A(n2654), .ZN(n2653) );
  INV_X1 U2609 ( .A(n5107), .ZN(n2657) );
  OAI22_X1 U2610 ( .A1(n4835), .A2(n2937), .B1(n4258), .B2(n4015), .ZN(n3465)
         );
  NAND2_X1 U2611 ( .A1(n2949), .A2(n3468), .ZN(n2935) );
  INV_X1 U2612 ( .A(n2509), .ZN(n2662) );
  NAND2_X1 U2613 ( .A1(n5182), .A2(n5183), .ZN(n5181) );
  AND2_X1 U2614 ( .A1(n3044), .A2(n3043), .ZN(n3541) );
  NOR2_X1 U2615 ( .A1(n2833), .A2(n2832), .ZN(n3871) );
  NAND2_X1 U2616 ( .A1(n4360), .A2(n4184), .ZN(n4353) );
  AND2_X1 U2617 ( .A1(n2577), .A2(n2581), .ZN(n2576) );
  NAND2_X1 U2618 ( .A1(n2579), .A2(n2580), .ZN(n2577) );
  NAND2_X1 U2619 ( .A1(n2501), .A2(n2590), .ZN(n2587) );
  INV_X1 U2620 ( .A(n3540), .ZN(n4149) );
  OR2_X1 U2621 ( .A1(n5219), .A2(n4840), .ZN(n4566) );
  NOR2_X1 U2622 ( .A1(n2860), .A2(IR_REG_28__SCAN_IN), .ZN(n2861) );
  INV_X1 U2623 ( .A(n4741), .ZN(n2627) );
  INV_X1 U2624 ( .A(n4762), .ZN(n2614) );
  INV_X1 U2625 ( .A(n4782), .ZN(n2618) );
  NAND2_X1 U2626 ( .A1(n4436), .A2(n4096), .ZN(n2549) );
  XNOR2_X1 U2627 ( .A(n3472), .B(n3968), .ZN(n3474) );
  NAND2_X1 U2628 ( .A1(n2644), .A2(n2515), .ZN(n4077) );
  NAND2_X1 U2629 ( .A1(n2645), .A2(n2647), .ZN(n2643) );
  AND3_X1 U2630 ( .A1(n2876), .A2(n2919), .A3(n2913), .ZN(n2964) );
  AND2_X1 U2631 ( .A1(n2704), .A2(n4685), .ZN(n2706) );
  NOR2_X1 U2632 ( .A1(n4677), .A2(n2805), .ZN(n2806) );
  NOR2_X1 U2633 ( .A1(n4688), .A2(n2809), .ZN(n2810) );
  INV_X1 U2634 ( .A(n2808), .ZN(n2809) );
  INV_X1 U2635 ( .A(n2714), .ZN(n2715) );
  AND3_X1 U2636 ( .A1(n2620), .A2(n2721), .A3(n2619), .ZN(n2725) );
  AND2_X1 U2637 ( .A1(n4410), .A2(n4096), .ZN(n4182) );
  NOR2_X1 U2638 ( .A1(n4410), .A2(n4096), .ZN(n4178) );
  AND2_X1 U2639 ( .A1(n4482), .A2(n4475), .ZN(n4177) );
  AND2_X1 U2640 ( .A1(n2587), .A2(n2586), .ZN(n2585) );
  INV_X1 U2641 ( .A(n4229), .ZN(n2586) );
  NAND2_X1 U2642 ( .A1(n4325), .A2(n3605), .ZN(n2590) );
  NAND2_X1 U2643 ( .A1(n4624), .A2(n4625), .ZN(n2955) );
  INV_X1 U2644 ( .A(n2978), .ZN(n2979) );
  NAND2_X1 U2645 ( .A1(n2768), .A2(n2763), .ZN(n2764) );
  NAND2_X1 U2646 ( .A1(n2785), .A2(IR_REG_31__SCAN_IN), .ZN(n2771) );
  NAND2_X1 U2647 ( .A1(n2771), .A2(n3382), .ZN(n2773) );
  NAND2_X1 U2648 ( .A1(n2782), .A2(n2768), .ZN(n2785) );
  AND2_X1 U2649 ( .A1(n4622), .A2(n3461), .ZN(n2770) );
  AND2_X1 U2650 ( .A1(n2510), .A2(n4004), .ZN(n2671) );
  NOR2_X1 U2651 ( .A1(n4031), .A2(n2669), .ZN(n2668) );
  INV_X1 U2652 ( .A(n2671), .ZN(n2669) );
  INV_X1 U2653 ( .A(n5004), .ZN(n2661) );
  INV_X2 U2654 ( .A(n3468), .ZN(n4015) );
  INV_X1 U2655 ( .A(n4998), .ZN(n2663) );
  NAND2_X1 U2656 ( .A1(n3897), .A2(n3896), .ZN(n4049) );
  NAND2_X1 U2657 ( .A1(n4049), .A2(n3901), .ZN(n5001) );
  XNOR2_X1 U2658 ( .A(n3501), .B(n3502), .ZN(n4141) );
  INV_X1 U2659 ( .A(n4320), .ZN(n5070) );
  OR2_X1 U2660 ( .A1(n2917), .A2(n2901), .ZN(n2921) );
  INV_X1 U2661 ( .A(n4625), .ZN(n4243) );
  AND2_X1 U2662 ( .A1(n3592), .A2(n3591), .ZN(n3889) );
  XNOR2_X1 U2663 ( .A(n2692), .B(REG1_REG_1__SCAN_IN), .ZN(n4666) );
  NAND2_X1 U2664 ( .A1(n2603), .A2(n2602), .ZN(n4792) );
  INV_X1 U2665 ( .A(n4795), .ZN(n2603) );
  NAND2_X1 U2666 ( .A1(n2697), .A2(n2696), .ZN(n2698) );
  XNOR2_X1 U2667 ( .A(n2806), .B(n4892), .ZN(n4817) );
  XNOR2_X1 U2668 ( .A(n2810), .B(n4706), .ZN(n4698) );
  OR2_X1 U2669 ( .A1(n4702), .A2(n2622), .ZN(n2619) );
  OR2_X1 U2670 ( .A1(n4716), .A2(n4701), .ZN(n2622) );
  NAND2_X1 U2671 ( .A1(n2719), .A2(n2621), .ZN(n2620) );
  INV_X1 U2672 ( .A(n4716), .ZN(n2621) );
  OR2_X1 U2673 ( .A1(n4702), .A2(n4701), .ZN(n2624) );
  OR2_X1 U2674 ( .A1(n2854), .A2(n2517), .ZN(n2596) );
  OR2_X1 U2675 ( .A1(n2491), .A2(n4721), .ZN(n2597) );
  OR2_X1 U2676 ( .A1(n2851), .A2(n2636), .ZN(n2635) );
  OR2_X1 U2677 ( .A1(n4725), .A2(n2852), .ZN(n2636) );
  OR2_X1 U2678 ( .A1(n2492), .A2(n4725), .ZN(n2637) );
  OR2_X1 U2679 ( .A1(n2851), .A2(n2852), .ZN(n2638) );
  NOR2_X1 U2680 ( .A1(n4731), .A2(n4732), .ZN(n4730) );
  NAND2_X1 U2681 ( .A1(n4783), .A2(n2825), .ZN(n2826) );
  XNOR2_X1 U2682 ( .A(n2826), .B(n5105), .ZN(n4334) );
  NAND2_X1 U2683 ( .A1(n2631), .A2(n2529), .ZN(n2630) );
  INV_X1 U2684 ( .A(n4347), .ZN(n2633) );
  AOI21_X1 U2685 ( .B1(n2567), .B2(n2565), .A(n3810), .ZN(n4381) );
  NOR2_X1 U2686 ( .A1(n3806), .A2(n2566), .ZN(n2565) );
  NAND2_X1 U2687 ( .A1(n2568), .A2(n2499), .ZN(n2567) );
  OAI22_X1 U2688 ( .A1(n4443), .A2(n4450), .B1(n4452), .B2(n4410), .ZN(n4432)
         );
  OR2_X1 U2689 ( .A1(n3771), .A2(n3770), .ZN(n3782) );
  AND2_X1 U2690 ( .A1(n5200), .A2(n4169), .ZN(n4532) );
  NAND2_X1 U2691 ( .A1(n3726), .A2(n2508), .ZN(n2580) );
  NOR2_X1 U2692 ( .A1(n3723), .A2(n3722), .ZN(n3724) );
  NOR2_X1 U2693 ( .A1(n4319), .A2(n5089), .ZN(n3722) );
  INV_X1 U2694 ( .A(n5057), .ZN(n3924) );
  NAND2_X1 U2695 ( .A1(n3555), .A2(n2590), .ZN(n2588) );
  AND2_X1 U2696 ( .A1(n3565), .A2(n3564), .ZN(n4238) );
  NAND2_X1 U2697 ( .A1(n3047), .A2(n4232), .ZN(n3069) );
  AND2_X1 U2698 ( .A1(n2999), .A2(n2975), .ZN(n2556) );
  NAND2_X1 U2699 ( .A1(n2977), .A2(n3306), .ZN(n2609) );
  OR2_X1 U2700 ( .A1(n2977), .A2(n4673), .ZN(n2555) );
  NAND2_X1 U2701 ( .A1(n3855), .A2(n3854), .ZN(n3865) );
  NOR2_X1 U2702 ( .A1(n2563), .A2(n2560), .ZN(n2559) );
  NAND2_X1 U2703 ( .A1(n4234), .A2(n2561), .ZN(n2560) );
  INV_X1 U2704 ( .A(n3542), .ZN(n2561) );
  AND2_X1 U2705 ( .A1(n2876), .A2(n4628), .ZN(n2910) );
  NAND2_X1 U2706 ( .A1(n2848), .A2(n4622), .ZN(n2966) );
  NAND2_X1 U2707 ( .A1(n2865), .A2(n2868), .ZN(n2869) );
  INV_X1 U2708 ( .A(IR_REG_13__SCAN_IN), .ZN(n2673) );
  NAND2_X1 U2709 ( .A1(n2640), .A2(n2639), .ZN(n2641) );
  INV_X1 U2710 ( .A(IR_REG_0__SCAN_IN), .ZN(n2640) );
  INV_X1 U2711 ( .A(IR_REG_1__SCAN_IN), .ZN(n2639) );
  INV_X1 U2712 ( .A(n3827), .ZN(n4355) );
  AOI22_X1 U2713 ( .A1(n5074), .A2(n3935), .B1(n3934), .B2(n5071), .ZN(n5108)
         );
  AND2_X1 U2714 ( .A1(n5190), .A2(n5177), .ZN(n4148) );
  CLKBUF_X1 U2715 ( .A(U4043), .Z(n4328) );
  INV_X1 U2716 ( .A(n4824), .ZN(n4798) );
  NOR2_X1 U2717 ( .A1(n3871), .A2(n3870), .ZN(n3874) );
  NAND2_X1 U2718 ( .A1(n4558), .A2(n4981), .ZN(n5103) );
  NAND2_X1 U2719 ( .A1(n2905), .A2(n2904), .ZN(n4840) );
  NAND2_X1 U2720 ( .A1(n4564), .A2(n2536), .ZN(n4608) );
  INV_X1 U2721 ( .A(n4563), .ZN(n4564) );
  NOR2_X1 U2722 ( .A1(n2496), .A2(n2538), .ZN(n2537) );
  INV_X1 U2723 ( .A(n4114), .ZN(n2646) );
  INV_X1 U2724 ( .A(IR_REG_18__SCAN_IN), .ZN(n3180) );
  INV_X1 U2725 ( .A(n2576), .ZN(n2573) );
  INV_X1 U2726 ( .A(n5157), .ZN(n2654) );
  OR2_X1 U2727 ( .A1(n5125), .A2(n2507), .ZN(n2658) );
  NOR2_X1 U2728 ( .A1(n3938), .A2(n3937), .ZN(n2655) );
  INV_X1 U2729 ( .A(n2929), .ZN(n2875) );
  NAND2_X1 U2730 ( .A1(n4792), .A2(n2802), .ZN(n2803) );
  AND2_X1 U2731 ( .A1(n2803), .A2(n4685), .ZN(n2805) );
  AND3_X1 U2732 ( .A1(n2637), .A2(n2635), .A3(n2520), .ZN(n2726) );
  NOR2_X1 U2733 ( .A1(n4743), .A2(n2817), .ZN(n2819) );
  AND2_X1 U2734 ( .A1(n4995), .A2(REG1_REG_11__SCAN_IN), .ZN(n2817) );
  NAND2_X1 U2735 ( .A1(n2626), .A2(n2625), .ZN(n2628) );
  AOI21_X1 U2736 ( .B1(n2493), .B2(n2627), .A(n2730), .ZN(n2625) );
  NAND2_X1 U2737 ( .A1(n4730), .A2(n2627), .ZN(n2626) );
  NAND2_X1 U2738 ( .A1(n2613), .A2(n2611), .ZN(n2615) );
  AOI21_X1 U2739 ( .B1(n2735), .B2(n2614), .A(n2612), .ZN(n2611) );
  INV_X1 U2740 ( .A(n2738), .ZN(n2612) );
  NOR2_X1 U2741 ( .A1(n4763), .A2(n2822), .ZN(n2823) );
  INV_X1 U2742 ( .A(n2821), .ZN(n2822) );
  NAND2_X1 U2743 ( .A1(n2617), .A2(n2616), .ZN(n2750) );
  NOR2_X1 U2744 ( .A1(n4575), .A2(n3827), .ZN(n4373) );
  INV_X1 U2745 ( .A(n4374), .ZN(n4372) );
  NAND2_X1 U2746 ( .A1(n4486), .A2(n3779), .ZN(n2568) );
  AND2_X1 U2747 ( .A1(n4425), .A2(n4415), .ZN(n4209) );
  INV_X1 U2748 ( .A(n4522), .ZN(n3840) );
  AND2_X1 U2749 ( .A1(n4221), .A2(n3718), .ZN(n3719) );
  INV_X1 U2750 ( .A(n5079), .ZN(n3723) );
  NOR2_X1 U2751 ( .A1(n4321), .A2(n5039), .ZN(n3720) );
  INV_X1 U2752 ( .A(REG3_REG_12__SCAN_IN), .ZN(n3625) );
  INV_X1 U2753 ( .A(n2955), .ZN(n2922) );
  NAND2_X1 U2754 ( .A1(n3180), .A2(n3376), .ZN(n2842) );
  INV_X1 U2755 ( .A(n2966), .ZN(n2899) );
  INV_X1 U2756 ( .A(n4362), .ZN(n3855) );
  NAND2_X1 U2757 ( .A1(n2548), .A2(n4415), .ZN(n2547) );
  INV_X1 U2758 ( .A(n2549), .ZN(n2548) );
  NOR2_X1 U2759 ( .A1(n4473), .A2(n2549), .ZN(n4434) );
  AND2_X1 U2760 ( .A1(n2954), .A2(n4243), .ZN(n2906) );
  INV_X1 U2761 ( .A(IR_REG_26__SCAN_IN), .ZN(n3192) );
  INV_X1 U2762 ( .A(REG3_REG_14__SCAN_IN), .ZN(n3668) );
  AND2_X1 U2763 ( .A1(n3981), .A2(n4039), .ZN(n4042) );
  NAND2_X1 U2764 ( .A1(n2642), .A2(n2645), .ZN(n4043) );
  AND2_X1 U2765 ( .A1(n4199), .A2(DATAI_28_), .ZN(n3827) );
  INV_X1 U2766 ( .A(n4313), .ZN(n4025) );
  INV_X1 U2767 ( .A(n4424), .ZN(n4436) );
  NAND2_X1 U2768 ( .A1(n4104), .A2(n3491), .ZN(n4908) );
  AND2_X1 U2769 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n3003) );
  AND2_X1 U2770 ( .A1(n2883), .A2(n2882), .ZN(n2932) );
  NOR2_X1 U2771 ( .A1(n3626), .A2(n3625), .ZN(n3648) );
  NAND2_X1 U2772 ( .A1(n3648), .A2(REG3_REG_13__SCAN_IN), .ZN(n3669) );
  INV_X1 U2773 ( .A(n4480), .ZN(n4489) );
  NAND2_X1 U2774 ( .A1(n3608), .A2(REG3_REG_11__SCAN_IN), .ZN(n3626) );
  INV_X1 U2775 ( .A(n4317), .ZN(n4549) );
  OAI21_X1 U2776 ( .B1(n5108), .B2(n5107), .A(n2652), .ZN(n5126) );
  INV_X1 U2777 ( .A(n2655), .ZN(n2652) );
  NOR2_X1 U2778 ( .A1(n3041), .A2(n3040), .ZN(n3059) );
  INV_X1 U2780 ( .A(n2921), .ZN(n2908) );
  AND4_X1 U2781 ( .A1(n3862), .A2(n3861), .A3(n3860), .A4(n3859), .ZN(n4201)
         );
  AND4_X1 U2782 ( .A1(n3805), .A2(n3804), .A3(n3803), .A4(n3802), .ZN(n4386)
         );
  AND4_X1 U2783 ( .A1(n3797), .A2(n3796), .A3(n3795), .A4(n3794), .ZN(n4097)
         );
  AND2_X1 U2784 ( .A1(n3769), .A2(n3768), .ZN(n4071) );
  AND2_X1 U2785 ( .A1(n3731), .A2(n3730), .ZN(n5122) );
  NAND2_X1 U2786 ( .A1(n4667), .A2(n2801), .ZN(n2602) );
  AND2_X1 U2787 ( .A1(n4663), .A2(n2693), .ZN(n4801) );
  NOR2_X1 U2788 ( .A1(n2805), .A2(n2804), .ZN(n4676) );
  NOR2_X1 U2789 ( .A1(n2803), .A2(n4685), .ZN(n2804) );
  NOR2_X1 U2790 ( .A1(n2706), .A2(n2705), .ZN(n4679) );
  AND2_X1 U2791 ( .A1(n4679), .A2(REG2_REG_3__SCAN_IN), .ZN(n4680) );
  OR2_X1 U2792 ( .A1(n4817), .A2(n4898), .ZN(n2594) );
  NOR2_X1 U2793 ( .A1(n4698), .A2(n4929), .ZN(n4697) );
  OR2_X1 U2794 ( .A1(n2854), .A2(n4959), .ZN(n2598) );
  AND3_X1 U2795 ( .A1(n2597), .A2(n2596), .A3(n2519), .ZN(n2814) );
  XNOR2_X1 U2796 ( .A(n2628), .B(n5017), .ZN(n4754) );
  XNOR2_X1 U2797 ( .A(n2819), .B(n2818), .ZN(n4751) );
  NOR2_X1 U2798 ( .A1(n4751), .A2(n5031), .ZN(n4750) );
  NOR2_X1 U2799 ( .A1(n4754), .A2(n3659), .ZN(n4753) );
  XNOR2_X1 U2800 ( .A(n2615), .B(n3682), .ZN(n4774) );
  NOR2_X1 U2801 ( .A1(n4774), .A2(n4773), .ZN(n4772) );
  OR2_X1 U2802 ( .A1(n4786), .A2(n4785), .ZN(n4783) );
  XNOR2_X1 U2803 ( .A(n2750), .B(n5105), .ZN(n4337) );
  NAND2_X1 U2804 ( .A1(n4337), .A2(n4553), .ZN(n4336) );
  NAND2_X1 U2805 ( .A1(n2634), .A2(n2753), .ZN(n2632) );
  AND2_X1 U2806 ( .A1(n2632), .A2(n2532), .ZN(n2629) );
  AND2_X1 U2807 ( .A1(n4199), .A2(DATAI_30_), .ZN(n5240) );
  AND2_X1 U2808 ( .A1(n4199), .A2(DATAI_29_), .ZN(n4374) );
  AND2_X1 U2809 ( .A1(n4192), .A2(n4185), .ZN(n4382) );
  INV_X1 U2810 ( .A(n4161), .ZN(n4415) );
  OR2_X1 U2811 ( .A1(n4432), .A2(n4433), .ZN(n4430) );
  AND2_X1 U2812 ( .A1(n4199), .A2(DATAI_25_), .ZN(n4424) );
  AND2_X1 U2813 ( .A1(n4402), .A2(n4180), .ZN(n4433) );
  NOR2_X1 U2814 ( .A1(n3782), .A2(n4095), .ZN(n3793) );
  NAND2_X1 U2815 ( .A1(n4449), .A2(n4450), .ZN(n4448) );
  NOR2_X1 U2816 ( .A1(n4473), .A2(n4452), .ZN(n4444) );
  AOI21_X1 U2817 ( .B1(n4459), .B2(n4409), .A(n3781), .ZN(n4443) );
  NOR2_X1 U2818 ( .A1(n4178), .A2(n4182), .ZN(n4450) );
  NAND2_X1 U2819 ( .A1(n4487), .A2(n4489), .ZN(n4488) );
  OR2_X1 U2820 ( .A1(n4177), .A2(n3845), .ZN(n4465) );
  AND2_X1 U2821 ( .A1(n4199), .A2(DATAI_22_), .ZN(n4480) );
  AND2_X1 U2822 ( .A1(n3777), .A2(n3776), .ZN(n4482) );
  AND2_X1 U2823 ( .A1(n3751), .A2(REG3_REG_20__SCAN_IN), .ZN(n3753) );
  NAND2_X1 U2824 ( .A1(n4199), .A2(DATAI_20_), .ZN(n4522) );
  AND2_X1 U2825 ( .A1(n4165), .A2(n4174), .ZN(n4515) );
  INV_X1 U2826 ( .A(REG3_REG_19__SCAN_IN), .ZN(n3880) );
  INV_X1 U2827 ( .A(n5204), .ZN(n5193) );
  INV_X1 U2828 ( .A(n5161), .ZN(n4539) );
  INV_X1 U2829 ( .A(n5127), .ZN(n5142) );
  INV_X1 U2830 ( .A(REG3_REG_17__SCAN_IN), .ZN(n3732) );
  INV_X1 U2831 ( .A(n3712), .ZN(n3728) );
  NAND2_X1 U2832 ( .A1(n4555), .A2(n3829), .ZN(n2546) );
  NOR2_X2 U2833 ( .A1(n3676), .A2(n5039), .ZN(n3706) );
  NAND2_X1 U2834 ( .A1(n3696), .A2(n5081), .ZN(n5085) );
  INV_X1 U2835 ( .A(n4221), .ZN(n5081) );
  OR2_X1 U2836 ( .A1(n4322), .A2(n5022), .ZN(n3663) );
  AOI21_X1 U2837 ( .B1(n2585), .B2(n2588), .A(n2583), .ZN(n2582) );
  INV_X1 U2838 ( .A(n2585), .ZN(n2584) );
  NOR2_X1 U2839 ( .A1(n3887), .A2(n3889), .ZN(n2583) );
  AND2_X1 U2840 ( .A1(n3589), .A2(REG3_REG_10__SCAN_IN), .ZN(n3608) );
  INV_X1 U2841 ( .A(n4053), .ZN(n3887) );
  OR2_X1 U2842 ( .A1(n4657), .A2(n2955), .ZN(n5175) );
  NAND2_X1 U2843 ( .A1(n3607), .A2(n4278), .ZN(n3623) );
  NOR2_X1 U2844 ( .A1(n3561), .A2(n3595), .ZN(n3589) );
  NAND2_X1 U2845 ( .A1(n4950), .A2(n4969), .ZN(n2554) );
  OR2_X1 U2846 ( .A1(n3513), .A2(n3512), .ZN(n3561) );
  AND2_X1 U2847 ( .A1(n4965), .A2(n3602), .ZN(n4228) );
  NOR2_X1 U2848 ( .A1(n3558), .A2(n3577), .ZN(n4963) );
  INV_X1 U2849 ( .A(n4272), .ZN(n3528) );
  NAND2_X1 U2850 ( .A1(n2542), .A2(n2528), .ZN(n3049) );
  INV_X1 U2851 ( .A(n4878), .ZN(n2542) );
  OR2_X1 U2852 ( .A1(n4878), .A2(n4879), .ZN(n4876) );
  INV_X1 U2853 ( .A(n5237), .ZN(n5229) );
  OR2_X1 U2854 ( .A1(n2874), .A2(n4832), .ZN(n5237) );
  INV_X1 U2855 ( .A(n5175), .ZN(n4511) );
  INV_X1 U2856 ( .A(n2906), .ZN(n4832) );
  INV_X1 U2857 ( .A(n4370), .ZN(n2538) );
  NOR2_X1 U2858 ( .A1(n2523), .A2(n2589), .ZN(n4962) );
  INV_X1 U2859 ( .A(n3600), .ZN(n2589) );
  NOR2_X1 U2860 ( .A1(n2563), .A2(n3542), .ZN(n2558) );
  INV_X1 U2861 ( .A(n5221), .ZN(n5169) );
  NAND2_X1 U2862 ( .A1(n4561), .A2(n4861), .ZN(n5221) );
  NOR2_X1 U2863 ( .A1(n4569), .A2(n4568), .ZN(n4607) );
  NAND2_X1 U2864 ( .A1(n2779), .A2(n3192), .ZN(n2776) );
  XNOR2_X1 U2865 ( .A(n2766), .B(n3387), .ZN(n2895) );
  XNOR2_X1 U2866 ( .A(n2769), .B(n3188), .ZN(n2849) );
  NAND2_X1 U2867 ( .A1(n2773), .A2(IR_REG_31__SCAN_IN), .ZN(n2769) );
  NAND2_X1 U2868 ( .A1(n2774), .A2(n2773), .ZN(n2913) );
  INV_X1 U2869 ( .A(IR_REG_10__SCAN_IN), .ZN(n2557) );
  AND2_X1 U2870 ( .A1(n2535), .A2(n2534), .ZN(n2651) );
  NOR2_X1 U2871 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_2__SCAN_IN), .ZN(n2535)
         );
  NOR2_X1 U2872 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2534)
         );
  INV_X1 U2873 ( .A(IR_REG_2__SCAN_IN), .ZN(n2683) );
  INV_X1 U2874 ( .A(IR_REG_4__SCAN_IN), .ZN(n2708) );
  INV_X1 U2875 ( .A(IR_REG_3__SCAN_IN), .ZN(n3155) );
  XNOR2_X1 U2876 ( .A(n2691), .B(n3339), .ZN(n2692) );
  INV_X1 U2877 ( .A(n3508), .ZN(n3506) );
  AOI21_X1 U2878 ( .B1(n4079), .B2(n2671), .A(n2670), .ZN(n4032) );
  AND2_X1 U2879 ( .A1(n3820), .A2(n3813), .ZN(n4392) );
  INV_X1 U2880 ( .A(n2667), .ZN(n2666) );
  OAI22_X1 U2881 ( .A1(n4031), .A2(n4008), .B1(n4013), .B2(n4014), .ZN(n2667)
         );
  OAI22_X1 U2882 ( .A1(n2933), .A2(n2932), .B1(n4016), .B2(n2931), .ZN(n3466)
         );
  INV_X1 U2883 ( .A(n3465), .ZN(n2938) );
  NAND2_X1 U2884 ( .A1(n4116), .A2(n4114), .ZN(n2650) );
  INV_X1 U2885 ( .A(n2664), .ZN(n5021) );
  INV_X1 U2886 ( .A(n2660), .ZN(n2659) );
  OAI21_X1 U2887 ( .B1(n3896), .B2(n2662), .A(n2661), .ZN(n2660) );
  OAI21_X2 U2888 ( .B1(n2482), .B2(n2878), .A(n2877), .ZN(n2950) );
  INV_X1 U2889 ( .A(IR_REG_0__SCAN_IN), .ZN(n2878) );
  NAND2_X1 U2890 ( .A1(n2482), .A2(DATAI_0_), .ZN(n2877) );
  MUX2_X1 U2891 ( .A(n5034), .B(DATAI_13_), .S(n2977), .Z(n5039) );
  AND2_X1 U2892 ( .A1(n4049), .A2(n2509), .ZN(n4999) );
  AOI21_X1 U2893 ( .B1(n5126), .B2(n5125), .A(n2507), .ZN(n5159) );
  INV_X1 U2894 ( .A(n4026), .ZN(n4151) );
  NAND2_X1 U2895 ( .A1(n4079), .A2(n4004), .ZN(n4158) );
  AND2_X1 U2896 ( .A1(n4199), .A2(DATAI_26_), .ZN(n4161) );
  OR2_X1 U2897 ( .A1(n3926), .A2(n3925), .ZN(n3927) );
  NOR2_X2 U2898 ( .A1(n2921), .A2(n2920), .ZN(n5190) );
  INV_X1 U2899 ( .A(n5185), .ZN(n5160) );
  INV_X1 U2900 ( .A(n5186), .ZN(n5162) );
  INV_X1 U2901 ( .A(n4201), .ZN(n4311) );
  INV_X1 U2902 ( .A(n4097), .ZN(n4453) );
  NAND2_X1 U2903 ( .A1(n3790), .A2(n3789), .ZN(n4410) );
  INV_X1 U2904 ( .A(n4482), .ZN(n4314) );
  INV_X1 U2905 ( .A(n4071), .ZN(n4315) );
  NAND4_X1 U2906 ( .A1(n3717), .A2(n3716), .A3(n3715), .A4(n3714), .ZN(n4520)
         );
  INV_X1 U2907 ( .A(n4238), .ZN(n4325) );
  INV_X1 U2908 ( .A(n3541), .ZN(n4329) );
  AOI21_X1 U2909 ( .B1(REG0_REG_2__SCAN_IN), .B2(n2939), .A(n2940), .ZN(n2943)
         );
  INV_X1 U2910 ( .A(n2602), .ZN(n4796) );
  AND2_X1 U2911 ( .A1(n4676), .A2(REG1_REG_3__SCAN_IN), .ZN(n4677) );
  INV_X1 U2912 ( .A(n2594), .ZN(n4816) );
  OAI21_X1 U2913 ( .B1(n4817), .B2(n2592), .A(n2591), .ZN(n4688) );
  NAND2_X1 U2914 ( .A1(n2595), .A2(REG1_REG_4__SCAN_IN), .ZN(n2592) );
  INV_X1 U2915 ( .A(n4689), .ZN(n2595) );
  INV_X1 U2916 ( .A(n2807), .ZN(n2593) );
  NAND2_X1 U2917 ( .A1(n2606), .A2(REG1_REG_6__SCAN_IN), .ZN(n2605) );
  NAND2_X1 U2918 ( .A1(n2811), .A2(n2606), .ZN(n2604) );
  INV_X1 U2919 ( .A(n4712), .ZN(n2606) );
  NAND2_X1 U2920 ( .A1(n2619), .A2(n2620), .ZN(n4715) );
  NAND2_X1 U2921 ( .A1(n2597), .A2(n2596), .ZN(n4720) );
  NAND2_X1 U2922 ( .A1(n2637), .A2(n2635), .ZN(n4724) );
  NOR2_X1 U2923 ( .A1(n4742), .A2(n4741), .ZN(n4740) );
  NOR2_X1 U2924 ( .A1(n4730), .A2(n2493), .ZN(n4742) );
  OAI21_X1 U2925 ( .B1(n4751), .B2(n2600), .A(n2599), .ZN(n4763) );
  NAND2_X1 U2926 ( .A1(n2601), .A2(REG1_REG_12__SCAN_IN), .ZN(n2600) );
  NAND2_X1 U2927 ( .A1(n2820), .A2(n2601), .ZN(n2599) );
  INV_X1 U2928 ( .A(n4764), .ZN(n2601) );
  NOR2_X1 U2929 ( .A1(n2745), .A2(n4772), .ZN(n4781) );
  OAI211_X1 U2930 ( .C1(n2828), .C2(n4343), .A(n2607), .B(n2829), .ZN(n2833)
         );
  NAND2_X1 U2931 ( .A1(n4334), .A2(n2608), .ZN(n2607) );
  NOR2_X1 U2932 ( .A1(n4343), .A2(REG1_REG_16__SCAN_IN), .ZN(n2608) );
  NAND2_X1 U2933 ( .A1(n2630), .A2(n2632), .ZN(n3875) );
  OR2_X1 U2934 ( .A1(n2831), .A2(n4808), .ZN(n4827) );
  XNOR2_X1 U2935 ( .A(n3879), .B(n3878), .ZN(n3884) );
  NAND2_X1 U2936 ( .A1(n2630), .A2(n2629), .ZN(n3879) );
  INV_X1 U2937 ( .A(n4363), .ZN(n4357) );
  NAND2_X1 U2938 ( .A1(n4371), .A2(n4370), .ZN(n4565) );
  NAND2_X1 U2939 ( .A1(n2516), .A2(n2576), .ZN(n4530) );
  INV_X1 U2940 ( .A(n2574), .ZN(n5139) );
  AOI21_X1 U2941 ( .B1(n3727), .B2(n2575), .A(n2500), .ZN(n2574) );
  INV_X1 U2942 ( .A(n2580), .ZN(n2575) );
  OAI21_X1 U2943 ( .B1(n3557), .B2(n2588), .A(n2587), .ZN(n3635) );
  NAND2_X1 U2944 ( .A1(n3069), .A2(n3068), .ZN(n3544) );
  INV_X1 U2945 ( .A(n5103), .ZN(n5144) );
  INV_X1 U2946 ( .A(n5216), .ZN(n5136) );
  NAND2_X1 U2947 ( .A1(n2976), .A2(n2975), .ZN(n3022) );
  INV_X1 U2948 ( .A(n4566), .ZN(n2909) );
  AND2_X2 U2949 ( .A1(n4607), .A2(n4570), .ZN(n5253) );
  AOI21_X1 U2950 ( .B1(n5233), .B2(n5249), .A(n5232), .ZN(n5236) );
  AND2_X2 U2951 ( .A1(n4607), .A2(n4606), .ZN(n5257) );
  NAND2_X1 U2952 ( .A1(n2966), .A2(n2910), .ZN(n4652) );
  INV_X1 U2953 ( .A(IR_REG_29__SCAN_IN), .ZN(n2862) );
  XNOR2_X1 U2954 ( .A(n2779), .B(IR_REG_26__SCAN_IN), .ZN(n4622) );
  INV_X1 U2955 ( .A(n2895), .ZN(n3461) );
  INV_X1 U2956 ( .A(n2954), .ZN(n4624) );
  XNOR2_X1 U2957 ( .A(n2787), .B(IR_REG_21__SCAN_IN), .ZN(n4625) );
  INV_X1 U2958 ( .A(n4840), .ZN(n4626) );
  XNOR2_X1 U2959 ( .A(n2755), .B(IR_REG_18__SCAN_IN), .ZN(n5154) );
  INV_X1 U2960 ( .A(n3572), .ZN(n4727) );
  XNOR2_X1 U2961 ( .A(n2695), .B(IR_REG_2__SCAN_IN), .ZN(n4858) );
  INV_X1 U2962 ( .A(n2692), .ZN(n4673) );
  INV_X1 U2963 ( .A(n4628), .ZN(n2837) );
  NAND2_X1 U2964 ( .A1(n3828), .A2(n4840), .ZN(n3867) );
  NAND2_X1 U2965 ( .A1(n2541), .A2(n2539), .ZN(U3515) );
  OR2_X1 U2966 ( .A1(n5257), .A2(n2540), .ZN(n2539) );
  INV_X1 U2967 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2540) );
  INV_X1 U2968 ( .A(n2874), .ZN(n4841) );
  XNOR2_X2 U2969 ( .A(n2845), .B(n3374), .ZN(n2874) );
  INV_X1 U2970 ( .A(n4108), .ZN(n2544) );
  AND2_X1 U2971 ( .A1(n2658), .A2(n2522), .ZN(n2488) );
  NOR2_X1 U2972 ( .A1(n4753), .A2(n2735), .ZN(n4761) );
  OR2_X1 U2973 ( .A1(n4316), .A2(n5161), .ZN(n2489) );
  AND2_X1 U2974 ( .A1(n2648), .A2(n2646), .ZN(n2490) );
  OR2_X1 U2975 ( .A1(n2813), .A2(n4942), .ZN(n2491) );
  OR2_X1 U2976 ( .A1(n2725), .A2(n4942), .ZN(n2492) );
  AND2_X1 U2977 ( .A1(n2727), .A2(n4737), .ZN(n2493) );
  OR2_X1 U2978 ( .A1(n4473), .A2(n2547), .ZN(n2494) );
  NOR2_X1 U2979 ( .A1(n4680), .A2(n2706), .ZN(n2710) );
  NOR2_X1 U2980 ( .A1(n4396), .A2(n2494), .ZN(n2550) );
  AND2_X1 U2981 ( .A1(n4572), .A2(n3866), .ZN(n2495) );
  AND2_X1 U2982 ( .A1(n4562), .A2(n5221), .ZN(n2496) );
  NOR2_X1 U2983 ( .A1(n4907), .A2(n4141), .ZN(n2497) );
  NOR2_X1 U2984 ( .A1(n4781), .A2(n4782), .ZN(n2498) );
  INV_X1 U2985 ( .A(n2572), .ZN(n2571) );
  NOR2_X1 U2986 ( .A1(n4532), .A2(n2573), .ZN(n2572) );
  AND2_X1 U2987 ( .A1(n3792), .A2(n3791), .ZN(n2499) );
  NOR2_X1 U2988 ( .A1(n4318), .A2(n5109), .ZN(n2500) );
  INV_X1 U2989 ( .A(IR_REG_25__SCAN_IN), .ZN(n3387) );
  INV_X1 U2990 ( .A(IR_REG_9__SCAN_IN), .ZN(n2685) );
  NAND2_X1 U2991 ( .A1(n3600), .A2(n3601), .ZN(n2501) );
  AND2_X1 U2992 ( .A1(n4232), .A2(n3543), .ZN(n2502) );
  NOR2_X1 U2993 ( .A1(n4346), .A2(n2753), .ZN(n2503) );
  AND2_X1 U2994 ( .A1(n2676), .A2(n2760), .ZN(n2504) );
  INV_X1 U2995 ( .A(n2615), .ZN(n2744) );
  NAND2_X1 U2996 ( .A1(n2694), .A2(n2683), .ZN(n2701) );
  AND2_X1 U2997 ( .A1(n2504), .A2(n2861), .ZN(n2505) );
  NOR2_X1 U2998 ( .A1(n2767), .A2(n2764), .ZN(n2506) );
  NAND2_X1 U2999 ( .A1(n2687), .A2(n2685), .ZN(n2736) );
  AND2_X1 U3000 ( .A1(n3945), .A2(n3944), .ZN(n2507) );
  AND2_X1 U3001 ( .A1(n4498), .A2(n3970), .ZN(n4487) );
  OR2_X1 U3002 ( .A1(n5122), .A2(n4555), .ZN(n2508) );
  AND2_X1 U3003 ( .A1(n3901), .A2(n2663), .ZN(n2509) );
  AND2_X1 U3004 ( .A1(n2716), .A2(n2684), .ZN(n2687) );
  AND2_X1 U3005 ( .A1(n2687), .A2(n2672), .ZN(n2742) );
  OR2_X1 U3006 ( .A1(n4156), .A2(n4155), .ZN(n2510) );
  NOR2_X1 U3007 ( .A1(n3826), .A2(n2546), .ZN(n2545) );
  OR2_X1 U3008 ( .A1(n4389), .A2(n4355), .ZN(n2511) );
  NOR2_X1 U3009 ( .A1(n4750), .A2(n2820), .ZN(n2512) );
  NAND2_X1 U3010 ( .A1(n2687), .A2(n2674), .ZN(n2739) );
  OR2_X1 U3011 ( .A1(n2507), .A2(n2655), .ZN(n2513) );
  INV_X1 U3012 ( .A(n2757), .ZN(n2761) );
  INV_X1 U3013 ( .A(n4555), .ZN(n5109) );
  NAND2_X1 U3014 ( .A1(n3977), .A2(n4123), .ZN(n2514) );
  AND2_X1 U3015 ( .A1(n3993), .A2(n2643), .ZN(n2515) );
  INV_X1 U3016 ( .A(n2579), .ZN(n2578) );
  NOR2_X1 U3017 ( .A1(n3738), .A2(n2500), .ZN(n2579) );
  INV_X1 U3018 ( .A(n4008), .ZN(n2670) );
  OR2_X1 U3019 ( .A1(n3727), .A2(n2578), .ZN(n2516) );
  OR2_X1 U3020 ( .A1(n4721), .A2(n4959), .ZN(n2517) );
  NOR2_X1 U3021 ( .A1(n4761), .A2(n4762), .ZN(n2518) );
  NAND2_X1 U3022 ( .A1(n4727), .A2(REG1_REG_9__SCAN_IN), .ZN(n2519) );
  NAND2_X1 U3023 ( .A1(n4727), .A2(REG2_REG_9__SCAN_IN), .ZN(n2520) );
  INV_X1 U3024 ( .A(IR_REG_31__SCAN_IN), .ZN(n2765) );
  AND2_X2 U3025 ( .A1(n2969), .A2(n5216), .ZN(n5246) );
  NAND2_X1 U3026 ( .A1(n2562), .A2(n2559), .ZN(n3554) );
  NOR2_X1 U3027 ( .A1(n3826), .A2(n5089), .ZN(n2521) );
  NOR2_X1 U3028 ( .A1(n3558), .A2(n2554), .ZN(n3618) );
  OR2_X1 U3029 ( .A1(n3949), .A2(n3950), .ZN(n2522) );
  INV_X1 U3030 ( .A(n4096), .ZN(n4452) );
  AND2_X1 U3031 ( .A1(n3556), .A2(n3555), .ZN(n2523) );
  AND2_X1 U3032 ( .A1(n2562), .A2(n2558), .ZN(n2524) );
  AND2_X1 U3033 ( .A1(n2598), .A2(n2491), .ZN(n2525) );
  AND2_X1 U3034 ( .A1(n2638), .A2(n2492), .ZN(n2526) );
  AND2_X1 U3035 ( .A1(n4258), .A2(n4833), .ZN(n3012) );
  OR2_X1 U3036 ( .A1(n2743), .A2(n2761), .ZN(n5052) );
  INV_X1 U3037 ( .A(IR_REG_1__SCAN_IN), .ZN(n3339) );
  NOR2_X1 U3038 ( .A1(n4697), .A2(n2811), .ZN(n2527) );
  AND2_X1 U3039 ( .A1(n3013), .A2(n2544), .ZN(n2528) );
  AND2_X1 U3040 ( .A1(n2634), .A2(n2633), .ZN(n2529) );
  AND2_X1 U3041 ( .A1(n2594), .A2(n2593), .ZN(n2530) );
  AND2_X1 U3042 ( .A1(n4789), .A2(REG2_REG_15__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U3043 ( .A1(n5154), .A2(REG2_REG_18__SCAN_IN), .ZN(n2532) );
  AND2_X1 U3044 ( .A1(n2624), .A2(n2623), .ZN(n2533) );
  NAND2_X1 U3045 ( .A1(n4608), .A2(n5257), .ZN(n2541) );
  NOR2_X2 U3046 ( .A1(n4878), .A2(n2543), .ZN(n3070) );
  NAND3_X1 U3047 ( .A1(n3013), .A2(n2544), .A3(n3051), .ZN(n2543) );
  INV_X1 U3048 ( .A(n2550), .ZN(n4575) );
  NAND2_X1 U3049 ( .A1(n2504), .A2(n2761), .ZN(n2552) );
  OR2_X2 U3050 ( .A1(n3636), .A2(n5006), .ZN(n3656) );
  NAND2_X1 U3051 ( .A1(n3618), .A2(n3887), .ZN(n3636) );
  XNOR2_X2 U3052 ( .A(n2949), .B(n4258), .ZN(n2996) );
  XNOR2_X2 U3053 ( .A(n2780), .B(IR_REG_28__SCAN_IN), .ZN(n2791) );
  NAND2_X1 U3054 ( .A1(n2556), .A2(n2976), .ZN(n3020) );
  NAND2_X1 U3055 ( .A1(n3020), .A2(n2980), .ZN(n4868) );
  NAND3_X1 U3056 ( .A1(n3166), .A2(n3170), .A3(n2557), .ZN(n2675) );
  NAND2_X1 U3057 ( .A1(n3047), .A2(n2502), .ZN(n2562) );
  INV_X1 U3058 ( .A(n2569), .ZN(n5199) );
  NAND2_X1 U3059 ( .A1(n3727), .A2(n3726), .ZN(n4546) );
  OR2_X1 U3060 ( .A1(n4549), .A2(n5142), .ZN(n2581) );
  NAND2_X1 U3061 ( .A1(n2807), .A2(n2595), .ZN(n2591) );
  INV_X1 U3062 ( .A(n2598), .ZN(n2853) );
  OAI21_X1 U3063 ( .B1(n4698), .B2(n2605), .A(n2604), .ZN(n4711) );
  NAND2_X1 U3064 ( .A1(n4333), .A2(n2828), .ZN(n4344) );
  NAND2_X1 U3065 ( .A1(n4334), .A2(n5118), .ZN(n4333) );
  NAND2_X1 U3066 ( .A1(n4797), .A2(n2700), .ZN(n2704) );
  NAND2_X1 U3067 ( .A1(n2610), .A2(n2699), .ZN(n4797) );
  INV_X1 U3068 ( .A(n4800), .ZN(n2610) );
  NAND2_X1 U3069 ( .A1(n4753), .A2(n2614), .ZN(n2613) );
  NAND2_X1 U3070 ( .A1(n4772), .A2(n2618), .ZN(n2616) );
  AOI21_X1 U3071 ( .B1(n2745), .B2(n2618), .A(n2531), .ZN(n2617) );
  INV_X1 U3072 ( .A(n2624), .ZN(n4700) );
  INV_X1 U3073 ( .A(n2719), .ZN(n2623) );
  INV_X1 U3074 ( .A(n2628), .ZN(n2734) );
  INV_X1 U3075 ( .A(n4348), .ZN(n2631) );
  NOR2_X1 U3076 ( .A1(n4348), .A2(n4347), .ZN(n4346) );
  INV_X1 U3077 ( .A(n2792), .ZN(n2634) );
  INV_X1 U3078 ( .A(n2638), .ZN(n2850) );
  NAND2_X1 U3079 ( .A1(n2641), .A2(IR_REG_31__SCAN_IN), .ZN(n2695) );
  INV_X1 U3080 ( .A(n2641), .ZN(n2694) );
  OR2_X1 U3081 ( .A1(n4116), .A2(n2647), .ZN(n2642) );
  NAND2_X1 U3082 ( .A1(n4116), .A2(n2645), .ZN(n2644) );
  NAND4_X1 U3083 ( .A1(n2694), .A2(n3155), .A3(n2683), .A4(n2708), .ZN(n2712)
         );
  AND2_X2 U3084 ( .A1(n2651), .A2(n2694), .ZN(n2716) );
  NAND2_X1 U3085 ( .A1(n4079), .A2(n2668), .ZN(n2665) );
  NAND2_X1 U3086 ( .A1(n2665), .A2(n2666), .ZN(n4021) );
  NAND3_X1 U3087 ( .A1(n4104), .A2(n3491), .A3(n2497), .ZN(n3509) );
  NAND2_X1 U3088 ( .A1(n2761), .A2(n2505), .ZN(n2866) );
  NAND2_X1 U3089 ( .A1(n2761), .A2(n2760), .ZN(n2767) );
  XNOR2_X1 U3090 ( .A(n4414), .B(n4413), .ZN(n4579) );
  NAND2_X1 U3091 ( .A1(n4430), .A2(n4411), .ZN(n4414) );
  INV_X1 U3092 ( .A(n4332), .ZN(n3477) );
  NAND2_X1 U3093 ( .A1(n3853), .A2(n4353), .ZN(n3854) );
  NAND2_X1 U3094 ( .A1(n3012), .A2(n3029), .ZN(n4878) );
  NOR2_X1 U3095 ( .A1(n5241), .A2(n5240), .ZN(n5242) );
  AND2_X1 U3096 ( .A1(n2951), .A2(n2950), .ZN(n2952) );
  NAND2_X1 U3097 ( .A1(n3468), .A2(n2950), .ZN(n2883) );
  NOR2_X2 U3098 ( .A1(n3853), .A2(n4353), .ZN(n4362) );
  OR2_X1 U3099 ( .A1(n3864), .A2(n3863), .ZN(n2677) );
  AND2_X1 U3100 ( .A1(n2948), .A2(n2947), .ZN(n5091) );
  INV_X1 U3101 ( .A(n5091), .ZN(n5207) );
  AND2_X1 U3102 ( .A1(n3465), .A2(n3464), .ZN(n2678) );
  AND2_X1 U3103 ( .A1(n2799), .A2(n2798), .ZN(n2679) );
  NAND2_X1 U3104 ( .A1(n4317), .A2(n5142), .ZN(n2680) );
  OR2_X1 U3105 ( .A1(n3778), .A2(n4465), .ZN(n4408) );
  INV_X1 U3106 ( .A(n5017), .ZN(n2818) );
  CLKBUF_X3 U3107 ( .A(n2939), .Z(n3858) );
  AND2_X1 U3108 ( .A1(n4331), .A2(n4108), .ZN(n2681) );
  NOR2_X1 U3109 ( .A1(n4822), .A2(n4821), .ZN(n4820) );
  INV_X1 U3110 ( .A(n2485), .ZN(n3762) );
  AND2_X1 U3111 ( .A1(n2942), .A2(n2941), .ZN(n2682) );
  AND2_X1 U3112 ( .A1(n4995), .A2(REG2_REG_11__SCAN_IN), .ZN(n2730) );
  INV_X1 U3113 ( .A(n3899), .ZN(n3900) );
  AND2_X1 U3114 ( .A1(n4627), .A2(REG2_REG_17__SCAN_IN), .ZN(n2753) );
  INV_X1 U3115 ( .A(n4234), .ZN(n3530) );
  NAND2_X1 U3116 ( .A1(n3510), .A2(n3511), .ZN(n3505) );
  NAND2_X1 U3117 ( .A1(n3488), .A2(n3490), .ZN(n3491) );
  OR2_X1 U3118 ( .A1(n3913), .A2(n3912), .ZN(n3914) );
  INV_X1 U3119 ( .A(n4801), .ZN(n2699) );
  NAND2_X1 U3120 ( .A1(n4319), .A2(n5089), .ZN(n3726) );
  INV_X1 U3121 ( .A(n4879), .ZN(n3013) );
  INV_X1 U3122 ( .A(IR_REG_22__SCAN_IN), .ZN(n2762) );
  NOR2_X1 U3123 ( .A1(n3506), .A2(n3505), .ZN(n3507) );
  INV_X1 U3124 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3770) );
  INV_X1 U3125 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3040) );
  AND2_X1 U3126 ( .A1(n3857), .A2(n3821), .ZN(n4023) );
  OR2_X1 U3127 ( .A1(n4627), .A2(REG1_REG_17__SCAN_IN), .ZN(n2829) );
  AND2_X1 U3128 ( .A1(n3753), .A2(REG3_REG_21__SCAN_IN), .ZN(n3766) );
  INV_X1 U3129 ( .A(n4228), .ZN(n3555) );
  AND2_X1 U3130 ( .A1(n4199), .A2(DATAI_27_), .ZN(n4396) );
  INV_X1 U3131 ( .A(n5082), .ZN(n5086) );
  INV_X1 U3132 ( .A(n4137), .ZN(n3029) );
  INV_X1 U3133 ( .A(IR_REG_27__SCAN_IN), .ZN(n3391) );
  AND2_X1 U3134 ( .A1(n4050), .A2(n4048), .ZN(n3896) );
  INV_X1 U3135 ( .A(REG3_REG_8__SCAN_IN), .ZN(n3512) );
  NAND2_X1 U3136 ( .A1(n4199), .A2(DATAI_21_), .ZN(n3970) );
  NAND2_X1 U3137 ( .A1(n4199), .A2(DATAI_24_), .ZN(n4096) );
  AND2_X1 U3138 ( .A1(n4103), .A2(n4105), .ZN(n3487) );
  AOI22_X1 U3139 ( .A1(n4010), .A2(n2951), .B1(n2881), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2882) );
  NAND2_X1 U3140 ( .A1(n3766), .A2(REG3_REG_22__SCAN_IN), .ZN(n3771) );
  AND2_X1 U3141 ( .A1(n2911), .A2(n5216), .ZN(n5185) );
  AOI21_X1 U3142 ( .B1(n4737), .B2(n2815), .A(n4733), .ZN(n4745) );
  INV_X1 U3143 ( .A(n3877), .ZN(n3878) );
  INV_X1 U3144 ( .A(n4412), .ZN(n4413) );
  AND2_X1 U3145 ( .A1(n4463), .A2(n3842), .ZN(n4485) );
  OR2_X1 U3146 ( .A1(n4512), .A2(n5193), .ZN(n3750) );
  INV_X1 U3147 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3595) );
  OR2_X1 U31480 ( .A1(n2969), .A2(n2968), .ZN(n5196) );
  AND2_X1 U31490 ( .A1(n4657), .A2(n2922), .ZN(n5177) );
  AND2_X1 U3150 ( .A1(n3689), .A2(n3686), .ZN(n4230) );
  INV_X1 U3151 ( .A(n5177), .ZN(n5121) );
  INV_X1 U3152 ( .A(IR_REG_15__SCAN_IN), .ZN(n2758) );
  AND2_X1 U3153 ( .A1(n4199), .A2(DATAI_23_), .ZN(n4475) );
  INV_X1 U3154 ( .A(n3970), .ZN(n4506) );
  NAND2_X1 U3155 ( .A1(n3728), .A2(REG3_REG_16__SCAN_IN), .ZN(n3733) );
  NOR2_X1 U3156 ( .A1(n3733), .A2(n3732), .ZN(n3739) );
  INV_X1 U3157 ( .A(n5192), .ZN(n4160) );
  NOR2_X1 U3158 ( .A1(n3669), .A2(n3668), .ZN(n3698) );
  AND4_X1 U3159 ( .A1(n3825), .A2(n3824), .A3(n3823), .A4(n3822), .ZN(n4389)
         );
  AND2_X1 U3160 ( .A1(n3741), .A2(n3740), .ZN(n5176) );
  INV_X1 U3161 ( .A(n4827), .ZN(n4804) );
  AND2_X1 U3162 ( .A1(n4660), .A2(n4305), .ZN(n4824) );
  NOR2_X1 U3163 ( .A1(n3742), .A2(n3880), .ZN(n3751) );
  AND2_X1 U3164 ( .A1(n4251), .A2(n3685), .ZN(n4229) );
  INV_X1 U3166 ( .A(n5196), .ZN(n5244) );
  AOI21_X1 U3167 ( .B1(n2899), .B2(n3399), .A(n2884), .ZN(n4570) );
  INV_X1 U3168 ( .A(n5219), .ZN(n5249) );
  INV_X1 U3169 ( .A(n4570), .ZN(n4606) );
  AND2_X1 U3170 ( .A1(n2795), .A2(n2794), .ZN(n4815) );
  NAND2_X1 U3171 ( .A1(n2908), .A2(n2907), .ZN(n5186) );
  NAND2_X1 U3172 ( .A1(n3520), .A2(STATE_REG_SCAN_IN), .ZN(n5192) );
  INV_X1 U3173 ( .A(n4386), .ZN(n4425) );
  INV_X1 U3174 ( .A(n5122), .ZN(n4318) );
  OR2_X1 U3175 ( .A1(n2831), .A2(n4658), .ZN(n4793) );
  NAND2_X1 U3176 ( .A1(n2910), .A2(n2909), .ZN(n5216) );
  INV_X1 U3178 ( .A(n5253), .ZN(n5251) );
  INV_X1 U3179 ( .A(n5257), .ZN(n5254) );
  AND2_X1 U3180 ( .A1(n2896), .A2(n2849), .ZN(n2884) );
  AND2_X1 U3181 ( .A1(n2913), .A2(STATE_REG_SCAN_IN), .ZN(n4628) );
  AND2_X1 U3182 ( .A1(n2752), .A2(n2747), .ZN(n4789) );
  AND2_X1 U3183 ( .A1(n2707), .A2(n2703), .ZN(n4685) );
  INV_X4 U3184 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X2 U3185 ( .A(IR_REG_8__SCAN_IN), .ZN(n3351) );
  NAND2_X1 U3186 ( .A1(n2736), .A2(IR_REG_31__SCAN_IN), .ZN(n2686) );
  XNOR2_X1 U3187 ( .A(n2686), .B(IR_REG_10__SCAN_IN), .ZN(n4737) );
  NOR2_X1 U3188 ( .A1(n2687), .A2(n2765), .ZN(n2688) );
  MUX2_X1 U3189 ( .A(n2765), .B(n2688), .S(IR_REG_9__SCAN_IN), .Z(n2689) );
  INV_X1 U3190 ( .A(n2689), .ZN(n2690) );
  NAND2_X1 U3191 ( .A1(n2690), .A2(n2736), .ZN(n3572) );
  NAND2_X1 U3192 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2691)
         );
  XNOR2_X1 U3193 ( .A(n2692), .B(REG2_REG_1__SCAN_IN), .ZN(n4664) );
  AND2_X1 U3194 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4807)
         );
  NAND2_X1 U3195 ( .A1(n4664), .A2(n4807), .ZN(n4663) );
  NAND2_X1 U3196 ( .A1(n4673), .A2(REG2_REG_1__SCAN_IN), .ZN(n2693) );
  NAND2_X1 U3197 ( .A1(n4858), .A2(REG2_REG_2__SCAN_IN), .ZN(n2700) );
  INV_X1 U3198 ( .A(n4858), .ZN(n2697) );
  INV_X1 U3199 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2696) );
  NAND2_X1 U3200 ( .A1(n2700), .A2(n2698), .ZN(n4800) );
  NAND2_X1 U3201 ( .A1(n2701), .A2(IR_REG_31__SCAN_IN), .ZN(n2702) );
  NAND2_X1 U3202 ( .A1(n2702), .A2(n3155), .ZN(n2707) );
  OR2_X1 U3203 ( .A1(n2702), .A2(n3155), .ZN(n2703) );
  NOR2_X1 U3204 ( .A1(n2704), .A2(n4685), .ZN(n2705) );
  NAND2_X1 U3205 ( .A1(n2707), .A2(IR_REG_31__SCAN_IN), .ZN(n2709) );
  XNOR2_X1 U3206 ( .A(n2709), .B(n2708), .ZN(n4892) );
  NOR2_X1 U3207 ( .A1(n2710), .A2(n4892), .ZN(n2711) );
  XNOR2_X1 U3208 ( .A(n2710), .B(n4892), .ZN(n4822) );
  INV_X1 U3209 ( .A(REG2_REG_4__SCAN_IN), .ZN(n4821) );
  NOR2_X1 U32100 ( .A1(n2711), .A2(n4820), .ZN(n4693) );
  NAND2_X1 U32110 ( .A1(n2712), .A2(IR_REG_31__SCAN_IN), .ZN(n2713) );
  XNOR2_X1 U32120 ( .A(n2713), .B(IR_REG_5__SCAN_IN), .ZN(n4901) );
  NAND2_X1 U32130 ( .A1(n4901), .A2(REG2_REG_5__SCAN_IN), .ZN(n2714) );
  OAI21_X1 U32140 ( .B1(n4901), .B2(REG2_REG_5__SCAN_IN), .A(n2714), .ZN(n4692) );
  NOR2_X1 U32150 ( .A1(n4693), .A2(n4692), .ZN(n4691) );
  NOR2_X1 U32160 ( .A1(n4691), .A2(n2715), .ZN(n2718) );
  OR2_X1 U32170 ( .A1(n2716), .A2(n2765), .ZN(n2717) );
  XNOR2_X1 U32180 ( .A(n2717), .B(IR_REG_6__SCAN_IN), .ZN(n4923) );
  INV_X1 U32190 ( .A(n4923), .ZN(n4706) );
  NOR2_X1 U32200 ( .A1(n2718), .A2(n4706), .ZN(n2719) );
  INV_X1 U32210 ( .A(REG2_REG_6__SCAN_IN), .ZN(n4701) );
  XNOR2_X1 U32220 ( .A(n2718), .B(n4706), .ZN(n4702) );
  NAND2_X1 U32230 ( .A1(n2716), .A2(n3352), .ZN(n2720) );
  NAND2_X1 U32240 ( .A1(n2720), .A2(IR_REG_31__SCAN_IN), .ZN(n2722) );
  XNOR2_X1 U32250 ( .A(n2722), .B(IR_REG_7__SCAN_IN), .ZN(n4932) );
  NAND2_X1 U32260 ( .A1(n4932), .A2(REG2_REG_7__SCAN_IN), .ZN(n2721) );
  OAI21_X1 U32270 ( .B1(n4932), .B2(REG2_REG_7__SCAN_IN), .A(n2721), .ZN(n4716) );
  NAND2_X1 U32280 ( .A1(n2722), .A2(n3348), .ZN(n2723) );
  NAND2_X1 U32290 ( .A1(n2723), .A2(IR_REG_31__SCAN_IN), .ZN(n2724) );
  XNOR2_X1 U32300 ( .A(n2724), .B(n3351), .ZN(n4942) );
  INV_X1 U32310 ( .A(REG2_REG_8__SCAN_IN), .ZN(n2852) );
  XNOR2_X1 U32320 ( .A(n2725), .B(n4942), .ZN(n2851) );
  XNOR2_X1 U32330 ( .A(n4727), .B(REG2_REG_9__SCAN_IN), .ZN(n4725) );
  INV_X1 U32340 ( .A(n2726), .ZN(n2727) );
  XOR2_X1 U32350 ( .A(n4737), .B(n2726), .Z(n4731) );
  INV_X1 U32360 ( .A(REG2_REG_10__SCAN_IN), .ZN(n4732) );
  OR2_X1 U32370 ( .A1(n2736), .A2(IR_REG_10__SCAN_IN), .ZN(n2728) );
  NAND2_X1 U32380 ( .A1(n2728), .A2(IR_REG_31__SCAN_IN), .ZN(n2731) );
  XNOR2_X1 U32390 ( .A(n2731), .B(IR_REG_11__SCAN_IN), .ZN(n4995) );
  NAND2_X1 U32400 ( .A1(n4995), .A2(REG2_REG_11__SCAN_IN), .ZN(n2729) );
  OAI21_X1 U32410 ( .B1(n4995), .B2(REG2_REG_11__SCAN_IN), .A(n2729), .ZN(
        n4741) );
  NAND2_X1 U32420 ( .A1(n2731), .A2(n3166), .ZN(n2732) );
  NAND2_X1 U32430 ( .A1(n2732), .A2(IR_REG_31__SCAN_IN), .ZN(n2733) );
  XNOR2_X1 U32440 ( .A(n2733), .B(IR_REG_12__SCAN_IN), .ZN(n5017) );
  NOR2_X1 U32450 ( .A1(n2734), .A2(n2818), .ZN(n2735) );
  NAND2_X1 U32460 ( .A1(n2739), .A2(IR_REG_31__SCAN_IN), .ZN(n2737) );
  XNOR2_X1 U32470 ( .A(n2737), .B(IR_REG_13__SCAN_IN), .ZN(n5034) );
  NAND2_X1 U32480 ( .A1(n5034), .A2(REG2_REG_13__SCAN_IN), .ZN(n2738) );
  OAI21_X1 U32490 ( .B1(n5034), .B2(REG2_REG_13__SCAN_IN), .A(n2738), .ZN(
        n4762) );
  NOR2_X1 U32500 ( .A1(n2742), .A2(n2765), .ZN(n2740) );
  MUX2_X1 U32510 ( .A(n2765), .B(n2740), .S(IR_REG_14__SCAN_IN), .Z(n2743) );
  INV_X1 U32520 ( .A(IR_REG_14__SCAN_IN), .ZN(n2741) );
  INV_X1 U32530 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4773) );
  NOR2_X1 U32540 ( .A1(n2744), .A2(n5052), .ZN(n2745) );
  NAND2_X1 U32550 ( .A1(n2757), .A2(IR_REG_31__SCAN_IN), .ZN(n2746) );
  NAND2_X1 U32560 ( .A1(n2746), .A2(n2758), .ZN(n2752) );
  OR2_X1 U32570 ( .A1(n2746), .A2(n2758), .ZN(n2747) );
  XNOR2_X1 U32580 ( .A(n4789), .B(REG2_REG_15__SCAN_IN), .ZN(n4782) );
  INV_X1 U32590 ( .A(n2750), .ZN(n2749) );
  NAND2_X1 U32600 ( .A1(n2752), .A2(IR_REG_31__SCAN_IN), .ZN(n2748) );
  XNOR2_X1 U32610 ( .A(n2748), .B(n3179), .ZN(n5105) );
  NAND2_X1 U32620 ( .A1(n2749), .A2(n5105), .ZN(n2751) );
  INV_X1 U32630 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4553) );
  NAND2_X1 U32640 ( .A1(n2751), .A2(n4336), .ZN(n4348) );
  XNOR2_X1 U32650 ( .A(n2844), .B(IR_REG_17__SCAN_IN), .ZN(n4627) );
  XNOR2_X1 U32660 ( .A(n4627), .B(REG2_REG_17__SCAN_IN), .ZN(n4347) );
  NAND2_X1 U32670 ( .A1(n2844), .A2(n3376), .ZN(n2754) );
  NAND2_X1 U32680 ( .A1(n2754), .A2(IR_REG_31__SCAN_IN), .ZN(n2755) );
  NAND2_X1 U32690 ( .A1(REG2_REG_18__SCAN_IN), .A2(n5154), .ZN(n2756) );
  OAI21_X1 U32700 ( .B1(n5154), .B2(REG2_REG_18__SCAN_IN), .A(n2756), .ZN(
        n2792) );
  OR2_X1 U32710 ( .A1(n2506), .A2(n2765), .ZN(n2766) );
  INV_X1 U32720 ( .A(n2849), .ZN(n4623) );
  INV_X1 U32730 ( .A(n2771), .ZN(n2772) );
  NAND2_X1 U32740 ( .A1(n2772), .A2(IR_REG_23__SCAN_IN), .ZN(n2774) );
  INV_X1 U32750 ( .A(n2910), .ZN(n2901) );
  INV_X1 U32760 ( .A(n2913), .ZN(n2775) );
  NAND2_X1 U32770 ( .A1(n2775), .A2(STATE_REG_SCAN_IN), .ZN(n4309) );
  NAND2_X1 U32780 ( .A1(n2901), .A2(n4309), .ZN(n2795) );
  NAND2_X1 U32790 ( .A1(n3192), .A2(n3391), .ZN(n2860) );
  NAND2_X1 U32800 ( .A1(n2860), .A2(IR_REG_31__SCAN_IN), .ZN(n2778) );
  NAND2_X1 U32810 ( .A1(n2779), .A2(n2778), .ZN(n2780) );
  NAND2_X1 U32820 ( .A1(n2782), .A2(n2781), .ZN(n2783) );
  NAND2_X1 U32830 ( .A1(n2783), .A2(IR_REG_31__SCAN_IN), .ZN(n2784) );
  MUX2_X1 U32840 ( .A(IR_REG_31__SCAN_IN), .B(n2784), .S(IR_REG_22__SCAN_IN), 
        .Z(n2786) );
  NAND2_X1 U32850 ( .A1(n2786), .A2(n2785), .ZN(n2954) );
  NAND2_X1 U32860 ( .A1(n2767), .A2(IR_REG_31__SCAN_IN), .ZN(n2787) );
  NAND2_X1 U32870 ( .A1(n2922), .A2(n2913), .ZN(n2788) );
  NAND2_X1 U32880 ( .A1(n4199), .A2(n2788), .ZN(n2794) );
  INV_X1 U32890 ( .A(n2794), .ZN(n2789) );
  NAND2_X1 U32900 ( .A1(n2795), .A2(n2789), .ZN(n2831) );
  INV_X1 U32910 ( .A(n2831), .ZN(n4660) );
  NOR2_X1 U32920 ( .A1(n4805), .A2(n4657), .ZN(n4305) );
  AOI211_X1 U32930 ( .C1(n2503), .C2(n2792), .A(n4798), .B(n3875), .ZN(n2793)
         );
  INV_X1 U32940 ( .A(n2793), .ZN(n2799) );
  INV_X1 U32950 ( .A(n4657), .ZN(n4808) );
  AOI22_X1 U32960 ( .A1(REG3_REG_18__SCAN_IN), .A2(U3149), .B1(n4815), .B2(
        ADDR_REG_18__SCAN_IN), .ZN(n2796) );
  INV_X1 U32970 ( .A(n2796), .ZN(n2797) );
  AOI21_X1 U32980 ( .B1(n5154), .B2(n4804), .A(n2797), .ZN(n2798) );
  NAND2_X1 U32990 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(
        n4670) );
  INV_X1 U33000 ( .A(n4670), .ZN(n2800) );
  NAND2_X1 U33010 ( .A1(n4666), .A2(n2800), .ZN(n4667) );
  NAND2_X1 U33020 ( .A1(n4673), .A2(REG1_REG_1__SCAN_IN), .ZN(n2801) );
  NAND2_X1 U33030 ( .A1(n4858), .A2(REG1_REG_2__SCAN_IN), .ZN(n2802) );
  OAI21_X1 U33040 ( .B1(n4858), .B2(REG1_REG_2__SCAN_IN), .A(n2802), .ZN(n4795) );
  INV_X1 U33050 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4898) );
  NOR2_X1 U33060 ( .A1(n2806), .A2(n4892), .ZN(n2807) );
  NAND2_X1 U33070 ( .A1(n4901), .A2(REG1_REG_5__SCAN_IN), .ZN(n2808) );
  OAI21_X1 U33080 ( .B1(n4901), .B2(REG1_REG_5__SCAN_IN), .A(n2808), .ZN(n4689) );
  NOR2_X1 U33090 ( .A1(n2810), .A2(n4706), .ZN(n2811) );
  INV_X1 U33100 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4929) );
  NAND2_X1 U33110 ( .A1(n4932), .A2(REG1_REG_7__SCAN_IN), .ZN(n2812) );
  OAI21_X1 U33120 ( .B1(n4932), .B2(REG1_REG_7__SCAN_IN), .A(n2812), .ZN(n4712) );
  AOI21_X1 U33130 ( .B1(REG1_REG_7__SCAN_IN), .B2(n4932), .A(n4711), .ZN(n2813) );
  INV_X1 U33140 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4959) );
  XNOR2_X1 U33150 ( .A(n4942), .B(n2813), .ZN(n2854) );
  XOR2_X1 U33160 ( .A(REG1_REG_9__SCAN_IN), .B(n3572), .Z(n4721) );
  INV_X1 U33170 ( .A(n2814), .ZN(n2815) );
  XOR2_X1 U33180 ( .A(n4737), .B(n2814), .Z(n4734) );
  INV_X1 U33190 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4992) );
  NOR2_X1 U33200 ( .A1(n4734), .A2(n4992), .ZN(n4733) );
  NAND2_X1 U33210 ( .A1(n4995), .A2(REG1_REG_11__SCAN_IN), .ZN(n2816) );
  OAI21_X1 U33220 ( .B1(n4995), .B2(REG1_REG_11__SCAN_IN), .A(n2816), .ZN(
        n4744) );
  NOR2_X1 U33230 ( .A1(n4745), .A2(n4744), .ZN(n4743) );
  INV_X1 U33240 ( .A(REG1_REG_12__SCAN_IN), .ZN(n5031) );
  NOR2_X1 U33250 ( .A1(n2819), .A2(n2818), .ZN(n2820) );
  NAND2_X1 U33260 ( .A1(n5034), .A2(REG1_REG_13__SCAN_IN), .ZN(n2821) );
  OAI21_X1 U33270 ( .B1(n5034), .B2(REG1_REG_13__SCAN_IN), .A(n2821), .ZN(
        n4764) );
  XNOR2_X1 U33280 ( .A(n2823), .B(n5052), .ZN(n4770) );
  INV_X1 U33290 ( .A(REG1_REG_14__SCAN_IN), .ZN(n5067) );
  NOR2_X1 U33300 ( .A1(n4770), .A2(n5067), .ZN(n4769) );
  NOR2_X1 U33310 ( .A1(n2823), .A2(n5052), .ZN(n2824) );
  NOR2_X1 U33320 ( .A1(n4769), .A2(n2824), .ZN(n4786) );
  XNOR2_X1 U33330 ( .A(n4789), .B(REG1_REG_15__SCAN_IN), .ZN(n4785) );
  NAND2_X1 U33340 ( .A1(n4789), .A2(REG1_REG_15__SCAN_IN), .ZN(n2825) );
  INV_X1 U33350 ( .A(REG1_REG_16__SCAN_IN), .ZN(n5118) );
  INV_X1 U33360 ( .A(n2826), .ZN(n2827) );
  NAND2_X1 U33370 ( .A1(n2827), .A2(n5105), .ZN(n2828) );
  XNOR2_X1 U33380 ( .A(n4627), .B(REG1_REG_17__SCAN_IN), .ZN(n4343) );
  NAND2_X1 U33390 ( .A1(REG1_REG_18__SCAN_IN), .A2(n5154), .ZN(n2830) );
  OAI21_X1 U33400 ( .B1(n5154), .B2(REG1_REG_18__SCAN_IN), .A(n2830), .ZN(
        n2832) );
  INV_X1 U33410 ( .A(n3871), .ZN(n2835) );
  INV_X1 U33420 ( .A(n4805), .ZN(n4658) );
  AOI21_X1 U33430 ( .B1(n2833), .B2(n2832), .A(n4793), .ZN(n2834) );
  NAND2_X1 U33440 ( .A1(n2835), .A2(n2834), .ZN(n2836) );
  NAND2_X1 U33450 ( .A1(n2679), .A2(n2836), .ZN(U3258) );
  NOR2_X2 U33460 ( .A1(n2876), .A2(n2837), .ZN(U4043) );
  INV_X1 U33470 ( .A(DATAI_28_), .ZN(n2838) );
  MUX2_X1 U33480 ( .A(n2838), .B(n4657), .S(STATE_REG_SCAN_IN), .Z(n2839) );
  INV_X1 U33490 ( .A(n2839), .ZN(U3324) );
  INV_X1 U33500 ( .A(DATAI_27_), .ZN(n2840) );
  MUX2_X1 U33510 ( .A(n2840), .B(n4805), .S(STATE_REG_SCAN_IN), .Z(n2841) );
  INV_X1 U33520 ( .A(n2841), .ZN(U3325) );
  INV_X1 U3353 ( .A(DATAI_20_), .ZN(n3275) );
  NAND2_X1 U33540 ( .A1(n2842), .A2(IR_REG_31__SCAN_IN), .ZN(n2843) );
  NAND2_X1 U3355 ( .A1(n2844), .A2(n2843), .ZN(n2903) );
  MUX2_X1 U3356 ( .A(n3275), .B(n2874), .S(STATE_REG_SCAN_IN), .Z(n2846) );
  INV_X1 U3357 ( .A(n2846), .ZN(U3332) );
  NAND2_X1 U3358 ( .A1(n2895), .A2(n2849), .ZN(n2847) );
  MUX2_X1 U3359 ( .A(n2849), .B(n2847), .S(B_REG_SCAN_IN), .Z(n2848) );
  INV_X1 U3360 ( .A(D_REG_0__SCAN_IN), .ZN(n3399) );
  INV_X1 U3361 ( .A(n4622), .ZN(n2896) );
  AOI22_X1 U3362 ( .A1(n4652), .A2(n3399), .B1(n2884), .B2(n4628), .ZN(U3458)
         );
  NOR2_X1 U3363 ( .A1(n4815), .A2(n4328), .ZN(U3148) );
  AOI21_X1 U3364 ( .B1(n2852), .B2(n2851), .A(n2850), .ZN(n2858) );
  AOI211_X1 U3365 ( .C1(n2854), .C2(n4959), .A(n2853), .B(n4793), .ZN(n2857)
         );
  NOR2_X1 U3366 ( .A1(STATE_REG_SCAN_IN), .A2(n3512), .ZN(n4947) );
  AOI21_X1 U3367 ( .B1(n4815), .B2(ADDR_REG_8__SCAN_IN), .A(n4947), .ZN(n2855)
         );
  OAI21_X1 U3368 ( .B1(n4942), .B2(n4827), .A(n2855), .ZN(n2856) );
  AOI211_X1 U3369 ( .C1(n2858), .C2(n4824), .A(n2857), .B(n2856), .ZN(n2859)
         );
  INV_X1 U3370 ( .A(n2859), .ZN(U3248) );
  INV_X1 U3371 ( .A(n2876), .ZN(n2881) );
  INV_X1 U3372 ( .A(n2866), .ZN(n2863) );
  NAND2_X1 U3373 ( .A1(n2863), .A2(n2862), .ZN(n2865) );
  XNOR2_X2 U3374 ( .A(n2864), .B(IR_REG_30__SCAN_IN), .ZN(n4620) );
  NAND2_X1 U3375 ( .A1(n2866), .A2(IR_REG_31__SCAN_IN), .ZN(n2867) );
  MUX2_X1 U3376 ( .A(IR_REG_31__SCAN_IN), .B(n2867), .S(IR_REG_29__SCAN_IN), 
        .Z(n2868) );
  INV_X1 U3377 ( .A(n2869), .ZN(n4621) );
  NAND2_X1 U3378 ( .A1(n2939), .A2(REG0_REG_0__SCAN_IN), .ZN(n2873) );
  INV_X2 U3379 ( .A(n3785), .ZN(n2982) );
  NAND2_X1 U3380 ( .A1(n2487), .A2(REG3_REG_0__SCAN_IN), .ZN(n2872) );
  NAND2_X1 U3381 ( .A1(n2983), .A2(REG1_REG_0__SCAN_IN), .ZN(n2871) );
  NAND2_X1 U3382 ( .A1(n2485), .A2(REG2_REG_0__SCAN_IN), .ZN(n2870) );
  INV_X1 U3383 ( .A(n2951), .ZN(n2879) );
  AND2_X4 U3384 ( .A1(n2875), .A2(n2876), .ZN(n3468) );
  OAI22_X1 U3385 ( .A1(n2879), .A2(n4015), .B1(n2880), .B2(n4833), .ZN(n2931)
         );
  AOI21_X1 U3386 ( .B1(REG1_REG_0__SCAN_IN), .B2(n2881), .A(n2931), .ZN(n2933)
         );
  INV_X1 U3387 ( .A(n2880), .ZN(n3469) );
  XNOR2_X1 U3388 ( .A(n2933), .B(n2932), .ZN(n4806) );
  NOR4_X1 U3389 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_23__SCAN_IN), .ZN(n2888) );
  NOR4_X1 U3390 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2887) );
  NOR4_X1 U3391 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2886) );
  NOR4_X1 U3392 ( .A1(D_REG_24__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2885) );
  NAND4_X1 U3393 ( .A1(n2888), .A2(n2887), .A3(n2886), .A4(n2885), .ZN(n2963)
         );
  INV_X1 U3394 ( .A(n2963), .ZN(n2894) );
  NOR2_X1 U3395 ( .A1(D_REG_3__SCAN_IN), .A2(D_REG_10__SCAN_IN), .ZN(n2892) );
  NOR4_X1 U3396 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_27__SCAN_IN), .ZN(n2891) );
  NOR4_X1 U3397 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2890) );
  NOR4_X1 U3398 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2889) );
  NAND4_X1 U3399 ( .A1(n2892), .A2(n2891), .A3(n2890), .A4(n2889), .ZN(n2962)
         );
  INV_X1 U3400 ( .A(n2962), .ZN(n2893) );
  NAND3_X1 U3401 ( .A1(n2894), .A2(n2893), .A3(D_REG_1__SCAN_IN), .ZN(n2898)
         );
  NAND2_X1 U3402 ( .A1(n2896), .A2(n2895), .ZN(n4618) );
  INV_X1 U3403 ( .A(n4618), .ZN(n2897) );
  AOI21_X1 U3404 ( .B1(n2899), .B2(n2898), .A(n2897), .ZN(n2900) );
  NAND2_X1 U3405 ( .A1(n4570), .A2(n2900), .ZN(n2917) );
  INV_X1 U3406 ( .A(n2902), .ZN(n2905) );
  NAND2_X1 U3407 ( .A1(n2903), .A2(IR_REG_19__SCAN_IN), .ZN(n2904) );
  OAI211_X1 U3408 ( .C1(n4840), .C2(n4832), .A(n5237), .B(n2955), .ZN(n2915)
         );
  INV_X1 U3409 ( .A(n2915), .ZN(n2907) );
  NAND2_X1 U3410 ( .A1(n2908), .A2(n5229), .ZN(n2911) );
  NAND2_X1 U3411 ( .A1(n2874), .A2(n4840), .ZN(n2912) );
  NAND2_X1 U3412 ( .A1(n2912), .A2(n2922), .ZN(n2919) );
  NOR2_X1 U3413 ( .A1(n2955), .A2(U3149), .ZN(n2914) );
  NAND2_X1 U3414 ( .A1(n2964), .A2(n2914), .ZN(n4304) );
  NAND3_X1 U3415 ( .A1(n4304), .A2(n5237), .A3(n2915), .ZN(n2916) );
  NAND2_X1 U3416 ( .A1(n2917), .A2(n2916), .ZN(n2918) );
  NAND2_X1 U3417 ( .A1(n2918), .A2(n2964), .ZN(n3520) );
  OR2_X1 U3418 ( .A1(n3520), .A2(U3149), .ZN(n4136) );
  AOI22_X1 U3419 ( .A1(n5160), .A2(n2950), .B1(REG3_REG_0__SCAN_IN), .B2(n4136), .ZN(n2928) );
  INV_X1 U3420 ( .A(n2919), .ZN(n2920) );
  NAND2_X1 U3421 ( .A1(n2939), .A2(REG0_REG_1__SCAN_IN), .ZN(n2926) );
  NAND2_X1 U3422 ( .A1(n2487), .A2(REG3_REG_1__SCAN_IN), .ZN(n2925) );
  NAND2_X1 U3423 ( .A1(n2484), .A2(REG2_REG_1__SCAN_IN), .ZN(n2924) );
  NAND2_X1 U3424 ( .A1(n2983), .A2(REG1_REG_1__SCAN_IN), .ZN(n2923) );
  NAND4_X2 U3425 ( .A1(n2926), .A2(n2925), .A3(n2924), .A4(n2923), .ZN(n2949)
         );
  NAND2_X1 U3426 ( .A1(n4148), .A2(n2949), .ZN(n2927) );
  OAI211_X1 U3427 ( .C1(n4806), .C2(n5186), .A(n2928), .B(n2927), .ZN(U3229)
         );
  NAND2_X1 U3428 ( .A1(n4840), .A2(n4624), .ZN(n2930) );
  INV_X1 U3429 ( .A(DATAI_1_), .ZN(n3306) );
  OR2_X1 U3430 ( .A1(n4258), .A2(n2486), .ZN(n2934) );
  NAND2_X1 U3431 ( .A1(n2935), .A2(n2934), .ZN(n2936) );
  XNOR2_X1 U3432 ( .A(n2936), .B(n4016), .ZN(n3464) );
  INV_X1 U3433 ( .A(n2949), .ZN(n4835) );
  XNOR2_X1 U3434 ( .A(n3464), .B(n2938), .ZN(n3467) );
  XNOR2_X1 U3435 ( .A(n3466), .B(n3467), .ZN(n2946) );
  INV_X1 U3436 ( .A(n4258), .ZN(n2997) );
  AOI22_X1 U3437 ( .A1(n5160), .A2(n2997), .B1(REG3_REG_1__SCAN_IN), .B2(n4136), .ZN(n2945) );
  NAND2_X1 U3438 ( .A1(n5190), .A2(n4511), .ZN(n4026) );
  AND2_X1 U3439 ( .A1(n2484), .A2(REG2_REG_2__SCAN_IN), .ZN(n2940) );
  NAND2_X1 U3440 ( .A1(n2487), .A2(REG3_REG_2__SCAN_IN), .ZN(n2942) );
  NAND2_X1 U3441 ( .A1(n2983), .A2(REG1_REG_2__SCAN_IN), .ZN(n2941) );
  AOI22_X1 U3442 ( .A1(n4151), .A2(n2951), .B1(n4148), .B2(n2978), .ZN(n2944)
         );
  OAI211_X1 U3443 ( .C1(n2946), .C2(n5186), .A(n2945), .B(n2944), .ZN(U3219)
         );
  OR2_X1 U3444 ( .A1(n2874), .A2(n4243), .ZN(n2948) );
  NAND2_X1 U3445 ( .A1(n4626), .A2(n4624), .ZN(n2947) );
  INV_X1 U3446 ( .A(n2996), .ZN(n4239) );
  XNOR2_X1 U3447 ( .A(n4239), .B(n4260), .ZN(n2961) );
  NAND2_X1 U3448 ( .A1(n2952), .A2(n2996), .ZN(n2976) );
  OAI21_X1 U3449 ( .B1(n2996), .B2(n2952), .A(n2976), .ZN(n2953) );
  INV_X1 U3450 ( .A(n2953), .ZN(n4854) );
  NAND2_X1 U3451 ( .A1(n2929), .A2(n2954), .ZN(n2957) );
  AND2_X1 U3452 ( .A1(n2955), .A2(n4840), .ZN(n2956) );
  NAND2_X1 U3453 ( .A1(n2957), .A2(n2956), .ZN(n4561) );
  INV_X1 U3454 ( .A(n4561), .ZN(n4875) );
  NAND2_X1 U3455 ( .A1(n4854), .A2(n4875), .ZN(n2959) );
  AOI22_X1 U3456 ( .A1(n4511), .A2(n2951), .B1(n2978), .B2(n5177), .ZN(n2958)
         );
  OAI211_X1 U3457 ( .C1(n5237), .C2(n4258), .A(n2959), .B(n2958), .ZN(n2960)
         );
  AOI21_X1 U34580 ( .B1(n5207), .B2(n2961), .A(n2960), .ZN(n4851) );
  NOR2_X1 U34590 ( .A1(n2963), .A2(n2962), .ZN(n2965) );
  OAI21_X1 U3460 ( .B1(n2966), .B2(D_REG_1__SCAN_IN), .A(n4618), .ZN(n4567) );
  NOR2_X1 U3461 ( .A1(n4568), .A2(n4567), .ZN(n2967) );
  NAND2_X1 U3462 ( .A1(n4606), .A2(n2967), .ZN(n2969) );
  OR2_X1 U3463 ( .A1(n2929), .A2(n4840), .ZN(n3048) );
  INV_X1 U3464 ( .A(n3048), .ZN(n4847) );
  NAND2_X1 U3465 ( .A1(n4558), .A2(n4847), .ZN(n3034) );
  INV_X1 U3466 ( .A(n3034), .ZN(n4886) );
  INV_X1 U34670 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2972) );
  NOR2_X1 U3468 ( .A1(n4833), .A2(n4258), .ZN(n4850) );
  OR2_X1 U34690 ( .A1(n5219), .A2(n4626), .ZN(n2968) );
  NOR3_X1 U3470 ( .A1(n4850), .A2(n5196), .A3(n3012), .ZN(n2970) );
  AOI21_X1 U34710 ( .B1(n5136), .B2(REG3_REG_1__SCAN_IN), .A(n2970), .ZN(n2971) );
  OAI21_X1 U3472 ( .B1(n2972), .B2(n4558), .A(n2971), .ZN(n2973) );
  AOI21_X1 U34730 ( .B1(n4886), .B2(n4854), .A(n2973), .ZN(n2974) );
  OAI21_X1 U3474 ( .B1(n4851), .B2(n5246), .A(n2974), .ZN(U3289) );
  NAND2_X1 U34750 ( .A1(n2949), .A2(n2997), .ZN(n2975) );
  MUX2_X1 U3476 ( .A(n4858), .B(DATAI_2_), .S(n2977), .Z(n4137) );
  NAND2_X1 U34770 ( .A1(n2979), .A2(n4137), .ZN(n3000) );
  NAND2_X1 U3478 ( .A1(n2978), .A2(n3029), .ZN(n4264) );
  NAND2_X1 U34790 ( .A1(n3000), .A2(n4264), .ZN(n2999) );
  NAND2_X1 U3480 ( .A1(n2979), .A2(n3029), .ZN(n2980) );
  NAND2_X1 U34810 ( .A1(n2485), .A2(REG2_REG_3__SCAN_IN), .ZN(n2987) );
  INV_X1 U3482 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4884) );
  NAND2_X1 U34830 ( .A1(n2982), .A2(n4884), .ZN(n2986) );
  NAND2_X1 U3484 ( .A1(n2939), .A2(REG0_REG_3__SCAN_IN), .ZN(n2985) );
  NAND2_X1 U34850 ( .A1(n2483), .A2(REG1_REG_3__SCAN_IN), .ZN(n2984) );
  MUX2_X1 U3486 ( .A(n4685), .B(DATAI_3_), .S(n2482), .Z(n4879) );
  NOR2_X1 U34870 ( .A1(n4332), .A2(n4879), .ZN(n2988) );
  OAI22_X1 U3488 ( .A1(n4868), .A2(n2988), .B1(n3477), .B2(n3013), .ZN(n3046)
         );
  NAND2_X1 U34890 ( .A1(n2485), .A2(REG2_REG_4__SCAN_IN), .ZN(n2993) );
  NOR2_X1 U3490 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2989) );
  NOR2_X1 U34910 ( .A1(n3003), .A2(n2989), .ZN(n4107) );
  NAND2_X1 U3492 ( .A1(n2982), .A2(n4107), .ZN(n2992) );
  NAND2_X1 U34930 ( .A1(n2939), .A2(REG0_REG_4__SCAN_IN), .ZN(n2991) );
  NAND2_X1 U3494 ( .A1(n4188), .A2(REG1_REG_4__SCAN_IN), .ZN(n2990) );
  INV_X1 U34950 ( .A(n4331), .ZN(n3485) );
  INV_X1 U3496 ( .A(n4892), .ZN(n2994) );
  MUX2_X1 U34970 ( .A(n2994), .B(DATAI_4_), .S(n2977), .Z(n4108) );
  NAND2_X1 U3498 ( .A1(n3485), .A2(n4108), .ZN(n4267) );
  NAND2_X1 U34990 ( .A1(n4331), .A2(n2544), .ZN(n4269) );
  NAND2_X1 U3500 ( .A1(n4267), .A2(n4269), .ZN(n4233) );
  XNOR2_X1 U35010 ( .A(n3046), .B(n4233), .ZN(n4893) );
  INV_X1 U3502 ( .A(n4260), .ZN(n2995) );
  OR2_X1 U35030 ( .A1(n2996), .A2(n2995), .ZN(n2998) );
  NAND2_X1 U3504 ( .A1(n4835), .A2(n2997), .ZN(n4261) );
  NAND2_X1 U35050 ( .A1(n2998), .A2(n4261), .ZN(n3023) );
  INV_X1 U35060 ( .A(n2999), .ZN(n3019) );
  NAND2_X1 U35070 ( .A1(n3023), .A2(n3019), .ZN(n3001) );
  NAND2_X1 U35080 ( .A1(n3001), .A2(n3000), .ZN(n4869) );
  NAND2_X1 U35090 ( .A1(n3477), .A2(n4879), .ZN(n4266) );
  NAND2_X1 U35100 ( .A1(n4332), .A2(n3013), .ZN(n4263) );
  AND2_X1 U35110 ( .A1(n4266), .A2(n4263), .ZN(n4219) );
  NAND2_X1 U35120 ( .A1(n4869), .A2(n4219), .ZN(n3002) );
  NAND2_X1 U35130 ( .A1(n3002), .A2(n4266), .ZN(n3037) );
  XOR2_X1 U35140 ( .A(n3037), .B(n4233), .Z(n3010) );
  NAND2_X1 U35150 ( .A1(n3003), .A2(REG3_REG_5__SCAN_IN), .ZN(n3041) );
  OAI21_X1 U35160 ( .B1(n3003), .B2(REG3_REG_5__SCAN_IN), .A(n3041), .ZN(n4915) );
  INV_X1 U35170 ( .A(n4915), .ZN(n3053) );
  NAND2_X1 U35180 ( .A1(n2982), .A2(n3053), .ZN(n3007) );
  NAND2_X1 U35190 ( .A1(n2485), .A2(REG2_REG_5__SCAN_IN), .ZN(n3006) );
  NAND2_X1 U35200 ( .A1(n2483), .A2(REG1_REG_5__SCAN_IN), .ZN(n3005) );
  NAND2_X1 U35210 ( .A1(n3858), .A2(REG0_REG_5__SCAN_IN), .ZN(n3004) );
  NAND4_X1 U35220 ( .A1(n3007), .A2(n3006), .A3(n3005), .A4(n3004), .ZN(n4330)
         );
  AOI22_X1 U35230 ( .A1(n4511), .A2(n4332), .B1(n4330), .B2(n5177), .ZN(n3008)
         );
  OAI21_X1 U35240 ( .B1(n2544), .B2(n5237), .A(n3008), .ZN(n3009) );
  AOI21_X1 U35250 ( .B1(n3010), .B2(n5207), .A(n3009), .ZN(n3011) );
  OAI21_X1 U35260 ( .B1(n4893), .B2(n4561), .A(n3011), .ZN(n4894) );
  NAND2_X1 U35270 ( .A1(n4894), .A2(n4558), .ZN(n3018) );
  AOI21_X1 U35280 ( .B1(n4876), .B2(n4108), .A(n5219), .ZN(n3014) );
  AND2_X1 U35290 ( .A1(n3014), .A2(n3049), .ZN(n4895) );
  NOR2_X1 U35300 ( .A1(n5246), .A2(n4626), .ZN(n4524) );
  INV_X1 U35310 ( .A(n4107), .ZN(n3015) );
  OAI22_X1 U35320 ( .A1(n4558), .A2(n4821), .B1(n3015), .B2(n5216), .ZN(n3016)
         );
  AOI21_X1 U35330 ( .B1(n4895), .B2(n4524), .A(n3016), .ZN(n3017) );
  OAI211_X1 U35340 ( .C1(n4893), .C2(n3034), .A(n3018), .B(n3017), .ZN(U3286)
         );
  INV_X1 U35350 ( .A(n3020), .ZN(n3021) );
  AOI21_X1 U35360 ( .B1(n3019), .B2(n3022), .A(n3021), .ZN(n4862) );
  XNOR2_X1 U35370 ( .A(n3023), .B(n2999), .ZN(n3028) );
  INV_X1 U35380 ( .A(n4862), .ZN(n3026) );
  AOI22_X1 U35390 ( .A1(n4511), .A2(n2949), .B1(n4332), .B2(n5177), .ZN(n3024)
         );
  OAI21_X1 U35400 ( .B1(n3029), .B2(n5237), .A(n3024), .ZN(n3025) );
  AOI21_X1 U35410 ( .B1(n3026), .B2(n4875), .A(n3025), .ZN(n3027) );
  OAI21_X1 U35420 ( .B1(n5091), .B2(n3028), .A(n3027), .ZN(n4863) );
  NAND2_X1 U35430 ( .A1(n4863), .A2(n4558), .ZN(n3033) );
  OAI21_X1 U35440 ( .B1(n3012), .B2(n3029), .A(n4878), .ZN(n4860) );
  INV_X1 U35450 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3030) );
  OAI22_X1 U35460 ( .A1(n4860), .A2(n5196), .B1(n3030), .B2(n5216), .ZN(n3031)
         );
  AOI21_X1 U35470 ( .B1(REG2_REG_2__SCAN_IN), .B2(n5246), .A(n3031), .ZN(n3032) );
  OAI211_X1 U35480 ( .C1(n4862), .C2(n3034), .A(n3033), .B(n3032), .ZN(U3288)
         );
  MUX2_X1 U35490 ( .A(n4901), .B(DATAI_5_), .S(n2482), .Z(n4913) );
  INV_X1 U35500 ( .A(n4913), .ZN(n3051) );
  INV_X1 U35510 ( .A(n4330), .ZN(n3035) );
  NAND2_X1 U35520 ( .A1(n3035), .A2(n4913), .ZN(n4249) );
  NAND2_X1 U35530 ( .A1(n4330), .A2(n3051), .ZN(n3527) );
  NAND2_X1 U35540 ( .A1(n4249), .A2(n3527), .ZN(n4232) );
  INV_X1 U35550 ( .A(n4232), .ZN(n3039) );
  INV_X1 U35560 ( .A(n4267), .ZN(n3036) );
  OAI21_X1 U35570 ( .B1(n3037), .B2(n3036), .A(n4269), .ZN(n3038) );
  NAND2_X1 U35580 ( .A1(n3038), .A2(n3039), .ZN(n3529) );
  OAI211_X1 U35590 ( .C1(n3039), .C2(n3038), .A(n3529), .B(n5207), .ZN(n3045)
         );
  AOI22_X1 U35600 ( .A1(n2485), .A2(REG2_REG_6__SCAN_IN), .B1(n4188), .B2(
        REG1_REG_6__SCAN_IN), .ZN(n3044) );
  AND2_X1 U35610 ( .A1(n3041), .A2(n3040), .ZN(n3042) );
  NOR2_X1 U35620 ( .A1(n3059), .A2(n3042), .ZN(n4147) );
  AOI22_X1 U35630 ( .A1(n2982), .A2(n4147), .B1(n3858), .B2(
        REG0_REG_6__SCAN_IN), .ZN(n3043) );
  AOI22_X1 U35640 ( .A1(n4329), .A2(n5177), .B1(n4511), .B2(n4331), .ZN(n4906)
         );
  OAI211_X1 U35650 ( .C1(n5237), .C2(n3051), .A(n3045), .B(n4906), .ZN(n4917)
         );
  INV_X1 U35660 ( .A(n4917), .ZN(n3057) );
  AOI21_X1 U35670 ( .B1(n3046), .B2(n4233), .A(n2681), .ZN(n3047) );
  OAI21_X1 U35680 ( .B1(n3047), .B2(n4232), .A(n3069), .ZN(n4919) );
  NAND2_X1 U35690 ( .A1(n4561), .A2(n3048), .ZN(n4981) );
  INV_X1 U35700 ( .A(n3049), .ZN(n3052) );
  INV_X1 U35710 ( .A(n3070), .ZN(n3050) );
  OAI21_X1 U35720 ( .B1(n3052), .B2(n3051), .A(n3050), .ZN(n4916) );
  AOI22_X1 U35730 ( .A1(n5246), .A2(REG2_REG_5__SCAN_IN), .B1(n3053), .B2(
        n5136), .ZN(n3054) );
  OAI21_X1 U35740 ( .B1(n4916), .B2(n5196), .A(n3054), .ZN(n3055) );
  AOI21_X1 U35750 ( .B1(n4919), .B2(n5144), .A(n3055), .ZN(n3056) );
  OAI21_X1 U35760 ( .B1(n5246), .B2(n3057), .A(n3056), .ZN(U3285) );
  NAND2_X1 U35770 ( .A1(n3529), .A2(n3527), .ZN(n3058) );
  MUX2_X1 U35780 ( .A(n4923), .B(DATAI_6_), .S(n2482), .Z(n3540) );
  NAND2_X1 U35790 ( .A1(n3541), .A2(n3540), .ZN(n4272) );
  NAND2_X1 U35800 ( .A1(n4329), .A2(n4149), .ZN(n4247) );
  NAND2_X1 U35810 ( .A1(n4272), .A2(n4247), .ZN(n4225) );
  XNOR2_X1 U3582 ( .A(n3058), .B(n4225), .ZN(n3067) );
  NAND2_X1 U3583 ( .A1(n2485), .A2(REG2_REG_7__SCAN_IN), .ZN(n3064) );
  NAND2_X1 U3584 ( .A1(n3059), .A2(REG3_REG_7__SCAN_IN), .ZN(n3513) );
  OR2_X1 U3585 ( .A1(n3059), .A2(REG3_REG_7__SCAN_IN), .ZN(n3060) );
  AND2_X1 U3586 ( .A1(n3513), .A2(n3060), .ZN(n3537) );
  NAND2_X1 U3587 ( .A1(n2982), .A2(n3537), .ZN(n3063) );
  NAND2_X1 U3588 ( .A1(n3858), .A2(REG0_REG_7__SCAN_IN), .ZN(n3062) );
  NAND2_X1 U3589 ( .A1(n4188), .A2(REG1_REG_7__SCAN_IN), .ZN(n3061) );
  NAND4_X1 U3590 ( .A1(n3064), .A2(n3063), .A3(n3062), .A4(n3061), .ZN(n4327)
         );
  AOI22_X1 U3591 ( .A1(n4511), .A2(n4330), .B1(n4327), .B2(n5177), .ZN(n3065)
         );
  OAI21_X1 U3592 ( .B1(n4149), .B2(n5237), .A(n3065), .ZN(n3066) );
  AOI21_X1 U3593 ( .B1(n3067), .B2(n5207), .A(n3066), .ZN(n4925) );
  OR2_X1 U3594 ( .A1(n4330), .A2(n4913), .ZN(n3068) );
  XNOR2_X1 U3595 ( .A(n3544), .B(n4225), .ZN(n4928) );
  NAND2_X1 U3596 ( .A1(n3070), .A2(n4149), .ZN(n3534) );
  OAI21_X1 U3597 ( .B1(n3070), .B2(n4149), .A(n3534), .ZN(n4926) );
  NOR2_X1 U3598 ( .A1(n4926), .A2(n5196), .ZN(n3073) );
  INV_X1 U3599 ( .A(n4147), .ZN(n3071) );
  OAI22_X1 U3600 ( .A1(n4558), .A2(n4701), .B1(n3071), .B2(n5216), .ZN(n3072)
         );
  AOI211_X1 U3601 ( .C1(n4928), .C2(n5144), .A(n3073), .B(n3072), .ZN(n3074)
         );
  OAI21_X1 U3602 ( .B1(n5246), .B2(n4925), .A(n3074), .ZN(U3284) );
  XOR2_X1 U3603 ( .A(DATAI_31_), .B(keyinput_128), .Z(n3078) );
  XOR2_X1 U3604 ( .A(DATAI_29_), .B(keyinput_130), .Z(n3077) );
  XOR2_X1 U3605 ( .A(DATAI_30_), .B(keyinput_129), .Z(n3076) );
  XNOR2_X1 U3606 ( .A(DATAI_28_), .B(keyinput_131), .ZN(n3075) );
  NAND4_X1 U3607 ( .A1(n3078), .A2(n3077), .A3(n3076), .A4(n3075), .ZN(n3081)
         );
  XOR2_X1 U3608 ( .A(DATAI_27_), .B(keyinput_132), .Z(n3080) );
  XOR2_X1 U3609 ( .A(DATAI_26_), .B(keyinput_133), .Z(n3079) );
  AOI21_X1 U3610 ( .B1(n3081), .B2(n3080), .A(n3079), .ZN(n3085) );
  XOR2_X1 U3611 ( .A(DATAI_25_), .B(keyinput_134), .Z(n3084) );
  XOR2_X1 U3612 ( .A(DATAI_23_), .B(keyinput_136), .Z(n3083) );
  XNOR2_X1 U3613 ( .A(DATAI_24_), .B(keyinput_135), .ZN(n3082) );
  OAI211_X1 U3614 ( .C1(n3085), .C2(n3084), .A(n3083), .B(n3082), .ZN(n3087)
         );
  XNOR2_X1 U3615 ( .A(DATAI_22_), .B(keyinput_137), .ZN(n3086) );
  NAND2_X1 U3616 ( .A1(n3087), .A2(n3086), .ZN(n3094) );
  INV_X1 U3617 ( .A(DATAI_21_), .ZN(n3089) );
  OAI22_X1 U3618 ( .A1(n3089), .A2(keyinput_138), .B1(DATAI_20_), .B2(
        keyinput_139), .ZN(n3088) );
  AOI221_X1 U3619 ( .B1(n3089), .B2(keyinput_138), .C1(keyinput_139), .C2(
        DATAI_20_), .A(n3088), .ZN(n3093) );
  XOR2_X1 U3620 ( .A(DATAI_17_), .B(keyinput_142), .Z(n3092) );
  OAI22_X1 U3621 ( .A1(DATAI_19_), .A2(keyinput_140), .B1(DATAI_18_), .B2(
        keyinput_141), .ZN(n3090) );
  AOI221_X1 U3622 ( .B1(DATAI_19_), .B2(keyinput_140), .C1(keyinput_141), .C2(
        DATAI_18_), .A(n3090), .ZN(n3091) );
  NAND4_X1 U3623 ( .A1(n3094), .A2(n3093), .A3(n3092), .A4(n3091), .ZN(n3098)
         );
  INV_X1 U3624 ( .A(DATAI_16_), .ZN(n5104) );
  XNOR2_X1 U3625 ( .A(n5104), .B(keyinput_143), .ZN(n3097) );
  INV_X1 U3626 ( .A(DATAI_14_), .ZN(n5051) );
  XNOR2_X1 U3627 ( .A(n5051), .B(keyinput_145), .ZN(n3096) );
  XOR2_X1 U3628 ( .A(DATAI_15_), .B(keyinput_144), .Z(n3095) );
  AOI211_X1 U3629 ( .C1(n3098), .C2(n3097), .A(n3096), .B(n3095), .ZN(n3101)
         );
  XNOR2_X1 U3630 ( .A(DATAI_13_), .B(keyinput_146), .ZN(n3100) );
  XNOR2_X1 U3631 ( .A(DATAI_12_), .B(keyinput_147), .ZN(n3099) );
  NOR3_X1 U3632 ( .A1(n3101), .A2(n3100), .A3(n3099), .ZN(n3107) );
  INV_X1 U3633 ( .A(DATAI_10_), .ZN(n3291) );
  AOI22_X1 U3634 ( .A1(DATAI_7_), .A2(keyinput_152), .B1(n3291), .B2(
        keyinput_149), .ZN(n3102) );
  OAI221_X1 U3635 ( .B1(DATAI_7_), .B2(keyinput_152), .C1(n3291), .C2(
        keyinput_149), .A(n3102), .ZN(n3106) );
  AOI22_X1 U3636 ( .A1(DATAI_8_), .A2(keyinput_151), .B1(DATAI_9_), .B2(
        keyinput_150), .ZN(n3103) );
  OAI221_X1 U3637 ( .B1(DATAI_8_), .B2(keyinput_151), .C1(DATAI_9_), .C2(
        keyinput_150), .A(n3103), .ZN(n3105) );
  XNOR2_X1 U3638 ( .A(DATAI_11_), .B(keyinput_148), .ZN(n3104) );
  NOR4_X1 U3639 ( .A1(n3107), .A2(n3106), .A3(n3105), .A4(n3104), .ZN(n3110)
         );
  XNOR2_X1 U3640 ( .A(DATAI_6_), .B(keyinput_153), .ZN(n3109) );
  XOR2_X1 U3641 ( .A(DATAI_5_), .B(keyinput_154), .Z(n3108) );
  OAI21_X1 U3642 ( .B1(n3110), .B2(n3109), .A(n3108), .ZN(n3114) );
  XNOR2_X1 U3643 ( .A(DATAI_4_), .B(keyinput_155), .ZN(n3113) );
  XOR2_X1 U3644 ( .A(DATAI_2_), .B(keyinput_157), .Z(n3112) );
  XOR2_X1 U3645 ( .A(DATAI_3_), .B(keyinput_156), .Z(n3111) );
  AOI211_X1 U3646 ( .C1(n3114), .C2(n3113), .A(n3112), .B(n3111), .ZN(n3121)
         );
  XNOR2_X1 U3647 ( .A(n3306), .B(keyinput_158), .ZN(n3120) );
  XOR2_X1 U3648 ( .A(DATAI_0_), .B(keyinput_159), .Z(n3118) );
  XOR2_X1 U3649 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_161), .Z(n3117) );
  XNOR2_X1 U3650 ( .A(U3149), .B(keyinput_160), .ZN(n3116) );
  INV_X1 U3651 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4033) );
  XNOR2_X1 U3652 ( .A(n4033), .B(keyinput_162), .ZN(n3115) );
  NOR4_X1 U3653 ( .A1(n3118), .A2(n3117), .A3(n3116), .A4(n3115), .ZN(n3119)
         );
  OAI21_X1 U3654 ( .B1(n3121), .B2(n3120), .A(n3119), .ZN(n3124) );
  XOR2_X1 U3655 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput_163), .Z(n3123) );
  XNOR2_X1 U3656 ( .A(n3770), .B(keyinput_164), .ZN(n3122) );
  AOI21_X1 U3657 ( .B1(n3124), .B2(n3123), .A(n3122), .ZN(n3129) );
  XOR2_X1 U3658 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput_165), .Z(n3126) );
  XNOR2_X1 U3659 ( .A(n4884), .B(keyinput_166), .ZN(n3125) );
  NAND2_X1 U3660 ( .A1(n3126), .A2(n3125), .ZN(n3128) );
  XNOR2_X1 U3661 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput_167), .ZN(n3127) );
  OAI21_X1 U3662 ( .B1(n3129), .B2(n3128), .A(n3127), .ZN(n3136) );
  INV_X1 U3663 ( .A(REG3_REG_28__SCAN_IN), .ZN(n4022) );
  XNOR2_X1 U3664 ( .A(n4022), .B(keyinput_168), .ZN(n3135) );
  XOR2_X1 U3665 ( .A(REG3_REG_21__SCAN_IN), .B(keyinput_171), .Z(n3133) );
  XOR2_X1 U3666 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_170), .Z(n3132) );
  XNOR2_X1 U3667 ( .A(n3512), .B(keyinput_169), .ZN(n3131) );
  XNOR2_X1 U3668 ( .A(REG3_REG_12__SCAN_IN), .B(keyinput_172), .ZN(n3130) );
  NAND4_X1 U3669 ( .A1(n3133), .A2(n3132), .A3(n3131), .A4(n3130), .ZN(n3134)
         );
  AOI21_X1 U3670 ( .B1(n3136), .B2(n3135), .A(n3134), .ZN(n3140) );
  XOR2_X1 U3671 ( .A(REG3_REG_25__SCAN_IN), .B(keyinput_173), .Z(n3139) );
  XOR2_X1 U3672 ( .A(REG3_REG_5__SCAN_IN), .B(keyinput_175), .Z(n3138) );
  XOR2_X1 U3673 ( .A(REG3_REG_16__SCAN_IN), .B(keyinput_174), .Z(n3137) );
  OAI211_X1 U3674 ( .C1(n3140), .C2(n3139), .A(n3138), .B(n3137), .ZN(n3143)
         );
  XOR2_X1 U3675 ( .A(REG3_REG_17__SCAN_IN), .B(keyinput_176), .Z(n3142) );
  XNOR2_X1 U3676 ( .A(REG3_REG_24__SCAN_IN), .B(keyinput_177), .ZN(n3141) );
  AOI21_X1 U3677 ( .B1(n3143), .B2(n3142), .A(n3141), .ZN(n3146) );
  XNOR2_X1 U3678 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_178), .ZN(n3145) );
  XNOR2_X1 U3679 ( .A(n3595), .B(keyinput_179), .ZN(n3144) );
  OAI21_X1 U3680 ( .B1(n3146), .B2(n3145), .A(n3144), .ZN(n3153) );
  XOR2_X1 U3681 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_180), .Z(n3152) );
  XOR2_X1 U3682 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_183), .Z(n3150) );
  XOR2_X1 U3683 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput_181), .Z(n3149) );
  XNOR2_X1 U3684 ( .A(REG3_REG_13__SCAN_IN), .B(keyinput_182), .ZN(n3148) );
  XNOR2_X1 U3685 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_184), .ZN(n3147) );
  NAND4_X1 U3686 ( .A1(n3150), .A2(n3149), .A3(n3148), .A4(n3147), .ZN(n3151)
         );
  AOI21_X1 U3687 ( .B1(n3153), .B2(n3152), .A(n3151), .ZN(n3165) );
  XNOR2_X1 U3688 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_185), .ZN(n3164) );
  OAI22_X1 U3689 ( .A1(IR_REG_6__SCAN_IN), .A2(keyinput_189), .B1(keyinput_190), .B2(IR_REG_7__SCAN_IN), .ZN(n3154) );
  AOI221_X1 U3690 ( .B1(IR_REG_6__SCAN_IN), .B2(keyinput_189), .C1(
        IR_REG_7__SCAN_IN), .C2(keyinput_190), .A(n3154), .ZN(n3163) );
  XNOR2_X1 U3691 ( .A(n3155), .B(keyinput_186), .ZN(n3158) );
  XNOR2_X1 U3692 ( .A(n3351), .B(keyinput_191), .ZN(n3157) );
  XNOR2_X1 U3693 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_192), .ZN(n3156) );
  NAND3_X1 U3694 ( .A1(n3158), .A2(n3157), .A3(n3156), .ZN(n3161) );
  XNOR2_X1 U3695 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_187), .ZN(n3160) );
  XNOR2_X1 U3696 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_188), .ZN(n3159) );
  NOR3_X1 U3697 ( .A1(n3161), .A2(n3160), .A3(n3159), .ZN(n3162) );
  OAI211_X1 U3698 ( .C1(n3165), .C2(n3164), .A(n3163), .B(n3162), .ZN(n3169)
         );
  XNOR2_X1 U3699 ( .A(n3166), .B(keyinput_194), .ZN(n3168) );
  XNOR2_X1 U3700 ( .A(IR_REG_10__SCAN_IN), .B(keyinput_193), .ZN(n3167) );
  NAND3_X1 U3701 ( .A1(n3169), .A2(n3168), .A3(n3167), .ZN(n3174) );
  XNOR2_X1 U3702 ( .A(n3170), .B(keyinput_195), .ZN(n3173) );
  XOR2_X1 U3703 ( .A(IR_REG_13__SCAN_IN), .B(keyinput_196), .Z(n3172) );
  XNOR2_X1 U3704 ( .A(IR_REG_14__SCAN_IN), .B(keyinput_197), .ZN(n3171) );
  AOI211_X1 U3705 ( .C1(n3174), .C2(n3173), .A(n3172), .B(n3171), .ZN(n3187)
         );
  XNOR2_X1 U3706 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_204), .ZN(n3178) );
  XNOR2_X1 U3707 ( .A(IR_REG_22__SCAN_IN), .B(keyinput_205), .ZN(n3177) );
  XNOR2_X1 U3708 ( .A(IR_REG_17__SCAN_IN), .B(keyinput_200), .ZN(n3176) );
  XNOR2_X1 U3709 ( .A(IR_REG_19__SCAN_IN), .B(keyinput_202), .ZN(n3175) );
  NAND4_X1 U3710 ( .A1(n3178), .A2(n3177), .A3(n3176), .A4(n3175), .ZN(n3186)
         );
  XNOR2_X1 U3711 ( .A(n3179), .B(keyinput_199), .ZN(n3184) );
  XNOR2_X1 U3712 ( .A(n3374), .B(keyinput_203), .ZN(n3183) );
  XNOR2_X1 U3713 ( .A(n3180), .B(keyinput_201), .ZN(n3182) );
  XNOR2_X1 U3714 ( .A(IR_REG_15__SCAN_IN), .B(keyinput_198), .ZN(n3181) );
  NAND4_X1 U3715 ( .A1(n3184), .A2(n3183), .A3(n3182), .A4(n3181), .ZN(n3185)
         );
  NOR3_X1 U3716 ( .A1(n3187), .A2(n3186), .A3(n3185), .ZN(n3191) );
  XNOR2_X1 U3717 ( .A(n3188), .B(keyinput_207), .ZN(n3190) );
  XNOR2_X1 U3718 ( .A(IR_REG_23__SCAN_IN), .B(keyinput_206), .ZN(n3189) );
  NOR3_X1 U3719 ( .A1(n3191), .A2(n3190), .A3(n3189), .ZN(n3195) );
  XNOR2_X1 U3720 ( .A(n3387), .B(keyinput_208), .ZN(n3194) );
  XNOR2_X1 U3721 ( .A(n3192), .B(keyinput_209), .ZN(n3193) );
  OAI21_X1 U3722 ( .B1(n3195), .B2(n3194), .A(n3193), .ZN(n3202) );
  XOR2_X1 U3723 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_214), .Z(n3198) );
  XOR2_X1 U3724 ( .A(IR_REG_30__SCAN_IN), .B(keyinput_213), .Z(n3197) );
  XNOR2_X1 U3725 ( .A(n3391), .B(keyinput_210), .ZN(n3196) );
  NOR3_X1 U3726 ( .A1(n3198), .A2(n3197), .A3(n3196), .ZN(n3201) );
  XNOR2_X1 U3727 ( .A(IR_REG_29__SCAN_IN), .B(keyinput_212), .ZN(n3200) );
  XNOR2_X1 U3728 ( .A(IR_REG_28__SCAN_IN), .B(keyinput_211), .ZN(n3199) );
  NAND4_X1 U3729 ( .A1(n3202), .A2(n3201), .A3(n3200), .A4(n3199), .ZN(n3210)
         );
  XNOR2_X1 U3730 ( .A(D_REG_2__SCAN_IN), .B(keyinput_217), .ZN(n3206) );
  OAI22_X1 U3731 ( .A1(n3399), .A2(keyinput_215), .B1(keyinput_216), .B2(
        D_REG_1__SCAN_IN), .ZN(n3203) );
  AOI21_X1 U3732 ( .B1(n3399), .B2(keyinput_215), .A(n3203), .ZN(n3204) );
  INV_X1 U3733 ( .A(n3204), .ZN(n3205) );
  AOI211_X1 U3734 ( .C1(D_REG_1__SCAN_IN), .C2(keyinput_216), .A(n3206), .B(
        n3205), .ZN(n3209) );
  INV_X1 U3735 ( .A(D_REG_3__SCAN_IN), .ZN(n4630) );
  XNOR2_X1 U3736 ( .A(n4630), .B(keyinput_218), .ZN(n3208) );
  XNOR2_X1 U3737 ( .A(D_REG_4__SCAN_IN), .B(keyinput_219), .ZN(n3207) );
  AOI211_X1 U3738 ( .C1(n3210), .C2(n3209), .A(n3208), .B(n3207), .ZN(n3213)
         );
  INV_X1 U3739 ( .A(D_REG_6__SCAN_IN), .ZN(n4633) );
  XNOR2_X1 U3740 ( .A(n4633), .B(keyinput_221), .ZN(n3212) );
  XNOR2_X1 U3741 ( .A(D_REG_5__SCAN_IN), .B(keyinput_220), .ZN(n3211) );
  NOR3_X1 U3742 ( .A1(n3213), .A2(n3212), .A3(n3211), .ZN(n3216) );
  INV_X1 U3743 ( .A(D_REG_7__SCAN_IN), .ZN(n4634) );
  XNOR2_X1 U3744 ( .A(n4634), .B(keyinput_222), .ZN(n3215) );
  XNOR2_X1 U3745 ( .A(D_REG_8__SCAN_IN), .B(keyinput_223), .ZN(n3214) );
  OAI21_X1 U3746 ( .B1(n3216), .B2(n3215), .A(n3214), .ZN(n3219) );
  INV_X1 U3747 ( .A(D_REG_9__SCAN_IN), .ZN(n4636) );
  XNOR2_X1 U3748 ( .A(n4636), .B(keyinput_224), .ZN(n3218) );
  XNOR2_X1 U3749 ( .A(D_REG_10__SCAN_IN), .B(keyinput_225), .ZN(n3217) );
  NAND3_X1 U3750 ( .A1(n3219), .A2(n3218), .A3(n3217), .ZN(n3223) );
  XOR2_X1 U3751 ( .A(D_REG_13__SCAN_IN), .B(keyinput_228), .Z(n3222) );
  XOR2_X1 U3752 ( .A(D_REG_11__SCAN_IN), .B(keyinput_226), .Z(n3221) );
  XNOR2_X1 U3753 ( .A(D_REG_12__SCAN_IN), .B(keyinput_227), .ZN(n3220) );
  NAND4_X1 U3754 ( .A1(n3223), .A2(n3222), .A3(n3221), .A4(n3220), .ZN(n3226)
         );
  XNOR2_X1 U3755 ( .A(D_REG_14__SCAN_IN), .B(keyinput_229), .ZN(n3225) );
  XNOR2_X1 U3756 ( .A(D_REG_15__SCAN_IN), .B(keyinput_230), .ZN(n3224) );
  NAND3_X1 U3757 ( .A1(n3226), .A2(n3225), .A3(n3224), .ZN(n3229) );
  XNOR2_X1 U3758 ( .A(D_REG_16__SCAN_IN), .B(keyinput_231), .ZN(n3228) );
  XNOR2_X1 U3759 ( .A(D_REG_17__SCAN_IN), .B(keyinput_232), .ZN(n3227) );
  AOI21_X1 U3760 ( .B1(n3229), .B2(n3228), .A(n3227), .ZN(n3235) );
  INV_X1 U3761 ( .A(D_REG_18__SCAN_IN), .ZN(n4642) );
  XNOR2_X1 U3762 ( .A(n4642), .B(keyinput_233), .ZN(n3234) );
  INV_X1 U3763 ( .A(D_REG_21__SCAN_IN), .ZN(n4645) );
  XNOR2_X1 U3764 ( .A(n4645), .B(keyinput_236), .ZN(n3232) );
  XNOR2_X1 U3765 ( .A(D_REG_20__SCAN_IN), .B(keyinput_235), .ZN(n3231) );
  XNOR2_X1 U3766 ( .A(D_REG_19__SCAN_IN), .B(keyinput_234), .ZN(n3230) );
  NOR3_X1 U3767 ( .A1(n3232), .A2(n3231), .A3(n3230), .ZN(n3233) );
  OAI21_X1 U3768 ( .B1(n3235), .B2(n3234), .A(n3233), .ZN(n3238) );
  XNOR2_X1 U3769 ( .A(D_REG_22__SCAN_IN), .B(keyinput_237), .ZN(n3237) );
  XNOR2_X1 U3770 ( .A(D_REG_23__SCAN_IN), .B(keyinput_238), .ZN(n3236) );
  AOI21_X1 U3771 ( .B1(n3238), .B2(n3237), .A(n3236), .ZN(n3241) );
  INV_X1 U3772 ( .A(D_REG_24__SCAN_IN), .ZN(n4648) );
  XNOR2_X1 U3773 ( .A(n4648), .B(keyinput_239), .ZN(n3240) );
  INV_X1 U3774 ( .A(D_REG_25__SCAN_IN), .ZN(n4649) );
  XNOR2_X1 U3775 ( .A(n4649), .B(keyinput_240), .ZN(n3239) );
  NOR3_X1 U3776 ( .A1(n3241), .A2(n3240), .A3(n3239), .ZN(n3244) );
  INV_X1 U3777 ( .A(D_REG_27__SCAN_IN), .ZN(n4651) );
  XNOR2_X1 U3778 ( .A(n4651), .B(keyinput_242), .ZN(n3243) );
  XNOR2_X1 U3779 ( .A(D_REG_26__SCAN_IN), .B(keyinput_241), .ZN(n3242) );
  NOR3_X1 U3780 ( .A1(n3244), .A2(n3243), .A3(n3242), .ZN(n3251) );
  XOR2_X1 U3781 ( .A(D_REG_28__SCAN_IN), .B(keyinput_243), .Z(n3250) );
  XOR2_X1 U3782 ( .A(REG0_REG_0__SCAN_IN), .B(keyinput_247), .Z(n3248) );
  INV_X1 U3783 ( .A(D_REG_31__SCAN_IN), .ZN(n4655) );
  XNOR2_X1 U3784 ( .A(n4655), .B(keyinput_246), .ZN(n3247) );
  XNOR2_X1 U3785 ( .A(D_REG_29__SCAN_IN), .B(keyinput_244), .ZN(n3246) );
  XNOR2_X1 U3786 ( .A(D_REG_30__SCAN_IN), .B(keyinput_245), .ZN(n3245) );
  NOR4_X1 U3787 ( .A1(n3248), .A2(n3247), .A3(n3246), .A4(n3245), .ZN(n3249)
         );
  OAI21_X1 U3788 ( .B1(n3251), .B2(n3250), .A(n3249), .ZN(n3254) );
  XNOR2_X1 U3789 ( .A(REG0_REG_1__SCAN_IN), .B(keyinput_248), .ZN(n3253) );
  XOR2_X1 U3790 ( .A(REG0_REG_2__SCAN_IN), .B(keyinput_249), .Z(n3252) );
  AOI21_X1 U3791 ( .B1(n3254), .B2(n3253), .A(n3252), .ZN(n3260) );
  INV_X1 U3792 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4939) );
  AOI22_X1 U3793 ( .A1(REG0_REG_4__SCAN_IN), .A2(keyinput_251), .B1(n4939), 
        .B2(keyinput_254), .ZN(n3255) );
  OAI221_X1 U3794 ( .B1(REG0_REG_4__SCAN_IN), .B2(keyinput_251), .C1(n4939), 
        .C2(keyinput_254), .A(n3255), .ZN(n3259) );
  INV_X1 U3795 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4921) );
  AOI22_X1 U3796 ( .A1(REG0_REG_3__SCAN_IN), .A2(keyinput_250), .B1(n4921), 
        .B2(keyinput_252), .ZN(n3256) );
  OAI221_X1 U3797 ( .B1(REG0_REG_3__SCAN_IN), .B2(keyinput_250), .C1(n4921), 
        .C2(keyinput_252), .A(n3256), .ZN(n3258) );
  XNOR2_X1 U3798 ( .A(REG0_REG_6__SCAN_IN), .B(keyinput_253), .ZN(n3257) );
  NOR4_X1 U3799 ( .A1(n3260), .A2(n3259), .A3(n3258), .A4(n3257), .ZN(n3460)
         );
  XNOR2_X1 U3800 ( .A(REG0_REG_8__SCAN_IN), .B(keyinput_255), .ZN(n3459) );
  XNOR2_X1 U3801 ( .A(REG0_REG_8__SCAN_IN), .B(keyinput_127), .ZN(n3458) );
  XOR2_X1 U3802 ( .A(DATAI_29_), .B(keyinput_2), .Z(n3264) );
  XNOR2_X1 U3803 ( .A(DATAI_31_), .B(keyinput_0), .ZN(n3263) );
  XNOR2_X1 U3804 ( .A(DATAI_30_), .B(keyinput_1), .ZN(n3262) );
  XNOR2_X1 U3805 ( .A(DATAI_28_), .B(keyinput_3), .ZN(n3261) );
  NOR4_X1 U3806 ( .A1(n3264), .A2(n3263), .A3(n3262), .A4(n3261), .ZN(n3267)
         );
  XNOR2_X1 U3807 ( .A(DATAI_27_), .B(keyinput_4), .ZN(n3266) );
  XOR2_X1 U3808 ( .A(DATAI_26_), .B(keyinput_5), .Z(n3265) );
  OAI21_X1 U3809 ( .B1(n3267), .B2(n3266), .A(n3265), .ZN(n3271) );
  XOR2_X1 U3810 ( .A(DATAI_25_), .B(keyinput_6), .Z(n3270) );
  XOR2_X1 U3811 ( .A(DATAI_23_), .B(keyinput_8), .Z(n3269) );
  XNOR2_X1 U3812 ( .A(DATAI_24_), .B(keyinput_7), .ZN(n3268) );
  AOI211_X1 U3813 ( .C1(n3271), .C2(n3270), .A(n3269), .B(n3268), .ZN(n3273)
         );
  XOR2_X1 U3814 ( .A(DATAI_22_), .B(keyinput_9), .Z(n3272) );
  NOR2_X1 U3815 ( .A1(n3273), .A2(n3272), .ZN(n3281) );
  AOI22_X1 U3816 ( .A1(DATAI_17_), .A2(keyinput_14), .B1(n3275), .B2(
        keyinput_11), .ZN(n3274) );
  OAI221_X1 U3817 ( .B1(DATAI_17_), .B2(keyinput_14), .C1(n3275), .C2(
        keyinput_11), .A(n3274), .ZN(n3280) );
  INV_X1 U3818 ( .A(DATAI_18_), .ZN(n3277) );
  AOI22_X1 U3819 ( .A1(DATAI_21_), .A2(keyinput_10), .B1(n3277), .B2(
        keyinput_13), .ZN(n3276) );
  OAI221_X1 U3820 ( .B1(DATAI_21_), .B2(keyinput_10), .C1(n3277), .C2(
        keyinput_13), .A(n3276), .ZN(n3279) );
  XNOR2_X1 U3821 ( .A(DATAI_19_), .B(keyinput_12), .ZN(n3278) );
  NOR4_X1 U3822 ( .A1(n3281), .A2(n3280), .A3(n3279), .A4(n3278), .ZN(n3285)
         );
  XNOR2_X1 U3823 ( .A(DATAI_16_), .B(keyinput_15), .ZN(n3284) );
  XNOR2_X1 U3824 ( .A(n5051), .B(keyinput_17), .ZN(n3283) );
  XNOR2_X1 U3825 ( .A(DATAI_15_), .B(keyinput_16), .ZN(n3282) );
  OAI211_X1 U3826 ( .C1(n3285), .C2(n3284), .A(n3283), .B(n3282), .ZN(n3288)
         );
  XOR2_X1 U3827 ( .A(DATAI_13_), .B(keyinput_18), .Z(n3287) );
  XOR2_X1 U3828 ( .A(DATAI_12_), .B(keyinput_19), .Z(n3286) );
  NAND3_X1 U3829 ( .A1(n3288), .A2(n3287), .A3(n3286), .ZN(n3298) );
  INV_X1 U3830 ( .A(DATAI_9_), .ZN(n3290) );
  OAI22_X1 U3831 ( .A1(n3290), .A2(keyinput_22), .B1(DATAI_11_), .B2(
        keyinput_20), .ZN(n3289) );
  AOI221_X1 U3832 ( .B1(n3290), .B2(keyinput_22), .C1(keyinput_20), .C2(
        DATAI_11_), .A(n3289), .ZN(n3297) );
  INV_X1 U3833 ( .A(keyinput_21), .ZN(n3295) );
  XNOR2_X1 U3834 ( .A(DATAI_7_), .B(keyinput_24), .ZN(n3294) );
  INV_X1 U3835 ( .A(DATAI_8_), .ZN(n4941) );
  AOI22_X1 U3836 ( .A1(n4941), .A2(keyinput_23), .B1(n3291), .B2(keyinput_21), 
        .ZN(n3292) );
  OAI21_X1 U3837 ( .B1(n4941), .B2(keyinput_23), .A(n3292), .ZN(n3293) );
  AOI211_X1 U3838 ( .C1(DATAI_10_), .C2(n3295), .A(n3294), .B(n3293), .ZN(
        n3296) );
  NAND3_X1 U3839 ( .A1(n3298), .A2(n3297), .A3(n3296), .ZN(n3301) );
  XOR2_X1 U3840 ( .A(DATAI_6_), .B(keyinput_25), .Z(n3300) );
  XOR2_X1 U3841 ( .A(DATAI_5_), .B(keyinput_26), .Z(n3299) );
  AOI21_X1 U3842 ( .B1(n3301), .B2(n3300), .A(n3299), .ZN(n3305) );
  XNOR2_X1 U3843 ( .A(DATAI_4_), .B(keyinput_27), .ZN(n3304) );
  XOR2_X1 U3844 ( .A(DATAI_2_), .B(keyinput_29), .Z(n3303) );
  XNOR2_X1 U3845 ( .A(DATAI_3_), .B(keyinput_28), .ZN(n3302) );
  OAI211_X1 U3846 ( .C1(n3305), .C2(n3304), .A(n3303), .B(n3302), .ZN(n3313)
         );
  XNOR2_X1 U3847 ( .A(n3306), .B(keyinput_30), .ZN(n3312) );
  XOR2_X1 U3848 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_33), .Z(n3310) );
  XOR2_X1 U3849 ( .A(DATAI_0_), .B(keyinput_31), .Z(n3309) );
  XNOR2_X1 U3850 ( .A(U3149), .B(keyinput_32), .ZN(n3308) );
  XNOR2_X1 U3851 ( .A(n4033), .B(keyinput_34), .ZN(n3307) );
  NAND4_X1 U3852 ( .A1(n3310), .A2(n3309), .A3(n3308), .A4(n3307), .ZN(n3311)
         );
  AOI21_X1 U3853 ( .B1(n3313), .B2(n3312), .A(n3311), .ZN(n3316) );
  XNOR2_X1 U3854 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput_35), .ZN(n3315) );
  XNOR2_X1 U3855 ( .A(n3770), .B(keyinput_36), .ZN(n3314) );
  OAI21_X1 U3856 ( .B1(n3316), .B2(n3315), .A(n3314), .ZN(n3321) );
  XNOR2_X1 U3857 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_38), .ZN(n3318) );
  XNOR2_X1 U3858 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput_37), .ZN(n3317) );
  NOR2_X1 U3859 ( .A1(n3318), .A2(n3317), .ZN(n3320) );
  XNOR2_X1 U3860 ( .A(n3880), .B(keyinput_39), .ZN(n3319) );
  AOI21_X1 U3861 ( .B1(n3321), .B2(n3320), .A(n3319), .ZN(n3328) );
  XNOR2_X1 U3862 ( .A(n4022), .B(keyinput_40), .ZN(n3327) );
  XOR2_X1 U3863 ( .A(REG3_REG_12__SCAN_IN), .B(keyinput_44), .Z(n3325) );
  XOR2_X1 U3864 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_42), .Z(n3324) );
  XNOR2_X1 U3865 ( .A(n3512), .B(keyinput_41), .ZN(n3323) );
  XNOR2_X1 U3866 ( .A(REG3_REG_21__SCAN_IN), .B(keyinput_43), .ZN(n3322) );
  NOR4_X1 U3867 ( .A1(n3325), .A2(n3324), .A3(n3323), .A4(n3322), .ZN(n3326)
         );
  OAI21_X1 U3868 ( .B1(n3328), .B2(n3327), .A(n3326), .ZN(n3332) );
  XNOR2_X1 U3869 ( .A(REG3_REG_25__SCAN_IN), .B(keyinput_45), .ZN(n3331) );
  XNOR2_X1 U3870 ( .A(REG3_REG_16__SCAN_IN), .B(keyinput_46), .ZN(n3330) );
  XNOR2_X1 U3871 ( .A(REG3_REG_5__SCAN_IN), .B(keyinput_47), .ZN(n3329) );
  AOI211_X1 U3872 ( .C1(n3332), .C2(n3331), .A(n3330), .B(n3329), .ZN(n3335)
         );
  XOR2_X1 U3873 ( .A(REG3_REG_17__SCAN_IN), .B(keyinput_48), .Z(n3334) );
  INV_X1 U3874 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4095) );
  XNOR2_X1 U3875 ( .A(n4095), .B(keyinput_49), .ZN(n3333) );
  OAI21_X1 U3876 ( .B1(n3335), .B2(n3334), .A(n3333), .ZN(n3338) );
  XNOR2_X1 U3877 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_50), .ZN(n3337) );
  XNOR2_X1 U3878 ( .A(n3595), .B(keyinput_51), .ZN(n3336) );
  AOI21_X1 U3879 ( .B1(n3338), .B2(n3337), .A(n3336), .ZN(n3346) );
  XNOR2_X1 U3880 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_52), .ZN(n3345) );
  XNOR2_X1 U3881 ( .A(n3339), .B(keyinput_56), .ZN(n3343) );
  XNOR2_X1 U3882 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput_53), .ZN(n3342) );
  XOR2_X1 U3883 ( .A(REG3_REG_13__SCAN_IN), .B(keyinput_54), .Z(n3341) );
  XNOR2_X1 U3884 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_55), .ZN(n3340) );
  NOR4_X1 U3885 ( .A1(n3343), .A2(n3342), .A3(n3341), .A4(n3340), .ZN(n3344)
         );
  OAI21_X1 U3886 ( .B1(n3346), .B2(n3345), .A(n3344), .ZN(n3360) );
  XNOR2_X1 U3887 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_57), .ZN(n3359) );
  AOI22_X1 U3888 ( .A1(IR_REG_5__SCAN_IN), .A2(keyinput_60), .B1(n3348), .B2(
        keyinput_62), .ZN(n3347) );
  OAI221_X1 U3889 ( .B1(IR_REG_5__SCAN_IN), .B2(keyinput_60), .C1(n3348), .C2(
        keyinput_62), .A(n3347), .ZN(n3358) );
  OAI22_X1 U3890 ( .A1(IR_REG_4__SCAN_IN), .A2(keyinput_59), .B1(keyinput_64), 
        .B2(IR_REG_9__SCAN_IN), .ZN(n3350) );
  AND2_X1 U3891 ( .A1(IR_REG_4__SCAN_IN), .A2(keyinput_59), .ZN(n3349) );
  AOI211_X1 U3892 ( .C1(keyinput_64), .C2(IR_REG_9__SCAN_IN), .A(n3350), .B(
        n3349), .ZN(n3356) );
  XNOR2_X1 U3893 ( .A(n3351), .B(keyinput_63), .ZN(n3355) );
  XNOR2_X1 U3894 ( .A(n3352), .B(keyinput_61), .ZN(n3354) );
  XNOR2_X1 U3895 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_58), .ZN(n3353) );
  NAND4_X1 U3896 ( .A1(n3356), .A2(n3355), .A3(n3354), .A4(n3353), .ZN(n3357)
         );
  AOI211_X1 U3897 ( .C1(n3360), .C2(n3359), .A(n3358), .B(n3357), .ZN(n3363)
         );
  XNOR2_X1 U3898 ( .A(IR_REG_10__SCAN_IN), .B(keyinput_65), .ZN(n3362) );
  XNOR2_X1 U3899 ( .A(IR_REG_11__SCAN_IN), .B(keyinput_66), .ZN(n3361) );
  NOR3_X1 U3900 ( .A1(n3363), .A2(n3362), .A3(n3361), .ZN(n3367) );
  XNOR2_X1 U3901 ( .A(IR_REG_12__SCAN_IN), .B(keyinput_67), .ZN(n3366) );
  XNOR2_X1 U3902 ( .A(IR_REG_13__SCAN_IN), .B(keyinput_68), .ZN(n3365) );
  XNOR2_X1 U3903 ( .A(IR_REG_14__SCAN_IN), .B(keyinput_69), .ZN(n3364) );
  OAI211_X1 U3904 ( .C1(n3367), .C2(n3366), .A(n3365), .B(n3364), .ZN(n3386)
         );
  INV_X1 U3905 ( .A(keyinput_75), .ZN(n3373) );
  AOI22_X1 U3906 ( .A1(n3377), .A2(keyinput_74), .B1(n2762), .B2(keyinput_77), 
        .ZN(n3371) );
  AOI22_X1 U3907 ( .A1(IR_REG_16__SCAN_IN), .A2(keyinput_71), .B1(n3376), .B2(
        keyinput_72), .ZN(n3370) );
  AOI22_X1 U3908 ( .A1(IR_REG_18__SCAN_IN), .A2(keyinput_73), .B1(
        IR_REG_20__SCAN_IN), .B2(keyinput_75), .ZN(n3369) );
  AOI22_X1 U3909 ( .A1(IR_REG_15__SCAN_IN), .A2(keyinput_70), .B1(
        IR_REG_21__SCAN_IN), .B2(keyinput_76), .ZN(n3368) );
  NAND4_X1 U3910 ( .A1(n3371), .A2(n3370), .A3(n3369), .A4(n3368), .ZN(n3372)
         );
  AOI21_X1 U3911 ( .B1(n3374), .B2(n3373), .A(n3372), .ZN(n3375) );
  OAI21_X1 U3912 ( .B1(IR_REG_16__SCAN_IN), .B2(keyinput_71), .A(n3375), .ZN(
        n3381) );
  OAI22_X1 U3913 ( .A1(keyinput_72), .A2(n3376), .B1(n2762), .B2(keyinput_77), 
        .ZN(n3380) );
  OAI22_X1 U3914 ( .A1(n3377), .A2(keyinput_74), .B1(IR_REG_21__SCAN_IN), .B2(
        keyinput_76), .ZN(n3379) );
  OAI22_X1 U3915 ( .A1(IR_REG_18__SCAN_IN), .A2(keyinput_73), .B1(
        IR_REG_15__SCAN_IN), .B2(keyinput_70), .ZN(n3378) );
  NOR4_X1 U3916 ( .A1(n3381), .A2(n3380), .A3(n3379), .A4(n3378), .ZN(n3385)
         );
  XNOR2_X1 U3917 ( .A(n3382), .B(keyinput_78), .ZN(n3384) );
  XNOR2_X1 U3918 ( .A(IR_REG_24__SCAN_IN), .B(keyinput_79), .ZN(n3383) );
  AOI211_X1 U3919 ( .C1(n3386), .C2(n3385), .A(n3384), .B(n3383), .ZN(n3390)
         );
  XNOR2_X1 U3920 ( .A(n3387), .B(keyinput_80), .ZN(n3389) );
  XNOR2_X1 U3921 ( .A(IR_REG_26__SCAN_IN), .B(keyinput_81), .ZN(n3388) );
  OAI21_X1 U3922 ( .B1(n3390), .B2(n3389), .A(n3388), .ZN(n3398) );
  XOR2_X1 U3923 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_86), .Z(n3394) );
  XNOR2_X1 U3924 ( .A(n3391), .B(keyinput_82), .ZN(n3393) );
  XNOR2_X1 U3925 ( .A(IR_REG_29__SCAN_IN), .B(keyinput_84), .ZN(n3392) );
  NOR3_X1 U3926 ( .A1(n3394), .A2(n3393), .A3(n3392), .ZN(n3397) );
  XNOR2_X1 U3927 ( .A(IR_REG_30__SCAN_IN), .B(keyinput_85), .ZN(n3396) );
  XNOR2_X1 U3928 ( .A(IR_REG_28__SCAN_IN), .B(keyinput_83), .ZN(n3395) );
  NAND4_X1 U3929 ( .A1(n3398), .A2(n3397), .A3(n3396), .A4(n3395), .ZN(n3403)
         );
  XNOR2_X1 U3930 ( .A(n3399), .B(keyinput_87), .ZN(n3402) );
  XOR2_X1 U3931 ( .A(D_REG_2__SCAN_IN), .B(keyinput_89), .Z(n3401) );
  XNOR2_X1 U3932 ( .A(D_REG_1__SCAN_IN), .B(keyinput_88), .ZN(n3400) );
  NAND4_X1 U3933 ( .A1(n3403), .A2(n3402), .A3(n3401), .A4(n3400), .ZN(n3406)
         );
  XNOR2_X1 U3934 ( .A(D_REG_4__SCAN_IN), .B(keyinput_91), .ZN(n3405) );
  XNOR2_X1 U3935 ( .A(D_REG_3__SCAN_IN), .B(keyinput_90), .ZN(n3404) );
  NAND3_X1 U3936 ( .A1(n3406), .A2(n3405), .A3(n3404), .ZN(n3409) );
  XNOR2_X1 U3937 ( .A(n4633), .B(keyinput_93), .ZN(n3408) );
  XNOR2_X1 U3938 ( .A(D_REG_5__SCAN_IN), .B(keyinput_92), .ZN(n3407) );
  NAND3_X1 U3939 ( .A1(n3409), .A2(n3408), .A3(n3407), .ZN(n3412) );
  XNOR2_X1 U3940 ( .A(n4634), .B(keyinput_94), .ZN(n3411) );
  XNOR2_X1 U3941 ( .A(D_REG_8__SCAN_IN), .B(keyinput_95), .ZN(n3410) );
  AOI21_X1 U3942 ( .B1(n3412), .B2(n3411), .A(n3410), .ZN(n3415) );
  XNOR2_X1 U3943 ( .A(n4636), .B(keyinput_96), .ZN(n3414) );
  INV_X1 U3944 ( .A(D_REG_10__SCAN_IN), .ZN(n4637) );
  XNOR2_X1 U3945 ( .A(n4637), .B(keyinput_97), .ZN(n3413) );
  NOR3_X1 U3946 ( .A1(n3415), .A2(n3414), .A3(n3413), .ZN(n3419) );
  XNOR2_X1 U3947 ( .A(D_REG_11__SCAN_IN), .B(keyinput_98), .ZN(n3418) );
  XNOR2_X1 U3948 ( .A(D_REG_13__SCAN_IN), .B(keyinput_100), .ZN(n3417) );
  XNOR2_X1 U3949 ( .A(D_REG_12__SCAN_IN), .B(keyinput_99), .ZN(n3416) );
  NOR4_X1 U3950 ( .A1(n3419), .A2(n3418), .A3(n3417), .A4(n3416), .ZN(n3422)
         );
  INV_X1 U3951 ( .A(D_REG_15__SCAN_IN), .ZN(n4639) );
  XNOR2_X1 U3952 ( .A(n4639), .B(keyinput_102), .ZN(n3421) );
  XNOR2_X1 U3953 ( .A(D_REG_14__SCAN_IN), .B(keyinput_101), .ZN(n3420) );
  NOR3_X1 U3954 ( .A1(n3422), .A2(n3421), .A3(n3420), .ZN(n3425) );
  XNOR2_X1 U3955 ( .A(D_REG_16__SCAN_IN), .B(keyinput_103), .ZN(n3424) );
  INV_X1 U3956 ( .A(D_REG_17__SCAN_IN), .ZN(n4641) );
  XNOR2_X1 U3957 ( .A(n4641), .B(keyinput_104), .ZN(n3423) );
  OAI21_X1 U3958 ( .B1(n3425), .B2(n3424), .A(n3423), .ZN(n3431) );
  XNOR2_X1 U3959 ( .A(D_REG_18__SCAN_IN), .B(keyinput_105), .ZN(n3430) );
  XNOR2_X1 U3960 ( .A(n4645), .B(keyinput_108), .ZN(n3428) );
  XNOR2_X1 U3961 ( .A(D_REG_19__SCAN_IN), .B(keyinput_106), .ZN(n3427) );
  XNOR2_X1 U3962 ( .A(D_REG_20__SCAN_IN), .B(keyinput_107), .ZN(n3426) );
  NAND3_X1 U3963 ( .A1(n3428), .A2(n3427), .A3(n3426), .ZN(n3429) );
  AOI21_X1 U3964 ( .B1(n3431), .B2(n3430), .A(n3429), .ZN(n3434) );
  INV_X1 U3965 ( .A(D_REG_22__SCAN_IN), .ZN(n4646) );
  XNOR2_X1 U3966 ( .A(n4646), .B(keyinput_109), .ZN(n3433) );
  INV_X1 U3967 ( .A(D_REG_23__SCAN_IN), .ZN(n4647) );
  XNOR2_X1 U3968 ( .A(n4647), .B(keyinput_110), .ZN(n3432) );
  OAI21_X1 U3969 ( .B1(n3434), .B2(n3433), .A(n3432), .ZN(n3437) );
  XNOR2_X1 U3970 ( .A(n4649), .B(keyinput_112), .ZN(n3436) );
  XNOR2_X1 U3971 ( .A(n4648), .B(keyinput_111), .ZN(n3435) );
  NAND3_X1 U3972 ( .A1(n3437), .A2(n3436), .A3(n3435), .ZN(n3440) );
  XNOR2_X1 U3973 ( .A(D_REG_26__SCAN_IN), .B(keyinput_113), .ZN(n3439) );
  XNOR2_X1 U3974 ( .A(D_REG_27__SCAN_IN), .B(keyinput_114), .ZN(n3438) );
  NAND3_X1 U3975 ( .A1(n3440), .A2(n3439), .A3(n3438), .ZN(n3447) );
  XNOR2_X1 U3976 ( .A(D_REG_28__SCAN_IN), .B(keyinput_115), .ZN(n3446) );
  XNOR2_X1 U3977 ( .A(D_REG_30__SCAN_IN), .B(keyinput_117), .ZN(n3444) );
  XNOR2_X1 U3978 ( .A(D_REG_29__SCAN_IN), .B(keyinput_116), .ZN(n3443) );
  XNOR2_X1 U3979 ( .A(D_REG_31__SCAN_IN), .B(keyinput_118), .ZN(n3442) );
  XNOR2_X1 U3980 ( .A(REG0_REG_0__SCAN_IN), .B(keyinput_119), .ZN(n3441) );
  NAND4_X1 U3981 ( .A1(n3444), .A2(n3443), .A3(n3442), .A4(n3441), .ZN(n3445)
         );
  AOI21_X1 U3982 ( .B1(n3447), .B2(n3446), .A(n3445), .ZN(n3450) );
  XNOR2_X1 U3983 ( .A(REG0_REG_1__SCAN_IN), .B(keyinput_120), .ZN(n3449) );
  XNOR2_X1 U3984 ( .A(REG0_REG_2__SCAN_IN), .B(keyinput_121), .ZN(n3448) );
  OAI21_X1 U3985 ( .B1(n3450), .B2(n3449), .A(n3448), .ZN(n3456) );
  OAI22_X1 U3986 ( .A1(n4939), .A2(keyinput_126), .B1(REG0_REG_3__SCAN_IN), 
        .B2(keyinput_122), .ZN(n3451) );
  AOI221_X1 U3987 ( .B1(n4939), .B2(keyinput_126), .C1(keyinput_122), .C2(
        REG0_REG_3__SCAN_IN), .A(n3451), .ZN(n3455) );
  XOR2_X1 U3988 ( .A(REG0_REG_4__SCAN_IN), .B(keyinput_123), .Z(n3454) );
  OAI22_X1 U3989 ( .A1(n4921), .A2(keyinput_124), .B1(keyinput_125), .B2(
        REG0_REG_6__SCAN_IN), .ZN(n3452) );
  AOI221_X1 U3990 ( .B1(n4921), .B2(keyinput_124), .C1(REG0_REG_6__SCAN_IN), 
        .C2(keyinput_125), .A(n3452), .ZN(n3453) );
  NAND4_X1 U3991 ( .A1(n3456), .A2(n3455), .A3(n3454), .A4(n3453), .ZN(n3457)
         );
  OAI211_X1 U3992 ( .C1(n3460), .C2(n3459), .A(n3458), .B(n3457), .ZN(n3463)
         );
  MUX2_X1 U3993 ( .A(n3461), .B(DATAI_25_), .S(U3149), .Z(n3462) );
  XNOR2_X1 U3994 ( .A(n3463), .B(n3462), .ZN(U3327) );
  NAND2_X1 U3995 ( .A1(n2978), .A2(n3468), .ZN(n3471) );
  NAND2_X1 U3996 ( .A1(n4137), .A2(n3987), .ZN(n3470) );
  NAND2_X1 U3997 ( .A1(n3471), .A2(n3470), .ZN(n3472) );
  AOI22_X1 U3998 ( .A1(n2978), .A2(n4010), .B1(n4137), .B2(n3468), .ZN(n3473)
         );
  NAND2_X1 U3999 ( .A1(n3474), .A2(n3473), .ZN(n3476) );
  OAI21_X1 U4000 ( .B1(n3474), .B2(n3473), .A(n3476), .ZN(n3475) );
  INV_X1 U4001 ( .A(n3475), .ZN(n4134) );
  NAND2_X1 U4002 ( .A1(n4133), .A2(n4134), .ZN(n4132) );
  NAND2_X1 U4003 ( .A1(n4132), .A2(n3476), .ZN(n4059) );
  OAI22_X1 U4004 ( .A1(n3477), .A2(n2937), .B1(n3013), .B2(n4015), .ZN(n3482)
         );
  NAND2_X1 U4005 ( .A1(n4332), .A2(n3468), .ZN(n3479) );
  NAND2_X1 U4006 ( .A1(n4879), .A2(n3987), .ZN(n3478) );
  NAND2_X1 U4007 ( .A1(n3479), .A2(n3478), .ZN(n3480) );
  XNOR2_X1 U4008 ( .A(n3480), .B(n4016), .ZN(n3481) );
  XOR2_X1 U4009 ( .A(n3482), .B(n3481), .Z(n4060) );
  NAND2_X1 U4010 ( .A1(n4059), .A2(n4060), .ZN(n4058) );
  INV_X1 U4011 ( .A(n3481), .ZN(n3484) );
  INV_X1 U4012 ( .A(n3482), .ZN(n3483) );
  NAND2_X1 U4013 ( .A1(n3484), .A2(n3483), .ZN(n4103) );
  OAI22_X1 U4014 ( .A1(n3485), .A2(n4015), .B1(n2544), .B2(n2880), .ZN(n3486)
         );
  XNOR2_X1 U4015 ( .A(n3486), .B(n4016), .ZN(n3488) );
  AOI22_X1 U4016 ( .A1(n4331), .A2(n4010), .B1(n4108), .B2(n3468), .ZN(n3489)
         );
  XNOR2_X1 U4017 ( .A(n3488), .B(n3489), .ZN(n4105) );
  INV_X1 U4018 ( .A(n3489), .ZN(n3490) );
  NAND2_X1 U4019 ( .A1(n4330), .A2(n3468), .ZN(n3493) );
  NAND2_X1 U4020 ( .A1(n4913), .A2(n3987), .ZN(n3492) );
  NAND2_X1 U4021 ( .A1(n3493), .A2(n3492), .ZN(n3494) );
  XNOR2_X1 U4022 ( .A(n3494), .B(n3968), .ZN(n3496) );
  AOI22_X1 U4023 ( .A1(n4330), .A2(n4010), .B1(n4913), .B2(n3468), .ZN(n3495)
         );
  NAND2_X1 U4024 ( .A1(n3496), .A2(n3495), .ZN(n4142) );
  OAI21_X1 U4025 ( .B1(n3496), .B2(n3495), .A(n4142), .ZN(n4907) );
  OAI22_X1 U4026 ( .A1(n3541), .A2(n4015), .B1(n4149), .B2(n2880), .ZN(n3497)
         );
  XNOR2_X1 U4027 ( .A(n3497), .B(n4016), .ZN(n3501) );
  OAI22_X1 U4028 ( .A1(n3541), .A2(n2937), .B1(n4149), .B2(n4015), .ZN(n3502)
         );
  OR2_X1 U4029 ( .A1(n4141), .A2(n4142), .ZN(n3508) );
  NAND2_X1 U4030 ( .A1(n4327), .A2(n3468), .ZN(n3499) );
  MUX2_X1 U4031 ( .A(n4932), .B(DATAI_7_), .S(n2482), .Z(n3536) );
  NAND2_X1 U4032 ( .A1(n3536), .A2(n3987), .ZN(n3498) );
  NAND2_X1 U4033 ( .A1(n3499), .A2(n3498), .ZN(n3500) );
  XNOR2_X1 U4034 ( .A(n3500), .B(n4016), .ZN(n3583) );
  AOI22_X1 U4035 ( .A1(n4327), .A2(n4010), .B1(n3536), .B2(n3468), .ZN(n3581)
         );
  XNOR2_X1 U4036 ( .A(n3583), .B(n3581), .ZN(n3510) );
  INV_X1 U4037 ( .A(n3501), .ZN(n3504) );
  INV_X1 U4038 ( .A(n3502), .ZN(n3503) );
  NAND2_X1 U4039 ( .A1(n3504), .A2(n3503), .ZN(n3511) );
  NAND2_X1 U4040 ( .A1(n3509), .A2(n3507), .ZN(n3584) );
  NAND2_X1 U4041 ( .A1(n3584), .A2(n5162), .ZN(n3526) );
  AND2_X1 U4042 ( .A1(n3509), .A2(n3508), .ZN(n4143) );
  AOI21_X1 U40430 ( .B1(n4143), .B2(n3511), .A(n3510), .ZN(n3525) );
  NAND2_X1 U4044 ( .A1(n2485), .A2(REG2_REG_8__SCAN_IN), .ZN(n3519) );
  NAND2_X1 U4045 ( .A1(n3513), .A2(n3512), .ZN(n3514) );
  NAND2_X1 U4046 ( .A1(n3561), .A2(n3514), .ZN(n4954) );
  INV_X1 U4047 ( .A(n4954), .ZN(n3515) );
  NAND2_X1 U4048 ( .A1(n2982), .A2(n3515), .ZN(n3518) );
  NAND2_X1 U4049 ( .A1(n3858), .A2(REG0_REG_8__SCAN_IN), .ZN(n3517) );
  NAND2_X1 U4050 ( .A1(n4188), .A2(REG1_REG_8__SCAN_IN), .ZN(n3516) );
  NAND4_X1 U4051 ( .A1(n3519), .A2(n3518), .A3(n3517), .A4(n3516), .ZN(n4326)
         );
  AOI22_X1 U4052 ( .A1(n4148), .A2(n4326), .B1(n4160), .B2(n3537), .ZN(n3524)
         );
  INV_X1 U4053 ( .A(REG3_REG_7__SCAN_IN), .ZN(n3521) );
  NOR2_X1 U4054 ( .A1(STATE_REG_SCAN_IN), .A2(n3521), .ZN(n4713) );
  INV_X1 U4055 ( .A(n3536), .ZN(n3552) );
  NOR2_X1 U4056 ( .A1(n5185), .A2(n3552), .ZN(n3522) );
  AOI211_X1 U4057 ( .C1(n4151), .C2(n4329), .A(n4713), .B(n3522), .ZN(n3523)
         );
  OAI211_X1 U4058 ( .C1(n3526), .C2(n3525), .A(n3524), .B(n3523), .ZN(U3210)
         );
  AND2_X1 U4059 ( .A1(n3527), .A2(n4247), .ZN(n4270) );
  AOI21_X2 U4060 ( .B1(n3529), .B2(n4270), .A(n3528), .ZN(n3531) );
  INV_X1 U4061 ( .A(n4327), .ZN(n3551) );
  NAND2_X1 U4062 ( .A1(n3551), .A2(n3536), .ZN(n4273) );
  NAND2_X1 U4063 ( .A1(n4327), .A2(n3552), .ZN(n3603) );
  NAND2_X1 U4064 ( .A1(n4273), .A2(n3603), .ZN(n4234) );
  NAND2_X1 U4065 ( .A1(n3531), .A2(n3530), .ZN(n3604) );
  OAI211_X1 U4066 ( .C1(n3531), .C2(n3530), .A(n3604), .B(n5207), .ZN(n3533)
         );
  AOI22_X1 U4067 ( .A1(n4329), .A2(n4511), .B1(n5177), .B2(n4326), .ZN(n3532)
         );
  OAI211_X1 U4068 ( .C1(n5237), .C2(n3552), .A(n3533), .B(n3532), .ZN(n4935)
         );
  INV_X1 U4069 ( .A(n4935), .ZN(n3549) );
  INV_X1 U4070 ( .A(n3558), .ZN(n3535) );
  AOI211_X1 U4071 ( .C1(n3536), .C2(n3534), .A(n5219), .B(n3535), .ZN(n4936)
         );
  INV_X1 U4072 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3539) );
  INV_X1 U4073 ( .A(n3537), .ZN(n3538) );
  OAI22_X1 U4074 ( .A1(n4558), .A2(n3539), .B1(n3538), .B2(n5216), .ZN(n3547)
         );
  NAND2_X1 U4075 ( .A1(n4329), .A2(n3540), .ZN(n3543) );
  NOR2_X1 U4076 ( .A1(n2524), .A2(n4234), .ZN(n4934) );
  INV_X1 U4077 ( .A(n3554), .ZN(n3545) );
  NOR3_X1 U4078 ( .A1(n4934), .A2(n3545), .A3(n5103), .ZN(n3546) );
  AOI211_X1 U4079 ( .C1(n4524), .C2(n4936), .A(n3547), .B(n3546), .ZN(n3548)
         );
  OAI21_X1 U4080 ( .B1(n5246), .B2(n3549), .A(n3548), .ZN(U3283) );
  INV_X1 U4081 ( .A(n4326), .ZN(n3599) );
  INV_X1 U4082 ( .A(n4942), .ZN(n3550) );
  MUX2_X1 U4083 ( .A(n3550), .B(DATAI_8_), .S(n2977), .Z(n3577) );
  NAND2_X1 U4084 ( .A1(n3599), .A2(n3577), .ZN(n4965) );
  INV_X1 U4085 ( .A(n3577), .ZN(n4950) );
  NAND2_X1 U4086 ( .A1(n4326), .A2(n4950), .ZN(n3602) );
  NAND2_X1 U4087 ( .A1(n4327), .A2(n3536), .ZN(n3553) );
  NAND2_X1 U4088 ( .A1(n3554), .A2(n3553), .ZN(n3557) );
  INV_X1 U4089 ( .A(n3557), .ZN(n3556) );
  AOI21_X1 U4090 ( .B1(n4228), .B2(n3557), .A(n2523), .ZN(n4955) );
  AOI21_X1 U4091 ( .B1(n3577), .B2(n3558), .A(n4963), .ZN(n4958) );
  OAI22_X1 U4092 ( .A1(n4558), .A2(n2852), .B1(n4954), .B2(n5216), .ZN(n3559)
         );
  AOI21_X1 U4093 ( .B1(n4958), .B2(n5244), .A(n3559), .ZN(n3571) );
  NAND2_X1 U4094 ( .A1(n3604), .A2(n3603), .ZN(n3560) );
  XNOR2_X1 U4095 ( .A(n3560), .B(n4228), .ZN(n3569) );
  AND2_X1 U4096 ( .A1(n3561), .A2(n3595), .ZN(n3562) );
  OR2_X1 U4097 ( .A1(n3562), .A2(n3589), .ZN(n4987) );
  INV_X1 U4098 ( .A(n4987), .ZN(n3563) );
  AOI22_X1 U4099 ( .A1(n2982), .A2(n3563), .B1(n2483), .B2(REG1_REG_9__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4100 ( .A1(n2485), .A2(REG2_REG_9__SCAN_IN), .B1(n3858), .B2(
        REG0_REG_9__SCAN_IN), .ZN(n3564) );
  OR2_X1 U4101 ( .A1(n4238), .A2(n5121), .ZN(n3567) );
  NAND2_X1 U4102 ( .A1(n4327), .A2(n4511), .ZN(n3566) );
  NAND2_X1 U4103 ( .A1(n3567), .A2(n3566), .ZN(n4948) );
  AOI21_X1 U4104 ( .B1(n3577), .B2(n5229), .A(n4948), .ZN(n3568) );
  OAI21_X1 U4105 ( .B1(n3569), .B2(n5091), .A(n3568), .ZN(n4957) );
  NAND2_X1 U4106 ( .A1(n4957), .A2(n4558), .ZN(n3570) );
  OAI211_X1 U4107 ( .C1(n4955), .C2(n5103), .A(n3571), .B(n3570), .ZN(U3282)
         );
  MUX2_X1 U4108 ( .A(n3572), .B(n3290), .S(n2977), .Z(n4969) );
  OAI22_X1 U4109 ( .A1(n4238), .A2(n2937), .B1(n4969), .B2(n4015), .ZN(n3893)
         );
  OAI22_X1 U4110 ( .A1(n4238), .A2(n4015), .B1(n4969), .B2(n2880), .ZN(n3573)
         );
  XNOR2_X1 U4111 ( .A(n3573), .B(n4016), .ZN(n3892) );
  XOR2_X1 U4112 ( .A(n3893), .B(n3892), .Z(n3587) );
  NAND2_X1 U4113 ( .A1(n4326), .A2(n3468), .ZN(n3575) );
  NAND2_X1 U4114 ( .A1(n3577), .A2(n3987), .ZN(n3574) );
  NAND2_X1 U4115 ( .A1(n3575), .A2(n3574), .ZN(n3576) );
  XNOR2_X1 U4116 ( .A(n3576), .B(n3968), .ZN(n3579) );
  AOI22_X1 U4117 ( .A1(n4326), .A2(n4010), .B1(n3577), .B2(n3468), .ZN(n3578)
         );
  NAND2_X1 U4118 ( .A1(n3579), .A2(n3578), .ZN(n3585) );
  OAI21_X1 U4119 ( .B1(n3579), .B2(n3578), .A(n3585), .ZN(n3580) );
  INV_X1 U4120 ( .A(n3580), .ZN(n4945) );
  INV_X1 U4121 ( .A(n3581), .ZN(n3582) );
  NAND2_X1 U4122 ( .A1(n3583), .A2(n3582), .ZN(n4943) );
  NAND3_X1 U4123 ( .A1(n3584), .A2(n4945), .A3(n4943), .ZN(n4944) );
  NAND2_X1 U4124 ( .A1(n4944), .A2(n3585), .ZN(n3586) );
  NAND2_X1 U4125 ( .A1(n3586), .A2(n3587), .ZN(n3897) );
  OAI21_X1 U4126 ( .B1(n3587), .B2(n3586), .A(n3897), .ZN(n3588) );
  NAND2_X1 U4127 ( .A1(n3588), .A2(n5162), .ZN(n3598) );
  AOI22_X1 U4128 ( .A1(n2485), .A2(REG2_REG_10__SCAN_IN), .B1(n4188), .B2(
        REG1_REG_10__SCAN_IN), .ZN(n3592) );
  NOR2_X1 U4129 ( .A1(n3589), .A2(REG3_REG_10__SCAN_IN), .ZN(n3590) );
  OR2_X1 U4130 ( .A1(n3608), .A2(n3590), .ZN(n3619) );
  INV_X1 U4131 ( .A(n3619), .ZN(n4052) );
  AOI22_X1 U4132 ( .A1(n2982), .A2(n4052), .B1(n3858), .B2(
        REG0_REG_10__SCAN_IN), .ZN(n3591) );
  OR2_X1 U4133 ( .A1(n3889), .A2(n5121), .ZN(n3594) );
  NAND2_X1 U4134 ( .A1(n4326), .A2(n4511), .ZN(n3593) );
  NAND2_X1 U4135 ( .A1(n3594), .A2(n3593), .ZN(n4970) );
  NOR2_X1 U4136 ( .A1(STATE_REG_SCAN_IN), .A2(n3595), .ZN(n4722) );
  OAI22_X1 U4137 ( .A1(n5185), .A2(n4969), .B1(n4987), .B2(n5192), .ZN(n3596)
         );
  AOI211_X1 U4138 ( .C1(n5190), .C2(n4970), .A(n4722), .B(n3596), .ZN(n3597)
         );
  NAND2_X1 U4139 ( .A1(n3598), .A2(n3597), .ZN(U3228) );
  NAND2_X1 U4140 ( .A1(n3599), .A2(n4950), .ZN(n3600) );
  NAND2_X1 U4141 ( .A1(n4238), .A2(n4969), .ZN(n3601) );
  INV_X1 U4142 ( .A(n4969), .ZN(n3605) );
  MUX2_X1 U4143 ( .A(n4737), .B(DATAI_10_), .S(n2482), .Z(n4053) );
  NAND2_X1 U4144 ( .A1(n3889), .A2(n4053), .ZN(n4251) );
  INV_X1 U4145 ( .A(n3889), .ZN(n4324) );
  NAND2_X1 U4146 ( .A1(n4324), .A2(n3887), .ZN(n3685) );
  XNOR2_X1 U4147 ( .A(n3635), .B(n4229), .ZN(n4989) );
  AND2_X1 U4148 ( .A1(n3603), .A2(n3602), .ZN(n4246) );
  NAND2_X1 U4149 ( .A1(n3604), .A2(n4246), .ZN(n4966) );
  NAND2_X1 U4150 ( .A1(n4238), .A2(n3605), .ZN(n3606) );
  AND2_X1 U4151 ( .A1(n4965), .A2(n3606), .ZN(n4275) );
  NAND2_X1 U4152 ( .A1(n4966), .A2(n4275), .ZN(n3607) );
  NAND2_X1 U4153 ( .A1(n4325), .A2(n4969), .ZN(n4278) );
  XNOR2_X1 U4154 ( .A(n3623), .B(n4229), .ZN(n3617) );
  NAND2_X1 U4155 ( .A1(n2485), .A2(REG2_REG_11__SCAN_IN), .ZN(n3614) );
  OR2_X1 U4156 ( .A1(n3608), .A2(REG3_REG_11__SCAN_IN), .ZN(n3609) );
  NAND2_X1 U4157 ( .A1(n3609), .A2(n3626), .ZN(n5009) );
  INV_X1 U4158 ( .A(n5009), .ZN(n3610) );
  NAND2_X1 U4159 ( .A1(n2982), .A2(n3610), .ZN(n3613) );
  NAND2_X1 U4160 ( .A1(n3858), .A2(REG0_REG_11__SCAN_IN), .ZN(n3612) );
  NAND2_X1 U4161 ( .A1(n4188), .A2(REG1_REG_11__SCAN_IN), .ZN(n3611) );
  NAND4_X1 U4162 ( .A1(n3614), .A2(n3613), .A3(n3612), .A4(n3611), .ZN(n4323)
         );
  INV_X1 U4163 ( .A(n4323), .ZN(n3653) );
  OAI22_X1 U4164 ( .A1(n4238), .A2(n5175), .B1(n3653), .B2(n5121), .ZN(n3615)
         );
  AOI21_X1 U4165 ( .B1(n4053), .B2(n5229), .A(n3615), .ZN(n3616) );
  OAI21_X1 U4166 ( .B1(n3617), .B2(n5091), .A(n3616), .ZN(n4991) );
  OAI21_X1 U4167 ( .B1(n3618), .B2(n3887), .A(n3636), .ZN(n4988) );
  NOR2_X1 U4168 ( .A1(n4988), .A2(n5196), .ZN(n3621) );
  OAI22_X1 U4169 ( .A1(n4558), .A2(n4732), .B1(n3619), .B2(n5216), .ZN(n3620)
         );
  AOI211_X1 U4170 ( .C1(n4991), .C2(n4558), .A(n3621), .B(n3620), .ZN(n3622)
         );
  OAI21_X1 U4171 ( .B1(n4989), .B2(n5103), .A(n3622), .ZN(U3280) );
  MUX2_X1 U4172 ( .A(n4995), .B(DATAI_11_), .S(n2977), .Z(n5006) );
  NAND2_X1 U4173 ( .A1(n3653), .A2(n5006), .ZN(n3689) );
  INV_X1 U4174 ( .A(n5006), .ZN(n3624) );
  NAND2_X1 U4175 ( .A1(n4323), .A2(n3624), .ZN(n3686) );
  NAND2_X1 U4176 ( .A1(n3623), .A2(n4251), .ZN(n3688) );
  NAND2_X1 U4177 ( .A1(n3688), .A2(n3685), .ZN(n3647) );
  XOR2_X1 U4178 ( .A(n4230), .B(n3647), .Z(n3634) );
  NOR2_X1 U4179 ( .A1(n3624), .A2(n5237), .ZN(n3633) );
  OR2_X1 U4180 ( .A1(n3889), .A2(n5175), .ZN(n3632) );
  AOI21_X1 U4181 ( .B1(n3626), .B2(n3625), .A(n3648), .ZN(n3658) );
  NAND2_X1 U4182 ( .A1(n2982), .A2(n3658), .ZN(n3630) );
  NAND2_X1 U4183 ( .A1(n2485), .A2(REG2_REG_12__SCAN_IN), .ZN(n3629) );
  NAND2_X1 U4184 ( .A1(n2483), .A2(REG1_REG_12__SCAN_IN), .ZN(n3628) );
  NAND2_X1 U4185 ( .A1(n3858), .A2(REG0_REG_12__SCAN_IN), .ZN(n3627) );
  NAND4_X1 U4186 ( .A1(n3630), .A2(n3629), .A3(n3628), .A4(n3627), .ZN(n4322)
         );
  NAND2_X1 U4187 ( .A1(n4322), .A2(n5177), .ZN(n3631) );
  NAND2_X1 U4188 ( .A1(n3632), .A2(n3631), .ZN(n4997) );
  AOI211_X1 U4189 ( .C1(n3634), .C2(n5207), .A(n3633), .B(n4997), .ZN(n5010)
         );
  XNOR2_X1 U4190 ( .A(n3643), .B(n4230), .ZN(n5013) );
  NAND2_X1 U4191 ( .A1(n5013), .A2(n5144), .ZN(n3642) );
  NAND2_X1 U4192 ( .A1(n3636), .A2(n5006), .ZN(n3637) );
  NAND2_X1 U4193 ( .A1(n3656), .A2(n3637), .ZN(n5011) );
  INV_X1 U4194 ( .A(n5011), .ZN(n3640) );
  INV_X1 U4195 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3638) );
  OAI22_X1 U4196 ( .A1(n4558), .A2(n3638), .B1(n5009), .B2(n5216), .ZN(n3639)
         );
  AOI21_X1 U4197 ( .B1(n3640), .B2(n5244), .A(n3639), .ZN(n3641) );
  OAI211_X1 U4198 ( .C1(n5246), .C2(n5010), .A(n3642), .B(n3641), .ZN(U3279)
         );
  OAI22_X1 U4199 ( .A1(n3643), .A2(n4230), .B1(n5006), .B2(n4323), .ZN(n3644)
         );
  INV_X1 U4200 ( .A(n4322), .ZN(n3911) );
  MUX2_X1 U4201 ( .A(n5017), .B(DATAI_12_), .S(n2482), .Z(n5022) );
  NAND2_X1 U4202 ( .A1(n3911), .A2(n5022), .ZN(n3690) );
  INV_X1 U4203 ( .A(n5022), .ZN(n3910) );
  NAND2_X1 U4204 ( .A1(n4322), .A2(n3910), .ZN(n3684) );
  NAND2_X1 U4205 ( .A1(n3690), .A2(n3684), .ZN(n4227) );
  NAND2_X1 U4206 ( .A1(n3644), .A2(n4227), .ZN(n3664) );
  OAI21_X1 U4207 ( .B1(n3644), .B2(n4227), .A(n3664), .ZN(n3645) );
  INV_X1 U4208 ( .A(n3645), .ZN(n5028) );
  INV_X1 U4209 ( .A(n3686), .ZN(n3646) );
  AOI21_X1 U4210 ( .B1(n3647), .B2(n4230), .A(n3646), .ZN(n3666) );
  XNOR2_X1 U4211 ( .A(n3666), .B(n4227), .ZN(n3655) );
  OAI21_X1 U4212 ( .B1(n3648), .B2(REG3_REG_13__SCAN_IN), .A(n3669), .ZN(n5043) );
  INV_X1 U4213 ( .A(n5043), .ZN(n3677) );
  NAND2_X1 U4214 ( .A1(n2982), .A2(n3677), .ZN(n3652) );
  NAND2_X1 U4215 ( .A1(n2485), .A2(REG2_REG_13__SCAN_IN), .ZN(n3651) );
  NAND2_X1 U4216 ( .A1(n2483), .A2(REG1_REG_13__SCAN_IN), .ZN(n3650) );
  NAND2_X1 U4217 ( .A1(n3858), .A2(REG0_REG_13__SCAN_IN), .ZN(n3649) );
  NAND4_X1 U4218 ( .A1(n3652), .A2(n3651), .A3(n3650), .A4(n3649), .ZN(n4321)
         );
  INV_X1 U4219 ( .A(n4321), .ZN(n3703) );
  OAI22_X1 U4220 ( .A1(n3653), .A2(n5175), .B1(n3703), .B2(n5121), .ZN(n5019)
         );
  AOI21_X1 U4221 ( .B1(n5022), .B2(n5229), .A(n5019), .ZN(n3654) );
  OAI21_X1 U4222 ( .B1(n3655), .B2(n5091), .A(n3654), .ZN(n5030) );
  INV_X1 U4223 ( .A(n3656), .ZN(n3657) );
  OAI21_X1 U4224 ( .B1(n3657), .B2(n3910), .A(n3676), .ZN(n5027) );
  NOR2_X1 U4225 ( .A1(n5027), .A2(n5196), .ZN(n3661) );
  INV_X1 U4226 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3659) );
  INV_X1 U4227 ( .A(n3658), .ZN(n5026) );
  OAI22_X1 U4228 ( .A1(n4558), .A2(n3659), .B1(n5026), .B2(n5216), .ZN(n3660)
         );
  AOI211_X1 U4229 ( .C1(n5030), .C2(n4558), .A(n3661), .B(n3660), .ZN(n3662)
         );
  OAI21_X1 U4230 ( .B1(n5028), .B2(n5103), .A(n3662), .ZN(U3278) );
  NAND2_X1 U4231 ( .A1(n3664), .A2(n3663), .ZN(n3721) );
  NAND2_X1 U4232 ( .A1(n4321), .A2(n5039), .ZN(n3718) );
  INV_X1 U4233 ( .A(n3718), .ZN(n3665) );
  OR2_X1 U4234 ( .A1(n3665), .A2(n3720), .ZN(n4224) );
  XNOR2_X1 U4235 ( .A(n3721), .B(n4224), .ZN(n5044) );
  OAI21_X1 U4236 ( .B1(n3666), .B2(n4227), .A(n3684), .ZN(n3667) );
  XNOR2_X1 U4237 ( .A(n3667), .B(n4224), .ZN(n3675) );
  NAND2_X1 U4238 ( .A1(n2485), .A2(REG2_REG_14__SCAN_IN), .ZN(n3673) );
  AOI21_X1 U4239 ( .B1(n3669), .B2(n3668), .A(n3698), .ZN(n5053) );
  NAND2_X1 U4240 ( .A1(n2982), .A2(n5053), .ZN(n3672) );
  NAND2_X1 U4241 ( .A1(n3858), .A2(REG0_REG_14__SCAN_IN), .ZN(n3671) );
  NAND2_X1 U4242 ( .A1(n2483), .A2(REG1_REG_14__SCAN_IN), .ZN(n3670) );
  NAND4_X1 U4243 ( .A1(n3673), .A2(n3672), .A3(n3671), .A4(n3670), .ZN(n4320)
         );
  OAI22_X1 U4244 ( .A1(n5070), .A2(n5121), .B1(n3911), .B2(n5175), .ZN(n5036)
         );
  AOI21_X1 U4245 ( .B1(n5039), .B2(n5229), .A(n5036), .ZN(n3674) );
  OAI21_X1 U4246 ( .B1(n3675), .B2(n5091), .A(n3674), .ZN(n5046) );
  AOI21_X1 U4247 ( .B1(n5039), .B2(n3676), .A(n3706), .ZN(n5047) );
  INV_X1 U4248 ( .A(n5047), .ZN(n3679) );
  AOI22_X1 U4249 ( .A1(n5246), .A2(REG2_REG_13__SCAN_IN), .B1(n5136), .B2(
        n3677), .ZN(n3678) );
  OAI21_X1 U4250 ( .B1(n3679), .B2(n5196), .A(n3678), .ZN(n3680) );
  AOI21_X1 U4251 ( .B1(n5046), .B2(n4558), .A(n3680), .ZN(n3681) );
  OAI21_X1 U4252 ( .B1(n5044), .B2(n5103), .A(n3681), .ZN(U3277) );
  AOI21_X1 U4253 ( .B1(n3721), .B2(n3718), .A(n3720), .ZN(n5080) );
  INV_X1 U4254 ( .A(n5052), .ZN(n3682) );
  MUX2_X1 U4255 ( .A(n3682), .B(DATAI_14_), .S(n4199), .Z(n5057) );
  NAND2_X1 U4256 ( .A1(n5070), .A2(n5057), .ZN(n5084) );
  NAND2_X1 U4257 ( .A1(n4320), .A2(n3924), .ZN(n3831) );
  NAND2_X1 U4258 ( .A1(n5084), .A2(n3831), .ZN(n4221) );
  XNOR2_X1 U4259 ( .A(n5080), .B(n5081), .ZN(n5066) );
  INV_X1 U4260 ( .A(n5066), .ZN(n3711) );
  INV_X1 U4261 ( .A(n5039), .ZN(n3691) );
  NAND2_X1 U4262 ( .A1(n4321), .A2(n3691), .ZN(n3683) );
  AND2_X1 U4263 ( .A1(n3684), .A2(n3683), .ZN(n3693) );
  AND2_X1 U4264 ( .A1(n3686), .A2(n3685), .ZN(n3687) );
  AND2_X1 U4265 ( .A1(n3693), .A2(n3687), .ZN(n4279) );
  NAND2_X1 U4266 ( .A1(n3688), .A2(n4279), .ZN(n3695) );
  NAND2_X1 U4267 ( .A1(n3690), .A2(n3689), .ZN(n3694) );
  NOR2_X1 U4268 ( .A1(n4321), .A2(n3691), .ZN(n3692) );
  AOI21_X1 U4269 ( .B1(n3694), .B2(n3693), .A(n3692), .ZN(n4254) );
  NAND2_X1 U4270 ( .A1(n3695), .A2(n4254), .ZN(n3696) );
  OAI21_X1 U4271 ( .B1(n5081), .B2(n3696), .A(n5085), .ZN(n3697) );
  NAND2_X1 U4272 ( .A1(n3697), .A2(n5207), .ZN(n3705) );
  NAND2_X1 U4273 ( .A1(n3698), .A2(REG3_REG_15__SCAN_IN), .ZN(n3712) );
  OAI21_X1 U4274 ( .B1(n3698), .B2(REG3_REG_15__SCAN_IN), .A(n3712), .ZN(n5078) );
  INV_X1 U4275 ( .A(n5078), .ZN(n5097) );
  NAND2_X1 U4276 ( .A1(n2982), .A2(n5097), .ZN(n3702) );
  NAND2_X1 U4277 ( .A1(n2485), .A2(REG2_REG_15__SCAN_IN), .ZN(n3701) );
  NAND2_X1 U4278 ( .A1(n4188), .A2(REG1_REG_15__SCAN_IN), .ZN(n3700) );
  NAND2_X1 U4279 ( .A1(n3858), .A2(REG0_REG_15__SCAN_IN), .ZN(n3699) );
  NAND4_X1 U4280 ( .A1(n3702), .A2(n3701), .A3(n3700), .A4(n3699), .ZN(n4319)
         );
  INV_X1 U4281 ( .A(n4319), .ZN(n4550) );
  OAI22_X1 U4282 ( .A1(n3703), .A2(n5175), .B1(n4550), .B2(n5121), .ZN(n5054)
         );
  INV_X1 U4283 ( .A(n5054), .ZN(n3704) );
  OAI211_X1 U4284 ( .C1(n5237), .C2(n3924), .A(n3705), .B(n3704), .ZN(n5062)
         );
  NAND2_X1 U4285 ( .A1(n3706), .A2(n3924), .ZN(n3826) );
  OR2_X1 U4286 ( .A1(n3706), .A2(n3924), .ZN(n3707) );
  NAND2_X1 U4287 ( .A1(n3826), .A2(n3707), .ZN(n5064) );
  AOI22_X1 U4288 ( .A1(n5246), .A2(REG2_REG_14__SCAN_IN), .B1(n5136), .B2(
        n5053), .ZN(n3708) );
  OAI21_X1 U4289 ( .B1(n5064), .B2(n5196), .A(n3708), .ZN(n3709) );
  AOI21_X1 U4290 ( .B1(n5062), .B2(n4558), .A(n3709), .ZN(n3710) );
  OAI21_X1 U4291 ( .B1(n3711), .B2(n5103), .A(n3710), .ZN(U3276) );
  NAND2_X1 U4292 ( .A1(n3739), .A2(REG3_REG_18__SCAN_IN), .ZN(n3742) );
  NOR2_X1 U4293 ( .A1(n3753), .A2(REG3_REG_21__SCAN_IN), .ZN(n3713) );
  OR2_X1 U4294 ( .A1(n3766), .A2(n3713), .ZN(n4499) );
  INV_X1 U4295 ( .A(n4499), .ZN(n4072) );
  NAND2_X1 U4296 ( .A1(n4072), .A2(n2487), .ZN(n3717) );
  NAND2_X1 U4297 ( .A1(n2483), .A2(REG1_REG_21__SCAN_IN), .ZN(n3716) );
  NAND2_X1 U4298 ( .A1(n3858), .A2(REG0_REG_21__SCAN_IN), .ZN(n3715) );
  NAND2_X1 U4299 ( .A1(n2485), .A2(REG2_REG_21__SCAN_IN), .ZN(n3714) );
  OAI21_X1 U4300 ( .B1(n3721), .B2(n3720), .A(n3719), .ZN(n3725) );
  NAND2_X1 U4301 ( .A1(n5070), .A2(n3924), .ZN(n5079) );
  MUX2_X1 U4302 ( .A(n4789), .B(DATAI_15_), .S(n4199), .Z(n5089) );
  NAND2_X1 U4303 ( .A1(n3725), .A2(n3724), .ZN(n3727) );
  INV_X1 U4304 ( .A(n5089), .ZN(n3829) );
  OAI21_X1 U4305 ( .B1(n3728), .B2(REG3_REG_16__SCAN_IN), .A(n3733), .ZN(n5113) );
  INV_X1 U4306 ( .A(n5113), .ZN(n3729) );
  AOI22_X1 U4307 ( .A1(n2487), .A2(n3729), .B1(n4188), .B2(
        REG1_REG_16__SCAN_IN), .ZN(n3731) );
  AOI22_X1 U4308 ( .A1(n2485), .A2(REG2_REG_16__SCAN_IN), .B1(n3858), .B2(
        REG0_REG_16__SCAN_IN), .ZN(n3730) );
  MUX2_X1 U4309 ( .A(n5105), .B(n5104), .S(n4199), .Z(n4555) );
  AOI21_X1 U4310 ( .B1(n3733), .B2(n3732), .A(n3739), .ZN(n5137) );
  NAND2_X1 U4311 ( .A1(n2982), .A2(n5137), .ZN(n3737) );
  NAND2_X1 U4312 ( .A1(n2485), .A2(REG2_REG_17__SCAN_IN), .ZN(n3736) );
  NAND2_X1 U4313 ( .A1(n4188), .A2(REG1_REG_17__SCAN_IN), .ZN(n3735) );
  NAND2_X1 U4314 ( .A1(n3858), .A2(REG0_REG_17__SCAN_IN), .ZN(n3734) );
  NAND4_X1 U4315 ( .A1(n3737), .A2(n3736), .A3(n3735), .A4(n3734), .ZN(n4317)
         );
  MUX2_X1 U4316 ( .A(n4627), .B(DATAI_17_), .S(n4199), .Z(n5127) );
  NOR2_X1 U4317 ( .A1(n4317), .A2(n5127), .ZN(n3738) );
  OAI21_X1 U4318 ( .B1(n3739), .B2(REG3_REG_18__SCAN_IN), .A(n3742), .ZN(n5166) );
  INV_X1 U4319 ( .A(n5166), .ZN(n4540) );
  AOI22_X1 U4320 ( .A1(n2487), .A2(n4540), .B1(n2483), .B2(
        REG1_REG_18__SCAN_IN), .ZN(n3741) );
  AOI22_X1 U4321 ( .A1(n2485), .A2(REG2_REG_18__SCAN_IN), .B1(n3858), .B2(
        REG0_REG_18__SCAN_IN), .ZN(n3740) );
  MUX2_X1 U4322 ( .A(n5154), .B(DATAI_18_), .S(n4199), .Z(n5161) );
  OR2_X1 U4323 ( .A1(n5176), .A2(n5161), .ZN(n5200) );
  NAND2_X1 U4324 ( .A1(n5176), .A2(n5161), .ZN(n4169) );
  INV_X1 U4325 ( .A(n5176), .ZN(n4316) );
  NAND2_X1 U4326 ( .A1(n2485), .A2(REG2_REG_19__SCAN_IN), .ZN(n3748) );
  AND2_X1 U4327 ( .A1(n3742), .A2(n3880), .ZN(n3743) );
  OR2_X1 U4328 ( .A1(n3743), .A2(n3751), .ZN(n5215) );
  INV_X1 U4329 ( .A(n5215), .ZN(n3744) );
  NAND2_X1 U4330 ( .A1(n2982), .A2(n3744), .ZN(n3747) );
  NAND2_X1 U4331 ( .A1(n4188), .A2(REG1_REG_19__SCAN_IN), .ZN(n3746) );
  NAND2_X1 U4332 ( .A1(n3858), .A2(REG0_REG_19__SCAN_IN), .ZN(n3745) );
  NAND4_X1 U4333 ( .A1(n3748), .A2(n3747), .A3(n3746), .A4(n3745), .ZN(n4512)
         );
  INV_X1 U4334 ( .A(n4512), .ZN(n4531) );
  INV_X1 U4335 ( .A(DATAI_19_), .ZN(n3749) );
  MUX2_X1 U4336 ( .A(n4840), .B(n3749), .S(n4199), .Z(n5204) );
  NAND2_X1 U4337 ( .A1(n4531), .A2(n5193), .ZN(n4166) );
  NAND2_X1 U4338 ( .A1(n4512), .A2(n5204), .ZN(n3838) );
  NAND2_X1 U4339 ( .A1(n4166), .A2(n3838), .ZN(n5202) );
  NAND2_X1 U4340 ( .A1(n5199), .A2(n5202), .ZN(n5198) );
  NAND2_X1 U4341 ( .A1(n5198), .A2(n3750), .ZN(n4510) );
  NAND2_X1 U4342 ( .A1(n2485), .A2(REG2_REG_20__SCAN_IN), .ZN(n3757) );
  NOR2_X1 U4343 ( .A1(n3751), .A2(REG3_REG_20__SCAN_IN), .ZN(n3752) );
  NOR2_X1 U4344 ( .A1(n3753), .A2(n3752), .ZN(n4525) );
  NAND2_X1 U4345 ( .A1(n2982), .A2(n4525), .ZN(n3756) );
  NAND2_X1 U4346 ( .A1(n3858), .A2(REG0_REG_20__SCAN_IN), .ZN(n3755) );
  NAND2_X1 U4347 ( .A1(n4188), .A2(REG1_REG_20__SCAN_IN), .ZN(n3754) );
  NAND4_X1 U4348 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n5178)
         );
  NAND2_X1 U4349 ( .A1(n5178), .A2(n3840), .ZN(n3759) );
  NOR2_X1 U4350 ( .A1(n5178), .A2(n3840), .ZN(n3758) );
  AOI21_X1 U4351 ( .B1(n4510), .B2(n3759), .A(n3758), .ZN(n4497) );
  OAI21_X1 U4352 ( .B1(n4506), .B2(n4520), .A(n4497), .ZN(n3761) );
  NAND2_X1 U4353 ( .A1(n4520), .A2(n4506), .ZN(n3760) );
  NAND2_X1 U4354 ( .A1(n3761), .A2(n3760), .ZN(n4486) );
  INV_X1 U4355 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4492) );
  NAND2_X1 U4356 ( .A1(n2483), .A2(REG1_REG_22__SCAN_IN), .ZN(n3764) );
  NAND2_X1 U4357 ( .A1(n3858), .A2(REG0_REG_22__SCAN_IN), .ZN(n3763) );
  OAI211_X1 U4358 ( .C1(n3762), .C2(n4492), .A(n3764), .B(n3763), .ZN(n3765)
         );
  INV_X1 U4359 ( .A(n3765), .ZN(n3769) );
  OR2_X1 U4360 ( .A1(n3766), .A2(REG3_REG_22__SCAN_IN), .ZN(n3767) );
  AND2_X1 U4361 ( .A1(n3771), .A2(n3767), .ZN(n4490) );
  NAND2_X1 U4362 ( .A1(n4490), .A2(n2982), .ZN(n3768) );
  NAND2_X1 U4363 ( .A1(n4071), .A2(n4480), .ZN(n4463) );
  NAND2_X1 U4364 ( .A1(n4315), .A2(n4489), .ZN(n3842) );
  INV_X1 U4365 ( .A(n4485), .ZN(n4407) );
  NAND2_X1 U4366 ( .A1(n3771), .A2(n3770), .ZN(n3772) );
  AND2_X1 U4367 ( .A1(n3782), .A2(n3772), .ZN(n4469) );
  NAND2_X1 U4368 ( .A1(n4469), .A2(n2982), .ZN(n3777) );
  INV_X1 U4369 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4471) );
  NAND2_X1 U4370 ( .A1(n2983), .A2(REG1_REG_23__SCAN_IN), .ZN(n3774) );
  NAND2_X1 U4371 ( .A1(n3858), .A2(REG0_REG_23__SCAN_IN), .ZN(n3773) );
  OAI211_X1 U4372 ( .C1(n3762), .C2(n4471), .A(n3774), .B(n3773), .ZN(n3775)
         );
  INV_X1 U4373 ( .A(n3775), .ZN(n3776) );
  NAND2_X1 U4374 ( .A1(n4314), .A2(n4475), .ZN(n3780) );
  INV_X1 U4375 ( .A(n3780), .ZN(n3778) );
  NOR2_X1 U4376 ( .A1(n4482), .A2(n4475), .ZN(n3845) );
  AND2_X1 U4377 ( .A1(n4407), .A2(n4408), .ZN(n3779) );
  INV_X1 U4378 ( .A(n4408), .ZN(n3781) );
  NAND2_X1 U4379 ( .A1(n4315), .A2(n4480), .ZN(n4458) );
  AND2_X1 U4380 ( .A1(n4458), .A2(n3780), .ZN(n4409) );
  OR2_X1 U4381 ( .A1(n3781), .A2(n4409), .ZN(n3792) );
  NAND2_X1 U4382 ( .A1(n3782), .A2(n4095), .ZN(n3784) );
  INV_X1 U4383 ( .A(n3793), .ZN(n3783) );
  NAND2_X1 U4384 ( .A1(n3784), .A2(n3783), .ZN(n4445) );
  OR2_X1 U4385 ( .A1(n4445), .A2(n3785), .ZN(n3790) );
  INV_X1 U4386 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4446) );
  NAND2_X1 U4387 ( .A1(n2483), .A2(REG1_REG_24__SCAN_IN), .ZN(n3787) );
  NAND2_X1 U4388 ( .A1(n3858), .A2(REG0_REG_24__SCAN_IN), .ZN(n3786) );
  OAI211_X1 U4389 ( .C1(n3762), .C2(n4446), .A(n3787), .B(n3786), .ZN(n3788)
         );
  INV_X1 U4390 ( .A(n3788), .ZN(n3789) );
  INV_X1 U4391 ( .A(n4450), .ZN(n3791) );
  NAND2_X1 U4392 ( .A1(n2483), .A2(REG1_REG_25__SCAN_IN), .ZN(n3797) );
  NAND2_X1 U4393 ( .A1(REG3_REG_25__SCAN_IN), .A2(n3793), .ZN(n3800) );
  OAI21_X1 U4394 ( .B1(REG3_REG_25__SCAN_IN), .B2(n3793), .A(n3800), .ZN(n4437) );
  INV_X1 U4395 ( .A(n4437), .ZN(n4083) );
  NAND2_X1 U4396 ( .A1(n2487), .A2(n4083), .ZN(n3796) );
  NAND2_X1 U4397 ( .A1(n2485), .A2(REG2_REG_25__SCAN_IN), .ZN(n3795) );
  NAND2_X1 U4398 ( .A1(n3858), .A2(REG0_REG_25__SCAN_IN), .ZN(n3794) );
  NAND2_X1 U4399 ( .A1(n4097), .A2(n4424), .ZN(n4402) );
  NAND2_X1 U4400 ( .A1(n4453), .A2(n4436), .ZN(n4180) );
  NAND2_X1 U4401 ( .A1(n2483), .A2(REG1_REG_26__SCAN_IN), .ZN(n3805) );
  INV_X1 U4402 ( .A(n3800), .ZN(n3798) );
  NAND2_X1 U4403 ( .A1(n3798), .A2(REG3_REG_26__SCAN_IN), .ZN(n3812) );
  INV_X1 U4404 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3799) );
  NAND2_X1 U4405 ( .A1(n3800), .A2(n3799), .ZN(n3801) );
  AND2_X1 U4406 ( .A1(n3812), .A2(n3801), .ZN(n4416) );
  NAND2_X1 U4407 ( .A1(n2487), .A2(n4416), .ZN(n3804) );
  NAND2_X1 U4408 ( .A1(n2485), .A2(REG2_REG_26__SCAN_IN), .ZN(n3803) );
  NAND2_X1 U4409 ( .A1(n3858), .A2(REG0_REG_26__SCAN_IN), .ZN(n3802) );
  AND2_X1 U4410 ( .A1(n4386), .A2(n4415), .ZN(n3809) );
  OR2_X1 U4411 ( .A1(n4433), .A2(n3809), .ZN(n3806) );
  OR2_X1 U4412 ( .A1(n4386), .A2(n4415), .ZN(n3807) );
  NAND2_X1 U4413 ( .A1(n4453), .A2(n4424), .ZN(n4411) );
  AND2_X1 U4414 ( .A1(n3807), .A2(n4411), .ZN(n3808) );
  NOR2_X1 U4415 ( .A1(n3809), .A2(n3808), .ZN(n3810) );
  INV_X1 U4416 ( .A(n3812), .ZN(n3811) );
  NAND2_X1 U4417 ( .A1(n3811), .A2(REG3_REG_27__SCAN_IN), .ZN(n3820) );
  NAND2_X1 U4418 ( .A1(n3812), .A2(n4033), .ZN(n3813) );
  NAND2_X1 U4419 ( .A1(n2487), .A2(n4392), .ZN(n3817) );
  NAND2_X1 U4420 ( .A1(n2483), .A2(REG1_REG_27__SCAN_IN), .ZN(n3816) );
  NAND2_X1 U4421 ( .A1(n2485), .A2(REG2_REG_27__SCAN_IN), .ZN(n3815) );
  NAND2_X1 U4422 ( .A1(n3858), .A2(REG0_REG_27__SCAN_IN), .ZN(n3814) );
  NAND4_X1 U4423 ( .A1(n3817), .A2(n3816), .A3(n3815), .A4(n3814), .ZN(n4313)
         );
  NOR2_X1 U4424 ( .A1(n4313), .A2(n4396), .ZN(n3818) );
  INV_X1 U4425 ( .A(n4396), .ZN(n4034) );
  OAI22_X1 U4426 ( .A1(n4381), .A2(n3818), .B1(n4025), .B2(n4034), .ZN(n4354)
         );
  INV_X1 U4427 ( .A(n3820), .ZN(n3819) );
  NAND2_X1 U4428 ( .A1(n3819), .A2(REG3_REG_28__SCAN_IN), .ZN(n3857) );
  NAND2_X1 U4429 ( .A1(n3820), .A2(n4022), .ZN(n3821) );
  NAND2_X1 U4430 ( .A1(n2487), .A2(n4023), .ZN(n3825) );
  NAND2_X1 U4431 ( .A1(n2483), .A2(REG1_REG_28__SCAN_IN), .ZN(n3824) );
  NAND2_X1 U4432 ( .A1(n2485), .A2(REG2_REG_28__SCAN_IN), .ZN(n3823) );
  NAND2_X1 U4433 ( .A1(n3858), .A2(REG0_REG_28__SCAN_IN), .ZN(n3822) );
  NAND2_X1 U4434 ( .A1(n4389), .A2(n3827), .ZN(n4360) );
  INV_X1 U4435 ( .A(n4389), .ZN(n4312) );
  NAND2_X1 U4436 ( .A1(n4312), .A2(n4355), .ZN(n4184) );
  XNOR2_X1 U4437 ( .A(n4354), .B(n4353), .ZN(n4573) );
  NAND2_X1 U4438 ( .A1(n5140), .A2(n4539), .ZN(n4538) );
  OR2_X2 U4439 ( .A1(n4538), .A2(n5193), .ZN(n5195) );
  NOR2_X2 U4440 ( .A1(n5195), .A2(n3840), .ZN(n4498) );
  INV_X1 U4441 ( .A(n4373), .ZN(n4375) );
  OAI211_X1 U4442 ( .C1(n2550), .C2(n4355), .A(n4375), .B(n5249), .ZN(n4571)
         );
  INV_X1 U4443 ( .A(n4571), .ZN(n3828) );
  INV_X1 U4444 ( .A(n3696), .ZN(n3833) );
  NAND2_X1 U4445 ( .A1(n4550), .A2(n5089), .ZN(n3832) );
  AND2_X1 U4446 ( .A1(n5084), .A2(n3832), .ZN(n4255) );
  NAND2_X1 U4447 ( .A1(n4319), .A2(n3829), .ZN(n3830) );
  NAND2_X1 U4448 ( .A1(n3831), .A2(n3830), .ZN(n4282) );
  AND2_X1 U4449 ( .A1(n4282), .A2(n3832), .ZN(n4284) );
  AOI21_X1 U4450 ( .B1(n3833), .B2(n4255), .A(n4284), .ZN(n4176) );
  INV_X1 U4451 ( .A(n4176), .ZN(n4548) );
  XNOR2_X1 U4452 ( .A(n4318), .B(n5109), .ZN(n4547) );
  NAND2_X1 U4453 ( .A1(n4548), .A2(n4547), .ZN(n3834) );
  NAND2_X1 U4454 ( .A1(n4318), .A2(n4555), .ZN(n4173) );
  NAND2_X1 U4455 ( .A1(n3834), .A2(n4173), .ZN(n5132) );
  INV_X1 U4456 ( .A(n5132), .ZN(n3835) );
  NAND2_X1 U4457 ( .A1(n3835), .A2(n2680), .ZN(n3836) );
  NAND2_X1 U4458 ( .A1(n4549), .A2(n5127), .ZN(n4220) );
  NAND2_X1 U4459 ( .A1(n3836), .A2(n4220), .ZN(n4535) );
  INV_X1 U4460 ( .A(n4535), .ZN(n3837) );
  NAND2_X1 U4461 ( .A1(n3837), .A2(n4169), .ZN(n5201) );
  NAND2_X1 U4462 ( .A1(n5200), .A2(n3838), .ZN(n4167) );
  INV_X1 U4463 ( .A(n4167), .ZN(n4175) );
  INV_X1 U4464 ( .A(n4166), .ZN(n3839) );
  AOI21_X2 U4465 ( .B1(n5201), .B2(n4175), .A(n3839), .ZN(n4516) );
  INV_X1 U4466 ( .A(n5178), .ZN(n4070) );
  NAND2_X1 U4467 ( .A1(n4070), .A2(n3840), .ZN(n4165) );
  NAND2_X1 U4468 ( .A1(n5178), .A2(n4522), .ZN(n4174) );
  NAND2_X1 U4469 ( .A1(n4516), .A2(n4515), .ZN(n4514) );
  NAND2_X1 U4470 ( .A1(n4514), .A2(n4174), .ZN(n4461) );
  OR2_X1 U4471 ( .A1(n4520), .A2(n3970), .ZN(n4215) );
  NAND2_X1 U4472 ( .A1(n4463), .A2(n4215), .ZN(n4170) );
  INV_X1 U4473 ( .A(n4170), .ZN(n3841) );
  NAND2_X1 U4474 ( .A1(n4461), .A2(n3841), .ZN(n3847) );
  AND2_X1 U4475 ( .A1(n4520), .A2(n3970), .ZN(n4462) );
  NAND2_X1 U4476 ( .A1(n4463), .A2(n4462), .ZN(n3843) );
  NAND2_X1 U4477 ( .A1(n3843), .A2(n3842), .ZN(n3844) );
  OR2_X1 U4478 ( .A1(n3845), .A2(n3844), .ZN(n4291) );
  INV_X1 U4479 ( .A(n4291), .ZN(n3846) );
  NAND2_X1 U4480 ( .A1(n3847), .A2(n3846), .ZN(n3849) );
  INV_X1 U4481 ( .A(n4177), .ZN(n3848) );
  NAND2_X1 U4482 ( .A1(n3849), .A2(n3848), .ZN(n4449) );
  INV_X1 U4483 ( .A(n4178), .ZN(n3850) );
  NAND2_X1 U4484 ( .A1(n4448), .A2(n3850), .ZN(n4423) );
  NAND2_X1 U4485 ( .A1(n4386), .A2(n4161), .ZN(n4210) );
  NAND2_X1 U4486 ( .A1(n4402), .A2(n4210), .ZN(n4295) );
  INV_X1 U4487 ( .A(n4295), .ZN(n3851) );
  NAND2_X1 U4488 ( .A1(n4025), .A2(n4396), .ZN(n4192) );
  NAND2_X1 U4489 ( .A1(n4313), .A2(n4034), .ZN(n4185) );
  INV_X1 U4490 ( .A(n4192), .ZN(n3852) );
  NOR2_X1 U4491 ( .A1(n4385), .A2(n3852), .ZN(n3853) );
  NAND2_X1 U4492 ( .A1(n4313), .A2(n4511), .ZN(n3856) );
  OAI21_X1 U4493 ( .B1(n5237), .B2(n4355), .A(n3856), .ZN(n3864) );
  INV_X1 U4494 ( .A(n3857), .ZN(n4359) );
  NAND2_X1 U4495 ( .A1(n2487), .A2(n4359), .ZN(n3862) );
  NAND2_X1 U4496 ( .A1(n2483), .A2(REG1_REG_29__SCAN_IN), .ZN(n3861) );
  NAND2_X1 U4497 ( .A1(n2485), .A2(REG2_REG_29__SCAN_IN), .ZN(n3860) );
  NAND2_X1 U4498 ( .A1(n3858), .A2(REG0_REG_29__SCAN_IN), .ZN(n3859) );
  AND2_X1 U4499 ( .A1(n4311), .A2(n5177), .ZN(n3863) );
  AOI21_X2 U4500 ( .B1(n3865), .B2(n5207), .A(n2677), .ZN(n4572) );
  NAND2_X1 U4501 ( .A1(n4023), .A2(n5136), .ZN(n3866) );
  AOI21_X1 U4502 ( .B1(n3867), .B2(n2495), .A(n5246), .ZN(n3868) );
  AOI21_X1 U4503 ( .B1(n5246), .B2(REG2_REG_28__SCAN_IN), .A(n3868), .ZN(n3869) );
  OAI21_X1 U4504 ( .B1(n4573), .B2(n5103), .A(n3869), .ZN(U3262) );
  AND2_X1 U4505 ( .A1(n5154), .A2(REG1_REG_18__SCAN_IN), .ZN(n3870) );
  INV_X1 U4506 ( .A(REG1_REG_19__SCAN_IN), .ZN(n5223) );
  MUX2_X1 U4507 ( .A(n5223), .B(REG1_REG_19__SCAN_IN), .S(n4840), .Z(n3872) );
  INV_X1 U4508 ( .A(n3872), .ZN(n3873) );
  XNOR2_X1 U4509 ( .A(n3874), .B(n3873), .ZN(n3886) );
  INV_X1 U4510 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3876) );
  MUX2_X1 U4511 ( .A(n3876), .B(REG2_REG_19__SCAN_IN), .S(n4840), .Z(n3877) );
  NOR2_X1 U4512 ( .A1(STATE_REG_SCAN_IN), .A2(n3880), .ZN(n5189) );
  INV_X1 U4513 ( .A(n5189), .ZN(n3882) );
  NAND2_X1 U4514 ( .A1(n4815), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3881) );
  OAI211_X1 U4515 ( .C1(n4827), .C2(n4840), .A(n3882), .B(n3881), .ZN(n3883)
         );
  AOI21_X1 U4516 ( .B1(n3884), .B2(n4824), .A(n3883), .ZN(n3885) );
  OAI21_X1 U4517 ( .B1(n3886), .B2(n4793), .A(n3885), .ZN(U3259) );
  OAI22_X1 U4518 ( .A1(n3889), .A2(n4015), .B1(n3887), .B2(n2486), .ZN(n3888)
         );
  XNOR2_X1 U4519 ( .A(n3888), .B(n3968), .ZN(n3899) );
  OR2_X1 U4520 ( .A1(n3889), .A2(n2937), .ZN(n3891) );
  NAND2_X1 U4521 ( .A1(n4053), .A2(n3468), .ZN(n3890) );
  NAND2_X1 U4522 ( .A1(n3891), .A2(n3890), .ZN(n3898) );
  XNOR2_X1 U4523 ( .A(n3899), .B(n3898), .ZN(n4050) );
  INV_X1 U4524 ( .A(n3892), .ZN(n3895) );
  INV_X1 U4525 ( .A(n3893), .ZN(n3894) );
  NAND2_X1 U4526 ( .A1(n3895), .A2(n3894), .ZN(n4048) );
  NAND2_X1 U4527 ( .A1(n4323), .A2(n3468), .ZN(n3903) );
  NAND2_X1 U4528 ( .A1(n5006), .A2(n3987), .ZN(n3902) );
  NAND2_X1 U4529 ( .A1(n3903), .A2(n3902), .ZN(n3904) );
  XNOR2_X1 U4530 ( .A(n3904), .B(n3968), .ZN(n3906) );
  AOI22_X1 U4531 ( .A1(n4323), .A2(n4010), .B1(n5006), .B2(n3468), .ZN(n3905)
         );
  NOR2_X1 U4532 ( .A1(n3906), .A2(n3905), .ZN(n4998) );
  AND2_X1 U4533 ( .A1(n3906), .A2(n3905), .ZN(n5004) );
  NAND2_X1 U4534 ( .A1(n4322), .A2(n3468), .ZN(n3908) );
  NAND2_X1 U4535 ( .A1(n5022), .A2(n3987), .ZN(n3907) );
  NAND2_X1 U4536 ( .A1(n3908), .A2(n3907), .ZN(n3909) );
  XNOR2_X1 U4537 ( .A(n3909), .B(n4016), .ZN(n3913) );
  OAI22_X1 U4538 ( .A1(n3911), .A2(n2937), .B1(n4015), .B2(n3910), .ZN(n3912)
         );
  XNOR2_X1 U4539 ( .A(n3913), .B(n3912), .ZN(n5020) );
  OAI21_X1 U4540 ( .B1(n5021), .B2(n5020), .A(n3914), .ZN(n5037) );
  NAND2_X1 U4541 ( .A1(n4321), .A2(n3468), .ZN(n3916) );
  NAND2_X1 U4542 ( .A1(n5039), .A2(n3987), .ZN(n3915) );
  NAND2_X1 U4543 ( .A1(n3916), .A2(n3915), .ZN(n3917) );
  XNOR2_X1 U4544 ( .A(n3917), .B(n4016), .ZN(n3918) );
  AOI22_X1 U4545 ( .A1(n4321), .A2(n4010), .B1(n3468), .B2(n5039), .ZN(n3919)
         );
  XNOR2_X1 U4546 ( .A(n3918), .B(n3919), .ZN(n5038) );
  INV_X1 U4547 ( .A(n3918), .ZN(n3920) );
  NAND2_X1 U4548 ( .A1(n4320), .A2(n3468), .ZN(n3922) );
  NAND2_X1 U4549 ( .A1(n5057), .A2(n3987), .ZN(n3921) );
  NAND2_X1 U4550 ( .A1(n3922), .A2(n3921), .ZN(n3923) );
  XNOR2_X1 U4551 ( .A(n3923), .B(n4016), .ZN(n3926) );
  OAI22_X1 U4552 ( .A1(n5070), .A2(n2937), .B1(n4015), .B2(n3924), .ZN(n3925)
         );
  XNOR2_X1 U4553 ( .A(n3926), .B(n3925), .ZN(n5055) );
  NAND2_X1 U4554 ( .A1(n4319), .A2(n3468), .ZN(n3929) );
  NAND2_X1 U4555 ( .A1(n5089), .A2(n3987), .ZN(n3928) );
  NAND2_X1 U4556 ( .A1(n3929), .A2(n3928), .ZN(n3930) );
  XNOR2_X1 U4557 ( .A(n3930), .B(n4016), .ZN(n5072) );
  NAND2_X1 U4558 ( .A1(n4319), .A2(n4010), .ZN(n3932) );
  NAND2_X1 U4559 ( .A1(n5089), .A2(n3468), .ZN(n3931) );
  NAND2_X1 U4560 ( .A1(n3932), .A2(n3931), .ZN(n3933) );
  NAND2_X1 U4561 ( .A1(n5072), .A2(n3933), .ZN(n3935) );
  INV_X1 U4562 ( .A(n5072), .ZN(n3934) );
  INV_X1 U4563 ( .A(n3933), .ZN(n5071) );
  OAI22_X1 U4564 ( .A1(n5122), .A2(n4015), .B1(n2486), .B2(n4555), .ZN(n3936)
         );
  XNOR2_X1 U4565 ( .A(n3936), .B(n4016), .ZN(n3938) );
  OAI22_X1 U4566 ( .A1(n5122), .A2(n2937), .B1(n4015), .B2(n4555), .ZN(n3937)
         );
  XNOR2_X1 U4567 ( .A(n3938), .B(n3937), .ZN(n5107) );
  NAND2_X1 U4568 ( .A1(n4317), .A2(n3468), .ZN(n3940) );
  NAND2_X1 U4569 ( .A1(n5127), .A2(n3987), .ZN(n3939) );
  NAND2_X1 U4570 ( .A1(n3940), .A2(n3939), .ZN(n3941) );
  XNOR2_X1 U4571 ( .A(n3941), .B(n4016), .ZN(n3942) );
  OAI22_X1 U4572 ( .A1(n4549), .A2(n2937), .B1(n4015), .B2(n5142), .ZN(n3943)
         );
  XOR2_X1 U4573 ( .A(n3942), .B(n3943), .Z(n5125) );
  INV_X1 U4574 ( .A(n3942), .ZN(n3945) );
  INV_X1 U4575 ( .A(n3943), .ZN(n3944) );
  OAI22_X1 U4576 ( .A1(n5176), .A2(n4015), .B1(n4539), .B2(n2880), .ZN(n3946)
         );
  XNOR2_X1 U4577 ( .A(n3946), .B(n3968), .ZN(n3949) );
  OR2_X1 U4578 ( .A1(n5176), .A2(n2937), .ZN(n3948) );
  NAND2_X1 U4579 ( .A1(n5161), .A2(n3468), .ZN(n3947) );
  AND2_X1 U4580 ( .A1(n3948), .A2(n3947), .ZN(n3950) );
  NAND2_X1 U4581 ( .A1(n3950), .A2(n3949), .ZN(n5157) );
  NAND2_X1 U4582 ( .A1(n4512), .A2(n3468), .ZN(n3952) );
  OR2_X1 U4583 ( .A1(n5204), .A2(n2880), .ZN(n3951) );
  NAND2_X1 U4584 ( .A1(n3952), .A2(n3951), .ZN(n3953) );
  XNOR2_X1 U4585 ( .A(n3953), .B(n4016), .ZN(n3957) );
  NAND2_X1 U4586 ( .A1(n4512), .A2(n4010), .ZN(n3955) );
  OR2_X1 U4587 ( .A1(n5204), .A2(n4015), .ZN(n3954) );
  NAND2_X1 U4588 ( .A1(n3955), .A2(n3954), .ZN(n3956) );
  NOR2_X1 U4589 ( .A1(n3957), .A2(n3956), .ZN(n3958) );
  AOI21_X1 U4590 ( .B1(n3957), .B2(n3956), .A(n3958), .ZN(n5183) );
  INV_X1 U4591 ( .A(n3958), .ZN(n3959) );
  NAND2_X1 U4592 ( .A1(n5181), .A2(n3959), .ZN(n4116) );
  NAND2_X1 U4593 ( .A1(n5178), .A2(n3468), .ZN(n3961) );
  OR2_X1 U4594 ( .A1(n4522), .A2(n2486), .ZN(n3960) );
  NAND2_X1 U4595 ( .A1(n3961), .A2(n3960), .ZN(n3962) );
  XNOR2_X1 U4596 ( .A(n3962), .B(n3968), .ZN(n3965) );
  NOR2_X1 U4597 ( .A1(n4522), .A2(n4015), .ZN(n3963) );
  AOI21_X1 U4598 ( .B1(n5178), .B2(n4010), .A(n3963), .ZN(n3964) );
  OR2_X1 U4599 ( .A1(n3965), .A2(n3964), .ZN(n4114) );
  NAND2_X1 U4600 ( .A1(n3965), .A2(n3964), .ZN(n4113) );
  NAND2_X1 U4601 ( .A1(n4520), .A2(n3468), .ZN(n3967) );
  OR2_X1 U4602 ( .A1(n3970), .A2(n2486), .ZN(n3966) );
  NAND2_X1 U4603 ( .A1(n3967), .A2(n3966), .ZN(n3969) );
  XNOR2_X1 U4604 ( .A(n3969), .B(n3968), .ZN(n3973) );
  NOR2_X1 U4605 ( .A1(n3970), .A2(n4015), .ZN(n3971) );
  AOI21_X1 U4606 ( .B1(n4520), .B2(n4010), .A(n3971), .ZN(n3974) );
  AND2_X1 U4607 ( .A1(n3973), .A2(n3974), .ZN(n4122) );
  OAI22_X1 U4608 ( .A1(n4071), .A2(n4015), .B1(n2486), .B2(n4489), .ZN(n3972)
         );
  XNOR2_X1 U4609 ( .A(n3972), .B(n4016), .ZN(n3980) );
  OAI22_X1 U4610 ( .A1(n4071), .A2(n2937), .B1(n4015), .B2(n4489), .ZN(n3979)
         );
  XNOR2_X1 U4611 ( .A(n3980), .B(n3979), .ZN(n4126) );
  INV_X1 U4612 ( .A(n4126), .ZN(n3977) );
  INV_X1 U4613 ( .A(n3973), .ZN(n3976) );
  INV_X1 U4614 ( .A(n3974), .ZN(n3975) );
  NAND2_X1 U4615 ( .A1(n3976), .A2(n3975), .ZN(n4123) );
  AOI22_X1 U4616 ( .A1(n4314), .A2(n3468), .B1(n3987), .B2(n4475), .ZN(n3978)
         );
  XNOR2_X1 U4617 ( .A(n3978), .B(n4016), .ZN(n3983) );
  AOI22_X1 U4618 ( .A1(n4314), .A2(n4010), .B1(n3468), .B2(n4475), .ZN(n3984)
         );
  XNOR2_X1 U4619 ( .A(n3983), .B(n3984), .ZN(n4040) );
  INV_X1 U4620 ( .A(n4040), .ZN(n3981) );
  OR2_X1 U4621 ( .A1(n3980), .A2(n3979), .ZN(n4039) );
  INV_X1 U4622 ( .A(n4410), .ZN(n4427) );
  OAI22_X1 U4623 ( .A1(n4427), .A2(n2937), .B1(n4015), .B2(n4096), .ZN(n4094)
         );
  AND2_X1 U4624 ( .A1(n4042), .A2(n4094), .ZN(n3982) );
  NAND2_X1 U4625 ( .A1(n4043), .A2(n3982), .ZN(n3991) );
  INV_X1 U4626 ( .A(n4094), .ZN(n3989) );
  INV_X1 U4627 ( .A(n3983), .ZN(n3986) );
  INV_X1 U4628 ( .A(n3984), .ZN(n3985) );
  NAND2_X1 U4629 ( .A1(n3986), .A2(n3985), .ZN(n3994) );
  AOI22_X1 U4630 ( .A1(n4410), .A2(n3468), .B1(n3987), .B2(n4452), .ZN(n3988)
         );
  XOR2_X1 U4631 ( .A(n4016), .B(n3988), .Z(n3992) );
  INV_X1 U4632 ( .A(n3992), .ZN(n3995) );
  AND2_X1 U4633 ( .A1(n3994), .A2(n3995), .ZN(n4089) );
  OR2_X1 U4634 ( .A1(n3989), .A2(n4089), .ZN(n3990) );
  AND2_X1 U4635 ( .A1(n4042), .A2(n3992), .ZN(n3993) );
  OR2_X1 U4636 ( .A1(n3995), .A2(n3994), .ZN(n4076) );
  OAI22_X1 U4637 ( .A1(n4097), .A2(n4015), .B1(n2880), .B2(n4436), .ZN(n3996)
         );
  XNOR2_X1 U4638 ( .A(n3996), .B(n4016), .ZN(n4003) );
  OR2_X1 U4639 ( .A1(n4097), .A2(n2937), .ZN(n3998) );
  NAND2_X1 U4640 ( .A1(n4424), .A2(n3468), .ZN(n3997) );
  NAND2_X1 U4641 ( .A1(n3998), .A2(n3997), .ZN(n4002) );
  XNOR2_X1 U4642 ( .A(n4003), .B(n4002), .ZN(n4082) );
  INV_X1 U4643 ( .A(n4082), .ZN(n3999) );
  AND2_X1 U4644 ( .A1(n4076), .A2(n3999), .ZN(n4000) );
  AND2_X1 U4645 ( .A1(n4077), .A2(n4000), .ZN(n4001) );
  NAND2_X1 U4646 ( .A1(n4078), .A2(n4001), .ZN(n4079) );
  OR2_X1 U4647 ( .A1(n4003), .A2(n4002), .ZN(n4004) );
  OAI22_X1 U4648 ( .A1(n4386), .A2(n4015), .B1(n2486), .B2(n4415), .ZN(n4005)
         );
  XNOR2_X1 U4649 ( .A(n4005), .B(n4016), .ZN(n4156) );
  OR2_X1 U4650 ( .A1(n4386), .A2(n2937), .ZN(n4007) );
  NAND2_X1 U4651 ( .A1(n4161), .A2(n3468), .ZN(n4006) );
  NAND2_X1 U4652 ( .A1(n4007), .A2(n4006), .ZN(n4155) );
  NAND2_X1 U4653 ( .A1(n4156), .A2(n4155), .ZN(n4008) );
  AND2_X1 U4654 ( .A1(n4396), .A2(n3468), .ZN(n4009) );
  AOI21_X1 U4655 ( .B1(n4313), .B2(n4010), .A(n4009), .ZN(n4014) );
  OAI22_X1 U4656 ( .A1(n4025), .A2(n4015), .B1(n2880), .B2(n4034), .ZN(n4011)
         );
  XNOR2_X1 U4657 ( .A(n4011), .B(n4016), .ZN(n4012) );
  XOR2_X1 U4658 ( .A(n4014), .B(n4012), .Z(n4031) );
  INV_X1 U4659 ( .A(n4012), .ZN(n4013) );
  OAI22_X1 U4660 ( .A1(n4389), .A2(n4015), .B1(n4355), .B2(n2880), .ZN(n4019)
         );
  OAI22_X1 U4661 ( .A1(n4389), .A2(n2937), .B1(n4355), .B2(n4015), .ZN(n4017)
         );
  XNOR2_X1 U4662 ( .A(n4017), .B(n4016), .ZN(n4018) );
  XOR2_X1 U4663 ( .A(n4019), .B(n4018), .Z(n4020) );
  XNOR2_X1 U4664 ( .A(n4021), .B(n4020), .ZN(n4030) );
  OAI22_X1 U4665 ( .A1(n5185), .A2(n4355), .B1(STATE_REG_SCAN_IN), .B2(n4022), 
        .ZN(n4028) );
  INV_X1 U4666 ( .A(n4023), .ZN(n4024) );
  OAI22_X1 U4667 ( .A1(n4026), .A2(n4025), .B1(n4024), .B2(n5192), .ZN(n4027)
         );
  AOI211_X1 U4668 ( .C1(n4148), .C2(n4311), .A(n4028), .B(n4027), .ZN(n4029)
         );
  OAI21_X1 U4669 ( .B1(n4030), .B2(n5186), .A(n4029), .ZN(U3217) );
  XNOR2_X1 U4670 ( .A(n4032), .B(n4031), .ZN(n4038) );
  AOI22_X1 U4671 ( .A1(n4148), .A2(n4312), .B1(n4160), .B2(n4392), .ZN(n4037)
         );
  OAI22_X1 U4672 ( .A1(n5185), .A2(n4034), .B1(STATE_REG_SCAN_IN), .B2(n4033), 
        .ZN(n4035) );
  AOI21_X1 U4673 ( .B1(n4151), .B2(n4425), .A(n4035), .ZN(n4036) );
  OAI211_X1 U4674 ( .C1(n4038), .C2(n5186), .A(n4037), .B(n4036), .ZN(U3211)
         );
  NAND2_X1 U4675 ( .A1(n4043), .A2(n4039), .ZN(n4041) );
  AOI21_X1 U4676 ( .B1(n4041), .B2(n4040), .A(n5186), .ZN(n4044) );
  NAND2_X1 U4677 ( .A1(n4043), .A2(n4042), .ZN(n4090) );
  NAND2_X1 U4678 ( .A1(n4044), .A2(n4090), .ZN(n4047) );
  OAI22_X1 U4679 ( .A1(n4427), .A2(n5121), .B1(n4071), .B2(n5175), .ZN(n4466)
         );
  AOI22_X1 U4680 ( .A1(n4466), .A2(n5190), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n4046) );
  AOI22_X1 U4681 ( .A1(n5160), .A2(n4475), .B1(n4469), .B2(n4160), .ZN(n4045)
         );
  NAND3_X1 U4682 ( .A1(n4047), .A2(n4046), .A3(n4045), .ZN(U3213) );
  AND2_X1 U4683 ( .A1(n3897), .A2(n4048), .ZN(n4051) );
  OAI211_X1 U4684 ( .C1(n4051), .C2(n4050), .A(n5162), .B(n4049), .ZN(n4057)
         );
  AOI22_X1 U4685 ( .A1(n4148), .A2(n4323), .B1(n4160), .B2(n4052), .ZN(n4056)
         );
  AOI22_X1 U4686 ( .A1(n5160), .A2(n4053), .B1(REG3_REG_10__SCAN_IN), .B2(
        U3149), .ZN(n4055) );
  NAND2_X1 U4687 ( .A1(n4151), .A2(n4325), .ZN(n4054) );
  NAND4_X1 U4688 ( .A1(n4057), .A2(n4056), .A3(n4055), .A4(n4054), .ZN(U3214)
         );
  OAI21_X1 U4689 ( .B1(n4060), .B2(n4059), .A(n4058), .ZN(n4061) );
  NAND2_X1 U4690 ( .A1(n4061), .A2(n5162), .ZN(n4066) );
  NAND2_X1 U4691 ( .A1(n4331), .A2(n5177), .ZN(n4063) );
  NAND2_X1 U4692 ( .A1(n2978), .A2(n4511), .ZN(n4062) );
  NAND2_X1 U4693 ( .A1(n4063), .A2(n4062), .ZN(n4871) );
  AOI22_X1 U4694 ( .A1(n5160), .A2(n4879), .B1(n5190), .B2(n4871), .ZN(n4065)
         );
  MUX2_X1 U4695 ( .A(n5192), .B(STATE_REG_SCAN_IN), .S(REG3_REG_3__SCAN_IN), 
        .Z(n4064) );
  NAND3_X1 U4696 ( .A1(n4066), .A2(n4065), .A3(n4064), .ZN(U3215) );
  INV_X1 U4697 ( .A(n4122), .ZN(n4068) );
  NAND2_X1 U4698 ( .A1(n4068), .A2(n4123), .ZN(n4069) );
  XNOR2_X1 U4699 ( .A(n4067), .B(n4069), .ZN(n4075) );
  OAI22_X1 U4700 ( .A1(n4071), .A2(n5121), .B1(n4070), .B2(n5175), .ZN(n4505)
         );
  AOI22_X1 U4701 ( .A1(n4505), .A2(n5190), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n4074) );
  AOI22_X1 U4702 ( .A1(n5160), .A2(n4506), .B1(n4072), .B2(n4160), .ZN(n4073)
         );
  OAI211_X1 U4703 ( .C1(n4075), .C2(n5186), .A(n4074), .B(n4073), .ZN(U3220)
         );
  AND2_X1 U4704 ( .A1(n4077), .A2(n4076), .ZN(n4091) );
  NAND2_X1 U4705 ( .A1(n4078), .A2(n4091), .ZN(n4081) );
  INV_X1 U4706 ( .A(n4079), .ZN(n4080) );
  AOI21_X1 U4707 ( .B1(n4082), .B2(n4081), .A(n4080), .ZN(n4088) );
  AOI22_X1 U4708 ( .A1(n4148), .A2(n4425), .B1(n4160), .B2(n4083), .ZN(n4087)
         );
  INV_X1 U4709 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4084) );
  OAI22_X1 U4710 ( .A1(n5185), .A2(n4436), .B1(STATE_REG_SCAN_IN), .B2(n4084), 
        .ZN(n4085) );
  AOI21_X1 U4711 ( .B1(n4151), .B2(n4410), .A(n4085), .ZN(n4086) );
  OAI211_X1 U4712 ( .C1(n4088), .C2(n5186), .A(n4087), .B(n4086), .ZN(U3222)
         );
  NAND2_X1 U4713 ( .A1(n4090), .A2(n4089), .ZN(n4092) );
  NAND2_X1 U4714 ( .A1(n4092), .A2(n4091), .ZN(n4093) );
  XOR2_X1 U4715 ( .A(n4094), .B(n4093), .Z(n4102) );
  OAI22_X1 U4716 ( .A1(n5185), .A2(n4096), .B1(STATE_REG_SCAN_IN), .B2(n4095), 
        .ZN(n4100) );
  INV_X1 U4717 ( .A(n4148), .ZN(n4098) );
  OAI22_X1 U4718 ( .A1(n4098), .A2(n4097), .B1(n5192), .B2(n4445), .ZN(n4099)
         );
  AOI211_X1 U4719 ( .C1(n4151), .C2(n4314), .A(n4100), .B(n4099), .ZN(n4101)
         );
  OAI21_X1 U4720 ( .B1(n4102), .B2(n5186), .A(n4101), .ZN(U3226) );
  AND2_X1 U4721 ( .A1(n4058), .A2(n4103), .ZN(n4106) );
  OAI211_X1 U4722 ( .C1(n4106), .C2(n4105), .A(n5162), .B(n4104), .ZN(n4112)
         );
  AOI22_X1 U4723 ( .A1(n4148), .A2(n4330), .B1(n4160), .B2(n4107), .ZN(n4111)
         );
  AOI22_X1 U4724 ( .A1(n5160), .A2(n4108), .B1(REG3_REG_4__SCAN_IN), .B2(U3149), .ZN(n4110) );
  NAND2_X1 U4725 ( .A1(n4151), .A2(n4332), .ZN(n4109) );
  NAND4_X1 U4726 ( .A1(n4112), .A2(n4111), .A3(n4110), .A4(n4109), .ZN(U3227)
         );
  NAND2_X1 U4727 ( .A1(n4114), .A2(n4113), .ZN(n4115) );
  XNOR2_X1 U4728 ( .A(n4116), .B(n4115), .ZN(n4121) );
  AOI22_X1 U4729 ( .A1(n4148), .A2(n4520), .B1(n4160), .B2(n4525), .ZN(n4120)
         );
  INV_X1 U4730 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4117) );
  OAI22_X1 U4731 ( .A1(n5185), .A2(n4522), .B1(STATE_REG_SCAN_IN), .B2(n4117), 
        .ZN(n4118) );
  AOI21_X1 U4732 ( .B1(n4151), .B2(n4512), .A(n4118), .ZN(n4119) );
  OAI211_X1 U4733 ( .C1(n4121), .C2(n5186), .A(n4120), .B(n4119), .ZN(U3230)
         );
  OR2_X1 U4734 ( .A1(n4067), .A2(n4122), .ZN(n4124) );
  NAND2_X1 U4735 ( .A1(n4124), .A2(n4123), .ZN(n4125) );
  XOR2_X1 U4736 ( .A(n4126), .B(n4125), .Z(n4131) );
  AOI22_X1 U4737 ( .A1(n4151), .A2(n4520), .B1(n4490), .B2(n4160), .ZN(n4130)
         );
  INV_X1 U4738 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4127) );
  OAI22_X1 U4739 ( .A1(n5185), .A2(n4489), .B1(STATE_REG_SCAN_IN), .B2(n4127), 
        .ZN(n4128) );
  AOI21_X1 U4740 ( .B1(n4148), .B2(n4314), .A(n4128), .ZN(n4129) );
  OAI211_X1 U4741 ( .C1(n4131), .C2(n5186), .A(n4130), .B(n4129), .ZN(U3232)
         );
  OAI21_X1 U4742 ( .B1(n4134), .B2(n4133), .A(n4132), .ZN(n4135) );
  NAND2_X1 U4743 ( .A1(n4135), .A2(n5162), .ZN(n4140) );
  AOI22_X1 U4744 ( .A1(n5160), .A2(n4137), .B1(REG3_REG_2__SCAN_IN), .B2(n4136), .ZN(n4139) );
  AOI22_X1 U4745 ( .A1(n4151), .A2(n2949), .B1(n4148), .B2(n4332), .ZN(n4138)
         );
  NAND3_X1 U4746 ( .A1(n4140), .A2(n4139), .A3(n4138), .ZN(U3234) );
  INV_X1 U4747 ( .A(n4141), .ZN(n4145) );
  OR2_X1 U4748 ( .A1(n4908), .A2(n4907), .ZN(n4910) );
  NAND2_X1 U4749 ( .A1(n4910), .A2(n4142), .ZN(n4144) );
  OAI21_X1 U4750 ( .B1(n4145), .B2(n4144), .A(n4143), .ZN(n4146) );
  NAND2_X1 U4751 ( .A1(n4146), .A2(n5162), .ZN(n4154) );
  AOI22_X1 U4752 ( .A1(n4148), .A2(n4327), .B1(n4160), .B2(n4147), .ZN(n4153)
         );
  NAND2_X1 U4753 ( .A1(REG3_REG_6__SCAN_IN), .A2(U3149), .ZN(n4708) );
  OAI21_X1 U4754 ( .B1(n5185), .B2(n4149), .A(n4708), .ZN(n4150) );
  AOI21_X1 U4755 ( .B1(n4151), .B2(n4330), .A(n4150), .ZN(n4152) );
  NAND3_X1 U4756 ( .A1(n4154), .A2(n4153), .A3(n4152), .ZN(U3236) );
  XNOR2_X1 U4757 ( .A(n4156), .B(n4155), .ZN(n4157) );
  XNOR2_X1 U4758 ( .A(n4158), .B(n4157), .ZN(n4164) );
  AOI22_X1 U4759 ( .A1(n4453), .A2(n4511), .B1(n5177), .B2(n4313), .ZN(n4404)
         );
  INV_X1 U4760 ( .A(n4404), .ZN(n4159) );
  AOI22_X1 U4761 ( .A1(n4159), .A2(n5190), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n4163) );
  AOI22_X1 U4762 ( .A1(n5160), .A2(n4161), .B1(n4416), .B2(n4160), .ZN(n4162)
         );
  OAI211_X1 U4763 ( .C1(n4164), .C2(n5186), .A(n4163), .B(n4162), .ZN(U3237)
         );
  NAND2_X1 U4764 ( .A1(n4166), .A2(n4165), .ZN(n4172) );
  INV_X1 U4765 ( .A(n4174), .ZN(n4168) );
  AOI211_X1 U4766 ( .C1(n4169), .C2(n4220), .A(n4168), .B(n4167), .ZN(n4171)
         );
  AOI211_X1 U4767 ( .C1(n4174), .C2(n4172), .A(n4171), .B(n4170), .ZN(n4290)
         );
  AND2_X1 U4768 ( .A1(n5122), .A2(n5109), .ZN(n4287) );
  AND4_X1 U4769 ( .A1(n4175), .A2(n4174), .A3(n2680), .A4(n4173), .ZN(n4285)
         );
  OAI21_X1 U4770 ( .B1(n4176), .B2(n4287), .A(n4285), .ZN(n4179) );
  NOR2_X1 U4771 ( .A1(n4178), .A2(n4177), .ZN(n4288) );
  OAI221_X1 U4772 ( .B1(n4291), .B2(n4290), .C1(n4291), .C2(n4179), .A(n4288), 
        .ZN(n4183) );
  INV_X1 U4773 ( .A(n4180), .ZN(n4181) );
  NOR2_X1 U4774 ( .A1(n4182), .A2(n4181), .ZN(n4294) );
  AND2_X1 U4775 ( .A1(n4183), .A2(n4294), .ZN(n4187) );
  NAND2_X1 U4776 ( .A1(n4311), .A2(n4372), .ZN(n4212) );
  NAND2_X1 U4777 ( .A1(n4212), .A2(n4184), .ZN(n4193) );
  INV_X1 U4778 ( .A(n4185), .ZN(n4186) );
  NOR3_X1 U4779 ( .A1(n4193), .A2(n4186), .A3(n4209), .ZN(n4292) );
  OAI21_X1 U4780 ( .B1(n4187), .B2(n4295), .A(n4292), .ZN(n4208) );
  INV_X1 U4781 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4191) );
  NAND2_X1 U4782 ( .A1(n2483), .A2(REG1_REG_31__SCAN_IN), .ZN(n4190) );
  NAND2_X1 U4783 ( .A1(n3858), .A2(REG0_REG_31__SCAN_IN), .ZN(n4189) );
  OAI211_X1 U4784 ( .C1(n3762), .C2(n4191), .A(n4190), .B(n4189), .ZN(n5227)
         );
  INV_X1 U4785 ( .A(n5227), .ZN(n4204) );
  NAND2_X1 U4786 ( .A1(n4360), .A2(n4192), .ZN(n4195) );
  INV_X1 U4787 ( .A(n4193), .ZN(n4194) );
  NAND2_X1 U4788 ( .A1(n4195), .A2(n4194), .ZN(n4203) );
  INV_X1 U4789 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4198) );
  NAND2_X1 U4790 ( .A1(n2483), .A2(REG1_REG_30__SCAN_IN), .ZN(n4197) );
  NAND2_X1 U4791 ( .A1(n3858), .A2(REG0_REG_30__SCAN_IN), .ZN(n4196) );
  OAI211_X1 U4792 ( .C1(n3762), .C2(n4198), .A(n4197), .B(n4196), .ZN(n4369)
         );
  INV_X1 U4793 ( .A(n5240), .ZN(n4200) );
  NAND2_X1 U4794 ( .A1(n4199), .A2(DATAI_31_), .ZN(n5243) );
  NAND2_X1 U4795 ( .A1(n5227), .A2(n5243), .ZN(n4298) );
  OAI21_X1 U4796 ( .B1(n4369), .B2(n4200), .A(n4298), .ZN(n4214) );
  INV_X1 U4797 ( .A(n4214), .ZN(n4202) );
  NAND2_X1 U4798 ( .A1(n4201), .A2(n4374), .ZN(n4213) );
  NAND3_X1 U4799 ( .A1(n4203), .A2(n4202), .A3(n4213), .ZN(n4296) );
  AOI21_X1 U4800 ( .B1(n4204), .B2(n5240), .A(n4296), .ZN(n4207) );
  INV_X1 U4801 ( .A(n5243), .ZN(n4206) );
  INV_X1 U4802 ( .A(n4369), .ZN(n4205) );
  OAI22_X1 U4803 ( .A1(n4205), .A2(n5240), .B1(n5227), .B2(n5243), .ZN(n4297)
         );
  AOI22_X1 U4804 ( .A1(n4208), .A2(n4207), .B1(n4206), .B2(n4297), .ZN(n4245)
         );
  INV_X1 U4805 ( .A(n4209), .ZN(n4211) );
  NAND2_X1 U4806 ( .A1(n4211), .A2(n4210), .ZN(n4412) );
  NAND2_X1 U4807 ( .A1(n4213), .A2(n4212), .ZN(n4363) );
  OR4_X1 U4808 ( .A1(n4412), .A2(n4363), .A3(n4214), .A4(n4297), .ZN(n4218) );
  INV_X1 U4809 ( .A(n4433), .ZN(n4217) );
  INV_X1 U4810 ( .A(n4462), .ZN(n4216) );
  NAND2_X1 U4811 ( .A1(n4216), .A2(n4215), .ZN(n4502) );
  NOR4_X1 U4812 ( .A1(n4218), .A2(n4353), .A3(n4217), .A4(n4502), .ZN(n4223)
         );
  INV_X1 U4813 ( .A(n4219), .ZN(n4870) );
  NAND2_X1 U4814 ( .A1(n2680), .A2(n4220), .ZN(n5138) );
  AND2_X1 U4815 ( .A1(n2951), .A2(n4833), .ZN(n4257) );
  OR2_X1 U4816 ( .A1(n4257), .A2(n4260), .ZN(n4846) );
  NOR4_X1 U4817 ( .A1(n4870), .A2(n5138), .A3(n4846), .A4(n4221), .ZN(n4222)
         );
  NAND4_X1 U4818 ( .A1(n4223), .A2(n4485), .A3(n4532), .A4(n4222), .ZN(n4242)
         );
  NAND3_X1 U4819 ( .A1(n4224), .A2(n4382), .A3(n4515), .ZN(n4226) );
  NOR4_X1 U4820 ( .A1(n4465), .A2(n4226), .A3(n5202), .A4(n4225), .ZN(n4237)
         );
  INV_X1 U4821 ( .A(n4227), .ZN(n4231) );
  AND4_X1 U4822 ( .A1(n4231), .A2(n4230), .A3(n4229), .A4(n4228), .ZN(n4236)
         );
  NOR4_X1 U4823 ( .A1(n2999), .A2(n4234), .A3(n4233), .A4(n4232), .ZN(n4235)
         );
  NAND3_X1 U4824 ( .A1(n4237), .A2(n4236), .A3(n4235), .ZN(n4241) );
  XNOR2_X1 U4825 ( .A(n4319), .B(n5089), .ZN(n5082) );
  XNOR2_X1 U4826 ( .A(n4238), .B(n4969), .ZN(n4967) );
  NAND4_X1 U4827 ( .A1(n4239), .A2(n4450), .A3(n4547), .A4(n4967), .ZN(n4240)
         );
  NOR4_X1 U4828 ( .A1(n4242), .A2(n4241), .A3(n5086), .A4(n4240), .ZN(n4244)
         );
  MUX2_X1 U4829 ( .A(n4245), .B(n4244), .S(n4243), .Z(n4302) );
  INV_X1 U4830 ( .A(n4246), .ZN(n4276) );
  INV_X1 U4831 ( .A(n4247), .ZN(n4250) );
  INV_X1 U4832 ( .A(n4278), .ZN(n4248) );
  NOR4_X1 U4833 ( .A1(n4276), .A2(n4250), .A3(n4249), .A4(n4248), .ZN(n4253)
         );
  INV_X1 U4834 ( .A(n4251), .ZN(n4252) );
  OAI21_X1 U4835 ( .B1(n4253), .B2(n4252), .A(n4279), .ZN(n4256) );
  AND3_X1 U4836 ( .A1(n4256), .A2(n4255), .A3(n4254), .ZN(n4283) );
  AOI21_X1 U4837 ( .B1(n4258), .B2(n2949), .A(n4257), .ZN(n4259) );
  OAI21_X1 U4838 ( .B1(n4625), .B2(n4260), .A(n4259), .ZN(n4262) );
  NAND3_X1 U4839 ( .A1(n4262), .A2(n3000), .A3(n4261), .ZN(n4265) );
  NAND3_X1 U4840 ( .A1(n4265), .A2(n4264), .A3(n4263), .ZN(n4268) );
  NAND3_X1 U4841 ( .A1(n4268), .A2(n4267), .A3(n4266), .ZN(n4271) );
  NAND3_X1 U4842 ( .A1(n4271), .A2(n4270), .A3(n4269), .ZN(n4274) );
  AND3_X1 U4843 ( .A1(n4274), .A2(n4273), .A3(n4272), .ZN(n4277) );
  OAI21_X1 U4844 ( .B1(n4277), .B2(n4276), .A(n4275), .ZN(n4280) );
  NAND3_X1 U4845 ( .A1(n4280), .A2(n4279), .A3(n4278), .ZN(n4281) );
  OAI22_X1 U4846 ( .A1(n4284), .A2(n4283), .B1(n4282), .B2(n4281), .ZN(n4286)
         );
  OAI21_X1 U4847 ( .B1(n4287), .B2(n4286), .A(n4285), .ZN(n4289) );
  OAI221_X1 U4848 ( .B1(n4291), .B2(n4290), .C1(n4291), .C2(n4289), .A(n4288), 
        .ZN(n4293) );
  OAI221_X1 U4849 ( .B1(n4295), .B2(n4294), .C1(n4295), .C2(n4293), .A(n4292), 
        .ZN(n4300) );
  INV_X1 U4850 ( .A(n4296), .ZN(n4299) );
  AOI22_X1 U4851 ( .A1(n4300), .A2(n4299), .B1(n4298), .B2(n4297), .ZN(n4301)
         );
  MUX2_X1 U4852 ( .A(n4302), .B(n4301), .S(n2874), .Z(n4303) );
  XNOR2_X1 U4853 ( .A(n4303), .B(n4626), .ZN(n4310) );
  INV_X1 U4854 ( .A(n4304), .ZN(n4306) );
  NAND2_X1 U4855 ( .A1(n4306), .A2(n4305), .ZN(n4307) );
  OAI211_X1 U4856 ( .C1(n4624), .C2(n4309), .A(n4307), .B(B_REG_SCAN_IN), .ZN(
        n4308) );
  OAI21_X1 U4857 ( .B1(n4310), .B2(n4309), .A(n4308), .ZN(U3239) );
  MUX2_X1 U4858 ( .A(DATAO_REG_31__SCAN_IN), .B(n5227), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4859 ( .A(DATAO_REG_30__SCAN_IN), .B(n4369), .S(n4328), .Z(U3580)
         );
  MUX2_X1 U4860 ( .A(DATAO_REG_29__SCAN_IN), .B(n4311), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4861 ( .A(DATAO_REG_28__SCAN_IN), .B(n4312), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4862 ( .A(DATAO_REG_27__SCAN_IN), .B(n4313), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4863 ( .A(DATAO_REG_26__SCAN_IN), .B(n4425), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4864 ( .A(DATAO_REG_25__SCAN_IN), .B(n4453), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4865 ( .A(DATAO_REG_24__SCAN_IN), .B(n4410), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4866 ( .A(DATAO_REG_23__SCAN_IN), .B(n4314), .S(n4328), .Z(U3573)
         );
  MUX2_X1 U4867 ( .A(DATAO_REG_22__SCAN_IN), .B(n4315), .S(n4328), .Z(U3572)
         );
  MUX2_X1 U4868 ( .A(DATAO_REG_21__SCAN_IN), .B(n4520), .S(n4328), .Z(U3571)
         );
  MUX2_X1 U4869 ( .A(DATAO_REG_20__SCAN_IN), .B(n5178), .S(n4328), .Z(U3570)
         );
  MUX2_X1 U4870 ( .A(DATAO_REG_19__SCAN_IN), .B(n4512), .S(n4328), .Z(U3569)
         );
  MUX2_X1 U4871 ( .A(DATAO_REG_18__SCAN_IN), .B(n4316), .S(n4328), .Z(U3568)
         );
  MUX2_X1 U4872 ( .A(DATAO_REG_17__SCAN_IN), .B(n4317), .S(n4328), .Z(U3567)
         );
  MUX2_X1 U4873 ( .A(DATAO_REG_16__SCAN_IN), .B(n4318), .S(n4328), .Z(U3566)
         );
  MUX2_X1 U4874 ( .A(DATAO_REG_15__SCAN_IN), .B(n4319), .S(n4328), .Z(U3565)
         );
  MUX2_X1 U4875 ( .A(DATAO_REG_14__SCAN_IN), .B(n4320), .S(n4328), .Z(U3564)
         );
  MUX2_X1 U4876 ( .A(DATAO_REG_13__SCAN_IN), .B(n4321), .S(n4328), .Z(U3563)
         );
  MUX2_X1 U4877 ( .A(DATAO_REG_12__SCAN_IN), .B(n4322), .S(n4328), .Z(U3562)
         );
  MUX2_X1 U4878 ( .A(DATAO_REG_11__SCAN_IN), .B(n4323), .S(n4328), .Z(U3561)
         );
  MUX2_X1 U4879 ( .A(DATAO_REG_10__SCAN_IN), .B(n4324), .S(n4328), .Z(U3560)
         );
  MUX2_X1 U4880 ( .A(DATAO_REG_9__SCAN_IN), .B(n4325), .S(U4043), .Z(U3559) );
  MUX2_X1 U4881 ( .A(DATAO_REG_8__SCAN_IN), .B(n4326), .S(n4328), .Z(U3558) );
  MUX2_X1 U4882 ( .A(DATAO_REG_7__SCAN_IN), .B(n4327), .S(n4328), .Z(U3557) );
  MUX2_X1 U4883 ( .A(DATAO_REG_6__SCAN_IN), .B(n4329), .S(n4328), .Z(U3556) );
  MUX2_X1 U4884 ( .A(DATAO_REG_5__SCAN_IN), .B(n4330), .S(U4043), .Z(U3555) );
  MUX2_X1 U4885 ( .A(DATAO_REG_4__SCAN_IN), .B(n4331), .S(U4043), .Z(U3554) );
  MUX2_X1 U4886 ( .A(DATAO_REG_3__SCAN_IN), .B(n4332), .S(U4043), .Z(U3553) );
  MUX2_X1 U4887 ( .A(DATAO_REG_2__SCAN_IN), .B(n2978), .S(U4043), .Z(U3552) );
  MUX2_X1 U4888 ( .A(DATAO_REG_1__SCAN_IN), .B(n2949), .S(U4043), .Z(U3551) );
  MUX2_X1 U4889 ( .A(DATAO_REG_0__SCAN_IN), .B(n2951), .S(U4043), .Z(U3550) );
  OAI21_X1 U4890 ( .B1(n4334), .B2(n5118), .A(n4333), .ZN(n4335) );
  INV_X1 U4891 ( .A(n4335), .ZN(n4342) );
  OAI21_X1 U4892 ( .B1(n4337), .B2(n4553), .A(n4336), .ZN(n4340) );
  AOI22_X1 U4893 ( .A1(n4815), .A2(ADDR_REG_16__SCAN_IN), .B1(
        REG3_REG_16__SCAN_IN), .B2(U3149), .ZN(n4338) );
  OAI21_X1 U4894 ( .B1(n5105), .B2(n4827), .A(n4338), .ZN(n4339) );
  AOI21_X1 U4895 ( .B1(n4340), .B2(n4824), .A(n4339), .ZN(n4341) );
  OAI21_X1 U4896 ( .B1(n4342), .B2(n4793), .A(n4341), .ZN(U3256) );
  XNOR2_X1 U4897 ( .A(n4344), .B(n4343), .ZN(n4352) );
  AOI22_X1 U4898 ( .A1(n4815), .A2(ADDR_REG_17__SCAN_IN), .B1(
        REG3_REG_17__SCAN_IN), .B2(U3149), .ZN(n4345) );
  INV_X1 U4899 ( .A(n4345), .ZN(n4350) );
  AOI211_X1 U4900 ( .C1(n4348), .C2(n4347), .A(n4798), .B(n4346), .ZN(n4349)
         );
  AOI211_X1 U4901 ( .C1(n4804), .C2(n4627), .A(n4350), .B(n4349), .ZN(n4351)
         );
  OAI21_X1 U4902 ( .B1(n4352), .B2(n4793), .A(n4351), .ZN(U3257) );
  NAND2_X1 U4903 ( .A1(n4354), .A2(n4353), .ZN(n4356) );
  NAND2_X1 U4904 ( .A1(n4356), .A2(n2511), .ZN(n4358) );
  XNOR2_X1 U4905 ( .A(n4358), .B(n4357), .ZN(n4562) );
  NAND2_X1 U4906 ( .A1(n4562), .A2(n5144), .ZN(n4380) );
  AOI22_X1 U4907 ( .A1(n5246), .A2(REG2_REG_29__SCAN_IN), .B1(n4359), .B2(
        n5136), .ZN(n4379) );
  INV_X1 U4908 ( .A(n4360), .ZN(n4361) );
  NOR2_X1 U4909 ( .A1(n4362), .A2(n4361), .ZN(n4364) );
  XNOR2_X1 U4910 ( .A(n4364), .B(n4363), .ZN(n4365) );
  NAND2_X1 U4911 ( .A1(n4365), .A2(n5207), .ZN(n4371) );
  INV_X1 U4912 ( .A(B_REG_SCAN_IN), .ZN(n4366) );
  OR2_X1 U4913 ( .A1(n4805), .A2(n4366), .ZN(n4367) );
  AND2_X1 U4914 ( .A1(n5177), .A2(n4367), .ZN(n5226) );
  OAI22_X1 U4915 ( .A1(n4389), .A2(n5175), .B1(n4372), .B2(n5237), .ZN(n4368)
         );
  AOI21_X1 U4916 ( .B1(n5226), .B2(n4369), .A(n4368), .ZN(n4370) );
  NAND2_X1 U4917 ( .A1(n4565), .A2(n4558), .ZN(n4378) );
  NAND2_X1 U4918 ( .A1(n4373), .A2(n4372), .ZN(n5241) );
  AOI21_X1 U4919 ( .B1(n4375), .B2(n4374), .A(n5219), .ZN(n4376) );
  AND2_X1 U4920 ( .A1(n5241), .A2(n4376), .ZN(n4563) );
  NAND2_X1 U4921 ( .A1(n4563), .A2(n4524), .ZN(n4377) );
  NAND4_X1 U4922 ( .A1(n4380), .A2(n4379), .A3(n4378), .A4(n4377), .ZN(U3354)
         );
  XNOR2_X1 U4923 ( .A(n4381), .B(n4382), .ZN(n4578) );
  NOR2_X1 U4924 ( .A1(n4383), .A2(n4382), .ZN(n4384) );
  OR2_X1 U4925 ( .A1(n4385), .A2(n4384), .ZN(n4391) );
  OR2_X1 U4926 ( .A1(n4386), .A2(n5175), .ZN(n4388) );
  NAND2_X1 U4927 ( .A1(n4396), .A2(n5229), .ZN(n4387) );
  OAI211_X1 U4928 ( .C1(n4389), .C2(n5121), .A(n4388), .B(n4387), .ZN(n4390)
         );
  AOI21_X1 U4929 ( .B1(n4391), .B2(n5207), .A(n4390), .ZN(n4577) );
  INV_X1 U4930 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4394) );
  INV_X1 U4931 ( .A(n4392), .ZN(n4393) );
  OAI22_X1 U4932 ( .A1(n4558), .A2(n4394), .B1(n4393), .B2(n5216), .ZN(n4395)
         );
  INV_X1 U4933 ( .A(n4395), .ZN(n4398) );
  NAND2_X1 U4934 ( .A1(n2494), .A2(n4396), .ZN(n4574) );
  NAND3_X1 U4935 ( .A1(n4575), .A2(n5244), .A3(n4574), .ZN(n4397) );
  OAI211_X1 U4936 ( .C1(n4577), .C2(n5246), .A(n4398), .B(n4397), .ZN(n4399)
         );
  INV_X1 U4937 ( .A(n4399), .ZN(n4400) );
  OAI21_X1 U4938 ( .B1(n4578), .B2(n5103), .A(n4400), .ZN(U3263) );
  NAND2_X1 U4939 ( .A1(n4401), .A2(n4402), .ZN(n4403) );
  XOR2_X1 U4940 ( .A(n4412), .B(n4403), .Z(n4406) );
  OAI21_X1 U4941 ( .B1(n4415), .B2(n5237), .A(n4404), .ZN(n4405) );
  AOI21_X1 U4942 ( .B1(n4406), .B2(n5207), .A(n4405), .ZN(n4580) );
  NAND2_X1 U4943 ( .A1(n4486), .A2(n4407), .ZN(n4459) );
  NAND2_X1 U4944 ( .A1(n4579), .A2(n5144), .ZN(n4422) );
  OAI21_X1 U4945 ( .B1(n4434), .B2(n4415), .A(n2494), .ZN(n4582) );
  INV_X1 U4946 ( .A(n4582), .ZN(n4420) );
  INV_X1 U4947 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4418) );
  INV_X1 U4948 ( .A(n4416), .ZN(n4417) );
  OAI22_X1 U4949 ( .A1(n4558), .A2(n4418), .B1(n4417), .B2(n5216), .ZN(n4419)
         );
  AOI21_X1 U4950 ( .B1(n4420), .B2(n5244), .A(n4419), .ZN(n4421) );
  OAI211_X1 U4951 ( .C1(n5246), .C2(n4580), .A(n4422), .B(n4421), .ZN(U3264)
         );
  OAI21_X1 U4952 ( .B1(n4433), .B2(n4423), .A(n4401), .ZN(n4429) );
  AOI22_X1 U4953 ( .A1(n4425), .A2(n5177), .B1(n5229), .B2(n4424), .ZN(n4426)
         );
  OAI21_X1 U4954 ( .B1(n4427), .B2(n5175), .A(n4426), .ZN(n4428) );
  AOI21_X1 U4955 ( .B1(n4429), .B2(n5207), .A(n4428), .ZN(n4584) );
  INV_X1 U4956 ( .A(n4430), .ZN(n4431) );
  AOI21_X1 U4957 ( .B1(n4433), .B2(n4432), .A(n4431), .ZN(n4583) );
  NAND2_X1 U4958 ( .A1(n4583), .A2(n5144), .ZN(n4442) );
  INV_X1 U4959 ( .A(n4434), .ZN(n4435) );
  OAI21_X1 U4960 ( .B1(n4444), .B2(n4436), .A(n4435), .ZN(n4586) );
  INV_X1 U4961 ( .A(n4586), .ZN(n4440) );
  INV_X1 U4962 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4438) );
  OAI22_X1 U4963 ( .A1(n4558), .A2(n4438), .B1(n4437), .B2(n5216), .ZN(n4439)
         );
  AOI21_X1 U4964 ( .B1(n4440), .B2(n5244), .A(n4439), .ZN(n4441) );
  OAI211_X1 U4965 ( .C1(n5246), .C2(n4584), .A(n4442), .B(n4441), .ZN(U3265)
         );
  XOR2_X1 U4966 ( .A(n4450), .B(n4443), .Z(n4590) );
  AOI21_X1 U4967 ( .B1(n4452), .B2(n4473), .A(n4444), .ZN(n4588) );
  OAI22_X1 U4968 ( .A1(n4558), .A2(n4446), .B1(n4445), .B2(n5216), .ZN(n4447)
         );
  AOI21_X1 U4969 ( .B1(n4588), .B2(n5244), .A(n4447), .ZN(n4457) );
  OAI21_X1 U4970 ( .B1(n4450), .B2(n4449), .A(n4448), .ZN(n4451) );
  NAND2_X1 U4971 ( .A1(n4451), .A2(n5207), .ZN(n4455) );
  AOI22_X1 U4972 ( .A1(n4453), .A2(n5177), .B1(n5229), .B2(n4452), .ZN(n4454)
         );
  OAI211_X1 U4973 ( .C1(n4482), .C2(n5175), .A(n4455), .B(n4454), .ZN(n4587)
         );
  NAND2_X1 U4974 ( .A1(n4587), .A2(n4558), .ZN(n4456) );
  OAI211_X1 U4975 ( .C1(n4590), .C2(n5103), .A(n4457), .B(n4456), .ZN(U3266)
         );
  NAND2_X1 U4976 ( .A1(n4459), .A2(n4458), .ZN(n4460) );
  XNOR2_X1 U4977 ( .A(n4460), .B(n4465), .ZN(n4594) );
  INV_X1 U4978 ( .A(n4461), .ZN(n4503) );
  NOR2_X1 U4979 ( .A1(n4503), .A2(n4502), .ZN(n4501) );
  NOR2_X1 U4980 ( .A1(n4501), .A2(n4462), .ZN(n4479) );
  NAND2_X1 U4981 ( .A1(n4485), .A2(n4479), .ZN(n4478) );
  NAND2_X1 U4982 ( .A1(n4463), .A2(n4478), .ZN(n4464) );
  XNOR2_X1 U4983 ( .A(n4465), .B(n4464), .ZN(n4468) );
  AOI21_X1 U4984 ( .B1(n4475), .B2(n5229), .A(n4466), .ZN(n4467) );
  OAI21_X1 U4985 ( .B1(n4468), .B2(n5091), .A(n4467), .ZN(n4591) );
  INV_X1 U4986 ( .A(n4469), .ZN(n4470) );
  OAI22_X1 U4987 ( .A1(n4558), .A2(n4471), .B1(n4470), .B2(n5216), .ZN(n4472)
         );
  AOI21_X1 U4988 ( .B1(n4591), .B2(n4558), .A(n4472), .ZN(n4477) );
  INV_X1 U4989 ( .A(n4473), .ZN(n4474) );
  AOI21_X1 U4990 ( .B1(n4475), .B2(n4488), .A(n4474), .ZN(n4592) );
  NAND2_X1 U4991 ( .A1(n4592), .A2(n5244), .ZN(n4476) );
  OAI211_X1 U4992 ( .C1(n4594), .C2(n5103), .A(n4477), .B(n4476), .ZN(U3267)
         );
  OAI21_X1 U4993 ( .B1(n4479), .B2(n4485), .A(n4478), .ZN(n4484) );
  AOI22_X1 U4994 ( .A1(n4520), .A2(n4511), .B1(n4480), .B2(n5229), .ZN(n4481)
         );
  OAI21_X1 U4995 ( .B1(n4482), .B2(n5121), .A(n4481), .ZN(n4483) );
  AOI21_X1 U4996 ( .B1(n4484), .B2(n5207), .A(n4483), .ZN(n4596) );
  XNOR2_X1 U4997 ( .A(n4486), .B(n4485), .ZN(n4595) );
  NAND2_X1 U4998 ( .A1(n4595), .A2(n5144), .ZN(n4496) );
  OAI21_X1 U4999 ( .B1(n4487), .B2(n4489), .A(n4488), .ZN(n4598) );
  INV_X1 U5000 ( .A(n4598), .ZN(n4494) );
  INV_X1 U5001 ( .A(n4490), .ZN(n4491) );
  OAI22_X1 U5002 ( .A1(n4558), .A2(n4492), .B1(n4491), .B2(n5216), .ZN(n4493)
         );
  AOI21_X1 U5003 ( .B1(n4494), .B2(n5244), .A(n4493), .ZN(n4495) );
  OAI211_X1 U5004 ( .C1(n5246), .C2(n4596), .A(n4496), .B(n4495), .ZN(U3268)
         );
  XNOR2_X1 U5005 ( .A(n4497), .B(n4502), .ZN(n4602) );
  INV_X1 U5006 ( .A(n4498), .ZN(n4521) );
  AOI21_X1 U5007 ( .B1(n4506), .B2(n4521), .A(n4487), .ZN(n4599) );
  INV_X1 U5008 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4500) );
  OAI22_X1 U5009 ( .A1(n4558), .A2(n4500), .B1(n4499), .B2(n5216), .ZN(n4508)
         );
  AOI211_X1 U5010 ( .C1(n4503), .C2(n4502), .A(n5091), .B(n4501), .ZN(n4504)
         );
  AOI211_X1 U5011 ( .C1(n5229), .C2(n4506), .A(n4505), .B(n4504), .ZN(n4601)
         );
  NOR2_X1 U5012 ( .A1(n4601), .A2(n5246), .ZN(n4507) );
  AOI211_X1 U5013 ( .C1(n4599), .C2(n5244), .A(n4508), .B(n4507), .ZN(n4509)
         );
  OAI21_X1 U5014 ( .B1(n4602), .B2(n5103), .A(n4509), .ZN(U3269) );
  XNOR2_X1 U5015 ( .A(n4510), .B(n4515), .ZN(n4605) );
  NAND2_X1 U5016 ( .A1(n4512), .A2(n4511), .ZN(n4513) );
  OAI21_X1 U5017 ( .B1(n5237), .B2(n4522), .A(n4513), .ZN(n4519) );
  OAI211_X1 U5018 ( .C1(n4516), .C2(n4515), .A(n4514), .B(n5207), .ZN(n4517)
         );
  INV_X1 U5019 ( .A(n4517), .ZN(n4518) );
  AOI211_X1 U5020 ( .C1(n5177), .C2(n4520), .A(n4519), .B(n4518), .ZN(n4604)
         );
  INV_X1 U5021 ( .A(n4604), .ZN(n4528) );
  INV_X1 U5022 ( .A(n5195), .ZN(n4523) );
  OAI211_X1 U5023 ( .C1(n4523), .C2(n4522), .A(n4521), .B(n5249), .ZN(n4603)
         );
  INV_X1 U5024 ( .A(n4524), .ZN(n4542) );
  AOI22_X1 U5025 ( .A1(n5246), .A2(REG2_REG_20__SCAN_IN), .B1(n4525), .B2(
        n5136), .ZN(n4526) );
  OAI21_X1 U5026 ( .B1(n4603), .B2(n4542), .A(n4526), .ZN(n4527) );
  AOI21_X1 U5027 ( .B1(n4528), .B2(n4558), .A(n4527), .ZN(n4529) );
  OAI21_X1 U5028 ( .B1(n4605), .B2(n5103), .A(n4529), .ZN(U3270) );
  XOR2_X1 U5029 ( .A(n4532), .B(n4530), .Z(n5170) );
  OAI22_X1 U5030 ( .A1(n4549), .A2(n5175), .B1(n4531), .B2(n5121), .ZN(n5156)
         );
  INV_X1 U5031 ( .A(n4532), .ZN(n4536) );
  INV_X1 U5032 ( .A(n5200), .ZN(n4533) );
  NOR2_X1 U5033 ( .A1(n5201), .A2(n4533), .ZN(n4534) );
  AOI211_X1 U5034 ( .C1(n4536), .C2(n4535), .A(n5091), .B(n4534), .ZN(n4537)
         );
  AOI211_X1 U5035 ( .C1(n5229), .C2(n5161), .A(n5156), .B(n4537), .ZN(n5168)
         );
  INV_X1 U5036 ( .A(n5168), .ZN(n4544) );
  OAI211_X1 U5037 ( .C1(n5140), .C2(n4539), .A(n5249), .B(n4538), .ZN(n5167)
         );
  AOI22_X1 U5038 ( .A1(n5246), .A2(REG2_REG_18__SCAN_IN), .B1(n5136), .B2(
        n4540), .ZN(n4541) );
  OAI21_X1 U5039 ( .B1(n5167), .B2(n4542), .A(n4541), .ZN(n4543) );
  AOI21_X1 U5040 ( .B1(n4544), .B2(n4558), .A(n4543), .ZN(n4545) );
  OAI21_X1 U5041 ( .B1(n5170), .B2(n5103), .A(n4545), .ZN(U3272) );
  XOR2_X1 U5042 ( .A(n4546), .B(n4547), .Z(n5115) );
  XNOR2_X1 U5043 ( .A(n4548), .B(n4547), .ZN(n4552) );
  OAI22_X1 U5044 ( .A1(n4550), .A2(n5175), .B1(n4549), .B2(n5121), .ZN(n5106)
         );
  AOI21_X1 U5045 ( .B1(n5109), .B2(n5229), .A(n5106), .ZN(n4551) );
  OAI21_X1 U5046 ( .B1(n4552), .B2(n5091), .A(n4551), .ZN(n5117) );
  OAI22_X1 U5047 ( .A1(n4558), .A2(n4553), .B1(n5113), .B2(n5216), .ZN(n4557)
         );
  INV_X1 U5048 ( .A(n2545), .ZN(n4554) );
  OAI21_X1 U5049 ( .B1(n2521), .B2(n4555), .A(n4554), .ZN(n5114) );
  NOR2_X1 U5050 ( .A1(n5114), .A2(n5196), .ZN(n4556) );
  AOI211_X1 U5051 ( .C1(n5117), .C2(n4558), .A(n4557), .B(n4556), .ZN(n4559)
         );
  OAI21_X1 U5052 ( .B1(n5115), .B2(n5103), .A(n4559), .ZN(U3274) );
  NOR2_X1 U5053 ( .A1(n4840), .A2(n4624), .ZN(n4560) );
  NAND2_X1 U5054 ( .A1(n2874), .A2(n4560), .ZN(n4861) );
  NAND2_X1 U5055 ( .A1(n4567), .A2(n4566), .ZN(n4569) );
  MUX2_X1 U5056 ( .A(REG1_REG_29__SCAN_IN), .B(n4608), .S(n5253), .Z(U3547) );
  OAI211_X1 U5057 ( .C1(n4573), .C2(n5169), .A(n4572), .B(n4571), .ZN(n4609)
         );
  MUX2_X1 U5058 ( .A(REG1_REG_28__SCAN_IN), .B(n4609), .S(n5253), .Z(U3546) );
  NAND3_X1 U5059 ( .A1(n4575), .A2(n5249), .A3(n4574), .ZN(n4576) );
  OAI211_X1 U5060 ( .C1(n4578), .C2(n5169), .A(n4577), .B(n4576), .ZN(n4610)
         );
  MUX2_X1 U5061 ( .A(REG1_REG_27__SCAN_IN), .B(n4610), .S(n5253), .Z(U3545) );
  NAND2_X1 U5062 ( .A1(n4579), .A2(n5221), .ZN(n4581) );
  OAI211_X1 U5063 ( .C1(n5219), .C2(n4582), .A(n4581), .B(n4580), .ZN(n4611)
         );
  MUX2_X1 U5064 ( .A(REG1_REG_26__SCAN_IN), .B(n4611), .S(n5253), .Z(U3544) );
  NAND2_X1 U5065 ( .A1(n4583), .A2(n5221), .ZN(n4585) );
  OAI211_X1 U5066 ( .C1(n5219), .C2(n4586), .A(n4585), .B(n4584), .ZN(n4612)
         );
  MUX2_X1 U5067 ( .A(REG1_REG_25__SCAN_IN), .B(n4612), .S(n5253), .Z(U3543) );
  AOI21_X1 U5068 ( .B1(n5249), .B2(n4588), .A(n4587), .ZN(n4589) );
  OAI21_X1 U5069 ( .B1(n4590), .B2(n5169), .A(n4589), .ZN(n4613) );
  MUX2_X1 U5070 ( .A(REG1_REG_24__SCAN_IN), .B(n4613), .S(n5253), .Z(U3542) );
  AOI21_X1 U5071 ( .B1(n4592), .B2(n5249), .A(n4591), .ZN(n4593) );
  OAI21_X1 U5072 ( .B1(n4594), .B2(n5169), .A(n4593), .ZN(n4614) );
  MUX2_X1 U5073 ( .A(REG1_REG_23__SCAN_IN), .B(n4614), .S(n5253), .Z(U3541) );
  NAND2_X1 U5074 ( .A1(n4595), .A2(n5221), .ZN(n4597) );
  OAI211_X1 U5075 ( .C1(n5219), .C2(n4598), .A(n4597), .B(n4596), .ZN(n4615)
         );
  MUX2_X1 U5076 ( .A(REG1_REG_22__SCAN_IN), .B(n4615), .S(n5253), .Z(U3540) );
  NAND2_X1 U5077 ( .A1(n4599), .A2(n5249), .ZN(n4600) );
  OAI211_X1 U5078 ( .C1(n4602), .C2(n5169), .A(n4601), .B(n4600), .ZN(n4616)
         );
  MUX2_X1 U5079 ( .A(REG1_REG_21__SCAN_IN), .B(n4616), .S(n5253), .Z(U3539) );
  OAI211_X1 U5080 ( .C1(n4605), .C2(n5169), .A(n4604), .B(n4603), .ZN(n4617)
         );
  MUX2_X1 U5081 ( .A(REG1_REG_20__SCAN_IN), .B(n4617), .S(n5253), .Z(U3538) );
  MUX2_X1 U5082 ( .A(REG0_REG_28__SCAN_IN), .B(n4609), .S(n5257), .Z(U3514) );
  MUX2_X1 U5083 ( .A(REG0_REG_27__SCAN_IN), .B(n4610), .S(n5257), .Z(U3513) );
  MUX2_X1 U5084 ( .A(REG0_REG_26__SCAN_IN), .B(n4611), .S(n5257), .Z(U3512) );
  MUX2_X1 U5085 ( .A(REG0_REG_25__SCAN_IN), .B(n4612), .S(n5257), .Z(U3511) );
  MUX2_X1 U5086 ( .A(REG0_REG_24__SCAN_IN), .B(n4613), .S(n5257), .Z(U3510) );
  MUX2_X1 U5087 ( .A(REG0_REG_23__SCAN_IN), .B(n4614), .S(n5257), .Z(U3509) );
  MUX2_X1 U5088 ( .A(REG0_REG_22__SCAN_IN), .B(n4615), .S(n5257), .Z(U3508) );
  MUX2_X1 U5089 ( .A(REG0_REG_21__SCAN_IN), .B(n4616), .S(n5257), .Z(U3507) );
  MUX2_X1 U5090 ( .A(REG0_REG_20__SCAN_IN), .B(n4617), .S(n5257), .Z(U3506) );
  MUX2_X1 U5091 ( .A(n4618), .B(D_REG_1__SCAN_IN), .S(n4652), .Z(U3459) );
  NOR3_X1 U5092 ( .A1(n2865), .A2(IR_REG_30__SCAN_IN), .A3(n2765), .ZN(n4619)
         );
  MUX2_X1 U5093 ( .A(DATAI_31_), .B(n4619), .S(STATE_REG_SCAN_IN), .Z(U3321)
         );
  MUX2_X1 U5094 ( .A(DATAI_30_), .B(n4620), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U5095 ( .A(n4621), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5096 ( .A(DATAI_26_), .B(n4622), .S(STATE_REG_SCAN_IN), .Z(U3326)
         );
  MUX2_X1 U5097 ( .A(n4623), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U5098 ( .A(n4624), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U5099 ( .A(n4625), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5100 ( .A(DATAI_19_), .B(n4626), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U5101 ( .A(DATAI_17_), .B(n4627), .S(STATE_REG_SCAN_IN), .Z(U3335)
         );
  MUX2_X1 U5102 ( .A(n4789), .B(DATAI_15_), .S(U3149), .Z(U3337) );
  MUX2_X1 U5103 ( .A(DATAI_10_), .B(n4737), .S(STATE_REG_SCAN_IN), .Z(U3342)
         );
  MUX2_X1 U5104 ( .A(DATAI_9_), .B(n4727), .S(STATE_REG_SCAN_IN), .Z(U3343) );
  MUX2_X1 U5105 ( .A(n4685), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5106 ( .A(n4673), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U5107 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(STATE_REG_SCAN_IN), 
        .Z(U3352) );
  INV_X1 U5108 ( .A(DATAI_23_), .ZN(n4629) );
  AOI21_X1 U5109 ( .B1(U3149), .B2(n4629), .A(n4628), .ZN(U3329) );
  AND2_X1 U5110 ( .A1(n4652), .A2(D_REG_2__SCAN_IN), .ZN(U3320) );
  NOR2_X1 U5111 ( .A1(n4656), .A2(n4630), .ZN(U3319) );
  INV_X1 U5112 ( .A(D_REG_4__SCAN_IN), .ZN(n4631) );
  NOR2_X1 U5113 ( .A1(n4656), .A2(n4631), .ZN(U3318) );
  INV_X1 U5114 ( .A(D_REG_5__SCAN_IN), .ZN(n4632) );
  NOR2_X1 U5115 ( .A1(n4656), .A2(n4632), .ZN(U3317) );
  NOR2_X1 U5116 ( .A1(n4656), .A2(n4633), .ZN(U3316) );
  NOR2_X1 U5117 ( .A1(n4656), .A2(n4634), .ZN(U3315) );
  INV_X1 U5118 ( .A(D_REG_8__SCAN_IN), .ZN(n4635) );
  NOR2_X1 U5119 ( .A1(n4656), .A2(n4635), .ZN(U3314) );
  NOR2_X1 U5120 ( .A1(n4656), .A2(n4636), .ZN(U3313) );
  NOR2_X1 U5121 ( .A1(n4656), .A2(n4637), .ZN(U3312) );
  AND2_X1 U5122 ( .A1(n4652), .A2(D_REG_11__SCAN_IN), .ZN(U3311) );
  AND2_X1 U5123 ( .A1(n4652), .A2(D_REG_12__SCAN_IN), .ZN(U3310) );
  AND2_X1 U5124 ( .A1(n4652), .A2(D_REG_13__SCAN_IN), .ZN(U3309) );
  INV_X1 U5125 ( .A(D_REG_14__SCAN_IN), .ZN(n4638) );
  NOR2_X1 U5126 ( .A1(n4656), .A2(n4638), .ZN(U3308) );
  NOR2_X1 U5127 ( .A1(n4656), .A2(n4639), .ZN(U3307) );
  INV_X1 U5128 ( .A(D_REG_16__SCAN_IN), .ZN(n4640) );
  NOR2_X1 U5129 ( .A1(n4656), .A2(n4640), .ZN(U3306) );
  NOR2_X1 U5130 ( .A1(n4656), .A2(n4641), .ZN(U3305) );
  NOR2_X1 U5131 ( .A1(n4656), .A2(n4642), .ZN(U3304) );
  INV_X1 U5132 ( .A(D_REG_19__SCAN_IN), .ZN(n4643) );
  NOR2_X1 U5133 ( .A1(n4656), .A2(n4643), .ZN(U3303) );
  INV_X1 U5134 ( .A(D_REG_20__SCAN_IN), .ZN(n4644) );
  NOR2_X1 U5135 ( .A1(n4656), .A2(n4644), .ZN(U3302) );
  NOR2_X1 U5136 ( .A1(n4656), .A2(n4645), .ZN(U3301) );
  NOR2_X1 U5137 ( .A1(n4656), .A2(n4646), .ZN(U3300) );
  NOR2_X1 U5138 ( .A1(n4656), .A2(n4647), .ZN(U3299) );
  NOR2_X1 U5139 ( .A1(n4656), .A2(n4648), .ZN(U3298) );
  NOR2_X1 U5140 ( .A1(n4656), .A2(n4649), .ZN(U3297) );
  INV_X1 U5141 ( .A(D_REG_26__SCAN_IN), .ZN(n4650) );
  NOR2_X1 U5142 ( .A1(n4656), .A2(n4650), .ZN(U3296) );
  NOR2_X1 U5143 ( .A1(n4656), .A2(n4651), .ZN(U3295) );
  AND2_X1 U5144 ( .A1(n4652), .A2(D_REG_28__SCAN_IN), .ZN(U3294) );
  INV_X1 U5145 ( .A(D_REG_29__SCAN_IN), .ZN(n4653) );
  NOR2_X1 U5146 ( .A1(n4656), .A2(n4653), .ZN(U3293) );
  INV_X1 U5147 ( .A(D_REG_30__SCAN_IN), .ZN(n4654) );
  NOR2_X1 U5148 ( .A1(n4656), .A2(n4654), .ZN(U3292) );
  NOR2_X1 U5149 ( .A1(n4656), .A2(n4655), .ZN(U3291) );
  INV_X1 U5150 ( .A(REG3_REG_0__SCAN_IN), .ZN(n4843) );
  INV_X1 U5151 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4849) );
  AOI21_X1 U5152 ( .B1(n4658), .B2(n4849), .A(n4657), .ZN(n4812) );
  OAI21_X1 U5153 ( .B1(n4658), .B2(REG1_REG_0__SCAN_IN), .A(n4812), .ZN(n4659)
         );
  XNOR2_X1 U5154 ( .A(n4659), .B(IR_REG_0__SCAN_IN), .ZN(n4661) );
  AOI22_X1 U5155 ( .A1(n4661), .A2(n4660), .B1(n4815), .B2(ADDR_REG_0__SCAN_IN), .ZN(n4662) );
  OAI21_X1 U5156 ( .B1(STATE_REG_SCAN_IN), .B2(n4843), .A(n4662), .ZN(U3240)
         );
  AOI22_X1 U5157 ( .A1(ADDR_REG_1__SCAN_IN), .A2(n4815), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4675) );
  OAI211_X1 U5158 ( .C1(n4807), .C2(n4664), .A(n4824), .B(n4663), .ZN(n4665)
         );
  INV_X1 U5159 ( .A(n4665), .ZN(n4672) );
  INV_X1 U5160 ( .A(n4666), .ZN(n4669) );
  INV_X1 U5161 ( .A(n4667), .ZN(n4668) );
  AOI211_X1 U5162 ( .C1(n4670), .C2(n4669), .A(n4668), .B(n4793), .ZN(n4671)
         );
  AOI211_X1 U5163 ( .C1(n4804), .C2(n4673), .A(n4672), .B(n4671), .ZN(n4674)
         );
  NAND2_X1 U5164 ( .A1(n4675), .A2(n4674), .ZN(U3241) );
  AOI22_X1 U5165 ( .A1(REG3_REG_3__SCAN_IN), .A2(U3149), .B1(n4815), .B2(
        ADDR_REG_3__SCAN_IN), .ZN(n4687) );
  INV_X1 U5166 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4881) );
  INV_X1 U5167 ( .A(n4676), .ZN(n4678) );
  AOI211_X1 U5168 ( .C1(n4881), .C2(n4678), .A(n4677), .B(n4793), .ZN(n4684)
         );
  INV_X1 U5169 ( .A(REG2_REG_3__SCAN_IN), .ZN(n4682) );
  INV_X1 U5170 ( .A(n4679), .ZN(n4681) );
  AOI211_X1 U5171 ( .C1(n4682), .C2(n4681), .A(n4680), .B(n4798), .ZN(n4683)
         );
  AOI211_X1 U5172 ( .C1(n4804), .C2(n4685), .A(n4684), .B(n4683), .ZN(n4686)
         );
  NAND2_X1 U5173 ( .A1(n4687), .A2(n4686), .ZN(U3243) );
  AOI211_X1 U5174 ( .C1(n2530), .C2(n4689), .A(n4688), .B(n4793), .ZN(n4690)
         );
  AND2_X1 U5175 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n4903) );
  AOI211_X1 U5176 ( .C1(n4815), .C2(ADDR_REG_5__SCAN_IN), .A(n4690), .B(n4903), 
        .ZN(n4696) );
  AOI211_X1 U5177 ( .C1(n4693), .C2(n4692), .A(n4691), .B(n4798), .ZN(n4694)
         );
  AOI21_X1 U5178 ( .B1(n4804), .B2(n4901), .A(n4694), .ZN(n4695) );
  NAND2_X1 U5179 ( .A1(n4696), .A2(n4695), .ZN(U3245) );
  NAND2_X1 U5180 ( .A1(ADDR_REG_6__SCAN_IN), .A2(n4815), .ZN(n4710) );
  INV_X1 U5181 ( .A(n4793), .ZN(n4819) );
  AOI21_X1 U5182 ( .B1(n4698), .B2(n4929), .A(n4697), .ZN(n4699) );
  NAND2_X1 U5183 ( .A1(n4819), .A2(n4699), .ZN(n4705) );
  AOI21_X1 U5184 ( .B1(n4702), .B2(n4701), .A(n4700), .ZN(n4703) );
  NAND2_X1 U5185 ( .A1(n4824), .A2(n4703), .ZN(n4704) );
  OAI211_X1 U5186 ( .C1(n4827), .C2(n4706), .A(n4705), .B(n4704), .ZN(n4707)
         );
  INV_X1 U5187 ( .A(n4707), .ZN(n4709) );
  NAND3_X1 U5188 ( .A1(n4710), .A2(n4709), .A3(n4708), .ZN(U3246) );
  AOI211_X1 U5189 ( .C1(n2527), .C2(n4712), .A(n4711), .B(n4793), .ZN(n4714)
         );
  AOI211_X1 U5190 ( .C1(n4815), .C2(ADDR_REG_7__SCAN_IN), .A(n4714), .B(n4713), 
        .ZN(n4719) );
  AOI211_X1 U5191 ( .C1(n2533), .C2(n4716), .A(n4715), .B(n4798), .ZN(n4717)
         );
  AOI21_X1 U5192 ( .B1(n4804), .B2(n4932), .A(n4717), .ZN(n4718) );
  NAND2_X1 U5193 ( .A1(n4719), .A2(n4718), .ZN(U3247) );
  AOI211_X1 U5194 ( .C1(n2525), .C2(n4721), .A(n4793), .B(n4720), .ZN(n4723)
         );
  AOI211_X1 U5195 ( .C1(n4815), .C2(ADDR_REG_9__SCAN_IN), .A(n4723), .B(n4722), 
        .ZN(n4729) );
  AOI211_X1 U5196 ( .C1(n2526), .C2(n4725), .A(n4798), .B(n4724), .ZN(n4726)
         );
  AOI21_X1 U5197 ( .B1(n4804), .B2(n4727), .A(n4726), .ZN(n4728) );
  NAND2_X1 U5198 ( .A1(n4729), .A2(n4728), .ZN(U3249) );
  AOI22_X1 U5199 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .B1(n4815), .B2(
        ADDR_REG_10__SCAN_IN), .ZN(n4739) );
  AOI211_X1 U5200 ( .C1(n4732), .C2(n4731), .A(n4798), .B(n4730), .ZN(n4736)
         );
  AOI211_X1 U5201 ( .C1(n4992), .C2(n4734), .A(n4793), .B(n4733), .ZN(n4735)
         );
  AOI211_X1 U5202 ( .C1(n4804), .C2(n4737), .A(n4736), .B(n4735), .ZN(n4738)
         );
  NAND2_X1 U5203 ( .A1(n4739), .A2(n4738), .ZN(U3250) );
  AOI22_X1 U5204 ( .A1(REG3_REG_11__SCAN_IN), .A2(U3149), .B1(n4815), .B2(
        ADDR_REG_11__SCAN_IN), .ZN(n4749) );
  AOI211_X1 U5205 ( .C1(n4742), .C2(n4741), .A(n4740), .B(n4798), .ZN(n4747)
         );
  AOI211_X1 U5206 ( .C1(n4745), .C2(n4744), .A(n4743), .B(n4793), .ZN(n4746)
         );
  AOI211_X1 U5207 ( .C1(n4804), .C2(n4995), .A(n4747), .B(n4746), .ZN(n4748)
         );
  NAND2_X1 U5208 ( .A1(n4749), .A2(n4748), .ZN(U3251) );
  AOI22_X1 U5209 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .B1(n4815), .B2(
        ADDR_REG_12__SCAN_IN), .ZN(n4760) );
  AOI21_X1 U5210 ( .B1(n4751), .B2(n5031), .A(n4750), .ZN(n4752) );
  NAND2_X1 U5211 ( .A1(n4819), .A2(n4752), .ZN(n4757) );
  AOI21_X1 U5212 ( .B1(n4754), .B2(n3659), .A(n4753), .ZN(n4755) );
  NAND2_X1 U5213 ( .A1(n4824), .A2(n4755), .ZN(n4756) );
  OAI211_X1 U5214 ( .C1(n4827), .C2(n2818), .A(n4757), .B(n4756), .ZN(n4758)
         );
  INV_X1 U5215 ( .A(n4758), .ZN(n4759) );
  NAND2_X1 U5216 ( .A1(n4760), .A2(n4759), .ZN(U3252) );
  AOI22_X1 U5217 ( .A1(REG3_REG_13__SCAN_IN), .A2(U3149), .B1(n4815), .B2(
        ADDR_REG_13__SCAN_IN), .ZN(n4768) );
  AOI211_X1 U5218 ( .C1(n4761), .C2(n4762), .A(n2518), .B(n4798), .ZN(n4766)
         );
  AOI211_X1 U5219 ( .C1(n2512), .C2(n4764), .A(n4763), .B(n4793), .ZN(n4765)
         );
  AOI211_X1 U5220 ( .C1(n4804), .C2(n5034), .A(n4766), .B(n4765), .ZN(n4767)
         );
  NAND2_X1 U5221 ( .A1(n4768), .A2(n4767), .ZN(U3253) );
  AOI22_X1 U5222 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .B1(n4815), .B2(
        ADDR_REG_14__SCAN_IN), .ZN(n4780) );
  AOI21_X1 U5223 ( .B1(n4770), .B2(n5067), .A(n4769), .ZN(n4771) );
  NAND2_X1 U5224 ( .A1(n4819), .A2(n4771), .ZN(n4777) );
  AOI21_X1 U5225 ( .B1(n4774), .B2(n4773), .A(n4772), .ZN(n4775) );
  NAND2_X1 U5226 ( .A1(n4824), .A2(n4775), .ZN(n4776) );
  OAI211_X1 U5227 ( .C1(n4827), .C2(n5052), .A(n4777), .B(n4776), .ZN(n4778)
         );
  INV_X1 U5228 ( .A(n4778), .ZN(n4779) );
  NAND2_X1 U5229 ( .A1(n4780), .A2(n4779), .ZN(U3254) );
  AOI22_X1 U5230 ( .A1(REG3_REG_15__SCAN_IN), .A2(U3149), .B1(n4815), .B2(
        ADDR_REG_15__SCAN_IN), .ZN(n4791) );
  AOI211_X1 U5231 ( .C1(n4781), .C2(n4782), .A(n4798), .B(n2498), .ZN(n4788)
         );
  INV_X1 U5232 ( .A(n4783), .ZN(n4784) );
  AOI211_X1 U5233 ( .C1(n4786), .C2(n4785), .A(n4793), .B(n4784), .ZN(n4787)
         );
  AOI211_X1 U5234 ( .C1(n4804), .C2(n4789), .A(n4788), .B(n4787), .ZN(n4790)
         );
  NAND2_X1 U5235 ( .A1(n4791), .A2(n4790), .ZN(U3255) );
  AOI22_X1 U5236 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4815), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4814) );
  INV_X1 U5237 ( .A(n4792), .ZN(n4794) );
  AOI211_X1 U5238 ( .C1(n4796), .C2(n4795), .A(n4794), .B(n4793), .ZN(n4803)
         );
  INV_X1 U5239 ( .A(n4797), .ZN(n4799) );
  AOI211_X1 U5240 ( .C1(n4801), .C2(n4800), .A(n4799), .B(n4798), .ZN(n4802)
         );
  AOI211_X1 U5241 ( .C1(n4804), .C2(n4858), .A(n4803), .B(n4802), .ZN(n4813)
         );
  MUX2_X1 U5242 ( .A(n4807), .B(n4806), .S(n4805), .Z(n4809) );
  NAND2_X1 U5243 ( .A1(n4809), .A2(n4808), .ZN(n4811) );
  OAI211_X1 U5244 ( .C1(IR_REG_0__SCAN_IN), .C2(n4812), .A(n4811), .B(U4043), 
        .ZN(n4829) );
  NAND3_X1 U5245 ( .A1(n4814), .A2(n4813), .A3(n4829), .ZN(U3242) );
  AOI22_X1 U5246 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .B1(n4815), .B2(
        ADDR_REG_4__SCAN_IN), .ZN(n4831) );
  AOI21_X1 U5247 ( .B1(n4817), .B2(n4898), .A(n4816), .ZN(n4818) );
  NAND2_X1 U5248 ( .A1(n4819), .A2(n4818), .ZN(n4826) );
  AOI21_X1 U5249 ( .B1(n4822), .B2(n4821), .A(n4820), .ZN(n4823) );
  NAND2_X1 U5250 ( .A1(n4824), .A2(n4823), .ZN(n4825) );
  OAI211_X1 U5251 ( .C1(n4827), .C2(n4892), .A(n4826), .B(n4825), .ZN(n4828)
         );
  INV_X1 U5252 ( .A(n4828), .ZN(n4830) );
  NAND3_X1 U5253 ( .A1(n4831), .A2(n4830), .A3(n4829), .ZN(U3244) );
  INV_X1 U5254 ( .A(n4861), .ZN(n4896) );
  NOR2_X1 U5255 ( .A1(n4833), .A2(n4832), .ZN(n4839) );
  OAI21_X1 U5256 ( .B1(n4875), .B2(n5207), .A(n4846), .ZN(n4834) );
  OAI21_X1 U5257 ( .B1(n4835), .B2(n5121), .A(n4834), .ZN(n4844) );
  AOI211_X1 U5258 ( .C1(n4896), .C2(n4846), .A(n4839), .B(n4844), .ZN(n4838)
         );
  INV_X1 U5259 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4836) );
  AOI22_X1 U5260 ( .A1(n5253), .A2(n4838), .B1(n4836), .B2(n5251), .ZN(U3518)
         );
  INV_X1 U5261 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4837) );
  AOI22_X1 U5262 ( .A1(n5257), .A2(n4838), .B1(n4837), .B2(n5254), .ZN(U3467)
         );
  OAI21_X1 U5263 ( .B1(n4841), .B2(n4840), .A(n4839), .ZN(n4842) );
  OAI21_X1 U5264 ( .B1(n5216), .B2(n4843), .A(n4842), .ZN(n4845) );
  AOI211_X1 U5265 ( .C1(n4847), .C2(n4846), .A(n4845), .B(n4844), .ZN(n4848)
         );
  AOI22_X1 U5266 ( .A1(n5246), .A2(n4849), .B1(n4848), .B2(n4558), .ZN(U3290)
         );
  NOR3_X1 U5267 ( .A1(n4850), .A2(n3012), .A3(n5219), .ZN(n4853) );
  INV_X1 U5268 ( .A(n4851), .ZN(n4852) );
  AOI211_X1 U5269 ( .C1(n4854), .C2(n4896), .A(n4853), .B(n4852), .ZN(n4857)
         );
  INV_X1 U5270 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4855) );
  AOI22_X1 U5271 ( .A1(n5253), .A2(n4857), .B1(n4855), .B2(n5251), .ZN(U3519)
         );
  INV_X1 U5272 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4856) );
  AOI22_X1 U5273 ( .A1(n5257), .A2(n4857), .B1(n4856), .B2(n5254), .ZN(U3469)
         );
  OAI22_X1 U5274 ( .A1(U3149), .A2(n4858), .B1(DATAI_2_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4859) );
  INV_X1 U5275 ( .A(n4859), .ZN(U3350) );
  OAI22_X1 U5276 ( .A1(n4862), .A2(n4861), .B1(n5219), .B2(n4860), .ZN(n4864)
         );
  NOR2_X1 U5277 ( .A1(n4864), .A2(n4863), .ZN(n4867) );
  INV_X1 U5278 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4865) );
  AOI22_X1 U5279 ( .A1(n5253), .A2(n4867), .B1(n4865), .B2(n5251), .ZN(U3520)
         );
  INV_X1 U5280 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4866) );
  AOI22_X1 U5281 ( .A1(n5257), .A2(n4867), .B1(n4866), .B2(n5254), .ZN(U3471)
         );
  XNOR2_X1 U5282 ( .A(n4868), .B(n4870), .ZN(n4887) );
  XNOR2_X1 U5283 ( .A(n4869), .B(n4870), .ZN(n4873) );
  AOI21_X1 U5284 ( .B1(n4879), .B2(n5229), .A(n4871), .ZN(n4872) );
  OAI21_X1 U5285 ( .B1(n4873), .B2(n5091), .A(n4872), .ZN(n4874) );
  AOI21_X1 U5286 ( .B1(n4875), .B2(n4887), .A(n4874), .ZN(n4890) );
  INV_X1 U5287 ( .A(n4876), .ZN(n4877) );
  AOI21_X1 U5288 ( .B1(n4879), .B2(n4878), .A(n4877), .ZN(n4885) );
  AOI22_X1 U5289 ( .A1(n4887), .A2(n4896), .B1(n5249), .B2(n4885), .ZN(n4880)
         );
  AND2_X1 U5290 ( .A1(n4890), .A2(n4880), .ZN(n4883) );
  AOI22_X1 U5291 ( .A1(n5253), .A2(n4883), .B1(n4881), .B2(n5251), .ZN(U3521)
         );
  INV_X1 U5292 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4882) );
  AOI22_X1 U5293 ( .A1(n5257), .A2(n4883), .B1(n4882), .B2(n5254), .ZN(U3473)
         );
  AOI22_X1 U5294 ( .A1(n5246), .A2(REG2_REG_3__SCAN_IN), .B1(n5136), .B2(n4884), .ZN(n4889) );
  AOI22_X1 U5295 ( .A1(n4887), .A2(n4886), .B1(n5244), .B2(n4885), .ZN(n4888)
         );
  OAI211_X1 U5296 ( .C1(n5246), .C2(n4890), .A(n4889), .B(n4888), .ZN(U3287)
         );
  INV_X1 U5297 ( .A(DATAI_4_), .ZN(n4891) );
  AOI22_X1 U5298 ( .A1(STATE_REG_SCAN_IN), .A2(n4892), .B1(n4891), .B2(U3149), 
        .ZN(U3348) );
  INV_X1 U5299 ( .A(n4893), .ZN(n4897) );
  AOI211_X1 U5300 ( .C1(n4897), .C2(n4896), .A(n4895), .B(n4894), .ZN(n4900)
         );
  AOI22_X1 U5301 ( .A1(n5253), .A2(n4900), .B1(n4898), .B2(n5251), .ZN(U3522)
         );
  INV_X1 U5302 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4899) );
  AOI22_X1 U5303 ( .A1(n5257), .A2(n4900), .B1(n4899), .B2(n5254), .ZN(U3475)
         );
  OAI22_X1 U5304 ( .A1(U3149), .A2(n4901), .B1(DATAI_5_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4902) );
  INV_X1 U5305 ( .A(n4902), .ZN(U3347) );
  INV_X1 U5306 ( .A(n5190), .ZN(n4905) );
  INV_X1 U5307 ( .A(n4903), .ZN(n4904) );
  OAI21_X1 U5308 ( .B1(n4906), .B2(n4905), .A(n4904), .ZN(n4912) );
  NAND2_X1 U5309 ( .A1(n4908), .A2(n4907), .ZN(n4909) );
  AOI21_X1 U5310 ( .B1(n4910), .B2(n4909), .A(n5186), .ZN(n4911) );
  AOI211_X1 U5311 ( .C1(n4913), .C2(n5160), .A(n4912), .B(n4911), .ZN(n4914)
         );
  OAI21_X1 U5312 ( .B1(n5192), .B2(n4915), .A(n4914), .ZN(U3224) );
  NOR2_X1 U5313 ( .A1(n4916), .A2(n5219), .ZN(n4918) );
  AOI211_X1 U5314 ( .C1(n5221), .C2(n4919), .A(n4918), .B(n4917), .ZN(n4922)
         );
  INV_X1 U5315 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4920) );
  AOI22_X1 U5316 ( .A1(n5253), .A2(n4922), .B1(n4920), .B2(n5251), .ZN(U3523)
         );
  AOI22_X1 U5317 ( .A1(n5257), .A2(n4922), .B1(n4921), .B2(n5254), .ZN(U3477)
         );
  OAI22_X1 U5318 ( .A1(U3149), .A2(n4923), .B1(DATAI_6_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4924) );
  INV_X1 U5319 ( .A(n4924), .ZN(U3346) );
  OAI21_X1 U5320 ( .B1(n5219), .B2(n4926), .A(n4925), .ZN(n4927) );
  AOI21_X1 U5321 ( .B1(n5221), .B2(n4928), .A(n4927), .ZN(n4931) );
  AOI22_X1 U5322 ( .A1(n5253), .A2(n4931), .B1(n4929), .B2(n5251), .ZN(U3524)
         );
  INV_X1 U5323 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4930) );
  AOI22_X1 U5324 ( .A1(n5257), .A2(n4931), .B1(n4930), .B2(n5254), .ZN(U3479)
         );
  OAI22_X1 U5325 ( .A1(U3149), .A2(n4932), .B1(DATAI_7_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4933) );
  INV_X1 U5326 ( .A(n4933), .ZN(U3345) );
  NOR2_X1 U5327 ( .A1(n4934), .A2(n5169), .ZN(n4937) );
  AOI211_X1 U5328 ( .C1(n4937), .C2(n3554), .A(n4936), .B(n4935), .ZN(n4940)
         );
  INV_X1 U5329 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4938) );
  AOI22_X1 U5330 ( .A1(n5253), .A2(n4940), .B1(n4938), .B2(n5251), .ZN(U3525)
         );
  AOI22_X1 U5331 ( .A1(n5257), .A2(n4940), .B1(n4939), .B2(n5254), .ZN(U3481)
         );
  AOI22_X1 U5332 ( .A1(STATE_REG_SCAN_IN), .A2(n4942), .B1(n4941), .B2(U3149), 
        .ZN(U3344) );
  AND2_X1 U5333 ( .A1(n3584), .A2(n4943), .ZN(n4946) );
  OAI21_X1 U5334 ( .B1(n4946), .B2(n4945), .A(n4944), .ZN(n4952) );
  AOI21_X1 U5335 ( .B1(n5190), .B2(n4948), .A(n4947), .ZN(n4949) );
  OAI21_X1 U5336 ( .B1(n5185), .B2(n4950), .A(n4949), .ZN(n4951) );
  AOI21_X1 U5337 ( .B1(n4952), .B2(n5162), .A(n4951), .ZN(n4953) );
  OAI21_X1 U5338 ( .B1(n5192), .B2(n4954), .A(n4953), .ZN(U3218) );
  NOR2_X1 U5339 ( .A1(n4955), .A2(n5169), .ZN(n4956) );
  AOI211_X1 U5340 ( .C1(n5249), .C2(n4958), .A(n4957), .B(n4956), .ZN(n4961)
         );
  AOI22_X1 U5341 ( .A1(n5253), .A2(n4961), .B1(n4959), .B2(n5251), .ZN(U3526)
         );
  INV_X1 U5342 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4960) );
  AOI22_X1 U5343 ( .A1(n5257), .A2(n4961), .B1(n4960), .B2(n5254), .ZN(U3483)
         );
  XNOR2_X1 U5344 ( .A(n4962), .B(n4967), .ZN(n4980) );
  NOR2_X1 U5345 ( .A1(n4963), .A2(n4969), .ZN(n4964) );
  OR2_X1 U5346 ( .A1(n3618), .A2(n4964), .ZN(n4978) );
  NAND2_X1 U5347 ( .A1(n4966), .A2(n4965), .ZN(n4968) );
  XNOR2_X1 U5348 ( .A(n4968), .B(n4967), .ZN(n4972) );
  NOR2_X1 U5349 ( .A1(n4969), .A2(n5237), .ZN(n4971) );
  AOI211_X1 U5350 ( .C1(n4972), .C2(n5207), .A(n4971), .B(n4970), .ZN(n4982)
         );
  OAI21_X1 U5351 ( .B1(n5219), .B2(n4978), .A(n4982), .ZN(n4973) );
  AOI21_X1 U5352 ( .B1(n4980), .B2(n5221), .A(n4973), .ZN(n4976) );
  INV_X1 U5353 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4974) );
  AOI22_X1 U5354 ( .A1(n5253), .A2(n4976), .B1(n4974), .B2(n5251), .ZN(U3527)
         );
  INV_X1 U5355 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4975) );
  AOI22_X1 U5356 ( .A1(n5257), .A2(n4976), .B1(n4975), .B2(n5254), .ZN(U3485)
         );
  INV_X1 U5357 ( .A(REG2_REG_9__SCAN_IN), .ZN(n4977) );
  OAI22_X1 U5358 ( .A1(n4978), .A2(n5196), .B1(n4977), .B2(n4558), .ZN(n4979)
         );
  INV_X1 U5359 ( .A(n4979), .ZN(n4986) );
  INV_X1 U5360 ( .A(n4980), .ZN(n4983) );
  INV_X1 U5361 ( .A(n4981), .ZN(n5209) );
  OAI21_X1 U5362 ( .B1(n4983), .B2(n5209), .A(n4982), .ZN(n4984) );
  NAND2_X1 U5363 ( .A1(n4984), .A2(n4558), .ZN(n4985) );
  OAI211_X1 U5364 ( .C1(n5216), .C2(n4987), .A(n4986), .B(n4985), .ZN(U3281)
         );
  OAI22_X1 U5365 ( .A1(n4989), .A2(n5169), .B1(n4988), .B2(n5219), .ZN(n4990)
         );
  NOR2_X1 U5366 ( .A1(n4991), .A2(n4990), .ZN(n4994) );
  AOI22_X1 U5367 ( .A1(n5253), .A2(n4994), .B1(n4992), .B2(n5251), .ZN(U3528)
         );
  INV_X1 U5368 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4993) );
  AOI22_X1 U5369 ( .A1(n5257), .A2(n4994), .B1(n4993), .B2(n5254), .ZN(U3487)
         );
  OAI22_X1 U5370 ( .A1(U3149), .A2(n4995), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4996) );
  INV_X1 U5371 ( .A(n4996), .ZN(U3341) );
  AOI22_X1 U5372 ( .A1(n5190), .A2(n4997), .B1(REG3_REG_11__SCAN_IN), .B2(
        U3149), .ZN(n5008) );
  INV_X1 U5373 ( .A(n5001), .ZN(n5003) );
  OR2_X1 U5374 ( .A1(n4998), .A2(n5004), .ZN(n5000) );
  AOI21_X1 U5375 ( .B1(n5001), .B2(n5000), .A(n4999), .ZN(n5002) );
  AOI211_X1 U5376 ( .C1(n5004), .C2(n5003), .A(n5186), .B(n5002), .ZN(n5005)
         );
  AOI21_X1 U5377 ( .B1(n5006), .B2(n5160), .A(n5005), .ZN(n5007) );
  OAI211_X1 U5378 ( .C1(n5192), .C2(n5009), .A(n5008), .B(n5007), .ZN(U3233)
         );
  OAI21_X1 U5379 ( .B1(n5219), .B2(n5011), .A(n5010), .ZN(n5012) );
  AOI21_X1 U5380 ( .B1(n5013), .B2(n5221), .A(n5012), .ZN(n5016) );
  INV_X1 U5381 ( .A(REG1_REG_11__SCAN_IN), .ZN(n5014) );
  AOI22_X1 U5382 ( .A1(n5253), .A2(n5016), .B1(n5014), .B2(n5251), .ZN(U3529)
         );
  INV_X1 U5383 ( .A(REG0_REG_11__SCAN_IN), .ZN(n5015) );
  AOI22_X1 U5384 ( .A1(n5257), .A2(n5016), .B1(n5015), .B2(n5254), .ZN(U3489)
         );
  OAI22_X1 U5385 ( .A1(U3149), .A2(n5017), .B1(DATAI_12_), .B2(
        STATE_REG_SCAN_IN), .ZN(n5018) );
  INV_X1 U5386 ( .A(n5018), .ZN(U3340) );
  AOI22_X1 U5387 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .B1(n5190), .B2(
        n5019), .ZN(n5025) );
  XNOR2_X1 U5388 ( .A(n5021), .B(n5020), .ZN(n5023) );
  AOI22_X1 U5389 ( .A1(n5023), .A2(n5162), .B1(n5022), .B2(n5160), .ZN(n5024)
         );
  OAI211_X1 U5390 ( .C1(n5192), .C2(n5026), .A(n5025), .B(n5024), .ZN(U3221)
         );
  OAI22_X1 U5391 ( .A1(n5028), .A2(n5169), .B1(n5027), .B2(n5219), .ZN(n5029)
         );
  NOR2_X1 U5392 ( .A1(n5030), .A2(n5029), .ZN(n5033) );
  AOI22_X1 U5393 ( .A1(n5253), .A2(n5033), .B1(n5031), .B2(n5251), .ZN(U3530)
         );
  INV_X1 U5394 ( .A(REG0_REG_12__SCAN_IN), .ZN(n5032) );
  AOI22_X1 U5395 ( .A1(n5257), .A2(n5033), .B1(n5032), .B2(n5254), .ZN(U3491)
         );
  OAI22_X1 U5396 ( .A1(U3149), .A2(n5034), .B1(DATAI_13_), .B2(
        STATE_REG_SCAN_IN), .ZN(n5035) );
  INV_X1 U5397 ( .A(n5035), .ZN(U3339) );
  AOI22_X1 U5398 ( .A1(REG3_REG_13__SCAN_IN), .A2(U3149), .B1(n5190), .B2(
        n5036), .ZN(n5042) );
  XNOR2_X1 U5399 ( .A(n5037), .B(n5038), .ZN(n5040) );
  AOI22_X1 U5400 ( .A1(n5040), .A2(n5162), .B1(n5039), .B2(n5160), .ZN(n5041)
         );
  OAI211_X1 U5401 ( .C1(n5192), .C2(n5043), .A(n5042), .B(n5041), .ZN(U3231)
         );
  NOR2_X1 U5402 ( .A1(n5044), .A2(n5169), .ZN(n5045) );
  AOI211_X1 U5403 ( .C1(n5249), .C2(n5047), .A(n5046), .B(n5045), .ZN(n5050)
         );
  INV_X1 U5404 ( .A(REG1_REG_13__SCAN_IN), .ZN(n5048) );
  AOI22_X1 U5405 ( .A1(n5253), .A2(n5050), .B1(n5048), .B2(n5251), .ZN(U3531)
         );
  INV_X1 U5406 ( .A(REG0_REG_13__SCAN_IN), .ZN(n5049) );
  AOI22_X1 U5407 ( .A1(n5257), .A2(n5050), .B1(n5049), .B2(n5254), .ZN(U3493)
         );
  AOI22_X1 U5408 ( .A1(STATE_REG_SCAN_IN), .A2(n5052), .B1(n5051), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5409 ( .A(n5053), .ZN(n5061) );
  AOI22_X1 U5410 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .B1(n5190), .B2(
        n5054), .ZN(n5060) );
  XNOR2_X1 U5411 ( .A(n5056), .B(n5055), .ZN(n5058) );
  AOI22_X1 U5412 ( .A1(n5058), .A2(n5162), .B1(n5057), .B2(n5160), .ZN(n5059)
         );
  OAI211_X1 U5413 ( .C1(n5192), .C2(n5061), .A(n5060), .B(n5059), .ZN(U3212)
         );
  INV_X1 U5414 ( .A(n5062), .ZN(n5063) );
  OAI21_X1 U5415 ( .B1(n5219), .B2(n5064), .A(n5063), .ZN(n5065) );
  AOI21_X1 U5416 ( .B1(n5221), .B2(n5066), .A(n5065), .ZN(n5069) );
  AOI22_X1 U5417 ( .A1(n5253), .A2(n5069), .B1(n5067), .B2(n5251), .ZN(U3532)
         );
  INV_X1 U5418 ( .A(REG0_REG_14__SCAN_IN), .ZN(n5068) );
  AOI22_X1 U5419 ( .A1(n5257), .A2(n5069), .B1(n5068), .B2(n5254), .ZN(U3495)
         );
  OAI22_X1 U5420 ( .A1(n5122), .A2(n5121), .B1(n5070), .B2(n5175), .ZN(n5088)
         );
  AOI22_X1 U5421 ( .A1(REG3_REG_15__SCAN_IN), .A2(U3149), .B1(n5190), .B2(
        n5088), .ZN(n5077) );
  XNOR2_X1 U5422 ( .A(n5072), .B(n5071), .ZN(n5073) );
  XNOR2_X1 U5423 ( .A(n5074), .B(n5073), .ZN(n5075) );
  AOI22_X1 U5424 ( .A1(n5075), .A2(n5162), .B1(n5089), .B2(n5160), .ZN(n5076)
         );
  OAI211_X1 U5425 ( .C1(n5192), .C2(n5078), .A(n5077), .B(n5076), .ZN(U3238)
         );
  AOI21_X1 U5426 ( .B1(n5089), .B2(n3826), .A(n2521), .ZN(n5098) );
  OAI21_X1 U5427 ( .B1(n5081), .B2(n5080), .A(n5079), .ZN(n5083) );
  XNOR2_X1 U5428 ( .A(n5083), .B(n5082), .ZN(n5102) );
  NOR2_X1 U5429 ( .A1(n5169), .A2(n5102), .ZN(n5093) );
  NAND2_X1 U5430 ( .A1(n5085), .A2(n5084), .ZN(n5087) );
  XNOR2_X1 U5431 ( .A(n5087), .B(n5086), .ZN(n5092) );
  AOI21_X1 U5432 ( .B1(n5089), .B2(n5229), .A(n5088), .ZN(n5090) );
  OAI21_X1 U5433 ( .B1(n5092), .B2(n5091), .A(n5090), .ZN(n5099) );
  AOI211_X1 U5434 ( .C1(n5098), .C2(n5249), .A(n5093), .B(n5099), .ZN(n5096)
         );
  INV_X1 U5435 ( .A(REG1_REG_15__SCAN_IN), .ZN(n5094) );
  AOI22_X1 U5436 ( .A1(n5253), .A2(n5096), .B1(n5094), .B2(n5251), .ZN(U3533)
         );
  INV_X1 U5437 ( .A(REG0_REG_15__SCAN_IN), .ZN(n5095) );
  AOI22_X1 U5438 ( .A1(n5257), .A2(n5096), .B1(n5095), .B2(n5254), .ZN(U3497)
         );
  AOI22_X1 U5439 ( .A1(REG2_REG_15__SCAN_IN), .A2(n5246), .B1(n5097), .B2(
        n5136), .ZN(n5101) );
  AOI22_X1 U5440 ( .A1(n5099), .A2(n4558), .B1(n5098), .B2(n5244), .ZN(n5100)
         );
  OAI211_X1 U5441 ( .C1(n5103), .C2(n5102), .A(n5101), .B(n5100), .ZN(U3275)
         );
  AOI22_X1 U5442 ( .A1(STATE_REG_SCAN_IN), .A2(n5105), .B1(n5104), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5443 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .B1(n5190), .B2(
        n5106), .ZN(n5112) );
  XNOR2_X1 U5444 ( .A(n5108), .B(n5107), .ZN(n5110) );
  AOI22_X1 U5445 ( .A1(n5110), .A2(n5162), .B1(n5109), .B2(n5160), .ZN(n5111)
         );
  OAI211_X1 U5446 ( .C1(n5192), .C2(n5113), .A(n5112), .B(n5111), .ZN(U3223)
         );
  OAI22_X1 U5447 ( .A1(n5115), .A2(n5169), .B1(n5114), .B2(n5219), .ZN(n5116)
         );
  NOR2_X1 U5448 ( .A1(n5117), .A2(n5116), .ZN(n5120) );
  AOI22_X1 U5449 ( .A1(n5253), .A2(n5120), .B1(n5118), .B2(n5251), .ZN(U3534)
         );
  INV_X1 U5450 ( .A(REG0_REG_16__SCAN_IN), .ZN(n5119) );
  AOI22_X1 U5451 ( .A1(n5257), .A2(n5120), .B1(n5119), .B2(n5254), .ZN(U3499)
         );
  INV_X1 U5452 ( .A(n5137), .ZN(n5131) );
  OR2_X1 U5453 ( .A1(n5176), .A2(n5121), .ZN(n5124) );
  OR2_X1 U5454 ( .A1(n5122), .A2(n5175), .ZN(n5123) );
  NAND2_X1 U5455 ( .A1(n5124), .A2(n5123), .ZN(n5133) );
  AOI22_X1 U5456 ( .A1(REG3_REG_17__SCAN_IN), .A2(U3149), .B1(n5190), .B2(
        n5133), .ZN(n5130) );
  XNOR2_X1 U5457 ( .A(n5126), .B(n5125), .ZN(n5128) );
  AOI22_X1 U5458 ( .A1(n5128), .A2(n5162), .B1(n5127), .B2(n5160), .ZN(n5129)
         );
  OAI211_X1 U5459 ( .C1(n5192), .C2(n5131), .A(n5130), .B(n5129), .ZN(U3225)
         );
  XNOR2_X1 U5460 ( .A(n5132), .B(n5138), .ZN(n5135) );
  NOR2_X1 U5461 ( .A1(n5142), .A2(n5237), .ZN(n5134) );
  AOI211_X1 U5462 ( .C1(n5135), .C2(n5207), .A(n5134), .B(n5133), .ZN(n5147)
         );
  AOI22_X1 U5463 ( .A1(REG2_REG_17__SCAN_IN), .A2(n5246), .B1(n5137), .B2(
        n5136), .ZN(n5146) );
  XNOR2_X1 U5464 ( .A(n5139), .B(n5138), .ZN(n5150) );
  INV_X1 U5465 ( .A(n5140), .ZN(n5141) );
  OAI21_X1 U5466 ( .B1(n2545), .B2(n5142), .A(n5141), .ZN(n5148) );
  INV_X1 U5467 ( .A(n5148), .ZN(n5143) );
  AOI22_X1 U5468 ( .A1(n5150), .A2(n5144), .B1(n5244), .B2(n5143), .ZN(n5145)
         );
  OAI211_X1 U5469 ( .C1(n5246), .C2(n5147), .A(n5146), .B(n5145), .ZN(U3273)
         );
  OAI21_X1 U5470 ( .B1(n5219), .B2(n5148), .A(n5147), .ZN(n5149) );
  AOI21_X1 U5471 ( .B1(n5150), .B2(n5221), .A(n5149), .ZN(n5153) );
  INV_X1 U5472 ( .A(REG1_REG_17__SCAN_IN), .ZN(n5151) );
  AOI22_X1 U5473 ( .A1(n5253), .A2(n5153), .B1(n5151), .B2(n5251), .ZN(U3535)
         );
  INV_X1 U5474 ( .A(REG0_REG_17__SCAN_IN), .ZN(n5152) );
  AOI22_X1 U5475 ( .A1(n5257), .A2(n5153), .B1(n5152), .B2(n5254), .ZN(U3501)
         );
  OAI22_X1 U5476 ( .A1(U3149), .A2(n5154), .B1(DATAI_18_), .B2(
        STATE_REG_SCAN_IN), .ZN(n5155) );
  INV_X1 U5477 ( .A(n5155), .ZN(U3334) );
  AOI22_X1 U5478 ( .A1(REG3_REG_18__SCAN_IN), .A2(U3149), .B1(n5190), .B2(
        n5156), .ZN(n5165) );
  NAND2_X1 U5479 ( .A1(n2522), .A2(n5157), .ZN(n5158) );
  XNOR2_X1 U5480 ( .A(n5159), .B(n5158), .ZN(n5163) );
  AOI22_X1 U5481 ( .A1(n5163), .A2(n5162), .B1(n5161), .B2(n5160), .ZN(n5164)
         );
  OAI211_X1 U5482 ( .C1(n5192), .C2(n5166), .A(n5165), .B(n5164), .ZN(U3235)
         );
  OAI211_X1 U5483 ( .C1(n5170), .C2(n5169), .A(n5168), .B(n5167), .ZN(n5171)
         );
  INV_X1 U5484 ( .A(n5171), .ZN(n5174) );
  INV_X1 U5485 ( .A(REG1_REG_18__SCAN_IN), .ZN(n5172) );
  AOI22_X1 U5486 ( .A1(n5253), .A2(n5174), .B1(n5172), .B2(n5251), .ZN(U3536)
         );
  INV_X1 U5487 ( .A(REG0_REG_18__SCAN_IN), .ZN(n5173) );
  AOI22_X1 U5488 ( .A1(n5257), .A2(n5174), .B1(n5173), .B2(n5254), .ZN(U3503)
         );
  OR2_X1 U5489 ( .A1(n5176), .A2(n5175), .ZN(n5180) );
  NAND2_X1 U5490 ( .A1(n5178), .A2(n5177), .ZN(n5179) );
  NAND2_X1 U5491 ( .A1(n5180), .A2(n5179), .ZN(n5205) );
  OAI21_X1 U5492 ( .B1(n5183), .B2(n5182), .A(n5181), .ZN(n5184) );
  INV_X1 U5493 ( .A(n5184), .ZN(n5187) );
  OAI22_X1 U5494 ( .A1(n5187), .A2(n5186), .B1(n5185), .B2(n5204), .ZN(n5188)
         );
  AOI211_X1 U5495 ( .C1(n5190), .C2(n5205), .A(n5189), .B(n5188), .ZN(n5191)
         );
  OAI21_X1 U5496 ( .B1(n5192), .B2(n5215), .A(n5191), .ZN(U3216) );
  NAND2_X1 U5497 ( .A1(n4538), .A2(n5193), .ZN(n5194) );
  NAND2_X1 U5498 ( .A1(n5195), .A2(n5194), .ZN(n5218) );
  OAI22_X1 U5499 ( .A1(n5218), .A2(n5196), .B1(n3876), .B2(n4558), .ZN(n5197)
         );
  INV_X1 U5500 ( .A(n5197), .ZN(n5214) );
  OAI21_X1 U5501 ( .B1(n5199), .B2(n5202), .A(n5198), .ZN(n5222) );
  INV_X1 U5502 ( .A(n5222), .ZN(n5210) );
  NAND2_X1 U5503 ( .A1(n5201), .A2(n5200), .ZN(n5203) );
  XNOR2_X1 U5504 ( .A(n5203), .B(n5202), .ZN(n5208) );
  NOR2_X1 U5505 ( .A1(n5204), .A2(n5237), .ZN(n5206) );
  AOI211_X1 U5506 ( .C1(n5208), .C2(n5207), .A(n5206), .B(n5205), .ZN(n5217)
         );
  OAI21_X1 U5507 ( .B1(n5210), .B2(n5209), .A(n5217), .ZN(n5212) );
  NAND2_X1 U5508 ( .A1(n5212), .A2(n4558), .ZN(n5213) );
  OAI211_X1 U5509 ( .C1(n5216), .C2(n5215), .A(n5214), .B(n5213), .ZN(U3271)
         );
  OAI21_X1 U5510 ( .B1(n5219), .B2(n5218), .A(n5217), .ZN(n5220) );
  AOI21_X1 U5511 ( .B1(n5222), .B2(n5221), .A(n5220), .ZN(n5225) );
  AOI22_X1 U5512 ( .A1(n5253), .A2(n5225), .B1(n5223), .B2(n5251), .ZN(U3537)
         );
  INV_X1 U5513 ( .A(REG0_REG_19__SCAN_IN), .ZN(n5224) );
  AOI22_X1 U5514 ( .A1(n5257), .A2(n5225), .B1(n5224), .B2(n5254), .ZN(U3505)
         );
  NAND2_X1 U5515 ( .A1(n5227), .A2(n5226), .ZN(n5239) );
  INV_X1 U5516 ( .A(n5239), .ZN(n5228) );
  AOI21_X1 U5517 ( .B1(n5240), .B2(n5229), .A(n5228), .ZN(n5231) );
  XOR2_X1 U5518 ( .A(n5240), .B(n5241), .Z(n5233) );
  AOI22_X1 U5519 ( .A1(n5233), .A2(n5244), .B1(REG2_REG_30__SCAN_IN), .B2(
        n5246), .ZN(n5230) );
  OAI21_X1 U5520 ( .B1(n5246), .B2(n5231), .A(n5230), .ZN(U3261) );
  INV_X1 U5521 ( .A(n5231), .ZN(n5232) );
  INV_X1 U5522 ( .A(REG1_REG_30__SCAN_IN), .ZN(n5234) );
  AOI22_X1 U5523 ( .A1(n5253), .A2(n5236), .B1(n5234), .B2(n5251), .ZN(U3548)
         );
  INV_X1 U5524 ( .A(REG0_REG_30__SCAN_IN), .ZN(n5235) );
  AOI22_X1 U5525 ( .A1(n5257), .A2(n5236), .B1(n5235), .B2(n5254), .ZN(U3516)
         );
  OR2_X1 U5526 ( .A1(n5243), .A2(n5237), .ZN(n5238) );
  AND2_X1 U5527 ( .A1(n5239), .A2(n5238), .ZN(n5247) );
  XOR2_X1 U5528 ( .A(n5243), .B(n5242), .Z(n5250) );
  AOI22_X1 U5529 ( .A1(n5250), .A2(n5244), .B1(n5246), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n5245) );
  OAI21_X1 U5530 ( .B1(n5246), .B2(n5247), .A(n5245), .ZN(U3260) );
  INV_X1 U5531 ( .A(n5247), .ZN(n5248) );
  AOI21_X1 U5532 ( .B1(n5250), .B2(n5249), .A(n5248), .ZN(n5256) );
  INV_X1 U5533 ( .A(REG1_REG_31__SCAN_IN), .ZN(n5252) );
  AOI22_X1 U5534 ( .A1(n5253), .A2(n5256), .B1(n5252), .B2(n5251), .ZN(U3549)
         );
  INV_X1 U5535 ( .A(REG0_REG_31__SCAN_IN), .ZN(n5255) );
  AOI22_X1 U5536 ( .A1(n5257), .A2(n5256), .B1(n5255), .B2(n5254), .ZN(U3517)
         );
  CLKBUF_X1 U2523 ( .A(n3469), .Z(n3987) );
  CLKBUF_X1 U2779 ( .A(n2977), .Z(n4199) );
  INV_X2 U3165 ( .A(n5246), .ZN(n4558) );
endmodule

