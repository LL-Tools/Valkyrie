

module b22_C_AntiSAT_k_128_3 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, 
        SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, 
        SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, 
        SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, 
        U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, 
        P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, 
        P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, 
        P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, 
        P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, 
        P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, 
        P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, 
        P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, 
        P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, 
        P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, 
        P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, 
        P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, 
        P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, 
        P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, 
        P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, 
        P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, 
        P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, 
        P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, 
        P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, 
        P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, 
        P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, 
        P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, 
        P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, 
        P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, 
        P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, 
        P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, 
        P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, 
        P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, 
        P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, 
        P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, 
        P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, 
        P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, 
        P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, 
        P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, 
        P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, 
        P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, 
        P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, 
        P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, 
        P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457;

  INV_X1 U7221 ( .A(n14896), .ZN(n14894) );
  AND2_X1 U7222 ( .A1(n13986), .A2(n13985), .ZN(n14191) );
  AND2_X1 U7223 ( .A1(n13437), .A2(n13436), .ZN(n13438) );
  NAND2_X1 U7224 ( .A1(n11620), .A2(n14582), .ZN(n11726) );
  INV_X1 U7226 ( .A(n10712), .ZN(n10963) );
  CLKBUF_X2 U7227 ( .A(n7846), .Z(n8211) );
  CLKBUF_X2 U7228 ( .A(n7853), .Z(n6474) );
  CLKBUF_X2 U7229 ( .A(n8614), .Z(n9967) );
  INV_X1 U7230 ( .A(n9744), .ZN(n9552) );
  CLKBUF_X2 U7231 ( .A(n7824), .Z(n10356) );
  INV_X1 U7232 ( .A(n12002), .ZN(n6476) );
  NOR4_X1 U7233 ( .A1(n9174), .A2(n12202), .A3(n8422), .A4(n12567), .ZN(n8424)
         );
  INV_X1 U7234 ( .A(n8307), .ZN(n9184) );
  INV_X1 U7235 ( .A(n12968), .ZN(n12937) );
  INV_X1 U7236 ( .A(n9290), .ZN(n9551) );
  NAND2_X1 U7237 ( .A1(n13997), .A2(n13996), .ZN(n9021) );
  NAND2_X1 U7238 ( .A1(n8450), .A2(n6488), .ZN(n7824) );
  INV_X1 U7239 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n7929) );
  AND3_X1 U7240 ( .A1(n9291), .A2(n7763), .A3(n9292), .ZN(n9786) );
  OAI21_X1 U7241 ( .B1(n14134), .B2(n12115), .A(n12113), .ZN(n14113) );
  NAND2_X1 U7242 ( .A1(n13972), .A2(n13973), .ZN(n14185) );
  NAND2_X1 U7243 ( .A1(n8635), .A2(n7237), .ZN(n7236) );
  OAI21_X1 U7244 ( .B1(n9939), .B2(n9286), .A(n9383), .ZN(n11222) );
  XNOR2_X1 U7245 ( .A(n6485), .B(n7029), .ZN(n13269) );
  OAI211_X1 U7246 ( .C1(n14185), .C2(n14273), .A(n14184), .B(n14186), .ZN(
        n14287) );
  INV_X1 U7247 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6920) );
  AND4_X1 U7248 ( .A1(n9198), .A2(n9197), .A3(n9457), .A4(n9476), .ZN(n6473)
         );
  AND2_X1 U7249 ( .A1(n7824), .A2(n9211), .ZN(n7853) );
  NAND2_X2 U7250 ( .A1(n11386), .A2(n11403), .ZN(n11385) );
  OR2_X2 U7251 ( .A1(n9492), .A2(n9493), .ZN(n7162) );
  NAND2_X2 U7252 ( .A1(n9072), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7059) );
  NAND2_X2 U7253 ( .A1(n8631), .A2(n8630), .ZN(n8635) );
  NAND2_X2 U7254 ( .A1(n11253), .A2(n11252), .ZN(n11255) );
  NAND2_X2 U7255 ( .A1(n11220), .A2(n11219), .ZN(n11253) );
  AOI21_X2 U7256 ( .B1(n12580), .B2(n8519), .A(n8518), .ZN(n12568) );
  OAI21_X2 U7257 ( .B1(n12623), .B2(n7678), .A(n6798), .ZN(n12580) );
  NAND2_X2 U7258 ( .A1(n8621), .A2(n6529), .ZN(n8631) );
  NAND4_X2 U7259 ( .A1(n7819), .A2(n7818), .A3(n7817), .A4(n7816), .ZN(n15201)
         );
  NAND2_X2 U7260 ( .A1(n9630), .A2(n9629), .ZN(n13488) );
  NAND2_X2 U7261 ( .A1(n14405), .A2(n14406), .ZN(n14453) );
  AND3_X4 U7262 ( .A1(n9277), .A2(n9278), .A3(n7760), .ZN(n6766) );
  AND2_X2 U7263 ( .A1(n11944), .A2(n12085), .ZN(n11942) );
  AND2_X2 U7264 ( .A1(n12085), .A2(n9124), .ZN(n11941) );
  NAND2_X2 U7265 ( .A1(n8573), .A2(n7748), .ZN(n7060) );
  OAI21_X2 U7266 ( .B1(n9041), .B2(n9040), .A(n9039), .ZN(n9053) );
  NOR2_X2 U7267 ( .A1(n8109), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8120) );
  AOI21_X2 U7268 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n13922), .A(n14754), .ZN(
        n13924) );
  AND2_X2 U7269 ( .A1(n14751), .A2(n14750), .ZN(n14754) );
  NAND2_X2 U7270 ( .A1(n13912), .A2(n7050), .ZN(n14693) );
  INV_X2 U7271 ( .A(n8918), .ZN(n6475) );
  INV_X1 U7272 ( .A(n8918), .ZN(n8594) );
  NOR2_X2 U7273 ( .A1(n11579), .A2(n11582), .ZN(n11753) );
  NAND2_X2 U7274 ( .A1(n6879), .A2(n8855), .ZN(n14134) );
  OAI21_X2 U7275 ( .B1(n9821), .B2(n6602), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9207) );
  AOI21_X4 U7276 ( .B1(n14454), .B2(n14407), .A(n14451), .ZN(n15453) );
  XNOR2_X2 U7277 ( .A(n7174), .B(n7052), .ZN(n10156) );
  NAND2_X1 U7278 ( .A1(n8977), .A2(n8976), .ZN(n14211) );
  OAI21_X1 U7279 ( .B1(n11654), .B2(n7629), .A(n7627), .ZN(n14543) );
  NOR2_X1 U7280 ( .A1(n13546), .A2(n13076), .ZN(n6607) );
  NOR2_X1 U7281 ( .A1(n14559), .A2(n13077), .ZN(n6610) );
  NAND2_X1 U7282 ( .A1(n10993), .A2(n10992), .ZN(n11129) );
  NAND2_X1 U7283 ( .A1(n9412), .A2(n9411), .ZN(n11465) );
  NAND2_X1 U7284 ( .A1(n9360), .A2(n9359), .ZN(n15048) );
  NAND2_X1 U7285 ( .A1(n8407), .A2(n8406), .ZN(n8482) );
  INV_X1 U7286 ( .A(n10631), .ZN(n10637) );
  INV_X1 U7287 ( .A(n12374), .ZN(n7815) );
  NOR2_X1 U7288 ( .A1(n14675), .A2(n14671), .ZN(n14749) );
  NOR2_X1 U7289 ( .A1(n14675), .A2(n10301), .ZN(n14778) );
  INV_X2 U7290 ( .A(n10276), .ZN(n14861) );
  NAND2_X2 U7291 ( .A1(n10183), .A2(n10182), .ZN(n13615) );
  CLKBUF_X2 U7292 ( .A(n10220), .Z(n7054) );
  CLKBUF_X2 U7293 ( .A(n7844), .Z(n8212) );
  NAND2_X1 U7294 ( .A1(n10565), .A2(n9248), .ZN(n6526) );
  BUF_X2 U7295 ( .A(n9281), .Z(n9713) );
  CLKBUF_X2 U7296 ( .A(n6525), .Z(n9656) );
  INV_X4 U7297 ( .A(n14837), .ZN(n10182) );
  INV_X1 U7298 ( .A(n9413), .ZN(n9293) );
  NAND2_X2 U7300 ( .A1(n9290), .A2(n9211), .ZN(n9744) );
  NAND2_X2 U7301 ( .A1(n9290), .A2(n9676), .ZN(n9286) );
  AND2_X1 U7302 ( .A1(n9077), .A2(n9155), .ZN(n14348) );
  NAND2_X1 U7303 ( .A1(n9676), .A2(P1_U3086), .ZN(n14347) );
  NAND3_X1 U7304 ( .A1(n9199), .A2(n9212), .A3(n9204), .ZN(n9821) );
  AOI21_X1 U7305 ( .B1(n14287), .B2(n14896), .A(n7001), .ZN(n14187) );
  OAI21_X1 U7306 ( .B1(n14178), .B2(n14889), .A(n7058), .ZN(n9164) );
  NAND2_X1 U7307 ( .A1(n6484), .A2(n6483), .ZN(n13552) );
  AND2_X1 U7308 ( .A1(n13457), .A2(n13271), .ZN(n6483) );
  NOR2_X1 U7309 ( .A1(n12769), .A2(n6732), .ZN(n12830) );
  AOI21_X1 U7310 ( .B1(n7529), .B2(n12547), .A(n7526), .ZN(n12525) );
  NAND2_X1 U7311 ( .A1(n7579), .A2(n7577), .ZN(n14019) );
  NAND2_X1 U7312 ( .A1(n7178), .A2(n7177), .ZN(n13452) );
  NAND2_X1 U7313 ( .A1(n12566), .A2(n7700), .ZN(n9166) );
  NAND2_X1 U7314 ( .A1(n13277), .A2(n13267), .ZN(n13263) );
  NAND2_X1 U7315 ( .A1(n13327), .A2(n6481), .ZN(n13311) );
  OAI21_X1 U7316 ( .B1(n14044), .B2(n7457), .A(n7455), .ZN(n14000) );
  AOI21_X1 U7317 ( .B1(n6876), .B2(n7576), .A(n6502), .ZN(n6874) );
  XNOR2_X1 U7318 ( .A(n13201), .B(n13200), .ZN(n9802) );
  NAND2_X1 U7319 ( .A1(n7186), .A2(n7185), .ZN(n13288) );
  NAND2_X1 U7320 ( .A1(n6482), .A2(n7355), .ZN(n13327) );
  NAND2_X1 U7321 ( .A1(n13353), .A2(n7357), .ZN(n6482) );
  NAND2_X1 U7322 ( .A1(n9746), .A2(n9745), .ZN(n13204) );
  CLKBUF_X1 U7323 ( .A(n11938), .Z(n14323) );
  AOI21_X1 U7324 ( .B1(n13929), .B2(n14749), .A(n14778), .ZN(n7173) );
  INV_X1 U7325 ( .A(n12652), .ZN(n12653) );
  NAND2_X1 U7326 ( .A1(n12652), .A2(n8513), .ZN(n12639) );
  NOR2_X1 U7327 ( .A1(n12430), .A2(n12748), .ZN(n12457) );
  NAND2_X1 U7328 ( .A1(n9043), .A2(n9042), .ZN(n14288) );
  NAND2_X1 U7329 ( .A1(n6917), .A2(n6915), .ZN(n14046) );
  OR2_X1 U7330 ( .A1(n13335), .A2(n13251), .ZN(n6481) );
  NAND2_X1 U7331 ( .A1(n13243), .A2(n13242), .ZN(n13381) );
  NOR2_X1 U7332 ( .A1(n12407), .A2(n12409), .ZN(n12428) );
  NOR2_X1 U7333 ( .A1(n12383), .A2(n12385), .ZN(n12405) );
  NAND2_X1 U7334 ( .A1(n7051), .A2(n7587), .ZN(n14144) );
  OR2_X1 U7335 ( .A1(n7510), .A2(n14663), .ZN(n7505) );
  AND2_X1 U7336 ( .A1(n7290), .A2(n7288), .ZN(n12406) );
  NOR2_X1 U7337 ( .A1(n12471), .A2(n12470), .ZN(n12488) );
  NAND2_X1 U7338 ( .A1(n13235), .A2(n13234), .ZN(n13430) );
  OR2_X1 U7339 ( .A1(n14439), .A2(n14438), .ZN(n7510) );
  AND2_X1 U7340 ( .A1(n14439), .A2(n14438), .ZN(n14659) );
  OR2_X1 U7341 ( .A1(n12575), .A2(n8523), .ZN(n8389) );
  NAND2_X1 U7342 ( .A1(n6646), .A2(n6515), .ZN(n12753) );
  NAND2_X1 U7343 ( .A1(n11923), .A2(n11922), .ZN(n13235) );
  NOR2_X1 U7344 ( .A1(n12443), .A2(n12444), .ZN(n12468) );
  AND2_X1 U7345 ( .A1(n8264), .A2(n8263), .ZN(n12602) );
  NAND2_X1 U7346 ( .A1(n13421), .A2(n13404), .ZN(n13398) );
  OR2_X1 U7347 ( .A1(n12469), .A2(n12442), .ZN(n12443) );
  NAND2_X1 U7348 ( .A1(n11469), .A2(n11468), .ZN(n11467) );
  AND2_X1 U7349 ( .A1(n13904), .A2(n14720), .ZN(n14738) );
  XNOR2_X1 U7350 ( .A(n8956), .B(SI_22_), .ZN(n9598) );
  NAND2_X1 U7351 ( .A1(n11443), .A2(n12130), .ZN(n11442) );
  OR2_X1 U7352 ( .A1(n11577), .A2(n11576), .ZN(n11578) );
  NAND2_X1 U7353 ( .A1(n8162), .A2(n8163), .ZN(n8175) );
  NAND2_X1 U7354 ( .A1(n6699), .A2(n11720), .ZN(n11878) );
  NAND2_X1 U7355 ( .A1(n8910), .A2(n8909), .ZN(n8945) );
  NAND2_X1 U7356 ( .A1(n11559), .A2(n12128), .ZN(n11564) );
  NAND2_X1 U7357 ( .A1(n11529), .A2(n7018), .ZN(n11532) );
  OAI21_X1 U7358 ( .B1(n10870), .B2(n7460), .A(n6918), .ZN(n11375) );
  OR2_X1 U7359 ( .A1(n14559), .A2(n14573), .ZN(n6478) );
  NAND2_X1 U7360 ( .A1(n8128), .A2(n8127), .ZN(n8129) );
  AOI21_X1 U7361 ( .B1(n14976), .B2(n14426), .A(n14463), .ZN(n14427) );
  NAND2_X1 U7362 ( .A1(n11129), .A2(n6486), .ZN(n11220) );
  NAND2_X1 U7363 ( .A1(n9461), .A2(n9460), .ZN(n14573) );
  NAND2_X1 U7364 ( .A1(n8860), .A2(n8859), .ZN(n8874) );
  NAND2_X1 U7365 ( .A1(n9216), .A2(n9215), .ZN(n14559) );
  OR2_X1 U7366 ( .A1(n11229), .A2(n11274), .ZN(n11260) );
  NAND2_X1 U7367 ( .A1(n9443), .A2(n9442), .ZN(n11722) );
  AND2_X1 U7368 ( .A1(n11130), .A2(n11128), .ZN(n6486) );
  XNOR2_X1 U7369 ( .A(n11982), .B(n9093), .ZN(n12125) );
  OR2_X1 U7370 ( .A1(n8189), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8200) );
  NAND2_X1 U7371 ( .A1(n9396), .A2(n9395), .ZN(n11274) );
  NAND2_X2 U7372 ( .A1(n8692), .A2(n8691), .ZN(n11982) );
  INV_X1 U7373 ( .A(n6803), .ZN(n10754) );
  NAND2_X1 U7374 ( .A1(n6803), .A2(n7179), .ZN(n11003) );
  NAND2_X1 U7375 ( .A1(n8076), .A2(n7092), .ZN(n8093) );
  NAND2_X1 U7376 ( .A1(n8675), .A2(n8674), .ZN(n11979) );
  NAND2_X1 U7377 ( .A1(n8689), .A2(n8701), .ZN(n9939) );
  NAND2_X1 U7378 ( .A1(n8722), .A2(n8706), .ZN(n9945) );
  AND2_X1 U7379 ( .A1(n7180), .A2(n10756), .ZN(n6803) );
  OR2_X1 U7380 ( .A1(n8154), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8167) );
  NAND2_X1 U7381 ( .A1(n8639), .A2(n8638), .ZN(n14813) );
  NAND2_X1 U7382 ( .A1(n8593), .A2(n8592), .ZN(n10855) );
  NAND2_X1 U7383 ( .A1(n8658), .A2(n8657), .ZN(n11976) );
  NAND2_X1 U7384 ( .A1(n9345), .A2(n9344), .ZN(n10997) );
  NOR2_X1 U7385 ( .A1(n11806), .A2(n15195), .ZN(n12660) );
  NAND2_X1 U7386 ( .A1(n6965), .A2(n6963), .ZN(n8049) );
  NAND2_X1 U7387 ( .A1(n7514), .A2(n14417), .ZN(n14419) );
  OAI21_X1 U7388 ( .B1(n8653), .B2(n8652), .A(n8667), .ZN(n9927) );
  INV_X1 U7389 ( .A(n10657), .ZN(n15099) );
  AOI21_X1 U7390 ( .B1(n10690), .B2(n15208), .A(n10689), .ZN(n12334) );
  AND2_X1 U7391 ( .A1(n8299), .A2(n8297), .ZN(n10738) );
  OR2_X1 U7392 ( .A1(n9328), .A2(n9327), .ZN(n10657) );
  AND2_X1 U7393 ( .A1(n8628), .A2(n8627), .ZN(n10928) );
  NAND2_X1 U7394 ( .A1(n7184), .A2(n9786), .ZN(n10437) );
  INV_X1 U7395 ( .A(n9786), .ZN(n9785) );
  NAND2_X1 U7396 ( .A1(n8022), .A2(n8021), .ZN(n8038) );
  NAND2_X1 U7397 ( .A1(n7025), .A2(n7024), .ZN(n10631) );
  AOI21_X1 U7398 ( .B1(n10553), .B2(n10518), .A(n10519), .ZN(n10521) );
  INV_X1 U7399 ( .A(n7184), .ZN(n10336) );
  NAND4_X1 U7400 ( .A1(n9310), .A2(n9309), .A3(n9308), .A4(n9307), .ZN(n9780)
         );
  NAND4_X1 U7401 ( .A1(n9322), .A2(n9321), .A3(n9320), .A4(n9319), .ZN(n13088)
         );
  INV_X2 U7402 ( .A(n8215), .ZN(n8224) );
  OR2_X1 U7403 ( .A1(n10551), .A2(n7827), .ZN(n10553) );
  AND2_X1 U7404 ( .A1(n6766), .A2(n15067), .ZN(n7184) );
  NAND2_X2 U7405 ( .A1(n10200), .A2(n9267), .ZN(n12968) );
  AND2_X2 U7406 ( .A1(n10185), .A2(n11941), .ZN(n10220) );
  NAND4_X1 U7407 ( .A1(n9285), .A2(n9284), .A3(n9283), .A4(n9282), .ZN(n9784)
         );
  NAND4_X1 U7408 ( .A1(n9265), .A2(n9264), .A3(n9263), .A4(n9262), .ZN(n9782)
         );
  OR2_X1 U7409 ( .A1(n12088), .A2(n9901), .ZN(n8590) );
  INV_X1 U7410 ( .A(n6895), .ZN(n6894) );
  OR2_X1 U7411 ( .A1(n9286), .A2(n9930), .ZN(n9278) );
  BUF_X2 U7412 ( .A(n9306), .Z(n9749) );
  INV_X1 U7413 ( .A(n11941), .ZN(n11952) );
  NAND2_X1 U7414 ( .A1(n9154), .A2(n9153), .ZN(n10185) );
  CLKBUF_X3 U7415 ( .A(n8610), .Z(n9966) );
  INV_X1 U7416 ( .A(n9806), .ZN(n9267) );
  AND2_X1 U7417 ( .A1(n9242), .A2(n9241), .ZN(n9281) );
  XNOR2_X1 U7418 ( .A(n8250), .B(n8249), .ZN(n11084) );
  INV_X1 U7419 ( .A(n8549), .ZN(n8551) );
  XNOR2_X1 U7420 ( .A(n7785), .B(n7784), .ZN(n12223) );
  AND2_X2 U7421 ( .A1(n9747), .A2(n11328), .ZN(n9806) );
  AND2_X1 U7422 ( .A1(n9240), .A2(n13577), .ZN(n9540) );
  OR2_X1 U7423 ( .A1(n9744), .A2(n9896), .ZN(n9277) );
  INV_X1 U7424 ( .A(n9286), .ZN(n7011) );
  NAND2_X2 U7425 ( .A1(n7039), .A2(n7037), .ZN(n14331) );
  XNOR2_X1 U7426 ( .A(n9237), .B(n9236), .ZN(n13577) );
  XNOR2_X1 U7427 ( .A(n9235), .B(n9234), .ZN(n9240) );
  INV_X1 U7428 ( .A(n10379), .ZN(n12506) );
  INV_X1 U7429 ( .A(n8550), .ZN(n14325) );
  NAND2_X1 U7430 ( .A1(n7057), .A2(n7055), .ZN(n12100) );
  NAND2_X1 U7431 ( .A1(n7568), .A2(n7569), .ZN(n8549) );
  NAND2_X2 U7432 ( .A1(n9233), .A2(n9232), .ZN(n11328) );
  INV_X2 U7433 ( .A(n12889), .ZN(n12903) );
  INV_X2 U7434 ( .A(n14322), .ZN(n14327) );
  OR2_X1 U7435 ( .A1(n9068), .A2(n7498), .ZN(n7057) );
  NAND2_X1 U7436 ( .A1(n13569), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9235) );
  OAI21_X1 U7437 ( .B1(n9155), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9131) );
  OR2_X1 U7438 ( .A1(n8548), .A2(n8545), .ZN(n7569) );
  CLKBUF_X1 U7439 ( .A(n8435), .Z(n8441) );
  OR2_X1 U7440 ( .A1(n9228), .A2(n9208), .ZN(n9222) );
  NAND2_X1 U7441 ( .A1(n7163), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9225) );
  NAND2_X1 U7442 ( .A1(n9076), .A2(n9075), .ZN(n9155) );
  NAND2_X1 U7443 ( .A1(n14320), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8546) );
  MUX2_X1 U7444 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9074), .S(
        P1_IR_REG_22__SCAN_IN), .Z(n9077) );
  NAND2_X1 U7445 ( .A1(n7801), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7803) );
  OR2_X1 U7446 ( .A1(n9067), .A2(n8672), .ZN(n9071) );
  AND2_X1 U7447 ( .A1(n7840), .A2(n7857), .ZN(n10558) );
  AND2_X1 U7448 ( .A1(n7563), .A2(n8841), .ZN(n9133) );
  AND2_X1 U7449 ( .A1(n7917), .A2(n7916), .ZN(n7938) );
  NOR3_X1 U7450 ( .A1(n7446), .A2(n7780), .A3(n7346), .ZN(n7345) );
  AND2_X1 U7451 ( .A1(n9213), .A2(n6473), .ZN(n9199) );
  AND2_X1 U7452 ( .A1(n7588), .A2(n8541), .ZN(n6959) );
  AND2_X1 U7453 ( .A1(n6491), .A2(n7756), .ZN(n8841) );
  NAND2_X1 U7454 ( .A1(n7758), .A2(n7447), .ZN(n7446) );
  AND3_X1 U7455 ( .A1(n6477), .A2(n6480), .A3(n6479), .ZN(n9213) );
  AND2_X1 U7456 ( .A1(n6503), .A2(n8544), .ZN(n7588) );
  NAND2_X1 U7457 ( .A1(n6793), .A2(n7591), .ZN(n6704) );
  XOR2_X1 U7458 ( .A(n14402), .B(n14403), .Z(n14404) );
  AND3_X1 U7459 ( .A1(n7752), .A2(n8584), .A3(n8844), .ZN(n7496) );
  AND3_X1 U7460 ( .A1(n7397), .A2(n9276), .A3(n9288), .ZN(n9194) );
  AND2_X1 U7461 ( .A1(n7117), .A2(n9196), .ZN(n6477) );
  NAND3_X1 U7462 ( .A1(n8430), .A2(n8438), .A3(n7779), .ZN(n7780) );
  NAND2_X1 U7463 ( .A1(n15422), .A2(n7781), .ZN(n7346) );
  NOR2_X2 U7464 ( .A1(n15157), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n14403) );
  AND2_X1 U7465 ( .A1(n7774), .A2(n7698), .ZN(n6495) );
  CLKBUF_X1 U7466 ( .A(n10361), .Z(n7016) );
  AND4_X1 U7467 ( .A1(n7776), .A2(n7775), .A3(n7981), .A4(n7963), .ZN(n7762)
         );
  NOR2_X2 U7468 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n8584) );
  NOR2_X1 U7469 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n7776) );
  NOR2_X1 U7470 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), .ZN(
        n7775) );
  NOR2_X1 U7471 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n7752) );
  INV_X1 U7472 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n9476) );
  NOR2_X1 U7473 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6479) );
  NOR2_X1 U7474 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n6480) );
  INV_X1 U7475 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n9457) );
  INV_X4 U7476 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7477 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9288) );
  INV_X1 U7478 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9193) );
  INV_X1 U7479 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8248) );
  INV_X1 U7480 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n9323) );
  INV_X1 U7481 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8078) );
  INV_X1 U7482 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8624) );
  INV_X1 U7483 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9234) );
  NOR2_X1 U7484 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n8816) );
  INV_X1 U7485 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n9224) );
  NOR2_X1 U7486 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7772) );
  NOR2_X1 U7487 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n7771) );
  NOR2_X1 U7488 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n9219) );
  INV_X1 U7489 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n9221) );
  INV_X1 U7490 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9812) );
  NOR2_X1 U7491 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n10361) );
  INV_X4 U7492 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7493 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n14475) );
  NOR2_X2 U7494 ( .A1(n13288), .A2(n13282), .ZN(n13277) );
  NOR2_X2 U7495 ( .A1(n13312), .A2(n13476), .ZN(n7186) );
  NOR2_X2 U7496 ( .A1(n11003), .A2(n15048), .ZN(n11137) );
  NOR2_X2 U7497 ( .A1(n11726), .A2(n6478), .ZN(n6820) );
  AND2_X2 U7498 ( .A1(n11335), .A2(n11367), .ZN(n11620) );
  NOR2_X2 U7499 ( .A1(n11260), .A2(n11465), .ZN(n11335) );
  NOR2_X2 U7500 ( .A1(n13398), .A2(n13387), .ZN(n6819) );
  AND2_X2 U7501 ( .A1(n13438), .A2(n13525), .ZN(n13421) );
  NAND2_X2 U7502 ( .A1(n9825), .A2(n13584), .ZN(n9290) );
  XNOR2_X1 U7503 ( .A(n7371), .B(n9210), .ZN(n13584) );
  XNOR2_X2 U7504 ( .A(n9207), .B(n9206), .ZN(n9825) );
  AOI21_X2 U7505 ( .B1(n11921), .B2(n11920), .A(n6607), .ZN(n11923) );
  AOI21_X2 U7506 ( .B1(n13430), .B2(n13429), .A(n13237), .ZN(n13410) );
  OAI21_X2 U7507 ( .B1(n13371), .B2(n13370), .A(n6701), .ZN(n13353) );
  NAND2_X1 U7508 ( .A1(n13269), .A2(n14570), .ZN(n6484) );
  NAND2_X1 U7509 ( .A1(n13272), .A2(n13259), .ZN(n6485) );
  OAI21_X2 U7510 ( .B1(n14558), .B2(n6610), .A(n11879), .ZN(n11918) );
  OAI21_X2 U7511 ( .B1(n11878), .B2(n11877), .A(n6698), .ZN(n14558) );
  NOR2_X2 U7512 ( .A1(n10125), .A2(n10126), .ZN(n10136) );
  OAI21_X2 U7513 ( .B1(n10124), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10123), .ZN(
        n10125) );
  CLKBUF_X1 U7514 ( .A(n14334), .Z(n6487) );
  XNOR2_X1 U7515 ( .A(n8562), .B(n8561), .ZN(n14334) );
  INV_X4 U7516 ( .A(n13687), .ZN(n10183) );
  OAI21_X2 U7517 ( .B1(n13381), .B2(n13244), .A(n13246), .ZN(n13371) );
  XNOR2_X1 U7518 ( .A(n7803), .B(n7802), .ZN(n6488) );
  INV_X1 U7519 ( .A(n12539), .ZN(n10379) );
  AOI21_X2 U7520 ( .B1(n10137), .B2(P1_REG1_REG_6__SCAN_IN), .A(n10136), .ZN(
        n10140) );
  NOR2_X1 U7521 ( .A1(n10437), .A2(n10631), .ZN(n10641) );
  AOI21_X2 U7522 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(n10086), .A(n10306), .ZN(
        n10109) );
  AOI211_X2 U7523 ( .C1(n14146), .C2(n14181), .A(n13975), .B(n13974), .ZN(
        n13976) );
  AOI21_X2 U7524 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n10103), .A(n10107), .ZN(
        n10316) );
  XNOR2_X2 U7525 ( .A(n7059), .B(n6920), .ZN(n12085) );
  AND2_X1 U7526 ( .A1(n15090), .A2(n11328), .ZN(n6489) );
  NAND2_X4 U7527 ( .A1(n7824), .A2(n9676), .ZN(n7833) );
  INV_X1 U7528 ( .A(n12097), .ZN(n7493) );
  OR2_X1 U7529 ( .A1(n12792), .A2(n12667), .ZN(n8272) );
  OAI21_X1 U7530 ( .B1(n9053), .B2(n7619), .A(n7617), .ZN(n9742) );
  AOI21_X1 U7531 ( .B1(n7620), .B2(n7618), .A(n6666), .ZN(n7617) );
  INV_X1 U7532 ( .A(n7620), .ZN(n7619) );
  INV_X1 U7533 ( .A(n9056), .ZN(n7618) );
  OAI21_X1 U7534 ( .B1(n9005), .B2(n7610), .A(n7606), .ZN(n9041) );
  NOR2_X1 U7535 ( .A1(n7611), .A2(n7612), .ZN(n7610) );
  AND2_X1 U7536 ( .A1(n7609), .A2(n7607), .ZN(n7606) );
  NAND2_X1 U7537 ( .A1(n7611), .A2(n7259), .ZN(n7609) );
  NAND2_X1 U7538 ( .A1(n7594), .A2(n7592), .ZN(n8761) );
  AOI21_X1 U7539 ( .B1(n7595), .B2(n7597), .A(n7593), .ZN(n7592) );
  INV_X1 U7540 ( .A(n8738), .ZN(n7593) );
  NAND2_X1 U7541 ( .A1(n7283), .A2(n7282), .ZN(n7281) );
  INV_X1 U7542 ( .A(n12460), .ZN(n7282) );
  INV_X1 U7543 ( .A(n13081), .ZN(n11356) );
  NAND2_X1 U7544 ( .A1(n14546), .A2(n7628), .ZN(n7627) );
  INV_X1 U7545 ( .A(n7631), .ZN(n7630) );
  OR2_X1 U7546 ( .A1(n13375), .A2(n13247), .ZN(n6701) );
  INV_X1 U7547 ( .A(n13894), .ZN(n10801) );
  NAND2_X1 U7548 ( .A1(n9021), .A2(n7575), .ZN(n13984) );
  INV_X1 U7549 ( .A(n8727), .ZN(n12087) );
  NAND2_X1 U7550 ( .A1(n11977), .A2(n6856), .ZN(n6855) );
  INV_X1 U7551 ( .A(n11980), .ZN(n7481) );
  NAND2_X1 U7552 ( .A1(n6962), .A2(n6961), .ZN(n12023) );
  NAND2_X1 U7553 ( .A1(n13883), .A2(n6476), .ZN(n6961) );
  NAND2_X1 U7554 ( .A1(n14604), .A2(n12002), .ZN(n6962) );
  OAI22_X1 U7555 ( .A1(n7467), .A2(n6536), .B1(n6845), .B2(n12051), .ZN(n12054) );
  NAND2_X1 U7556 ( .A1(n12049), .A2(n12048), .ZN(n7467) );
  INV_X1 U7557 ( .A(n9628), .ZN(n7707) );
  INV_X1 U7558 ( .A(n8872), .ZN(n8875) );
  NAND2_X1 U7559 ( .A1(n12382), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7292) );
  AND2_X1 U7560 ( .A1(n9709), .A2(n9802), .ZN(n9769) );
  NAND2_X1 U7561 ( .A1(n8974), .A2(n8973), .ZN(n8988) );
  XNOR2_X1 U7562 ( .A(n10963), .B(n7086), .ZN(n11677) );
  NAND2_X1 U7563 ( .A1(n12252), .A2(n12183), .ZN(n12185) );
  INV_X1 U7564 ( .A(n12223), .ZN(n7789) );
  OR2_X1 U7565 ( .A1(n10521), .A2(n6594), .ZN(n6870) );
  NAND2_X1 U7566 ( .A1(n6870), .A2(n7218), .ZN(n7046) );
  OR2_X1 U7567 ( .A1(n10782), .A2(n10781), .ZN(n10783) );
  NAND2_X1 U7568 ( .A1(n6867), .A2(n6643), .ZN(n11392) );
  INV_X1 U7569 ( .A(n11390), .ZN(n6867) );
  NAND2_X1 U7570 ( .A1(n11756), .A2(n7292), .ZN(n7291) );
  NAND2_X1 U7571 ( .A1(n7048), .A2(n7047), .ZN(n7290) );
  AND2_X1 U7572 ( .A1(n11752), .A2(n7292), .ZN(n7047) );
  INV_X1 U7573 ( .A(n11753), .ZN(n7048) );
  NOR2_X1 U7574 ( .A1(n12612), .A2(n7682), .ZN(n7681) );
  INV_X1 U7575 ( .A(n8515), .ZN(n7682) );
  INV_X1 U7576 ( .A(n8516), .ZN(n7679) );
  NAND2_X1 U7577 ( .A1(n7693), .A2(n7692), .ZN(n12652) );
  NOR2_X1 U7578 ( .A1(n12654), .A2(n7694), .ZN(n7692) );
  OR2_X1 U7579 ( .A1(n12369), .A2(n11664), .ZN(n8322) );
  OR2_X1 U7580 ( .A1(n12371), .A2(n11647), .ZN(n8314) );
  OR2_X1 U7581 ( .A1(n12217), .A2(n12205), .ZN(n8403) );
  AND2_X1 U7582 ( .A1(n8051), .A2(n7342), .ZN(n8435) );
  NOR2_X1 U7583 ( .A1(n7446), .A2(n7343), .ZN(n7342) );
  NAND2_X1 U7584 ( .A1(n7344), .A2(n15422), .ZN(n7343) );
  INV_X1 U7585 ( .A(n7780), .ZN(n7344) );
  NAND2_X1 U7586 ( .A1(n6737), .A2(n7927), .ZN(n6736) );
  INV_X1 U7587 ( .A(n7924), .ZN(n6737) );
  INV_X1 U7588 ( .A(n7927), .ZN(n6738) );
  INV_X1 U7589 ( .A(n7947), .ZN(n7105) );
  INV_X1 U7590 ( .A(n13577), .ZN(n9241) );
  AND2_X1 U7591 ( .A1(n6790), .A2(n7064), .ZN(n13274) );
  AND2_X1 U7592 ( .A1(n7375), .A2(n7373), .ZN(n7064) );
  INV_X1 U7593 ( .A(n13275), .ZN(n7373) );
  INV_X1 U7594 ( .A(n13354), .ZN(n7362) );
  OR2_X1 U7595 ( .A1(n13533), .A2(n9792), .ZN(n13213) );
  NOR2_X1 U7596 ( .A1(n11883), .A2(n11920), .ZN(n6791) );
  NAND2_X1 U7597 ( .A1(n6558), .A2(n6492), .ZN(n7368) );
  NAND2_X1 U7598 ( .A1(n13357), .A2(n13494), .ZN(n13342) );
  AND2_X1 U7599 ( .A1(n9220), .A2(n9201), .ZN(n7661) );
  INV_X1 U7600 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n9198) );
  INV_X1 U7601 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n9197) );
  INV_X1 U7602 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9195) );
  OR2_X1 U7603 ( .A1(n13687), .A2(n14873), .ZN(n10798) );
  NAND2_X1 U7604 ( .A1(n13894), .A2(n10220), .ZN(n10799) );
  NAND2_X1 U7605 ( .A1(n7493), .A2(n12084), .ZN(n7491) );
  AND2_X1 U7606 ( .A1(n14708), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7168) );
  AND2_X1 U7607 ( .A1(n14030), .A2(n9111), .ZN(n7459) );
  NAND2_X1 U7608 ( .A1(n14074), .A2(n8938), .ZN(n14067) );
  INV_X1 U7609 ( .A(n14348), .ZN(n11944) );
  AND3_X1 U7610 ( .A1(n7563), .A2(n8841), .A3(n8541), .ZN(n8543) );
  NOR2_X1 U7611 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n9066) );
  NAND2_X1 U7612 ( .A1(n7234), .A2(SI_3_), .ZN(n8619) );
  NAND2_X1 U7613 ( .A1(n12884), .A2(n10709), .ZN(n6692) );
  AND2_X1 U7614 ( .A1(n7426), .A2(n7428), .ZN(n7424) );
  AOI21_X1 U7615 ( .B1(n8244), .B2(n8243), .A(n8242), .ZN(n8423) );
  AND2_X1 U7616 ( .A1(n11084), .A2(n9185), .ZN(n10709) );
  NAND2_X1 U7617 ( .A1(n7790), .A2(n7789), .ZN(n7846) );
  NAND2_X2 U7618 ( .A1(n7789), .A2(n12895), .ZN(n7844) );
  NAND2_X1 U7619 ( .A1(n7518), .A2(n12410), .ZN(n7517) );
  OR2_X1 U7620 ( .A1(n12457), .A2(n12458), .ZN(n7283) );
  NAND2_X1 U7621 ( .A1(n7225), .A2(n7224), .ZN(n7525) );
  INV_X1 U7622 ( .A(n12453), .ZN(n7224) );
  NAND2_X1 U7623 ( .A1(n7326), .A2(n7331), .ZN(n7320) );
  AOI21_X1 U7624 ( .B1(n12727), .B2(n7301), .A(n7300), .ZN(n7299) );
  INV_X1 U7625 ( .A(n8357), .ZN(n7300) );
  INV_X1 U7626 ( .A(n8356), .ZN(n7301) );
  NOR2_X1 U7627 ( .A1(n11314), .A2(n7676), .ZN(n7675) );
  INV_X1 U7628 ( .A(n8490), .ZN(n7676) );
  NAND2_X1 U7629 ( .A1(n7031), .A2(n7030), .ZN(n8219) );
  NAND2_X1 U7630 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n14333), .ZN(n7030) );
  NAND2_X1 U7631 ( .A1(n7032), .A2(n6679), .ZN(n7031) );
  AND2_X1 U7632 ( .A1(n8435), .A2(n6501), .ZN(n7799) );
  AOI21_X1 U7633 ( .B1(n8175), .B2(n8174), .A(n6967), .ZN(n8183) );
  AND2_X1 U7634 ( .A1(n14342), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6967) );
  AND2_X1 U7635 ( .A1(n7111), .A2(n6556), .ZN(n8128) );
  NAND2_X1 U7636 ( .A1(n8116), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7111) );
  NAND2_X1 U7637 ( .A1(n8049), .A2(n8050), .ZN(n7096) );
  OR2_X1 U7638 ( .A1(n7839), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n7857) );
  OAI21_X1 U7639 ( .B1(n7537), .B2(n7536), .A(n7534), .ZN(n7872) );
  AOI21_X1 U7640 ( .B1(n7535), .B2(n7854), .A(n6601), .ZN(n7534) );
  INV_X1 U7641 ( .A(n7836), .ZN(n7535) );
  NAND2_X1 U7642 ( .A1(n7835), .A2(n7834), .ZN(n7537) );
  INV_X1 U7643 ( .A(n6711), .ZN(n6710) );
  NAND2_X1 U7644 ( .A1(n11842), .A2(n6708), .ZN(n6707) );
  OAI21_X1 U7645 ( .B1(n7638), .B2(n6712), .A(n6713), .ZN(n6711) );
  OAI211_X1 U7646 ( .C1(n10827), .C2(n6719), .A(n11104), .B(n6718), .ZN(n11070) );
  INV_X1 U7647 ( .A(n11063), .ZN(n6719) );
  NAND2_X1 U7648 ( .A1(n7653), .A2(n11063), .ZN(n6718) );
  INV_X1 U7649 ( .A(n13074), .ZN(n13251) );
  NAND2_X1 U7650 ( .A1(n9247), .A2(n11328), .ZN(n9880) );
  AOI21_X1 U7651 ( .B1(n13324), .B2(n13323), .A(n7034), .ZN(n13320) );
  AND2_X1 U7652 ( .A1(n13488), .A2(n13251), .ZN(n7034) );
  NAND2_X1 U7653 ( .A1(n7361), .A2(n13250), .ZN(n7360) );
  INV_X1 U7654 ( .A(n7364), .ZN(n7361) );
  OAI21_X1 U7655 ( .B1(n13395), .B2(n6644), .A(n13219), .ZN(n13383) );
  NAND2_X1 U7656 ( .A1(n7395), .A2(n6562), .ZN(n7392) );
  INV_X1 U7657 ( .A(n9286), .ZN(n9743) );
  NAND2_X1 U7658 ( .A1(n7399), .A2(n7400), .ZN(n6792) );
  OAI21_X1 U7659 ( .B1(n11226), .B2(n7402), .A(n11329), .ZN(n7401) );
  AND2_X1 U7660 ( .A1(n15090), .A2(n11328), .ZN(n14562) );
  AND2_X1 U7661 ( .A1(n11439), .A2(n9248), .ZN(n15090) );
  OR2_X1 U7662 ( .A1(n9930), .A2(n9676), .ZN(n7751) );
  OR2_X1 U7663 ( .A1(n13786), .A2(n6975), .ZN(n6974) );
  AND2_X1 U7664 ( .A1(n13629), .A2(n13630), .ZN(n6975) );
  INV_X1 U7665 ( .A(n7767), .ZN(n7746) );
  XNOR2_X1 U7666 ( .A(n10266), .B(n11048), .ZN(n10794) );
  INV_X1 U7667 ( .A(n13615), .ZN(n13759) );
  NAND2_X1 U7668 ( .A1(n8614), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8563) );
  AND2_X1 U7669 ( .A1(n8549), .A2(n8550), .ZN(n8610) );
  NAND2_X1 U7670 ( .A1(n13998), .A2(n9116), .ZN(n13978) );
  NAND2_X1 U7671 ( .A1(n14019), .A2(n9003), .ZN(n13997) );
  NAND2_X1 U7672 ( .A1(n14043), .A2(n7582), .ZN(n7579) );
  NAND2_X1 U7673 ( .A1(n14102), .A2(n7464), .ZN(n14086) );
  AND2_X1 U7674 ( .A1(n14096), .A2(n12039), .ZN(n7464) );
  NAND2_X1 U7675 ( .A1(n14144), .A2(n12021), .ZN(n6879) );
  OR2_X1 U7676 ( .A1(n14597), .A2(n8806), .ZN(n12008) );
  NAND2_X1 U7677 ( .A1(n11442), .A2(n9098), .ZN(n11469) );
  NOR2_X2 U7678 ( .A1(n10943), .A2(n11982), .ZN(n11421) );
  OR2_X1 U7679 ( .A1(n10907), .A2(n9086), .ZN(n9089) );
  NOR2_X1 U7680 ( .A1(n7574), .A2(n8629), .ZN(n7573) );
  INV_X1 U7681 ( .A(n8608), .ZN(n7574) );
  NAND2_X1 U7682 ( .A1(n12090), .A2(n12089), .ZN(n13942) );
  NAND2_X1 U7683 ( .A1(n8705), .A2(n8704), .ZN(n8722) );
  OAI21_X1 U7684 ( .B1(n8670), .B2(n6896), .A(n8687), .ZN(n6895) );
  INV_X1 U7685 ( .A(n8683), .ZN(n6896) );
  NOR2_X1 U7686 ( .A1(n14657), .A2(n6759), .ZN(n14439) );
  NOR2_X1 U7687 ( .A1(n14656), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6759) );
  AOI22_X1 U7688 ( .A1(n14384), .A2(n14383), .B1(P1_ADDR_REG_14__SCAN_IN), 
        .B2(n14382), .ZN(n14440) );
  NOR2_X1 U7689 ( .A1(n12426), .A2(n12427), .ZN(n12451) );
  NOR2_X1 U7690 ( .A1(n12481), .A2(n12717), .ZN(n12502) );
  NAND2_X1 U7691 ( .A1(n7528), .A2(n7527), .ZN(n7526) );
  INV_X1 U7692 ( .A(n12523), .ZN(n7527) );
  NAND2_X1 U7693 ( .A1(n12524), .A2(n15173), .ZN(n7528) );
  AOI21_X1 U7694 ( .B1(n9166), .B2(n6802), .A(n8524), .ZN(n12563) );
  NAND2_X1 U7695 ( .A1(n6734), .A2(n6733), .ZN(n12769) );
  INV_X1 U7696 ( .A(n6993), .ZN(n6734) );
  NAND2_X1 U7697 ( .A1(n12569), .A2(n14499), .ZN(n6733) );
  NAND2_X1 U7698 ( .A1(n11513), .A2(n11512), .ZN(n11654) );
  INV_X1 U7699 ( .A(n13204), .ZN(n13453) );
  NAND2_X1 U7700 ( .A1(n9027), .A2(n9026), .ZN(n13988) );
  NOR2_X1 U7701 ( .A1(n13787), .A2(n13788), .ZN(n13786) );
  INV_X1 U7702 ( .A(n9317), .ZN(n7715) );
  INV_X1 U7703 ( .A(n9316), .ZN(n7713) );
  INV_X1 U7704 ( .A(n9341), .ZN(n7140) );
  NOR2_X1 U7705 ( .A1(n6544), .A2(n7140), .ZN(n7139) );
  NAND2_X1 U7706 ( .A1(n7021), .A2(n7020), .ZN(n11971) );
  OR2_X1 U7707 ( .A1(n7478), .A2(n11974), .ZN(n7014) );
  INV_X1 U7708 ( .A(n11973), .ZN(n7478) );
  INV_X1 U7709 ( .A(n11981), .ZN(n7480) );
  NAND2_X1 U7710 ( .A1(n6539), .A2(n6851), .ZN(n6853) );
  NOR2_X1 U7711 ( .A1(n6579), .A2(n6852), .ZN(n6851) );
  INV_X1 U7712 ( .A(n6855), .ZN(n6852) );
  NAND2_X1 U7713 ( .A1(n11992), .A2(n7476), .ZN(n7475) );
  NOR2_X1 U7714 ( .A1(n7476), .A2(n11992), .ZN(n7477) );
  AOI21_X1 U7715 ( .B1(n6500), .B2(n7151), .A(n6586), .ZN(n7149) );
  OR2_X1 U7716 ( .A1(n12115), .A2(n14264), .ZN(n12025) );
  NAND2_X1 U7717 ( .A1(n12003), .A2(n6981), .ZN(n6980) );
  AOI21_X1 U7718 ( .B1(n12002), .B2(n12022), .A(n12027), .ZN(n12031) );
  INV_X1 U7719 ( .A(n12035), .ZN(n7488) );
  INV_X1 U7720 ( .A(n6846), .ZN(n6850) );
  OAI21_X1 U7721 ( .B1(n12137), .B2(n12038), .A(n12041), .ZN(n6846) );
  NAND2_X1 U7722 ( .A1(n12137), .A2(n12041), .ZN(n6847) );
  NAND2_X1 U7723 ( .A1(n7022), .A2(n6850), .ZN(n6849) );
  AOI21_X1 U7724 ( .B1(n9547), .B2(n9546), .A(n9545), .ZN(n9549) );
  AOI21_X1 U7725 ( .B1(n12054), .B2(n12053), .A(n12052), .ZN(n7469) );
  NAND2_X1 U7726 ( .A1(n12056), .A2(n6864), .ZN(n6863) );
  INV_X1 U7727 ( .A(n12055), .ZN(n6864) );
  INV_X1 U7728 ( .A(n9582), .ZN(n7146) );
  NAND2_X1 U7729 ( .A1(n12065), .A2(n6858), .ZN(n6857) );
  NAND2_X1 U7730 ( .A1(n12066), .A2(n6861), .ZN(n6860) );
  INV_X1 U7731 ( .A(n9100), .ZN(n7454) );
  AND2_X1 U7732 ( .A1(n7600), .A2(n7247), .ZN(n7246) );
  NAND2_X1 U7733 ( .A1(n8760), .A2(n8759), .ZN(n7247) );
  INV_X1 U7734 ( .A(n11688), .ZN(n6682) );
  OR2_X1 U7735 ( .A1(n8150), .A2(n7549), .ZN(n7544) );
  NAND2_X1 U7736 ( .A1(n11796), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6750) );
  INV_X1 U7737 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n6817) );
  NAND2_X1 U7738 ( .A1(n6636), .A2(n7707), .ZN(n7704) );
  NOR2_X1 U7739 ( .A1(n6636), .A2(n7707), .ZN(n7706) );
  OAI21_X1 U7740 ( .B1(n14398), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6593), .ZN(
        n7499) );
  AND2_X1 U7741 ( .A1(n12244), .A2(n7433), .ZN(n7432) );
  OR2_X1 U7742 ( .A1(n12325), .A2(n7434), .ZN(n7433) );
  INV_X1 U7743 ( .A(n7340), .ZN(n7334) );
  NAND2_X1 U7744 ( .A1(n6604), .A2(n8393), .ZN(n7337) );
  AND2_X1 U7745 ( .A1(n8399), .A2(n8241), .ZN(n7532) );
  NAND2_X1 U7746 ( .A1(n7519), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7194) );
  NAND2_X1 U7747 ( .A1(n7279), .A2(n15174), .ZN(n7277) );
  INV_X1 U7748 ( .A(n11392), .ZN(n7279) );
  NOR2_X1 U7749 ( .A1(n7289), .A2(n12414), .ZN(n7288) );
  INV_X1 U7750 ( .A(n7291), .ZN(n7289) );
  NOR2_X1 U7751 ( .A1(n12618), .A2(n12626), .ZN(n8516) );
  AND2_X1 U7752 ( .A1(n7320), .A2(n12621), .ZN(n7317) );
  OAI22_X1 U7753 ( .A1(n8511), .A2(n7695), .B1(n12855), .B2(n12679), .ZN(n7694) );
  INV_X1 U7754 ( .A(n8509), .ZN(n7695) );
  INV_X1 U7755 ( .A(n8505), .ZN(n7670) );
  INV_X1 U7756 ( .A(n7671), .ZN(n7666) );
  INV_X1 U7757 ( .A(n8500), .ZN(n7690) );
  INV_X1 U7758 ( .A(n7305), .ZN(n7304) );
  NOR2_X1 U7759 ( .A1(n11799), .A2(n7306), .ZN(n7305) );
  INV_X1 U7760 ( .A(n7952), .ZN(n7306) );
  OR2_X1 U7761 ( .A1(n12372), .A2(n11210), .ZN(n8305) );
  OR2_X1 U7762 ( .A1(n15201), .A2(n10724), .ZN(n8291) );
  INV_X1 U7763 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7447) );
  INV_X1 U7764 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8430) );
  NOR2_X1 U7765 ( .A1(n8063), .A2(n7446), .ZN(n7347) );
  NOR2_X1 U7766 ( .A1(n8247), .A2(P3_IR_REG_19__SCAN_IN), .ZN(n8251) );
  NOR2_X1 U7767 ( .A1(n8063), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n7087) );
  INV_X1 U7768 ( .A(n7094), .ZN(n6747) );
  INV_X1 U7769 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7976) );
  NAND2_X1 U7770 ( .A1(n7975), .A2(n7974), .ZN(n7978) );
  INV_X1 U7771 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7962) );
  INV_X1 U7772 ( .A(n7104), .ZN(n7103) );
  OAI21_X1 U7773 ( .B1(n7944), .B2(n7105), .A(n7960), .ZN(n7104) );
  INV_X1 U7774 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7926) );
  OAI21_X1 U7775 ( .B1(n7269), .B2(n7016), .A(n7267), .ZN(n7266) );
  NAND2_X1 U7776 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7269) );
  NAND2_X1 U7777 ( .A1(n7929), .A2(n7268), .ZN(n7267) );
  NOR2_X1 U7778 ( .A1(n6712), .A2(n6709), .ZN(n6708) );
  INV_X1 U7779 ( .A(n7640), .ZN(n6709) );
  AND2_X1 U7780 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n9633), .ZN(n9643) );
  NAND2_X1 U7781 ( .A1(n9778), .A2(n6554), .ZN(n7130) );
  AND2_X1 U7782 ( .A1(n9769), .A2(n9734), .ZN(n7134) );
  NOR2_X1 U7783 ( .A1(n6971), .A2(n9768), .ZN(n9773) );
  INV_X1 U7784 ( .A(n7130), .ZN(n7129) );
  INV_X1 U7785 ( .A(n7134), .ZN(n7126) );
  OAI21_X1 U7786 ( .B1(n7131), .B2(n7129), .A(n11328), .ZN(n7128) );
  AOI21_X1 U7787 ( .B1(n7377), .B2(n7376), .A(n6603), .ZN(n7375) );
  INV_X1 U7788 ( .A(n7381), .ZN(n7376) );
  NAND2_X1 U7789 ( .A1(n7027), .A2(n7377), .ZN(n6790) );
  NAND2_X1 U7790 ( .A1(n13476), .A2(n13257), .ZN(n7384) );
  INV_X1 U7791 ( .A(n13227), .ZN(n13258) );
  NOR2_X1 U7792 ( .A1(n7394), .A2(n13211), .ZN(n7393) );
  INV_X1 U7793 ( .A(n11933), .ZN(n7394) );
  NOR2_X1 U7794 ( .A1(n6564), .A2(n6784), .ZN(n6783) );
  INV_X1 U7795 ( .A(n11723), .ZN(n6784) );
  NOR2_X1 U7796 ( .A1(n11126), .A2(n6772), .ZN(n6771) );
  INV_X1 U7797 ( .A(n10998), .ZN(n6772) );
  INV_X1 U7798 ( .A(n10994), .ZN(n6768) );
  OR2_X1 U7799 ( .A1(n9379), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n9381) );
  OR2_X1 U7800 ( .A1(n9381), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n9407) );
  INV_X1 U7801 ( .A(n13713), .ZN(n7729) );
  INV_X1 U7802 ( .A(n13685), .ZN(n6956) );
  INV_X1 U7803 ( .A(n13692), .ZN(n7733) );
  AND2_X1 U7804 ( .A1(n13729), .A2(n7732), .ZN(n7731) );
  OR2_X1 U7805 ( .A1(n13841), .A2(n7733), .ZN(n7732) );
  INV_X1 U7806 ( .A(n11946), .ZN(n11947) );
  AOI21_X1 U7807 ( .B1(n6985), .B2(n6905), .A(n6553), .ZN(n6904) );
  INV_X1 U7808 ( .A(n9118), .ZN(n6905) );
  AND2_X1 U7809 ( .A1(n7226), .A2(n6826), .ZN(n9122) );
  INV_X1 U7810 ( .A(n14288), .ZN(n6826) );
  NOR2_X1 U7811 ( .A1(n14001), .A2(n13988), .ZN(n7226) );
  NOR2_X1 U7812 ( .A1(n9109), .A2(n6913), .ZN(n6912) );
  NAND2_X1 U7813 ( .A1(n6914), .A2(n9106), .ZN(n6913) );
  INV_X1 U7814 ( .A(n9108), .ZN(n6914) );
  NOR2_X1 U7815 ( .A1(n14073), .A2(n9108), .ZN(n6916) );
  NOR2_X1 U7816 ( .A1(n14264), .A2(n14150), .ZN(n12115) );
  INV_X1 U7817 ( .A(n6909), .ZN(n6908) );
  OAI21_X1 U7818 ( .B1(n12133), .B2(n6910), .A(n12134), .ZN(n6909) );
  OR2_X1 U7819 ( .A1(n11856), .A2(n6910), .ZN(n6907) );
  INV_X1 U7820 ( .A(n12125), .ZN(n7461) );
  OR2_X1 U7821 ( .A1(n7463), .A2(n12126), .ZN(n6919) );
  INV_X1 U7822 ( .A(n9094), .ZN(n7463) );
  NAND2_X1 U7823 ( .A1(n14348), .A2(n14138), .ZN(n11945) );
  AND2_X1 U7824 ( .A1(n11945), .A2(n11952), .ZN(n11048) );
  NAND2_X1 U7825 ( .A1(n6911), .A2(n7450), .ZN(n14114) );
  INV_X1 U7826 ( .A(n7451), .ZN(n7450) );
  NAND2_X1 U7827 ( .A1(n6907), .A2(n6580), .ZN(n6911) );
  OAI21_X1 U7828 ( .B1(n6532), .B2(n7452), .A(n9101), .ZN(n7451) );
  OR2_X1 U7829 ( .A1(n11558), .A2(n14630), .ZN(n11556) );
  NAND2_X1 U7830 ( .A1(n11421), .A2(n6831), .ZN(n11558) );
  AND2_X1 U7831 ( .A1(n14787), .A2(n14797), .ZN(n6831) );
  XNOR2_X1 U7832 ( .A(n8988), .B(n11824), .ZN(n8987) );
  AND2_X1 U7833 ( .A1(n8899), .A2(n8898), .ZN(n9067) );
  OAI21_X1 U7834 ( .B1(n8874), .B2(n8873), .A(n6528), .ZN(n8890) );
  AND2_X1 U7835 ( .A1(n7253), .A2(n7250), .ZN(n7249) );
  INV_X1 U7836 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8540) );
  NOR2_X1 U7837 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n7562) );
  NOR2_X1 U7838 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n7561) );
  OAI21_X1 U7839 ( .B1(n8761), .B2(n8760), .A(n8759), .ZN(n8773) );
  INV_X1 U7840 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8707) );
  NAND2_X1 U7841 ( .A1(n7236), .A2(n6705), .ZN(n8671) );
  AND2_X1 U7842 ( .A1(n7235), .A2(n8666), .ZN(n6705) );
  OAI21_X1 U7843 ( .B1(n9211), .B2(n6883), .A(n6882), .ZN(n8650) );
  NAND2_X1 U7844 ( .A1(n9211), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6882) );
  OAI21_X1 U7845 ( .B1(n9211), .B2(n6881), .A(n6880), .ZN(n8632) );
  NAND2_X1 U7846 ( .A1(n9211), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n6880) );
  NAND2_X1 U7847 ( .A1(n6809), .A2(SI_4_), .ZN(n8630) );
  NAND2_X1 U7848 ( .A1(n8580), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7065) );
  NAND2_X1 U7849 ( .A1(n6755), .A2(n6754), .ZN(n14352) );
  NAND2_X1 U7850 ( .A1(n6548), .A2(n14401), .ZN(n6754) );
  XNOR2_X1 U7851 ( .A(n7499), .B(P3_ADDR_REG_5__SCAN_IN), .ZN(n14411) );
  INV_X1 U7852 ( .A(n7499), .ZN(n14358) );
  OAI22_X1 U7853 ( .A1(n14415), .A2(n14364), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n14363), .ZN(n14365) );
  INV_X1 U7854 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14363) );
  AOI22_X1 U7855 ( .A1(P3_ADDR_REG_12__SCAN_IN), .A2(n14379), .B1(n14430), 
        .B2(n14378), .ZN(n14433) );
  NAND2_X1 U7856 ( .A1(n6689), .A2(n6572), .ZN(n12252) );
  INV_X1 U7857 ( .A(n12255), .ZN(n7070) );
  INV_X1 U7858 ( .A(n11211), .ZN(n7426) );
  INV_X1 U7859 ( .A(n10965), .ZN(n7425) );
  AND2_X1 U7860 ( .A1(n12273), .A2(n7419), .ZN(n7418) );
  NAND2_X1 U7861 ( .A1(n7420), .A2(n12169), .ZN(n7419) );
  INV_X1 U7862 ( .A(n12167), .ZN(n7420) );
  NAND2_X1 U7863 ( .A1(n7429), .A2(n10960), .ZN(n7428) );
  NOR2_X1 U7864 ( .A1(n11686), .A2(n11685), .ZN(n11687) );
  NAND2_X1 U7865 ( .A1(n12281), .A2(n12280), .ZN(n12174) );
  INV_X1 U7866 ( .A(n10709), .ZN(n8472) );
  NAND2_X1 U7867 ( .A1(n7532), .A2(n8402), .ZN(n8255) );
  AND4_X1 U7868 ( .A1(n8182), .A2(n8181), .A3(n8180), .A4(n8179), .ZN(n8517)
         );
  NAND2_X1 U7869 ( .A1(n6872), .A2(n10362), .ZN(n10531) );
  NAND2_X1 U7870 ( .A1(n10369), .A2(n10370), .ZN(n10401) );
  NAND2_X1 U7871 ( .A1(n7046), .A2(n7045), .ZN(n10415) );
  INV_X1 U7872 ( .A(n6870), .ZN(n10414) );
  OR2_X1 U7873 ( .A1(n10769), .A2(n10768), .ZN(n10770) );
  NAND2_X1 U7874 ( .A1(n6869), .A2(n6868), .ZN(n11390) );
  NAND2_X1 U7875 ( .A1(n11151), .A2(n7287), .ZN(n6869) );
  AND2_X1 U7876 ( .A1(n6671), .A2(n7285), .ZN(n11150) );
  NAND2_X1 U7877 ( .A1(n7277), .A2(n11391), .ZN(n15161) );
  OR2_X1 U7878 ( .A1(n11384), .A2(n11383), .ZN(n11386) );
  AND3_X1 U7879 ( .A1(n7198), .A2(n11385), .A3(P3_REG1_REG_9__SCAN_IN), .ZN(
        n15158) );
  AND3_X1 U7880 ( .A1(n7277), .A2(n11391), .A3(P3_REG2_REG_9__SCAN_IN), .ZN(
        n15160) );
  NAND2_X1 U7881 ( .A1(n7200), .A2(n15174), .ZN(n7198) );
  INV_X1 U7882 ( .A(n11386), .ZN(n7200) );
  OR2_X1 U7883 ( .A1(n11573), .A2(n11572), .ZN(n11574) );
  OR2_X1 U7884 ( .A1(n12379), .A2(n12378), .ZN(n12380) );
  OR2_X1 U7885 ( .A1(n12522), .A2(n12521), .ZN(n7531) );
  OAI21_X1 U7886 ( .B1(n12608), .B2(n7098), .A(n7097), .ZN(n12578) );
  NAND2_X1 U7887 ( .A1(n6609), .A2(n8264), .ZN(n7097) );
  NAND2_X1 U7888 ( .A1(n8264), .A2(n12612), .ZN(n7098) );
  AOI21_X1 U7889 ( .B1(n7677), .B2(n6799), .A(n6591), .ZN(n6798) );
  NAND2_X1 U7890 ( .A1(n12623), .A2(n7681), .ZN(n7680) );
  INV_X1 U7891 ( .A(n7680), .ZN(n12610) );
  OR2_X1 U7892 ( .A1(n8374), .A2(n8270), .ZN(n12637) );
  NAND2_X1 U7893 ( .A1(n7330), .A2(n8271), .ZN(n7116) );
  NOR2_X1 U7894 ( .A1(n12670), .A2(n8126), .ZN(n7329) );
  INV_X1 U7895 ( .A(n8271), .ZN(n8126) );
  NAND2_X1 U7896 ( .A1(n12688), .A2(n6571), .ZN(n7693) );
  NOR2_X1 U7897 ( .A1(n8511), .A2(n8404), .ZN(n7696) );
  INV_X1 U7898 ( .A(n8273), .ZN(n7330) );
  AOI21_X1 U7899 ( .B1(n8105), .B2(n8104), .A(n8103), .ZN(n12671) );
  AOI21_X1 U7900 ( .B1(n7299), .B2(n12722), .A(n7298), .ZN(n7297) );
  INV_X1 U7901 ( .A(n12711), .ZN(n7298) );
  AND2_X1 U7902 ( .A1(n8277), .A2(n12696), .ZN(n12711) );
  INV_X1 U7903 ( .A(n12691), .ZN(n12725) );
  NAND2_X1 U7904 ( .A1(n12736), .A2(n8504), .ZN(n8506) );
  OAI21_X1 U7905 ( .B1(n8003), .B2(n7311), .A(n7308), .ZN(n12742) );
  INV_X1 U7906 ( .A(n7312), .ZN(n7311) );
  AOI21_X1 U7907 ( .B1(n7312), .B2(n7310), .A(n7309), .ZN(n7308) );
  NOR2_X1 U7908 ( .A1(n6515), .A2(n8347), .ZN(n7312) );
  INV_X1 U7909 ( .A(n8418), .ZN(n12741) );
  NOR2_X1 U7910 ( .A1(n8346), .A2(n7315), .ZN(n7314) );
  INV_X1 U7911 ( .A(n8341), .ZN(n7315) );
  NOR2_X1 U7912 ( .A1(n11485), .A2(n6807), .ZN(n6806) );
  INV_X1 U7913 ( .A(n8493), .ZN(n6807) );
  AND2_X1 U7914 ( .A1(n8530), .A2(n9183), .ZN(n12586) );
  NAND2_X1 U7915 ( .A1(n11287), .A2(n11599), .ZN(n11286) );
  AND2_X1 U7916 ( .A1(n11242), .A2(n8491), .ZN(n7673) );
  NAND2_X1 U7917 ( .A1(n10740), .A2(n8489), .ZN(n10841) );
  NAND2_X1 U7918 ( .A1(n10841), .A2(n10840), .ZN(n10839) );
  INV_X1 U7919 ( .A(n11084), .ZN(n11310) );
  NAND2_X1 U7920 ( .A1(n10705), .A2(n8307), .ZN(n15183) );
  OR2_X1 U7921 ( .A1(n15202), .A2(n10694), .ZN(n15198) );
  AND3_X1 U7922 ( .A1(n8002), .A2(n8001), .A3(n8000), .ZN(n14520) );
  NOR2_X1 U7923 ( .A1(n9179), .A2(n8476), .ZN(n10692) );
  AND2_X1 U7924 ( .A1(n10673), .A2(n12883), .ZN(n10688) );
  NAND2_X1 U7925 ( .A1(n11200), .A2(n11084), .ZN(n15195) );
  AND2_X1 U7926 ( .A1(n8522), .A2(n8307), .ZN(n15200) );
  AOI21_X1 U7927 ( .B1(n8455), .B2(n12904), .A(n7017), .ZN(n10033) );
  XNOR2_X1 U7928 ( .A(n7787), .B(n7786), .ZN(n7788) );
  NAND2_X1 U7929 ( .A1(n12885), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7787) );
  AOI21_X1 U7930 ( .B1(n8195), .B2(n8196), .A(n7543), .ZN(n8207) );
  AND2_X1 U7931 ( .A1(n14336), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7543) );
  NAND2_X1 U7932 ( .A1(n6978), .A2(n6977), .ZN(n8437) );
  NAND2_X1 U7933 ( .A1(n7929), .A2(n7781), .ZN(n6977) );
  NAND2_X1 U7934 ( .A1(n8161), .A2(n14346), .ZN(n8162) );
  NAND2_X1 U7935 ( .A1(n7347), .A2(n8430), .ZN(n8444) );
  XNOR2_X1 U7936 ( .A(n8160), .B(n13598), .ZN(n8161) );
  NOR2_X1 U7937 ( .A1(n8140), .A2(n7548), .ZN(n7547) );
  INV_X1 U7938 ( .A(n7550), .ZN(n7548) );
  NAND2_X1 U7939 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n11438), .ZN(n7550) );
  XNOR2_X1 U7940 ( .A(n8115), .B(n11327), .ZN(n8116) );
  NAND2_X1 U7941 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n7090), .ZN(n7089) );
  NAND2_X1 U7942 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n7093), .ZN(n7092) );
  NAND2_X1 U7943 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n7095), .ZN(n7094) );
  NAND2_X1 U7944 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n6964), .ZN(n6963) );
  NAND2_X1 U7945 ( .A1(n8038), .A2(n8039), .ZN(n6965) );
  INV_X1 U7946 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6964) );
  INV_X1 U7947 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7996) );
  NAND2_X1 U7948 ( .A1(n7978), .A2(n7977), .ZN(n7995) );
  XNOR2_X1 U7949 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n7994) );
  XNOR2_X1 U7950 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n7960) );
  INV_X1 U7951 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7946) );
  XNOR2_X1 U7952 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n7944) );
  NAND2_X1 U7953 ( .A1(n6735), .A2(n7927), .ZN(n7945) );
  NAND2_X1 U7954 ( .A1(n7925), .A2(n7924), .ZN(n6735) );
  NAND2_X1 U7955 ( .A1(n6725), .A2(n6723), .ZN(n7907) );
  AOI21_X1 U7956 ( .B1(n6727), .B2(n6724), .A(n6509), .ZN(n6723) );
  OR2_X1 U7957 ( .A1(n7872), .A2(n6726), .ZN(n6725) );
  CLKBUF_X1 U7958 ( .A(n7892), .Z(n7893) );
  NAND2_X1 U7959 ( .A1(n7820), .A2(n7821), .ZN(n7088) );
  NOR2_X1 U7960 ( .A1(n7633), .A2(n11831), .ZN(n7628) );
  AND2_X1 U7961 ( .A1(n11832), .A2(n7634), .ZN(n7633) );
  NAND2_X1 U7962 ( .A1(n11655), .A2(n7635), .ZN(n7634) );
  INV_X1 U7963 ( .A(n11653), .ZN(n7635) );
  NAND2_X1 U7964 ( .A1(n13027), .A2(n6992), .ZN(n12923) );
  OR2_X1 U7965 ( .A1(n12920), .A2(n6527), .ZN(n6992) );
  NOR2_X1 U7966 ( .A1(n7643), .A2(n12999), .ZN(n7642) );
  AND2_X1 U7967 ( .A1(n12906), .A2(n11843), .ZN(n7643) );
  NAND2_X1 U7968 ( .A1(n12979), .A2(n6720), .ZN(n12919) );
  NAND2_X1 U7969 ( .A1(n12917), .A2(n6721), .ZN(n6720) );
  INV_X1 U7970 ( .A(n12918), .ZN(n6721) );
  OR2_X1 U7971 ( .A1(n11461), .A2(n11462), .ZN(n11459) );
  XNOR2_X1 U7972 ( .A(n9835), .B(n9837), .ZN(n7624) );
  INV_X1 U7973 ( .A(n9248), .ZN(n9834) );
  NAND2_X1 U7974 ( .A1(n9281), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9273) );
  NAND2_X1 U7975 ( .A1(n6525), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9263) );
  AND2_X1 U7976 ( .A1(n9241), .A2(n9240), .ZN(n9306) );
  NAND2_X1 U7977 ( .A1(n9681), .A2(n9680), .ZN(n13201) );
  NAND2_X1 U7978 ( .A1(n6790), .A2(n7375), .ZN(n6788) );
  AND2_X1 U7979 ( .A1(n13259), .A2(n9779), .ZN(n13275) );
  NAND2_X1 U7980 ( .A1(n13476), .A2(n13256), .ZN(n7350) );
  NOR2_X1 U7981 ( .A1(n13476), .A2(n13256), .ZN(n7349) );
  INV_X1 U7982 ( .A(n13301), .ZN(n6700) );
  NOR2_X1 U7983 ( .A1(n7374), .A2(n7382), .ZN(n7381) );
  INV_X1 U7984 ( .A(n7384), .ZN(n7382) );
  NAND2_X1 U7985 ( .A1(n7264), .A2(n7384), .ZN(n7380) );
  NAND2_X1 U7986 ( .A1(n13300), .A2(n7265), .ZN(n7264) );
  NAND2_X1 U7987 ( .A1(n7385), .A2(n13319), .ZN(n7265) );
  AND2_X1 U7988 ( .A1(n13328), .A2(n7356), .ZN(n7355) );
  NAND2_X1 U7989 ( .A1(n7359), .A2(n7357), .ZN(n7356) );
  OAI21_X1 U7990 ( .B1(n6778), .B2(n6497), .A(n6774), .ZN(n13324) );
  INV_X1 U7991 ( .A(n6775), .ZN(n6774) );
  OAI21_X1 U7992 ( .B1(n6776), .B2(n6497), .A(n6560), .ZN(n6775) );
  OR2_X1 U7993 ( .A1(n13354), .A2(n6777), .ZN(n6776) );
  INV_X1 U7994 ( .A(n6780), .ZN(n6777) );
  NAND2_X1 U7995 ( .A1(n13223), .A2(n6779), .ZN(n6778) );
  AND2_X1 U7996 ( .A1(n6780), .A2(n7396), .ZN(n6779) );
  OR2_X1 U7997 ( .A1(n13375), .A2(n13224), .ZN(n7396) );
  NAND2_X1 U7998 ( .A1(n6819), .A2(n6818), .ZN(n13373) );
  NAND2_X1 U7999 ( .A1(n13414), .A2(n13214), .ZN(n13217) );
  NAND2_X1 U8000 ( .A1(n11934), .A2(n7393), .ZN(n7388) );
  INV_X1 U8001 ( .A(n7392), .ZN(n7391) );
  OR2_X1 U8002 ( .A1(n9464), .A2(n9238), .ZN(n9481) );
  INV_X1 U8003 ( .A(n6791), .ZN(n11934) );
  OR2_X1 U8004 ( .A1(n14573), .A2(n13078), .ZN(n6698) );
  OR2_X1 U8005 ( .A1(n11615), .A2(n11718), .ZN(n11724) );
  NAND2_X1 U8006 ( .A1(n6792), .A2(n6576), .ZN(n11614) );
  OAI22_X1 U8007 ( .A1(n11224), .A2(n11223), .B1(n15115), .B2(n13084), .ZN(
        n11225) );
  NAND2_X1 U8008 ( .A1(n7403), .A2(n11226), .ZN(n11258) );
  INV_X1 U8009 ( .A(n11225), .ZN(n7403) );
  NAND2_X1 U8010 ( .A1(n15115), .A2(n11137), .ZN(n11229) );
  XNOR2_X1 U8011 ( .A(n11222), .B(n13084), .ZN(n11131) );
  OAI22_X1 U8012 ( .A1(n10991), .A2(n10994), .B1(n10997), .B2(n13086), .ZN(
        n10993) );
  OAI21_X1 U8013 ( .B1(n10644), .B2(n7406), .A(n10757), .ZN(n7405) );
  INV_X1 U8014 ( .A(n10664), .ZN(n7180) );
  XNOR2_X1 U8015 ( .A(n13088), .B(n15099), .ZN(n10654) );
  NAND2_X1 U8016 ( .A1(n10331), .A2(n10330), .ZN(n10333) );
  OR2_X1 U8017 ( .A1(n9782), .A2(n15067), .ZN(n10327) );
  NAND2_X1 U8018 ( .A1(n9711), .A2(n9710), .ZN(n13469) );
  NAND2_X1 U8019 ( .A1(n9427), .A2(n9426), .ZN(n15122) );
  OR2_X1 U8020 ( .A1(n9290), .A2(n10006), .ZN(n7760) );
  AND2_X1 U8021 ( .A1(n13586), .A2(n9856), .ZN(n15077) );
  NAND2_X1 U8022 ( .A1(n9818), .A2(n9814), .ZN(n9996) );
  AND2_X1 U8023 ( .A1(n9210), .A2(n9206), .ZN(n7721) );
  INV_X1 U8024 ( .A(n7407), .ZN(n7370) );
  MUX2_X1 U8025 ( .A(n9227), .B(P2_IR_REG_31__SCAN_IN), .S(n9226), .Z(n9229)
         );
  NAND2_X1 U8026 ( .A1(n9217), .A2(n7165), .ZN(n9533) );
  AOI21_X1 U8027 ( .B1(n6954), .B2(n6957), .A(n6953), .ZN(n6952) );
  INV_X1 U8028 ( .A(n13813), .ZN(n6953) );
  AOI21_X1 U8029 ( .B1(n6934), .B2(n6933), .A(n6649), .ZN(n6932) );
  INV_X1 U8030 ( .A(n13853), .ZN(n6933) );
  NAND2_X1 U8031 ( .A1(n13770), .A2(n13685), .ZN(n13840) );
  INV_X1 U8032 ( .A(n11781), .ZN(n6927) );
  AND2_X1 U8033 ( .A1(n14612), .A2(n14609), .ZN(n13625) );
  NOR2_X1 U8034 ( .A1(n7745), .A2(n6927), .ZN(n6926) );
  AOI21_X1 U8035 ( .B1(n7744), .B2(n11533), .A(n6605), .ZN(n7743) );
  OR2_X1 U8036 ( .A1(n11530), .A2(n11531), .ZN(n7018) );
  NAND2_X1 U8037 ( .A1(n12079), .A2(n6575), .ZN(n6838) );
  AOI21_X1 U8038 ( .B1(n12083), .B2(n6567), .A(n6837), .ZN(n6836) );
  AND4_X1 U8039 ( .A1(n8618), .A2(n8617), .A3(n8616), .A4(n8615), .ZN(n10929)
         );
  OR2_X1 U8040 ( .A1(n8915), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8597) );
  AND2_X1 U8041 ( .A1(n9152), .A2(n9151), .ZN(n9153) );
  XNOR2_X1 U8042 ( .A(n10156), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n10146) );
  INV_X1 U8043 ( .A(n10156), .ZN(n10084) );
  AND2_X1 U8044 ( .A1(n14699), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7169) );
  INV_X1 U8045 ( .A(n13902), .ZN(n13903) );
  INV_X1 U8046 ( .A(n7456), .ZN(n7455) );
  OAI21_X1 U8047 ( .B1(n7459), .B2(n7457), .A(n9115), .ZN(n7456) );
  NOR2_X1 U8048 ( .A1(n7580), .A2(n7578), .ZN(n7577) );
  INV_X1 U8049 ( .A(n14020), .ZN(n7578) );
  NAND2_X1 U8050 ( .A1(n14044), .A2(n7459), .ZN(n14028) );
  NOR2_X1 U8051 ( .A1(n14030), .A2(n7583), .ZN(n7582) );
  INV_X1 U8052 ( .A(n8967), .ZN(n7583) );
  OR2_X1 U8053 ( .A1(n14043), .A2(n8968), .ZN(n7584) );
  NAND2_X1 U8054 ( .A1(n14086), .A2(n9106), .ZN(n14072) );
  NAND2_X1 U8055 ( .A1(n14101), .A2(n12137), .ZN(n6884) );
  NAND2_X1 U8056 ( .A1(n6640), .A2(n6960), .ZN(n14102) );
  NOR2_X1 U8057 ( .A1(n14147), .A2(n14264), .ZN(n14135) );
  OR2_X1 U8058 ( .A1(n14622), .A2(n8830), .ZN(n12026) );
  NAND2_X1 U8059 ( .A1(n11810), .A2(n6532), .ZN(n14145) );
  INV_X1 U8060 ( .A(n12134), .ZN(n8831) );
  NAND2_X1 U8061 ( .A1(n8808), .A2(n8807), .ZN(n11850) );
  INV_X1 U8062 ( .A(n11852), .ZN(n8808) );
  AND2_X1 U8063 ( .A1(n12026), .A2(n12020), .ZN(n12134) );
  NAND2_X1 U8064 ( .A1(n6907), .A2(n6908), .ZN(n11810) );
  NAND2_X1 U8065 ( .A1(n11856), .A2(n12133), .ZN(n11855) );
  NAND2_X1 U8066 ( .A1(n11564), .A2(n9097), .ZN(n11443) );
  NAND2_X1 U8067 ( .A1(n11554), .A2(n8756), .ZN(n11449) );
  INV_X1 U8068 ( .A(n8682), .ZN(n7567) );
  AND2_X1 U8069 ( .A1(n6887), .A2(n12125), .ZN(n7566) );
  NAND2_X1 U8070 ( .A1(n11087), .A2(n8665), .ZN(n10942) );
  NAND2_X1 U8071 ( .A1(n10942), .A2(n12124), .ZN(n10941) );
  NAND2_X1 U8072 ( .A1(n7228), .A2(n7227), .ZN(n10943) );
  NAND2_X1 U8073 ( .A1(n11088), .A2(n11091), .ZN(n11087) );
  NAND2_X1 U8074 ( .A1(n7571), .A2(n14882), .ZN(n7570) );
  NOR2_X1 U8075 ( .A1(n10342), .A2(n10888), .ZN(n11950) );
  NAND2_X1 U8076 ( .A1(n8902), .A2(n8901), .ZN(n14251) );
  INV_X1 U8077 ( .A(n14269), .ZN(n14885) );
  OR2_X1 U8078 ( .A1(n8727), .A2(n9902), .ZN(n8607) );
  NAND3_X1 U8079 ( .A1(n9140), .A2(n9139), .A3(n9151), .ZN(n9953) );
  AND2_X1 U8080 ( .A1(n10185), .A2(n9958), .ZN(n10192) );
  NOR2_X1 U8081 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n7038) );
  INV_X1 U8082 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8542) );
  OAI21_X1 U8083 ( .B1(n9598), .B2(n7615), .A(n8957), .ZN(n8971) );
  INV_X1 U8084 ( .A(n9597), .ZN(n7615) );
  AND2_X1 U8085 ( .A1(n6618), .A2(n8898), .ZN(n7497) );
  NOR2_X1 U8086 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n7056) );
  INV_X1 U8087 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8819) );
  INV_X1 U8088 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n8815) );
  OR3_X1 U8089 ( .A1(n8743), .A2(P1_IR_REG_8__SCAN_IN), .A3(n8742), .ZN(n8818)
         );
  XNOR2_X1 U8090 ( .A(n8761), .B(n8760), .ZN(n9973) );
  INV_X1 U8091 ( .A(n7596), .ZN(n7595) );
  OAI21_X1 U8092 ( .B1(n8704), .B2(n7597), .A(n8725), .ZN(n7596) );
  INV_X1 U8093 ( .A(n8721), .ZN(n7597) );
  NAND2_X1 U8094 ( .A1(n8701), .A2(n8700), .ZN(n8705) );
  NAND2_X1 U8095 ( .A1(n7237), .A2(n7239), .ZN(n7235) );
  NAND2_X1 U8096 ( .A1(n8671), .A2(n8670), .ZN(n8684) );
  INV_X1 U8097 ( .A(n8648), .ZN(n7239) );
  INV_X1 U8098 ( .A(n7238), .ZN(n7237) );
  OAI21_X1 U8099 ( .B1(n8634), .B2(n7239), .A(n8652), .ZN(n7238) );
  NAND2_X1 U8100 ( .A1(n8635), .A2(n8634), .ZN(n8649) );
  OR2_X1 U8101 ( .A1(n7234), .A2(SI_3_), .ZN(n6983) );
  OAI21_X1 U8102 ( .B1(n6702), .B2(SI_2_), .A(n6892), .ZN(n8581) );
  NAND2_X1 U8103 ( .A1(n8579), .A2(n7605), .ZN(n6893) );
  NAND2_X1 U8104 ( .A1(n6893), .A2(n6891), .ZN(n8599) );
  INV_X1 U8105 ( .A(n8581), .ZN(n6891) );
  NAND2_X1 U8106 ( .A1(n8580), .A2(n9965), .ZN(n6989) );
  INV_X1 U8107 ( .A(n6758), .ZN(n14402) );
  NAND2_X1 U8108 ( .A1(n7067), .A2(n14410), .ZN(n14413) );
  AOI21_X1 U8109 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n15398), .A(n14369), .ZN(
        n14424) );
  NOR2_X1 U8110 ( .A1(n14397), .A2(n14396), .ZN(n14369) );
  AOI21_X1 U8111 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n14376), .A(n14375), .ZN(
        n14430) );
  NOR2_X1 U8112 ( .A1(n14393), .A2(n14392), .ZN(n14375) );
  OR2_X1 U8113 ( .A1(n14663), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7504) );
  INV_X1 U8114 ( .A(n12754), .ZN(n12726) );
  NAND2_X1 U8115 ( .A1(n6695), .A2(n7410), .ZN(n12230) );
  AOI21_X1 U8116 ( .B1(n6493), .B2(n7413), .A(n7411), .ZN(n7410) );
  INV_X1 U8117 ( .A(n12231), .ZN(n7411) );
  NAND3_X1 U8118 ( .A1(n10952), .A2(n10953), .A3(n10951), .ZN(n10961) );
  INV_X1 U8119 ( .A(n12360), .ZN(n12340) );
  INV_X1 U8120 ( .A(n11200), .ZN(n8471) );
  NAND2_X1 U8121 ( .A1(n8426), .A2(n10709), .ZN(n8427) );
  OR2_X1 U8122 ( .A1(n7540), .A2(n9186), .ZN(n7538) );
  INV_X1 U8123 ( .A(n8517), .ZN(n12597) );
  OR2_X1 U8124 ( .A1(n7846), .A2(n10723), .ZN(n7807) );
  NAND2_X1 U8125 ( .A1(n7804), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7808) );
  OR2_X1 U8126 ( .A1(n12451), .A2(n12452), .ZN(n7225) );
  INV_X1 U8127 ( .A(n7283), .ZN(n12461) );
  INV_X1 U8128 ( .A(n7281), .ZN(n12480) );
  INV_X1 U8129 ( .A(n7525), .ZN(n12482) );
  NOR2_X1 U8130 ( .A1(n12502), .A2(n12503), .ZN(n12505) );
  NAND2_X1 U8131 ( .A1(n7531), .A2(n7530), .ZN(n7529) );
  NAND2_X1 U8132 ( .A1(n12522), .A2(n12521), .ZN(n7530) );
  NAND2_X1 U8133 ( .A1(n6997), .A2(n15173), .ZN(n7220) );
  XNOR2_X1 U8134 ( .A(n12542), .B(n6998), .ZN(n6997) );
  INV_X1 U8135 ( .A(n12541), .ZN(n6998) );
  INV_X1 U8136 ( .A(n12546), .ZN(n7219) );
  INV_X1 U8137 ( .A(n12540), .ZN(n7272) );
  NAND2_X1 U8138 ( .A1(n7270), .A2(n6866), .ZN(n7273) );
  AOI21_X1 U8139 ( .B1(n12503), .B2(n7271), .A(n12528), .ZN(n7270) );
  XNOR2_X1 U8140 ( .A(n7223), .B(n7222), .ZN(n7221) );
  INV_X1 U8141 ( .A(n12537), .ZN(n7222) );
  NAND2_X1 U8142 ( .A1(n7531), .A2(n12530), .ZN(n7223) );
  AOI21_X1 U8143 ( .B1(n12890), .B2(n6474), .A(n8234), .ZN(n14512) );
  NAND2_X1 U8144 ( .A1(n8210), .A2(n8209), .ZN(n12217) );
  OR2_X1 U8145 ( .A1(n7833), .A2(n12159), .ZN(n8187) );
  INV_X1 U8146 ( .A(n12836), .ZN(n12590) );
  OR2_X1 U8147 ( .A1(n7833), .A2(n11305), .ZN(n8142) );
  NAND2_X1 U8148 ( .A1(n8133), .A2(n8132), .ZN(n12646) );
  NAND2_X1 U8149 ( .A1(n8119), .A2(n8118), .ZN(n12792) );
  OR2_X1 U8150 ( .A1(n7833), .A2(n11085), .ZN(n8118) );
  NOR2_X1 U8151 ( .A1(n6494), .A2(n12766), .ZN(n7685) );
  AND2_X1 U8152 ( .A1(n7766), .A2(n7688), .ZN(n7686) );
  NAND2_X1 U8153 ( .A1(n8532), .A2(n8531), .ZN(n8533) );
  NOR2_X1 U8154 ( .A1(n12768), .A2(n15222), .ZN(n6732) );
  OR2_X1 U8155 ( .A1(n10356), .A2(n10558), .ZN(n7841) );
  OR2_X1 U8156 ( .A1(n15244), .A2(n15195), .ZN(n12880) );
  INV_X1 U8157 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n7784) );
  OR2_X1 U8158 ( .A1(n7799), .A2(n7929), .ZN(n6821) );
  XNOR2_X1 U8159 ( .A(n8258), .B(n8257), .ZN(n11200) );
  INV_X1 U8160 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8257) );
  OAI21_X1 U8161 ( .B1(n8256), .B2(P3_IR_REG_21__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8258) );
  INV_X1 U8162 ( .A(n12459), .ZN(n12483) );
  NAND2_X1 U8163 ( .A1(n7636), .A2(n11655), .ZN(n7631) );
  INV_X1 U8164 ( .A(n7628), .ZN(n7626) );
  OR2_X1 U8165 ( .A1(n9961), .A2(n9286), .ZN(n9412) );
  NAND2_X1 U8166 ( .A1(n14911), .A2(n9842), .ZN(n9870) );
  OAI21_X1 U8167 ( .B1(n13045), .B2(n7657), .A(n7655), .ZN(n12972) );
  AOI21_X1 U8168 ( .B1(n7658), .B2(n7656), .A(n12966), .ZN(n7655) );
  INV_X1 U8169 ( .A(n7658), .ZN(n7657) );
  INV_X1 U8170 ( .A(n7659), .ZN(n7656) );
  OAI22_X1 U8171 ( .A1(n14543), .A2(n11841), .B1(n13063), .B2(n11840), .ZN(
        n11842) );
  NAND2_X1 U8172 ( .A1(n9499), .A2(n9498), .ZN(n13538) );
  OAI211_X1 U8173 ( .C1(n6717), .C2(n14911), .A(n10451), .B(n6715), .ZN(n10452) );
  INV_X1 U8174 ( .A(n10448), .ZN(n6717) );
  NAND2_X1 U8175 ( .A1(n14911), .A2(n7660), .ZN(n10483) );
  NAND2_X1 U8176 ( .A1(n9600), .A2(n9599), .ZN(n13501) );
  NAND2_X1 U8177 ( .A1(n6706), .A2(n7654), .ZN(n11513) );
  AOI21_X1 U8178 ( .B1(n11462), .B2(n11358), .A(n6657), .ZN(n7654) );
  NAND2_X1 U8179 ( .A1(n11461), .A2(n11358), .ZN(n6706) );
  OR2_X1 U8180 ( .A1(n9744), .A2(n9905), .ZN(n9292) );
  OR2_X1 U8181 ( .A1(n9290), .A2(n14929), .ZN(n7763) );
  NAND2_X1 U8182 ( .A1(n7624), .A2(n7623), .ZN(n14909) );
  AND2_X1 U8183 ( .A1(n10499), .A2(n14899), .ZN(n7623) );
  INV_X1 U8184 ( .A(n14903), .ZN(n14912) );
  AND2_X1 U8185 ( .A1(n9882), .A2(n9881), .ZN(n14914) );
  NAND2_X1 U8186 ( .A1(n10500), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14551) );
  NAND2_X1 U8187 ( .A1(n9479), .A2(n9478), .ZN(n13546) );
  NAND2_X1 U8188 ( .A1(n9611), .A2(n9610), .ZN(n13248) );
  OR2_X1 U8189 ( .A1(n13206), .A2(n13453), .ZN(n7178) );
  OR2_X1 U8190 ( .A1(n15076), .A2(n15066), .ZN(n15055) );
  OR2_X1 U8191 ( .A1(n9902), .A2(n9286), .ZN(n7025) );
  AND2_X1 U8192 ( .A1(n9313), .A2(n6552), .ZN(n7024) );
  NAND2_X1 U8193 ( .A1(n15082), .A2(n9878), .ZN(n15070) );
  NOR2_X1 U8194 ( .A1(n13456), .A2(n13455), .ZN(n13457) );
  AND2_X1 U8195 ( .A1(n13454), .A2(n15123), .ZN(n13455) );
  AOI21_X1 U8196 ( .B1(n11113), .B2(n11112), .A(n11111), .ZN(n11118) );
  AND2_X1 U8197 ( .A1(n13633), .A2(n13634), .ZN(n7734) );
  NAND2_X1 U8198 ( .A1(n8947), .A2(n7749), .ZN(n7748) );
  OR2_X1 U8199 ( .A1(n8947), .A2(n10156), .ZN(n8573) );
  NAND2_X1 U8200 ( .A1(n7751), .A2(n7750), .ZN(n7749) );
  NAND2_X1 U8201 ( .A1(n13821), .A2(n13680), .ZN(n13772) );
  NAND2_X1 U8202 ( .A1(n8930), .A2(n8929), .ZN(n14076) );
  OR2_X1 U8203 ( .A1(n13626), .A2(n13627), .ZN(n6990) );
  NAND2_X1 U8204 ( .A1(n8847), .A2(n8846), .ZN(n14604) );
  OAI21_X1 U8205 ( .B1(n8947), .B2(n7044), .A(n6834), .ZN(n10259) );
  INV_X1 U8206 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7044) );
  NAND2_X1 U8207 ( .A1(n8947), .A2(n14350), .ZN(n6834) );
  AND2_X1 U8208 ( .A1(n7739), .A2(n13662), .ZN(n7738) );
  NAND2_X1 U8209 ( .A1(n9009), .A2(n9008), .ZN(n13866) );
  NAND4_X1 U8210 ( .A1(n8645), .A2(n8644), .A3(n8643), .A4(n8642), .ZN(n13893)
         );
  OR2_X1 U8211 ( .A1(n8918), .A2(n8565), .ZN(n8566) );
  NOR2_X1 U8212 ( .A1(n10471), .A2(n10470), .ZN(n11032) );
  NAND2_X1 U8213 ( .A1(n10094), .A2(n10093), .ZN(n14767) );
  INV_X1 U8214 ( .A(n14138), .ZN(n13930) );
  OR2_X1 U8215 ( .A1(n13934), .A2(n10182), .ZN(n6824) );
  NAND2_X1 U8216 ( .A1(n13984), .A2(n6876), .ZN(n13973) );
  NAND2_X1 U8217 ( .A1(n8798), .A2(n8797), .ZN(n14597) );
  OR2_X1 U8218 ( .A1(n14896), .A2(n14173), .ZN(n7042) );
  NAND2_X1 U8219 ( .A1(n14288), .A2(n14230), .ZN(n7004) );
  NAND2_X1 U8220 ( .A1(n8731), .A2(n8730), .ZN(n11995) );
  NAND2_X1 U8221 ( .A1(n8713), .A2(n8712), .ZN(n11991) );
  OR2_X1 U8222 ( .A1(n9945), .A2(n8727), .ZN(n8713) );
  AND2_X1 U8223 ( .A1(n14896), .A2(n14881), .ZN(n14230) );
  AND2_X1 U8224 ( .A1(n6824), .A2(n13937), .ZN(n14280) );
  NAND2_X1 U8225 ( .A1(n6878), .A2(n9130), .ZN(n14178) );
  NAND2_X1 U8226 ( .A1(n9058), .A2(n9057), .ZN(n14180) );
  AND2_X1 U8227 ( .A1(n14288), .A2(n14306), .ZN(n6986) );
  OR2_X1 U8228 ( .A1(n9939), .A2(n8727), .ZN(n8692) );
  AND2_X1 U8229 ( .A1(n6959), .A2(n8545), .ZN(n6958) );
  NOR2_X1 U8230 ( .A1(n14458), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7511) );
  OR2_X1 U8231 ( .A1(n14654), .A2(n14653), .ZN(n6763) );
  OR2_X1 U8232 ( .A1(n14659), .A2(n7504), .ZN(n7500) );
  OR2_X1 U8233 ( .A1(n14659), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7503) );
  OR2_X1 U8234 ( .A1(n7510), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n7509) );
  OR2_X1 U8235 ( .A1(n14663), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n7508) );
  NOR2_X1 U8236 ( .A1(n14667), .A2(n14668), .ZN(n14666) );
  NAND2_X1 U8237 ( .A1(n13897), .A2(n7060), .ZN(n11949) );
  OAI21_X1 U8238 ( .B1(n7716), .B2(n7714), .A(n7712), .ZN(n9335) );
  AND2_X1 U8239 ( .A1(n9316), .A2(n9317), .ZN(n7714) );
  NAND2_X1 U8240 ( .A1(n7713), .A2(n7715), .ZN(n7712) );
  NAND2_X1 U8241 ( .A1(n11966), .A2(n11965), .ZN(n11970) );
  INV_X1 U8242 ( .A(n11969), .ZN(n7020) );
  NAND2_X1 U8243 ( .A1(n7136), .A2(n7722), .ZN(n9373) );
  NAND2_X1 U8244 ( .A1(n9355), .A2(n7723), .ZN(n7722) );
  INV_X1 U8245 ( .A(n9356), .ZN(n7723) );
  NAND2_X1 U8246 ( .A1(n7480), .A2(n11980), .ZN(n7479) );
  NAND2_X1 U8247 ( .A1(n6539), .A2(n6855), .ZN(n6854) );
  NAND2_X1 U8248 ( .A1(n7718), .A2(n6563), .ZN(n7717) );
  NOR2_X1 U8249 ( .A1(n6534), .A2(n7121), .ZN(n7120) );
  INV_X1 U8250 ( .A(n9436), .ZN(n7009) );
  NAND2_X1 U8251 ( .A1(n6535), .A2(n7152), .ZN(n7150) );
  NOR2_X1 U8252 ( .A1(n6535), .A2(n7152), .ZN(n7151) );
  AOI21_X1 U8253 ( .B1(n7477), .B2(n7475), .A(n7473), .ZN(n7472) );
  INV_X1 U8254 ( .A(n11999), .ZN(n7473) );
  OR2_X1 U8255 ( .A1(n12018), .A2(n7487), .ZN(n7486) );
  INV_X1 U8256 ( .A(n12031), .ZN(n7487) );
  MUX2_X1 U8257 ( .A(n12029), .B(n12028), .S(n12002), .Z(n12030) );
  AND2_X1 U8258 ( .A1(n12005), .A2(n6980), .ZN(n6840) );
  NOR2_X1 U8259 ( .A1(n12006), .A2(n6844), .ZN(n6843) );
  AND2_X1 U8260 ( .A1(n7485), .A2(n7488), .ZN(n7484) );
  AND2_X1 U8261 ( .A1(n12010), .A2(n12031), .ZN(n7485) );
  NAND2_X1 U8262 ( .A1(n12005), .A2(n12007), .ZN(n6841) );
  NOR2_X1 U8263 ( .A1(n7161), .A2(n7160), .ZN(n7159) );
  OAI21_X1 U8264 ( .B1(n7022), .B2(n12137), .A(n6850), .ZN(n12044) );
  NAND2_X1 U8265 ( .A1(n6849), .A2(n6848), .ZN(n12043) );
  AND2_X1 U8266 ( .A1(n12045), .A2(n6847), .ZN(n6848) );
  INV_X1 U8267 ( .A(n12050), .ZN(n6845) );
  INV_X1 U8268 ( .A(n9548), .ZN(n7155) );
  INV_X1 U8269 ( .A(n9549), .ZN(n7156) );
  NAND2_X1 U8270 ( .A1(n6862), .A2(n6865), .ZN(n12059) );
  NAND2_X1 U8271 ( .A1(n6987), .A2(n12055), .ZN(n6865) );
  INV_X1 U8272 ( .A(n9581), .ZN(n7147) );
  NAND2_X1 U8273 ( .A1(n12067), .A2(n12069), .ZN(n7495) );
  NAND2_X1 U8274 ( .A1(n6859), .A2(n6508), .ZN(n7494) );
  AND2_X1 U8275 ( .A1(n9006), .A2(SI_26_), .ZN(n7614) );
  INV_X1 U8276 ( .A(n8775), .ZN(n7602) );
  INV_X1 U8277 ( .A(n7601), .ZN(n7600) );
  OAI21_X1 U8278 ( .B1(n8772), .B2(n7602), .A(n8792), .ZN(n7601) );
  INV_X1 U8279 ( .A(n7997), .ZN(n7110) );
  INV_X1 U8280 ( .A(n7977), .ZN(n6742) );
  AND4_X1 U8281 ( .A1(n9802), .A2(n9767), .A3(n9766), .A4(n9765), .ZN(n9768)
         );
  AND2_X1 U8282 ( .A1(n9762), .A2(n9761), .ZN(n6971) );
  NAND2_X1 U8283 ( .A1(n9769), .A2(n7616), .ZN(n9772) );
  NOR2_X1 U8284 ( .A1(n9770), .A2(n9771), .ZN(n7616) );
  AND2_X1 U8285 ( .A1(n7380), .A2(n7378), .ZN(n7377) );
  INV_X1 U8286 ( .A(n13286), .ZN(n7378) );
  INV_X1 U8287 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n7117) );
  OAI21_X1 U8288 ( .B1(n14348), .B2(n14138), .A(n11945), .ZN(n11946) );
  INV_X1 U8289 ( .A(n12008), .ZN(n6910) );
  INV_X1 U8290 ( .A(n9671), .ZN(n7621) );
  AOI21_X1 U8291 ( .B1(n9004), .B2(n7614), .A(n7613), .ZN(n7612) );
  INV_X1 U8292 ( .A(n9022), .ZN(n7613) );
  AOI21_X1 U8293 ( .B1(n9004), .B2(n9006), .A(SI_26_), .ZN(n7611) );
  NAND2_X1 U8294 ( .A1(n7612), .A2(n7608), .ZN(n7607) );
  INV_X1 U8295 ( .A(n7614), .ZN(n7608) );
  INV_X1 U8296 ( .A(n8888), .ZN(n7250) );
  AOI21_X1 U8297 ( .B1(n7242), .B2(n7245), .A(n6608), .ZN(n7240) );
  AOI21_X1 U8298 ( .B1(n7246), .B2(n7244), .A(n7243), .ZN(n7242) );
  INV_X1 U8299 ( .A(n8759), .ZN(n7244) );
  INV_X1 U8300 ( .A(n7598), .ZN(n7243) );
  AOI21_X1 U8301 ( .B1(n7600), .B2(n7602), .A(n6597), .ZN(n7598) );
  INV_X1 U8302 ( .A(n7246), .ZN(n7245) );
  INV_X1 U8303 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n15325) );
  INV_X1 U8304 ( .A(P1_RD_REG_SCAN_IN), .ZN(n6794) );
  INV_X1 U8305 ( .A(P2_RD_REG_SCAN_IN), .ZN(n6797) );
  NOR2_X1 U8306 ( .A1(n14354), .A2(n14355), .ZN(n14356) );
  INV_X1 U8307 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n14357) );
  OR2_X1 U8308 ( .A1(n11682), .A2(n6696), .ZN(n11683) );
  OR2_X1 U8309 ( .A1(n11681), .A2(n12371), .ZN(n6697) );
  INV_X1 U8310 ( .A(n12177), .ZN(n7434) );
  OAI21_X1 U8311 ( .B1(n11687), .B2(n6683), .A(n6681), .ZN(n11905) );
  INV_X1 U8312 ( .A(n7414), .ZN(n6683) );
  AOI21_X1 U8313 ( .B1(n7414), .B2(n6682), .A(n6595), .ZN(n6681) );
  NOR2_X1 U8314 ( .A1(n10517), .A2(n6549), .ZN(n10404) );
  AND2_X1 U8315 ( .A1(n7215), .A2(n7214), .ZN(n10605) );
  INV_X1 U8316 ( .A(n11153), .ZN(n7287) );
  INV_X1 U8317 ( .A(n11395), .ZN(n7278) );
  NOR2_X1 U8318 ( .A1(n12428), .A2(n7049), .ZN(n12455) );
  AND2_X1 U8319 ( .A1(n12436), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7049) );
  AND2_X1 U8320 ( .A1(n7525), .A2(n7524), .ZN(n12516) );
  NAND2_X1 U8321 ( .A1(n12483), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7524) );
  NAND2_X1 U8322 ( .A1(n7672), .A2(n15441), .ZN(n7671) );
  NAND2_X1 U8323 ( .A1(n8506), .A2(n7668), .ZN(n7667) );
  INV_X1 U8324 ( .A(n7314), .ZN(n7310) );
  INV_X1 U8325 ( .A(n8350), .ZN(n7309) );
  INV_X1 U8326 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n7916) );
  NAND2_X1 U8327 ( .A1(n15178), .A2(n8485), .ZN(n8487) );
  NAND2_X1 U8328 ( .A1(n6969), .A2(n6968), .ZN(n8299) );
  INV_X1 U8329 ( .A(n8207), .ZN(n7032) );
  INV_X1 U8330 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7779) );
  OR2_X1 U8331 ( .A1(n8441), .A2(n6979), .ZN(n6978) );
  NAND2_X1 U8332 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), 
        .ZN(n6979) );
  INV_X1 U8333 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8438) );
  AOI21_X1 U8334 ( .B1(n8129), .B2(n6658), .A(n6749), .ZN(n8160) );
  NAND2_X1 U8335 ( .A1(n7544), .A2(n6750), .ZN(n6749) );
  INV_X1 U8336 ( .A(n8150), .ZN(n7545) );
  OAI21_X1 U8337 ( .B1(n7091), .B2(n6745), .A(n6743), .ZN(n8115) );
  AOI21_X1 U8338 ( .B1(n8107), .B2(n6744), .A(n6521), .ZN(n6743) );
  INV_X1 U8339 ( .A(n8107), .ZN(n6745) );
  INV_X1 U8340 ( .A(n7089), .ZN(n6744) );
  OAI21_X1 U8341 ( .B1(n7978), .B2(n7109), .A(n6740), .ZN(n8020) );
  AND2_X1 U8342 ( .A1(n7106), .A2(n6741), .ZN(n6740) );
  NAND2_X1 U8343 ( .A1(n7108), .A2(n6742), .ZN(n6741) );
  AOI21_X1 U8344 ( .B1(n7108), .B2(n7110), .A(n6516), .ZN(n7106) );
  INV_X1 U8345 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n7981) );
  INV_X1 U8346 ( .A(n6727), .ZN(n6726) );
  NOR2_X1 U8347 ( .A1(n6728), .A2(n7887), .ZN(n6727) );
  AND2_X1 U8348 ( .A1(n6881), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7887) );
  INV_X1 U8349 ( .A(n7873), .ZN(n6728) );
  INV_X1 U8350 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7773) );
  INV_X1 U8351 ( .A(n13035), .ZN(n6712) );
  NAND2_X1 U8352 ( .A1(n12913), .A2(n12914), .ZN(n6713) );
  OR4_X1 U8353 ( .A1(n13298), .A2(n13319), .A3(n13328), .A4(n9797), .ZN(n9798)
         );
  NOR2_X1 U8354 ( .A1(n13342), .A2(n13488), .ZN(n7187) );
  NOR2_X1 U8355 ( .A1(n9602), .A2(n9601), .ZN(n9621) );
  OR2_X1 U8356 ( .A1(n9385), .A2(n9384), .ZN(n9398) );
  INV_X1 U8357 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9397) );
  NOR2_X1 U8358 ( .A1(n9398), .A2(n9397), .ZN(n9414) );
  OR2_X1 U8359 ( .A1(n9362), .A2(n9361), .ZN(n9385) );
  INV_X1 U8360 ( .A(n10659), .ZN(n7406) );
  NAND2_X1 U8361 ( .A1(n10646), .A2(n9781), .ZN(n10636) );
  NAND2_X1 U8362 ( .A1(n9687), .A2(n9686), .ZN(n13454) );
  NAND2_X1 U8363 ( .A1(n9205), .A2(n7408), .ZN(n7407) );
  INV_X1 U8364 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n7408) );
  INV_X1 U8365 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9200) );
  OR2_X1 U8366 ( .A1(n9439), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n9456) );
  NAND2_X1 U8367 ( .A1(n6948), .A2(n6541), .ZN(n6947) );
  INV_X1 U8368 ( .A(n13757), .ZN(n6948) );
  INV_X1 U8370 ( .A(n7490), .ZN(n6837) );
  AOI21_X1 U8371 ( .B1(n6499), .B2(n7492), .A(n6589), .ZN(n7490) );
  NOR2_X1 U8372 ( .A1(n7493), .A2(n12084), .ZN(n7492) );
  OR2_X1 U8373 ( .A1(n14020), .A2(n7458), .ZN(n7457) );
  INV_X1 U8374 ( .A(n9113), .ZN(n7458) );
  NOR2_X1 U8375 ( .A1(n14221), .A2(n14305), .ZN(n7231) );
  NOR2_X1 U8376 ( .A1(n13837), .A2(n14597), .ZN(n6825) );
  OR2_X1 U8377 ( .A1(n8765), .A2(n8764), .ZN(n8785) );
  NAND2_X1 U8378 ( .A1(n7567), .A2(n12125), .ZN(n6886) );
  AND2_X1 U8379 ( .A1(n10931), .A2(n10912), .ZN(n10911) );
  AND2_X1 U8380 ( .A1(n6827), .A2(n6828), .ZN(n10857) );
  NOR2_X1 U8381 ( .A1(n13742), .A2(n10276), .ZN(n6827) );
  NAND2_X1 U8382 ( .A1(n10267), .A2(n10276), .ZN(n11959) );
  AND2_X1 U8383 ( .A1(n14348), .A2(n9124), .ZN(n11943) );
  NAND2_X1 U8384 ( .A1(n6830), .A2(n6829), .ZN(n14089) );
  NOR2_X1 U8385 ( .A1(n9004), .A2(n8986), .ZN(n7260) );
  INV_X1 U8386 ( .A(n9004), .ZN(n7261) );
  NAND2_X1 U8387 ( .A1(n7256), .A2(n8989), .ZN(n9005) );
  AND2_X1 U8388 ( .A1(n8909), .A2(n8894), .ZN(n8895) );
  AOI21_X1 U8389 ( .B1(n8873), .B2(n6528), .A(n7254), .ZN(n7253) );
  NOR2_X1 U8390 ( .A1(n8876), .A2(n10354), .ZN(n7254) );
  INV_X1 U8391 ( .A(n8873), .ZN(n7255) );
  OAI21_X1 U8392 ( .B1(n8761), .B2(n7245), .A(n7242), .ZN(n8834) );
  XNOR2_X1 U8393 ( .A(n8834), .B(n9948), .ZN(n8811) );
  NAND2_X1 U8394 ( .A1(n7061), .A2(n6810), .ZN(n6809) );
  NAND2_X1 U8395 ( .A1(n8580), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7061) );
  OAI21_X1 U8396 ( .B1(n9211), .B2(n9903), .A(n6984), .ZN(n7234) );
  NAND2_X1 U8397 ( .A1(n9211), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6984) );
  XNOR2_X1 U8398 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n6758) );
  INV_X1 U8399 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n14353) );
  XNOR2_X1 U8400 ( .A(n14356), .B(n14357), .ZN(n14398) );
  INV_X1 U8401 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15398) );
  NOR2_X1 U8402 ( .A1(n14368), .A2(n14367), .ZN(n14397) );
  NOR2_X1 U8403 ( .A1(n14418), .A2(n14366), .ZN(n14367) );
  AOI21_X1 U8404 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(n14374), .A(n14373), .ZN(
        n14393) );
  NOR2_X1 U8405 ( .A1(n14372), .A2(n14394), .ZN(n14373) );
  OAI22_X1 U8406 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14381), .B1(n14433), 
        .B2(n14380), .ZN(n14436) );
  NAND2_X1 U8407 ( .A1(n11906), .A2(n12367), .ZN(n6694) );
  OR2_X1 U8408 ( .A1(n11908), .A2(n7413), .ZN(n7412) );
  NAND2_X1 U8409 ( .A1(n12162), .A2(n6672), .ZN(n7413) );
  AND2_X1 U8410 ( .A1(n7084), .A2(n7445), .ZN(n7083) );
  AND2_X1 U8411 ( .A1(n11740), .A2(n11738), .ZN(n7414) );
  AOI21_X1 U8412 ( .B1(n12224), .B2(n12198), .A(n12201), .ZN(n7441) );
  INV_X1 U8413 ( .A(n7441), .ZN(n7438) );
  XNOR2_X1 U8414 ( .A(n11677), .B(n7085), .ZN(n11673) );
  NAND2_X1 U8415 ( .A1(n7071), .A2(n7073), .ZN(n6689) );
  AOI21_X1 U8416 ( .B1(n7075), .B2(n7078), .A(n7074), .ZN(n7073) );
  INV_X1 U8417 ( .A(n12300), .ZN(n7074) );
  AND2_X1 U8418 ( .A1(n6694), .A2(n6555), .ZN(n11907) );
  NOR2_X1 U8419 ( .A1(n8056), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8067) );
  XNOR2_X1 U8420 ( .A(n10712), .B(n6691), .ZN(n11495) );
  NAND2_X1 U8421 ( .A1(n7081), .A2(n12186), .ZN(n12288) );
  NAND2_X1 U8422 ( .A1(n12317), .A2(n7445), .ZN(n7081) );
  AND2_X1 U8423 ( .A1(n12267), .A2(n12190), .ZN(n12289) );
  OR2_X1 U8424 ( .A1(n8144), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8154) );
  NAND2_X1 U8425 ( .A1(n11687), .A2(n11688), .ZN(n11739) );
  AND2_X1 U8426 ( .A1(n7430), .A2(n7076), .ZN(n7075) );
  NAND2_X1 U8427 ( .A1(n7432), .A2(n7077), .ZN(n7076) );
  AOI21_X1 U8428 ( .B1(n7432), .B2(n7434), .A(n6566), .ZN(n7430) );
  INV_X1 U8429 ( .A(n12173), .ZN(n7077) );
  INV_X1 U8430 ( .A(n7432), .ZN(n7078) );
  NAND2_X1 U8431 ( .A1(n11907), .A2(n11908), .ZN(n12163) );
  NAND2_X1 U8432 ( .A1(n8134), .A2(n12319), .ZN(n8144) );
  AND2_X1 U8433 ( .A1(n8120), .A2(n12256), .ZN(n8134) );
  NAND2_X1 U8434 ( .A1(n12185), .A2(n12184), .ZN(n7445) );
  NAND2_X1 U8435 ( .A1(n7069), .A2(n7444), .ZN(n7443) );
  INV_X1 U8436 ( .A(n12184), .ZN(n7444) );
  XNOR2_X1 U8437 ( .A(n11905), .B(n11903), .ZN(n11906) );
  OAI211_X1 U8438 ( .C1(n7833), .C2(SI_2_), .A(n7826), .B(n7825), .ZN(n10724)
         );
  OR2_X1 U8439 ( .A1(n10356), .A2(n10406), .ZN(n7825) );
  AND2_X1 U8440 ( .A1(n10706), .A2(n10705), .ZN(n12330) );
  NAND2_X1 U8441 ( .A1(n7335), .A2(n7006), .ZN(n9173) );
  NOR2_X1 U8442 ( .A1(n7337), .A2(n7336), .ZN(n7335) );
  OR2_X1 U8443 ( .A1(n6511), .A2(n7099), .ZN(n7006) );
  NAND2_X1 U8444 ( .A1(n7542), .A2(n7541), .ZN(n7540) );
  NAND2_X1 U8445 ( .A1(n8401), .A2(n8400), .ZN(n7542) );
  OR2_X1 U8446 ( .A1(n8236), .A2(n10378), .ZN(n7805) );
  INV_X1 U8447 ( .A(n7194), .ZN(n7193) );
  NAND2_X1 U8448 ( .A1(n10368), .A2(n7519), .ZN(n10534) );
  NAND2_X1 U8449 ( .A1(n6871), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n10533) );
  NAND2_X1 U8450 ( .A1(n7191), .A2(n7190), .ZN(n10370) );
  OAI21_X1 U8451 ( .B1(n7837), .B2(n7266), .A(n10399), .ZN(n7190) );
  INV_X1 U8452 ( .A(n7266), .ZN(n7192) );
  NAND2_X1 U8453 ( .A1(n10403), .A2(n10514), .ZN(n10549) );
  OR2_X1 U8454 ( .A1(n10549), .A2(n7828), .ZN(n10547) );
  AOI21_X1 U8455 ( .B1(n10547), .B2(n10514), .A(n10515), .ZN(n10517) );
  NAND2_X1 U8456 ( .A1(n7216), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7215) );
  INV_X1 U8457 ( .A(n7046), .ZN(n10598) );
  INV_X1 U8458 ( .A(n11148), .ZN(n7213) );
  INV_X1 U8459 ( .A(n11389), .ZN(n7199) );
  NOR2_X1 U8460 ( .A1(n11753), .A2(n11754), .ZN(n11755) );
  AOI21_X1 U8461 ( .B1(n7290), .B2(n7291), .A(n12388), .ZN(n6873) );
  OR2_X1 U8462 ( .A1(n12401), .A2(n12402), .ZN(n7518) );
  INV_X1 U8463 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7698) );
  XNOR2_X1 U8464 ( .A(n12455), .B(n12456), .ZN(n12430) );
  AND2_X1 U8465 ( .A1(n7517), .A2(n7516), .ZN(n12450) );
  NAND2_X1 U8466 ( .A1(n12436), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7516) );
  NAND2_X1 U8467 ( .A1(n12483), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7280) );
  XNOR2_X1 U8468 ( .A(n12516), .B(n12517), .ZN(n12484) );
  INV_X1 U8469 ( .A(n12504), .ZN(n7271) );
  NAND2_X1 U8470 ( .A1(n12502), .A2(n7271), .ZN(n6866) );
  AND4_X1 U8471 ( .A1(n8206), .A2(n8205), .A3(n8204), .A4(n8203), .ZN(n12226)
         );
  NOR2_X1 U8472 ( .A1(n8200), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n12549) );
  AND4_X1 U8473 ( .A1(n8194), .A2(n8193), .A3(n8192), .A4(n8191), .ZN(n8523)
         );
  NAND2_X1 U8474 ( .A1(n6801), .A2(n14499), .ZN(n6800) );
  NAND2_X1 U8475 ( .A1(n8527), .A2(n6569), .ZN(n6801) );
  NAND2_X1 U8476 ( .A1(n8262), .A2(n7339), .ZN(n7338) );
  NAND2_X1 U8477 ( .A1(n8261), .A2(n8264), .ZN(n7339) );
  NOR2_X1 U8478 ( .A1(n8260), .A2(n7341), .ZN(n7340) );
  INV_X1 U8479 ( .A(n8263), .ZN(n7341) );
  NAND3_X1 U8480 ( .A1(n8261), .A2(n12578), .A3(n6753), .ZN(n6752) );
  AND2_X1 U8481 ( .A1(n8262), .A2(n8261), .ZN(n12579) );
  NAND2_X1 U8482 ( .A1(n7316), .A2(n7318), .ZN(n12608) );
  AOI21_X1 U8483 ( .B1(n7317), .B2(n7324), .A(n7319), .ZN(n7318) );
  INV_X1 U8484 ( .A(n8265), .ZN(n7319) );
  OR2_X1 U8485 ( .A1(n12608), .A2(n12609), .ZN(n7100) );
  NAND2_X1 U8486 ( .A1(n8512), .A2(n12667), .ZN(n8513) );
  INV_X1 U8487 ( .A(n7694), .ZN(n7691) );
  AOI21_X1 U8488 ( .B1(n12677), .B2(n8510), .A(n8509), .ZN(n12665) );
  OR2_X1 U8489 ( .A1(n8097), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8109) );
  INV_X1 U8490 ( .A(n12365), .ZN(n12679) );
  NOR2_X1 U8491 ( .A1(n6805), .A2(n6804), .ZN(n12677) );
  INV_X1 U8492 ( .A(n8508), .ZN(n6804) );
  INV_X1 U8493 ( .A(n12688), .ZN(n6805) );
  INV_X1 U8494 ( .A(n7664), .ZN(n7662) );
  AOI21_X1 U8495 ( .B1(n7665), .B2(n7669), .A(n7757), .ZN(n7664) );
  AND2_X1 U8496 ( .A1(n8280), .A2(n8279), .ZN(n12695) );
  NOR2_X1 U8497 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(n8068), .ZN(n8086) );
  NOR2_X1 U8498 ( .A1(n6647), .A2(n7690), .ZN(n7689) );
  AND2_X1 U8499 ( .A1(n8012), .A2(n15429), .ZN(n8031) );
  OR2_X1 U8500 ( .A1(n7968), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7988) );
  NAND2_X1 U8501 ( .A1(n11798), .A2(n8496), .ZN(n14495) );
  NOR2_X1 U8502 ( .A1(n7303), .A2(n6590), .ZN(n7302) );
  NOR2_X1 U8503 ( .A1(n7304), .A2(n7951), .ZN(n7303) );
  NAND2_X1 U8504 ( .A1(n11703), .A2(n7951), .ZN(n7307) );
  NAND2_X1 U8505 ( .A1(n7307), .A2(n7305), .ZN(n14501) );
  NAND2_X1 U8506 ( .A1(n11286), .A2(n8493), .ZN(n11484) );
  NOR2_X1 U8507 ( .A1(n7899), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7917) );
  OR2_X1 U8508 ( .A1(n7880), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7899) );
  NAND2_X1 U8509 ( .A1(n7293), .A2(n8305), .ZN(n11240) );
  NAND2_X1 U8510 ( .A1(n10836), .A2(n8301), .ZN(n11309) );
  AND2_X1 U8511 ( .A1(n8305), .A2(n8306), .ZN(n11314) );
  INV_X1 U8512 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10416) );
  INV_X1 U8513 ( .A(n8485), .ZN(n15180) );
  AND2_X1 U8514 ( .A1(n10688), .A2(n15188), .ZN(n11192) );
  NOR2_X1 U8515 ( .A1(n8527), .A2(n6569), .ZN(n7700) );
  XNOR2_X1 U8516 ( .A(n9173), .B(n9167), .ZN(n12214) );
  AND2_X1 U8517 ( .A1(n8307), .A2(n9182), .ZN(n10615) );
  INV_X1 U8518 ( .A(n7559), .ZN(n7558) );
  OAI21_X1 U8519 ( .B1(n8220), .B2(n6524), .A(n7560), .ZN(n7559) );
  INV_X1 U8520 ( .A(n8231), .ZN(n7560) );
  NAND2_X1 U8521 ( .A1(n7557), .A2(n7554), .ZN(n7553) );
  OR2_X1 U8522 ( .A1(n7558), .A2(n8233), .ZN(n7554) );
  AOI21_X1 U8523 ( .B1(n7558), .B2(n6524), .A(n6680), .ZN(n7557) );
  INV_X1 U8524 ( .A(n8233), .ZN(n7556) );
  OAI22_X1 U8525 ( .A1(n8183), .A2(n8184), .B1(P2_DATAO_REG_26__SCAN_IN), .B2(
        n13587), .ZN(n8195) );
  INV_X1 U8526 ( .A(n7347), .ZN(n8429) );
  XNOR2_X1 U8527 ( .A(n8253), .B(P3_IR_REG_20__SCAN_IN), .ZN(n9185) );
  XNOR2_X1 U8528 ( .A(n8095), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12531) );
  INV_X1 U8529 ( .A(n7087), .ZN(n8080) );
  NAND2_X1 U8530 ( .A1(n7087), .A2(n8078), .ZN(n8247) );
  OAI21_X1 U8531 ( .B1(n7096), .B2(n6748), .A(n6746), .ZN(n8074) );
  AOI21_X1 U8532 ( .B1(n6747), .B2(n8062), .A(n6522), .ZN(n6746) );
  INV_X1 U8533 ( .A(n8062), .ZN(n6748) );
  OR2_X1 U8534 ( .A1(n8006), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n8023) );
  XNOR2_X1 U8535 ( .A(n8020), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8019) );
  INV_X1 U8536 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n7963) );
  NAND2_X1 U8537 ( .A1(n6739), .A2(n7101), .ZN(n7975) );
  AOI21_X1 U8538 ( .B1(n7103), .B2(n7105), .A(n6651), .ZN(n7101) );
  OAI21_X1 U8539 ( .B1(n7925), .B2(n6738), .A(n6599), .ZN(n6739) );
  XNOR2_X1 U8540 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n7974) );
  XNOR2_X1 U8541 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n7924) );
  XNOR2_X1 U8542 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n7906) );
  AND2_X1 U8543 ( .A1(n7772), .A2(n7771), .ZN(n7442) );
  XNOR2_X1 U8544 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7820) );
  NAND2_X1 U8545 ( .A1(n6498), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7523) );
  AND2_X1 U8546 ( .A1(n9965), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7821) );
  AND2_X1 U8547 ( .A1(n12940), .A2(n12936), .ZN(n7658) );
  INV_X1 U8548 ( .A(n6766), .ZN(n10502) );
  INV_X1 U8549 ( .A(n12958), .ZN(n7650) );
  AND2_X1 U8550 ( .A1(n12916), .A2(n12915), .ZN(n7651) );
  NAND2_X1 U8551 ( .A1(n6716), .A2(n10448), .ZN(n6715) );
  INV_X1 U8552 ( .A(n7660), .ZN(n6716) );
  AND2_X1 U8553 ( .A1(n9500), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9514) );
  AND2_X1 U8554 ( .A1(n9867), .A2(n9842), .ZN(n7660) );
  INV_X1 U8555 ( .A(n9869), .ZN(n9867) );
  INV_X1 U8556 ( .A(n7648), .ZN(n13017) );
  XNOR2_X1 U8557 ( .A(n10502), .B(n12968), .ZN(n9835) );
  OR2_X1 U8558 ( .A1(n9538), .A2(n9537), .ZN(n9556) );
  NAND2_X1 U8559 ( .A1(n9514), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9538) );
  NOR2_X1 U8560 ( .A1(n12911), .A2(n7641), .ZN(n7640) );
  NAND2_X1 U8561 ( .A1(n7639), .A2(n12910), .ZN(n7638) );
  INV_X1 U8562 ( .A(n7642), .ZN(n7639) );
  INV_X1 U8563 ( .A(n10830), .ZN(n10828) );
  AND2_X1 U8564 ( .A1(n13046), .A2(n12932), .ZN(n7659) );
  NAND2_X1 U8565 ( .A1(n7127), .A2(n7130), .ZN(n9804) );
  NAND2_X1 U8566 ( .A1(n9735), .A2(n7134), .ZN(n6972) );
  NAND2_X1 U8567 ( .A1(n9736), .A2(n7125), .ZN(n7122) );
  NOR2_X1 U8568 ( .A1(n7129), .A2(n7126), .ZN(n7125) );
  AND3_X1 U8569 ( .A1(n9808), .A2(n9550), .A3(n11439), .ZN(n7702) );
  INV_X1 U8570 ( .A(n9713), .ZN(n9605) );
  OR2_X1 U8571 ( .A1(n14978), .A2(n14977), .ZN(n14980) );
  NOR2_X1 U8572 ( .A1(n13274), .A2(n7248), .ZN(n13228) );
  NOR2_X1 U8573 ( .A1(n13282), .A2(n13230), .ZN(n7248) );
  OR2_X1 U8574 ( .A1(n13230), .A2(n14541), .ZN(n7063) );
  NAND2_X1 U8575 ( .A1(n13465), .A2(n6578), .ZN(n13273) );
  AND2_X1 U8576 ( .A1(n9712), .A2(n9646), .ZN(n13303) );
  OR2_X1 U8577 ( .A1(n13482), .A2(n13252), .ZN(n13253) );
  NAND2_X1 U8578 ( .A1(n7187), .A2(n13317), .ZN(n13312) );
  INV_X1 U8579 ( .A(n7187), .ZN(n13330) );
  INV_X1 U8580 ( .A(n6819), .ZN(n13385) );
  OAI21_X1 U8581 ( .B1(n6791), .B2(n7390), .A(n7386), .ZN(n13414) );
  AOI21_X1 U8582 ( .B1(n7389), .B2(n7391), .A(n7387), .ZN(n7386) );
  INV_X1 U8583 ( .A(n13213), .ZN(n7387) );
  INV_X1 U8584 ( .A(n13238), .ZN(n13413) );
  NAND2_X1 U8585 ( .A1(n6820), .A2(n7181), .ZN(n11924) );
  INV_X1 U8586 ( .A(n13546), .ZN(n7181) );
  NOR2_X1 U8587 ( .A1(n9481), .A2(n9480), .ZN(n9500) );
  NAND2_X1 U8588 ( .A1(n6782), .A2(n6781), .ZN(n14552) );
  AOI21_X1 U8589 ( .B1(n6783), .B2(n11718), .A(n6551), .ZN(n6781) );
  NAND2_X1 U8590 ( .A1(n11615), .A2(n6783), .ZN(n6782) );
  NAND2_X1 U8591 ( .A1(n11719), .A2(n11718), .ZN(n6699) );
  OR2_X1 U8592 ( .A1(n9428), .A2(n11361), .ZN(n9445) );
  NOR2_X1 U8593 ( .A1(n9445), .A2(n9444), .ZN(n9462) );
  NAND2_X1 U8594 ( .A1(n6769), .A2(n6767), .ZN(n11224) );
  AOI21_X1 U8595 ( .B1(n6771), .B2(n6768), .A(n6588), .ZN(n6767) );
  OR2_X1 U8596 ( .A1(n10995), .A2(n6770), .ZN(n6769) );
  INV_X1 U8597 ( .A(n10997), .ZN(n7179) );
  INV_X1 U8598 ( .A(n14541), .ZN(n13049) );
  NAND2_X1 U8599 ( .A1(n10434), .A2(n10435), .ZN(n10647) );
  XNOR2_X1 U8600 ( .A(n9786), .B(n9784), .ZN(n7398) );
  INV_X1 U8601 ( .A(n9833), .ZN(n7033) );
  OAI21_X1 U8602 ( .B1(n9916), .B2(n9286), .A(n9259), .ZN(n15105) );
  INV_X1 U8603 ( .A(n9996), .ZN(n9831) );
  AND2_X1 U8604 ( .A1(n9217), .A2(n6625), .ZN(n9228) );
  AND2_X1 U8605 ( .A1(n9223), .A2(n7166), .ZN(n7165) );
  INV_X1 U8606 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7166) );
  OR2_X1 U8607 ( .A1(n9456), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n9475) );
  AND2_X1 U8608 ( .A1(n9382), .A2(n9407), .ZN(n10018) );
  INV_X1 U8609 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n9357) );
  AOI21_X1 U8610 ( .B1(n7727), .B2(n7729), .A(n6582), .ZN(n7724) );
  NOR2_X1 U8611 ( .A1(n8785), .A2(n8784), .ZN(n8799) );
  NAND2_X1 U8612 ( .A1(n13852), .A2(n13853), .ZN(n6936) );
  NAND2_X1 U8613 ( .A1(n13763), .A2(n6947), .ZN(n6946) );
  AND2_X1 U8614 ( .A1(n13859), .A2(n7728), .ZN(n7727) );
  OR2_X1 U8615 ( .A1(n13794), .A2(n7729), .ZN(n7728) );
  AND2_X1 U8616 ( .A1(n7724), .A2(n6541), .ZN(n6949) );
  AND2_X1 U8617 ( .A1(n6945), .A2(n6943), .ZN(n6942) );
  NAND2_X1 U8618 ( .A1(n6944), .A2(n6950), .ZN(n6943) );
  OR2_X1 U8619 ( .A1(n6949), .A2(n6946), .ZN(n6945) );
  INV_X1 U8620 ( .A(n6947), .ZN(n6944) );
  OR2_X1 U8621 ( .A1(n8676), .A2(n11119), .ZN(n8694) );
  NAND2_X1 U8622 ( .A1(n9676), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7750) );
  INV_X1 U8623 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10899) );
  OR2_X1 U8624 ( .A1(n8849), .A2(n8848), .ZN(n8866) );
  AND2_X1 U8625 ( .A1(n7730), .A2(n6955), .ZN(n6954) );
  AOI21_X1 U8626 ( .B1(n7731), .B2(n7733), .A(n6581), .ZN(n7730) );
  NAND2_X1 U8627 ( .A1(n7731), .A2(n6956), .ZN(n6955) );
  INV_X1 U8628 ( .A(n7731), .ZN(n6957) );
  NOR2_X1 U8629 ( .A1(n11532), .A2(n11533), .ZN(n11541) );
  NAND2_X1 U8630 ( .A1(n13840), .A2(n13841), .ZN(n13839) );
  INV_X1 U8631 ( .A(n8961), .ZN(n8960) );
  XNOR2_X1 U8632 ( .A(n7023), .B(n11048), .ZN(n10269) );
  NOR2_X1 U8633 ( .A1(n8866), .A2(n8865), .ZN(n8882) );
  NOR2_X1 U8634 ( .A1(n7741), .A2(n7737), .ZN(n7736) );
  INV_X1 U8635 ( .A(n14602), .ZN(n7737) );
  INV_X1 U8636 ( .A(n13803), .ZN(n7741) );
  NAND2_X1 U8637 ( .A1(n13803), .A2(n7740), .ZN(n7739) );
  INV_X1 U8638 ( .A(n13655), .ZN(n7740) );
  AND2_X1 U8639 ( .A1(n8799), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8823) );
  NAND2_X1 U8640 ( .A1(n8823), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8849) );
  NAND2_X1 U8641 ( .A1(n14594), .A2(n13641), .ZN(n13645) );
  NAND2_X1 U8642 ( .A1(n8594), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8575) );
  NOR2_X1 U8643 ( .A1(n10163), .A2(n6637), .ZN(n10167) );
  NOR2_X1 U8644 ( .A1(n10167), .A2(n10166), .ZN(n10286) );
  NOR2_X1 U8645 ( .A1(n11032), .A2(n6638), .ZN(n14684) );
  NOR2_X1 U8646 ( .A1(n14684), .A2(n14683), .ZN(n14682) );
  NAND2_X1 U8647 ( .A1(n11025), .A2(n11026), .ZN(n13912) );
  NOR2_X1 U8648 ( .A1(n14703), .A2(n14704), .ZN(n14705) );
  OR2_X1 U8649 ( .A1(n13910), .A2(n13909), .ZN(n14768) );
  AND2_X1 U8650 ( .A1(n13908), .A2(n14777), .ZN(n13910) );
  NAND2_X1 U8651 ( .A1(n9122), .A2(n9121), .ZN(n13941) );
  INV_X1 U8652 ( .A(n13981), .ZN(n9036) );
  NOR2_X1 U8653 ( .A1(n12141), .A2(n6899), .ZN(n6898) );
  INV_X1 U8654 ( .A(n6904), .ZN(n6899) );
  NAND2_X1 U8655 ( .A1(n12141), .A2(n6904), .ZN(n6901) );
  AND2_X1 U8656 ( .A1(n6904), .A2(n6906), .ZN(n6902) );
  INV_X1 U8657 ( .A(n9122), .ZN(n13963) );
  INV_X1 U8658 ( .A(n7226), .ZN(n13989) );
  AND2_X1 U8659 ( .A1(n13971), .A2(n9037), .ZN(n6876) );
  NOR2_X1 U8660 ( .A1(n14035), .A2(n14201), .ZN(n14012) );
  NAND2_X1 U8661 ( .A1(n7229), .A2(n14060), .ZN(n14035) );
  AND2_X1 U8662 ( .A1(n7231), .A2(n7230), .ZN(n7229) );
  NAND2_X1 U8663 ( .A1(n14044), .A2(n9111), .ZN(n14026) );
  AOI21_X1 U8664 ( .B1(n6916), .B2(n14066), .A(n6538), .ZN(n6915) );
  NAND2_X1 U8665 ( .A1(n14086), .A2(n6912), .ZN(n6917) );
  NAND2_X1 U8666 ( .A1(n14060), .A2(n7231), .ZN(n14047) );
  NAND2_X1 U8667 ( .A1(n14060), .A2(n14065), .ZN(n14061) );
  NOR2_X1 U8668 ( .A1(n14073), .A2(n7586), .ZN(n7585) );
  INV_X1 U8669 ( .A(n8923), .ZN(n7586) );
  AOI21_X1 U8670 ( .B1(n6490), .B2(n12133), .A(n6587), .ZN(n7587) );
  NAND2_X1 U8671 ( .A1(n11472), .A2(n14642), .ZN(n11853) );
  NAND2_X1 U8672 ( .A1(n7461), .A2(n9095), .ZN(n7460) );
  NAND2_X1 U8673 ( .A1(n6919), .A2(n9095), .ZN(n6918) );
  NAND2_X1 U8674 ( .A1(n11419), .A2(n8720), .ZN(n11372) );
  XNOR2_X1 U8675 ( .A(n11991), .B(n11545), .ZN(n12126) );
  OR2_X1 U8676 ( .A1(n8694), .A2(n8693), .ZN(n8715) );
  NOR2_X1 U8677 ( .A1(n8715), .A2(n8714), .ZN(n8750) );
  NAND2_X1 U8678 ( .A1(n10871), .A2(n7462), .ZN(n11423) );
  INV_X1 U8679 ( .A(n6919), .ZN(n7462) );
  OR2_X1 U8680 ( .A1(n10870), .A2(n12125), .ZN(n10871) );
  AOI21_X1 U8681 ( .B1(n12121), .B2(n7449), .A(n6568), .ZN(n7448) );
  INV_X1 U8682 ( .A(n9088), .ZN(n7449) );
  NAND2_X1 U8683 ( .A1(n6828), .A2(n14861), .ZN(n14836) );
  AND2_X1 U8684 ( .A1(n11421), .A2(n14797), .ZN(n6832) );
  NAND2_X1 U8685 ( .A1(n11427), .A2(n14868), .ZN(n14887) );
  OAI21_X1 U8686 ( .B1(n9742), .B2(n9740), .A(n9675), .ZN(n9679) );
  XNOR2_X1 U8687 ( .A(n9742), .B(n9741), .ZN(n13573) );
  XNOR2_X1 U8688 ( .A(n9053), .B(n9052), .ZN(n13578) );
  XNOR2_X1 U8689 ( .A(n9138), .B(P1_IR_REG_26__SCAN_IN), .ZN(n9151) );
  INV_X1 U8690 ( .A(n8543), .ZN(n9136) );
  XNOR2_X1 U8691 ( .A(n9005), .B(n9004), .ZN(n13590) );
  XNOR2_X1 U8692 ( .A(n9131), .B(P1_IR_REG_24__SCAN_IN), .ZN(n9154) );
  XNOR2_X1 U8693 ( .A(n8975), .B(n8986), .ZN(n13594) );
  XNOR2_X1 U8694 ( .A(n9157), .B(n9156), .ZN(n10175) );
  INV_X1 U8695 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9156) );
  XNOR2_X1 U8696 ( .A(n8928), .B(n8927), .ZN(n11437) );
  INV_X1 U8697 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8844) );
  XNOR2_X1 U8698 ( .A(n8811), .B(n8835), .ZN(n10423) );
  NAND2_X1 U8699 ( .A1(n7599), .A2(n8775), .ZN(n8793) );
  NAND2_X1 U8700 ( .A1(n8773), .A2(n8772), .ZN(n7599) );
  INV_X1 U8701 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8741) );
  INV_X1 U8702 ( .A(n7564), .ZN(n8842) );
  NAND2_X1 U8703 ( .A1(n8539), .A2(n8584), .ZN(n8587) );
  INV_X1 U8704 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8539) );
  INV_X1 U8705 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14351) );
  XNOR2_X1 U8706 ( .A(n6757), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n14401) );
  XNOR2_X1 U8707 ( .A(n14398), .B(n7053), .ZN(n14400) );
  INV_X1 U8708 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7053) );
  INV_X1 U8709 ( .A(n6760), .ZN(n14414) );
  NOR2_X1 U8710 ( .A1(n14361), .A2(n14360), .ZN(n14415) );
  NAND2_X1 U8711 ( .A1(n6764), .A2(n14420), .ZN(n14421) );
  NAND2_X1 U8712 ( .A1(n15450), .A2(n15451), .ZN(n6764) );
  AOI21_X1 U8713 ( .B1(n14371), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n14370), .ZN(
        n14395) );
  AND2_X1 U8714 ( .A1(n14425), .A2(n14424), .ZN(n14370) );
  NAND2_X1 U8715 ( .A1(n7512), .A2(n6763), .ZN(n14435) );
  OR2_X1 U8716 ( .A1(n14659), .A2(n7502), .ZN(n7501) );
  AND2_X1 U8717 ( .A1(n7504), .A2(n7506), .ZN(n7502) );
  NAND2_X1 U8718 ( .A1(n15002), .A2(n7507), .ZN(n7506) );
  INV_X1 U8719 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7507) );
  OR2_X1 U8720 ( .A1(n14390), .A2(n14389), .ZN(n14471) );
  XNOR2_X1 U8721 ( .A(n6688), .B(n12224), .ZN(n6687) );
  NAND2_X1 U8722 ( .A1(n12337), .A2(n12199), .ZN(n6688) );
  NAND2_X1 U8723 ( .A1(n11739), .A2(n7414), .ZN(n11867) );
  NAND2_X1 U8724 ( .A1(n7431), .A2(n12177), .ZN(n12245) );
  NAND2_X1 U8725 ( .A1(n12326), .A2(n12325), .ZN(n7431) );
  NAND2_X1 U8726 ( .A1(n12338), .A2(n12339), .ZN(n12337) );
  NAND2_X1 U8727 ( .A1(n6689), .A2(n12181), .ZN(n12254) );
  NAND2_X1 U8728 ( .A1(n7417), .A2(n12169), .ZN(n12274) );
  NAND2_X1 U8729 ( .A1(n12350), .A2(n12167), .ZN(n7417) );
  NAND2_X1 U8730 ( .A1(n11208), .A2(n7426), .ZN(n7422) );
  XNOR2_X1 U8731 ( .A(n11495), .B(n6690), .ZN(n11211) );
  NAND2_X1 U8732 ( .A1(n7415), .A2(n7416), .ZN(n12281) );
  AOI21_X1 U8733 ( .B1(n7418), .B2(n7421), .A(n6592), .ZN(n7416) );
  INV_X1 U8734 ( .A(n12169), .ZN(n7421) );
  NAND2_X1 U8735 ( .A1(n10961), .A2(n7428), .ZN(n10966) );
  NAND2_X1 U8736 ( .A1(n7072), .A2(n7075), .ZN(n12301) );
  OR2_X1 U8737 ( .A1(n12174), .A2(n7078), .ZN(n7072) );
  NAND2_X1 U8738 ( .A1(n12163), .A2(n12162), .ZN(n12310) );
  NAND2_X1 U8739 ( .A1(n7445), .A2(n7443), .ZN(n12318) );
  AND3_X1 U8740 ( .A1(n7987), .A2(n7986), .A3(n7985), .ZN(n11873) );
  NAND2_X1 U8741 ( .A1(n12174), .A2(n12173), .ZN(n12326) );
  OR2_X1 U8742 ( .A1(n10693), .A2(n10705), .ZN(n12328) );
  NAND2_X1 U8743 ( .A1(n10685), .A2(n10688), .ZN(n12360) );
  CLKBUF_X1 U8744 ( .A(n12332), .Z(n12356) );
  INV_X1 U8745 ( .A(n8523), .ZN(n12583) );
  OR2_X1 U8746 ( .A1(n7844), .A2(n7827), .ZN(n7830) );
  NAND4_X1 U8747 ( .A1(n7795), .A2(n7794), .A3(n7793), .A4(n7792), .ZN(n15202)
         );
  OR2_X1 U8748 ( .A1(n7844), .A2(n10360), .ZN(n7793) );
  INV_X1 U8749 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15157) );
  NAND2_X1 U8750 ( .A1(n7193), .A2(n10368), .ZN(n10536) );
  AOI22_X1 U8751 ( .A1(n10545), .A2(n10546), .B1(n10558), .B2(n10394), .ZN(
        n10512) );
  OAI22_X1 U8752 ( .A1(n10512), .A2(n10513), .B1(n10395), .B2(n10412), .ZN(
        n10397) );
  AND2_X1 U8753 ( .A1(n6677), .A2(n7211), .ZN(n11145) );
  INV_X1 U8754 ( .A(n11145), .ZN(n7209) );
  INV_X1 U8755 ( .A(n11150), .ZN(n7284) );
  NAND2_X1 U8756 ( .A1(n7198), .A2(n11385), .ZN(n15159) );
  INV_X1 U8757 ( .A(n15158), .ZN(n7196) );
  INV_X1 U8758 ( .A(n15160), .ZN(n7275) );
  AND2_X1 U8759 ( .A1(n6668), .A2(n7205), .ZN(n11749) );
  INV_X1 U8760 ( .A(n11749), .ZN(n7202) );
  NOR2_X1 U8761 ( .A1(n11751), .A2(n7967), .ZN(n7204) );
  NAND2_X1 U8762 ( .A1(n12400), .A2(n7188), .ZN(n12381) );
  NAND2_X1 U8763 ( .A1(n7189), .A2(n12414), .ZN(n7188) );
  INV_X1 U8764 ( .A(n12380), .ZN(n7189) );
  NOR2_X1 U8765 ( .A1(n12381), .A2(n8014), .ZN(n12401) );
  INV_X1 U8766 ( .A(n7517), .ZN(n12425) );
  INV_X1 U8767 ( .A(n7518), .ZN(n12404) );
  XNOR2_X1 U8768 ( .A(n12450), .B(n12456), .ZN(n12426) );
  AND2_X1 U8769 ( .A1(n8223), .A2(n8222), .ZN(n14515) );
  AND2_X1 U8770 ( .A1(n8200), .A2(n8190), .ZN(n12572) );
  NAND2_X1 U8771 ( .A1(n8166), .A2(n8165), .ZN(n12776) );
  OR2_X1 U8772 ( .A1(n7833), .A2(n12901), .ZN(n8165) );
  AND2_X1 U8773 ( .A1(n12599), .A2(n12598), .ZN(n12778) );
  NAND2_X1 U8774 ( .A1(n7680), .A2(n7677), .ZN(n12594) );
  NAND2_X1 U8775 ( .A1(n12623), .A2(n8515), .ZN(n12611) );
  NAND2_X1 U8776 ( .A1(n7321), .A2(n7320), .ZN(n12622) );
  NAND2_X1 U8777 ( .A1(n7323), .A2(n7322), .ZN(n7321) );
  NAND2_X1 U8778 ( .A1(n7325), .A2(n7328), .ZN(n12638) );
  NAND2_X1 U8779 ( .A1(n12671), .A2(n7329), .ZN(n7325) );
  AOI21_X1 U8780 ( .B1(n12671), .B2(n8511), .A(n7330), .ZN(n12650) );
  OAI21_X1 U8781 ( .B1(n12744), .B2(n12722), .A(n7299), .ZN(n12712) );
  NAND2_X1 U8782 ( .A1(n8506), .A2(n8505), .ZN(n12723) );
  NAND2_X1 U8783 ( .A1(n12744), .A2(n8356), .ZN(n12728) );
  NAND2_X1 U8784 ( .A1(n7313), .A2(n8345), .ZN(n12758) );
  NAND2_X1 U8785 ( .A1(n8003), .A2(n7314), .ZN(n7313) );
  NAND2_X1 U8786 ( .A1(n8501), .A2(n8500), .ZN(n14485) );
  NAND2_X1 U8787 ( .A1(n8003), .A2(n8341), .ZN(n14483) );
  AND2_X1 U8788 ( .A1(n11482), .A2(n8494), .ZN(n11706) );
  AND2_X1 U8789 ( .A1(n7674), .A2(n8491), .ZN(n11243) );
  INV_X1 U8790 ( .A(n12660), .ZN(n12761) );
  AND2_X1 U8791 ( .A1(n10977), .A2(n12531), .ZN(n15190) );
  AND2_X1 U8792 ( .A1(n11192), .A2(n15190), .ZN(n15209) );
  AND2_X1 U8793 ( .A1(n14513), .A2(n14514), .ZN(n14530) );
  INV_X1 U8794 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n7114) );
  AOI21_X1 U8795 ( .B1(n12896), .B2(n6474), .A(n6664), .ZN(n12836) );
  OR2_X1 U8796 ( .A1(n7833), .A2(n11824), .ZN(n8152) );
  INV_X1 U8797 ( .A(n12646), .ZN(n12849) );
  AOI21_X1 U8798 ( .B1(n10974), .B2(n6474), .A(n8108), .ZN(n12855) );
  NAND2_X1 U8799 ( .A1(n8028), .A2(n8027), .ZN(n12879) );
  AND3_X1 U8800 ( .A1(n7897), .A2(n7896), .A3(n7895), .ZN(n11647) );
  INV_X1 U8801 ( .A(n11196), .ZN(n10694) );
  AND2_X1 U8802 ( .A1(n8460), .A2(n8459), .ZN(n12882) );
  NAND2_X1 U8803 ( .A1(n10672), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12881) );
  AND2_X1 U8804 ( .A1(n6693), .A2(n6622), .ZN(n12884) );
  NAND2_X1 U8805 ( .A1(n10033), .A2(n8456), .ZN(n6693) );
  OAI211_X1 U8806 ( .C1(n8219), .C2(n7555), .A(n7552), .B(n7551), .ZN(n12890)
         );
  NAND2_X1 U8807 ( .A1(n7557), .A2(n7556), .ZN(n7555) );
  OAI21_X1 U8808 ( .B1(n8233), .B2(n7557), .A(n7553), .ZN(n7552) );
  AND2_X1 U8809 ( .A1(n6501), .A2(n7800), .ZN(n7699) );
  NAND2_X1 U8810 ( .A1(n7783), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7785) );
  AND2_X1 U8811 ( .A1(n7786), .A2(n7800), .ZN(n7782) );
  XNOR2_X1 U8812 ( .A(n8219), .B(n8208), .ZN(n12892) );
  AOI21_X1 U8813 ( .B1(n8129), .B2(n7547), .A(n7546), .ZN(n8151) );
  NAND2_X1 U8814 ( .A1(n8129), .A2(n7550), .ZN(n8141) );
  INV_X1 U8815 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8249) );
  XNOR2_X1 U8816 ( .A(n8128), .B(n8117), .ZN(n11083) );
  INV_X1 U8817 ( .A(SI_20_), .ZN(n10975) );
  INV_X1 U8818 ( .A(n9185), .ZN(n10977) );
  NAND2_X1 U8819 ( .A1(n7091), .A2(n7089), .ZN(n8106) );
  INV_X1 U8820 ( .A(SI_16_), .ZN(n10071) );
  NAND2_X1 U8821 ( .A1(n7096), .A2(n7094), .ZN(n8061) );
  INV_X1 U8822 ( .A(SI_15_), .ZN(n15386) );
  INV_X1 U8823 ( .A(SI_12_), .ZN(n9933) );
  NAND2_X1 U8824 ( .A1(n7107), .A2(n7997), .ZN(n8004) );
  NAND2_X1 U8825 ( .A1(n7995), .A2(n7994), .ZN(n7107) );
  INV_X1 U8826 ( .A(n12377), .ZN(n12382) );
  INV_X1 U8827 ( .A(SI_11_), .ZN(n9919) );
  NAND2_X1 U8828 ( .A1(n7102), .A2(n7947), .ZN(n7961) );
  NAND2_X1 U8829 ( .A1(n7945), .A2(n7944), .ZN(n7102) );
  NAND2_X1 U8830 ( .A1(n6729), .A2(n7873), .ZN(n7888) );
  NAND2_X1 U8831 ( .A1(n7872), .A2(n7871), .ZN(n6729) );
  NAND2_X1 U8832 ( .A1(n7537), .A2(n7836), .ZN(n7855) );
  NAND2_X1 U8833 ( .A1(n6496), .A2(n7523), .ZN(n10382) );
  AND2_X1 U8834 ( .A1(n13057), .A2(n12936), .ZN(n12941) );
  NAND2_X1 U8835 ( .A1(n13057), .A2(n7658), .ZN(n12967) );
  NAND2_X1 U8836 ( .A1(n9620), .A2(n9619), .ZN(n13225) );
  NAND2_X1 U8837 ( .A1(n11351), .A2(n11350), .ZN(n11461) );
  NAND2_X1 U8838 ( .A1(n9554), .A2(n9553), .ZN(n13518) );
  NAND2_X1 U8839 ( .A1(n7648), .A2(n7646), .ZN(n12979) );
  AND2_X1 U8840 ( .A1(n12980), .A2(n7647), .ZN(n7646) );
  INV_X1 U8841 ( .A(n7651), .ZN(n7647) );
  NOR2_X1 U8842 ( .A1(n13017), .A2(n7651), .ZN(n12981) );
  OAI21_X1 U8843 ( .B1(n13005), .B2(n12931), .A(n6598), .ZN(n13045) );
  OR2_X1 U8844 ( .A1(n13006), .A2(n12931), .ZN(n6722) );
  AND2_X1 U8845 ( .A1(n9659), .A2(n9658), .ZN(n13314) );
  NOR2_X1 U8846 ( .A1(n11842), .A2(n11843), .ZN(n12907) );
  NAND2_X1 U8847 ( .A1(n11842), .A2(n12906), .ZN(n7637) );
  NOR2_X1 U8848 ( .A1(n12907), .A2(n7641), .ZN(n13000) );
  NAND2_X1 U8849 ( .A1(n10483), .A2(n10448), .ZN(n10482) );
  NAND2_X1 U8850 ( .A1(n7649), .A2(n12958), .ZN(n13015) );
  NAND2_X1 U8851 ( .A1(n9567), .A2(n9566), .ZN(n13387) );
  NAND2_X1 U8852 ( .A1(n7632), .A2(n11655), .ZN(n11833) );
  NAND2_X1 U8853 ( .A1(n11654), .A2(n11653), .ZN(n7632) );
  NAND2_X1 U8854 ( .A1(n13026), .A2(n7759), .ZN(n13027) );
  XNOR2_X1 U8855 ( .A(n12919), .B(n6527), .ZN(n13026) );
  INV_X1 U8856 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n11361) );
  NAND2_X1 U8857 ( .A1(n9838), .A2(n14906), .ZN(n14911) );
  NAND2_X1 U8858 ( .A1(n6714), .A2(n7638), .ZN(n13036) );
  NAND2_X1 U8859 ( .A1(n11842), .A2(n7640), .ZN(n6714) );
  NAND2_X1 U8860 ( .A1(n10827), .A2(n10826), .ZN(n10829) );
  NAND2_X1 U8861 ( .A1(n13045), .A2(n7659), .ZN(n13057) );
  NAND2_X1 U8862 ( .A1(n9882), .A2(n9866), .ZN(n14903) );
  NAND2_X1 U8863 ( .A1(n9281), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9264) );
  AND2_X1 U8864 ( .A1(n6786), .A2(n6785), .ZN(n13463) );
  INV_X1 U8865 ( .A(n13276), .ZN(n6785) );
  NAND2_X1 U8866 ( .A1(n13287), .A2(n13286), .ZN(n13465) );
  NAND2_X1 U8867 ( .A1(n7379), .A2(n7380), .ZN(n13285) );
  NAND2_X1 U8868 ( .A1(n13320), .A2(n7381), .ZN(n7379) );
  NAND2_X1 U8869 ( .A1(n7383), .A2(n7385), .ZN(n13299) );
  OR2_X1 U8870 ( .A1(n13320), .A2(n13319), .ZN(n7383) );
  NAND2_X1 U8871 ( .A1(n7354), .A2(n7357), .ZN(n13329) );
  NAND2_X1 U8872 ( .A1(n7363), .A2(n7358), .ZN(n7354) );
  NAND2_X1 U8873 ( .A1(n6778), .A2(n6776), .ZN(n13341) );
  NOR2_X1 U8874 ( .A1(n6543), .A2(n7364), .ZN(n13339) );
  NAND2_X1 U8875 ( .A1(n13223), .A2(n7396), .ZN(n13350) );
  NAND2_X1 U8876 ( .A1(n9536), .A2(n9535), .ZN(n13424) );
  NAND2_X1 U8877 ( .A1(n9513), .A2(n9512), .ZN(n13533) );
  NAND2_X1 U8878 ( .A1(n7388), .A2(n7392), .ZN(n13433) );
  NAND2_X1 U8879 ( .A1(n11934), .A2(n11933), .ZN(n13212) );
  NAND2_X1 U8880 ( .A1(n11724), .A2(n11723), .ZN(n11880) );
  NAND2_X1 U8881 ( .A1(n6792), .A2(n11331), .ZN(n11334) );
  NAND2_X1 U8882 ( .A1(n7365), .A2(n6492), .ZN(n11609) );
  NAND2_X1 U8883 ( .A1(n6545), .A2(n11255), .ZN(n7365) );
  NAND2_X1 U8884 ( .A1(n11255), .A2(n11254), .ZN(n11343) );
  NAND2_X1 U8885 ( .A1(n11258), .A2(n11257), .ZN(n11330) );
  NAND2_X1 U8886 ( .A1(n11129), .A2(n11128), .ZN(n11132) );
  NAND2_X1 U8887 ( .A1(n6773), .A2(n10998), .ZN(n11127) );
  NAND2_X1 U8888 ( .A1(n10995), .A2(n10994), .ZN(n6773) );
  NAND2_X1 U8889 ( .A1(n7348), .A2(n10656), .ZN(n10749) );
  INV_X1 U8890 ( .A(n15055), .ZN(n14556) );
  NAND2_X1 U8891 ( .A1(n13427), .A2(n10567), .ZN(n15059) );
  AND2_X1 U8892 ( .A1(n10571), .A2(n10572), .ZN(n6765) );
  AND2_X2 U8893 ( .A1(n10621), .A2(n10211), .ZN(n15145) );
  INV_X1 U8894 ( .A(n7176), .ZN(n7175) );
  OAI21_X1 U8895 ( .B1(n13453), .B2(n15114), .A(n13451), .ZN(n7176) );
  OR2_X1 U8896 ( .A1(n13509), .A2(n13508), .ZN(n13560) );
  AND2_X1 U8897 ( .A1(n9873), .A2(n9824), .ZN(n15082) );
  AND2_X1 U8898 ( .A1(n7721), .A2(n9236), .ZN(n7720) );
  NAND2_X1 U8899 ( .A1(n6976), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9237) );
  NAND2_X1 U8900 ( .A1(n9209), .A2(n7721), .ZN(n6976) );
  XNOR2_X1 U8901 ( .A(n9820), .B(P2_IR_REG_26__SCAN_IN), .ZN(n13586) );
  XNOR2_X1 U8902 ( .A(n9822), .B(P2_IR_REG_25__SCAN_IN), .ZN(n13591) );
  XNOR2_X1 U8903 ( .A(n9819), .B(P2_IR_REG_24__SCAN_IN), .ZN(n13595) );
  INV_X1 U8904 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11796) );
  AND2_X1 U8905 ( .A1(n9676), .A2(P2_U3088), .ZN(n11792) );
  INV_X1 U8906 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11717) );
  INV_X1 U8907 ( .A(n9747), .ZN(n11439) );
  INV_X1 U8908 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9904) );
  NOR2_X1 U8909 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n9287) );
  NAND2_X1 U8910 ( .A1(n13839), .A2(n13692), .ZN(n13728) );
  NAND2_X1 U8911 ( .A1(n10797), .A2(n10796), .ZN(n13738) );
  AND2_X1 U8912 ( .A1(n6936), .A2(n6542), .ZN(n13748) );
  NAND2_X1 U8913 ( .A1(n6936), .A2(n6934), .ZN(n13746) );
  AND2_X1 U8914 ( .A1(n6941), .A2(n14623), .ZN(n6940) );
  NAND2_X1 U8915 ( .A1(n6942), .A2(n6946), .ZN(n6941) );
  NAND2_X1 U8916 ( .A1(n7742), .A2(n13655), .ZN(n13802) );
  NAND2_X1 U8917 ( .A1(n14603), .A2(n14602), .ZN(n7742) );
  OAI21_X1 U8918 ( .B1(n13770), .B2(n6957), .A(n6954), .ZN(n13812) );
  OR2_X1 U8919 ( .A1(n11541), .A2(n7745), .ZN(n11776) );
  NAND2_X1 U8920 ( .A1(n6932), .A2(n6935), .ZN(n6930) );
  NAND2_X1 U8921 ( .A1(n6929), .A2(n6932), .ZN(n13823) );
  OR2_X1 U8922 ( .A1(n13852), .A2(n6935), .ZN(n6929) );
  INV_X1 U8923 ( .A(n13833), .ZN(n6973) );
  INV_X1 U8924 ( .A(n6974), .ZN(n13834) );
  NAND2_X1 U8925 ( .A1(n6926), .A2(n11532), .ZN(n6923) );
  OAI211_X1 U8926 ( .C1(n6925), .C2(n11532), .A(n6924), .B(n11781), .ZN(n14610) );
  NAND2_X1 U8927 ( .A1(n7743), .A2(n7745), .ZN(n6924) );
  INV_X1 U8928 ( .A(n7743), .ZN(n6925) );
  NAND2_X1 U8929 ( .A1(n10273), .A2(n10274), .ZN(n10797) );
  NAND2_X1 U8930 ( .A1(n8881), .A2(n8880), .ZN(n14257) );
  AND2_X1 U8931 ( .A1(n11043), .A2(n11042), .ZN(n6991) );
  NAND2_X1 U8932 ( .A1(n7726), .A2(n13713), .ZN(n13858) );
  XNOR2_X1 U8933 ( .A(n13645), .B(n13646), .ZN(n14619) );
  NAND2_X1 U8934 ( .A1(n14619), .A2(n14620), .ZN(n14618) );
  AND2_X1 U8935 ( .A1(n10181), .A2(n10180), .ZN(n14621) );
  NAND2_X1 U8936 ( .A1(n10791), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14629) );
  OAI21_X1 U8937 ( .B1(n12152), .B2(n7761), .A(n12151), .ZN(n7471) );
  XNOR2_X1 U8938 ( .A(n10084), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n10151) );
  NOR2_X1 U8939 ( .A1(n10135), .A2(n10134), .ZN(n10163) );
  NOR2_X1 U8940 ( .A1(n10132), .A2(n7167), .ZN(n10135) );
  AND2_X1 U8941 ( .A1(n10137), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7167) );
  AOI21_X1 U8942 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n10164), .A(n10157), .ZN(
        n10160) );
  NOR2_X1 U8943 ( .A1(n10468), .A2(n6639), .ZN(n10471) );
  AOI21_X1 U8944 ( .B1(n11033), .B2(P1_REG1_REG_10__SCAN_IN), .A(n11023), .ZN(
        n14679) );
  OR2_X1 U8945 ( .A1(n13913), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7050) );
  NAND2_X1 U8946 ( .A1(n14741), .A2(n14740), .ZN(n14739) );
  OAI211_X1 U8947 ( .C1(n13977), .C2(n6903), .A(n6900), .B(n6897), .ZN(n13958)
         );
  NAND2_X1 U8948 ( .A1(n12141), .A2(n6985), .ZN(n6903) );
  OAI21_X1 U8949 ( .B1(n6902), .B2(n12141), .A(n6901), .ZN(n6900) );
  NAND2_X1 U8950 ( .A1(n13977), .A2(n6898), .ZN(n6897) );
  NAND2_X1 U8951 ( .A1(n13977), .A2(n9118), .ZN(n13961) );
  NAND2_X1 U8952 ( .A1(n9021), .A2(n9020), .ZN(n13982) );
  AND2_X1 U8953 ( .A1(n9046), .A2(n9031), .ZN(n13991) );
  NAND2_X1 U8954 ( .A1(n14028), .A2(n9113), .ZN(n14009) );
  AND2_X1 U8955 ( .A1(n7579), .A2(n7581), .ZN(n14021) );
  NAND2_X1 U8956 ( .A1(n7584), .A2(n8967), .ZN(n14031) );
  AOI21_X1 U8957 ( .B1(n14072), .B2(n14073), .A(n9108), .ZN(n14056) );
  NAND2_X1 U8958 ( .A1(n14102), .A2(n12039), .ZN(n14084) );
  NAND2_X1 U8959 ( .A1(n6884), .A2(n8908), .ZN(n14097) );
  NAND2_X1 U8960 ( .A1(n8864), .A2(n8863), .ZN(n14264) );
  NAND2_X1 U8961 ( .A1(n10465), .A2(n12087), .ZN(n8864) );
  NAND2_X1 U8962 ( .A1(n14145), .A2(n9100), .ZN(n14132) );
  NAND2_X1 U8963 ( .A1(n11850), .A2(n6490), .ZN(n11812) );
  NAND2_X1 U8964 ( .A1(n11855), .A2(n12008), .ZN(n11811) );
  OAI21_X1 U8965 ( .B1(n10942), .B2(n7567), .A(n7566), .ZN(n10866) );
  NAND2_X1 U8966 ( .A1(n10941), .A2(n8682), .ZN(n10867) );
  NAND2_X1 U8967 ( .A1(n9089), .A2(n9088), .ZN(n11092) );
  NAND2_X1 U8968 ( .A1(n7572), .A2(n7570), .ZN(n10906) );
  NAND2_X1 U8969 ( .A1(n8609), .A2(n8608), .ZN(n10938) );
  OR2_X1 U8970 ( .A1(n13950), .A2(n13930), .ZN(n14818) );
  NAND2_X1 U8971 ( .A1(n10177), .A2(n10192), .ZN(n14831) );
  OR2_X1 U8972 ( .A1(n14842), .A2(n10854), .ZN(n14161) );
  INV_X1 U8973 ( .A(n14845), .ZN(n14814) );
  OR2_X1 U8974 ( .A1(n10258), .A2(n11950), .ZN(n12118) );
  INV_X1 U8975 ( .A(n14143), .ZN(n14146) );
  INV_X1 U8976 ( .A(n10259), .ZN(n10888) );
  INV_X1 U8977 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7003) );
  INV_X1 U8978 ( .A(n13942), .ZN(n14286) );
  INV_X1 U8979 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n7589) );
  NAND2_X1 U8980 ( .A1(n8763), .A2(n8762), .ZN(n13791) );
  NAND2_X1 U8981 ( .A1(n8746), .A2(n8745), .ZN(n14630) );
  INV_X1 U8982 ( .A(n11995), .ZN(n14787) );
  INV_X1 U8983 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14330) );
  AND2_X1 U8984 ( .A1(n14320), .A2(n6611), .ZN(n7568) );
  OR2_X1 U8985 ( .A1(n8559), .A2(n8544), .ZN(n7039) );
  NOR2_X1 U8986 ( .A1(n8547), .A2(n7038), .ZN(n7037) );
  NAND2_X1 U8987 ( .A1(n6833), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8562) );
  INV_X1 U8988 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14342) );
  NOR2_X1 U8989 ( .A1(n9076), .A2(n7056), .ZN(n7055) );
  INV_X1 U8990 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11369) );
  INV_X1 U8991 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8814) );
  XNOR2_X1 U8992 ( .A(n8796), .B(P1_IR_REG_14__SCAN_IN), .ZN(n14708) );
  AND2_X1 U8993 ( .A1(n8795), .A2(n8781), .ZN(n14699) );
  OAI21_X1 U8994 ( .B1(n8726), .B2(n8725), .A(n8739), .ZN(n9961) );
  OR2_X1 U8995 ( .A1(n8705), .A2(n8704), .ZN(n8706) );
  NAND2_X1 U8996 ( .A1(n8684), .A2(n8683), .ZN(n8688) );
  NOR2_X1 U8997 ( .A1(n8670), .A2(n6890), .ZN(n6889) );
  INV_X1 U8998 ( .A(n8666), .ZN(n6890) );
  INV_X1 U8999 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9926) );
  NAND2_X1 U9000 ( .A1(n8649), .A2(n8648), .ZN(n8653) );
  INV_X1 U9001 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9917) );
  NAND2_X1 U9002 ( .A1(n8649), .A2(n6814), .ZN(n9916) );
  NAND2_X1 U9003 ( .A1(n6816), .A2(n8633), .ZN(n6814) );
  INV_X1 U9005 ( .A(n8635), .ZN(n6816) );
  OR2_X1 U9006 ( .A1(n8621), .A2(n6529), .ZN(n8622) );
  OR2_X1 U9007 ( .A1(n8600), .A2(n6559), .ZN(n8601) );
  INV_X1 U9008 ( .A(n6893), .ZN(n8582) );
  NAND2_X1 U9009 ( .A1(n7604), .A2(n8579), .ZN(n8571) );
  INV_X1 U9010 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7052) );
  NAND2_X1 U9011 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n7174) );
  OAI21_X1 U9012 ( .B1(n14409), .B2(n13105), .A(n15452), .ZN(n15445) );
  XNOR2_X1 U9013 ( .A(n14400), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15446) );
  XNOR2_X1 U9014 ( .A(n14414), .B(n7515), .ZN(n14457) );
  XNOR2_X1 U9015 ( .A(n14419), .B(n7066), .ZN(n15450) );
  OAI21_X1 U9016 ( .B1(n14460), .B2(n14461), .A(P2_ADDR_REG_9__SCAN_IN), .ZN(
        n7068) );
  AND2_X1 U9017 ( .A1(n14428), .A2(n14427), .ZN(n14649) );
  NOR2_X1 U9018 ( .A1(n14435), .A2(n14434), .ZN(n14656) );
  AND2_X1 U9019 ( .A1(n6762), .A2(n6761), .ZN(n14469) );
  NOR2_X1 U9020 ( .A1(n14469), .A2(n14468), .ZN(n14467) );
  NAND2_X1 U9021 ( .A1(n6686), .A2(n6684), .ZN(P3_U3154) );
  AND2_X1 U9022 ( .A1(n12229), .A2(n6685), .ZN(n6684) );
  NAND2_X1 U9023 ( .A1(n6687), .A2(n12340), .ZN(n6686) );
  NAND2_X1 U9024 ( .A1(n12575), .A2(n12334), .ZN(n6685) );
  OAI21_X1 U9025 ( .B1(n7026), .B2(n8434), .A(n8433), .ZN(n8454) );
  INV_X1 U9026 ( .A(n7225), .ZN(n12454) );
  NOR2_X1 U9027 ( .A1(n12505), .A2(n12504), .ZN(n12529) );
  NAND2_X1 U9028 ( .A1(n7221), .A2(n12547), .ZN(n6999) );
  NOR2_X1 U9029 ( .A1(n9191), .A2(n6494), .ZN(n7683) );
  AND2_X1 U9030 ( .A1(n7686), .A2(n7685), .ZN(n7684) );
  NAND2_X1 U9031 ( .A1(n6813), .A2(n6812), .ZN(P3_U3487) );
  AOI21_X1 U9032 ( .B1(n12767), .B2(n12823), .A(n6667), .ZN(n6812) );
  NAND2_X1 U9033 ( .A1(n12765), .A2(n15254), .ZN(n6813) );
  NAND2_X1 U9034 ( .A1(n6731), .A2(n6730), .ZN(n12770) );
  NAND2_X1 U9035 ( .A1(n12766), .A2(n15259), .ZN(n6730) );
  NAND2_X1 U9036 ( .A1(n12830), .A2(n15254), .ZN(n6731) );
  INV_X1 U9037 ( .A(n7295), .ZN(n7294) );
  OAI21_X1 U9038 ( .B1(n7687), .B2(n15244), .A(n9177), .ZN(n7295) );
  NAND2_X1 U9039 ( .A1(n7115), .A2(n7112), .ZN(P3_U3455) );
  INV_X1 U9040 ( .A(n7113), .ZN(n7112) );
  NAND2_X1 U9041 ( .A1(n12765), .A2(n15246), .ZN(n7115) );
  OAI22_X1 U9042 ( .A1(n8534), .A2(n12880), .B1(n15246), .B2(n7114), .ZN(n7113) );
  INV_X1 U9043 ( .A(n6995), .ZN(n6994) );
  OAI22_X1 U9044 ( .A1(n12832), .A2(n12880), .B1(n15246), .B2(n12831), .ZN(
        n6995) );
  OAI21_X1 U9045 ( .B1(n11654), .B2(n7631), .A(n7626), .ZN(n14545) );
  OR2_X1 U9046 ( .A1(n15145), .A2(n7352), .ZN(n7351) );
  INV_X1 U9047 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7352) );
  NAND2_X1 U9048 ( .A1(n15132), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7262) );
  AOI21_X1 U9049 ( .B1(n7172), .B2(n13930), .A(n7171), .ZN(n7170) );
  OAI21_X1 U9050 ( .B1(n14781), .B2(n7591), .A(n13933), .ZN(n7171) );
  INV_X1 U9051 ( .A(n7041), .ZN(n7040) );
  OAI21_X1 U9052 ( .B1(n14282), .B2(n14210), .A(n7042), .ZN(n7041) );
  AOI21_X1 U9053 ( .B1(n14180), .B2(n14230), .A(n6676), .ZN(n7465) );
  NAND2_X1 U9054 ( .A1(n7004), .A2(n7002), .ZN(n7001) );
  OR2_X1 U9055 ( .A1(n14896), .A2(n7003), .ZN(n7002) );
  OAI21_X1 U9056 ( .B1(n14280), .B2(n14889), .A(n6822), .ZN(P1_U3527) );
  AOI21_X1 U9057 ( .B1(n12107), .B2(n14306), .A(n6823), .ZN(n6822) );
  NOR2_X1 U9058 ( .A1(n14891), .A2(n14281), .ZN(n6823) );
  OR2_X1 U9059 ( .A1(n14891), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7058) );
  NAND2_X1 U9060 ( .A1(n7590), .A2(n6970), .ZN(P1_U3524) );
  NOR2_X1 U9061 ( .A1(n6986), .A2(n6674), .ZN(n6970) );
  NAND2_X1 U9062 ( .A1(n14287), .A2(n14891), .ZN(n7590) );
  INV_X1 U9063 ( .A(n6763), .ZN(n14652) );
  INV_X1 U9064 ( .A(n7510), .ZN(n14660) );
  AND2_X1 U9065 ( .A1(n7503), .A2(n7510), .ZN(n14664) );
  NAND2_X1 U9066 ( .A1(n7505), .A2(n7500), .ZN(n14662) );
  NAND2_X2 U9067 ( .A1(n11948), .A2(n12093), .ZN(n12002) );
  NAND2_X2 U9068 ( .A1(n6489), .A2(n9247), .ZN(n10457) );
  AND2_X1 U9069 ( .A1(n8831), .A2(n8809), .ZN(n6490) );
  AND3_X1 U9070 ( .A1(n8816), .A2(n7562), .A3(n7561), .ZN(n6491) );
  INV_X1 U9071 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8672) );
  NAND2_X4 U9072 ( .A1(n6692), .A2(n10711), .ZN(n10712) );
  INV_X1 U9073 ( .A(n6474), .ZN(n8055) );
  NAND2_X1 U9074 ( .A1(n8199), .A2(n8198), .ZN(n12767) );
  AND2_X1 U9075 ( .A1(n12008), .A2(n12019), .ZN(n12133) );
  OR2_X1 U9076 ( .A1(n11465), .A2(n13081), .ZN(n6492) );
  AND2_X1 U9077 ( .A1(n7412), .A2(n12308), .ZN(n6493) );
  NOR2_X1 U9078 ( .A1(n9192), .A2(n12829), .ZN(n6494) );
  AND2_X1 U9079 ( .A1(n7521), .A2(n7520), .ZN(n6496) );
  NOR2_X1 U9080 ( .A1(n13225), .A2(n12921), .ZN(n6497) );
  OAI211_X1 U9081 ( .C1(n7833), .C2(SI_3_), .A(n7842), .B(n7841), .ZN(n11640)
         );
  INV_X1 U9082 ( .A(n11640), .ZN(n6968) );
  AND2_X1 U9083 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n6498) );
  OR2_X1 U9084 ( .A1(n12590), .A2(n8517), .ZN(n8261) );
  AND2_X1 U9085 ( .A1(n7491), .A2(n12096), .ZN(n6499) );
  AND2_X1 U9086 ( .A1(n6583), .A2(n7150), .ZN(n6500) );
  NAND3_X1 U9087 ( .A1(n7443), .A2(n12656), .A3(n7445), .ZN(n12317) );
  AND2_X1 U9088 ( .A1(n7781), .A2(n7802), .ZN(n6501) );
  AND2_X1 U9089 ( .A1(n14288), .A2(n13872), .ZN(n6502) );
  AND2_X1 U9090 ( .A1(n8542), .A2(n8561), .ZN(n6503) );
  NAND2_X1 U9091 ( .A1(n8959), .A2(n8958), .ZN(n14221) );
  OR2_X1 U9092 ( .A1(n7445), .A2(n7084), .ZN(n6504) );
  AND2_X1 U9093 ( .A1(n6495), .A2(n6817), .ZN(n6505) );
  AND2_X1 U9094 ( .A1(n8624), .A2(n8540), .ZN(n6506) );
  NAND2_X2 U9095 ( .A1(n11952), .A2(n10185), .ZN(n13687) );
  AND2_X1 U9096 ( .A1(n6886), .A2(n6585), .ZN(n6507) );
  OR2_X1 U9097 ( .A1(n12776), .A2(n12614), .ZN(n8264) );
  AND2_X1 U9098 ( .A1(n6606), .A2(n6857), .ZN(n6508) );
  INV_X1 U9099 ( .A(n12107), .ZN(n14282) );
  OR2_X1 U9100 ( .A1(n12767), .A2(n12226), .ZN(n8393) );
  INV_X1 U9101 ( .A(n10929), .ZN(n7571) );
  INV_X1 U9102 ( .A(n7645), .ZN(n13013) );
  NAND2_X1 U9103 ( .A1(n6707), .A2(n6710), .ZN(n7645) );
  AND2_X1 U9104 ( .A1(n9917), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n6509) );
  INV_X1 U9105 ( .A(n12066), .ZN(n6858) );
  NAND2_X1 U9106 ( .A1(n14351), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n6510) );
  INV_X1 U9107 ( .A(n14622), .ZN(n7233) );
  INV_X1 U9108 ( .A(n12004), .ZN(n6981) );
  OR2_X1 U9109 ( .A1(n8394), .A2(n7334), .ZN(n6511) );
  AND2_X1 U9110 ( .A1(n7213), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n6512) );
  NAND2_X1 U9111 ( .A1(n6942), .A2(n6628), .ZN(n6513) );
  INV_X1 U9112 ( .A(n7328), .ZN(n7327) );
  AND2_X1 U9113 ( .A1(n7116), .A2(n8272), .ZN(n7328) );
  XOR2_X1 U9114 ( .A(n14604), .B(n13805), .Z(n6514) );
  INV_X1 U9115 ( .A(n12137), .ZN(n6960) );
  INV_X1 U9116 ( .A(n11751), .ZN(n7206) );
  INV_X1 U9117 ( .A(n6830), .ZN(n14103) );
  NOR2_X1 U9118 ( .A1(n14121), .A2(n14251), .ZN(n6830) );
  NOR2_X1 U9119 ( .A1(n14148), .A2(n14604), .ZN(n7232) );
  NAND2_X1 U9120 ( .A1(n8350), .A2(n8354), .ZN(n6515) );
  INV_X1 U9121 ( .A(n12575), .ZN(n12832) );
  NAND2_X1 U9122 ( .A1(n8188), .A2(n8187), .ZN(n12575) );
  AND2_X1 U9123 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n7533), .ZN(n6516) );
  NAND2_X1 U9124 ( .A1(n11472), .A2(n6825), .ZN(n6517) );
  AND2_X1 U9125 ( .A1(n7199), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n6518) );
  AND2_X1 U9126 ( .A1(n7278), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n6519) );
  NAND2_X1 U9127 ( .A1(n7063), .A2(n6678), .ZN(n6520) );
  INV_X1 U9128 ( .A(n14559), .ZN(n7182) );
  INV_X1 U9129 ( .A(n12906), .ZN(n7641) );
  NAND2_X1 U9130 ( .A1(n14325), .A2(n8551), .ZN(n8918) );
  AND2_X1 U9131 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n7005), .ZN(n6521) );
  AND2_X1 U9132 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n10446), .ZN(n6522) );
  NAND2_X1 U9133 ( .A1(n7625), .A2(n9247), .ZN(n10200) );
  INV_X1 U9134 ( .A(n11979), .ZN(n7227) );
  OR2_X1 U9135 ( .A1(n10602), .A2(n7215), .ZN(n6523) );
  AND2_X1 U9136 ( .A1(n14330), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6524) );
  AND2_X1 U9137 ( .A1(n9242), .A2(n13577), .ZN(n6525) );
  INV_X1 U9138 ( .A(n7745), .ZN(n7744) );
  NAND2_X1 U9139 ( .A1(n11547), .A2(n7746), .ZN(n7745) );
  XOR2_X1 U9140 ( .A(n13501), .B(n12968), .Z(n6527) );
  INV_X1 U9141 ( .A(n9540), .ZN(n9589) );
  INV_X1 U9142 ( .A(n12372), .ZN(n6690) );
  NAND2_X1 U9143 ( .A1(n12625), .A2(n12624), .ZN(n12623) );
  NAND2_X1 U9144 ( .A1(n7697), .A2(n6495), .ZN(n7932) );
  INV_X1 U9145 ( .A(n14115), .ZN(n7483) );
  INV_X1 U9146 ( .A(n11210), .ZN(n6691) );
  AND2_X1 U9147 ( .A1(n8876), .A2(n10354), .ZN(n6528) );
  NAND3_X2 U9148 ( .A1(n10204), .A2(n9806), .A3(n9880), .ZN(n9413) );
  NOR2_X1 U9149 ( .A1(n7893), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n7911) );
  NAND2_X1 U9150 ( .A1(n9194), .A2(n9193), .ZN(n9256) );
  AND2_X1 U9151 ( .A1(n12223), .A2(n12895), .ZN(n7843) );
  INV_X1 U9152 ( .A(n7843), .ZN(n8215) );
  AND2_X1 U9153 ( .A1(n8630), .A2(n6808), .ZN(n6529) );
  NAND2_X1 U9154 ( .A1(n13005), .A2(n13006), .ZN(n6530) );
  OR2_X1 U9155 ( .A1(n12492), .A2(n12493), .ZN(n6531) );
  INV_X1 U9156 ( .A(n13260), .ZN(n7029) );
  INV_X1 U9157 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7397) );
  AND2_X1 U9158 ( .A1(n6514), .A2(n12026), .ZN(n6532) );
  NAND4_X1 U9159 ( .A1(n7808), .A2(n7807), .A3(n7806), .A4(n7805), .ZN(n12374)
         );
  NAND3_X1 U9160 ( .A1(n8590), .A2(n8591), .A3(n8589), .ZN(n10276) );
  AND2_X1 U9161 ( .A1(n9250), .A2(n9249), .ZN(n6533) );
  AND2_X1 U9162 ( .A1(n9404), .A2(n9403), .ZN(n6534) );
  AND2_X1 U9163 ( .A1(n9470), .A2(n9469), .ZN(n6535) );
  AND2_X1 U9164 ( .A1(n6845), .A2(n12051), .ZN(n6536) );
  NOR2_X1 U9165 ( .A1(n14211), .A2(n13876), .ZN(n6537) );
  NOR2_X1 U9166 ( .A1(n14065), .A2(n13878), .ZN(n6538) );
  NAND2_X1 U9167 ( .A1(n7481), .A2(n11981), .ZN(n6539) );
  XNOR2_X1 U9168 ( .A(n11979), .B(n11114), .ZN(n12124) );
  INV_X1 U9169 ( .A(n12124), .ZN(n6885) );
  NAND2_X1 U9170 ( .A1(n14618), .A2(n13648), .ZN(n14603) );
  AND2_X1 U9171 ( .A1(n7832), .A2(n7831), .ZN(n6540) );
  NAND2_X1 U9172 ( .A1(n13756), .A2(n13755), .ZN(n6541) );
  OR2_X1 U9173 ( .A1(n13668), .A2(n13667), .ZN(n6542) );
  INV_X1 U9174 ( .A(n6935), .ZN(n6934) );
  NAND2_X1 U9175 ( .A1(n13747), .A2(n6542), .ZN(n6935) );
  NAND3_X1 U9176 ( .A1(n6540), .A2(n7830), .A3(n7829), .ZN(n10960) );
  INV_X1 U9177 ( .A(n10960), .ZN(n6969) );
  AND2_X1 U9178 ( .A1(n7363), .A2(n7362), .ZN(n6543) );
  AND2_X1 U9179 ( .A1(n9261), .A2(n9260), .ZN(n6544) );
  NOR2_X1 U9180 ( .A1(n11342), .A2(n7369), .ZN(n6545) );
  NOR4_X1 U9181 ( .A1(n9794), .A2(n13429), .A3(n14557), .A4(n11922), .ZN(n6546) );
  AND2_X1 U9182 ( .A1(n6756), .A2(n6510), .ZN(n6547) );
  NAND2_X1 U9183 ( .A1(n6757), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n6548) );
  AND3_X1 U9184 ( .A1(n7936), .A2(n7935), .A3(n7934), .ZN(n11664) );
  INV_X1 U9185 ( .A(n11664), .ZN(n7086) );
  INV_X1 U9186 ( .A(n9167), .ZN(n9174) );
  AND2_X1 U9187 ( .A1(n8403), .A2(n8402), .ZN(n9167) );
  NAND2_X1 U9188 ( .A1(n9584), .A2(n9583), .ZN(n13375) );
  INV_X1 U9189 ( .A(n13375), .ZN(n6818) );
  AND2_X1 U9190 ( .A1(n10412), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U9191 ( .A1(n7752), .A2(n8584), .ZN(n8603) );
  OR2_X1 U9192 ( .A1(n13087), .A2(n15105), .ZN(n6550) );
  INV_X1 U9193 ( .A(n13469), .ZN(n7185) );
  NAND2_X2 U9194 ( .A1(n8551), .A2(n8550), .ZN(n8915) );
  XNOR2_X1 U9195 ( .A(n8874), .B(n8861), .ZN(n10465) );
  NAND2_X1 U9196 ( .A1(n8783), .A2(n8782), .ZN(n13837) );
  AND2_X1 U9197 ( .A1(n14573), .A2(n14542), .ZN(n6551) );
  OR2_X1 U9198 ( .A1(n9290), .A2(n13103), .ZN(n6552) );
  AND2_X1 U9199 ( .A1(n14288), .A2(n9119), .ZN(n6553) );
  NAND2_X1 U9200 ( .A1(n7815), .A2(n7814), .ZN(n8407) );
  NAND2_X1 U9201 ( .A1(n7693), .A2(n7691), .ZN(n12651) );
  AND2_X1 U9202 ( .A1(n8393), .A2(n8259), .ZN(n8527) );
  AND2_X1 U9203 ( .A1(n9775), .A2(n9774), .ZN(n6554) );
  INV_X1 U9204 ( .A(n14096), .ZN(n8922) );
  INV_X1 U9205 ( .A(n11978), .ZN(n6856) );
  INV_X1 U9206 ( .A(n11994), .ZN(n7476) );
  NAND2_X1 U9207 ( .A1(n11905), .A2(n11904), .ZN(n6555) );
  OR2_X1 U9208 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n8115), .ZN(n6556) );
  AND2_X1 U9209 ( .A1(n13822), .A2(n6930), .ZN(n6557) );
  OR2_X1 U9210 ( .A1(n15122), .A2(n13080), .ZN(n6558) );
  NOR2_X1 U9211 ( .A1(n13317), .A2(n13252), .ZN(n7374) );
  AND2_X1 U9212 ( .A1(n8619), .A2(n6983), .ZN(n6559) );
  NAND2_X1 U9213 ( .A1(n8899), .A2(n7497), .ZN(n9073) );
  OR2_X1 U9214 ( .A1(n13494), .A2(n13226), .ZN(n6560) );
  OR2_X1 U9215 ( .A1(n12925), .A2(n12924), .ZN(n6561) );
  NOR2_X1 U9216 ( .A1(n13538), .A2(n13210), .ZN(n6562) );
  AND2_X1 U9217 ( .A1(n9392), .A2(n9391), .ZN(n6563) );
  NAND2_X1 U9218 ( .A1(n7442), .A2(n7016), .ZN(n7890) );
  NOR2_X1 U9219 ( .A1(n14573), .A2(n14542), .ZN(n6564) );
  INV_X1 U9220 ( .A(n9194), .ZN(n9311) );
  AND2_X1 U9221 ( .A1(n9421), .A2(n9420), .ZN(n6565) );
  AND2_X1 U9222 ( .A1(n12179), .A2(n12692), .ZN(n6566) );
  NAND2_X1 U9223 ( .A1(n8389), .A2(n8525), .ZN(n12567) );
  INV_X1 U9224 ( .A(n12567), .ZN(n6753) );
  AND2_X1 U9225 ( .A1(n6499), .A2(n12082), .ZN(n6567) );
  AND2_X1 U9226 ( .A1(n8153), .A2(n8152), .ZN(n12841) );
  INV_X1 U9227 ( .A(n7186), .ZN(n13302) );
  AND2_X1 U9228 ( .A1(n11976), .A2(n9090), .ZN(n6568) );
  NOR2_X1 U9229 ( .A1(n12575), .A2(n12583), .ZN(n6569) );
  AND2_X1 U9230 ( .A1(n6550), .A2(n10656), .ZN(n6570) );
  AND2_X1 U9231 ( .A1(n7696), .A2(n8508), .ZN(n6571) );
  INV_X1 U9232 ( .A(n7576), .ZN(n7575) );
  NAND2_X1 U9233 ( .A1(n9036), .A2(n9020), .ZN(n7576) );
  AND2_X1 U9234 ( .A1(n7070), .A2(n12181), .ZN(n6572) );
  INV_X1 U9235 ( .A(n7324), .ZN(n7322) );
  NAND2_X1 U9236 ( .A1(n7328), .A2(n7331), .ZN(n7324) );
  INV_X1 U9237 ( .A(n12621), .ZN(n12624) );
  AND2_X1 U9238 ( .A1(n8922), .A2(n8908), .ZN(n6573) );
  AND2_X1 U9239 ( .A1(n13682), .A2(n13680), .ZN(n6574) );
  AND2_X1 U9240 ( .A1(n6499), .A2(n12078), .ZN(n6575) );
  INV_X1 U9241 ( .A(n6985), .ZN(n6906) );
  AND2_X1 U9242 ( .A1(n11332), .A2(n11331), .ZN(n6576) );
  INV_X1 U9243 ( .A(n7453), .ZN(n7452) );
  NOR2_X1 U9244 ( .A1(n9102), .A2(n7454), .ZN(n7453) );
  AND2_X1 U9245 ( .A1(n9398), .A2(n9397), .ZN(n6577) );
  OR2_X1 U9246 ( .A1(n7185), .A2(n13258), .ZN(n6578) );
  INV_X1 U9247 ( .A(n7669), .ZN(n7668) );
  OR2_X1 U9248 ( .A1(n8507), .A2(n7670), .ZN(n7669) );
  OR2_X1 U9249 ( .A1(n6856), .A2(n11977), .ZN(n6579) );
  AND2_X1 U9250 ( .A1(n6908), .A2(n7453), .ZN(n6580) );
  AND2_X1 U9251 ( .A1(n13698), .A2(n13697), .ZN(n6581) );
  AND2_X1 U9252 ( .A1(n13720), .A2(n13719), .ZN(n6582) );
  NAND2_X1 U9253 ( .A1(n13249), .A2(n7360), .ZN(n7357) );
  AND2_X1 U9254 ( .A1(n8322), .A2(n8321), .ZN(n11485) );
  INV_X1 U9255 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n9226) );
  INV_X1 U9256 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7802) );
  INV_X1 U9257 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8561) );
  INV_X1 U9258 ( .A(n14065), .ZN(n14305) );
  INV_X1 U9259 ( .A(n12633), .ZN(n12845) );
  NAND2_X1 U9260 ( .A1(n8143), .A2(n8142), .ZN(n12633) );
  OR2_X1 U9261 ( .A1(n6533), .A2(n9474), .ZN(n6583) );
  AND2_X1 U9262 ( .A1(n8272), .A2(n8271), .ZN(n12654) );
  AND2_X1 U9263 ( .A1(n11705), .A2(n8494), .ZN(n6584) );
  OR2_X1 U9264 ( .A1(n11982), .A2(n13890), .ZN(n6585) );
  AND2_X1 U9265 ( .A1(n6533), .A2(n9474), .ZN(n6586) );
  NOR2_X1 U9266 ( .A1(n14622), .A2(n14151), .ZN(n6587) );
  NOR2_X1 U9267 ( .A1(n15048), .A2(n11125), .ZN(n6588) );
  NOR2_X1 U9268 ( .A1(n12099), .A2(n12098), .ZN(n6589) );
  OR2_X1 U9269 ( .A1(n14502), .A2(n14503), .ZN(n6590) );
  AND2_X1 U9270 ( .A1(n12776), .A2(n12582), .ZN(n6591) );
  AND2_X1 U9271 ( .A1(n12171), .A2(n12353), .ZN(n6592) );
  OR2_X1 U9272 ( .A1(n14356), .A2(n14357), .ZN(n6593) );
  INV_X1 U9273 ( .A(n7390), .ZN(n7389) );
  OAI21_X1 U9274 ( .B1(n7393), .B2(n7391), .A(n13432), .ZN(n7390) );
  AND2_X1 U9275 ( .A1(n10412), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6594) );
  NOR2_X1 U9276 ( .A1(n11868), .A2(n11870), .ZN(n6595) );
  INV_X1 U9277 ( .A(n11831), .ZN(n7636) );
  NAND2_X1 U9278 ( .A1(n7584), .A2(n7582), .ZN(n6596) );
  NAND3_X1 U9279 ( .A1(n7604), .A2(n8579), .A3(n7603), .ZN(n7605) );
  AND2_X1 U9280 ( .A1(n8794), .A2(n9944), .ZN(n6597) );
  INV_X1 U9281 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n9210) );
  AND2_X1 U9282 ( .A1(n6722), .A2(n12986), .ZN(n6598) );
  AND2_X1 U9283 ( .A1(n7103), .A2(n6736), .ZN(n6599) );
  INV_X1 U9284 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9903) );
  AND3_X1 U9285 ( .A1(n9070), .A2(n6920), .A3(n8898), .ZN(n6600) );
  AND2_X1 U9286 ( .A1(n9903), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6601) );
  OR2_X1 U9287 ( .A1(n7407), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n6602) );
  AND2_X1 U9288 ( .A1(n12590), .A2(n8517), .ZN(n8260) );
  NOR2_X1 U9289 ( .A1(n7185), .A2(n13227), .ZN(n6603) );
  OR2_X1 U9290 ( .A1(n8394), .A2(n6753), .ZN(n6604) );
  AND2_X1 U9291 ( .A1(n11775), .A2(n7747), .ZN(n6605) );
  OR2_X1 U9292 ( .A1(n12069), .A2(n12067), .ZN(n6606) );
  OAI21_X1 U9293 ( .B1(n7329), .B2(n7327), .A(n8375), .ZN(n7326) );
  INV_X1 U9294 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6881) );
  INV_X1 U9295 ( .A(n12065), .ZN(n6861) );
  NAND2_X1 U9296 ( .A1(n8837), .A2(n8833), .ZN(n6608) );
  INV_X1 U9297 ( .A(n7359), .ZN(n7358) );
  NAND2_X1 U9298 ( .A1(n13249), .A2(n7362), .ZN(n7359) );
  INV_X1 U9299 ( .A(n7653), .ZN(n7652) );
  NAND2_X1 U9300 ( .A1(n10828), .A2(n10826), .ZN(n7653) );
  INV_X1 U9301 ( .A(n12056), .ZN(n6987) );
  NAND2_X1 U9302 ( .A1(n8268), .A2(n8263), .ZN(n6609) );
  INV_X1 U9303 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7533) );
  OR2_X1 U9304 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n6611) );
  INV_X1 U9305 ( .A(n8374), .ZN(n7331) );
  OR2_X1 U9306 ( .A1(n14480), .A2(n14479), .ZN(n6612) );
  OR2_X1 U9307 ( .A1(n14413), .A2(n14412), .ZN(n6613) );
  OR2_X1 U9308 ( .A1(n10360), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n6614) );
  AND3_X1 U9309 ( .A1(n9195), .A2(n9323), .A3(n9193), .ZN(n6615) );
  OR2_X1 U9310 ( .A1(n9423), .A2(n6565), .ZN(n6616) );
  AND2_X1 U9311 ( .A1(n9594), .A2(n9593), .ZN(n6617) );
  AND2_X1 U9312 ( .A1(n9066), .A2(n7498), .ZN(n6618) );
  NOR2_X1 U9313 ( .A1(n12711), .A2(n7666), .ZN(n7665) );
  INV_X1 U9314 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7268) );
  INV_X1 U9315 ( .A(n7581), .ZN(n7580) );
  AOI21_X1 U9316 ( .B1(n7582), .B2(n8968), .A(n6537), .ZN(n7581) );
  AND2_X1 U9317 ( .A1(n8527), .A2(n12567), .ZN(n6619) );
  AND2_X1 U9318 ( .A1(n13984), .A2(n9037), .ZN(n6620) );
  OR2_X1 U9319 ( .A1(n12054), .A2(n12053), .ZN(n6621) );
  OR2_X1 U9320 ( .A1(n8458), .A2(n8448), .ZN(n6622) );
  AND2_X1 U9321 ( .A1(n14095), .A2(n8923), .ZN(n6623) );
  INV_X1 U9322 ( .A(n11257), .ZN(n7402) );
  AND2_X1 U9323 ( .A1(n7501), .A2(n7508), .ZN(n6624) );
  AND2_X1 U9324 ( .A1(n7661), .A2(n9226), .ZN(n6625) );
  OR2_X1 U9325 ( .A1(n11975), .A2(n11973), .ZN(n6626) );
  OR2_X1 U9326 ( .A1(n6981), .A2(n12003), .ZN(n6627) );
  NOR2_X1 U9327 ( .A1(n7133), .A2(n7132), .ZN(n7131) );
  NAND2_X1 U9328 ( .A1(n6949), .A2(n6950), .ZN(n6628) );
  OR2_X1 U9329 ( .A1(n12118), .A2(n11952), .ZN(n6629) );
  AND2_X1 U9330 ( .A1(n7165), .A2(n7164), .ZN(n6630) );
  INV_X1 U9331 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7800) );
  OR2_X1 U9332 ( .A1(n7718), .A2(n6563), .ZN(n6631) );
  AND2_X1 U9333 ( .A1(n7015), .A2(n7014), .ZN(n6632) );
  AND2_X1 U9334 ( .A1(n7255), .A2(SI_18_), .ZN(n6633) );
  INV_X1 U9335 ( .A(n7099), .ZN(n12603) );
  NAND2_X1 U9336 ( .A1(n7100), .A2(n8268), .ZN(n7099) );
  INV_X1 U9337 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n9236) );
  INV_X1 U9338 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9201) );
  AND2_X1 U9339 ( .A1(n7220), .A2(n7219), .ZN(n6634) );
  INV_X1 U9340 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7786) );
  INV_X1 U9341 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8544) );
  INV_X1 U9342 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8545) );
  INV_X1 U9343 ( .A(n7678), .ZN(n7677) );
  NAND2_X1 U9344 ( .A1(n12595), .A2(n7679), .ZN(n7678) );
  INV_X1 U9345 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7164) );
  OR2_X1 U9346 ( .A1(n13016), .A2(n7650), .ZN(n6635) );
  INV_X1 U9347 ( .A(n10220), .ZN(n13686) );
  INV_X1 U9348 ( .A(n10457), .ZN(n11062) );
  INV_X1 U9349 ( .A(n7854), .ZN(n7536) );
  NAND2_X1 U9350 ( .A1(n9217), .A2(n9223), .ZN(n9495) );
  AND2_X1 U9351 ( .A1(n9627), .A2(n9626), .ZN(n6636) );
  NAND2_X1 U9352 ( .A1(n12230), .A2(n12166), .ZN(n12350) );
  AND2_X1 U9353 ( .A1(n10164), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6637) );
  AND2_X1 U9354 ( .A1(n11033), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6638) );
  XNOR2_X1 U9355 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n7871) );
  INV_X1 U9356 ( .A(n7871), .ZN(n6724) );
  INV_X1 U9357 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7093) );
  INV_X1 U9358 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7095) );
  INV_X1 U9359 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9070) );
  INV_X1 U9360 ( .A(n14211), .ZN(n7230) );
  INV_X1 U9361 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n14359) );
  OR2_X1 U9362 ( .A1(n7984), .A2(n7983), .ZN(n11762) );
  AND2_X1 U9363 ( .A1(n10474), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6639) );
  INV_X1 U9364 ( .A(n15174), .ZN(n11403) );
  NAND2_X1 U9365 ( .A1(n7667), .A2(n7671), .ZN(n12705) );
  AND2_X1 U9366 ( .A1(n9104), .A2(n9103), .ZN(n6640) );
  AND2_X1 U9367 ( .A1(n11810), .A2(n12026), .ZN(n6641) );
  AND2_X1 U9368 ( .A1(n7307), .A2(n7952), .ZN(n6642) );
  NAND2_X1 U9369 ( .A1(n11406), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n6643) );
  NOR2_X1 U9370 ( .A1(n13518), .A2(n13218), .ZN(n6644) );
  AND2_X1 U9371 ( .A1(n7637), .A2(n7642), .ZN(n6645) );
  INV_X1 U9372 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7781) );
  AND2_X1 U9373 ( .A1(n6811), .A2(n8502), .ZN(n6646) );
  INV_X1 U9374 ( .A(n12186), .ZN(n7084) );
  AND2_X1 U9375 ( .A1(n14490), .A2(n12755), .ZN(n6647) );
  INV_X1 U9376 ( .A(n7109), .ZN(n7108) );
  OAI21_X1 U9377 ( .B1(n7994), .B2(n7110), .A(n8005), .ZN(n7109) );
  NAND2_X1 U9378 ( .A1(n8841), .A2(n8842), .ZN(n6648) );
  AND2_X1 U9379 ( .A1(n13673), .A2(n13672), .ZN(n6649) );
  NAND2_X1 U9380 ( .A1(n7667), .A2(n7665), .ZN(n6650) );
  AND2_X1 U9381 ( .A1(n7962), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n6651) );
  INV_X1 U9382 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10102) );
  INV_X1 U9383 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10464) );
  OR2_X1 U9384 ( .A1(n7185), .A2(n12998), .ZN(n6652) );
  NOR2_X1 U9385 ( .A1(n11755), .A2(n11756), .ZN(n6653) );
  AND2_X1 U9386 ( .A1(n11850), .A2(n8809), .ZN(n6654) );
  NAND2_X1 U9387 ( .A1(n7645), .A2(n12959), .ZN(n7649) );
  AND2_X1 U9388 ( .A1(n7287), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n6655) );
  INV_X1 U9389 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7498) );
  NAND2_X1 U9390 ( .A1(n9879), .A2(n15070), .ZN(n14916) );
  INV_X1 U9391 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7005) );
  XNOR2_X1 U9392 ( .A(n9071), .B(n9070), .ZN(n14138) );
  AND2_X1 U9393 ( .A1(n10366), .A2(n12506), .ZN(n12547) );
  NAND2_X1 U9394 ( .A1(n11286), .A2(n6806), .ZN(n11482) );
  NAND2_X1 U9395 ( .A1(n8912), .A2(n8911), .ZN(n14240) );
  INV_X1 U9396 ( .A(n14240), .ZN(n6829) );
  AND2_X1 U9397 ( .A1(n10827), .A2(n7652), .ZN(n6656) );
  NOR2_X1 U9398 ( .A1(n8437), .A2(n8436), .ZN(n8458) );
  INV_X1 U9399 ( .A(n8458), .ZN(n7017) );
  INV_X1 U9400 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7090) );
  NAND2_X1 U9401 ( .A1(n11392), .A2(n11403), .ZN(n11391) );
  NAND2_X1 U9402 ( .A1(n10839), .A2(n8490), .ZN(n11313) );
  INV_X1 U9403 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11441) );
  XOR2_X1 U9404 ( .A(n11511), .B(n11509), .Z(n6657) );
  NAND2_X1 U9405 ( .A1(n8822), .A2(n8821), .ZN(n14622) );
  INV_X1 U9406 ( .A(n9006), .ZN(n7259) );
  AND2_X1 U9407 ( .A1(n7547), .A2(n7545), .ZN(n6658) );
  AND2_X1 U9408 ( .A1(n7427), .A2(n11207), .ZN(n6659) );
  INV_X1 U9409 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10446) );
  AND2_X1 U9410 ( .A1(n7275), .A2(n11391), .ZN(n6660) );
  AND2_X1 U9411 ( .A1(n7284), .A2(n11149), .ZN(n6661) );
  AND2_X1 U9412 ( .A1(n7196), .A2(n11385), .ZN(n6662) );
  AND2_X1 U9413 ( .A1(n7202), .A2(n11748), .ZN(n6663) );
  NOR2_X1 U9414 ( .A1(n7833), .A2(n12897), .ZN(n6664) );
  AND2_X2 U9415 ( .A1(n11191), .A2(n9190), .ZN(n15254) );
  OR2_X1 U9416 ( .A1(n9821), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n6665) );
  AND2_X1 U9417 ( .A1(n9673), .A2(n12893), .ZN(n6666) );
  INV_X1 U9418 ( .A(n7183), .ZN(n14560) );
  AND2_X1 U9419 ( .A1(n12766), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n6667) );
  INV_X1 U9420 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10443) );
  INV_X1 U9421 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11205) );
  INV_X1 U9422 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11021) );
  INV_X1 U9423 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10466) );
  INV_X1 U9424 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10497) );
  AND2_X1 U9425 ( .A1(n11748), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n6668) );
  NOR2_X1 U9426 ( .A1(n11541), .A2(n7767), .ZN(n6669) );
  AND2_X1 U9427 ( .A1(n10871), .A2(n9094), .ZN(n6670) );
  AND2_X1 U9428 ( .A1(n11149), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n6671) );
  INV_X1 U9429 ( .A(n7549), .ZN(n7546) );
  NAND2_X1 U9430 ( .A1(n11717), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7549) );
  INV_X1 U9431 ( .A(n12729), .ZN(n7672) );
  INV_X1 U9432 ( .A(n12369), .ZN(n7085) );
  INV_X1 U9433 ( .A(n13868), .ZN(n14623) );
  AND2_X2 U9434 ( .A1(n10257), .A2(n10852), .ZN(n14891) );
  AND2_X2 U9435 ( .A1(n10621), .A2(n10620), .ZN(n15134) );
  NAND2_X1 U9436 ( .A1(n10640), .A2(n10639), .ZN(n10655) );
  INV_X1 U9437 ( .A(n14499), .ZN(n15206) );
  NAND2_X1 U9438 ( .A1(n8521), .A2(n8520), .ZN(n14499) );
  OR2_X1 U9439 ( .A1(n12164), .A2(n12755), .ZN(n6672) );
  INV_X1 U9440 ( .A(n14835), .ZN(n6828) );
  INV_X1 U9441 ( .A(n11089), .ZN(n7228) );
  NAND2_X1 U9442 ( .A1(n8487), .A2(n8486), .ZN(n10737) );
  AND2_X1 U9443 ( .A1(n7214), .A2(n7216), .ZN(n6673) );
  NOR2_X1 U9444 ( .A1(n14891), .A2(n7589), .ZN(n6674) );
  AND2_X1 U9445 ( .A1(n7209), .A2(n11144), .ZN(n6675) );
  NOR2_X1 U9446 ( .A1(n14896), .A2(n14179), .ZN(n6676) );
  AND2_X1 U9447 ( .A1(n11144), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n6677) );
  OR2_X1 U9448 ( .A1(n13232), .A2(n13231), .ZN(n6678) );
  INV_X1 U9449 ( .A(SI_26_), .ZN(n12897) );
  INV_X1 U9450 ( .A(n12517), .ZN(n12509) );
  AND2_X1 U9451 ( .A1(n10204), .A2(n10203), .ZN(n15127) );
  INV_X1 U9452 ( .A(n15127), .ZN(n14579) );
  OR2_X1 U9453 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n14333), .ZN(n6679) );
  AND2_X1 U9454 ( .A1(n14328), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6680) );
  INV_X1 U9455 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7591) );
  INV_X1 U9456 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n6795) );
  INV_X1 U9457 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7062) );
  INV_X1 U9458 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6883) );
  INV_X1 U9459 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7515) );
  INV_X1 U9460 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7066) );
  NAND3_X1 U9461 ( .A1(n6694), .A2(n6493), .A3(n6555), .ZN(n6695) );
  NAND3_X1 U9462 ( .A1(n11680), .A2(n11673), .A3(n6697), .ZN(n6696) );
  AND3_X2 U9463 ( .A1(n7697), .A2(n6505), .A3(n7762), .ZN(n8051) );
  NAND4_X1 U9464 ( .A1(n7697), .A2(n6505), .A3(n7762), .A4(n15422), .ZN(n8063)
         );
  AOI21_X2 U9465 ( .B1(n6700), .B2(n7350), .A(n7349), .ZN(n13287) );
  NAND2_X1 U9466 ( .A1(n6702), .A2(SI_2_), .ZN(n6892) );
  MUX2_X1 U9467 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n8580), .Z(n6702) );
  NAND2_X4 U9468 ( .A1(n6704), .A2(n6703), .ZN(n8580) );
  NAND2_X2 U9469 ( .A1(n6796), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n6703) );
  NAND2_X1 U9470 ( .A1(n11069), .A2(n11070), .ZN(n11175) );
  XNOR2_X1 U9471 ( .A(n9806), .B(n9248), .ZN(n7625) );
  AND2_X2 U9472 ( .A1(n9229), .A2(n9811), .ZN(n9747) );
  AND2_X2 U9473 ( .A1(n9199), .A2(n9212), .ZN(n9217) );
  AND2_X2 U9474 ( .A1(n9194), .A2(n6615), .ZN(n9212) );
  NAND2_X1 U9475 ( .A1(n7907), .A2(n7906), .ZN(n7909) );
  NAND2_X1 U9476 ( .A1(n8074), .A2(n8075), .ZN(n8076) );
  NAND2_X1 U9477 ( .A1(n6752), .A2(n6751), .ZN(n12564) );
  NAND2_X1 U9478 ( .A1(n6753), .A2(n8260), .ZN(n6751) );
  NAND2_X1 U9479 ( .A1(n14403), .A2(n6758), .ZN(n6756) );
  NAND3_X1 U9480 ( .A1(n6548), .A2(n6510), .A3(n6756), .ZN(n6755) );
  INV_X1 U9481 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6757) );
  OAI21_X1 U9482 ( .B1(n15447), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6613), .ZN(
        n6760) );
  XNOR2_X1 U9483 ( .A(n14413), .B(n14412), .ZN(n15447) );
  AND3_X2 U9484 ( .A1(n7505), .A2(n6624), .A3(n7509), .ZN(n14667) );
  NAND2_X1 U9485 ( .A1(n14446), .A2(n15016), .ZN(n6761) );
  INV_X1 U9486 ( .A(n14666), .ZN(n6762) );
  NOR2_X2 U9487 ( .A1(n14429), .A2(n14650), .ZN(n14654) );
  XNOR2_X1 U9488 ( .A(n14421), .B(n14422), .ZN(n14458) );
  XNOR2_X2 U9489 ( .A(n7033), .B(n6766), .ZN(n10328) );
  NAND2_X1 U9490 ( .A1(n10334), .A2(n6766), .ZN(n10326) );
  OAI21_X1 U9491 ( .B1(n15114), .B2(n6766), .A(n10569), .ZN(n10206) );
  OAI211_X1 U9492 ( .C1(n6766), .C2(n15067), .A(n14562), .B(n10336), .ZN(
        n10569) );
  OAI21_X1 U9493 ( .B1(n15055), .B2(n6766), .A(n6765), .ZN(n10573) );
  INV_X1 U9494 ( .A(n6771), .ZN(n6770) );
  NAND2_X1 U9495 ( .A1(n13362), .A2(n13248), .ZN(n6780) );
  NAND3_X1 U9496 ( .A1(n6789), .A2(n6787), .A3(n14579), .ZN(n6786) );
  NAND2_X1 U9497 ( .A1(n6788), .A2(n13275), .ZN(n6787) );
  INV_X1 U9498 ( .A(n13274), .ZN(n6789) );
  NAND3_X1 U9499 ( .A1(n6795), .A2(P3_ADDR_REG_19__SCAN_IN), .A3(n6794), .ZN(
        n6793) );
  NAND3_X1 U9500 ( .A1(n14475), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(n6797), .ZN(
        n6796) );
  INV_X1 U9501 ( .A(n7681), .ZN(n6799) );
  NAND2_X1 U9502 ( .A1(n12568), .A2(n12567), .ZN(n12566) );
  AOI21_X1 U9503 ( .B1(n12568), .B2(n6619), .A(n6800), .ZN(n6802) );
  INV_X4 U9504 ( .A(n9211), .ZN(n9676) );
  OR2_X1 U9505 ( .A1(n6809), .A2(SI_4_), .ZN(n6808) );
  NAND2_X1 U9506 ( .A1(n9211), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6810) );
  XNOR2_X1 U9507 ( .A(n13205), .B(n13201), .ZN(n13195) );
  NOR2_X2 U9508 ( .A1(n13263), .A2(n13204), .ZN(n13205) );
  NAND2_X1 U9509 ( .A1(n8501), .A2(n7689), .ZN(n6811) );
  NAND3_X1 U9510 ( .A1(n7697), .A2(n7762), .A3(n6495), .ZN(n8040) );
  INV_X2 U9511 ( .A(n7892), .ZN(n7697) );
  NOR2_X2 U9512 ( .A1(n13373), .A2(n13501), .ZN(n13357) );
  NOR2_X1 U9513 ( .A1(n11726), .A2(n14573), .ZN(n7183) );
  INV_X1 U9514 ( .A(n6820), .ZN(n14561) );
  XNOR2_X2 U9515 ( .A(n6821), .B(n7800), .ZN(n8450) );
  INV_X1 U9516 ( .A(n6824), .ZN(n14172) );
  NAND3_X1 U9517 ( .A1(n11472), .A2(n6825), .A3(n7233), .ZN(n14148) );
  NOR2_X2 U9518 ( .A1(n13941), .A2(n13942), .ZN(n13940) );
  AND2_X1 U9519 ( .A1(n10857), .A2(n10928), .ZN(n10931) );
  NOR2_X2 U9520 ( .A1(n14076), .A2(n14089), .ZN(n14060) );
  OAI211_X1 U9521 ( .C1(n6832), .C2(n14787), .A(n11558), .B(n14837), .ZN(
        n11373) );
  NAND4_X1 U9522 ( .A1(n7563), .A2(n8841), .A3(n8541), .A4(n8542), .ZN(n6833)
         );
  NAND2_X2 U9523 ( .A1(n14334), .A2(n14331), .ZN(n8947) );
  NAND3_X1 U9524 ( .A1(n6835), .A2(n11951), .A3(n6629), .ZN(n11957) );
  NAND2_X1 U9525 ( .A1(n11953), .A2(n11949), .ZN(n6835) );
  MUX2_X1 U9526 ( .A(n7060), .B(n13897), .S(n12002), .Z(n11953) );
  NAND2_X1 U9527 ( .A1(n6838), .A2(n6836), .ZN(n12149) );
  NAND2_X1 U9528 ( .A1(n6982), .A2(n6840), .ZN(n6839) );
  NAND4_X1 U9529 ( .A1(n6842), .A2(n7484), .A3(n6841), .A4(n6839), .ZN(n7019)
         );
  NAND2_X1 U9530 ( .A1(n6982), .A2(n6843), .ZN(n6842) );
  INV_X1 U9531 ( .A(n6980), .ZN(n6844) );
  OAI211_X1 U9532 ( .C1(n6854), .C2(n6632), .A(n6853), .B(n7479), .ZN(n11985)
         );
  NAND3_X1 U9533 ( .A1(n12064), .A2(n12063), .A3(n6860), .ZN(n6859) );
  NAND3_X1 U9534 ( .A1(n7468), .A2(n6621), .A3(n6863), .ZN(n6862) );
  XNOR2_X2 U9535 ( .A(n12501), .B(n12517), .ZN(n12481) );
  NAND3_X1 U9536 ( .A1(n7285), .A2(n6655), .A3(n11149), .ZN(n6868) );
  NAND3_X1 U9537 ( .A1(n6496), .A2(n7523), .A3(n6614), .ZN(n6872) );
  INV_X1 U9538 ( .A(n10531), .ZN(n6871) );
  OR2_X2 U9539 ( .A1(n12406), .A2(n6873), .ZN(n12383) );
  OAI21_X1 U9540 ( .B1(n9021), .B2(n6875), .A(n6874), .ZN(n9065) );
  INV_X1 U9541 ( .A(n6876), .ZN(n6875) );
  NAND2_X1 U9542 ( .A1(n6877), .A2(n7465), .ZN(P1_U3557) );
  NAND2_X1 U9543 ( .A1(n14178), .A2(n14896), .ZN(n6877) );
  NAND2_X1 U9544 ( .A1(n13947), .A2(n14887), .ZN(n6878) );
  NAND2_X2 U9545 ( .A1(n8955), .A2(n8954), .ZN(n14043) );
  NAND2_X2 U9546 ( .A1(n6884), .A2(n6573), .ZN(n14095) );
  NAND2_X1 U9547 ( .A1(n6885), .A2(n8682), .ZN(n6887) );
  NAND2_X1 U9548 ( .A1(n8684), .A2(n6888), .ZN(n9935) );
  NAND3_X1 U9549 ( .A1(n7236), .A2(n6889), .A3(n7235), .ZN(n6888) );
  NAND2_X1 U9550 ( .A1(n8599), .A2(n6892), .ZN(n8600) );
  OAI21_X2 U9551 ( .B1(n8671), .B2(n6896), .A(n6894), .ZN(n8701) );
  OAI21_X1 U9552 ( .B1(n7743), .B2(n6927), .A(n13625), .ZN(n6922) );
  NAND2_X1 U9553 ( .A1(n6923), .A2(n6921), .ZN(n14611) );
  INV_X1 U9554 ( .A(n6922), .ZN(n6921) );
  NAND2_X1 U9555 ( .A1(n6928), .A2(n7743), .ZN(n11782) );
  NAND2_X1 U9556 ( .A1(n11532), .A2(n7744), .ZN(n6928) );
  NAND3_X1 U9557 ( .A1(n8551), .A2(n8550), .A3(P1_REG3_REG_1__SCAN_IN), .ZN(
        n8567) );
  XNOR2_X2 U9558 ( .A(n8546), .B(P1_IR_REG_30__SCAN_IN), .ZN(n8550) );
  NAND2_X1 U9559 ( .A1(n13852), .A2(n6932), .ZN(n6931) );
  NAND2_X2 U9560 ( .A1(n6931), .A2(n6557), .ZN(n13821) );
  INV_X1 U9561 ( .A(n7725), .ZN(n6938) );
  NAND3_X1 U9562 ( .A1(n6939), .A2(n6937), .A3(n13769), .ZN(P1_U3220) );
  NAND2_X1 U9563 ( .A1(n6940), .A2(n6938), .ZN(n6937) );
  NAND3_X1 U9564 ( .A1(n6513), .A2(n7725), .A3(n14623), .ZN(n6939) );
  NAND2_X1 U9565 ( .A1(n7725), .A2(n7724), .ZN(n13758) );
  INV_X1 U9566 ( .A(n13763), .ZN(n6950) );
  NAND2_X1 U9567 ( .A1(n13770), .A2(n6954), .ZN(n6951) );
  NAND2_X1 U9568 ( .A1(n6951), .A2(n6952), .ZN(n13706) );
  NOR2_X2 U9569 ( .A1(n13832), .A2(n7734), .ZN(n14595) );
  AND2_X2 U9570 ( .A1(n6974), .A2(n6973), .ZN(n13832) );
  NAND2_X1 U9571 ( .A1(n9133), .A2(n6959), .ZN(n8560) );
  NAND2_X1 U9572 ( .A1(n9133), .A2(n6958), .ZN(n14320) );
  NAND2_X2 U9573 ( .A1(n7735), .A2(n7738), .ZN(n13852) );
  NOR2_X1 U9574 ( .A1(n10807), .A2(n10806), .ZN(n10890) );
  AOI21_X1 U9575 ( .B1(n11045), .B2(n11044), .A(n6991), .ZN(n11113) );
  NAND2_X1 U9576 ( .A1(n10342), .A2(n10220), .ZN(n10190) );
  NAND2_X1 U9577 ( .A1(n10227), .A2(n10226), .ZN(n10272) );
  NAND2_X1 U9578 ( .A1(n11118), .A2(n11117), .ZN(n11529) );
  AOI21_X1 U9579 ( .B1(n10892), .B2(n10891), .A(n10890), .ZN(n11045) );
  NAND2_X1 U9580 ( .A1(n14000), .A2(n13999), .ZN(n13998) );
  NAND2_X1 U9581 ( .A1(n9092), .A2(n9091), .ZN(n10870) );
  NAND2_X1 U9582 ( .A1(n14611), .A2(n6990), .ZN(n13787) );
  NAND2_X1 U9583 ( .A1(n14046), .A2(n14045), .ZN(n14044) );
  OAI21_X1 U9584 ( .B1(n10930), .B2(n9084), .A(n9085), .ZN(n10907) );
  OAI21_X1 U9585 ( .B1(n13687), .B2(n14861), .A(n10265), .ZN(n10266) );
  NAND2_X1 U9586 ( .A1(n12077), .A2(n12076), .ZN(n12080) );
  AOI21_X1 U9587 ( .B1(n6988), .B2(n7488), .A(n7483), .ZN(n7482) );
  NAND2_X1 U9588 ( .A1(n8600), .A2(n6559), .ZN(n8620) );
  OAI21_X1 U9589 ( .B1(n14481), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n6612), .ZN(
        n7036) );
  NAND2_X1 U9590 ( .A1(n6966), .A2(n14499), .ZN(n7687) );
  XNOR2_X1 U9591 ( .A(n9168), .B(n9167), .ZN(n6966) );
  NAND2_X1 U9592 ( .A1(n11894), .A2(n11895), .ZN(n8501) );
  INV_X1 U9593 ( .A(n7338), .ZN(n7333) );
  NAND2_X1 U9594 ( .A1(n7674), .A2(n7673), .ZN(n11241) );
  NAND2_X1 U9595 ( .A1(n11482), .A2(n6584), .ZN(n11704) );
  OAI21_X1 U9596 ( .B1(n7686), .B2(n15244), .A(n7294), .ZN(P3_U3456) );
  AOI21_X1 U9597 ( .B1(n7663), .B2(n7665), .A(n7662), .ZN(n12690) );
  INV_X1 U9598 ( .A(n7332), .ZN(n12565) );
  OAI21_X1 U9599 ( .B1(n12768), .B2(n12586), .A(n12571), .ZN(n6993) );
  NOR2_X2 U9600 ( .A1(n7511), .A2(n14423), .ZN(n14460) );
  NAND2_X1 U9601 ( .A1(n8574), .A2(n11954), .ZN(n14824) );
  OAI21_X2 U9602 ( .B1(n14113), .B2(n8887), .A(n8886), .ZN(n14101) );
  NAND2_X1 U9603 ( .A1(n12117), .A2(n10339), .ZN(n8574) );
  INV_X2 U9604 ( .A(n13895), .ZN(n10267) );
  NAND2_X1 U9605 ( .A1(n8609), .A2(n7573), .ZN(n7572) );
  NAND2_X1 U9606 ( .A1(n11470), .A2(n8791), .ZN(n11852) );
  NAND2_X1 U9607 ( .A1(n11447), .A2(n8771), .ZN(n11471) );
  NAND2_X1 U9608 ( .A1(n11370), .A2(n8737), .ZN(n11555) );
  NAND2_X1 U9609 ( .A1(n7565), .A2(n6507), .ZN(n11420) );
  INV_X1 U9610 ( .A(n8874), .ZN(n7035) );
  NAND2_X1 U9611 ( .A1(n8857), .A2(n8856), .ZN(n8860) );
  NAND2_X1 U9612 ( .A1(n8620), .A2(n8619), .ZN(n8621) );
  NAND3_X1 U9613 ( .A1(n7131), .A2(n7124), .A3(n6972), .ZN(n7127) );
  NAND2_X1 U9614 ( .A1(n8840), .A2(n8839), .ZN(n8857) );
  AOI21_X1 U9615 ( .B1(n7028), .B2(n14579), .A(n6520), .ZN(n13271) );
  INV_X1 U9616 ( .A(n7401), .ZN(n7400) );
  AOI21_X1 U9617 ( .B1(n13383), .B2(n13382), .A(n13222), .ZN(n13366) );
  INV_X4 U9618 ( .A(n8580), .ZN(n9211) );
  OAI22_X1 U9619 ( .A1(n14552), .A2(n11882), .B1(n11881), .B2(n14559), .ZN(
        n11883) );
  OAI21_X1 U9620 ( .B1(n7405), .B2(n7404), .A(n10760), .ZN(n10995) );
  INV_X1 U9621 ( .A(n12185), .ZN(n7069) );
  NOR2_X1 U9622 ( .A1(n11684), .A2(n11683), .ZN(n11685) );
  OAI21_X1 U9623 ( .B1(n9089), .B2(n11091), .A(n7448), .ZN(n10945) );
  INV_X1 U9624 ( .A(n11970), .ZN(n7021) );
  NAND3_X1 U9625 ( .A1(n12000), .A2(n12001), .A3(n6627), .ZN(n6982) );
  NAND2_X1 U9626 ( .A1(n13217), .A2(n13216), .ZN(n13395) );
  NAND4_X1 U9627 ( .A1(n10361), .A2(n7772), .A3(n7771), .A4(n7773), .ZN(n7892)
         );
  NAND2_X1 U9628 ( .A1(n14181), .A2(n14269), .ZN(n14186) );
  NAND2_X1 U9629 ( .A1(n11241), .A2(n8492), .ZN(n11287) );
  NAND2_X1 U9630 ( .A1(n11704), .A2(n8495), .ZN(n11800) );
  OR2_X1 U9631 ( .A1(n14288), .A2(n9119), .ZN(n6985) );
  NAND2_X1 U9632 ( .A1(n8533), .A2(n12563), .ZN(n12765) );
  AOI21_X1 U9633 ( .B1(n12639), .B2(n8514), .A(n7755), .ZN(n12625) );
  NAND2_X1 U9634 ( .A1(n10839), .A2(n7675), .ZN(n7674) );
  NAND2_X1 U9635 ( .A1(n8705), .A2(n7595), .ZN(n7594) );
  NAND2_X1 U9636 ( .A1(n8761), .A2(n7242), .ZN(n7241) );
  NAND2_X1 U9637 ( .A1(n7241), .A2(n7240), .ZN(n8840) );
  NAND2_X1 U9638 ( .A1(n7486), .A2(n7489), .ZN(n6988) );
  NAND2_X1 U9639 ( .A1(n8568), .A2(n9892), .ZN(n7604) );
  OAI21_X2 U9640 ( .B1(n11255), .B2(n7368), .A(n7366), .ZN(n11719) );
  OAI211_X1 U9641 ( .C1(n8580), .C2(P2_DATAO_REG_0__SCAN_IN), .A(n6989), .B(
        SI_0_), .ZN(n8570) );
  INV_X1 U9642 ( .A(n11254), .ZN(n7369) );
  NAND2_X1 U9643 ( .A1(n13706), .A2(n13705), .ZN(n13793) );
  NAND2_X1 U9644 ( .A1(n10183), .A2(n7060), .ZN(n10218) );
  NAND4_X1 U9645 ( .A1(n6600), .A2(n8536), .A3(n8537), .A4(n8535), .ZN(n8538)
         );
  AND2_X1 U9646 ( .A1(n10187), .A2(n10186), .ZN(n10221) );
  NAND4_X1 U9647 ( .A1(n8595), .A2(n8596), .A3(n8597), .A4(n8598), .ZN(n13894)
         );
  OAI22_X1 U9648 ( .A1(n13615), .A2(n10341), .B1(n14844), .B2(n13686), .ZN(
        n10268) );
  NOR2_X2 U9649 ( .A1(n8877), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n8899) );
  NAND4_X1 U9650 ( .A1(n7496), .A2(n6491), .A3(n6506), .A4(n7756), .ZN(n8877)
         );
  NAND3_X1 U9651 ( .A1(n12947), .A2(n12946), .A3(n6652), .ZN(P2_U3186) );
  NAND2_X1 U9652 ( .A1(n10452), .A2(n10456), .ZN(n10827) );
  NAND2_X1 U9653 ( .A1(n6996), .A2(n6994), .ZN(P3_U3454) );
  OR2_X1 U9654 ( .A1(n12830), .A2(n15244), .ZN(n6996) );
  NAND3_X1 U9655 ( .A1(n7252), .A2(n7251), .A3(n7249), .ZN(n8891) );
  NAND2_X1 U9656 ( .A1(n13552), .A2(n15145), .ZN(n7353) );
  NAND2_X1 U9657 ( .A1(n10751), .A2(n10750), .ZN(n10991) );
  AND2_X1 U9658 ( .A1(n15149), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15153) );
  NOR2_X1 U9659 ( .A1(n11766), .A2(n11765), .ZN(n12389) );
  AOI21_X1 U9660 ( .B1(n12415), .B2(n12414), .A(n12413), .ZN(n12416) );
  NAND3_X1 U9661 ( .A1(n6634), .A2(n7000), .A3(n6999), .ZN(P3_U3201) );
  OR2_X2 U9662 ( .A1(n12548), .A2(n15162), .ZN(n7000) );
  NAND2_X1 U9663 ( .A1(n13273), .A2(n13275), .ZN(n13272) );
  NAND2_X1 U9664 ( .A1(n7348), .A2(n6570), .ZN(n10751) );
  NAND2_X1 U9665 ( .A1(n11852), .A2(n6490), .ZN(n7051) );
  NOR2_X1 U9666 ( .A1(n7338), .A2(n8394), .ZN(n7336) );
  AOI21_X1 U9667 ( .B1(n7684), .B2(n7687), .A(n7683), .ZN(P3_U3488) );
  NAND2_X1 U9668 ( .A1(n7007), .A2(n7717), .ZN(n9406) );
  NAND3_X1 U9669 ( .A1(n9378), .A2(n6631), .A3(n9377), .ZN(n7007) );
  INV_X1 U9670 ( .A(n13320), .ZN(n7027) );
  NAND2_X1 U9671 ( .A1(n9527), .A2(n9528), .ZN(n9526) );
  OAI21_X1 U9672 ( .B1(n9438), .B2(n9437), .A(n7008), .ZN(n7711) );
  NAND2_X1 U9673 ( .A1(n7010), .A2(n7009), .ZN(n7008) );
  NAND2_X1 U9674 ( .A1(n9438), .A2(n9437), .ZN(n7010) );
  INV_X1 U9675 ( .A(n9355), .ZN(n7137) );
  NAND2_X1 U9676 ( .A1(n7158), .A2(n7157), .ZN(n9580) );
  NAND2_X1 U9677 ( .A1(n7012), .A2(n7011), .ZN(n9291) );
  INV_X1 U9678 ( .A(n9906), .ZN(n7012) );
  NAND2_X1 U9679 ( .A1(n8599), .A2(n8583), .ZN(n9906) );
  AOI21_X1 U9680 ( .B1(n9491), .B2(n9490), .A(n9489), .ZN(n9493) );
  OAI211_X1 U9681 ( .C1(n9342), .C2(n7139), .A(n7135), .B(n7138), .ZN(n7136)
         );
  NOR2_X1 U9682 ( .A1(n9581), .A2(n7144), .ZN(n7143) );
  OR3_X1 U9683 ( .A1(n9618), .A2(n9617), .A3(n7706), .ZN(n7705) );
  NAND2_X1 U9684 ( .A1(n7705), .A2(n7704), .ZN(n9670) );
  NAND2_X1 U9685 ( .A1(n7013), .A2(n11960), .ZN(n11962) );
  NAND2_X1 U9686 ( .A1(n11957), .A2(n11956), .ZN(n7013) );
  NAND3_X1 U9687 ( .A1(n11972), .A2(n11971), .A3(n6626), .ZN(n7015) );
  AOI21_X1 U9688 ( .B1(n7645), .B2(n12960), .A(n6635), .ZN(n7644) );
  NAND2_X1 U9689 ( .A1(n12949), .A2(n12922), .ZN(n12948) );
  NAND2_X1 U9690 ( .A1(n7423), .A2(n7422), .ZN(n11684) );
  NAND2_X1 U9691 ( .A1(n7035), .A2(n6633), .ZN(n7252) );
  NAND2_X1 U9692 ( .A1(n9778), .A2(n9772), .ZN(n7133) );
  XNOR2_X1 U9693 ( .A(n9672), .B(n9671), .ZN(n13575) );
  OAI21_X1 U9694 ( .B1(n9817), .B2(n9816), .A(n9815), .ZN(n9830) );
  NAND2_X1 U9695 ( .A1(n8896), .A2(n8895), .ZN(n8910) );
  NAND4_X2 U9696 ( .A1(n8552), .A2(n8554), .A3(n8553), .A4(n8555), .ZN(n10342)
         );
  INV_X1 U9697 ( .A(n9773), .ZN(n7132) );
  NAND2_X1 U9698 ( .A1(n8971), .A2(n8970), .ZN(n8974) );
  OAI21_X2 U9699 ( .B1(n8945), .B2(n8944), .A(n8943), .ZN(n8956) );
  NAND2_X1 U9700 ( .A1(n7019), .A2(n7482), .ZN(n7022) );
  OR2_X1 U9701 ( .A1(n11998), .A2(n11999), .ZN(n12000) );
  NAND2_X1 U9702 ( .A1(n13739), .A2(n10805), .ZN(n10807) );
  XNOR2_X1 U9703 ( .A(n14352), .B(n14353), .ZN(n14408) );
  NAND2_X1 U9704 ( .A1(n10219), .A2(n10218), .ZN(n7023) );
  INV_X1 U9705 ( .A(n8560), .ZN(n8547) );
  NAND2_X1 U9706 ( .A1(n11449), .A2(n11448), .ZN(n11447) );
  XNOR2_X1 U9707 ( .A(n13228), .B(n7029), .ZN(n7028) );
  INV_X1 U9708 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13587) );
  NAND2_X1 U9709 ( .A1(n8093), .A2(n8094), .ZN(n7091) );
  NAND3_X1 U9710 ( .A1(n8427), .A2(n7538), .A3(n7539), .ZN(n7026) );
  NOR2_X1 U9711 ( .A1(n10645), .A2(n7406), .ZN(n7404) );
  XNOR2_X1 U9712 ( .A(n9679), .B(n9678), .ZN(n11938) );
  XNOR2_X1 U9713 ( .A(n14480), .B(n14479), .ZN(n14481) );
  XNOR2_X1 U9714 ( .A(n7036), .B(n14482), .ZN(SUB_1596_U4) );
  AOI21_X1 U9715 ( .B1(n15031), .B2(n14448), .A(n14467), .ZN(n14480) );
  NOR2_X1 U9716 ( .A1(n14408), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n14354) );
  NAND2_X1 U9717 ( .A1(n13897), .A2(n10220), .ZN(n10219) );
  NAND2_X1 U9718 ( .A1(n7043), .A2(n7040), .ZN(P1_U3559) );
  OR2_X1 U9719 ( .A1(n14280), .A2(n14894), .ZN(n7043) );
  INV_X1 U9720 ( .A(n7232), .ZN(n14147) );
  XNOR2_X1 U9721 ( .A(n7273), .B(n7272), .ZN(n12548) );
  NAND2_X1 U9722 ( .A1(n10414), .A2(n10413), .ZN(n7045) );
  NAND2_X1 U9723 ( .A1(n7522), .A2(n7809), .ZN(n7521) );
  NAND2_X1 U9724 ( .A1(n10221), .A2(n10222), .ZN(n10225) );
  INV_X1 U9725 ( .A(n7367), .ZN(n7366) );
  OAI21_X1 U9726 ( .B1(n6545), .B2(n7368), .A(n11610), .ZN(n7367) );
  NAND2_X1 U9727 ( .A1(n13552), .A2(n15134), .ZN(n7263) );
  XNOR2_X2 U9728 ( .A(n13917), .B(n13916), .ZN(n14727) );
  XNOR2_X2 U9729 ( .A(n13926), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n13927) );
  NAND2_X1 U9730 ( .A1(n8722), .A2(n8721), .ZN(n8726) );
  AOI21_X2 U9731 ( .B1(n14699), .B2(P1_REG1_REG_13__SCAN_IN), .A(n14691), .ZN(
        n14710) );
  OAI21_X1 U9732 ( .B1(n13928), .B2(n14767), .A(n7173), .ZN(n7172) );
  OAI21_X1 U9733 ( .B1(n13931), .B2(n13930), .A(n7170), .ZN(P1_U3262) );
  NAND4_X2 U9734 ( .A1(n8563), .A2(n8566), .A3(n8567), .A4(n8564), .ZN(n13897)
         );
  NAND2_X1 U9735 ( .A1(n7644), .A2(n7649), .ZN(n7648) );
  NAND2_X1 U9736 ( .A1(n14457), .A2(n14456), .ZN(n7514) );
  OAI21_X1 U9737 ( .B1(n10803), .B2(n10802), .A(n10805), .ZN(n13737) );
  INV_X1 U9738 ( .A(n12030), .ZN(n7489) );
  NAND2_X1 U9739 ( .A1(n7470), .A2(n12156), .ZN(P1_U3242) );
  NAND3_X1 U9740 ( .A1(n8646), .A2(n7570), .A3(n7572), .ZN(n10904) );
  NAND2_X1 U9741 ( .A1(n7513), .A2(n15387), .ZN(n7512) );
  INV_X2 U9742 ( .A(n7060), .ZN(n14844) );
  OAI21_X1 U9743 ( .B1(n7471), .B2(n12150), .A(n9949), .ZN(n7470) );
  NAND2_X1 U9744 ( .A1(n10272), .A2(n10271), .ZN(n10273) );
  NAND2_X1 U9745 ( .A1(n11375), .A2(n12127), .ZN(n11374) );
  AND2_X4 U9746 ( .A1(n11942), .A2(n12100), .ZN(n14837) );
  NAND2_X1 U9747 ( .A1(n9067), .A2(n9066), .ZN(n9069) );
  NAND2_X1 U9748 ( .A1(n14595), .A2(n14596), .ZN(n14594) );
  XNOR2_X1 U9749 ( .A(n10997), .B(n13086), .ZN(n10994) );
  NAND2_X1 U9750 ( .A1(n7353), .A2(n7351), .ZN(P2_U3528) );
  NAND2_X1 U9751 ( .A1(n11614), .A2(n11613), .ZN(n11615) );
  INV_X1 U9752 ( .A(n8570), .ZN(n7603) );
  OAI21_X2 U9753 ( .B1(n8580), .B2(n9929), .A(n7065), .ZN(n8569) );
  NAND2_X1 U9754 ( .A1(n7263), .A2(n7262), .ZN(P2_U3496) );
  NAND2_X1 U9755 ( .A1(n14459), .A2(n7068), .ZN(n14464) );
  NAND2_X2 U9756 ( .A1(n13821), .A2(n6574), .ZN(n13770) );
  NAND2_X1 U9757 ( .A1(n8543), .A2(n6503), .ZN(n7753) );
  NAND3_X1 U9758 ( .A1(n10797), .A2(n10804), .A3(n10796), .ZN(n13739) );
  NAND2_X1 U9759 ( .A1(n15446), .A2(n15445), .ZN(n7067) );
  NAND2_X1 U9760 ( .A1(n14654), .A2(n14653), .ZN(n7513) );
  NAND2_X1 U9761 ( .A1(n12174), .A2(n7075), .ZN(n7071) );
  INV_X1 U9762 ( .A(n12317), .ZN(n7079) );
  NAND4_X1 U9763 ( .A1(n7080), .A2(n12642), .A3(n6504), .A4(n7082), .ZN(n12237) );
  NAND2_X1 U9764 ( .A1(n7083), .A2(n12317), .ZN(n7082) );
  NAND2_X1 U9765 ( .A1(n7079), .A2(n12186), .ZN(n7080) );
  NAND3_X1 U9766 ( .A1(n7082), .A2(n6504), .A3(n7080), .ZN(n12238) );
  NAND2_X1 U9767 ( .A1(n12237), .A2(n12288), .ZN(n12191) );
  NAND2_X1 U9768 ( .A1(n7088), .A2(n7822), .ZN(n7835) );
  INV_X1 U9769 ( .A(n7100), .ZN(n12607) );
  OAI211_X1 U9770 ( .C1(n7120), .C2(n9406), .A(n6616), .B(n7119), .ZN(n7118)
         );
  NAND2_X1 U9771 ( .A1(n7118), .A2(n7719), .ZN(n9438) );
  NAND2_X1 U9772 ( .A1(n6534), .A2(n7121), .ZN(n7119) );
  INV_X1 U9773 ( .A(n9405), .ZN(n7121) );
  AOI21_X1 U9774 ( .B1(n9735), .B2(n7125), .A(n7128), .ZN(n7123) );
  NAND2_X1 U9775 ( .A1(n9736), .A2(n7134), .ZN(n7124) );
  NAND2_X1 U9776 ( .A1(n7123), .A2(n7122), .ZN(n7703) );
  NAND2_X1 U9777 ( .A1(n7137), .A2(n9356), .ZN(n7135) );
  NAND2_X1 U9778 ( .A1(n6544), .A2(n7140), .ZN(n7138) );
  NAND3_X1 U9779 ( .A1(n7145), .A2(n7142), .A3(n7141), .ZN(n9616) );
  NAND2_X1 U9780 ( .A1(n6617), .A2(n9596), .ZN(n7141) );
  NAND2_X1 U9781 ( .A1(n7146), .A2(n7143), .ZN(n7142) );
  INV_X1 U9782 ( .A(n9596), .ZN(n7144) );
  NAND3_X1 U9783 ( .A1(n7146), .A2(n7147), .A3(n6617), .ZN(n7145) );
  NAND2_X1 U9784 ( .A1(n9472), .A2(n6500), .ZN(n7148) );
  NAND2_X1 U9785 ( .A1(n7148), .A2(n7149), .ZN(n9491) );
  INV_X1 U9786 ( .A(n9471), .ZN(n7152) );
  NAND3_X1 U9787 ( .A1(n7154), .A2(n7153), .A3(n9563), .ZN(n7157) );
  NAND2_X1 U9788 ( .A1(n9548), .A2(n9564), .ZN(n7153) );
  NAND2_X1 U9789 ( .A1(n9549), .A2(n9564), .ZN(n7154) );
  NAND3_X1 U9790 ( .A1(n7156), .A2(n7155), .A3(n9565), .ZN(n7158) );
  OAI22_X2 U9791 ( .A1(n7162), .A2(n7159), .B1(n9510), .B2(n9509), .ZN(n9527)
         );
  INV_X1 U9792 ( .A(n9510), .ZN(n7160) );
  INV_X1 U9793 ( .A(n9509), .ZN(n7161) );
  NAND2_X1 U9794 ( .A1(n9217), .A2(n6630), .ZN(n7163) );
  NOR2_X2 U9795 ( .A1(n14705), .A2(n7168), .ZN(n13902) );
  NOR2_X2 U9796 ( .A1(n14694), .A2(n7169), .ZN(n14703) );
  NAND2_X1 U9797 ( .A1(n13452), .A2(n7175), .ZN(n13551) );
  NOR2_X1 U9798 ( .A1(n13205), .A2(n13459), .ZN(n7177) );
  NOR2_X2 U9799 ( .A1(n11924), .A2(n13538), .ZN(n13437) );
  NAND2_X1 U9800 ( .A1(n7194), .A2(n10368), .ZN(n10369) );
  NOR2_X2 U9801 ( .A1(n7837), .A2(n7266), .ZN(n10406) );
  NAND3_X1 U9802 ( .A1(n7839), .A2(n7192), .A3(P3_REG1_REG_2__SCAN_IN), .ZN(
        n7191) );
  NAND2_X1 U9803 ( .A1(n11387), .A2(n7199), .ZN(n7195) );
  NAND2_X1 U9804 ( .A1(n7197), .A2(n7195), .ZN(n11573) );
  NAND3_X1 U9805 ( .A1(n7198), .A2(n11385), .A3(n6518), .ZN(n7197) );
  NAND2_X1 U9806 ( .A1(n11750), .A2(n7206), .ZN(n7201) );
  NAND2_X1 U9807 ( .A1(n7201), .A2(n7203), .ZN(n12379) );
  NAND3_X1 U9808 ( .A1(n7205), .A2(n11748), .A3(n7204), .ZN(n7203) );
  INV_X1 U9809 ( .A(n11574), .ZN(n7207) );
  NAND2_X1 U9810 ( .A1(n7205), .A2(n11748), .ZN(n11575) );
  NAND2_X1 U9811 ( .A1(n7207), .A2(n11585), .ZN(n7205) );
  NAND2_X1 U9812 ( .A1(n11146), .A2(n7213), .ZN(n7208) );
  NAND2_X1 U9813 ( .A1(n7208), .A2(n7210), .ZN(n11384) );
  NAND3_X1 U9814 ( .A1(n7211), .A2(n11144), .A3(n6512), .ZN(n7210) );
  NAND2_X1 U9815 ( .A1(n7211), .A2(n11144), .ZN(n10771) );
  NAND2_X1 U9816 ( .A1(n7212), .A2(n10772), .ZN(n7211) );
  INV_X1 U9817 ( .A(n10770), .ZN(n7212) );
  INV_X1 U9818 ( .A(n10602), .ZN(n7214) );
  OR2_X1 U9819 ( .A1(n7217), .A2(n7218), .ZN(n7216) );
  INV_X1 U9820 ( .A(n10404), .ZN(n7217) );
  INV_X1 U9821 ( .A(n10413), .ZN(n7218) );
  OAI21_X1 U9822 ( .B1(n8635), .B2(n7239), .A(n7237), .ZN(n8667) );
  NAND2_X1 U9823 ( .A1(n8874), .A2(n6528), .ZN(n7251) );
  NAND3_X1 U9824 ( .A1(n7252), .A2(n7253), .A3(n7251), .ZN(n8889) );
  NAND2_X1 U9825 ( .A1(n8987), .A2(n8986), .ZN(n7256) );
  OAI21_X1 U9826 ( .B1(n8987), .B2(n7258), .A(n7257), .ZN(n9023) );
  AOI21_X1 U9827 ( .B1(n8989), .B2(n7260), .A(n7259), .ZN(n7257) );
  NAND2_X1 U9828 ( .A1(n8989), .A2(n7261), .ZN(n7258) );
  NAND2_X1 U9829 ( .A1(n11393), .A2(n7278), .ZN(n7274) );
  NAND2_X1 U9830 ( .A1(n7276), .A2(n7274), .ZN(n11577) );
  NAND3_X1 U9831 ( .A1(n7277), .A2(n11391), .A3(n6519), .ZN(n7276) );
  AND2_X2 U9832 ( .A1(n7281), .A2(n7280), .ZN(n12501) );
  NAND2_X1 U9833 ( .A1(n7285), .A2(n11149), .ZN(n10784) );
  NAND2_X1 U9834 ( .A1(n7286), .A2(n10772), .ZN(n7285) );
  INV_X1 U9835 ( .A(n10783), .ZN(n7286) );
  NAND2_X1 U9836 ( .A1(n11240), .A2(n11239), .ZN(n11238) );
  NAND2_X1 U9837 ( .A1(n11309), .A2(n11314), .ZN(n7293) );
  NAND2_X1 U9838 ( .A1(n12744), .A2(n7299), .ZN(n7296) );
  NAND2_X1 U9839 ( .A1(n7296), .A2(n7297), .ZN(n12714) );
  OAI21_X1 U9840 ( .B1(n11703), .B2(n7304), .A(n7302), .ZN(n14505) );
  INV_X1 U9841 ( .A(n12671), .ZN(n7323) );
  NAND2_X1 U9842 ( .A1(n7317), .A2(n12671), .ZN(n7316) );
  AOI21_X1 U9843 ( .B1(n12603), .B2(n7340), .A(n7333), .ZN(n7332) );
  NAND2_X1 U9844 ( .A1(n8051), .A2(n7345), .ZN(n7801) );
  NAND2_X1 U9845 ( .A1(n10655), .A2(n10654), .ZN(n7348) );
  INV_X1 U9846 ( .A(n13353), .ZN(n7363) );
  AND2_X1 U9847 ( .A1(n13501), .A2(n13248), .ZN(n7364) );
  INV_X1 U9848 ( .A(n7372), .ZN(n9209) );
  NAND4_X1 U9849 ( .A1(n9199), .A2(n9212), .A3(n9204), .A4(n7370), .ZN(n7372)
         );
  NAND2_X1 U9850 ( .A1(n7372), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7371) );
  INV_X1 U9851 ( .A(n7374), .ZN(n7385) );
  OAI21_X1 U9852 ( .B1(n11934), .B2(n7391), .A(n7389), .ZN(n13431) );
  INV_X1 U9853 ( .A(n13211), .ZN(n7395) );
  NAND2_X1 U9854 ( .A1(n10428), .A2(n7398), .ZN(n10430) );
  INV_X1 U9855 ( .A(n7398), .ZN(n10332) );
  XNOR2_X1 U9856 ( .A(n10428), .B(n7398), .ZN(n10701) );
  NAND2_X1 U9857 ( .A1(n11225), .A2(n11257), .ZN(n7399) );
  NAND2_X1 U9858 ( .A1(n10660), .A2(n10659), .ZN(n10758) );
  NAND2_X1 U9859 ( .A1(n10645), .A2(n10644), .ZN(n10660) );
  NAND2_X1 U9860 ( .A1(n10433), .A2(n10432), .ZN(n10434) );
  OAI21_X1 U9861 ( .B1(n10505), .B2(n10328), .A(n10326), .ZN(n10428) );
  NAND2_X1 U9862 ( .A1(n13412), .A2(n13240), .ZN(n13406) );
  OAI21_X1 U9863 ( .B1(n10729), .B2(n7409), .A(n10952), .ZN(n10730) );
  NAND2_X1 U9864 ( .A1(n10729), .A2(n7409), .ZN(n10952) );
  XNOR2_X1 U9865 ( .A(n10950), .B(n15201), .ZN(n7409) );
  OAI21_X1 U9866 ( .B1(n11907), .B2(n7413), .A(n6493), .ZN(n12232) );
  NAND2_X1 U9867 ( .A1(n12350), .A2(n7418), .ZN(n7415) );
  NAND3_X1 U9868 ( .A1(n7425), .A2(n10961), .A3(n7424), .ZN(n7423) );
  NAND3_X1 U9869 ( .A1(n7425), .A2(n7428), .A3(n10961), .ZN(n7427) );
  INV_X1 U9870 ( .A(n7427), .ZN(n11209) );
  INV_X1 U9871 ( .A(n10962), .ZN(n7429) );
  OAI211_X1 U9872 ( .C1(n12337), .C2(n7440), .A(n7437), .B(n7435), .ZN(n12209)
         );
  NAND2_X1 U9873 ( .A1(n12337), .A2(n7436), .ZN(n7435) );
  NOR2_X1 U9874 ( .A1(n12203), .A2(n7438), .ZN(n7436) );
  OAI22_X1 U9875 ( .A1(n7439), .A2(n7438), .B1(n12203), .B2(n7441), .ZN(n7437)
         );
  NOR2_X1 U9876 ( .A1(n12203), .A2(n12224), .ZN(n7439) );
  NAND2_X1 U9877 ( .A1(n12224), .A2(n12203), .ZN(n7440) );
  NAND2_X1 U9878 ( .A1(n10945), .A2(n6885), .ZN(n9092) );
  NAND2_X1 U9879 ( .A1(n7466), .A2(n11964), .ZN(n10930) );
  NAND2_X1 U9880 ( .A1(n10860), .A2(n11961), .ZN(n7466) );
  INV_X1 U9881 ( .A(n7469), .ZN(n7468) );
  OAI21_X1 U9882 ( .B1(n11993), .B2(n7477), .A(n7475), .ZN(n11998) );
  NAND2_X1 U9883 ( .A1(n7474), .A2(n7472), .ZN(n11997) );
  NAND2_X1 U9884 ( .A1(n11993), .A2(n7475), .ZN(n7474) );
  NAND2_X1 U9885 ( .A1(n7494), .A2(n7495), .ZN(n12072) );
  NAND3_X1 U9886 ( .A1(n6506), .A2(n7752), .A3(n8584), .ZN(n7564) );
  INV_X1 U9887 ( .A(n9073), .ZN(n9076) );
  NAND3_X1 U9888 ( .A1(n10367), .A2(n6496), .A3(n7523), .ZN(n7519) );
  NAND2_X1 U9889 ( .A1(n7809), .A2(n7929), .ZN(n7520) );
  INV_X1 U9890 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7522) );
  NAND3_X1 U9891 ( .A1(n7532), .A2(n8423), .A3(n8424), .ZN(n8425) );
  NAND2_X1 U9892 ( .A1(n7540), .A2(n15190), .ZN(n7539) );
  NAND2_X1 U9893 ( .A1(n8398), .A2(n8399), .ZN(n7541) );
  AOI21_X1 U9894 ( .B1(n8219), .B2(n8220), .A(n6524), .ZN(n8232) );
  NAND3_X1 U9895 ( .A1(n8219), .A2(n8233), .A3(n7558), .ZN(n7551) );
  NOR2_X1 U9896 ( .A1(n7564), .A2(n8538), .ZN(n7563) );
  NAND2_X1 U9897 ( .A1(n10942), .A2(n7566), .ZN(n7565) );
  NAND2_X1 U9898 ( .A1(n14095), .A2(n7585), .ZN(n14074) );
  OAI21_X1 U9899 ( .B1(n8705), .B2(n7597), .A(n7595), .ZN(n8739) );
  NAND2_X1 U9900 ( .A1(n8569), .A2(SI_1_), .ZN(n8579) );
  OAI21_X1 U9901 ( .B1(n9053), .B2(n9052), .A(n9056), .ZN(n9672) );
  AOI21_X1 U9902 ( .B1(n9052), .B2(n9056), .A(n7621), .ZN(n7620) );
  NAND2_X1 U9903 ( .A1(n14909), .A2(n7622), .ZN(n10509) );
  OR2_X1 U9904 ( .A1(n7624), .A2(n10499), .ZN(n7622) );
  NOR3_X1 U9905 ( .A1(n13012), .A2(n10506), .A3(n7624), .ZN(n10507) );
  NAND2_X1 U9906 ( .A1(n14546), .A2(n7630), .ZN(n7629) );
  NAND2_X1 U9907 ( .A1(n9217), .A2(n7661), .ZN(n9232) );
  NAND2_X1 U9908 ( .A1(n9217), .A2(n9220), .ZN(n9230) );
  INV_X1 U9909 ( .A(n8506), .ZN(n7663) );
  NOR2_X1 U9910 ( .A1(n12610), .A2(n8516), .ZN(n12596) );
  AND2_X1 U9911 ( .A1(n7688), .A2(n7687), .ZN(n12219) );
  INV_X1 U9912 ( .A(n9172), .ZN(n7688) );
  NAND2_X1 U9913 ( .A1(n8441), .A2(n7699), .ZN(n12885) );
  NAND2_X1 U9914 ( .A1(n9166), .A2(n9165), .ZN(n9168) );
  NAND3_X1 U9915 ( .A1(n8487), .A2(n8488), .A3(n8486), .ZN(n10740) );
  OAI21_X1 U9916 ( .B1(n7769), .B2(n9804), .A(n7701), .ZN(n9817) );
  NAND2_X1 U9917 ( .A1(n7703), .A2(n7702), .ZN(n7701) );
  OAI22_X1 U9918 ( .A1(n7711), .A2(n7709), .B1(n9455), .B2(n7708), .ZN(n9472)
         );
  INV_X1 U9919 ( .A(n9454), .ZN(n7708) );
  NOR2_X1 U9920 ( .A1(n9454), .A2(n7710), .ZN(n7709) );
  INV_X1 U9921 ( .A(n9455), .ZN(n7710) );
  OAI21_X1 U9922 ( .B1(n9304), .B2(n9303), .A(n9302), .ZN(n7716) );
  INV_X1 U9923 ( .A(n9393), .ZN(n7718) );
  NAND2_X1 U9924 ( .A1(n9423), .A2(n6565), .ZN(n7719) );
  NAND2_X1 U9925 ( .A1(n9209), .A2(n7720), .ZN(n13569) );
  NAND2_X1 U9926 ( .A1(n13793), .A2(n7727), .ZN(n7725) );
  NAND2_X1 U9927 ( .A1(n13793), .A2(n13794), .ZN(n7726) );
  NAND2_X1 U9928 ( .A1(n14603), .A2(n7736), .ZN(n7735) );
  INV_X1 U9929 ( .A(n11777), .ZN(n7747) );
  NAND2_X2 U9930 ( .A1(n8947), .A2(n9676), .ZN(n12088) );
  NAND2_X2 U9931 ( .A1(n8947), .A2(n9211), .ZN(n8727) );
  NAND2_X1 U9932 ( .A1(n7753), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8559) );
  INV_X4 U9933 ( .A(n9589), .ZN(n9750) );
  INV_X1 U9934 ( .A(n11918), .ZN(n11921) );
  NAND2_X1 U9935 ( .A1(n12047), .A2(n12046), .ZN(n12048) );
  NAND2_X1 U9936 ( .A1(n10184), .A2(n10342), .ZN(n10187) );
  OAI21_X1 U9937 ( .B1(n9811), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9813) );
  INV_X1 U9938 ( .A(n8899), .ZN(n8878) );
  INV_X1 U9939 ( .A(n7788), .ZN(n7790) );
  OR2_X1 U9940 ( .A1(n8236), .A2(n10399), .ZN(n7816) );
  NAND4_X2 U9941 ( .A1(n8578), .A2(n8575), .A3(n8576), .A4(n8577), .ZN(n13895)
         );
  NAND2_X1 U9942 ( .A1(n13645), .A2(n13647), .ZN(n13648) );
  INV_X1 U9943 ( .A(n9373), .ZN(n9376) );
  INV_X4 U9944 ( .A(n8915), .ZN(n9060) );
  INV_X1 U9945 ( .A(n12718), .ZN(n15214) );
  INV_X1 U9946 ( .A(n15194), .ZN(n12749) );
  OR2_X1 U9947 ( .A1(n13254), .A2(n13317), .ZN(n7754) );
  AND2_X1 U9948 ( .A1(n12849), .A2(n12656), .ZN(n7755) );
  AND4_X1 U9949 ( .A1(n8815), .A2(n8741), .A3(n8707), .A4(n8819), .ZN(n7756)
         );
  AND2_X1 U9950 ( .A1(n12866), .A2(n12691), .ZN(n7757) );
  AND4_X1 U9951 ( .A1(n7778), .A2(n8248), .A3(n7777), .A4(n8078), .ZN(n7758)
         );
  INV_X1 U9952 ( .A(n13198), .ZN(n14539) );
  NAND2_X1 U9953 ( .A1(n8447), .A2(n8446), .ZN(n11825) );
  AND2_X1 U9954 ( .A1(n13248), .A2(n10457), .ZN(n7759) );
  INV_X1 U9955 ( .A(SI_24_), .ZN(n11824) );
  OR2_X1 U9956 ( .A1(n12144), .A2(n12102), .ZN(n7761) );
  INV_X1 U9957 ( .A(n13226), .ZN(n12921) );
  INV_X1 U9958 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n14179) );
  INV_X1 U9959 ( .A(n12626), .ZN(n12187) );
  OR2_X1 U9960 ( .A1(n8941), .A2(SI_21_), .ZN(n7764) );
  INV_X1 U9961 ( .A(n14060), .ZN(n14075) );
  INV_X1 U9962 ( .A(n12792), .ZN(n8512) );
  INV_X1 U9963 ( .A(n15196), .ZN(n7814) );
  AND2_X1 U9964 ( .A1(n8715), .A2(n8714), .ZN(n7765) );
  OR2_X1 U9965 ( .A1(n12214), .A2(n14521), .ZN(n7766) );
  AND2_X1 U9966 ( .A1(n12586), .A2(n15222), .ZN(n14521) );
  INV_X1 U9967 ( .A(n14521), .ZN(n8531) );
  AND2_X1 U9968 ( .A1(n11540), .A2(n11539), .ZN(n7767) );
  OR2_X1 U9969 ( .A1(n8939), .A2(SI_20_), .ZN(n7768) );
  OR2_X1 U9970 ( .A1(n9803), .A2(n9247), .ZN(n7769) );
  NAND2_X1 U9971 ( .A1(n10568), .A2(n15070), .ZN(n13446) );
  OR4_X1 U9972 ( .A1(n15084), .A2(n14541), .A3(n13584), .A4(n9880), .ZN(n7770)
         );
  NAND3_X1 U9973 ( .A1(n9270), .A2(n9269), .A3(n9268), .ZN(n9299) );
  NAND2_X1 U9974 ( .A1(n9340), .A2(n9339), .ZN(n9342) );
  INV_X1 U9975 ( .A(n9374), .ZN(n9375) );
  OAI21_X1 U9976 ( .B1(n9293), .B2(n11356), .A(n9422), .ZN(n9423) );
  AND2_X1 U9977 ( .A1(n12017), .A2(n12009), .ZN(n12010) );
  NAND2_X1 U9978 ( .A1(n12062), .A2(n12061), .ZN(n12063) );
  AOI21_X1 U9979 ( .B1(n9580), .B2(n9579), .A(n9578), .ZN(n9582) );
  INV_X1 U9980 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7777) );
  INV_X1 U9981 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n9196) );
  INV_X1 U9982 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n15422) );
  INV_X1 U9983 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9206) );
  INV_X1 U9984 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n9223) );
  INV_X1 U9985 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8898) );
  INV_X1 U9986 ( .A(n8067), .ZN(n8068) );
  INV_X1 U9987 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n7774) );
  INV_X1 U9988 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9384) );
  INV_X1 U9989 ( .A(n9240), .ZN(n9242) );
  INV_X1 U9990 ( .A(n13079), .ZN(n11721) );
  INV_X1 U9991 ( .A(n10222), .ZN(n10223) );
  OR2_X1 U9992 ( .A1(n13640), .A2(n13639), .ZN(n13641) );
  INV_X1 U9993 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8764) );
  INV_X1 U9994 ( .A(n12120), .ZN(n8646) );
  NAND2_X1 U9995 ( .A1(n7768), .A2(n7764), .ZN(n8944) );
  INV_X1 U9996 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n8030) );
  OR2_X1 U9997 ( .A1(n11679), .A2(n11678), .ZN(n11686) );
  INV_X1 U9998 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n15410) );
  INV_X1 U9999 ( .A(n8364), .ZN(n8103) );
  NAND2_X1 U10000 ( .A1(n8043), .A2(n15410), .ZN(n8056) );
  INV_X1 U10001 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n15429) );
  NOR2_X1 U10002 ( .A1(n15246), .A2(n8214), .ZN(n9175) );
  NAND2_X1 U10003 ( .A1(n8301), .A2(n8300), .ZN(n10840) );
  AND2_X1 U10004 ( .A1(n9643), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n9644) );
  NOR2_X1 U10005 ( .A1(n9568), .A2(n13019), .ZN(n9585) );
  OR2_X1 U10006 ( .A1(n15010), .A2(n15009), .ZN(n15006) );
  INV_X1 U10007 ( .A(n9877), .ZN(n9878) );
  INV_X1 U10008 ( .A(n9247), .ZN(n9550) );
  INV_X1 U10009 ( .A(n11131), .ZN(n11130) );
  NAND2_X1 U10010 ( .A1(n14562), .A2(n9550), .ZN(n9877) );
  NAND2_X1 U10011 ( .A1(n9813), .A2(n9812), .ZN(n9818) );
  INV_X1 U10012 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8784) );
  NAND2_X1 U10013 ( .A1(n10223), .A2(n13604), .ZN(n10224) );
  INV_X1 U10014 ( .A(n13773), .ZN(n13682) );
  OR2_X1 U10015 ( .A1(n13654), .A2(n13653), .ZN(n13655) );
  NOR2_X1 U10016 ( .A1(n8913), .A2(n13826), .ZN(n8931) );
  OR2_X1 U10017 ( .A1(n9953), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9141) );
  INV_X1 U10018 ( .A(n14073), .ZN(n8937) );
  AOI21_X1 U10019 ( .B1(n13958), .B2(n14269), .A(n9129), .ZN(n9130) );
  OR2_X1 U10020 ( .A1(n9953), .A2(n10191), .ZN(n10172) );
  INV_X1 U10021 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8541) );
  AND2_X1 U10022 ( .A1(n8031), .A2(n8030), .ZN(n8043) );
  INV_X1 U10023 ( .A(n15441), .ZN(n12353) );
  INV_X1 U10024 ( .A(n12330), .ZN(n12351) );
  OR2_X1 U10025 ( .A1(n8211), .A2(n12572), .ZN(n8191) );
  INV_X1 U10026 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n11690) );
  INV_X1 U10027 ( .A(n12602), .ZN(n12595) );
  AND4_X1 U10028 ( .A1(n8060), .A2(n8059), .A3(n8058), .A4(n8057), .ZN(n15441)
         );
  OR2_X1 U10029 ( .A1(n14497), .A2(n14520), .ZN(n8341) );
  INV_X1 U10030 ( .A(n15209), .ZN(n12746) );
  INV_X1 U10031 ( .A(n12882), .ZN(n9188) );
  INV_X1 U10032 ( .A(n15200), .ZN(n15182) );
  NAND2_X1 U10033 ( .A1(n9644), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n9712) );
  INV_X1 U10034 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9238) );
  INV_X1 U10035 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10453) );
  AND2_X1 U10036 ( .A1(n9747), .A2(n9834), .ZN(n9997) );
  AND2_X1 U10037 ( .A1(n9700), .A2(n9699), .ZN(n12973) );
  OR2_X1 U10038 ( .A1(n9556), .A2(n9555), .ZN(n9568) );
  OR2_X1 U10039 ( .A1(n9994), .A2(n9995), .ZN(n10237) );
  AND2_X1 U10040 ( .A1(n10237), .A2(n10236), .ZN(n14985) );
  INV_X1 U10041 ( .A(n13225), .ZN(n13494) );
  INV_X1 U10042 ( .A(n11919), .ZN(n11920) );
  INV_X1 U10043 ( .A(n13078), .ZN(n14542) );
  INV_X1 U10044 ( .A(n14562), .ZN(n13459) );
  AND2_X1 U10045 ( .A1(n15090), .A2(n9880), .ZN(n15123) );
  NAND2_X1 U10046 ( .A1(n9818), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9819) );
  INV_X1 U10047 ( .A(n13737), .ZN(n10804) );
  INV_X1 U10048 ( .A(n14625), .ZN(n13846) );
  AND2_X1 U10049 ( .A1(n9141), .A2(n9954), .ZN(n10850) );
  AND2_X1 U10050 ( .A1(n13948), .A2(n9047), .ZN(n13764) );
  AND2_X1 U10051 ( .A1(n8882), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8903) );
  INV_X1 U10052 ( .A(n8947), .ZN(n9950) );
  INV_X1 U10053 ( .A(n9109), .ZN(n14066) );
  OR2_X1 U10054 ( .A1(n9953), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9160) );
  INV_X1 U10055 ( .A(n14872), .ZN(n14881) );
  AND2_X1 U10056 ( .A1(n10856), .A2(n9162), .ZN(n14872) );
  NOR2_X1 U10057 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n14411), .ZN(n14360) );
  OR2_X1 U10058 ( .A1(n7953), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7968) );
  NOR2_X1 U10059 ( .A1(n7988), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8012) );
  CLKBUF_X1 U10060 ( .A(n12334), .Z(n12358) );
  OR2_X1 U10061 ( .A1(n8211), .A2(n12213), .ZN(n8240) );
  AND4_X1 U10062 ( .A1(n8125), .A2(n8124), .A3(n8123), .A4(n8122), .ZN(n12667)
         );
  AND4_X1 U10063 ( .A1(n8091), .A2(n8090), .A3(n8089), .A4(n8088), .ZN(n12707)
         );
  INV_X1 U10064 ( .A(n15147), .ZN(n15175) );
  INV_X1 U10065 ( .A(n15150), .ZN(n15173) );
  INV_X1 U10066 ( .A(n15183), .ZN(n15203) );
  INV_X1 U10067 ( .A(n12663), .ZN(n14509) );
  NAND2_X1 U10068 ( .A1(n11195), .A2(n12746), .ZN(n12718) );
  AND3_X1 U10069 ( .A1(n9181), .A2(n9180), .A3(n9179), .ZN(n11191) );
  INV_X1 U10070 ( .A(n15195), .ZN(n15188) );
  INV_X1 U10071 ( .A(n15222), .ZN(n15242) );
  NAND2_X1 U10072 ( .A1(n8431), .A2(n8444), .ZN(n10672) );
  AND2_X1 U10073 ( .A1(n9634), .A2(n9657), .ZN(n13332) );
  AND3_X1 U10074 ( .A1(n9753), .A2(n9752), .A3(n9751), .ZN(n13231) );
  OR2_X1 U10075 ( .A1(n13358), .A2(n9605), .ZN(n9611) );
  INV_X1 U10076 ( .A(n15022), .ZN(n15035) );
  OR2_X1 U10077 ( .A1(n14947), .A2(P2_U3088), .ZN(n15037) );
  INV_X1 U10078 ( .A(n13171), .ZN(n15013) );
  INV_X1 U10079 ( .A(n13220), .ZN(n13382) );
  INV_X1 U10080 ( .A(n13310), .ZN(n13384) );
  INV_X1 U10081 ( .A(n15123), .ZN(n15114) );
  AND2_X1 U10082 ( .A1(n10200), .A2(n15107), .ZN(n14576) );
  AND2_X1 U10083 ( .A1(n11220), .A2(n11133), .ZN(n15118) );
  AND2_X1 U10084 ( .A1(n9996), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9824) );
  AND2_X1 U10085 ( .A1(n10197), .A2(n10851), .ZN(n14625) );
  AND4_X1 U10086 ( .A1(n8953), .A2(n8952), .A3(n8951), .A4(n8950), .ZN(n13774)
         );
  INV_X1 U10087 ( .A(n14749), .ZN(n14772) );
  INV_X1 U10088 ( .A(n14818), .ZN(n14849) );
  NAND2_X1 U10089 ( .A1(n13950), .A2(n14831), .ZN(n14165) );
  AND2_X1 U10090 ( .A1(n9160), .A2(n9957), .ZN(n10256) );
  INV_X1 U10091 ( .A(n14887), .ZN(n14273) );
  AND2_X1 U10092 ( .A1(n14891), .A2(n14881), .ZN(n14306) );
  INV_X1 U10093 ( .A(n10256), .ZN(n10852) );
  AND2_X1 U10094 ( .A1(n8728), .A2(n8711), .ZN(n10474) );
  AND2_X1 U10095 ( .A1(n14435), .A2(n14434), .ZN(n14657) );
  AND2_X1 U10096 ( .A1(n10373), .A2(n10372), .ZN(n15168) );
  AOI22_X1 U10097 ( .A1(n10680), .A2(P3_STATE_REG_SCAN_IN), .B1(n10691), .B2(
        n10679), .ZN(n12332) );
  AND4_X1 U10098 ( .A1(n8240), .A2(n8218), .A3(n8217), .A4(n8216), .ZN(n12205)
         );
  INV_X1 U10099 ( .A(n12707), .ZN(n12366) );
  INV_X1 U10100 ( .A(n12547), .ZN(n15164) );
  OR2_X1 U10101 ( .A1(n10365), .A2(n10359), .ZN(n15162) );
  NAND2_X1 U10102 ( .A1(n12749), .A2(n14489), .ZN(n12663) );
  INV_X1 U10103 ( .A(n12718), .ZN(n15194) );
  NAND2_X1 U10104 ( .A1(n15254), .A2(n15188), .ZN(n12829) );
  AND2_X1 U10105 ( .A1(n8481), .A2(n8480), .ZN(n15244) );
  INV_X2 U10106 ( .A(n15244), .ZN(n15246) );
  NAND2_X1 U10107 ( .A1(n8443), .A2(n8442), .ZN(n12904) );
  INV_X1 U10108 ( .A(SI_19_), .ZN(n10426) );
  INV_X1 U10109 ( .A(SI_13_), .ZN(n9944) );
  INV_X1 U10110 ( .A(n10558), .ZN(n10409) );
  INV_X1 U10111 ( .A(n13482), .ZN(n13317) );
  INV_X1 U10112 ( .A(n14916), .ZN(n12998) );
  OR2_X1 U10113 ( .A1(n9520), .A2(n9519), .ZN(n13236) );
  INV_X1 U10114 ( .A(P2_U3947), .ZN(n13083) );
  INV_X1 U10115 ( .A(n15043), .ZN(n15008) );
  OR2_X1 U10116 ( .A1(n10002), .A2(P2_U3088), .ZN(n15046) );
  OR2_X1 U10117 ( .A1(n15076), .A2(n10566), .ZN(n13427) );
  AND2_X1 U10118 ( .A1(n11619), .A2(n11618), .ZN(n14586) );
  INV_X1 U10119 ( .A(n15059), .ZN(n13448) );
  INV_X1 U10120 ( .A(n15145), .ZN(n15142) );
  AND2_X1 U10121 ( .A1(n14586), .A2(n14585), .ZN(n14593) );
  INV_X1 U10122 ( .A(n15134), .ZN(n15132) );
  NAND2_X1 U10123 ( .A1(n15082), .A2(n15078), .ZN(n15080) );
  INV_X1 U10124 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11327) );
  INV_X1 U10125 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10233) );
  INV_X1 U10126 ( .A(n11991), .ZN(n14797) );
  NAND2_X1 U10127 ( .A1(n10197), .A2(n10196), .ZN(n13868) );
  INV_X1 U10128 ( .A(n13774), .ZN(n13878) );
  OR2_X2 U10129 ( .A1(n9832), .A2(n10185), .ZN(n13896) );
  INV_X1 U10130 ( .A(n14673), .ZN(n14781) );
  OR2_X1 U10131 ( .A1(n14842), .A2(n10856), .ZN(n14845) );
  OR2_X1 U10132 ( .A1(n14842), .A2(n14885), .ZN(n14143) );
  INV_X1 U10133 ( .A(n14230), .ZN(n14210) );
  AND2_X2 U10134 ( .A1(n10257), .A2(n10256), .ZN(n14896) );
  INV_X1 U10135 ( .A(n14306), .ZN(n14297) );
  INV_X1 U10136 ( .A(n14891), .ZN(n14889) );
  AND2_X1 U10137 ( .A1(n10175), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9958) );
  INV_X1 U10138 ( .A(n9154), .ZN(n14344) );
  INV_X1 U10139 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10215) );
  NOR2_X2 U10140 ( .A1(n10673), .A2(n12881), .ZN(P3_U3897) );
  NAND2_X1 U10141 ( .A1(n8454), .A2(n8453), .ZN(P3_U3296) );
  AND2_X1 U10142 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10000), .ZN(P2_U3947) );
  INV_X1 U10143 ( .A(n13896), .ZN(P1_U4016) );
  NOR2_X1 U10144 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), 
        .ZN(n7778) );
  NAND2_X1 U10145 ( .A1(n7799), .A2(n7782), .ZN(n7783) );
  NAND2_X1 U10146 ( .A1(n7843), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n7795) );
  INV_X1 U10147 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n15146) );
  OR2_X1 U10148 ( .A1(n7846), .A2(n15146), .ZN(n7794) );
  INV_X1 U10149 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10360) );
  NAND2_X4 U10150 ( .A1(n7790), .A2(n12223), .ZN(n8236) );
  INV_X1 U10151 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n7791) );
  OR2_X1 U10152 ( .A1(n8236), .A2(n7791), .ZN(n7792) );
  INV_X1 U10153 ( .A(n7821), .ZN(n7797) );
  INV_X1 U10154 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U10155 ( .A1(n8557), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7796) );
  NAND2_X1 U10156 ( .A1(n7797), .A2(n7796), .ZN(n7798) );
  MUX2_X1 U10157 ( .A(n7798), .B(SI_0_), .S(n9676), .Z(n12905) );
  XNOR2_X2 U10158 ( .A(n7803), .B(n7802), .ZN(n12539) );
  MUX2_X1 U10159 ( .A(P3_IR_REG_0__SCAN_IN), .B(n12905), .S(n7824), .Z(n11196)
         );
  INV_X1 U10160 ( .A(n15198), .ZN(n7813) );
  INV_X1 U10161 ( .A(n7844), .ZN(n7804) );
  INV_X1 U10162 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10723) );
  NAND2_X1 U10163 ( .A1(n7843), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7806) );
  INV_X1 U10164 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10378) );
  XNOR2_X1 U10165 ( .A(n7820), .B(n7821), .ZN(n9891) );
  NAND2_X1 U10166 ( .A1(n7853), .A2(n9891), .ZN(n7812) );
  INV_X1 U10167 ( .A(SI_1_), .ZN(n9892) );
  OR2_X1 U10168 ( .A1(n7833), .A2(n9892), .ZN(n7811) );
  INV_X1 U10169 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7809) );
  OR2_X1 U10170 ( .A1(n7824), .A2(n10382), .ZN(n7810) );
  AND3_X2 U10171 ( .A1(n7812), .A2(n7811), .A3(n7810), .ZN(n15196) );
  NAND2_X1 U10172 ( .A1(n12374), .A2(n15196), .ZN(n8406) );
  NAND2_X1 U10173 ( .A1(n7813), .A2(n8406), .ZN(n10715) );
  NAND2_X1 U10174 ( .A1(n10715), .A2(n8407), .ZN(n15181) );
  NAND2_X1 U10175 ( .A1(n7843), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n7819) );
  INV_X1 U10176 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10733) );
  OR2_X1 U10177 ( .A1(n7846), .A2(n10733), .ZN(n7818) );
  INV_X1 U10178 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10405) );
  OR2_X1 U10179 ( .A1(n7844), .A2(n10405), .ZN(n7817) );
  INV_X1 U10180 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10399) );
  INV_X1 U10181 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9896) );
  NAND2_X1 U10182 ( .A1(n9896), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7822) );
  XNOR2_X1 U10183 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n7834) );
  INV_X1 U10184 ( .A(n7834), .ZN(n7823) );
  XNOR2_X1 U10185 ( .A(n7835), .B(n7823), .ZN(n9923) );
  NAND2_X1 U10186 ( .A1(n7853), .A2(n9923), .ZN(n7826) );
  AND2_X1 U10187 ( .A1(n10361), .A2(n7268), .ZN(n7837) );
  NAND2_X1 U10188 ( .A1(n15201), .A2(n10724), .ZN(n8295) );
  NAND2_X1 U10189 ( .A1(n8291), .A2(n8295), .ZN(n8485) );
  NAND2_X1 U10190 ( .A1(n15181), .A2(n15180), .ZN(n15179) );
  NAND2_X1 U10191 ( .A1(n15179), .A2(n8291), .ZN(n10736) );
  NAND2_X1 U10192 ( .A1(n7843), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n7832) );
  OR2_X1 U10193 ( .A1(n7846), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n7831) );
  INV_X1 U10194 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n7827) );
  INV_X1 U10195 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n7828) );
  OR2_X1 U10196 ( .A1(n8236), .A2(n7828), .ZN(n7829) );
  INV_X1 U10197 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9905) );
  NAND2_X1 U10198 ( .A1(n9905), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7836) );
  XNOR2_X1 U10199 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n7854) );
  XNOR2_X1 U10200 ( .A(n7855), .B(n7536), .ZN(n9925) );
  NAND2_X1 U10201 ( .A1(n7853), .A2(n9925), .ZN(n7842) );
  INV_X1 U10202 ( .A(n7837), .ZN(n7839) );
  NAND2_X1 U10203 ( .A1(n7839), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7838) );
  MUX2_X1 U10204 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7838), .S(
        P3_IR_REG_3__SCAN_IN), .Z(n7840) );
  NAND2_X1 U10205 ( .A1(n10960), .A2(n11640), .ZN(n8297) );
  NAND2_X1 U10206 ( .A1(n10736), .A2(n10738), .ZN(n10735) );
  NAND2_X1 U10207 ( .A1(n10735), .A2(n8299), .ZN(n10838) );
  NAND2_X1 U10208 ( .A1(n8224), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n7852) );
  INV_X1 U10209 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n7845) );
  OR2_X1 U10210 ( .A1(n7844), .A2(n7845), .ZN(n7851) );
  NOR2_X1 U10211 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n7864) );
  AND2_X1 U10212 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7847) );
  NOR2_X1 U10213 ( .A1(n7864), .A2(n7847), .ZN(n11626) );
  OR2_X1 U10214 ( .A1(n8211), .A2(n11626), .ZN(n7850) );
  INV_X1 U10215 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n7848) );
  OR2_X1 U10216 ( .A1(n8236), .A2(n7848), .ZN(n7849) );
  NAND4_X1 U10217 ( .A1(n7852), .A2(n7851), .A3(n7850), .A4(n7849), .ZN(n12373) );
  XNOR2_X1 U10218 ( .A(n7872), .B(n6724), .ZN(n9921) );
  NAND2_X1 U10219 ( .A1(n6474), .A2(n9921), .ZN(n7862) );
  NAND2_X1 U10220 ( .A1(n7857), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7856) );
  MUX2_X1 U10221 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7856), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n7860) );
  INV_X1 U10222 ( .A(n7857), .ZN(n7859) );
  INV_X1 U10223 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7858) );
  NAND2_X1 U10224 ( .A1(n7859), .A2(n7858), .ZN(n7875) );
  NAND2_X1 U10225 ( .A1(n7860), .A2(n7875), .ZN(n10412) );
  INV_X1 U10226 ( .A(n10412), .ZN(n10527) );
  OR2_X1 U10227 ( .A1(n10356), .A2(n10527), .ZN(n7861) );
  OAI211_X1 U10228 ( .C1(n7833), .C2(SI_4_), .A(n7862), .B(n7861), .ZN(n11627)
         );
  OR2_X1 U10229 ( .A1(n12373), .A2(n11627), .ZN(n8301) );
  NAND2_X1 U10230 ( .A1(n12373), .A2(n11627), .ZN(n8300) );
  INV_X1 U10231 ( .A(n10840), .ZN(n10837) );
  NAND2_X1 U10232 ( .A1(n10838), .A2(n10837), .ZN(n10836) );
  NAND2_X1 U10233 ( .A1(n8224), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n7870) );
  INV_X1 U10234 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n7863) );
  OR2_X1 U10235 ( .A1(n7844), .A2(n7863), .ZN(n7869) );
  NAND2_X1 U10236 ( .A1(n7864), .A2(n10416), .ZN(n7880) );
  OR2_X1 U10237 ( .A1(n7864), .A2(n10416), .ZN(n7865) );
  AND2_X1 U10238 ( .A1(n7880), .A2(n7865), .ZN(n11312) );
  OR2_X1 U10239 ( .A1(n7846), .A2(n11312), .ZN(n7868) );
  INV_X1 U10240 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n7866) );
  OR2_X1 U10241 ( .A1(n8236), .A2(n7866), .ZN(n7867) );
  NAND4_X1 U10242 ( .A1(n7870), .A2(n7869), .A3(n7868), .A4(n7867), .ZN(n12372) );
  NAND2_X1 U10243 ( .A1(n9904), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7873) );
  XNOR2_X1 U10244 ( .A(n6881), .B(P2_DATAO_REG_5__SCAN_IN), .ZN(n7874) );
  XNOR2_X1 U10245 ( .A(n7888), .B(n7874), .ZN(n9895) );
  NAND2_X1 U10246 ( .A1(n6474), .A2(n9895), .ZN(n7878) );
  NAND2_X1 U10247 ( .A1(n7875), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7876) );
  XNOR2_X1 U10248 ( .A(n7876), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10413) );
  OR2_X1 U10249 ( .A1(n10356), .A2(n10413), .ZN(n7877) );
  OAI211_X1 U10250 ( .C1(n7833), .C2(SI_5_), .A(n7878), .B(n7877), .ZN(n11210)
         );
  NAND2_X1 U10251 ( .A1(n12372), .A2(n11210), .ZN(n8306) );
  NAND2_X1 U10252 ( .A1(n8224), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n7886) );
  INV_X1 U10253 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n7879) );
  OR2_X1 U10254 ( .A1(n8212), .A2(n7879), .ZN(n7885) );
  NAND2_X1 U10255 ( .A1(n7880), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7881) );
  AND2_X1 U10256 ( .A1(n7899), .A2(n7881), .ZN(n11646) );
  OR2_X1 U10257 ( .A1(n8211), .A2(n11646), .ZN(n7884) );
  INV_X1 U10258 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n7882) );
  OR2_X1 U10259 ( .A1(n8236), .A2(n7882), .ZN(n7883) );
  NAND4_X1 U10260 ( .A1(n7886), .A2(n7885), .A3(n7884), .A4(n7883), .ZN(n12371) );
  INV_X1 U10261 ( .A(n7906), .ZN(n7889) );
  XNOR2_X1 U10262 ( .A(n7907), .B(n7889), .ZN(n9888) );
  NAND2_X1 U10263 ( .A1(n6474), .A2(n9888), .ZN(n7897) );
  INV_X1 U10264 ( .A(SI_6_), .ZN(n9889) );
  OR2_X1 U10265 ( .A1(n7833), .A2(n9889), .ZN(n7896) );
  NAND2_X1 U10266 ( .A1(n7890), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7891) );
  MUX2_X1 U10267 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7891), .S(
        P3_IR_REG_6__SCAN_IN), .Z(n7894) );
  NAND2_X1 U10268 ( .A1(n7894), .A2(n7893), .ZN(n10780) );
  OR2_X1 U10269 ( .A1(n10356), .A2(n10780), .ZN(n7895) );
  NAND2_X1 U10270 ( .A1(n12371), .A2(n11647), .ZN(n8313) );
  NAND2_X1 U10271 ( .A1(n8314), .A2(n8313), .ZN(n11242) );
  INV_X1 U10272 ( .A(n11242), .ZN(n11239) );
  NAND2_X1 U10273 ( .A1(n11238), .A2(n8314), .ZN(n11285) );
  NAND2_X1 U10274 ( .A1(n8224), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n7905) );
  INV_X1 U10275 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n7898) );
  OR2_X1 U10276 ( .A1(n8212), .A2(n7898), .ZN(n7904) );
  AND2_X1 U10277 ( .A1(n7899), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7900) );
  NOR2_X1 U10278 ( .A1(n7917), .A2(n7900), .ZN(n11633) );
  OR2_X1 U10279 ( .A1(n8211), .A2(n11633), .ZN(n7903) );
  INV_X1 U10280 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n7901) );
  OR2_X1 U10281 ( .A1(n8236), .A2(n7901), .ZN(n7902) );
  NAND4_X1 U10282 ( .A1(n7905), .A2(n7904), .A3(n7903), .A4(n7902), .ZN(n12370) );
  NAND2_X1 U10283 ( .A1(n9926), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7908) );
  NAND2_X1 U10284 ( .A1(n7909), .A2(n7908), .ZN(n7925) );
  XNOR2_X1 U10285 ( .A(n7925), .B(n7924), .ZN(n9909) );
  NAND2_X1 U10286 ( .A1(n6474), .A2(n9909), .ZN(n7915) );
  NAND2_X1 U10287 ( .A1(n7893), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7910) );
  MUX2_X1 U10288 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7910), .S(
        P3_IR_REG_7__SCAN_IN), .Z(n7913) );
  INV_X1 U10289 ( .A(n7911), .ZN(n7912) );
  NAND2_X1 U10290 ( .A1(n7913), .A2(n7912), .ZN(n11159) );
  INV_X1 U10291 ( .A(n11159), .ZN(n10772) );
  OR2_X1 U10292 ( .A1(n10356), .A2(n10772), .ZN(n7914) );
  OAI211_X1 U10293 ( .C1(n7833), .C2(SI_7_), .A(n7915), .B(n7914), .ZN(n11634)
         );
  OR2_X1 U10294 ( .A1(n12370), .A2(n11634), .ZN(n8318) );
  NAND2_X1 U10295 ( .A1(n12370), .A2(n11634), .ZN(n8317) );
  NAND2_X1 U10296 ( .A1(n8318), .A2(n8317), .ZN(n11599) );
  INV_X1 U10297 ( .A(n11599), .ZN(n11284) );
  NAND2_X1 U10298 ( .A1(n11285), .A2(n11284), .ZN(n11283) );
  NAND2_X1 U10299 ( .A1(n11283), .A2(n8318), .ZN(n11486) );
  NAND2_X1 U10300 ( .A1(n8224), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7923) );
  INV_X1 U10301 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11155) );
  OR2_X1 U10302 ( .A1(n8212), .A2(n11155), .ZN(n7922) );
  NOR2_X1 U10303 ( .A1(n7917), .A2(n7916), .ZN(n7918) );
  OR2_X1 U10304 ( .A1(n7938), .A2(n7918), .ZN(n11490) );
  INV_X1 U10305 ( .A(n11490), .ZN(n11672) );
  OR2_X1 U10306 ( .A1(n8211), .A2(n11672), .ZN(n7921) );
  INV_X1 U10307 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n7919) );
  OR2_X1 U10308 ( .A1(n8236), .A2(n7919), .ZN(n7920) );
  NAND4_X1 U10309 ( .A1(n7923), .A2(n7922), .A3(n7921), .A4(n7920), .ZN(n12369) );
  NAND2_X1 U10310 ( .A1(n7926), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7927) );
  INV_X1 U10311 ( .A(n7944), .ZN(n7928) );
  XNOR2_X1 U10312 ( .A(n7945), .B(n7928), .ZN(n9897) );
  NAND2_X1 U10313 ( .A1(n6474), .A2(n9897), .ZN(n7936) );
  INV_X1 U10314 ( .A(SI_8_), .ZN(n9898) );
  OR2_X1 U10315 ( .A1(n7833), .A2(n9898), .ZN(n7935) );
  NOR2_X1 U10316 ( .A1(n7911), .A2(n7929), .ZN(n7930) );
  MUX2_X1 U10317 ( .A(n7929), .B(n7930), .S(P3_IR_REG_8__SCAN_IN), .Z(n7931)
         );
  INV_X1 U10318 ( .A(n7931), .ZN(n7933) );
  NAND2_X1 U10319 ( .A1(n7933), .A2(n7932), .ZN(n11406) );
  OR2_X1 U10320 ( .A1(n10356), .A2(n11406), .ZN(n7934) );
  NAND2_X1 U10321 ( .A1(n12369), .A2(n11664), .ZN(n8321) );
  NAND2_X1 U10322 ( .A1(n11486), .A2(n11485), .ZN(n7937) );
  NAND2_X1 U10323 ( .A1(n7937), .A2(n8322), .ZN(n11703) );
  NAND2_X1 U10324 ( .A1(n8224), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7943) );
  INV_X1 U10325 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11402) );
  OR2_X1 U10326 ( .A1(n7844), .A2(n11402), .ZN(n7942) );
  INV_X1 U10327 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11401) );
  OR2_X1 U10328 ( .A1(n8236), .A2(n11401), .ZN(n7941) );
  NAND2_X1 U10329 ( .A1(n7938), .A2(n11690), .ZN(n7953) );
  OR2_X1 U10330 ( .A1(n7938), .A2(n11690), .ZN(n7939) );
  AND2_X1 U10331 ( .A1(n7953), .A2(n7939), .ZN(n11710) );
  OR2_X1 U10332 ( .A1(n8211), .A2(n11710), .ZN(n7940) );
  NAND4_X1 U10333 ( .A1(n7943), .A2(n7942), .A3(n7941), .A4(n7940), .ZN(n12368) );
  NAND2_X1 U10334 ( .A1(n7946), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7947) );
  XNOR2_X1 U10335 ( .A(n7961), .B(n7960), .ZN(n9913) );
  NAND2_X1 U10336 ( .A1(n6474), .A2(n9913), .ZN(n7950) );
  NAND2_X1 U10337 ( .A1(n7932), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7948) );
  XNOR2_X1 U10338 ( .A(n7948), .B(P3_IR_REG_9__SCAN_IN), .ZN(n15174) );
  OR2_X1 U10339 ( .A1(n10356), .A2(n15174), .ZN(n7949) );
  OAI211_X1 U10340 ( .C1(n7833), .C2(SI_9_), .A(n7950), .B(n7949), .ZN(n11709)
         );
  NAND2_X1 U10341 ( .A1(n12368), .A2(n11709), .ZN(n7951) );
  OR2_X1 U10342 ( .A1(n12368), .A2(n11709), .ZN(n7952) );
  NAND2_X1 U10343 ( .A1(n8224), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n7959) );
  INV_X1 U10344 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11397) );
  OR2_X1 U10345 ( .A1(n8212), .A2(n11397), .ZN(n7958) );
  NAND2_X1 U10346 ( .A1(n7953), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7954) );
  AND2_X1 U10347 ( .A1(n7968), .A2(n7954), .ZN(n11804) );
  OR2_X1 U10348 ( .A1(n8211), .A2(n11804), .ZN(n7957) );
  INV_X1 U10349 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n7955) );
  OR2_X1 U10350 ( .A1(n8236), .A2(n7955), .ZN(n7956) );
  NAND4_X1 U10351 ( .A1(n7959), .A2(n7958), .A3(n7957), .A4(n7956), .ZN(n14496) );
  XNOR2_X1 U10352 ( .A(n7975), .B(n7974), .ZN(n9907) );
  NAND2_X1 U10353 ( .A1(n6474), .A2(n9907), .ZN(n7966) );
  OR2_X1 U10354 ( .A1(n7932), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n7979) );
  NAND2_X1 U10355 ( .A1(n7979), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7964) );
  XNOR2_X1 U10356 ( .A(n7964), .B(n7963), .ZN(n11587) );
  INV_X1 U10357 ( .A(n11587), .ZN(n11400) );
  OR2_X1 U10358 ( .A1(n10356), .A2(n11400), .ZN(n7965) );
  OAI211_X1 U10359 ( .C1(n7833), .C2(SI_10_), .A(n7966), .B(n7965), .ZN(n11803) );
  NAND2_X1 U10360 ( .A1(n14496), .A2(n11803), .ZN(n8329) );
  OR2_X1 U10361 ( .A1(n14496), .A2(n11803), .ZN(n8330) );
  NAND2_X1 U10362 ( .A1(n8329), .A2(n8330), .ZN(n11799) );
  NAND2_X1 U10363 ( .A1(n8224), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n7973) );
  INV_X1 U10364 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11582) );
  OR2_X1 U10365 ( .A1(n8212), .A2(n11582), .ZN(n7972) );
  INV_X1 U10366 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n7967) );
  OR2_X1 U10367 ( .A1(n8236), .A2(n7967), .ZN(n7971) );
  NAND2_X1 U10368 ( .A1(n7968), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7969) );
  NAND2_X1 U10369 ( .A1(n7988), .A2(n7969), .ZN(n14500) );
  INV_X1 U10370 ( .A(n14500), .ZN(n11876) );
  OR2_X1 U10371 ( .A1(n8211), .A2(n11876), .ZN(n7970) );
  NAND4_X1 U10372 ( .A1(n7973), .A2(n7972), .A3(n7971), .A4(n7970), .ZN(n12367) );
  NAND2_X1 U10373 ( .A1(n7976), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7977) );
  XNOR2_X1 U10374 ( .A(n7995), .B(n7994), .ZN(n9918) );
  NAND2_X1 U10375 ( .A1(n6474), .A2(n9918), .ZN(n7987) );
  OR2_X1 U10376 ( .A1(n7833), .A2(SI_11_), .ZN(n7986) );
  NOR2_X1 U10377 ( .A1(n7979), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n7982) );
  NOR2_X1 U10378 ( .A1(n7982), .A2(n7929), .ZN(n7980) );
  MUX2_X1 U10379 ( .A(n7929), .B(n7980), .S(P3_IR_REG_11__SCAN_IN), .Z(n7984)
         );
  NAND2_X1 U10380 ( .A1(n7982), .A2(n7981), .ZN(n8006) );
  INV_X1 U10381 ( .A(n8006), .ZN(n7983) );
  INV_X1 U10382 ( .A(n11762), .ZN(n11585) );
  OR2_X1 U10383 ( .A1(n10356), .A2(n11585), .ZN(n7985) );
  INV_X1 U10384 ( .A(n11873), .ZN(n14507) );
  OR2_X1 U10385 ( .A1(n12367), .A2(n14507), .ZN(n8334) );
  NAND2_X1 U10386 ( .A1(n12367), .A2(n14507), .ZN(n8335) );
  NAND2_X1 U10387 ( .A1(n8334), .A2(n8335), .ZN(n14502) );
  INV_X1 U10388 ( .A(n8329), .ZN(n14503) );
  NAND2_X1 U10389 ( .A1(n14505), .A2(n8334), .ZN(n11893) );
  NAND2_X1 U10390 ( .A1(n8224), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n7993) );
  INV_X1 U10391 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11898) );
  OR2_X1 U10392 ( .A1(n8212), .A2(n11898), .ZN(n7992) );
  AND2_X1 U10393 ( .A1(n7988), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7989) );
  NOR2_X1 U10394 ( .A1(n8012), .A2(n7989), .ZN(n11917) );
  OR2_X1 U10395 ( .A1(n8211), .A2(n11917), .ZN(n7991) );
  INV_X1 U10396 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n12376) );
  OR2_X1 U10397 ( .A1(n8236), .A2(n12376), .ZN(n7990) );
  NAND4_X1 U10398 ( .A1(n7993), .A2(n7992), .A3(n7991), .A4(n7990), .ZN(n14497) );
  NAND2_X1 U10399 ( .A1(n7996), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7997) );
  XNOR2_X1 U10400 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n8005) );
  INV_X1 U10401 ( .A(n8005), .ZN(n7998) );
  XNOR2_X1 U10402 ( .A(n8004), .B(n7998), .ZN(n9931) );
  NAND2_X1 U10403 ( .A1(n6474), .A2(n9931), .ZN(n8002) );
  NAND2_X1 U10404 ( .A1(n8006), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7999) );
  XNOR2_X1 U10405 ( .A(n7999), .B(P3_IR_REG_12__SCAN_IN), .ZN(n12377) );
  OR2_X1 U10406 ( .A1(n10356), .A2(n12382), .ZN(n8001) );
  OR2_X1 U10407 ( .A1(n7833), .A2(n9933), .ZN(n8000) );
  NAND2_X1 U10408 ( .A1(n14497), .A2(n14520), .ZN(n8340) );
  NAND2_X1 U10409 ( .A1(n8341), .A2(n8340), .ZN(n11895) );
  INV_X1 U10410 ( .A(n11895), .ZN(n8414) );
  NAND2_X1 U10411 ( .A1(n11893), .A2(n8414), .ZN(n8003) );
  XNOR2_X1 U10412 ( .A(n8019), .B(n10233), .ZN(n9942) );
  NAND2_X1 U10413 ( .A1(n9942), .A2(n6474), .ZN(n8011) );
  NAND2_X1 U10414 ( .A1(n8023), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8008) );
  INV_X1 U10415 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8007) );
  XNOR2_X1 U10416 ( .A(n8008), .B(n8007), .ZN(n12388) );
  OAI22_X1 U10417 ( .A1(n7833), .A2(n9944), .B1(n10356), .B2(n12388), .ZN(
        n8009) );
  INV_X1 U10418 ( .A(n8009), .ZN(n8010) );
  NAND2_X1 U10419 ( .A1(n8011), .A2(n8010), .ZN(n14490) );
  NAND2_X1 U10420 ( .A1(n8224), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8018) );
  INV_X1 U10421 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12385) );
  OR2_X1 U10422 ( .A1(n8212), .A2(n12385), .ZN(n8017) );
  NOR2_X1 U10423 ( .A1(n8012), .A2(n15429), .ZN(n8013) );
  OR2_X1 U10424 ( .A1(n8031), .A2(n8013), .ZN(n14491) );
  INV_X1 U10425 ( .A(n14491), .ZN(n12313) );
  OR2_X1 U10426 ( .A1(n8211), .A2(n12313), .ZN(n8016) );
  INV_X1 U10427 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n8014) );
  OR2_X1 U10428 ( .A1(n8236), .A2(n8014), .ZN(n8015) );
  NAND4_X1 U10429 ( .A1(n8018), .A2(n8017), .A3(n8016), .A4(n8015), .ZN(n12755) );
  INV_X1 U10430 ( .A(n12755), .ZN(n11912) );
  AND2_X1 U10431 ( .A1(n14490), .A2(n11912), .ZN(n8346) );
  OR2_X1 U10432 ( .A1(n14490), .A2(n11912), .ZN(n8345) );
  NAND2_X1 U10433 ( .A1(n8019), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8022) );
  NAND2_X1 U10434 ( .A1(n10215), .A2(n8020), .ZN(n8021) );
  XNOR2_X1 U10435 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8039) );
  XNOR2_X1 U10436 ( .A(n8038), .B(n8039), .ZN(n9947) );
  NAND2_X1 U10437 ( .A1(n9947), .A2(n6474), .ZN(n8028) );
  OAI21_X1 U10438 ( .B1(n8023), .B2(P3_IR_REG_13__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8025) );
  INV_X1 U10439 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8024) );
  XNOR2_X1 U10440 ( .A(n8025), .B(n8024), .ZN(n12436) );
  INV_X1 U10441 ( .A(n12436), .ZN(n12422) );
  OAI22_X1 U10442 ( .A1(n7833), .A2(SI_14_), .B1(n12422), .B2(n10356), .ZN(
        n8026) );
  INV_X1 U10443 ( .A(n8026), .ZN(n8027) );
  NAND2_X1 U10444 ( .A1(n8224), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8037) );
  INV_X1 U10445 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n8029) );
  OR2_X1 U10446 ( .A1(n7844), .A2(n8029), .ZN(n8036) );
  NOR2_X1 U10447 ( .A1(n8031), .A2(n8030), .ZN(n8032) );
  OR2_X1 U10448 ( .A1(n8043), .A2(n8032), .ZN(n12759) );
  INV_X1 U10449 ( .A(n12759), .ZN(n8033) );
  OR2_X1 U10450 ( .A1(n8211), .A2(n8033), .ZN(n8035) );
  INV_X1 U10451 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12827) );
  OR2_X1 U10452 ( .A1(n8236), .A2(n12827), .ZN(n8034) );
  NAND4_X1 U10453 ( .A1(n8037), .A2(n8036), .A3(n8035), .A4(n8034), .ZN(n12737) );
  OR2_X1 U10454 ( .A1(n12879), .A2(n12737), .ZN(n8350) );
  NAND2_X1 U10455 ( .A1(n12879), .A2(n12737), .ZN(n8354) );
  AOI22_X1 U10456 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n10497), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n7095), .ZN(n8050) );
  XOR2_X1 U10457 ( .A(n8049), .B(n8050), .Z(n10068) );
  NAND2_X1 U10458 ( .A1(n8040), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8041) );
  XNOR2_X1 U10459 ( .A(n8041), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12456) );
  INV_X1 U10460 ( .A(n12456), .ZN(n12440) );
  OAI22_X1 U10461 ( .A1(n7833), .A2(n15386), .B1(n10356), .B2(n12440), .ZN(
        n8042) );
  AOI21_X1 U10462 ( .B1(n10068), .B2(n6474), .A(n8042), .ZN(n12745) );
  NAND2_X1 U10463 ( .A1(n8224), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8048) );
  INV_X1 U10464 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12748) );
  OR2_X1 U10465 ( .A1(n8212), .A2(n12748), .ZN(n8047) );
  INV_X1 U10466 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12427) );
  OR2_X1 U10467 ( .A1(n8236), .A2(n12427), .ZN(n8046) );
  OR2_X1 U10468 ( .A1(n8043), .A2(n15410), .ZN(n8044) );
  AND2_X1 U10469 ( .A1(n8044), .A2(n8056), .ZN(n12747) );
  OR2_X1 U10470 ( .A1(n8211), .A2(n12747), .ZN(n8045) );
  NAND4_X1 U10471 ( .A1(n8048), .A2(n8047), .A3(n8046), .A4(n8045), .ZN(n12754) );
  NAND2_X1 U10472 ( .A1(n12745), .A2(n12754), .ZN(n8351) );
  INV_X1 U10473 ( .A(n12745), .ZN(n12873) );
  NAND2_X1 U10474 ( .A1(n12873), .A2(n12726), .ZN(n8356) );
  NAND2_X1 U10475 ( .A1(n8351), .A2(n8356), .ZN(n8418) );
  NAND2_X1 U10476 ( .A1(n12742), .A2(n12741), .ZN(n12744) );
  AOI22_X1 U10477 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n10446), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10464), .ZN(n8062) );
  XNOR2_X1 U10478 ( .A(n8061), .B(n8062), .ZN(n10070) );
  OR2_X1 U10479 ( .A1(n8051), .A2(n7929), .ZN(n8052) );
  XNOR2_X1 U10480 ( .A(n8052), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12459) );
  OAI22_X1 U10481 ( .A1(n7833), .A2(n10071), .B1(n10356), .B2(n12483), .ZN(
        n8053) );
  INV_X1 U10482 ( .A(n8053), .ZN(n8054) );
  OAI21_X1 U10483 ( .B1(n10070), .B2(n8055), .A(n8054), .ZN(n12729) );
  NAND2_X1 U10484 ( .A1(n8224), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8060) );
  AOI21_X1 U10485 ( .B1(n8056), .B2(P3_REG3_REG_16__SCAN_IN), .A(n8067), .ZN(
        n12730) );
  OR2_X1 U10486 ( .A1(n8211), .A2(n12730), .ZN(n8059) );
  INV_X1 U10487 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12731) );
  OR2_X1 U10488 ( .A1(n8212), .A2(n12731), .ZN(n8058) );
  INV_X1 U10489 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12817) );
  OR2_X1 U10490 ( .A1(n8236), .A2(n12817), .ZN(n8057) );
  NAND2_X1 U10491 ( .A1(n12729), .A2(n15441), .ZN(n8357) );
  OR2_X1 U10492 ( .A1(n12729), .A2(n15441), .ZN(n8359) );
  NAND2_X1 U10493 ( .A1(n8357), .A2(n8359), .ZN(n12722) );
  INV_X1 U10494 ( .A(n12722), .ZN(n12727) );
  AOI22_X1 U10495 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n10466), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n7093), .ZN(n8075) );
  XOR2_X1 U10496 ( .A(n8074), .B(n8075), .Z(n10253) );
  INV_X1 U10497 ( .A(SI_17_), .ZN(n10255) );
  NAND2_X1 U10498 ( .A1(n8063), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8064) );
  MUX2_X1 U10499 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8064), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n8065) );
  AND2_X1 U10500 ( .A1(n8065), .A2(n8080), .ZN(n12517) );
  OAI22_X1 U10501 ( .A1(n7833), .A2(n10255), .B1(n10356), .B2(n12509), .ZN(
        n8066) );
  AOI21_X1 U10502 ( .B1(n10253), .B2(n6474), .A(n8066), .ZN(n12715) );
  NAND2_X1 U10503 ( .A1(n8224), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8073) );
  INV_X1 U10504 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12717) );
  OR2_X1 U10505 ( .A1(n8212), .A2(n12717), .ZN(n8072) );
  AND2_X1 U10506 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(n8068), .ZN(n8069) );
  NOR2_X1 U10507 ( .A1(n8086), .A2(n8069), .ZN(n12716) );
  OR2_X1 U10508 ( .A1(n8211), .A2(n12716), .ZN(n8071) );
  INV_X1 U10509 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12485) );
  OR2_X1 U10510 ( .A1(n8236), .A2(n12485), .ZN(n8070) );
  NAND4_X1 U10511 ( .A1(n8073), .A2(n8072), .A3(n8071), .A4(n8070), .ZN(n12691) );
  NAND2_X1 U10512 ( .A1(n12715), .A2(n12691), .ZN(n8277) );
  INV_X1 U10513 ( .A(n12715), .ZN(n12866) );
  NAND2_X1 U10514 ( .A1(n12866), .A2(n12725), .ZN(n12696) );
  AOI22_X1 U10515 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n11021), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n7090), .ZN(n8094) );
  INV_X1 U10516 ( .A(n8094), .ZN(n8077) );
  XNOR2_X1 U10517 ( .A(n8093), .B(n8077), .ZN(n10352) );
  NAND2_X1 U10518 ( .A1(n10352), .A2(n6474), .ZN(n8084) );
  INV_X1 U10519 ( .A(SI_18_), .ZN(n10354) );
  NAND2_X1 U10520 ( .A1(n8080), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8079) );
  MUX2_X1 U10521 ( .A(n8079), .B(P3_IR_REG_31__SCAN_IN), .S(n8078), .Z(n8081)
         );
  NAND2_X1 U10522 ( .A1(n8081), .A2(n8247), .ZN(n12520) );
  OAI22_X1 U10523 ( .A1(n7833), .A2(n10354), .B1(n10356), .B2(n12520), .ZN(
        n8082) );
  INV_X1 U10524 ( .A(n8082), .ZN(n8083) );
  NAND2_X1 U10525 ( .A1(n8084), .A2(n8083), .ZN(n12699) );
  NAND2_X1 U10526 ( .A1(n8224), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8091) );
  INV_X1 U10527 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12701) );
  OR2_X1 U10528 ( .A1(n8212), .A2(n12701), .ZN(n8090) );
  INV_X1 U10529 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n8085) );
  OR2_X1 U10530 ( .A1(n8086), .A2(n8085), .ZN(n8087) );
  NAND2_X1 U10531 ( .A1(n8086), .A2(n8085), .ZN(n8097) );
  AND2_X1 U10532 ( .A1(n8087), .A2(n8097), .ZN(n12700) );
  OR2_X1 U10533 ( .A1(n8211), .A2(n12700), .ZN(n8089) );
  INV_X1 U10534 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12808) );
  OR2_X1 U10535 ( .A1(n8236), .A2(n12808), .ZN(n8088) );
  OR2_X1 U10536 ( .A1(n12699), .A2(n12707), .ZN(n8280) );
  NAND2_X1 U10537 ( .A1(n12699), .A2(n12707), .ZN(n8279) );
  AND2_X1 U10538 ( .A1(n12695), .A2(n12696), .ZN(n8092) );
  NAND2_X1 U10539 ( .A1(n12714), .A2(n8092), .ZN(n12694) );
  NAND2_X1 U10540 ( .A1(n12694), .A2(n8280), .ZN(n12681) );
  INV_X1 U10541 ( .A(n12681), .ZN(n8105) );
  AOI22_X1 U10542 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n11205), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n7005), .ZN(n8107) );
  XNOR2_X1 U10543 ( .A(n8106), .B(n8107), .ZN(n10427) );
  NAND2_X1 U10544 ( .A1(n8247), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8095) );
  OAI22_X1 U10545 ( .A1(n7833), .A2(SI_19_), .B1(n12531), .B2(n10356), .ZN(
        n8096) );
  AOI21_X1 U10546 ( .B1(n10427), .B2(n6474), .A(n8096), .ZN(n12249) );
  INV_X1 U10547 ( .A(n12249), .ZN(n12859) );
  NAND2_X1 U10548 ( .A1(n8224), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8102) );
  INV_X1 U10549 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12683) );
  OR2_X1 U10550 ( .A1(n7844), .A2(n12683), .ZN(n8101) );
  NAND2_X1 U10551 ( .A1(n8097), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8098) );
  AND2_X1 U10552 ( .A1(n8109), .A2(n8098), .ZN(n12682) );
  OR2_X1 U10553 ( .A1(n8211), .A2(n12682), .ZN(n8100) );
  INV_X1 U10554 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12803) );
  OR2_X1 U10555 ( .A1(n8236), .A2(n12803), .ZN(n8099) );
  NAND4_X1 U10556 ( .A1(n8102), .A2(n8101), .A3(n8100), .A4(n8099), .ZN(n12692) );
  AND2_X1 U10557 ( .A1(n12859), .A2(n12692), .ZN(n8365) );
  INV_X1 U10558 ( .A(n8365), .ZN(n8104) );
  OR2_X1 U10559 ( .A1(n12859), .A2(n12692), .ZN(n8364) );
  XNOR2_X1 U10560 ( .A(n8116), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n10974) );
  NOR2_X1 U10561 ( .A1(n7833), .A2(n10975), .ZN(n8108) );
  NAND2_X1 U10562 ( .A1(n8224), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8114) );
  INV_X1 U10563 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12673) );
  OR2_X1 U10564 ( .A1(n8212), .A2(n12673), .ZN(n8113) );
  INV_X1 U10565 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n15280) );
  OR2_X1 U10566 ( .A1(n8236), .A2(n15280), .ZN(n8112) );
  AND2_X1 U10567 ( .A1(n8109), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8110) );
  NOR2_X1 U10568 ( .A1(n8120), .A2(n8110), .ZN(n12672) );
  OR2_X1 U10569 ( .A1(n8211), .A2(n12672), .ZN(n8111) );
  NAND4_X1 U10570 ( .A1(n8114), .A2(n8113), .A3(n8112), .A4(n8111), .ZN(n12365) );
  NAND2_X1 U10571 ( .A1(n12855), .A2(n12365), .ZN(n8273) );
  INV_X1 U10572 ( .A(n12855), .ZN(n12305) );
  NAND2_X1 U10573 ( .A1(n12305), .A2(n12679), .ZN(n8274) );
  NAND2_X1 U10574 ( .A1(n8273), .A2(n8274), .ZN(n12670) );
  INV_X1 U10575 ( .A(n12670), .ZN(n8511) );
  INV_X1 U10576 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11438) );
  AOI22_X1 U10577 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n11441), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n11438), .ZN(n8127) );
  INV_X1 U10578 ( .A(n8127), .ZN(n8117) );
  NAND2_X1 U10579 ( .A1(n11083), .A2(n6474), .ZN(n8119) );
  INV_X1 U10580 ( .A(SI_21_), .ZN(n11085) );
  NAND2_X1 U10581 ( .A1(n8224), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8125) );
  INV_X1 U10582 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12658) );
  OR2_X1 U10583 ( .A1(n8212), .A2(n12658), .ZN(n8124) );
  INV_X1 U10584 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12795) );
  OR2_X1 U10585 ( .A1(n8236), .A2(n12795), .ZN(n8123) );
  INV_X1 U10586 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n12256) );
  NOR2_X1 U10587 ( .A1(n8120), .A2(n12256), .ZN(n8121) );
  NOR2_X1 U10588 ( .A1(n8134), .A2(n8121), .ZN(n12657) );
  OR2_X1 U10589 ( .A1(n8211), .A2(n12657), .ZN(n8122) );
  NAND2_X1 U10590 ( .A1(n12792), .A2(n12667), .ZN(n8271) );
  INV_X1 U10591 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8130) );
  AOI22_X1 U10592 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(
        P1_DATAO_REG_22__SCAN_IN), .B1(n11717), .B2(n8130), .ZN(n8140) );
  XNOR2_X1 U10593 ( .A(n8141), .B(n8140), .ZN(n11202) );
  NAND2_X1 U10594 ( .A1(n11202), .A2(n6474), .ZN(n8133) );
  INV_X1 U10595 ( .A(SI_22_), .ZN(n8131) );
  OR2_X1 U10596 ( .A1(n7833), .A2(n8131), .ZN(n8132) );
  NAND2_X1 U10597 ( .A1(n8224), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8139) );
  INV_X1 U10598 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12644) );
  OR2_X1 U10599 ( .A1(n8212), .A2(n12644), .ZN(n8138) );
  INV_X1 U10600 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n12319) );
  OR2_X1 U10601 ( .A1(n8134), .A2(n12319), .ZN(n8135) );
  AND2_X1 U10602 ( .A1(n8144), .A2(n8135), .ZN(n12643) );
  OR2_X1 U10603 ( .A1(n8211), .A2(n12643), .ZN(n8137) );
  INV_X1 U10604 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12790) );
  OR2_X1 U10605 ( .A1(n8236), .A2(n12790), .ZN(n8136) );
  NAND4_X1 U10606 ( .A1(n8139), .A2(n8138), .A3(n8137), .A4(n8136), .ZN(n12627) );
  INV_X1 U10607 ( .A(n12627), .ZN(n12656) );
  NAND2_X1 U10608 ( .A1(n12646), .A2(n12656), .ZN(n8375) );
  AND2_X1 U10609 ( .A1(n12849), .A2(n12627), .ZN(n8374) );
  INV_X1 U10610 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11791) );
  AOI22_X1 U10611 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(
        P1_DATAO_REG_23__SCAN_IN), .B1(n11796), .B2(n11791), .ZN(n8150) );
  XNOR2_X1 U10612 ( .A(n8151), .B(n8150), .ZN(n11302) );
  NAND2_X1 U10613 ( .A1(n11302), .A2(n6474), .ZN(n8143) );
  INV_X1 U10614 ( .A(SI_23_), .ZN(n11305) );
  NAND2_X1 U10615 ( .A1(n8224), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8149) );
  INV_X1 U10616 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12631) );
  OR2_X1 U10617 ( .A1(n8212), .A2(n12631), .ZN(n8148) );
  NAND2_X1 U10618 ( .A1(n8144), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8145) );
  AND2_X1 U10619 ( .A1(n8154), .A2(n8145), .ZN(n12630) );
  OR2_X1 U10620 ( .A1(n8211), .A2(n12630), .ZN(n8147) );
  INV_X1 U10621 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n15390) );
  OR2_X1 U10622 ( .A1(n8236), .A2(n15390), .ZN(n8146) );
  NAND4_X1 U10623 ( .A1(n8149), .A2(n8148), .A3(n8147), .A4(n8146), .ZN(n12363) );
  XNOR2_X1 U10624 ( .A(n12633), .B(n12363), .ZN(n12621) );
  NAND2_X1 U10625 ( .A1(n12845), .A2(n12363), .ZN(n8265) );
  XNOR2_X1 U10626 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8161), .ZN(n11822) );
  NAND2_X1 U10627 ( .A1(n11822), .A2(n6474), .ZN(n8153) );
  NAND2_X1 U10628 ( .A1(n8224), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8159) );
  INV_X1 U10629 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12616) );
  OR2_X1 U10630 ( .A1(n7844), .A2(n12616), .ZN(n8158) );
  NAND2_X1 U10631 ( .A1(n8154), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8155) );
  NAND2_X1 U10632 ( .A1(n8167), .A2(n8155), .ZN(n12296) );
  INV_X1 U10633 ( .A(n12296), .ZN(n12615) );
  OR2_X1 U10634 ( .A1(n8211), .A2(n12615), .ZN(n8157) );
  INV_X1 U10635 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12783) );
  OR2_X1 U10636 ( .A1(n8236), .A2(n12783), .ZN(n8156) );
  NAND4_X1 U10637 ( .A1(n8159), .A2(n8158), .A3(n8157), .A4(n8156), .ZN(n12626) );
  NAND2_X1 U10638 ( .A1(n12841), .A2(n12626), .ZN(n8266) );
  INV_X1 U10639 ( .A(n12841), .ZN(n12618) );
  NAND2_X1 U10640 ( .A1(n12618), .A2(n12187), .ZN(n8268) );
  NAND2_X1 U10641 ( .A1(n8266), .A2(n8268), .ZN(n12609) );
  NAND2_X1 U10642 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n8160), .ZN(n8163) );
  INV_X1 U10643 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n14346) );
  INV_X1 U10644 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13593) );
  AOI22_X1 U10645 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .B1(n13593), .B2(n14342), .ZN(n8164) );
  XNOR2_X1 U10646 ( .A(n8175), .B(n8164), .ZN(n12899) );
  NAND2_X1 U10647 ( .A1(n12899), .A2(n6474), .ZN(n8166) );
  INV_X1 U10648 ( .A(SI_25_), .ZN(n12901) );
  NAND2_X1 U10649 ( .A1(n8224), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8173) );
  INV_X1 U10650 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n12601) );
  OR2_X1 U10651 ( .A1(n8212), .A2(n12601), .ZN(n8172) );
  NOR2_X2 U10652 ( .A1(n8167), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8177) );
  AND2_X1 U10653 ( .A1(n8167), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8168) );
  NOR2_X1 U10654 ( .A1(n8177), .A2(n8168), .ZN(n12600) );
  OR2_X1 U10655 ( .A1(n8211), .A2(n12600), .ZN(n8171) );
  INV_X1 U10656 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n8169) );
  OR2_X1 U10657 ( .A1(n8236), .A2(n8169), .ZN(n8170) );
  AND4_X2 U10658 ( .A1(n8173), .A2(n8172), .A3(n8171), .A4(n8170), .ZN(n12614)
         );
  NAND2_X1 U10659 ( .A1(n12776), .A2(n12614), .ZN(n8263) );
  NAND2_X1 U10660 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n13593), .ZN(n8174) );
  INV_X1 U10661 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14337) );
  AOI22_X1 U10662 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n13587), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n14337), .ZN(n8176) );
  XNOR2_X1 U10663 ( .A(n8183), .B(n8176), .ZN(n12896) );
  NAND2_X1 U10664 ( .A1(n8224), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8182) );
  INV_X1 U10665 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12588) );
  OR2_X1 U10666 ( .A1(n8212), .A2(n12588), .ZN(n8181) );
  INV_X1 U10667 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n12342) );
  OR2_X1 U10668 ( .A1(n8177), .A2(n12342), .ZN(n8178) );
  NAND2_X1 U10669 ( .A1(n8177), .A2(n12342), .ZN(n8189) );
  AND2_X1 U10670 ( .A1(n8178), .A2(n8189), .ZN(n12587) );
  OR2_X1 U10671 ( .A1(n8211), .A2(n12587), .ZN(n8180) );
  INV_X1 U10672 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12774) );
  OR2_X1 U10673 ( .A1(n8236), .A2(n12774), .ZN(n8179) );
  NOR2_X1 U10674 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n14337), .ZN(n8184) );
  INV_X1 U10675 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13583) );
  INV_X1 U10676 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14336) );
  AOI22_X1 U10677 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n13583), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n14336), .ZN(n8185) );
  INV_X1 U10678 ( .A(n8185), .ZN(n8186) );
  XNOR2_X1 U10679 ( .A(n8195), .B(n8186), .ZN(n12158) );
  NAND2_X1 U10680 ( .A1(n12158), .A2(n6474), .ZN(n8188) );
  INV_X1 U10681 ( .A(SI_27_), .ZN(n12159) );
  NAND2_X1 U10682 ( .A1(n8224), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8194) );
  INV_X1 U10683 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n12573) );
  OR2_X1 U10684 ( .A1(n8212), .A2(n12573), .ZN(n8193) );
  INV_X1 U10685 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n15259) );
  OR2_X1 U10686 ( .A1(n8236), .A2(n15259), .ZN(n8192) );
  NAND2_X1 U10687 ( .A1(n8189), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8190) );
  NAND2_X1 U10688 ( .A1(n12575), .A2(n8523), .ZN(n8525) );
  NAND2_X1 U10689 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n13583), .ZN(n8196) );
  INV_X1 U10690 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14333) );
  INV_X1 U10691 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n15389) );
  AOI22_X1 U10692 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n14333), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n15389), .ZN(n8197) );
  XNOR2_X1 U10693 ( .A(n8207), .B(n8197), .ZN(n12210) );
  NAND2_X1 U10694 ( .A1(n12210), .A2(n6474), .ZN(n8199) );
  INV_X1 U10695 ( .A(SI_28_), .ZN(n12212) );
  OR2_X1 U10696 ( .A1(n7833), .A2(n12212), .ZN(n8198) );
  NAND2_X1 U10697 ( .A1(n8224), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8206) );
  INV_X1 U10698 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12558) );
  OR2_X1 U10699 ( .A1(n7844), .A2(n12558), .ZN(n8205) );
  AND2_X1 U10700 ( .A1(n8200), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8201) );
  NOR2_X1 U10701 ( .A1(n12549), .A2(n8201), .ZN(n12557) );
  OR2_X1 U10702 ( .A1(n8211), .A2(n12557), .ZN(n8204) );
  INV_X1 U10703 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n8202) );
  OR2_X1 U10704 ( .A1(n8236), .A2(n8202), .ZN(n8203) );
  NAND2_X1 U10705 ( .A1(n12767), .A2(n12226), .ZN(n8259) );
  NAND2_X1 U10706 ( .A1(n8259), .A2(n8525), .ZN(n8394) );
  INV_X1 U10707 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13576) );
  AOI22_X1 U10708 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n13576), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n14330), .ZN(n8220) );
  INV_X1 U10709 ( .A(n8220), .ZN(n8208) );
  NAND2_X1 U10710 ( .A1(n12892), .A2(n6474), .ZN(n8210) );
  INV_X1 U10711 ( .A(SI_29_), .ZN(n12893) );
  OR2_X1 U10712 ( .A1(n7833), .A2(n12893), .ZN(n8209) );
  INV_X1 U10713 ( .A(n12549), .ZN(n12213) );
  INV_X1 U10714 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n15272) );
  OR2_X1 U10715 ( .A1(n8212), .A2(n15272), .ZN(n8218) );
  INV_X1 U10716 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8213) );
  OR2_X1 U10717 ( .A1(n8236), .A2(n8213), .ZN(n8217) );
  INV_X1 U10718 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8214) );
  OR2_X1 U10719 ( .A1(n8215), .A2(n8214), .ZN(n8216) );
  INV_X1 U10720 ( .A(n8403), .ZN(n8230) );
  INV_X1 U10721 ( .A(n8232), .ZN(n8221) );
  INV_X1 U10722 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14328) );
  INV_X1 U10723 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13574) );
  OAI22_X1 U10724 ( .A1(n14328), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n13574), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8231) );
  XNOR2_X1 U10725 ( .A(n8221), .B(n8231), .ZN(n12220) );
  NAND2_X1 U10726 ( .A1(n6474), .A2(n12220), .ZN(n8223) );
  INV_X1 U10727 ( .A(SI_30_), .ZN(n12222) );
  OR2_X1 U10728 ( .A1(n7833), .A2(n12222), .ZN(n8222) );
  NAND2_X1 U10729 ( .A1(n8224), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n8229) );
  INV_X1 U10730 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n8225) );
  OR2_X1 U10731 ( .A1(n8212), .A2(n8225), .ZN(n8228) );
  INV_X1 U10732 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n8226) );
  OR2_X1 U10733 ( .A1(n8236), .A2(n8226), .ZN(n8227) );
  NAND4_X1 U10734 ( .A1(n8240), .A2(n8229), .A3(n8228), .A4(n8227), .ZN(n12552) );
  OAI22_X1 U10735 ( .A1(n9173), .A2(n8230), .B1(n14515), .B2(n12552), .ZN(
        n8245) );
  INV_X1 U10736 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9972) );
  INV_X1 U10737 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14318) );
  AOI22_X1 U10738 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(
        P1_DATAO_REG_31__SCAN_IN), .B1(n9972), .B2(n14318), .ZN(n8233) );
  INV_X1 U10739 ( .A(SI_31_), .ZN(n12886) );
  NOR2_X1 U10740 ( .A1(n7833), .A2(n12886), .ZN(n8234) );
  NAND2_X1 U10741 ( .A1(n14512), .A2(n12552), .ZN(n8399) );
  NAND2_X1 U10742 ( .A1(n8224), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8239) );
  INV_X1 U10743 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n15412) );
  OR2_X1 U10744 ( .A1(n8212), .A2(n15412), .ZN(n8238) );
  INV_X1 U10745 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n8235) );
  OR2_X1 U10746 ( .A1(n8236), .A2(n8235), .ZN(n8237) );
  NAND4_X1 U10747 ( .A1(n8240), .A2(n8239), .A3(n8238), .A4(n8237), .ZN(n12362) );
  OR2_X1 U10748 ( .A1(n12362), .A2(n14515), .ZN(n8241) );
  NAND2_X1 U10749 ( .A1(n12217), .A2(n12205), .ZN(n8402) );
  INV_X1 U10750 ( .A(n14512), .ZN(n8244) );
  INV_X1 U10751 ( .A(n12552), .ZN(n8243) );
  AND2_X1 U10752 ( .A1(n12362), .A2(n14515), .ZN(n8242) );
  OAI22_X1 U10753 ( .A1(n8245), .A2(n8255), .B1(n14512), .B2(n8423), .ZN(n8246) );
  INV_X1 U10754 ( .A(n12531), .ZN(n12545) );
  XNOR2_X1 U10755 ( .A(n8246), .B(n12545), .ZN(n8254) );
  NAND2_X1 U10756 ( .A1(n8251), .A2(n8248), .ZN(n8256) );
  NAND2_X1 U10757 ( .A1(n8256), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8250) );
  INV_X1 U10758 ( .A(n8251), .ZN(n8252) );
  NAND2_X1 U10759 ( .A1(n8252), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8253) );
  NAND2_X1 U10760 ( .A1(n11310), .A2(n9185), .ZN(n8520) );
  NOR2_X1 U10761 ( .A1(n8254), .A2(n8520), .ZN(n8434) );
  NAND2_X1 U10762 ( .A1(n10977), .A2(n12545), .ZN(n9186) );
  INV_X1 U10763 ( .A(n9186), .ZN(n9182) );
  INV_X1 U10764 ( .A(n8255), .ZN(n8401) );
  INV_X1 U10765 ( .A(n8389), .ZN(n8392) );
  AND2_X2 U10766 ( .A1(n8471), .A2(n11310), .ZN(n8307) );
  NAND2_X1 U10767 ( .A1(n8260), .A2(n9184), .ZN(n8391) );
  INV_X1 U10768 ( .A(n8260), .ZN(n8262) );
  MUX2_X1 U10769 ( .A(n8263), .B(n8264), .S(n8307), .Z(n8384) );
  NAND2_X1 U10770 ( .A1(n8266), .A2(n8265), .ZN(n8267) );
  NAND2_X1 U10771 ( .A1(n8267), .A2(n8268), .ZN(n8269) );
  MUX2_X1 U10772 ( .A(n8269), .B(n8268), .S(n8307), .Z(n8382) );
  INV_X1 U10773 ( .A(n12609), .ZN(n12612) );
  INV_X1 U10774 ( .A(n8375), .ZN(n8270) );
  INV_X1 U10775 ( .A(n12637), .ZN(n12640) );
  MUX2_X1 U10776 ( .A(n8272), .B(n8271), .S(n8307), .Z(n8373) );
  MUX2_X1 U10777 ( .A(n8274), .B(n8273), .S(n8307), .Z(n8371) );
  INV_X1 U10778 ( .A(n12696), .ZN(n8275) );
  NAND2_X1 U10779 ( .A1(n12695), .A2(n8275), .ZN(n8276) );
  AND3_X1 U10780 ( .A1(n8276), .A2(n8364), .A3(n8279), .ZN(n8284) );
  INV_X1 U10781 ( .A(n8277), .ZN(n8278) );
  NAND2_X1 U10782 ( .A1(n8279), .A2(n8278), .ZN(n8281) );
  NAND2_X1 U10783 ( .A1(n8281), .A2(n8280), .ZN(n8282) );
  NOR2_X1 U10784 ( .A1(n8365), .A2(n8282), .ZN(n8283) );
  MUX2_X1 U10785 ( .A(n8284), .B(n8283), .S(n8307), .Z(n8368) );
  NAND2_X1 U10786 ( .A1(n15198), .A2(n11084), .ZN(n8285) );
  NAND2_X1 U10787 ( .A1(n15202), .A2(n10694), .ZN(n8409) );
  NAND2_X1 U10788 ( .A1(n8285), .A2(n8409), .ZN(n8287) );
  AND2_X1 U10789 ( .A1(n8406), .A2(n8409), .ZN(n8286) );
  MUX2_X1 U10790 ( .A(n8287), .B(n8286), .S(n8307), .Z(n8288) );
  NAND2_X1 U10791 ( .A1(n8288), .A2(n8407), .ZN(n8290) );
  MUX2_X1 U10792 ( .A(n8407), .B(n8406), .S(n9184), .Z(n8289) );
  NAND3_X1 U10793 ( .A1(n8290), .A2(n15180), .A3(n8289), .ZN(n8294) );
  NAND2_X1 U10794 ( .A1(n8299), .A2(n8291), .ZN(n8292) );
  NAND2_X1 U10795 ( .A1(n8292), .A2(n9184), .ZN(n8293) );
  NAND2_X1 U10796 ( .A1(n8294), .A2(n8293), .ZN(n8298) );
  AOI21_X1 U10797 ( .B1(n8297), .B2(n8295), .A(n9184), .ZN(n8296) );
  AOI21_X1 U10798 ( .B1(n8298), .B2(n8297), .A(n8296), .ZN(n8304) );
  OAI21_X1 U10799 ( .B1(n8299), .B2(n9184), .A(n10837), .ZN(n8303) );
  MUX2_X1 U10800 ( .A(n8301), .B(n8300), .S(n8307), .Z(n8302) );
  OAI211_X1 U10801 ( .C1(n8304), .C2(n8303), .A(n11314), .B(n8302), .ZN(n8312)
         );
  NAND2_X1 U10802 ( .A1(n8314), .A2(n8305), .ZN(n8309) );
  NAND2_X1 U10803 ( .A1(n8313), .A2(n8306), .ZN(n8308) );
  MUX2_X1 U10804 ( .A(n8309), .B(n8308), .S(n9184), .Z(n8310) );
  INV_X1 U10805 ( .A(n8310), .ZN(n8311) );
  NAND2_X1 U10806 ( .A1(n8312), .A2(n8311), .ZN(n8316) );
  MUX2_X1 U10807 ( .A(n8314), .B(n8313), .S(n8307), .Z(n8315) );
  NAND3_X1 U10808 ( .A1(n8316), .A2(n11284), .A3(n8315), .ZN(n8320) );
  MUX2_X1 U10809 ( .A(n8318), .B(n8317), .S(n9184), .Z(n8319) );
  NAND3_X1 U10810 ( .A1(n8320), .A2(n11485), .A3(n8319), .ZN(n8324) );
  XNOR2_X1 U10811 ( .A(n12368), .B(n11709), .ZN(n11705) );
  INV_X1 U10812 ( .A(n11705), .ZN(n8405) );
  MUX2_X1 U10813 ( .A(n8322), .B(n8321), .S(n8307), .Z(n8323) );
  NAND3_X1 U10814 ( .A1(n8324), .A2(n8405), .A3(n8323), .ZN(n8328) );
  OR2_X1 U10815 ( .A1(n11709), .A2(n9184), .ZN(n8326) );
  NAND2_X1 U10816 ( .A1(n11709), .A2(n9184), .ZN(n8325) );
  MUX2_X1 U10817 ( .A(n8326), .B(n8325), .S(n12368), .Z(n8327) );
  NAND2_X1 U10818 ( .A1(n8328), .A2(n8327), .ZN(n8333) );
  INV_X1 U10819 ( .A(n11799), .ZN(n11797) );
  MUX2_X1 U10820 ( .A(n8330), .B(n8329), .S(n9184), .Z(n8331) );
  INV_X1 U10821 ( .A(n14502), .ZN(n14494) );
  NAND2_X1 U10822 ( .A1(n8331), .A2(n14494), .ZN(n8332) );
  AOI21_X1 U10823 ( .B1(n8333), .B2(n11797), .A(n8332), .ZN(n8339) );
  NAND2_X1 U10824 ( .A1(n8341), .A2(n8334), .ZN(n8337) );
  NAND2_X1 U10825 ( .A1(n8340), .A2(n8335), .ZN(n8336) );
  MUX2_X1 U10826 ( .A(n8337), .B(n8336), .S(n8307), .Z(n8338) );
  OR2_X1 U10827 ( .A1(n8339), .A2(n8338), .ZN(n8344) );
  MUX2_X1 U10828 ( .A(n8341), .B(n8340), .S(n9184), .Z(n8343) );
  INV_X1 U10829 ( .A(n8346), .ZN(n8342) );
  NAND2_X1 U10830 ( .A1(n8342), .A2(n8345), .ZN(n14484) );
  AOI21_X1 U10831 ( .B1(n8344), .B2(n8343), .A(n14484), .ZN(n8349) );
  INV_X1 U10832 ( .A(n8345), .ZN(n8347) );
  MUX2_X1 U10833 ( .A(n8347), .B(n8346), .S(n8307), .Z(n8348) );
  OR3_X1 U10834 ( .A1(n8349), .A2(n8348), .A3(n6515), .ZN(n8355) );
  NAND3_X1 U10835 ( .A1(n8355), .A2(n12741), .A3(n8350), .ZN(n8352) );
  NAND3_X1 U10836 ( .A1(n8352), .A2(n8359), .A3(n8351), .ZN(n8353) );
  NAND2_X1 U10837 ( .A1(n8353), .A2(n8357), .ZN(n8362) );
  NAND3_X1 U10838 ( .A1(n8355), .A2(n12741), .A3(n8354), .ZN(n8358) );
  NAND3_X1 U10839 ( .A1(n8358), .A2(n8357), .A3(n8356), .ZN(n8360) );
  NAND2_X1 U10840 ( .A1(n8360), .A2(n8359), .ZN(n8361) );
  MUX2_X1 U10841 ( .A(n8362), .B(n8361), .S(n8307), .Z(n8363) );
  NAND3_X1 U10842 ( .A1(n8363), .A2(n12695), .A3(n12711), .ZN(n8367) );
  MUX2_X1 U10843 ( .A(n8365), .B(n8103), .S(n8307), .Z(n8366) );
  AOI21_X1 U10844 ( .B1(n8368), .B2(n8367), .A(n8366), .ZN(n8369) );
  NAND2_X1 U10845 ( .A1(n8511), .A2(n8369), .ZN(n8370) );
  NAND3_X1 U10846 ( .A1(n12654), .A2(n8371), .A3(n8370), .ZN(n8372) );
  NAND3_X1 U10847 ( .A1(n12640), .A2(n8373), .A3(n8372), .ZN(n8377) );
  MUX2_X1 U10848 ( .A(n8375), .B(n7331), .S(n8307), .Z(n8376) );
  NAND3_X1 U10849 ( .A1(n8377), .A2(n12621), .A3(n8376), .ZN(n8379) );
  INV_X1 U10850 ( .A(n12363), .ZN(n12642) );
  NAND3_X1 U10851 ( .A1(n12633), .A2(n12642), .A3(n8307), .ZN(n8378) );
  NAND2_X1 U10852 ( .A1(n8379), .A2(n8378), .ZN(n8380) );
  NAND2_X1 U10853 ( .A1(n12612), .A2(n8380), .ZN(n8381) );
  NAND3_X1 U10854 ( .A1(n12602), .A2(n8382), .A3(n8381), .ZN(n8383) );
  NAND2_X1 U10855 ( .A1(n8384), .A2(n8383), .ZN(n8385) );
  NAND2_X1 U10856 ( .A1(n12579), .A2(n8385), .ZN(n8387) );
  NAND3_X1 U10857 ( .A1(n12836), .A2(n8307), .A3(n12597), .ZN(n8386) );
  NAND3_X1 U10858 ( .A1(n6753), .A2(n8387), .A3(n8386), .ZN(n8388) );
  OAI21_X1 U10859 ( .B1(n8307), .B2(n8389), .A(n8388), .ZN(n8390) );
  OAI211_X1 U10860 ( .C1(n8392), .C2(n8391), .A(n8527), .B(n8390), .ZN(n8397)
         );
  OAI21_X1 U10861 ( .B1(n8394), .B2(n9184), .A(n8393), .ZN(n8395) );
  NAND2_X1 U10862 ( .A1(n8397), .A2(n8395), .ZN(n8396) );
  OAI211_X1 U10863 ( .C1(n8397), .C2(n8307), .A(n8396), .B(n8403), .ZN(n8400)
         );
  INV_X1 U10864 ( .A(n8423), .ZN(n8398) );
  INV_X1 U10865 ( .A(n8527), .ZN(n12202) );
  AND2_X1 U10866 ( .A1(n12249), .A2(n12692), .ZN(n8509) );
  INV_X1 U10867 ( .A(n12692), .ZN(n12327) );
  NAND2_X1 U10868 ( .A1(n12859), .A2(n12327), .ZN(n8510) );
  INV_X1 U10869 ( .A(n8510), .ZN(n8404) );
  NOR2_X1 U10870 ( .A1(n8509), .A2(n8404), .ZN(n12680) );
  INV_X1 U10871 ( .A(n14484), .ZN(n8415) );
  NAND4_X1 U10872 ( .A1(n8405), .A2(n10738), .A3(n11239), .A4(n11797), .ZN(
        n8412) );
  INV_X1 U10873 ( .A(n8482), .ZN(n8408) );
  NAND3_X1 U10874 ( .A1(n15180), .A2(n8408), .A3(n10837), .ZN(n8411) );
  AND2_X1 U10875 ( .A1(n15198), .A2(n8409), .ZN(n10686) );
  NAND4_X1 U10876 ( .A1(n11284), .A2(n11314), .A3(n11485), .A4(n10686), .ZN(
        n8410) );
  NOR3_X1 U10877 ( .A1(n8412), .A2(n8411), .A3(n8410), .ZN(n8413) );
  NAND4_X1 U10878 ( .A1(n8415), .A2(n14494), .A3(n8414), .A4(n8413), .ZN(n8416) );
  OR2_X1 U10879 ( .A1(n6515), .A2(n8416), .ZN(n8417) );
  NOR4_X1 U10880 ( .A1(n12722), .A2(n12680), .A3(n8418), .A4(n8417), .ZN(n8419) );
  NAND4_X1 U10881 ( .A1(n12654), .A2(n12695), .A3(n12711), .A4(n8419), .ZN(
        n8420) );
  NOR4_X1 U10882 ( .A1(n12609), .A2(n12670), .A3(n12637), .A4(n8420), .ZN(
        n8421) );
  NAND4_X1 U10883 ( .A1(n12602), .A2(n12621), .A3(n12579), .A4(n8421), .ZN(
        n8422) );
  XNOR2_X1 U10884 ( .A(n8425), .B(n12531), .ZN(n8426) );
  NAND2_X1 U10885 ( .A1(n8429), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8428) );
  MUX2_X1 U10886 ( .A(n8428), .B(P3_IR_REG_31__SCAN_IN), .S(n8430), .Z(n8431)
         );
  INV_X1 U10887 ( .A(n10672), .ZN(n8432) );
  NAND2_X1 U10888 ( .A1(n8432), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11303) );
  INV_X1 U10889 ( .A(n11303), .ZN(n8433) );
  INV_X1 U10890 ( .A(n7801), .ZN(n8436) );
  INV_X1 U10891 ( .A(n8444), .ZN(n8439) );
  NAND2_X1 U10892 ( .A1(n8439), .A2(n8438), .ZN(n8446) );
  NAND2_X1 U10893 ( .A1(n8446), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8440) );
  MUX2_X1 U10894 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8440), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8443) );
  INV_X1 U10895 ( .A(n8441), .ZN(n8442) );
  INV_X1 U10896 ( .A(n12904), .ZN(n8449) );
  NAND2_X1 U10897 ( .A1(n8444), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8445) );
  MUX2_X1 U10898 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8445), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8447) );
  INV_X1 U10899 ( .A(n11825), .ZN(n8448) );
  NAND3_X1 U10900 ( .A1(n8458), .A2(n8449), .A3(n8448), .ZN(n10673) );
  INV_X1 U10901 ( .A(n12881), .ZN(n12883) );
  NAND2_X1 U10902 ( .A1(n10615), .A2(n10688), .ZN(n10678) );
  NOR3_X1 U10903 ( .A1(n10678), .A2(n10379), .A3(n8450), .ZN(n8452) );
  OAI21_X1 U10904 ( .B1(n8471), .B2(n11303), .A(P3_B_REG_SCAN_IN), .ZN(n8451)
         );
  OR2_X1 U10905 ( .A1(n8452), .A2(n8451), .ZN(n8453) );
  XNOR2_X1 U10906 ( .A(n11825), .B(P3_B_REG_SCAN_IN), .ZN(n8455) );
  INV_X1 U10907 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8456) );
  INV_X1 U10908 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8457) );
  NAND2_X1 U10909 ( .A1(n10033), .A2(n8457), .ZN(n8460) );
  NAND2_X1 U10910 ( .A1(n7017), .A2(n12904), .ZN(n8459) );
  NAND2_X1 U10911 ( .A1(n12884), .A2(n12882), .ZN(n9181) );
  NOR2_X1 U10912 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_12__SCAN_IN), .ZN(
        n8464) );
  NOR4_X1 U10913 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_14__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n8463) );
  NOR4_X1 U10914 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8462) );
  NOR4_X1 U10915 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8461) );
  NAND4_X1 U10916 ( .A1(n8464), .A2(n8463), .A3(n8462), .A4(n8461), .ZN(n8470)
         );
  NOR4_X1 U10917 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n8468) );
  NOR4_X1 U10918 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_11__SCAN_IN), .ZN(n8467) );
  NOR4_X1 U10919 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8466) );
  NOR4_X1 U10920 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8465) );
  NAND4_X1 U10921 ( .A1(n8468), .A2(n8467), .A3(n8466), .A4(n8465), .ZN(n8469)
         );
  OAI21_X1 U10922 ( .B1(n8470), .B2(n8469), .A(n10033), .ZN(n9178) );
  INV_X1 U10923 ( .A(n9178), .ZN(n8476) );
  NOR2_X1 U10924 ( .A1(n9181), .A2(n8476), .ZN(n10687) );
  NAND2_X1 U10925 ( .A1(n8471), .A2(n12531), .ZN(n8521) );
  NOR2_X1 U10926 ( .A1(n8521), .A2(n8472), .ZN(n10682) );
  NAND2_X1 U10927 ( .A1(n10682), .A2(n10688), .ZN(n8473) );
  NAND2_X1 U10928 ( .A1(n10678), .A2(n8473), .ZN(n8474) );
  NAND2_X1 U10929 ( .A1(n10687), .A2(n8474), .ZN(n8481) );
  INV_X1 U10930 ( .A(n12884), .ZN(n8475) );
  NAND2_X1 U10931 ( .A1(n8475), .A2(n9188), .ZN(n9179) );
  OAI21_X1 U10932 ( .B1(n11200), .B2(n9185), .A(n12531), .ZN(n8477) );
  NAND2_X1 U10933 ( .A1(n8477), .A2(n11084), .ZN(n8479) );
  OAI21_X1 U10934 ( .B1(n9185), .B2(n11310), .A(n11200), .ZN(n8478) );
  NAND2_X1 U10935 ( .A1(n8479), .A2(n8478), .ZN(n10681) );
  NAND3_X1 U10936 ( .A1(n10692), .A2(n10688), .A3(n10681), .ZN(n8480) );
  INV_X1 U10937 ( .A(n12767), .ZN(n8534) );
  NAND2_X1 U10938 ( .A1(n15202), .A2(n11196), .ZN(n10718) );
  NAND2_X1 U10939 ( .A1(n8482), .A2(n10718), .ZN(n8484) );
  OR2_X1 U10940 ( .A1(n12374), .A2(n7814), .ZN(n8483) );
  NAND2_X1 U10941 ( .A1(n8484), .A2(n8483), .ZN(n15178) );
  INV_X1 U10942 ( .A(n10724), .ZN(n15189) );
  OR2_X1 U10943 ( .A1(n15201), .A2(n15189), .ZN(n8486) );
  INV_X1 U10944 ( .A(n10738), .ZN(n8488) );
  NAND2_X1 U10945 ( .A1(n10960), .A2(n6968), .ZN(n8489) );
  INV_X1 U10946 ( .A(n11627), .ZN(n10969) );
  NAND2_X1 U10947 ( .A1(n12373), .A2(n10969), .ZN(n8490) );
  OR2_X1 U10948 ( .A1(n12372), .A2(n6691), .ZN(n8491) );
  INV_X1 U10949 ( .A(n11647), .ZN(n11502) );
  NAND2_X1 U10950 ( .A1(n12371), .A2(n11502), .ZN(n8492) );
  INV_X1 U10951 ( .A(n11634), .ZN(n11606) );
  NAND2_X1 U10952 ( .A1(n12370), .A2(n11606), .ZN(n8493) );
  OR2_X1 U10953 ( .A1(n12369), .A2(n7086), .ZN(n8494) );
  INV_X1 U10954 ( .A(n11709), .ZN(n11692) );
  NAND2_X1 U10955 ( .A1(n12368), .A2(n11692), .ZN(n8495) );
  NAND2_X1 U10956 ( .A1(n11800), .A2(n11799), .ZN(n11798) );
  INV_X1 U10957 ( .A(n11803), .ZN(n11745) );
  NAND2_X1 U10958 ( .A1(n14496), .A2(n11745), .ZN(n8496) );
  OR2_X1 U10959 ( .A1(n12367), .A2(n11873), .ZN(n8497) );
  NAND2_X1 U10960 ( .A1(n14495), .A2(n8497), .ZN(n8499) );
  NAND2_X1 U10961 ( .A1(n12367), .A2(n11873), .ZN(n8498) );
  NAND2_X1 U10962 ( .A1(n8499), .A2(n8498), .ZN(n11894) );
  INV_X1 U10963 ( .A(n14520), .ZN(n11914) );
  NAND2_X1 U10964 ( .A1(n14497), .A2(n11914), .ZN(n8500) );
  OR2_X1 U10965 ( .A1(n14490), .A2(n12755), .ZN(n8502) );
  INV_X1 U10966 ( .A(n12737), .ZN(n14488) );
  OR2_X1 U10967 ( .A1(n12879), .A2(n14488), .ZN(n8503) );
  NAND2_X1 U10968 ( .A1(n12753), .A2(n8503), .ZN(n12736) );
  NAND2_X1 U10969 ( .A1(n12745), .A2(n12726), .ZN(n8504) );
  NAND2_X1 U10970 ( .A1(n12873), .A2(n12754), .ZN(n8505) );
  AND2_X1 U10971 ( .A1(n12729), .A2(n12353), .ZN(n8507) );
  INV_X1 U10972 ( .A(n12695), .ZN(n12689) );
  NAND2_X1 U10973 ( .A1(n12690), .A2(n12689), .ZN(n12688) );
  OR2_X1 U10974 ( .A1(n12699), .A2(n12366), .ZN(n8508) );
  INV_X1 U10975 ( .A(n12667), .ZN(n12364) );
  NAND2_X1 U10976 ( .A1(n12646), .A2(n12627), .ZN(n8514) );
  NAND2_X1 U10977 ( .A1(n12633), .A2(n12363), .ZN(n8515) );
  INV_X1 U10978 ( .A(n12614), .ZN(n12582) );
  NAND2_X1 U10979 ( .A1(n12836), .A2(n8517), .ZN(n8519) );
  NOR2_X1 U10980 ( .A1(n12836), .A2(n8517), .ZN(n8518) );
  OR2_X1 U10981 ( .A1(n8450), .A2(n12506), .ZN(n10359) );
  NAND2_X1 U10982 ( .A1(n10359), .A2(n10356), .ZN(n8522) );
  INV_X1 U10983 ( .A(n8522), .ZN(n10705) );
  OAI22_X1 U10984 ( .A1(n8523), .A2(n15183), .B1(n12205), .B2(n15182), .ZN(
        n8524) );
  INV_X1 U10985 ( .A(n8525), .ZN(n8526) );
  NOR2_X1 U10986 ( .A1(n12564), .A2(n8526), .ZN(n8528) );
  XNOR2_X1 U10987 ( .A(n8528), .B(n8527), .ZN(n12559) );
  INV_X1 U10988 ( .A(n12559), .ZN(n8532) );
  AND2_X1 U10989 ( .A1(n15195), .A2(n9182), .ZN(n8529) );
  NAND2_X1 U10990 ( .A1(n10681), .A2(n8529), .ZN(n8530) );
  OR3_X1 U10991 ( .A1(n11200), .A2(n12531), .A3(n10977), .ZN(n9183) );
  NAND2_X1 U10992 ( .A1(n11200), .A2(n15190), .ZN(n15222) );
  NOR2_X1 U10993 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), 
        .ZN(n8537) );
  NOR2_X1 U10994 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n8536) );
  NOR2_X1 U10995 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n8535) );
  NAND2_X1 U10996 ( .A1(n8560), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8548) );
  NAND2_X1 U10997 ( .A1(n8610), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8555) );
  NAND2_X1 U10998 ( .A1(n9060), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n8554) );
  AND2_X2 U10999 ( .A1(n14325), .A2(n8549), .ZN(n8614) );
  NAND2_X1 U11000 ( .A1(n8614), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8553) );
  NAND2_X1 U11001 ( .A1(n6475), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8552) );
  INV_X1 U11002 ( .A(SI_0_), .ZN(n8556) );
  NOR2_X1 U11003 ( .A1(n9676), .A2(n8556), .ZN(n8558) );
  XNOR2_X1 U11004 ( .A(n8558), .B(n8557), .ZN(n14350) );
  NAND2_X1 U11005 ( .A1(n10342), .A2(n10259), .ZN(n10339) );
  NAND2_X1 U11006 ( .A1(n8610), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8564) );
  INV_X1 U11007 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n8565) );
  INV_X1 U11008 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9929) );
  INV_X1 U11009 ( .A(n8569), .ZN(n8568) );
  NAND2_X1 U11010 ( .A1(n8571), .A2(n8570), .ZN(n8572) );
  NAND2_X1 U11011 ( .A1(n7605), .A2(n8572), .ZN(n9930) );
  XNOR2_X2 U11012 ( .A(n13897), .B(n14844), .ZN(n12117) );
  INV_X1 U11013 ( .A(n13897), .ZN(n10341) );
  NAND2_X1 U11014 ( .A1(n10341), .A2(n14844), .ZN(n11954) );
  NAND2_X1 U11015 ( .A1(n8610), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n8578) );
  NAND2_X1 U11016 ( .A1(n9060), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n8577) );
  NAND2_X1 U11017 ( .A1(n8614), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8576) );
  NAND2_X1 U11018 ( .A1(n8582), .A2(n8581), .ZN(n8583) );
  OR2_X1 U11019 ( .A1(n8727), .A2(n9906), .ZN(n8591) );
  INV_X1 U11020 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9901) );
  NOR2_X1 U11021 ( .A1(n8584), .A2(n8672), .ZN(n8585) );
  MUX2_X1 U11022 ( .A(n8672), .B(n8585), .S(P1_IR_REG_2__SCAN_IN), .Z(n8586)
         );
  INV_X1 U11023 ( .A(n8586), .ZN(n8588) );
  NAND2_X1 U11024 ( .A1(n8588), .A2(n8587), .ZN(n10310) );
  OR2_X1 U11025 ( .A1(n8947), .A2(n10310), .ZN(n8589) );
  NAND2_X1 U11026 ( .A1(n13895), .A2(n14861), .ZN(n11958) );
  NAND2_X2 U11027 ( .A1(n11959), .A2(n11958), .ZN(n14825) );
  NAND2_X1 U11028 ( .A1(n14824), .A2(n14825), .ZN(n8593) );
  NAND2_X1 U11029 ( .A1(n10267), .A2(n14861), .ZN(n8592) );
  NAND2_X1 U11030 ( .A1(n8610), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8598) );
  INV_X1 U11031 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n8612) );
  NAND2_X1 U11032 ( .A1(n8614), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8596) );
  NAND2_X1 U11033 ( .A1(n6475), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8595) );
  NAND2_X1 U11034 ( .A1(n8601), .A2(n8620), .ZN(n9902) );
  NAND2_X1 U11035 ( .A1(n8587), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8602) );
  MUX2_X1 U11036 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8602), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n8604) );
  NAND2_X1 U11037 ( .A1(n8604), .A2(n8603), .ZN(n10087) );
  OR2_X1 U11038 ( .A1(n8947), .A2(n10087), .ZN(n8606) );
  INV_X1 U11039 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9900) );
  OR2_X1 U11040 ( .A1(n12088), .A2(n9900), .ZN(n8605) );
  AND3_X2 U11041 ( .A1(n8607), .A2(n8606), .A3(n8605), .ZN(n14873) );
  INV_X1 U11042 ( .A(n14873), .ZN(n13742) );
  NAND2_X1 U11043 ( .A1(n10801), .A2(n13742), .ZN(n11964) );
  NAND2_X1 U11044 ( .A1(n13894), .A2(n14873), .ZN(n11963) );
  NAND2_X1 U11045 ( .A1(n11964), .A2(n11963), .ZN(n12116) );
  NAND2_X1 U11046 ( .A1(n10855), .A2(n12116), .ZN(n8609) );
  NAND2_X1 U11047 ( .A1(n10801), .A2(n14873), .ZN(n8608) );
  NAND2_X1 U11048 ( .A1(n6475), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8618) );
  NAND2_X1 U11049 ( .A1(n9966), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n8617) );
  INV_X1 U11050 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n8611) );
  NAND2_X1 U11051 ( .A1(n8612), .A2(n8611), .ZN(n8613) );
  NAND2_X1 U11052 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8640) );
  AND2_X1 U11053 ( .A1(n8613), .A2(n8640), .ZN(n10792) );
  NAND2_X1 U11054 ( .A1(n9060), .A2(n10792), .ZN(n8616) );
  NAND2_X1 U11055 ( .A1(n9967), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n8615) );
  NAND2_X1 U11056 ( .A1(n8631), .A2(n8622), .ZN(n9912) );
  OR2_X1 U11057 ( .A1(n9912), .A2(n8727), .ZN(n8628) );
  INV_X2 U11058 ( .A(n12088), .ZN(n8900) );
  NAND2_X1 U11059 ( .A1(n8603), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8623) );
  MUX2_X1 U11060 ( .A(n8623), .B(P1_IR_REG_31__SCAN_IN), .S(n8624), .Z(n8626)
         );
  INV_X1 U11061 ( .A(n8603), .ZN(n8625) );
  NAND2_X1 U11062 ( .A1(n8625), .A2(n8624), .ZN(n8636) );
  NAND2_X1 U11063 ( .A1(n8626), .A2(n8636), .ZN(n10321) );
  INV_X1 U11064 ( .A(n10321), .ZN(n10092) );
  AOI22_X1 U11065 ( .A1(n8900), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n9950), .B2(
        n10092), .ZN(n8627) );
  AND2_X1 U11066 ( .A1(n10929), .A2(n10928), .ZN(n8629) );
  NAND2_X1 U11067 ( .A1(n8632), .A2(SI_5_), .ZN(n8648) );
  OAI21_X1 U11068 ( .B1(n8632), .B2(SI_5_), .A(n8648), .ZN(n8633) );
  INV_X1 U11069 ( .A(n8633), .ZN(n8634) );
  OR2_X1 U11070 ( .A1(n9916), .A2(n8727), .ZN(n8639) );
  NAND2_X1 U11071 ( .A1(n8636), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8637) );
  XNOR2_X1 U11072 ( .A(n8637), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10124) );
  AOI22_X1 U11073 ( .A1(n8900), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9950), .B2(
        n10124), .ZN(n8638) );
  NAND2_X1 U11074 ( .A1(n9966), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8645) );
  NAND2_X1 U11075 ( .A1(n8614), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8644) );
  NOR2_X1 U11076 ( .A1(n8640), .A2(n10899), .ZN(n8659) );
  AND2_X1 U11077 ( .A1(n8640), .A2(n10899), .ZN(n8641) );
  NOR2_X1 U11078 ( .A1(n8659), .A2(n8641), .ZN(n14815) );
  NAND2_X1 U11079 ( .A1(n9060), .A2(n14815), .ZN(n8643) );
  NAND2_X1 U11080 ( .A1(n6475), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n8642) );
  XNOR2_X1 U11081 ( .A(n14813), .B(n13893), .ZN(n12120) );
  INV_X1 U11082 ( .A(n14813), .ZN(n10912) );
  INV_X1 U11083 ( .A(n13893), .ZN(n9087) );
  NAND2_X1 U11084 ( .A1(n10912), .A2(n9087), .ZN(n8647) );
  NAND2_X1 U11085 ( .A1(n10904), .A2(n8647), .ZN(n11088) );
  NAND2_X1 U11086 ( .A1(n8650), .A2(SI_6_), .ZN(n8666) );
  OAI21_X1 U11087 ( .B1(SI_6_), .B2(n8650), .A(n8666), .ZN(n8651) );
  INV_X1 U11088 ( .A(n8651), .ZN(n8652) );
  OR2_X1 U11089 ( .A1(n9927), .A2(n8727), .ZN(n8658) );
  NOR2_X1 U11090 ( .A1(n8842), .A2(n8672), .ZN(n8654) );
  MUX2_X1 U11091 ( .A(n8672), .B(n8654), .S(P1_IR_REG_6__SCAN_IN), .Z(n8656)
         );
  INV_X1 U11092 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8655) );
  AND2_X1 U11093 ( .A1(n8842), .A2(n8655), .ZN(n8690) );
  OR2_X1 U11094 ( .A1(n8656), .A2(n8690), .ZN(n10121) );
  INV_X1 U11095 ( .A(n10121), .ZN(n10137) );
  AOI22_X1 U11096 ( .A1(n8900), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9950), .B2(
        n10137), .ZN(n8657) );
  NAND2_X1 U11097 ( .A1(n6475), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8664) );
  NAND2_X1 U11098 ( .A1(n9966), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n8663) );
  NAND2_X1 U11099 ( .A1(n8659), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8676) );
  OR2_X1 U11100 ( .A1(n8659), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8660) );
  AND2_X1 U11101 ( .A1(n8676), .A2(n8660), .ZN(n11054) );
  NAND2_X1 U11102 ( .A1(n9060), .A2(n11054), .ZN(n8662) );
  NAND2_X1 U11103 ( .A1(n8614), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n8661) );
  NAND4_X1 U11104 ( .A1(n8664), .A2(n8663), .A3(n8662), .A4(n8661), .ZN(n13892) );
  INV_X1 U11105 ( .A(n13892), .ZN(n9090) );
  XNOR2_X1 U11106 ( .A(n11976), .B(n9090), .ZN(n11091) );
  OR2_X1 U11107 ( .A1(n11976), .A2(n13892), .ZN(n8665) );
  MUX2_X1 U11108 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9676), .Z(n8668) );
  NAND2_X1 U11109 ( .A1(n8668), .A2(SI_7_), .ZN(n8683) );
  OAI21_X1 U11110 ( .B1(n8668), .B2(SI_7_), .A(n8683), .ZN(n8669) );
  INV_X1 U11111 ( .A(n8669), .ZN(n8670) );
  OR2_X1 U11112 ( .A1(n9935), .A2(n8727), .ZN(n8675) );
  OR2_X1 U11113 ( .A1(n8690), .A2(n8672), .ZN(n8673) );
  XNOR2_X1 U11114 ( .A(n8673), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10164) );
  AOI22_X1 U11115 ( .A1(n8900), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9950), .B2(
        n10164), .ZN(n8674) );
  NAND2_X1 U11116 ( .A1(n6475), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8681) );
  NAND2_X1 U11117 ( .A1(n9966), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n8680) );
  INV_X1 U11118 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n11119) );
  NAND2_X1 U11119 ( .A1(n8676), .A2(n11119), .ZN(n8677) );
  AND2_X1 U11120 ( .A1(n8694), .A2(n8677), .ZN(n11122) );
  NAND2_X1 U11121 ( .A1(n9060), .A2(n11122), .ZN(n8679) );
  NAND2_X1 U11122 ( .A1(n9967), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n8678) );
  NAND4_X1 U11123 ( .A1(n8681), .A2(n8680), .A3(n8679), .A4(n8678), .ZN(n13891) );
  INV_X1 U11124 ( .A(n13891), .ZN(n11114) );
  OR2_X1 U11125 ( .A1(n11979), .A2(n13891), .ZN(n8682) );
  MUX2_X1 U11126 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9676), .Z(n8685) );
  NAND2_X1 U11127 ( .A1(n8685), .A2(SI_8_), .ZN(n8700) );
  OAI21_X1 U11128 ( .B1(SI_8_), .B2(n8685), .A(n8700), .ZN(n8686) );
  INV_X1 U11129 ( .A(n8686), .ZN(n8687) );
  OR2_X1 U11130 ( .A1(n8688), .A2(n8687), .ZN(n8689) );
  NAND2_X1 U11131 ( .A1(n8690), .A2(n15325), .ZN(n8743) );
  NAND2_X1 U11132 ( .A1(n8743), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8708) );
  XNOR2_X1 U11133 ( .A(n8708), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10287) );
  AOI22_X1 U11134 ( .A1(n8900), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9950), .B2(
        n10287), .ZN(n8691) );
  NAND2_X1 U11135 ( .A1(n9966), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8699) );
  NAND2_X1 U11136 ( .A1(n9967), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8698) );
  INV_X1 U11137 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8693) );
  NAND2_X1 U11138 ( .A1(n8694), .A2(n8693), .ZN(n8695) );
  NAND2_X1 U11139 ( .A1(n8715), .A2(n8695), .ZN(n11525) );
  INV_X1 U11140 ( .A(n11525), .ZN(n10875) );
  NAND2_X1 U11141 ( .A1(n9060), .A2(n10875), .ZN(n8697) );
  NAND2_X1 U11142 ( .A1(n6475), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8696) );
  NAND4_X1 U11143 ( .A1(n8699), .A2(n8698), .A3(n8697), .A4(n8696), .ZN(n13890) );
  INV_X1 U11144 ( .A(n13890), .ZN(n9093) );
  MUX2_X1 U11145 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9676), .Z(n8702) );
  NAND2_X1 U11146 ( .A1(n8702), .A2(SI_9_), .ZN(n8721) );
  OAI21_X1 U11147 ( .B1(SI_9_), .B2(n8702), .A(n8721), .ZN(n8703) );
  INV_X1 U11148 ( .A(n8703), .ZN(n8704) );
  NAND2_X1 U11149 ( .A1(n8708), .A2(n8707), .ZN(n8709) );
  NAND2_X1 U11150 ( .A1(n8709), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8710) );
  NAND2_X1 U11151 ( .A1(n8710), .A2(n8741), .ZN(n8728) );
  OR2_X1 U11152 ( .A1(n8710), .A2(n8741), .ZN(n8711) );
  AOI22_X1 U11153 ( .A1(n8900), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9950), .B2(
        n10474), .ZN(n8712) );
  NAND2_X1 U11154 ( .A1(n6475), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8719) );
  NAND2_X1 U11155 ( .A1(n9966), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n8718) );
  INV_X1 U11156 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8714) );
  NOR2_X1 U11157 ( .A1(n8750), .A2(n7765), .ZN(n14794) );
  NAND2_X1 U11158 ( .A1(n9060), .A2(n14794), .ZN(n8717) );
  NAND2_X1 U11159 ( .A1(n9967), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8716) );
  NAND4_X1 U11160 ( .A1(n8719), .A2(n8718), .A3(n8717), .A4(n8716), .ZN(n13889) );
  INV_X1 U11161 ( .A(n13889), .ZN(n11545) );
  NAND2_X1 U11162 ( .A1(n11420), .A2(n12126), .ZN(n11419) );
  OR2_X1 U11163 ( .A1(n11991), .A2(n13889), .ZN(n8720) );
  MUX2_X1 U11164 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9676), .Z(n8723) );
  NAND2_X1 U11165 ( .A1(n8723), .A2(SI_10_), .ZN(n8738) );
  OAI21_X1 U11166 ( .B1(n8723), .B2(SI_10_), .A(n8738), .ZN(n8724) );
  INV_X1 U11167 ( .A(n8724), .ZN(n8725) );
  OR2_X1 U11168 ( .A1(n9961), .A2(n8727), .ZN(n8731) );
  NAND2_X1 U11169 ( .A1(n8728), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8729) );
  XNOR2_X1 U11170 ( .A(n8729), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11033) );
  AOI22_X1 U11171 ( .A1(n8900), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n9950), 
        .B2(n11033), .ZN(n8730) );
  NAND2_X1 U11172 ( .A1(n6475), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8736) );
  NAND2_X1 U11173 ( .A1(n9966), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n8735) );
  INV_X1 U11174 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8732) );
  XNOR2_X1 U11175 ( .A(n8750), .B(n8732), .ZN(n14784) );
  NAND2_X1 U11176 ( .A1(n9060), .A2(n14784), .ZN(n8734) );
  NAND2_X1 U11177 ( .A1(n8614), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8733) );
  NAND4_X1 U11178 ( .A1(n8736), .A2(n8735), .A3(n8734), .A4(n8733), .ZN(n13888) );
  INV_X1 U11179 ( .A(n13888), .ZN(n11778) );
  XNOR2_X1 U11180 ( .A(n11995), .B(n11778), .ZN(n11371) );
  NAND2_X1 U11181 ( .A1(n11372), .A2(n11371), .ZN(n11370) );
  OR2_X1 U11182 ( .A1(n11995), .A2(n13888), .ZN(n8737) );
  MUX2_X1 U11183 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n9676), .Z(n8757) );
  XNOR2_X1 U11184 ( .A(n8757), .B(SI_11_), .ZN(n8760) );
  NAND2_X1 U11185 ( .A1(n9973), .A2(n12087), .ZN(n8746) );
  INV_X1 U11186 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n8740) );
  NAND2_X1 U11187 ( .A1(n8741), .A2(n8740), .ZN(n8742) );
  NAND2_X1 U11188 ( .A1(n8818), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8744) );
  XNOR2_X1 U11189 ( .A(n8744), .B(P1_IR_REG_11__SCAN_IN), .ZN(n14680) );
  AOI22_X1 U11190 ( .A1(n8900), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9950), 
        .B2(n14680), .ZN(n8745) );
  NAND2_X1 U11191 ( .A1(n9966), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U11192 ( .A1(n8750), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8748) );
  INV_X1 U11193 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8747) );
  NAND2_X1 U11194 ( .A1(n8748), .A2(n8747), .ZN(n8751) );
  AND2_X1 U11195 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n8749) );
  NAND2_X1 U11196 ( .A1(n8750), .A2(n8749), .ZN(n8765) );
  NAND2_X1 U11197 ( .A1(n8751), .A2(n8765), .ZN(n14617) );
  INV_X1 U11198 ( .A(n14617), .ZN(n14632) );
  NAND2_X1 U11199 ( .A1(n9060), .A2(n14632), .ZN(n8754) );
  NAND2_X1 U11200 ( .A1(n9967), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8753) );
  NAND2_X1 U11201 ( .A1(n6475), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8752) );
  NAND4_X1 U11202 ( .A1(n8755), .A2(n8754), .A3(n8753), .A4(n8752), .ZN(n13887) );
  INV_X1 U11203 ( .A(n13887), .ZN(n13614) );
  XNOR2_X1 U11204 ( .A(n14630), .B(n13614), .ZN(n11560) );
  NAND2_X1 U11205 ( .A1(n11555), .A2(n11560), .ZN(n11554) );
  OR2_X1 U11206 ( .A1(n14630), .A2(n13887), .ZN(n8756) );
  INV_X1 U11207 ( .A(n8757), .ZN(n8758) );
  NAND2_X1 U11208 ( .A1(n8758), .A2(n9919), .ZN(n8759) );
  MUX2_X1 U11209 ( .A(n7533), .B(n10102), .S(n9676), .Z(n8774) );
  XNOR2_X1 U11210 ( .A(n8774), .B(SI_12_), .ZN(n8772) );
  XNOR2_X1 U11211 ( .A(n8773), .B(n8772), .ZN(n10073) );
  NAND2_X1 U11212 ( .A1(n10073), .A2(n12087), .ZN(n8763) );
  OAI21_X1 U11213 ( .B1(n8818), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8777) );
  XNOR2_X1 U11214 ( .A(n8777), .B(P1_IR_REG_12__SCAN_IN), .ZN(n13913) );
  AOI22_X1 U11215 ( .A1(n8900), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n9950), 
        .B2(n13913), .ZN(n8762) );
  NAND2_X1 U11216 ( .A1(n6475), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8770) );
  NAND2_X1 U11217 ( .A1(n9966), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n8769) );
  NAND2_X1 U11218 ( .A1(n8765), .A2(n8764), .ZN(n8766) );
  AND2_X1 U11219 ( .A1(n8785), .A2(n8766), .ZN(n13782) );
  NAND2_X1 U11220 ( .A1(n9060), .A2(n13782), .ZN(n8768) );
  NAND2_X1 U11221 ( .A1(n9967), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8767) );
  NAND4_X1 U11222 ( .A1(n8770), .A2(n8769), .A3(n8768), .A4(n8767), .ZN(n13886) );
  INV_X1 U11223 ( .A(n13886), .ZN(n13609) );
  XNOR2_X1 U11224 ( .A(n13791), .B(n13609), .ZN(n11448) );
  OR2_X1 U11225 ( .A1(n13791), .A2(n13886), .ZN(n8771) );
  NAND2_X1 U11226 ( .A1(n8774), .A2(n9933), .ZN(n8775) );
  MUX2_X1 U11227 ( .A(n10215), .B(n10233), .S(n9676), .Z(n8794) );
  XNOR2_X1 U11228 ( .A(n8794), .B(SI_13_), .ZN(n8792) );
  XNOR2_X1 U11229 ( .A(n8793), .B(n8792), .ZN(n10213) );
  NAND2_X1 U11230 ( .A1(n10213), .A2(n12087), .ZN(n8783) );
  INV_X1 U11231 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8776) );
  NAND2_X1 U11232 ( .A1(n8777), .A2(n8776), .ZN(n8778) );
  NAND2_X1 U11233 ( .A1(n8778), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8780) );
  INV_X1 U11234 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8779) );
  NAND2_X1 U11235 ( .A1(n8780), .A2(n8779), .ZN(n8795) );
  OR2_X1 U11236 ( .A1(n8780), .A2(n8779), .ZN(n8781) );
  AOI22_X1 U11237 ( .A1(n8900), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n9950), 
        .B2(n14699), .ZN(n8782) );
  NAND2_X1 U11238 ( .A1(n9966), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8790) );
  AND2_X1 U11239 ( .A1(n8785), .A2(n8784), .ZN(n8786) );
  NOR2_X1 U11240 ( .A1(n8799), .A2(n8786), .ZN(n13830) );
  NAND2_X1 U11241 ( .A1(n9060), .A2(n13830), .ZN(n8789) );
  NAND2_X1 U11242 ( .A1(n9967), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8788) );
  NAND2_X1 U11243 ( .A1(n8594), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8787) );
  NAND4_X1 U11244 ( .A1(n8790), .A2(n8789), .A3(n8788), .A4(n8787), .ZN(n13885) );
  INV_X1 U11245 ( .A(n13885), .ZN(n13606) );
  XNOR2_X1 U11246 ( .A(n13837), .B(n13606), .ZN(n12132) );
  NAND2_X1 U11247 ( .A1(n11471), .A2(n12132), .ZN(n11470) );
  OR2_X1 U11248 ( .A1(n13837), .A2(n13885), .ZN(n8791) );
  INV_X1 U11249 ( .A(SI_14_), .ZN(n9948) );
  MUX2_X1 U11250 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n9676), .Z(n8835) );
  NAND2_X1 U11251 ( .A1(n10423), .A2(n12087), .ZN(n8798) );
  NAND2_X1 U11252 ( .A1(n8795), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8796) );
  AOI22_X1 U11253 ( .A1(n14708), .A2(n9950), .B1(n8900), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8797) );
  NAND2_X1 U11254 ( .A1(n9966), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8805) );
  NOR2_X1 U11255 ( .A1(n8799), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8800) );
  OR2_X1 U11256 ( .A1(n8823), .A2(n8800), .ZN(n14601) );
  INV_X1 U11257 ( .A(n14601), .ZN(n8801) );
  NAND2_X1 U11258 ( .A1(n9060), .A2(n8801), .ZN(n8804) );
  NAND2_X1 U11259 ( .A1(n9967), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8803) );
  NAND2_X1 U11260 ( .A1(n6475), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8802) );
  NAND4_X1 U11261 ( .A1(n8805), .A2(n8804), .A3(n8803), .A4(n8802), .ZN(n13884) );
  INV_X1 U11262 ( .A(n13884), .ZN(n8806) );
  NAND2_X1 U11263 ( .A1(n14597), .A2(n8806), .ZN(n12019) );
  INV_X1 U11264 ( .A(n12133), .ZN(n8807) );
  NAND2_X1 U11265 ( .A1(n14597), .A2(n13884), .ZN(n8809) );
  INV_X1 U11266 ( .A(n8834), .ZN(n8810) );
  OAI22_X1 U11267 ( .A1(n8811), .A2(n8835), .B1(n8810), .B2(SI_14_), .ZN(n8813) );
  MUX2_X1 U11268 ( .A(n7095), .B(n10497), .S(n9676), .Z(n8836) );
  XNOR2_X1 U11269 ( .A(n8836), .B(SI_15_), .ZN(n8812) );
  XNOR2_X1 U11270 ( .A(n8813), .B(n8812), .ZN(n10496) );
  NAND2_X1 U11271 ( .A1(n10496), .A2(n12087), .ZN(n8822) );
  NAND3_X1 U11272 ( .A1(n8816), .A2(n8815), .A3(n8814), .ZN(n8817) );
  OAI21_X1 U11273 ( .B1(n8818), .B2(n8817), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8820) );
  XNOR2_X1 U11274 ( .A(n8820), .B(n8819), .ZN(n13917) );
  INV_X1 U11275 ( .A(n13917), .ZN(n14724) );
  AOI22_X1 U11276 ( .A1(n8900), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9950), 
        .B2(n14724), .ZN(n8821) );
  NAND2_X1 U11277 ( .A1(n9966), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n8829) );
  OR2_X1 U11278 ( .A1(n8823), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8824) );
  NAND2_X1 U11279 ( .A1(n8849), .A2(n8824), .ZN(n14628) );
  INV_X1 U11280 ( .A(n14628), .ZN(n8825) );
  NAND2_X1 U11281 ( .A1(n9060), .A2(n8825), .ZN(n8828) );
  NAND2_X1 U11282 ( .A1(n9967), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8827) );
  NAND2_X1 U11283 ( .A1(n8594), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n8826) );
  NAND4_X1 U11284 ( .A1(n8829), .A2(n8828), .A3(n8827), .A4(n8826), .ZN(n14151) );
  INV_X1 U11285 ( .A(n14151), .ZN(n8830) );
  NAND2_X1 U11286 ( .A1(n14622), .A2(n8830), .ZN(n12020) );
  INV_X1 U11287 ( .A(n8836), .ZN(n8832) );
  NAND2_X1 U11288 ( .A1(n8832), .A2(SI_15_), .ZN(n8837) );
  NAND2_X1 U11289 ( .A1(n8835), .A2(SI_14_), .ZN(n8833) );
  NOR2_X1 U11290 ( .A1(n8835), .A2(SI_14_), .ZN(n8838) );
  AOI22_X1 U11291 ( .A1(n8838), .A2(n8837), .B1(n15386), .B2(n8836), .ZN(n8839) );
  MUX2_X1 U11292 ( .A(n10446), .B(n10464), .S(n9676), .Z(n8858) );
  XNOR2_X1 U11293 ( .A(n8858), .B(SI_16_), .ZN(n8856) );
  XNOR2_X1 U11294 ( .A(n8857), .B(n8856), .ZN(n10445) );
  NAND2_X1 U11295 ( .A1(n10445), .A2(n12087), .ZN(n8847) );
  NAND2_X1 U11296 ( .A1(n6648), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8843) );
  MUX2_X1 U11297 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8843), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n8845) );
  NAND2_X1 U11298 ( .A1(n8845), .A2(n8877), .ZN(n14744) );
  INV_X1 U11299 ( .A(n14744), .ZN(n13919) );
  AOI22_X1 U11300 ( .A1(n8900), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9950), 
        .B2(n13919), .ZN(n8846) );
  INV_X1 U11301 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8848) );
  NAND2_X1 U11302 ( .A1(n8849), .A2(n8848), .ZN(n8850) );
  NAND2_X1 U11303 ( .A1(n8866), .A2(n8850), .ZN(n14608) );
  INV_X1 U11304 ( .A(n14608), .ZN(n14154) );
  NAND2_X1 U11305 ( .A1(n9060), .A2(n14154), .ZN(n8854) );
  NAND2_X1 U11306 ( .A1(n8614), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8853) );
  NAND2_X1 U11307 ( .A1(n6475), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8852) );
  NAND2_X1 U11308 ( .A1(n9966), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8851) );
  NAND4_X1 U11309 ( .A1(n8854), .A2(n8853), .A3(n8852), .A4(n8851), .ZN(n13883) );
  NAND2_X1 U11310 ( .A1(n14604), .A2(n13883), .ZN(n12021) );
  OR2_X1 U11311 ( .A1(n14604), .A2(n13883), .ZN(n8855) );
  NAND2_X1 U11312 ( .A1(n8858), .A2(n10071), .ZN(n8859) );
  MUX2_X1 U11313 ( .A(n7093), .B(n10466), .S(n9676), .Z(n8872) );
  XNOR2_X1 U11314 ( .A(n8872), .B(SI_17_), .ZN(n8861) );
  NAND2_X1 U11315 ( .A1(n8877), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8862) );
  XNOR2_X1 U11316 ( .A(n8862), .B(P1_IR_REG_17__SCAN_IN), .ZN(n13922) );
  AOI22_X1 U11317 ( .A1(n8900), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9950), 
        .B2(n13922), .ZN(n8863) );
  INV_X1 U11318 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8865) );
  AND2_X1 U11319 ( .A1(n8866), .A2(n8865), .ZN(n8867) );
  OR2_X1 U11320 ( .A1(n8867), .A2(n8882), .ZN(n14136) );
  NAND2_X1 U11321 ( .A1(n6475), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8869) );
  NAND2_X1 U11322 ( .A1(n9966), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8868) );
  AND2_X1 U11323 ( .A1(n8869), .A2(n8868), .ZN(n8871) );
  NAND2_X1 U11324 ( .A1(n8614), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n8870) );
  OAI211_X1 U11325 ( .C1(n8915), .C2(n14136), .A(n8871), .B(n8870), .ZN(n14150) );
  NAND2_X1 U11326 ( .A1(n14264), .A2(n14150), .ZN(n12113) );
  NOR2_X1 U11327 ( .A1(n8875), .A2(SI_17_), .ZN(n8873) );
  NAND2_X1 U11328 ( .A1(n8875), .A2(SI_17_), .ZN(n8876) );
  MUX2_X1 U11329 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9676), .Z(n8888) );
  XNOR2_X1 U11330 ( .A(n8889), .B(n8888), .ZN(n10990) );
  NAND2_X1 U11331 ( .A1(n10990), .A2(n12087), .ZN(n8881) );
  NAND2_X1 U11332 ( .A1(n8878), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8879) );
  XNOR2_X1 U11333 ( .A(n8879), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14777) );
  AOI22_X1 U11334 ( .A1(n8900), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9950), 
        .B2(n14777), .ZN(n8880) );
  NOR2_X1 U11335 ( .A1(n8882), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8883) );
  OR2_X1 U11336 ( .A1(n8903), .A2(n8883), .ZN(n14124) );
  AOI22_X1 U11337 ( .A1(n6475), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n9966), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n8885) );
  NAND2_X1 U11338 ( .A1(n8614), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8884) );
  OAI211_X1 U11339 ( .C1(n14124), .C2(n8915), .A(n8885), .B(n8884), .ZN(n13882) );
  AND2_X1 U11340 ( .A1(n14257), .A2(n13882), .ZN(n8887) );
  OR2_X1 U11341 ( .A1(n14257), .A2(n13882), .ZN(n8886) );
  NAND2_X1 U11342 ( .A1(n8891), .A2(n8890), .ZN(n8896) );
  MUX2_X1 U11343 ( .A(n7005), .B(n11205), .S(n9676), .Z(n8892) );
  NAND2_X1 U11344 ( .A1(n8892), .A2(n10426), .ZN(n8909) );
  INV_X1 U11345 ( .A(n8892), .ZN(n8893) );
  NAND2_X1 U11346 ( .A1(n8893), .A2(SI_19_), .ZN(n8894) );
  OR2_X1 U11347 ( .A1(n8896), .A2(n8895), .ZN(n8897) );
  NAND2_X1 U11348 ( .A1(n8910), .A2(n8897), .ZN(n11204) );
  NAND2_X1 U11349 ( .A1(n11204), .A2(n12087), .ZN(n8902) );
  AOI22_X1 U11350 ( .A1(n8900), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9950), 
        .B2(n13930), .ZN(n8901) );
  NAND2_X1 U11351 ( .A1(n8903), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8913) );
  OR2_X1 U11352 ( .A1(n8903), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8904) );
  NAND2_X1 U11353 ( .A1(n8913), .A2(n8904), .ZN(n14105) );
  AOI22_X1 U11354 ( .A1(n8594), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n9966), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n8906) );
  NAND2_X1 U11355 ( .A1(n8614), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8905) );
  OAI211_X1 U11356 ( .C1(n14105), .C2(n8915), .A(n8906), .B(n8905), .ZN(n13881) );
  INV_X1 U11357 ( .A(n13881), .ZN(n8907) );
  OR2_X1 U11358 ( .A1(n14251), .A2(n8907), .ZN(n12040) );
  NAND2_X1 U11359 ( .A1(n14251), .A2(n8907), .ZN(n12039) );
  NAND2_X1 U11360 ( .A1(n12040), .A2(n12039), .ZN(n12137) );
  OR2_X1 U11361 ( .A1(n14251), .A2(n13881), .ZN(n8908) );
  XNOR2_X1 U11362 ( .A(n8945), .B(SI_20_), .ZN(n8924) );
  MUX2_X1 U11363 ( .A(n11369), .B(n11327), .S(n9676), .Z(n8940) );
  XNOR2_X1 U11364 ( .A(n8924), .B(n8940), .ZN(n11326) );
  NAND2_X1 U11365 ( .A1(n11326), .A2(n12087), .ZN(n8912) );
  OR2_X1 U11366 ( .A1(n12088), .A2(n11369), .ZN(n8911) );
  INV_X1 U11367 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13826) );
  NAND2_X1 U11368 ( .A1(n8913), .A2(n13826), .ZN(n8914) );
  INV_X1 U11369 ( .A(n8931), .ZN(n8932) );
  NAND2_X1 U11370 ( .A1(n8914), .A2(n8932), .ZN(n13824) );
  OR2_X1 U11371 ( .A1(n13824), .A2(n8915), .ZN(n8921) );
  INV_X1 U11372 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n14246) );
  NAND2_X1 U11373 ( .A1(n8614), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8917) );
  NAND2_X1 U11374 ( .A1(n9966), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8916) );
  OAI211_X1 U11375 ( .C1(n8918), .C2(n14246), .A(n8917), .B(n8916), .ZN(n8919)
         );
  INV_X1 U11376 ( .A(n8919), .ZN(n8920) );
  NAND2_X1 U11377 ( .A1(n8921), .A2(n8920), .ZN(n13880) );
  XNOR2_X1 U11378 ( .A(n14240), .B(n13880), .ZN(n14096) );
  NAND2_X1 U11379 ( .A1(n14240), .A2(n13880), .ZN(n8923) );
  INV_X1 U11380 ( .A(n8940), .ZN(n8939) );
  NAND2_X1 U11381 ( .A1(n8924), .A2(n8939), .ZN(n8926) );
  OR2_X1 U11382 ( .A1(n8945), .A2(n10975), .ZN(n8925) );
  NAND2_X1 U11383 ( .A1(n8926), .A2(n8925), .ZN(n8928) );
  MUX2_X1 U11384 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9676), .Z(n8941) );
  XNOR2_X1 U11385 ( .A(n8941), .B(SI_21_), .ZN(n8927) );
  NAND2_X1 U11386 ( .A1(n11437), .A2(n12087), .ZN(n8930) );
  OR2_X1 U11387 ( .A1(n12088), .A2(n11438), .ZN(n8929) );
  NAND2_X1 U11388 ( .A1(n6475), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8936) );
  NAND2_X1 U11389 ( .A1(n9966), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8935) );
  INV_X1 U11390 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13777) );
  NAND2_X1 U11391 ( .A1(n8931), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8949) );
  INV_X1 U11392 ( .A(n8949), .ZN(n8948) );
  AOI21_X1 U11393 ( .B1(n13777), .B2(n8932), .A(n8948), .ZN(n14077) );
  NAND2_X1 U11394 ( .A1(n9060), .A2(n14077), .ZN(n8934) );
  NAND2_X1 U11395 ( .A1(n8614), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8933) );
  NAND4_X1 U11396 ( .A1(n8936), .A2(n8935), .A3(n8934), .A4(n8933), .ZN(n13879) );
  XNOR2_X1 U11397 ( .A(n14076), .B(n13879), .ZN(n14073) );
  OR2_X1 U11398 ( .A1(n14076), .A2(n13879), .ZN(n8938) );
  NOR2_X1 U11399 ( .A1(n8940), .A2(n10975), .ZN(n8942) );
  AOI22_X1 U11400 ( .A1(n8942), .A2(n7764), .B1(n8941), .B2(SI_21_), .ZN(n8943) );
  OR2_X1 U11401 ( .A1(n9598), .A2(n9676), .ZN(n8946) );
  XNOR2_X1 U11402 ( .A(n8946), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14349) );
  NAND2_X1 U11403 ( .A1(n14349), .A2(n8947), .ZN(n14065) );
  NAND2_X1 U11404 ( .A1(n6475), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8953) );
  NAND2_X1 U11405 ( .A1(n9966), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8952) );
  INV_X1 U11406 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13845) );
  NAND2_X1 U11407 ( .A1(n8948), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8961) );
  AOI21_X1 U11408 ( .B1(n13845), .B2(n8949), .A(n8960), .ZN(n14063) );
  NAND2_X1 U11409 ( .A1(n9060), .A2(n14063), .ZN(n8951) );
  NAND2_X1 U11410 ( .A1(n8614), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8950) );
  XNOR2_X1 U11411 ( .A(n14065), .B(n13878), .ZN(n9109) );
  NAND2_X1 U11412 ( .A1(n14067), .A2(n9109), .ZN(n8955) );
  NAND2_X1 U11413 ( .A1(n14065), .A2(n13774), .ZN(n8954) );
  MUX2_X1 U11414 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9676), .Z(n9597) );
  NAND2_X1 U11415 ( .A1(n8956), .A2(SI_22_), .ZN(n8957) );
  MUX2_X1 U11416 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9676), .Z(n8972) );
  XNOR2_X1 U11417 ( .A(n8972), .B(SI_23_), .ZN(n8969) );
  XNOR2_X1 U11418 ( .A(n8971), .B(n8969), .ZN(n11793) );
  NAND2_X1 U11419 ( .A1(n11793), .A2(n12087), .ZN(n8959) );
  OR2_X1 U11420 ( .A1(n12088), .A2(n11791), .ZN(n8958) );
  NAND2_X1 U11421 ( .A1(n6475), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8966) );
  NAND2_X1 U11422 ( .A1(n9966), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8965) );
  INV_X1 U11423 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8962) );
  NAND2_X1 U11424 ( .A1(n8960), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8978) );
  INV_X1 U11425 ( .A(n8978), .ZN(n8980) );
  AOI21_X1 U11426 ( .B1(n8962), .B2(n8961), .A(n8980), .ZN(n14049) );
  NAND2_X1 U11427 ( .A1(n9060), .A2(n14049), .ZN(n8964) );
  NAND2_X1 U11428 ( .A1(n9967), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8963) );
  NAND4_X1 U11429 ( .A1(n8966), .A2(n8965), .A3(n8964), .A4(n8963), .ZN(n13877) );
  NOR2_X1 U11430 ( .A1(n14221), .A2(n13877), .ZN(n8968) );
  NAND2_X1 U11431 ( .A1(n14221), .A2(n13877), .ZN(n8967) );
  INV_X1 U11432 ( .A(n8969), .ZN(n8970) );
  NAND2_X1 U11433 ( .A1(n8972), .A2(SI_23_), .ZN(n8973) );
  INV_X1 U11434 ( .A(n8987), .ZN(n8975) );
  MUX2_X1 U11435 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9676), .Z(n8986) );
  NAND2_X1 U11436 ( .A1(n13594), .A2(n12087), .ZN(n8977) );
  OR2_X1 U11437 ( .A1(n12088), .A2(n14346), .ZN(n8976) );
  NAND2_X1 U11438 ( .A1(n9966), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8985) );
  NAND2_X1 U11439 ( .A1(n9967), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8984) );
  INV_X1 U11440 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8979) );
  NAND2_X1 U11441 ( .A1(n8979), .A2(n8978), .ZN(n8981) );
  NAND2_X1 U11442 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n8980), .ZN(n8997) );
  AND2_X1 U11443 ( .A1(n8981), .A2(n8997), .ZN(n14037) );
  NAND2_X1 U11444 ( .A1(n9060), .A2(n14037), .ZN(n8983) );
  NAND2_X1 U11445 ( .A1(n8594), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8982) );
  NAND4_X1 U11446 ( .A1(n8985), .A2(n8984), .A3(n8983), .A4(n8982), .ZN(n13876) );
  XNOR2_X1 U11447 ( .A(n14211), .B(n13876), .ZN(n14030) );
  NAND2_X1 U11448 ( .A1(n8988), .A2(SI_24_), .ZN(n8989) );
  MUX2_X1 U11449 ( .A(n14342), .B(n13593), .S(n9676), .Z(n8990) );
  NAND2_X1 U11450 ( .A1(n8990), .A2(n12901), .ZN(n9006) );
  INV_X1 U11451 ( .A(n8990), .ZN(n8991) );
  NAND2_X1 U11452 ( .A1(n8991), .A2(SI_25_), .ZN(n8992) );
  NAND2_X1 U11453 ( .A1(n9006), .A2(n8992), .ZN(n9004) );
  NAND2_X1 U11454 ( .A1(n13590), .A2(n12087), .ZN(n8994) );
  OR2_X1 U11455 ( .A1(n12088), .A2(n14342), .ZN(n8993) );
  NAND2_X2 U11456 ( .A1(n8994), .A2(n8993), .ZN(n14201) );
  NAND2_X1 U11457 ( .A1(n8594), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n9002) );
  NAND2_X1 U11458 ( .A1(n9966), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9001) );
  INV_X1 U11459 ( .A(n8997), .ZN(n8995) );
  NAND2_X1 U11460 ( .A1(n8995), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9012) );
  INV_X1 U11461 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8996) );
  NAND2_X1 U11462 ( .A1(n8997), .A2(n8996), .ZN(n8998) );
  AND2_X1 U11463 ( .A1(n9012), .A2(n8998), .ZN(n13795) );
  NAND2_X1 U11464 ( .A1(n9060), .A2(n13795), .ZN(n9000) );
  NAND2_X1 U11465 ( .A1(n9967), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8999) );
  NAND4_X1 U11466 ( .A1(n9002), .A2(n9001), .A3(n9000), .A4(n8999), .ZN(n13875) );
  INV_X1 U11467 ( .A(n13875), .ZN(n9114) );
  XNOR2_X1 U11468 ( .A(n14201), .B(n9114), .ZN(n14020) );
  NAND2_X1 U11469 ( .A1(n14201), .A2(n13875), .ZN(n9003) );
  MUX2_X1 U11470 ( .A(n14337), .B(n13587), .S(n9676), .Z(n9022) );
  XNOR2_X1 U11471 ( .A(n9022), .B(SI_26_), .ZN(n9007) );
  XNOR2_X1 U11472 ( .A(n9023), .B(n9007), .ZN(n13585) );
  NAND2_X1 U11473 ( .A1(n13585), .A2(n12087), .ZN(n9009) );
  OR2_X1 U11474 ( .A1(n12088), .A2(n14337), .ZN(n9008) );
  NAND2_X1 U11475 ( .A1(n9966), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9017) );
  NAND2_X1 U11476 ( .A1(n9967), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9016) );
  INV_X1 U11477 ( .A(n9012), .ZN(n9010) );
  NAND2_X1 U11478 ( .A1(n9010), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n9030) );
  INV_X1 U11479 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9011) );
  NAND2_X1 U11480 ( .A1(n9012), .A2(n9011), .ZN(n9013) );
  AND2_X1 U11481 ( .A1(n9030), .A2(n9013), .ZN(n13860) );
  NAND2_X1 U11482 ( .A1(n9060), .A2(n13860), .ZN(n9015) );
  NAND2_X1 U11483 ( .A1(n6475), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9014) );
  NAND4_X1 U11484 ( .A1(n9017), .A2(n9016), .A3(n9015), .A4(n9014), .ZN(n13874) );
  INV_X1 U11485 ( .A(n13874), .ZN(n9018) );
  NAND2_X1 U11486 ( .A1(n13866), .A2(n9018), .ZN(n9116) );
  OR2_X1 U11487 ( .A1(n13866), .A2(n9018), .ZN(n9019) );
  NAND2_X1 U11488 ( .A1(n9116), .A2(n9019), .ZN(n13996) );
  NAND2_X1 U11489 ( .A1(n13866), .A2(n13874), .ZN(n9020) );
  MUX2_X1 U11490 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n9676), .Z(n9038) );
  INV_X1 U11491 ( .A(n9038), .ZN(n9024) );
  XNOR2_X1 U11492 ( .A(n9024), .B(SI_27_), .ZN(n9025) );
  XNOR2_X1 U11493 ( .A(n9041), .B(n9025), .ZN(n13582) );
  NAND2_X1 U11494 ( .A1(n13582), .A2(n12087), .ZN(n9027) );
  OR2_X1 U11495 ( .A1(n12088), .A2(n14336), .ZN(n9026) );
  NAND2_X1 U11496 ( .A1(n9966), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9035) );
  NAND2_X1 U11497 ( .A1(n6475), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n9034) );
  INV_X1 U11498 ( .A(n9030), .ZN(n9028) );
  NAND2_X1 U11499 ( .A1(n9028), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9046) );
  INV_X1 U11500 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9029) );
  NAND2_X1 U11501 ( .A1(n9030), .A2(n9029), .ZN(n9031) );
  NAND2_X1 U11502 ( .A1(n9060), .A2(n13991), .ZN(n9033) );
  NAND2_X1 U11503 ( .A1(n8614), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9032) );
  NAND4_X1 U11504 ( .A1(n9035), .A2(n9034), .A3(n9033), .A4(n9032), .ZN(n13873) );
  XNOR2_X1 U11505 ( .A(n13988), .B(n13873), .ZN(n13981) );
  OR2_X1 U11506 ( .A1(n13988), .A2(n13873), .ZN(n9037) );
  NOR2_X1 U11507 ( .A1(n9038), .A2(SI_27_), .ZN(n9040) );
  NAND2_X1 U11508 ( .A1(n9038), .A2(SI_27_), .ZN(n9039) );
  MUX2_X1 U11509 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n9676), .Z(n9054) );
  XNOR2_X1 U11510 ( .A(n9054), .B(SI_28_), .ZN(n9052) );
  NAND2_X1 U11511 ( .A1(n13578), .A2(n12087), .ZN(n9043) );
  OR2_X1 U11512 ( .A1(n12088), .A2(n14333), .ZN(n9042) );
  NAND2_X1 U11513 ( .A1(n8594), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9051) );
  NAND2_X1 U11514 ( .A1(n9966), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9050) );
  INV_X1 U11515 ( .A(n9046), .ZN(n9044) );
  NAND2_X1 U11516 ( .A1(n9044), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n13948) );
  INV_X1 U11517 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9045) );
  NAND2_X1 U11518 ( .A1(n9046), .A2(n9045), .ZN(n9047) );
  NAND2_X1 U11519 ( .A1(n9060), .A2(n13764), .ZN(n9049) );
  NAND2_X1 U11520 ( .A1(n9967), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9048) );
  NAND4_X1 U11521 ( .A1(n9051), .A2(n9050), .A3(n9049), .A4(n9048), .ZN(n13872) );
  INV_X1 U11522 ( .A(n13872), .ZN(n9119) );
  XNOR2_X1 U11523 ( .A(n14288), .B(n9119), .ZN(n13971) );
  INV_X1 U11524 ( .A(n9054), .ZN(n9055) );
  NAND2_X1 U11525 ( .A1(n9055), .A2(n12212), .ZN(n9056) );
  MUX2_X1 U11526 ( .A(n14330), .B(n13576), .S(n9676), .Z(n9673) );
  XNOR2_X1 U11527 ( .A(n9673), .B(SI_29_), .ZN(n9671) );
  NAND2_X1 U11528 ( .A1(n13575), .A2(n12087), .ZN(n9058) );
  OR2_X1 U11529 ( .A1(n12088), .A2(n14330), .ZN(n9057) );
  NAND2_X1 U11530 ( .A1(n6475), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9064) );
  NAND2_X1 U11531 ( .A1(n9966), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9063) );
  INV_X1 U11532 ( .A(n13948), .ZN(n9059) );
  NAND2_X1 U11533 ( .A1(n9060), .A2(n9059), .ZN(n9062) );
  NAND2_X1 U11534 ( .A1(n9967), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9061) );
  NAND4_X1 U11535 ( .A1(n9064), .A2(n9063), .A3(n9062), .A4(n9061), .ZN(n13871) );
  XNOR2_X1 U11536 ( .A(n14180), .B(n13871), .ZN(n12141) );
  XNOR2_X1 U11537 ( .A(n9065), .B(n12141), .ZN(n13947) );
  NAND2_X1 U11538 ( .A1(n9069), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9068) );
  INV_X1 U11539 ( .A(n12100), .ZN(n9124) );
  NAND2_X1 U11540 ( .A1(n9071), .A2(n9070), .ZN(n9072) );
  NAND2_X1 U11541 ( .A1(n9073), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9074) );
  INV_X1 U11542 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9075) );
  NOR2_X1 U11543 ( .A1(n11952), .A2(n11945), .ZN(n9078) );
  NOR2_X1 U11544 ( .A1(n9078), .A2(n11048), .ZN(n10853) );
  NAND2_X1 U11545 ( .A1(n10853), .A2(n14138), .ZN(n11427) );
  NAND2_X1 U11546 ( .A1(n11942), .A2(n13930), .ZN(n14868) );
  NAND2_X1 U11547 ( .A1(n13897), .A2(n14844), .ZN(n9079) );
  NAND2_X1 U11548 ( .A1(n11950), .A2(n9079), .ZN(n9081) );
  NAND2_X1 U11549 ( .A1(n10341), .A2(n7060), .ZN(n9080) );
  NAND2_X1 U11550 ( .A1(n9081), .A2(n9080), .ZN(n14826) );
  INV_X1 U11551 ( .A(n14825), .ZN(n9082) );
  NAND2_X1 U11552 ( .A1(n14826), .A2(n9082), .ZN(n9083) );
  NAND2_X1 U11553 ( .A1(n9083), .A2(n11959), .ZN(n10860) );
  INV_X1 U11554 ( .A(n12116), .ZN(n11961) );
  INV_X1 U11555 ( .A(n10928), .ZN(n14882) );
  AND2_X1 U11556 ( .A1(n10929), .A2(n14882), .ZN(n9084) );
  NAND2_X1 U11557 ( .A1(n7571), .A2(n10928), .ZN(n9085) );
  NOR2_X1 U11558 ( .A1(n9087), .A2(n14813), .ZN(n9086) );
  NAND2_X1 U11559 ( .A1(n9087), .A2(n14813), .ZN(n9088) );
  INV_X1 U11560 ( .A(n11091), .ZN(n12121) );
  NAND2_X1 U11561 ( .A1(n11979), .A2(n11114), .ZN(n9091) );
  OR2_X1 U11562 ( .A1(n11982), .A2(n9093), .ZN(n9094) );
  INV_X1 U11563 ( .A(n12126), .ZN(n11424) );
  NAND2_X1 U11564 ( .A1(n11991), .A2(n11545), .ZN(n9095) );
  INV_X1 U11565 ( .A(n11371), .ZN(n12127) );
  OR2_X1 U11566 ( .A1(n11995), .A2(n11778), .ZN(n9096) );
  NAND2_X1 U11567 ( .A1(n11374), .A2(n9096), .ZN(n11559) );
  INV_X1 U11568 ( .A(n11560), .ZN(n12128) );
  OR2_X1 U11569 ( .A1(n14630), .A2(n13614), .ZN(n9097) );
  INV_X1 U11570 ( .A(n11448), .ZN(n12130) );
  OR2_X1 U11571 ( .A1(n13791), .A2(n13609), .ZN(n9098) );
  INV_X1 U11572 ( .A(n12132), .ZN(n11468) );
  OR2_X1 U11573 ( .A1(n13837), .A2(n13606), .ZN(n9099) );
  NAND2_X1 U11574 ( .A1(n11467), .A2(n9099), .ZN(n11856) );
  INV_X1 U11575 ( .A(n13883), .ZN(n13805) );
  NAND2_X1 U11576 ( .A1(n14604), .A2(n13805), .ZN(n9100) );
  INV_X1 U11577 ( .A(n14150), .ZN(n12032) );
  AND2_X1 U11578 ( .A1(n14264), .A2(n12032), .ZN(n9102) );
  OR2_X1 U11579 ( .A1(n14264), .A2(n12032), .ZN(n9101) );
  XNOR2_X1 U11580 ( .A(n14257), .B(n13882), .ZN(n14115) );
  NAND2_X1 U11581 ( .A1(n14114), .A2(n14115), .ZN(n9104) );
  INV_X1 U11582 ( .A(n13882), .ZN(n13807) );
  OR2_X1 U11583 ( .A1(n14257), .A2(n13807), .ZN(n9103) );
  INV_X1 U11584 ( .A(n13880), .ZN(n9105) );
  OR2_X1 U11585 ( .A1(n14240), .A2(n9105), .ZN(n9106) );
  INV_X1 U11586 ( .A(n13879), .ZN(n9107) );
  NOR2_X1 U11587 ( .A1(n14076), .A2(n9107), .ZN(n9108) );
  XNOR2_X1 U11588 ( .A(n14221), .B(n13877), .ZN(n14045) );
  INV_X1 U11589 ( .A(n13877), .ZN(n9110) );
  NAND2_X1 U11590 ( .A1(n14221), .A2(n9110), .ZN(n9111) );
  INV_X1 U11591 ( .A(n14030), .ZN(n14025) );
  INV_X1 U11592 ( .A(n13876), .ZN(n9112) );
  OR2_X1 U11593 ( .A1(n14211), .A2(n9112), .ZN(n9113) );
  NAND2_X1 U11594 ( .A1(n14201), .A2(n9114), .ZN(n9115) );
  INV_X1 U11595 ( .A(n13996), .ZN(n13999) );
  NAND2_X1 U11596 ( .A1(n13978), .A2(n13981), .ZN(n13977) );
  INV_X1 U11597 ( .A(n13873), .ZN(n9117) );
  NAND2_X1 U11598 ( .A1(n13988), .A2(n9117), .ZN(n9118) );
  OR2_X1 U11599 ( .A1(n12085), .A2(n12100), .ZN(n9120) );
  OAI21_X2 U11600 ( .B1(n11944), .B2(n14138), .A(n9120), .ZN(n14269) );
  INV_X1 U11601 ( .A(n13866), .ZN(n14196) );
  INV_X1 U11602 ( .A(n13837), .ZN(n14642) );
  NAND2_X1 U11603 ( .A1(n10888), .A2(n14844), .ZN(n14835) );
  INV_X1 U11604 ( .A(n11976), .ZN(n14805) );
  NAND2_X1 U11605 ( .A1(n10911), .A2(n14805), .ZN(n11089) );
  NOR2_X2 U11606 ( .A1(n13791), .A2(n11556), .ZN(n11472) );
  INV_X1 U11607 ( .A(n14257), .ZN(n14127) );
  NAND2_X1 U11608 ( .A1(n14135), .A2(n14127), .ZN(n14121) );
  INV_X1 U11609 ( .A(n14221), .ZN(n14052) );
  NAND2_X1 U11610 ( .A1(n14196), .A2(n14012), .ZN(n14001) );
  AOI21_X1 U11611 ( .B1(n14180), .B2(n13963), .A(n10182), .ZN(n9123) );
  INV_X1 U11612 ( .A(n14180), .ZN(n9121) );
  NAND2_X1 U11613 ( .A1(n9123), .A2(n13941), .ZN(n13956) );
  AND2_X2 U11614 ( .A1(n11943), .A2(n14331), .ZN(n14149) );
  INV_X1 U11615 ( .A(P1_B_REG_SCAN_IN), .ZN(n9132) );
  OR2_X1 U11616 ( .A1(n6487), .A2(n9132), .ZN(n9125) );
  AND2_X1 U11617 ( .A1(n14149), .A2(n9125), .ZN(n13936) );
  NAND2_X1 U11618 ( .A1(n8594), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9128) );
  NAND2_X1 U11619 ( .A1(n9966), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9127) );
  NAND2_X1 U11620 ( .A1(n9967), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9126) );
  NAND3_X1 U11621 ( .A1(n9128), .A2(n9127), .A3(n9126), .ZN(n13870) );
  NAND2_X1 U11622 ( .A1(n13936), .A2(n13870), .ZN(n13949) );
  INV_X1 U11623 ( .A(n14331), .ZN(n10301) );
  NAND2_X1 U11624 ( .A1(n11943), .A2(n10301), .ZN(n13804) );
  INV_X2 U11625 ( .A(n13804), .ZN(n13861) );
  NAND2_X1 U11626 ( .A1(n13872), .A2(n13861), .ZN(n13951) );
  NAND3_X1 U11627 ( .A1(n13956), .A2(n13949), .A3(n13951), .ZN(n9129) );
  NAND2_X1 U11628 ( .A1(n9154), .A2(n9132), .ZN(n9140) );
  INV_X1 U11629 ( .A(n9133), .ZN(n9134) );
  NAND2_X1 U11630 ( .A1(n9134), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9135) );
  MUX2_X1 U11631 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9135), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n9137) );
  NAND2_X1 U11632 ( .A1(n9137), .A2(n9136), .ZN(n14340) );
  NAND3_X1 U11633 ( .A1(n14344), .A2(P1_B_REG_SCAN_IN), .A3(n14340), .ZN(n9139) );
  NAND2_X1 U11634 ( .A1(n9136), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9138) );
  INV_X1 U11635 ( .A(n9151), .ZN(n14339) );
  NAND2_X1 U11636 ( .A1(n14339), .A2(n14340), .ZN(n9954) );
  NAND2_X1 U11637 ( .A1(n14837), .A2(n13930), .ZN(n10173) );
  INV_X1 U11638 ( .A(n10173), .ZN(n10177) );
  NOR2_X1 U11639 ( .A1(n10850), .A2(n10177), .ZN(n9159) );
  NOR4_X1 U11640 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n9150) );
  NOR4_X1 U11641 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n9149) );
  OR4_X1 U11642 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n9147) );
  NOR4_X1 U11643 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9145) );
  NOR4_X1 U11644 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9144) );
  NOR4_X1 U11645 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9143) );
  NOR4_X1 U11646 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9142) );
  NAND4_X1 U11647 ( .A1(n9145), .A2(n9144), .A3(n9143), .A4(n9142), .ZN(n9146)
         );
  NOR4_X1 U11648 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n9147), .A4(n9146), .ZN(n9148) );
  AND3_X1 U11649 ( .A1(n9150), .A2(n9149), .A3(n9148), .ZN(n10191) );
  INV_X1 U11650 ( .A(n14340), .ZN(n9152) );
  NAND2_X1 U11651 ( .A1(n9155), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9157) );
  NAND2_X1 U11652 ( .A1(n12085), .A2(n14138), .ZN(n9158) );
  NAND2_X1 U11653 ( .A1(n11943), .A2(n9158), .ZN(n10176) );
  AND3_X1 U11654 ( .A1(n10172), .A2(n10192), .A3(n10176), .ZN(n10851) );
  AND2_X1 U11655 ( .A1(n9159), .A2(n10851), .ZN(n10257) );
  NAND2_X1 U11656 ( .A1(n14344), .A2(n14339), .ZN(n9957) );
  NAND2_X1 U11657 ( .A1(n11944), .A2(n12100), .ZN(n9161) );
  NOR2_X1 U11658 ( .A1(n9161), .A2(n12085), .ZN(n10178) );
  INV_X1 U11659 ( .A(n10178), .ZN(n10856) );
  INV_X1 U11660 ( .A(n9161), .ZN(n10260) );
  NAND2_X1 U11661 ( .A1(n10260), .A2(n13930), .ZN(n9162) );
  NAND2_X1 U11662 ( .A1(n14180), .A2(n14306), .ZN(n9163) );
  NAND2_X1 U11663 ( .A1(n9164), .A2(n9163), .ZN(P1_U3525) );
  INV_X1 U11664 ( .A(n12226), .ZN(n12570) );
  NAND2_X1 U11665 ( .A1(n12767), .A2(n12570), .ZN(n9165) );
  INV_X1 U11666 ( .A(n12362), .ZN(n9171) );
  INV_X1 U11667 ( .A(n8450), .ZN(n9169) );
  NAND2_X1 U11668 ( .A1(n9169), .A2(P3_B_REG_SCAN_IN), .ZN(n9170) );
  NAND2_X1 U11669 ( .A1(n15200), .A2(n9170), .ZN(n12550) );
  OAI22_X1 U11670 ( .A1(n9171), .A2(n12550), .B1(n12226), .B2(n15183), .ZN(
        n9172) );
  INV_X1 U11671 ( .A(n12217), .ZN(n9192) );
  NOR2_X1 U11672 ( .A1(n9192), .A2(n12880), .ZN(n9176) );
  NOR2_X1 U11673 ( .A1(n9175), .A2(n9176), .ZN(n9177) );
  AND2_X1 U11674 ( .A1(n9178), .A2(n10688), .ZN(n9180) );
  OR2_X1 U11675 ( .A1(n9184), .A2(n9182), .ZN(n10674) );
  NAND2_X1 U11676 ( .A1(n9184), .A2(n9183), .ZN(n11186) );
  AND2_X1 U11677 ( .A1(n10674), .A2(n11186), .ZN(n11188) );
  OAI22_X1 U11678 ( .A1(n15195), .A2(n9185), .B1(n12531), .B2(n11200), .ZN(
        n9187) );
  AOI21_X1 U11679 ( .B1(n9187), .B2(n9186), .A(n8307), .ZN(n9189) );
  MUX2_X1 U11680 ( .A(n11188), .B(n9189), .S(n9188), .Z(n9190) );
  NAND2_X1 U11681 ( .A1(n12766), .A2(n8213), .ZN(n9191) );
  NAND4_X1 U11682 ( .A1(n9219), .A2(n9200), .A3(n9221), .A4(n9226), .ZN(n9203)
         );
  NAND4_X1 U11683 ( .A1(n9812), .A2(n9201), .A3(n7164), .A4(n9224), .ZN(n9202)
         );
  NOR2_X1 U11684 ( .A1(n9203), .A2(n9202), .ZN(n9204) );
  INV_X1 U11685 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9205) );
  INV_X1 U11686 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9208) );
  NAND2_X1 U11687 ( .A1(n10423), .A2(n9743), .ZN(n9216) );
  NAND2_X1 U11688 ( .A1(n9212), .A2(n9213), .ZN(n9439) );
  NAND2_X1 U11689 ( .A1(n9475), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9214) );
  XNOR2_X1 U11690 ( .A(n9214), .B(P2_IR_REG_14__SCAN_IN), .ZN(n13180) );
  AOI22_X1 U11691 ( .A1(n9552), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n9551), 
        .B2(n13180), .ZN(n9215) );
  NOR2_X1 U11692 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n9218) );
  AND2_X1 U11693 ( .A1(n9219), .A2(n9218), .ZN(n9220) );
  XNOR2_X2 U11694 ( .A(n9222), .B(n9221), .ZN(n9248) );
  XNOR2_X2 U11695 ( .A(n9225), .B(n9224), .ZN(n9247) );
  NAND2_X1 U11696 ( .A1(n9834), .A2(n9550), .ZN(n10204) );
  NAND2_X1 U11697 ( .A1(n9232), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9227) );
  INV_X1 U11698 ( .A(n9228), .ZN(n9811) );
  NAND2_X1 U11699 ( .A1(n9230), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9231) );
  MUX2_X1 U11700 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9231), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n9233) );
  NAND2_X1 U11701 ( .A1(n14559), .A2(n9718), .ZN(n9250) );
  NAND2_X1 U11702 ( .A1(n9750), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n9246) );
  NAND2_X1 U11703 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9318) );
  NOR2_X1 U11704 ( .A1(n9318), .A2(n10453), .ZN(n9346) );
  NAND2_X1 U11705 ( .A1(n9346), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9362) );
  INV_X1 U11706 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9361) );
  NAND2_X1 U11707 ( .A1(n9414), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9428) );
  INV_X1 U11708 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9444) );
  NAND2_X1 U11709 ( .A1(n9462), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9464) );
  NAND2_X1 U11710 ( .A1(n9464), .A2(n9238), .ZN(n9239) );
  NAND2_X1 U11711 ( .A1(n9481), .A2(n9239), .ZN(n14550) );
  INV_X1 U11712 ( .A(n14550), .ZN(n14555) );
  NAND2_X1 U11713 ( .A1(n9713), .A2(n14555), .ZN(n9245) );
  NAND2_X1 U11714 ( .A1(n9749), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n9244) );
  NAND2_X1 U11715 ( .A1(n9656), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n9243) );
  NAND4_X1 U11716 ( .A1(n9246), .A2(n9245), .A3(n9244), .A4(n9243), .ZN(n13077) );
  NOR2_X1 U11717 ( .A1(n9267), .A2(n9247), .ZN(n10565) );
  INV_X2 U11718 ( .A(n6526), .ZN(n9737) );
  NAND2_X1 U11719 ( .A1(n13077), .A2(n9737), .ZN(n9249) );
  NAND2_X1 U11720 ( .A1(n9750), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9255) );
  NAND2_X1 U11721 ( .A1(n9749), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9254) );
  AND2_X1 U11722 ( .A1(n9318), .A2(n10453), .ZN(n9251) );
  NOR2_X1 U11723 ( .A1(n9346), .A2(n9251), .ZN(n10665) );
  NAND2_X1 U11724 ( .A1(n9713), .A2(n10665), .ZN(n9253) );
  NAND2_X1 U11725 ( .A1(n9656), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9252) );
  NAND4_X1 U11726 ( .A1(n9255), .A2(n9254), .A3(n9253), .A4(n9252), .ZN(n13087) );
  NAND2_X1 U11727 ( .A1(n13087), .A2(n9413), .ZN(n9261) );
  INV_X1 U11728 ( .A(n9256), .ZN(n9257) );
  NAND2_X1 U11729 ( .A1(n9257), .A2(n9323), .ZN(n9325) );
  NAND2_X1 U11730 ( .A1(n9325), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9258) );
  XNOR2_X1 U11731 ( .A(n9258), .B(P2_IR_REG_5__SCAN_IN), .ZN(n13132) );
  AOI22_X1 U11732 ( .A1(n9552), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9551), .B2(
        n13132), .ZN(n9259) );
  NAND2_X1 U11733 ( .A1(n15105), .A2(n9756), .ZN(n9260) );
  NAND2_X1 U11734 ( .A1(n9306), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9265) );
  NAND2_X1 U11735 ( .A1(n9540), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n9262) );
  NAND2_X1 U11736 ( .A1(n9676), .A2(SI_0_), .ZN(n9266) );
  XNOR2_X1 U11737 ( .A(n9266), .B(n9965), .ZN(n13600) );
  MUX2_X1 U11738 ( .A(n7397), .B(n13600), .S(n9290), .Z(n15067) );
  NAND2_X1 U11739 ( .A1(n9782), .A2(n15067), .ZN(n9783) );
  INV_X4 U11740 ( .A(n6526), .ZN(n9756) );
  NAND2_X1 U11741 ( .A1(n9783), .A2(n9756), .ZN(n9270) );
  INV_X1 U11742 ( .A(n15067), .ZN(n15089) );
  NAND2_X1 U11743 ( .A1(n15067), .A2(n9267), .ZN(n9269) );
  OAI211_X1 U11744 ( .C1(n9267), .C2(n15067), .A(n9782), .B(n9413), .ZN(n9268)
         );
  NAND2_X1 U11745 ( .A1(n6525), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9274) );
  NAND2_X1 U11746 ( .A1(n9306), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9272) );
  NAND2_X1 U11747 ( .A1(n9540), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n9271) );
  NAND4_X1 U11748 ( .A1(n9274), .A2(n9273), .A3(n9272), .A4(n9271), .ZN(n9833)
         );
  NAND2_X1 U11749 ( .A1(n9833), .A2(n9413), .ZN(n9280) );
  INV_X1 U11750 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n9276) );
  NAND2_X1 U11751 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9275) );
  XNOR2_X1 U11752 ( .A(n9276), .B(n9275), .ZN(n10006) );
  NAND2_X1 U11753 ( .A1(n10502), .A2(n9756), .ZN(n9279) );
  NAND2_X1 U11754 ( .A1(n9280), .A2(n9279), .ZN(n9298) );
  NAND2_X1 U11755 ( .A1(n6525), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9285) );
  NAND2_X1 U11756 ( .A1(n9281), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n9284) );
  NAND2_X1 U11757 ( .A1(n9306), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9283) );
  NAND2_X1 U11758 ( .A1(n9540), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9282) );
  OR2_X1 U11759 ( .A1(n9287), .A2(n9208), .ZN(n9289) );
  XNOR2_X1 U11760 ( .A(n9289), .B(n9288), .ZN(n14929) );
  NOR2_X1 U11761 ( .A1(n9293), .A2(n9786), .ZN(n9294) );
  AOI21_X1 U11762 ( .B1(n9784), .B2(n9756), .A(n9294), .ZN(n9301) );
  NAND2_X1 U11763 ( .A1(n9785), .A2(n9756), .ZN(n9296) );
  NAND2_X1 U11764 ( .A1(n9784), .A2(n9413), .ZN(n9295) );
  NAND2_X1 U11765 ( .A1(n9296), .A2(n9295), .ZN(n9300) );
  OAI22_X1 U11766 ( .A1(n9299), .A2(n9298), .B1(n9301), .B2(n9300), .ZN(n9304)
         );
  AOI22_X1 U11767 ( .A1(n9833), .A2(n9756), .B1(n9413), .B2(n10502), .ZN(n9297) );
  AOI21_X1 U11768 ( .B1(n9299), .B2(n9298), .A(n9297), .ZN(n9303) );
  NAND2_X1 U11769 ( .A1(n9301), .A2(n9300), .ZN(n9302) );
  INV_X1 U11770 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9305) );
  NAND2_X1 U11771 ( .A1(n9713), .A2(n9305), .ZN(n9310) );
  NAND2_X1 U11772 ( .A1(n9750), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n9309) );
  NAND2_X1 U11773 ( .A1(n9306), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9308) );
  NAND2_X1 U11774 ( .A1(n6525), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9307) );
  NAND2_X1 U11775 ( .A1(n9780), .A2(n9413), .ZN(n9315) );
  NAND2_X1 U11776 ( .A1(n9311), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9312) );
  XNOR2_X1 U11777 ( .A(n9312), .B(n9193), .ZN(n13103) );
  OR2_X1 U11778 ( .A1(n9744), .A2(n9903), .ZN(n9313) );
  NAND2_X1 U11779 ( .A1(n10631), .A2(n9737), .ZN(n9314) );
  NAND2_X1 U11780 ( .A1(n9315), .A2(n9314), .ZN(n9317) );
  AOI22_X1 U11781 ( .A1(n9780), .A2(n9756), .B1(n9413), .B2(n10631), .ZN(n9316) );
  NAND2_X1 U11782 ( .A1(n9750), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9322) );
  NAND2_X1 U11783 ( .A1(n9749), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9321) );
  OAI21_X1 U11784 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n9318), .ZN(n10491) );
  INV_X1 U11785 ( .A(n10491), .ZN(n10642) );
  NAND2_X1 U11786 ( .A1(n9713), .A2(n10642), .ZN(n9320) );
  NAND2_X1 U11787 ( .A1(n9656), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9319) );
  NAND2_X1 U11788 ( .A1(n13088), .A2(n9756), .ZN(n9330) );
  NOR2_X1 U11789 ( .A1(n9912), .A2(n9286), .ZN(n9328) );
  NAND2_X1 U11790 ( .A1(n9256), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9324) );
  MUX2_X1 U11791 ( .A(n9324), .B(P2_IR_REG_31__SCAN_IN), .S(n9323), .Z(n9326)
         );
  NAND2_X1 U11792 ( .A1(n9326), .A2(n9325), .ZN(n10012) );
  OAI22_X1 U11793 ( .A1(n9744), .A2(n9904), .B1(n9290), .B2(n10012), .ZN(n9327) );
  NAND2_X1 U11794 ( .A1(n10657), .A2(n9718), .ZN(n9329) );
  NAND2_X1 U11795 ( .A1(n9330), .A2(n9329), .ZN(n9336) );
  NAND2_X1 U11796 ( .A1(n9335), .A2(n9336), .ZN(n9334) );
  NAND2_X1 U11797 ( .A1(n13088), .A2(n9413), .ZN(n9332) );
  NAND2_X1 U11798 ( .A1(n10657), .A2(n9756), .ZN(n9331) );
  NAND2_X1 U11799 ( .A1(n9332), .A2(n9331), .ZN(n9333) );
  NAND2_X1 U11800 ( .A1(n9334), .A2(n9333), .ZN(n9340) );
  INV_X1 U11801 ( .A(n9335), .ZN(n9338) );
  INV_X1 U11802 ( .A(n9336), .ZN(n9337) );
  NAND2_X1 U11803 ( .A1(n9338), .A2(n9337), .ZN(n9339) );
  AOI22_X1 U11804 ( .A1(n9737), .A2(n13087), .B1(n15105), .B2(n9718), .ZN(
        n9341) );
  OR2_X1 U11805 ( .A1(n9927), .A2(n9286), .ZN(n9345) );
  OR2_X1 U11806 ( .A1(n9212), .A2(n9208), .ZN(n9343) );
  XNOR2_X1 U11807 ( .A(n9343), .B(P2_IR_REG_6__SCAN_IN), .ZN(n13144) );
  AOI22_X1 U11808 ( .A1(n9552), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9551), .B2(
        n13144), .ZN(n9344) );
  NAND2_X1 U11809 ( .A1(n10997), .A2(n9413), .ZN(n9353) );
  NAND2_X1 U11810 ( .A1(n9656), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9351) );
  NAND2_X1 U11811 ( .A1(n9750), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n9350) );
  OR2_X1 U11812 ( .A1(n9346), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9347) );
  AND2_X1 U11813 ( .A1(n9362), .A2(n9347), .ZN(n10831) );
  NAND2_X1 U11814 ( .A1(n9713), .A2(n10831), .ZN(n9349) );
  NAND2_X1 U11815 ( .A1(n9749), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9348) );
  NAND4_X1 U11816 ( .A1(n9351), .A2(n9350), .A3(n9349), .A4(n9348), .ZN(n13086) );
  NAND2_X1 U11817 ( .A1(n13086), .A2(n9737), .ZN(n9352) );
  NAND2_X1 U11818 ( .A1(n9353), .A2(n9352), .ZN(n9356) );
  INV_X1 U11819 ( .A(n13086), .ZN(n10996) );
  NAND2_X1 U11820 ( .A1(n10997), .A2(n9737), .ZN(n9354) );
  OAI21_X1 U11821 ( .B1(n9293), .B2(n10996), .A(n9354), .ZN(n9355) );
  OR2_X1 U11822 ( .A1(n9935), .A2(n9286), .ZN(n9360) );
  NAND2_X1 U11823 ( .A1(n9212), .A2(n9357), .ZN(n9379) );
  NAND2_X1 U11824 ( .A1(n9379), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9358) );
  XNOR2_X1 U11825 ( .A(n9358), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13156) );
  AOI22_X1 U11826 ( .A1(n9552), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9551), .B2(
        n13156), .ZN(n9359) );
  NAND2_X1 U11827 ( .A1(n15048), .A2(n9756), .ZN(n9369) );
  NAND2_X1 U11828 ( .A1(n9656), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9367) );
  NAND2_X1 U11829 ( .A1(n9750), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9366) );
  NAND2_X1 U11830 ( .A1(n9362), .A2(n9361), .ZN(n9363) );
  AND2_X1 U11831 ( .A1(n9385), .A2(n9363), .ZN(n15052) );
  NAND2_X1 U11832 ( .A1(n9713), .A2(n15052), .ZN(n9365) );
  NAND2_X1 U11833 ( .A1(n9749), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9364) );
  NAND4_X1 U11834 ( .A1(n9367), .A2(n9366), .A3(n9365), .A4(n9364), .ZN(n13085) );
  NAND2_X1 U11835 ( .A1(n13085), .A2(n9413), .ZN(n9368) );
  NAND2_X1 U11836 ( .A1(n9369), .A2(n9368), .ZN(n9374) );
  NAND2_X1 U11837 ( .A1(n9373), .A2(n9374), .ZN(n9372) );
  INV_X1 U11838 ( .A(n13085), .ZN(n11125) );
  NAND2_X1 U11839 ( .A1(n15048), .A2(n9413), .ZN(n9370) );
  OAI21_X1 U11840 ( .B1(n11125), .B2(n6526), .A(n9370), .ZN(n9371) );
  NAND2_X1 U11841 ( .A1(n9372), .A2(n9371), .ZN(n9378) );
  NAND2_X1 U11842 ( .A1(n9376), .A2(n9375), .ZN(n9377) );
  NAND2_X1 U11843 ( .A1(n9381), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9380) );
  MUX2_X1 U11844 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9380), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n9382) );
  AOI22_X1 U11845 ( .A1(n9552), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9551), .B2(
        n10018), .ZN(n9383) );
  NAND2_X1 U11846 ( .A1(n11222), .A2(n9413), .ZN(n9392) );
  NAND2_X1 U11847 ( .A1(n9656), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9390) );
  NAND2_X1 U11848 ( .A1(n9750), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n9389) );
  NAND2_X1 U11849 ( .A1(n9385), .A2(n9384), .ZN(n9386) );
  NAND2_X1 U11850 ( .A1(n9398), .A2(n9386), .ZN(n11075) );
  INV_X1 U11851 ( .A(n11075), .ZN(n11138) );
  NAND2_X1 U11852 ( .A1(n9713), .A2(n11138), .ZN(n9388) );
  NAND2_X1 U11853 ( .A1(n9749), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9387) );
  NAND4_X1 U11854 ( .A1(n9390), .A2(n9389), .A3(n9388), .A4(n9387), .ZN(n13084) );
  NAND2_X1 U11855 ( .A1(n13084), .A2(n9756), .ZN(n9391) );
  AOI22_X1 U11856 ( .A1(n11222), .A2(n9756), .B1(n9718), .B2(n13084), .ZN(
        n9393) );
  OR2_X1 U11857 ( .A1(n9945), .A2(n9286), .ZN(n9396) );
  NAND2_X1 U11858 ( .A1(n9407), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9394) );
  XNOR2_X1 U11859 ( .A(n9394), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10020) );
  AOI22_X1 U11860 ( .A1(n9552), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n9551), .B2(
        n10020), .ZN(n9395) );
  NAND2_X1 U11861 ( .A1(n11274), .A2(n9756), .ZN(n9404) );
  NAND2_X1 U11862 ( .A1(n9750), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n9402) );
  NAND2_X1 U11863 ( .A1(n9656), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9401) );
  NOR2_X1 U11864 ( .A1(n9414), .A2(n6577), .ZN(n11231) );
  NAND2_X1 U11865 ( .A1(n9713), .A2(n11231), .ZN(n9400) );
  NAND2_X1 U11866 ( .A1(n9749), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n9399) );
  NAND4_X1 U11867 ( .A1(n9402), .A2(n9401), .A3(n9400), .A4(n9399), .ZN(n13082) );
  NAND2_X1 U11868 ( .A1(n13082), .A2(n9413), .ZN(n9403) );
  AOI22_X1 U11869 ( .A1(n11274), .A2(n9718), .B1(n9737), .B2(n13082), .ZN(
        n9405) );
  INV_X1 U11870 ( .A(n9407), .ZN(n9409) );
  INV_X1 U11871 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9408) );
  NAND2_X1 U11872 ( .A1(n9409), .A2(n9408), .ZN(n9424) );
  NAND2_X1 U11873 ( .A1(n9424), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9410) );
  XNOR2_X1 U11874 ( .A(n9410), .B(P2_IR_REG_10__SCAN_IN), .ZN(n14973) );
  AOI22_X1 U11875 ( .A1(n9552), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n9551), 
        .B2(n14973), .ZN(n9411) );
  NAND2_X1 U11876 ( .A1(n11465), .A2(n9413), .ZN(n9421) );
  NAND2_X1 U11877 ( .A1(n9656), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9419) );
  NAND2_X1 U11878 ( .A1(n9750), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n9418) );
  OR2_X1 U11879 ( .A1(n9414), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9415) );
  AND2_X1 U11880 ( .A1(n9415), .A2(n9428), .ZN(n11265) );
  NAND2_X1 U11881 ( .A1(n9713), .A2(n11265), .ZN(n9417) );
  NAND2_X1 U11882 ( .A1(n9749), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9416) );
  NAND4_X1 U11883 ( .A1(n9419), .A2(n9418), .A3(n9417), .A4(n9416), .ZN(n13081) );
  NAND2_X1 U11884 ( .A1(n13081), .A2(n9756), .ZN(n9420) );
  NAND2_X1 U11885 ( .A1(n11465), .A2(n9756), .ZN(n9422) );
  NAND2_X1 U11886 ( .A1(n9973), .A2(n9743), .ZN(n9427) );
  OAI21_X1 U11887 ( .B1(n9424), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9425) );
  XNOR2_X1 U11888 ( .A(n9425), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10241) );
  AOI22_X1 U11889 ( .A1(n9552), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n9551), 
        .B2(n10241), .ZN(n9426) );
  NAND2_X1 U11890 ( .A1(n15122), .A2(n9756), .ZN(n9435) );
  NAND2_X1 U11891 ( .A1(n9656), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n9433) );
  NAND2_X1 U11892 ( .A1(n9750), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n9432) );
  NAND2_X1 U11893 ( .A1(n9428), .A2(n11361), .ZN(n9429) );
  AND2_X1 U11894 ( .A1(n9445), .A2(n9429), .ZN(n11364) );
  NAND2_X1 U11895 ( .A1(n9713), .A2(n11364), .ZN(n9431) );
  NAND2_X1 U11896 ( .A1(n9749), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9430) );
  NAND4_X1 U11897 ( .A1(n9433), .A2(n9432), .A3(n9431), .A4(n9430), .ZN(n13080) );
  NAND2_X1 U11898 ( .A1(n13080), .A2(n9718), .ZN(n9434) );
  NAND2_X1 U11899 ( .A1(n9435), .A2(n9434), .ZN(n9437) );
  AOI22_X1 U11900 ( .A1(n15122), .A2(n9718), .B1(n9756), .B2(n13080), .ZN(
        n9436) );
  NAND2_X1 U11901 ( .A1(n10073), .A2(n9743), .ZN(n9443) );
  NAND2_X1 U11902 ( .A1(n9439), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9440) );
  MUX2_X1 U11903 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9440), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n9441) );
  AND2_X1 U11904 ( .A1(n9441), .A2(n9456), .ZN(n10244) );
  AOI22_X1 U11905 ( .A1(n9552), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n9551), 
        .B2(n10244), .ZN(n9442) );
  CLKBUF_X3 U11906 ( .A(n9413), .Z(n9718) );
  NAND2_X1 U11907 ( .A1(n11722), .A2(n9718), .ZN(n9452) );
  NAND2_X1 U11908 ( .A1(n9656), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n9450) );
  NAND2_X1 U11909 ( .A1(n9750), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9449) );
  AND2_X1 U11910 ( .A1(n9445), .A2(n9444), .ZN(n9446) );
  NOR2_X1 U11911 ( .A1(n9462), .A2(n9446), .ZN(n11621) );
  NAND2_X1 U11912 ( .A1(n9713), .A2(n11621), .ZN(n9448) );
  NAND2_X1 U11913 ( .A1(n9749), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n9447) );
  NAND4_X1 U11914 ( .A1(n9450), .A2(n9449), .A3(n9448), .A4(n9447), .ZN(n13079) );
  NAND2_X1 U11915 ( .A1(n13079), .A2(n9756), .ZN(n9451) );
  NAND2_X1 U11916 ( .A1(n9452), .A2(n9451), .ZN(n9455) );
  NAND2_X1 U11917 ( .A1(n11722), .A2(n9756), .ZN(n9453) );
  OAI21_X1 U11918 ( .B1(n9293), .B2(n11721), .A(n9453), .ZN(n9454) );
  NAND2_X1 U11919 ( .A1(n10213), .A2(n9743), .ZN(n9461) );
  NAND2_X1 U11920 ( .A1(n9456), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9458) );
  MUX2_X1 U11921 ( .A(n9458), .B(P2_IR_REG_31__SCAN_IN), .S(n9457), .Z(n9459)
         );
  AND2_X1 U11922 ( .A1(n9459), .A2(n9475), .ZN(n10583) );
  AOI22_X1 U11923 ( .A1(n9552), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n9551), 
        .B2(n10583), .ZN(n9460) );
  NAND2_X1 U11924 ( .A1(n14573), .A2(n9756), .ZN(n9470) );
  NAND2_X1 U11925 ( .A1(n9656), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9468) );
  NAND2_X1 U11926 ( .A1(n9750), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n9467) );
  OR2_X1 U11927 ( .A1(n9462), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9463) );
  AND2_X1 U11928 ( .A1(n9464), .A2(n9463), .ZN(n11656) );
  NAND2_X1 U11929 ( .A1(n9713), .A2(n11656), .ZN(n9466) );
  NAND2_X1 U11930 ( .A1(n9749), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9465) );
  NAND4_X1 U11931 ( .A1(n9468), .A2(n9467), .A3(n9466), .A4(n9465), .ZN(n13078) );
  NAND2_X1 U11932 ( .A1(n13078), .A2(n9718), .ZN(n9469) );
  AOI22_X1 U11933 ( .A1(n14573), .A2(n9718), .B1(n9737), .B2(n13078), .ZN(
        n9471) );
  INV_X1 U11934 ( .A(n13077), .ZN(n11881) );
  NAND2_X1 U11935 ( .A1(n14559), .A2(n9756), .ZN(n9473) );
  OAI21_X1 U11936 ( .B1(n9293), .B2(n11881), .A(n9473), .ZN(n9474) );
  NAND2_X1 U11937 ( .A1(n10496), .A2(n9743), .ZN(n9479) );
  OAI21_X1 U11938 ( .B1(n9475), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9477) );
  XNOR2_X1 U11939 ( .A(n9477), .B(n9476), .ZN(n13181) );
  INV_X1 U11940 ( .A(n13181), .ZN(n14999) );
  AOI22_X1 U11941 ( .A1(n9552), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n9551), 
        .B2(n14999), .ZN(n9478) );
  NAND2_X1 U11942 ( .A1(n13546), .A2(n9737), .ZN(n9488) );
  NAND2_X1 U11943 ( .A1(n9540), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n9486) );
  INV_X1 U11944 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9480) );
  AND2_X1 U11945 ( .A1(n9481), .A2(n9480), .ZN(n9482) );
  NOR2_X1 U11946 ( .A1(n9500), .A2(n9482), .ZN(n13058) );
  NAND2_X1 U11947 ( .A1(n9713), .A2(n13058), .ZN(n9485) );
  NAND2_X1 U11948 ( .A1(n9749), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n9484) );
  NAND2_X1 U11949 ( .A1(n9656), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n9483) );
  NAND4_X1 U11950 ( .A1(n9486), .A2(n9485), .A3(n9484), .A4(n9483), .ZN(n13076) );
  NAND2_X1 U11951 ( .A1(n13076), .A2(n9718), .ZN(n9487) );
  NAND2_X1 U11952 ( .A1(n9488), .A2(n9487), .ZN(n9490) );
  AOI22_X1 U11953 ( .A1(n13546), .A2(n9718), .B1(n9756), .B2(n13076), .ZN(
        n9489) );
  NOR2_X1 U11954 ( .A1(n9491), .A2(n9490), .ZN(n9492) );
  NAND2_X1 U11955 ( .A1(n10445), .A2(n9743), .ZN(n9499) );
  NOR2_X1 U11956 ( .A1(n9217), .A2(n9208), .ZN(n9494) );
  MUX2_X1 U11957 ( .A(n9208), .B(n9494), .S(P2_IR_REG_16__SCAN_IN), .Z(n9497)
         );
  INV_X1 U11958 ( .A(n9495), .ZN(n9496) );
  OR2_X1 U11959 ( .A1(n9497), .A2(n9496), .ZN(n13171) );
  AOI22_X1 U11960 ( .A1(n9552), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n9551), 
        .B2(n15013), .ZN(n9498) );
  NAND2_X1 U11961 ( .A1(n13538), .A2(n9718), .ZN(n9508) );
  NOR2_X1 U11962 ( .A1(n9500), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9501) );
  OR2_X1 U11963 ( .A1(n9514), .A2(n9501), .ZN(n11927) );
  INV_X1 U11964 ( .A(n11927), .ZN(n9502) );
  NAND2_X1 U11965 ( .A1(n9502), .A2(n9713), .ZN(n9506) );
  NAND2_X1 U11966 ( .A1(n9750), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n9505) );
  NAND2_X1 U11967 ( .A1(n9749), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n9504) );
  NAND2_X1 U11968 ( .A1(n9656), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n9503) );
  NAND4_X1 U11969 ( .A1(n9506), .A2(n9505), .A3(n9504), .A4(n9503), .ZN(n13233) );
  NAND2_X1 U11970 ( .A1(n13233), .A2(n9737), .ZN(n9507) );
  NAND2_X1 U11971 ( .A1(n9508), .A2(n9507), .ZN(n9510) );
  AOI22_X1 U11972 ( .A1(n13538), .A2(n9756), .B1(n9718), .B2(n13233), .ZN(
        n9509) );
  NAND2_X1 U11973 ( .A1(n10465), .A2(n9743), .ZN(n9513) );
  NAND2_X1 U11974 ( .A1(n9495), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9511) );
  XNOR2_X1 U11975 ( .A(n9511), .B(P2_IR_REG_17__SCAN_IN), .ZN(n15027) );
  AOI22_X1 U11976 ( .A1(n9552), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9551), 
        .B2(n15027), .ZN(n9512) );
  NAND2_X1 U11977 ( .A1(n13533), .A2(n9737), .ZN(n9522) );
  OR2_X1 U11978 ( .A1(n9514), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9515) );
  NAND2_X1 U11979 ( .A1(n9538), .A2(n9515), .ZN(n13441) );
  NAND2_X1 U11980 ( .A1(n9749), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9516) );
  OAI21_X1 U11981 ( .B1(n13441), .B2(n9605), .A(n9516), .ZN(n9520) );
  NAND2_X1 U11982 ( .A1(n9656), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9518) );
  NAND2_X1 U11983 ( .A1(n9750), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n9517) );
  NAND2_X1 U11984 ( .A1(n9518), .A2(n9517), .ZN(n9519) );
  NAND2_X1 U11985 ( .A1(n13236), .A2(n9718), .ZN(n9521) );
  NAND2_X1 U11986 ( .A1(n9522), .A2(n9521), .ZN(n9528) );
  NAND2_X1 U11987 ( .A1(n13533), .A2(n9718), .ZN(n9524) );
  NAND2_X1 U11988 ( .A1(n13236), .A2(n9737), .ZN(n9523) );
  NAND2_X1 U11989 ( .A1(n9524), .A2(n9523), .ZN(n9525) );
  NAND2_X1 U11990 ( .A1(n9526), .A2(n9525), .ZN(n9532) );
  INV_X1 U11991 ( .A(n9527), .ZN(n9530) );
  INV_X1 U11992 ( .A(n9528), .ZN(n9529) );
  NAND2_X1 U11993 ( .A1(n9530), .A2(n9529), .ZN(n9531) );
  NAND2_X1 U11994 ( .A1(n9532), .A2(n9531), .ZN(n9547) );
  NAND2_X1 U11995 ( .A1(n10990), .A2(n9743), .ZN(n9536) );
  NAND2_X1 U11996 ( .A1(n9533), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9534) );
  XNOR2_X1 U11997 ( .A(n9534), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13175) );
  AOI22_X1 U11998 ( .A1(n9552), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9551), 
        .B2(n13175), .ZN(n9535) );
  NAND2_X1 U11999 ( .A1(n13424), .A2(n9718), .ZN(n9544) );
  INV_X1 U12000 ( .A(n9749), .ZN(n9685) );
  INV_X1 U12001 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n13528) );
  INV_X1 U12002 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9537) );
  NAND2_X1 U12003 ( .A1(n9538), .A2(n9537), .ZN(n9539) );
  NAND2_X1 U12004 ( .A1(n9556), .A2(n9539), .ZN(n13419) );
  OR2_X1 U12005 ( .A1(n13419), .A2(n9605), .ZN(n9542) );
  AOI22_X1 U12006 ( .A1(n9656), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9540), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n9541) );
  OAI211_X1 U12007 ( .C1(n9685), .C2(n13528), .A(n9542), .B(n9541), .ZN(n13239) );
  NAND2_X1 U12008 ( .A1(n13239), .A2(n9737), .ZN(n9543) );
  NAND2_X1 U12009 ( .A1(n9544), .A2(n9543), .ZN(n9546) );
  AOI22_X1 U12010 ( .A1(n13424), .A2(n9756), .B1(n9718), .B2(n13239), .ZN(
        n9545) );
  NOR2_X1 U12011 ( .A1(n9547), .A2(n9546), .ZN(n9548) );
  NAND2_X1 U12012 ( .A1(n11204), .A2(n9743), .ZN(n9554) );
  AOI22_X1 U12013 ( .A1(n9552), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9550), 
        .B2(n9551), .ZN(n9553) );
  NAND2_X1 U12014 ( .A1(n13518), .A2(n9737), .ZN(n9561) );
  INV_X1 U12015 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9555) );
  NAND2_X1 U12016 ( .A1(n9556), .A2(n9555), .ZN(n9557) );
  NAND2_X1 U12017 ( .A1(n9568), .A2(n9557), .ZN(n13401) );
  AOI22_X1 U12018 ( .A1(n9749), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n9750), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n9559) );
  NAND2_X1 U12019 ( .A1(n9656), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n9558) );
  OAI211_X1 U12020 ( .C1(n13401), .C2(n9605), .A(n9559), .B(n9558), .ZN(n13075) );
  NAND2_X1 U12021 ( .A1(n13075), .A2(n9718), .ZN(n9560) );
  NAND2_X1 U12022 ( .A1(n9561), .A2(n9560), .ZN(n9564) );
  INV_X1 U12023 ( .A(n13075), .ZN(n13218) );
  NAND2_X1 U12024 ( .A1(n13518), .A2(n9718), .ZN(n9562) );
  OAI21_X1 U12025 ( .B1(n13218), .B2(n6526), .A(n9562), .ZN(n9563) );
  INV_X1 U12026 ( .A(n9564), .ZN(n9565) );
  NAND2_X1 U12027 ( .A1(n11326), .A2(n9743), .ZN(n9567) );
  OR2_X1 U12028 ( .A1(n9744), .A2(n11327), .ZN(n9566) );
  NAND2_X1 U12029 ( .A1(n13387), .A2(n9718), .ZN(n9577) );
  INV_X1 U12030 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13019) );
  AND2_X1 U12031 ( .A1(n9568), .A2(n13019), .ZN(n9569) );
  NOR2_X1 U12032 ( .A1(n9585), .A2(n9569), .ZN(n13018) );
  NAND2_X1 U12033 ( .A1(n13018), .A2(n9713), .ZN(n9575) );
  INV_X1 U12034 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9572) );
  NAND2_X1 U12035 ( .A1(n9656), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9571) );
  NAND2_X1 U12036 ( .A1(n9750), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n9570) );
  OAI211_X1 U12037 ( .C1(n9572), .C2(n9685), .A(n9571), .B(n9570), .ZN(n9573)
         );
  INV_X1 U12038 ( .A(n9573), .ZN(n9574) );
  NAND2_X1 U12039 ( .A1(n9575), .A2(n9574), .ZN(n13245) );
  NAND2_X1 U12040 ( .A1(n13245), .A2(n9737), .ZN(n9576) );
  NAND2_X1 U12041 ( .A1(n9577), .A2(n9576), .ZN(n9579) );
  AOI22_X1 U12042 ( .A1(n13387), .A2(n9756), .B1(n9718), .B2(n13245), .ZN(
        n9578) );
  NOR2_X1 U12043 ( .A1(n9580), .A2(n9579), .ZN(n9581) );
  NAND2_X1 U12044 ( .A1(n11437), .A2(n9743), .ZN(n9584) );
  OR2_X1 U12045 ( .A1(n9744), .A2(n11441), .ZN(n9583) );
  NAND2_X1 U12046 ( .A1(n13375), .A2(n9737), .ZN(n9594) );
  OR2_X1 U12047 ( .A1(n9585), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n9586) );
  NAND2_X1 U12048 ( .A1(n9585), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n9602) );
  AND2_X1 U12049 ( .A1(n9586), .A2(n9602), .ZN(n13374) );
  NAND2_X1 U12050 ( .A1(n13374), .A2(n9713), .ZN(n9592) );
  INV_X1 U12051 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n15261) );
  NAND2_X1 U12052 ( .A1(n9656), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9588) );
  NAND2_X1 U12053 ( .A1(n9749), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n9587) );
  OAI211_X1 U12054 ( .C1(n9589), .C2(n15261), .A(n9588), .B(n9587), .ZN(n9590)
         );
  INV_X1 U12055 ( .A(n9590), .ZN(n9591) );
  NAND2_X1 U12056 ( .A1(n9592), .A2(n9591), .ZN(n13247) );
  NAND2_X1 U12057 ( .A1(n13247), .A2(n9718), .ZN(n9593) );
  INV_X1 U12058 ( .A(n13247), .ZN(n13224) );
  NAND2_X1 U12059 ( .A1(n13375), .A2(n9718), .ZN(n9595) );
  OAI21_X1 U12060 ( .B1(n13224), .B2(n6526), .A(n9595), .ZN(n9596) );
  XNOR2_X1 U12061 ( .A(n9598), .B(n9597), .ZN(n11715) );
  NAND2_X1 U12062 ( .A1(n11715), .A2(n9743), .ZN(n9600) );
  OR2_X1 U12063 ( .A1(n9744), .A2(n11717), .ZN(n9599) );
  NAND2_X1 U12064 ( .A1(n13501), .A2(n9718), .ZN(n9613) );
  INV_X1 U12065 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9601) );
  NAND2_X1 U12066 ( .A1(n9602), .A2(n9601), .ZN(n9604) );
  INV_X1 U12067 ( .A(n9621), .ZN(n9603) );
  NAND2_X1 U12068 ( .A1(n9604), .A2(n9603), .ZN(n13358) );
  INV_X1 U12069 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9608) );
  NAND2_X1 U12070 ( .A1(n9750), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9607) );
  NAND2_X1 U12071 ( .A1(n9656), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9606) );
  OAI211_X1 U12072 ( .C1(n9685), .C2(n9608), .A(n9607), .B(n9606), .ZN(n9609)
         );
  INV_X1 U12073 ( .A(n9609), .ZN(n9610) );
  NAND2_X1 U12074 ( .A1(n13248), .A2(n9737), .ZN(n9612) );
  NAND2_X1 U12075 ( .A1(n9613), .A2(n9612), .ZN(n9615) );
  AOI22_X1 U12076 ( .A1(n13501), .A2(n9756), .B1(n9718), .B2(n13248), .ZN(
        n9614) );
  AOI21_X1 U12077 ( .B1(n9616), .B2(n9615), .A(n9614), .ZN(n9618) );
  NOR2_X1 U12078 ( .A1(n9616), .A2(n9615), .ZN(n9617) );
  NAND2_X1 U12079 ( .A1(n11793), .A2(n9743), .ZN(n9620) );
  OR2_X1 U12080 ( .A1(n9744), .A2(n11796), .ZN(n9619) );
  NAND2_X1 U12081 ( .A1(n13225), .A2(n9737), .ZN(n9627) );
  NAND2_X1 U12082 ( .A1(n9656), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9625) );
  NAND2_X1 U12083 ( .A1(n9750), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9624) );
  NAND2_X1 U12084 ( .A1(n9621), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n9632) );
  OAI21_X1 U12085 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(n9621), .A(n9632), .ZN(
        n12953) );
  INV_X1 U12086 ( .A(n12953), .ZN(n13345) );
  NAND2_X1 U12087 ( .A1(n9713), .A2(n13345), .ZN(n9623) );
  NAND2_X1 U12088 ( .A1(n9749), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n9622) );
  NAND4_X1 U12089 ( .A1(n9625), .A2(n9624), .A3(n9623), .A4(n9622), .ZN(n13226) );
  NAND2_X1 U12090 ( .A1(n13226), .A2(n9718), .ZN(n9626) );
  AOI22_X1 U12091 ( .A1(n13225), .A2(n9718), .B1(n9737), .B2(n13226), .ZN(
        n9628) );
  NAND2_X1 U12092 ( .A1(n13594), .A2(n9743), .ZN(n9630) );
  INV_X1 U12093 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13598) );
  OR2_X1 U12094 ( .A1(n9744), .A2(n13598), .ZN(n9629) );
  NAND2_X1 U12095 ( .A1(n13488), .A2(n9718), .ZN(n9640) );
  NAND2_X1 U12096 ( .A1(n9750), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9638) );
  NAND2_X1 U12097 ( .A1(n9656), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9637) );
  INV_X1 U12098 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9631) );
  NAND2_X1 U12099 ( .A1(n9631), .A2(n9632), .ZN(n9634) );
  INV_X1 U12100 ( .A(n9632), .ZN(n9633) );
  INV_X1 U12101 ( .A(n9643), .ZN(n9657) );
  NAND2_X1 U12102 ( .A1(n9713), .A2(n13332), .ZN(n9636) );
  NAND2_X1 U12103 ( .A1(n9749), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n9635) );
  NAND4_X1 U12104 ( .A1(n9638), .A2(n9637), .A3(n9636), .A4(n9635), .ZN(n13074) );
  NAND2_X1 U12105 ( .A1(n13074), .A2(n9737), .ZN(n9639) );
  NAND2_X1 U12106 ( .A1(n9640), .A2(n9639), .ZN(n9669) );
  NAND2_X1 U12107 ( .A1(n13585), .A2(n9743), .ZN(n9642) );
  OR2_X1 U12108 ( .A1(n9744), .A2(n13587), .ZN(n9641) );
  NAND2_X2 U12109 ( .A1(n9642), .A2(n9641), .ZN(n13476) );
  NAND2_X1 U12110 ( .A1(n9750), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9650) );
  NAND2_X1 U12111 ( .A1(n9749), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n9649) );
  INV_X1 U12112 ( .A(n9644), .ZN(n9659) );
  INV_X1 U12113 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9645) );
  NAND2_X1 U12114 ( .A1(n9659), .A2(n9645), .ZN(n9646) );
  NAND2_X1 U12115 ( .A1(n9713), .A2(n13303), .ZN(n9648) );
  NAND2_X1 U12116 ( .A1(n9656), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9647) );
  NAND4_X1 U12117 ( .A1(n9650), .A2(n9649), .A3(n9648), .A4(n9647), .ZN(n13256) );
  AND2_X1 U12118 ( .A1(n13256), .A2(n9737), .ZN(n9651) );
  AOI21_X1 U12119 ( .B1(n13476), .B2(n9718), .A(n9651), .ZN(n9727) );
  NAND2_X1 U12120 ( .A1(n13476), .A2(n9737), .ZN(n9653) );
  NAND2_X1 U12121 ( .A1(n13256), .A2(n9718), .ZN(n9652) );
  NAND2_X1 U12122 ( .A1(n9653), .A2(n9652), .ZN(n9726) );
  NAND2_X1 U12123 ( .A1(n9727), .A2(n9726), .ZN(n9731) );
  NAND2_X1 U12124 ( .A1(n13590), .A2(n9743), .ZN(n9655) );
  OR2_X1 U12125 ( .A1(n9744), .A2(n13593), .ZN(n9654) );
  NAND2_X2 U12126 ( .A1(n9655), .A2(n9654), .ZN(n13482) );
  NAND2_X1 U12127 ( .A1(n9656), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9663) );
  NAND2_X1 U12128 ( .A1(n9750), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9662) );
  INV_X1 U12129 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n12993) );
  NAND2_X1 U12130 ( .A1(n9657), .A2(n12993), .ZN(n9658) );
  NAND2_X1 U12131 ( .A1(n9713), .A2(n13314), .ZN(n9661) );
  NAND2_X1 U12132 ( .A1(n9749), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n9660) );
  NAND4_X1 U12133 ( .A1(n9663), .A2(n9662), .A3(n9661), .A4(n9660), .ZN(n13252) );
  AND2_X1 U12134 ( .A1(n13252), .A2(n9737), .ZN(n9664) );
  AOI21_X1 U12135 ( .B1(n13482), .B2(n9718), .A(n9664), .ZN(n9723) );
  NAND2_X1 U12136 ( .A1(n13482), .A2(n9737), .ZN(n9666) );
  NAND2_X1 U12137 ( .A1(n13252), .A2(n9718), .ZN(n9665) );
  NAND2_X1 U12138 ( .A1(n9666), .A2(n9665), .ZN(n9722) );
  NAND2_X1 U12139 ( .A1(n9723), .A2(n9722), .ZN(n9667) );
  OAI211_X1 U12140 ( .C1(n9670), .C2(n9669), .A(n9731), .B(n9667), .ZN(n9736)
         );
  AOI22_X1 U12141 ( .A1(n13488), .A2(n9737), .B1(n9718), .B2(n13074), .ZN(
        n9668) );
  AOI21_X1 U12142 ( .B1(n9670), .B2(n9669), .A(n9668), .ZN(n9735) );
  MUX2_X1 U12143 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9676), .Z(n9674) );
  XNOR2_X1 U12144 ( .A(n9674), .B(SI_30_), .ZN(n9740) );
  NAND2_X1 U12145 ( .A1(n9674), .A2(SI_30_), .ZN(n9675) );
  MUX2_X1 U12146 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9676), .Z(n9677) );
  XNOR2_X1 U12147 ( .A(n9677), .B(SI_31_), .ZN(n9678) );
  NAND2_X1 U12148 ( .A1(n11938), .A2(n9743), .ZN(n9681) );
  OR2_X1 U12149 ( .A1(n9744), .A2(n9972), .ZN(n9680) );
  INV_X1 U12150 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9684) );
  NAND2_X1 U12151 ( .A1(n9656), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9683) );
  NAND2_X1 U12152 ( .A1(n9750), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9682) );
  OAI211_X1 U12153 ( .C1(n9685), .C2(n9684), .A(n9683), .B(n9682), .ZN(n13200)
         );
  NAND2_X1 U12154 ( .A1(n13575), .A2(n9743), .ZN(n9687) );
  OR2_X1 U12155 ( .A1(n9744), .A2(n13576), .ZN(n9686) );
  NAND2_X1 U12156 ( .A1(n9656), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9692) );
  NAND2_X1 U12157 ( .A1(n9750), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9691) );
  NAND2_X1 U12158 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n9688) );
  NOR2_X1 U12159 ( .A1(n9712), .A2(n9688), .ZN(n13264) );
  NAND2_X1 U12160 ( .A1(n9713), .A2(n13264), .ZN(n9690) );
  NAND2_X1 U12161 ( .A1(n9749), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n9689) );
  NAND4_X1 U12162 ( .A1(n9692), .A2(n9691), .A3(n9690), .A4(n9689), .ZN(n13073) );
  AND2_X1 U12163 ( .A1(n13073), .A2(n9718), .ZN(n9693) );
  AOI21_X1 U12164 ( .B1(n13454), .B2(n9756), .A(n9693), .ZN(n9760) );
  NAND2_X1 U12165 ( .A1(n13454), .A2(n9718), .ZN(n9695) );
  NAND2_X1 U12166 ( .A1(n13073), .A2(n9737), .ZN(n9694) );
  NAND2_X1 U12167 ( .A1(n9695), .A2(n9694), .ZN(n9759) );
  NAND2_X1 U12168 ( .A1(n9760), .A2(n9759), .ZN(n9766) );
  NAND2_X1 U12169 ( .A1(n13578), .A2(n9743), .ZN(n9697) );
  OR2_X1 U12170 ( .A1(n9744), .A2(n15389), .ZN(n9696) );
  NAND2_X2 U12171 ( .A1(n9697), .A2(n9696), .ZN(n13282) );
  NAND2_X1 U12172 ( .A1(n9750), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9704) );
  NAND2_X1 U12173 ( .A1(n9749), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n9703) );
  INV_X1 U12174 ( .A(n13264), .ZN(n9700) );
  INV_X1 U12175 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n12944) );
  INV_X1 U12176 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9698) );
  OAI21_X1 U12177 ( .B1(n9712), .B2(n12944), .A(n9698), .ZN(n9699) );
  NAND2_X1 U12178 ( .A1(n9713), .A2(n12973), .ZN(n9702) );
  NAND2_X1 U12179 ( .A1(n9656), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9701) );
  NAND4_X1 U12180 ( .A1(n9704), .A2(n9703), .A3(n9702), .A4(n9701), .ZN(n13229) );
  AND2_X1 U12181 ( .A1(n13229), .A2(n9718), .ZN(n9705) );
  AOI21_X1 U12182 ( .B1(n13282), .B2(n9737), .A(n9705), .ZN(n9764) );
  NAND2_X1 U12183 ( .A1(n13282), .A2(n9718), .ZN(n9707) );
  NAND2_X1 U12184 ( .A1(n13229), .A2(n9737), .ZN(n9706) );
  NAND2_X1 U12185 ( .A1(n9707), .A2(n9706), .ZN(n9763) );
  NAND2_X1 U12186 ( .A1(n9764), .A2(n9763), .ZN(n9708) );
  AND2_X1 U12187 ( .A1(n9766), .A2(n9708), .ZN(n9709) );
  NAND2_X1 U12188 ( .A1(n13582), .A2(n9743), .ZN(n9711) );
  OR2_X1 U12189 ( .A1(n9744), .A2(n13583), .ZN(n9710) );
  NAND2_X1 U12190 ( .A1(n9656), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9717) );
  NAND2_X1 U12191 ( .A1(n9750), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9716) );
  XNOR2_X1 U12192 ( .A(n9712), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n13290) );
  NAND2_X1 U12193 ( .A1(n9713), .A2(n13290), .ZN(n9715) );
  NAND2_X1 U12194 ( .A1(n9749), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n9714) );
  NAND4_X1 U12195 ( .A1(n9717), .A2(n9716), .A3(n9715), .A4(n9714), .ZN(n13227) );
  AND2_X1 U12196 ( .A1(n13227), .A2(n9718), .ZN(n9719) );
  AOI21_X1 U12197 ( .B1(n13469), .B2(n9756), .A(n9719), .ZN(n9771) );
  NAND2_X1 U12198 ( .A1(n13469), .A2(n9718), .ZN(n9721) );
  NAND2_X1 U12199 ( .A1(n13227), .A2(n9737), .ZN(n9720) );
  NAND2_X1 U12200 ( .A1(n9721), .A2(n9720), .ZN(n9770) );
  NAND2_X1 U12201 ( .A1(n9771), .A2(n9770), .ZN(n9733) );
  INV_X1 U12202 ( .A(n9722), .ZN(n9725) );
  INV_X1 U12203 ( .A(n9723), .ZN(n9724) );
  AND2_X1 U12204 ( .A1(n9725), .A2(n9724), .ZN(n9730) );
  INV_X1 U12205 ( .A(n9726), .ZN(n9729) );
  INV_X1 U12206 ( .A(n9727), .ZN(n9728) );
  AOI22_X1 U12207 ( .A1(n9731), .A2(n9730), .B1(n9729), .B2(n9728), .ZN(n9732)
         );
  AND2_X1 U12208 ( .A1(n9733), .A2(n9732), .ZN(n9734) );
  MUX2_X1 U12209 ( .A(n13200), .B(n9293), .S(n13201), .Z(n9739) );
  NAND2_X1 U12210 ( .A1(n13200), .A2(n9737), .ZN(n9738) );
  NAND2_X1 U12211 ( .A1(n9739), .A2(n9738), .ZN(n9762) );
  INV_X1 U12212 ( .A(n9740), .ZN(n9741) );
  NAND2_X1 U12213 ( .A1(n13573), .A2(n9743), .ZN(n9746) );
  OR2_X1 U12214 ( .A1(n9744), .A2(n13574), .ZN(n9745) );
  INV_X1 U12215 ( .A(n11328), .ZN(n10202) );
  OAI211_X1 U12216 ( .C1(n10204), .C2(n10202), .A(n9747), .B(n9880), .ZN(n9748) );
  INV_X1 U12217 ( .A(n9748), .ZN(n9754) );
  NAND2_X1 U12218 ( .A1(n13200), .A2(n9718), .ZN(n9776) );
  NAND2_X1 U12219 ( .A1(n9749), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9753) );
  NAND2_X1 U12220 ( .A1(n9656), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9752) );
  NAND2_X1 U12221 ( .A1(n9750), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9751) );
  AOI21_X1 U12222 ( .B1(n9754), .B2(n9776), .A(n13231), .ZN(n9755) );
  AOI21_X1 U12223 ( .B1(n13204), .B2(n9756), .A(n9755), .ZN(n9775) );
  NAND2_X1 U12224 ( .A1(n13204), .A2(n9718), .ZN(n9758) );
  INV_X1 U12225 ( .A(n13231), .ZN(n13072) );
  NAND2_X1 U12226 ( .A1(n13072), .A2(n9756), .ZN(n9757) );
  NAND2_X1 U12227 ( .A1(n9758), .A2(n9757), .ZN(n9774) );
  OAI22_X1 U12228 ( .A1(n9775), .A2(n9774), .B1(n9760), .B2(n9759), .ZN(n9761)
         );
  INV_X1 U12229 ( .A(n9763), .ZN(n9767) );
  INV_X1 U12230 ( .A(n9764), .ZN(n9765) );
  MUX2_X1 U12231 ( .A(n13200), .B(n6526), .S(n13201), .Z(n9777) );
  NAND2_X1 U12232 ( .A1(n9777), .A2(n9776), .ZN(n9778) );
  XNOR2_X1 U12233 ( .A(n13204), .B(n13231), .ZN(n9800) );
  INV_X1 U12234 ( .A(n13073), .ZN(n12974) );
  XNOR2_X1 U12235 ( .A(n13454), .B(n12974), .ZN(n13260) );
  XNOR2_X1 U12236 ( .A(n13469), .B(n13258), .ZN(n13286) );
  NAND2_X1 U12237 ( .A1(n13282), .A2(n13229), .ZN(n13259) );
  OR2_X1 U12238 ( .A1(n13282), .A2(n13229), .ZN(n9779) );
  INV_X1 U12239 ( .A(n13256), .ZN(n13257) );
  XNOR2_X1 U12240 ( .A(n13476), .B(n13257), .ZN(n13298) );
  INV_X1 U12241 ( .A(n13252), .ZN(n13254) );
  XNOR2_X1 U12242 ( .A(n13482), .B(n13254), .ZN(n13319) );
  XNOR2_X1 U12243 ( .A(n13488), .B(n13251), .ZN(n13328) );
  OR2_X1 U12244 ( .A1(n13225), .A2(n13226), .ZN(n13249) );
  NAND2_X1 U12245 ( .A1(n13225), .A2(n13226), .ZN(n13250) );
  NAND2_X1 U12246 ( .A1(n13249), .A2(n13250), .ZN(n13340) );
  INV_X1 U12247 ( .A(n13245), .ZN(n13221) );
  XNOR2_X1 U12248 ( .A(n13387), .B(n13221), .ZN(n13220) );
  OR2_X1 U12249 ( .A1(n13518), .A2(n13075), .ZN(n13242) );
  NAND2_X1 U12250 ( .A1(n13518), .A2(n13075), .ZN(n13241) );
  NAND2_X1 U12251 ( .A1(n13242), .A2(n13241), .ZN(n13405) );
  XNOR2_X1 U12252 ( .A(n14573), .B(n14542), .ZN(n11725) );
  XNOR2_X1 U12253 ( .A(n11722), .B(n11721), .ZN(n11718) );
  INV_X1 U12254 ( .A(n13080), .ZN(n11612) );
  XNOR2_X1 U12255 ( .A(n15122), .B(n11612), .ZN(n11344) );
  XNOR2_X1 U12256 ( .A(n11465), .B(n11356), .ZN(n11259) );
  INV_X1 U12257 ( .A(n13082), .ZN(n11256) );
  XNOR2_X1 U12258 ( .A(n11274), .B(n11256), .ZN(n11252) );
  OR2_X1 U12259 ( .A1(n9780), .A2(n10637), .ZN(n10646) );
  NAND2_X1 U12260 ( .A1(n9780), .A2(n10637), .ZN(n9781) );
  NOR2_X1 U12261 ( .A1(n10636), .A2(n11328), .ZN(n9787) );
  NAND2_X1 U12262 ( .A1(n10327), .A2(n9783), .ZN(n15072) );
  INV_X1 U12263 ( .A(n15072), .ZN(n15086) );
  NAND4_X1 U12264 ( .A1(n9787), .A2(n15086), .A3(n10328), .A4(n10332), .ZN(
        n9788) );
  INV_X1 U12265 ( .A(n15105), .ZN(n10756) );
  XNOR2_X1 U12266 ( .A(n10756), .B(n13087), .ZN(n10661) );
  NOR3_X1 U12267 ( .A1(n9788), .A2(n10661), .A3(n10654), .ZN(n9789) );
  XNOR2_X1 U12268 ( .A(n15048), .B(n13085), .ZN(n10999) );
  NAND4_X1 U12269 ( .A1(n11131), .A2(n9789), .A3(n10999), .A4(n10994), .ZN(
        n9790) );
  OR4_X1 U12270 ( .A1(n11344), .A2(n11259), .A3(n11252), .A4(n9790), .ZN(n9791) );
  OR3_X1 U12271 ( .A1(n11725), .A2(n11718), .A3(n9791), .ZN(n9794) );
  INV_X1 U12272 ( .A(n13236), .ZN(n9792) );
  NAND2_X1 U12273 ( .A1(n13533), .A2(n9792), .ZN(n9793) );
  NAND2_X1 U12274 ( .A1(n13213), .A2(n9793), .ZN(n13429) );
  XNOR2_X1 U12275 ( .A(n14559), .B(n11881), .ZN(n14557) );
  INV_X1 U12276 ( .A(n13233), .ZN(n13210) );
  XNOR2_X1 U12277 ( .A(n13538), .B(n13210), .ZN(n11922) );
  XNOR2_X1 U12278 ( .A(n13424), .B(n13239), .ZN(n13238) );
  XNOR2_X1 U12279 ( .A(n13546), .B(n13076), .ZN(n11919) );
  NAND4_X1 U12280 ( .A1(n13405), .A2(n6546), .A3(n13238), .A4(n11919), .ZN(
        n9795) );
  NOR2_X1 U12281 ( .A1(n13220), .A2(n9795), .ZN(n9796) );
  XNOR2_X1 U12282 ( .A(n13375), .B(n13247), .ZN(n13370) );
  XNOR2_X1 U12283 ( .A(n13501), .B(n13248), .ZN(n13354) );
  NAND4_X1 U12284 ( .A1(n13340), .A2(n9796), .A3(n13370), .A4(n13354), .ZN(
        n9797) );
  OR4_X1 U12285 ( .A1(n13260), .A2(n13286), .A3(n13275), .A4(n9798), .ZN(n9799) );
  NOR2_X1 U12286 ( .A1(n9800), .A2(n9799), .ZN(n9801) );
  NAND2_X1 U12287 ( .A1(n9802), .A2(n9801), .ZN(n9808) );
  MUX2_X1 U12288 ( .A(n11439), .B(n9248), .S(n11328), .Z(n9803) );
  INV_X1 U12289 ( .A(n9804), .ZN(n9810) );
  OAI21_X1 U12290 ( .B1(n9550), .B2(n11439), .A(n9880), .ZN(n9805) );
  AOI21_X1 U12291 ( .B1(n9806), .B2(n9248), .A(n9805), .ZN(n9809) );
  NAND2_X1 U12292 ( .A1(n11439), .A2(n9247), .ZN(n9807) );
  OAI22_X1 U12293 ( .A1(n9810), .A2(n9809), .B1(n9808), .B2(n9807), .ZN(n9816)
         );
  OR2_X1 U12294 ( .A1(n9813), .A2(n9812), .ZN(n9814) );
  NAND2_X1 U12295 ( .A1(n9831), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11794) );
  INV_X1 U12296 ( .A(n11794), .ZN(n9815) );
  NAND2_X1 U12297 ( .A1(n6665), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9820) );
  NAND2_X1 U12298 ( .A1(n9821), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9822) );
  AND2_X1 U12299 ( .A1(n13586), .A2(n13591), .ZN(n9823) );
  NAND2_X1 U12300 ( .A1(n13595), .A2(n9823), .ZN(n9873) );
  INV_X1 U12301 ( .A(n15082), .ZN(n15084) );
  INV_X1 U12302 ( .A(n9825), .ZN(n9826) );
  NAND2_X1 U12303 ( .A1(n9826), .A2(n9997), .ZN(n14541) );
  OAI21_X1 U12304 ( .B1(n11794), .B2(n9834), .A(P2_B_REG_SCAN_IN), .ZN(n9827)
         );
  INV_X1 U12305 ( .A(n9827), .ZN(n9828) );
  NAND2_X1 U12306 ( .A1(n7770), .A2(n9828), .ZN(n9829) );
  NAND2_X1 U12307 ( .A1(n9830), .A2(n9829), .ZN(P2_U3328) );
  NOR2_X1 U12308 ( .A1(n9873), .A2(n9831), .ZN(n10000) );
  INV_X1 U12309 ( .A(n9958), .ZN(n9832) );
  INV_X2 U12310 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NAND2_X1 U12311 ( .A1(n9833), .A2(n10457), .ZN(n9837) );
  NAND2_X1 U12312 ( .A1(n15067), .A2(n12937), .ZN(n10499) );
  AND2_X1 U12313 ( .A1(n9782), .A2(n15089), .ZN(n10505) );
  NAND2_X1 U12314 ( .A1(n10505), .A2(n10457), .ZN(n14899) );
  INV_X1 U12315 ( .A(n9835), .ZN(n9836) );
  NAND2_X1 U12316 ( .A1(n9837), .A2(n9836), .ZN(n14907) );
  NAND2_X1 U12317 ( .A1(n14909), .A2(n14907), .ZN(n9838) );
  NAND2_X1 U12318 ( .A1(n9784), .A2(n10457), .ZN(n9841) );
  XNOR2_X1 U12319 ( .A(n9785), .B(n12968), .ZN(n9839) );
  XNOR2_X1 U12320 ( .A(n9841), .B(n9839), .ZN(n14906) );
  INV_X1 U12321 ( .A(n9839), .ZN(n9840) );
  NAND2_X1 U12322 ( .A1(n9841), .A2(n9840), .ZN(n9842) );
  AND2_X1 U12323 ( .A1(n9780), .A2(n10457), .ZN(n9843) );
  XNOR2_X1 U12324 ( .A(n10631), .B(n12968), .ZN(n10485) );
  NAND2_X1 U12325 ( .A1(n9843), .A2(n10485), .ZN(n10447) );
  INV_X1 U12326 ( .A(n9843), .ZN(n9845) );
  INV_X1 U12327 ( .A(n10485), .ZN(n9844) );
  NAND2_X1 U12328 ( .A1(n9845), .A2(n9844), .ZN(n9846) );
  NAND2_X1 U12329 ( .A1(n10447), .A2(n9846), .ZN(n9869) );
  NOR4_X1 U12330 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n9850) );
  NOR4_X1 U12331 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n9849) );
  NOR4_X1 U12332 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9848) );
  NOR4_X1 U12333 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n9847) );
  NAND4_X1 U12334 ( .A1(n9850), .A2(n9849), .A3(n9848), .A4(n9847), .ZN(n9858)
         );
  NOR2_X1 U12335 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n9854) );
  NOR4_X1 U12336 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n9853) );
  NOR4_X1 U12337 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n9852) );
  NOR4_X1 U12338 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9851) );
  NAND4_X1 U12339 ( .A1(n9854), .A2(n9853), .A3(n9852), .A4(n9851), .ZN(n9857)
         );
  XNOR2_X1 U12340 ( .A(n13595), .B(P2_B_REG_SCAN_IN), .ZN(n9855) );
  OR2_X1 U12341 ( .A1(n13591), .A2(n9855), .ZN(n9856) );
  OAI21_X1 U12342 ( .B1(n9858), .B2(n9857), .A(n15077), .ZN(n10210) );
  INV_X1 U12343 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9859) );
  NAND2_X1 U12344 ( .A1(n15077), .A2(n9859), .ZN(n9861) );
  OR2_X1 U12345 ( .A1(n13586), .A2(n13591), .ZN(n9860) );
  NAND2_X1 U12346 ( .A1(n9861), .A2(n9860), .ZN(n9872) );
  INV_X1 U12347 ( .A(n9872), .ZN(n10561) );
  AND2_X1 U12348 ( .A1(n15082), .A2(n10561), .ZN(n15083) );
  OR2_X1 U12349 ( .A1(n13595), .A2(n13586), .ZN(n9864) );
  INV_X1 U12350 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9862) );
  NAND2_X1 U12351 ( .A1(n15077), .A2(n9862), .ZN(n9863) );
  NAND2_X1 U12352 ( .A1(n9864), .A2(n9863), .ZN(n15081) );
  INV_X1 U12353 ( .A(n15081), .ZN(n10619) );
  AND2_X1 U12354 ( .A1(n15083), .A2(n10619), .ZN(n9865) );
  AND2_X1 U12355 ( .A1(n10210), .A2(n9865), .ZN(n9882) );
  NOR2_X1 U12356 ( .A1(n15123), .A2(n9997), .ZN(n9866) );
  INV_X1 U12357 ( .A(n10483), .ZN(n9868) );
  AOI211_X1 U12358 ( .C1(n9870), .C2(n9869), .A(n14903), .B(n9868), .ZN(n9887)
         );
  NAND2_X1 U12359 ( .A1(n10210), .A2(n10619), .ZN(n9871) );
  NAND2_X1 U12360 ( .A1(n9871), .A2(n9877), .ZN(n9875) );
  NAND2_X1 U12361 ( .A1(n9877), .A2(n9872), .ZN(n10618) );
  NAND2_X1 U12362 ( .A1(n9997), .A2(n9880), .ZN(n10208) );
  AND4_X1 U12363 ( .A1(n10618), .A2(n9873), .A3(n9996), .A4(n10208), .ZN(n9874) );
  NAND2_X1 U12364 ( .A1(n9875), .A2(n9874), .ZN(n10500) );
  INV_X1 U12365 ( .A(n14551), .ZN(n13007) );
  MUX2_X1 U12366 ( .A(n13007), .B(P2_U3088), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n9886) );
  NAND2_X1 U12367 ( .A1(n15090), .A2(n10202), .ZN(n15066) );
  INV_X1 U12368 ( .A(n15066), .ZN(n9876) );
  NAND2_X1 U12369 ( .A1(n9882), .A2(n9876), .ZN(n9879) );
  INV_X1 U12370 ( .A(n9880), .ZN(n9881) );
  INV_X1 U12371 ( .A(n14914), .ZN(n13038) );
  NAND2_X1 U12372 ( .A1(n9784), .A2(n13049), .ZN(n9884) );
  AND2_X2 U12373 ( .A1(n9997), .A2(n9825), .ZN(n13198) );
  NAND2_X1 U12374 ( .A1(n13088), .A2(n13198), .ZN(n9883) );
  AND2_X1 U12375 ( .A1(n9884), .A2(n9883), .ZN(n10627) );
  OAI22_X1 U12376 ( .A1(n10637), .A2(n12998), .B1(n13038), .B2(n10627), .ZN(
        n9885) );
  OR3_X1 U12377 ( .A1(n9887), .A2(n9886), .A3(n9885), .ZN(P2_U3190) );
  NOR2_X1 U12378 ( .A1(n9676), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12889) );
  INV_X1 U12379 ( .A(n9888), .ZN(n9890) );
  NAND2_X2 U12380 ( .A1(n9676), .A2(P3_U3151), .ZN(n12900) );
  OAI222_X1 U12381 ( .A1(n12903), .A2(n9890), .B1(n12900), .B2(n9889), .C1(
        P3_U3151), .C2(n10780), .ZN(P3_U3289) );
  INV_X1 U12382 ( .A(n9891), .ZN(n9893) );
  OAI222_X1 U12383 ( .A1(n12903), .A2(n9893), .B1(n12900), .B2(n9892), .C1(
        P3_U3151), .C2(n10382), .ZN(P3_U3294) );
  INV_X1 U12384 ( .A(SI_5_), .ZN(n9894) );
  OAI222_X1 U12385 ( .A1(n7218), .A2(P3_U3151), .B1(n12903), .B2(n9895), .C1(
        n9894), .C2(n12900), .ZN(P3_U3290) );
  INV_X2 U12386 ( .A(n11792), .ZN(n13597) );
  NOR2_X1 U12387 ( .A1(n9676), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13580) );
  INV_X2 U12388 ( .A(n13580), .ZN(n13599) );
  OAI222_X1 U12389 ( .A1(n13597), .A2(n9930), .B1(n10006), .B2(P2_U3088), .C1(
        n9896), .C2(n13599), .ZN(P2_U3326) );
  INV_X1 U12390 ( .A(n9897), .ZN(n9899) );
  OAI222_X1 U12391 ( .A1(n12903), .A2(n9899), .B1(n12900), .B2(n9898), .C1(
        P3_U3151), .C2(n11406), .ZN(P3_U3287) );
  NOR2_X1 U12392 ( .A1(n9676), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14322) );
  OAI222_X1 U12393 ( .A1(n14347), .A2(n9900), .B1(n14327), .B2(n9902), .C1(
        n10087), .C2(P1_U3086), .ZN(P1_U3352) );
  OAI222_X1 U12394 ( .A1(n14347), .A2(n9901), .B1(n14327), .B2(n9906), .C1(
        n10310), .C2(P1_U3086), .ZN(P1_U3353) );
  OAI222_X1 U12395 ( .A1(n13599), .A2(n9903), .B1(n13103), .B2(P2_U3088), .C1(
        n13597), .C2(n9902), .ZN(P2_U3324) );
  OAI222_X1 U12396 ( .A1(n13599), .A2(n9904), .B1(n10012), .B2(P2_U3088), .C1(
        n13597), .C2(n9912), .ZN(P2_U3323) );
  OAI222_X1 U12397 ( .A1(n13597), .A2(n9906), .B1(n14929), .B2(P2_U3088), .C1(
        n9905), .C2(n13599), .ZN(P2_U3325) );
  INV_X1 U12398 ( .A(SI_10_), .ZN(n9908) );
  OAI222_X1 U12399 ( .A1(P3_U3151), .A2(n11587), .B1(n12900), .B2(n9908), .C1(
        n12903), .C2(n9907), .ZN(P3_U3285) );
  INV_X1 U12400 ( .A(SI_7_), .ZN(n9910) );
  OAI222_X1 U12401 ( .A1(P3_U3151), .A2(n11159), .B1(n12900), .B2(n9910), .C1(
        n12903), .C2(n9909), .ZN(P3_U3288) );
  INV_X1 U12402 ( .A(n13132), .ZN(n9911) );
  OAI222_X1 U12403 ( .A1(n13599), .A2(n6881), .B1(n9911), .B2(P2_U3088), .C1(
        n13597), .C2(n9916), .ZN(P2_U3322) );
  OAI222_X1 U12404 ( .A1(n14347), .A2(n7062), .B1(n14327), .B2(n9912), .C1(
        n10321), .C2(P1_U3086), .ZN(P1_U3351) );
  INV_X1 U12405 ( .A(SI_9_), .ZN(n9914) );
  OAI222_X1 U12406 ( .A1(P3_U3151), .A2(n11403), .B1(n12900), .B2(n9914), .C1(
        n9913), .C2(n12903), .ZN(P3_U3286) );
  INV_X1 U12407 ( .A(n10124), .ZN(n9915) );
  OAI222_X1 U12408 ( .A1(n14347), .A2(n9917), .B1(n14327), .B2(n9916), .C1(
        n9915), .C2(P1_U3086), .ZN(P1_U3350) );
  OAI222_X1 U12409 ( .A1(P3_U3151), .A2(n11762), .B1(n12900), .B2(n9919), .C1(
        n12903), .C2(n9918), .ZN(P3_U3284) );
  INV_X1 U12410 ( .A(SI_4_), .ZN(n9920) );
  OAI222_X1 U12411 ( .A1(n10412), .A2(P3_U3151), .B1(n12903), .B2(n9921), .C1(
        n9920), .C2(n12900), .ZN(P3_U3291) );
  INV_X1 U12412 ( .A(n10406), .ZN(n10390) );
  INV_X1 U12413 ( .A(SI_2_), .ZN(n9922) );
  OAI222_X1 U12414 ( .A1(n10390), .A2(P3_U3151), .B1(n12903), .B2(n9923), .C1(
        n9922), .C2(n12900), .ZN(P3_U3293) );
  INV_X1 U12415 ( .A(SI_3_), .ZN(n9924) );
  OAI222_X1 U12416 ( .A1(n10409), .A2(P3_U3151), .B1(n12903), .B2(n9925), .C1(
        n9924), .C2(n12900), .ZN(P3_U3292) );
  OAI222_X1 U12417 ( .A1(n14347), .A2(n9926), .B1(n14327), .B2(n9927), .C1(
        n10121), .C2(P1_U3086), .ZN(P1_U3349) );
  INV_X1 U12418 ( .A(n13144), .ZN(n9928) );
  OAI222_X1 U12419 ( .A1(n13599), .A2(n6883), .B1(n9928), .B2(P2_U3088), .C1(
        n13597), .C2(n9927), .ZN(P2_U3321) );
  OAI222_X1 U12420 ( .A1(P1_U3086), .A2(n10156), .B1(n14327), .B2(n9930), .C1(
        n9929), .C2(n14347), .ZN(P1_U3354) );
  INV_X1 U12421 ( .A(n9931), .ZN(n9932) );
  OAI222_X1 U12422 ( .A1(n12900), .A2(n9933), .B1(n12903), .B2(n9932), .C1(
        n12382), .C2(P3_U3151), .ZN(P3_U3283) );
  INV_X1 U12423 ( .A(n14347), .ZN(n10424) );
  AOI22_X1 U12424 ( .A1(n10164), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10424), .ZN(n9934) );
  OAI21_X1 U12425 ( .B1(n9935), .B2(n14327), .A(n9934), .ZN(P1_U3348) );
  INV_X1 U12426 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9937) );
  INV_X1 U12427 ( .A(n13156), .ZN(n9936) );
  OAI222_X1 U12428 ( .A1(n13599), .A2(n9937), .B1(n9936), .B2(P2_U3088), .C1(
        n13597), .C2(n9935), .ZN(P2_U3320) );
  AOI22_X1 U12429 ( .A1(n10287), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10424), .ZN(n9938) );
  OAI21_X1 U12430 ( .B1(n9939), .B2(n14327), .A(n9938), .ZN(P1_U3347) );
  INV_X1 U12431 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9940) );
  INV_X1 U12432 ( .A(n10018), .ZN(n14941) );
  OAI222_X1 U12433 ( .A1(n13599), .A2(n9940), .B1(n14941), .B2(P2_U3088), .C1(
        n13597), .C2(n9939), .ZN(P2_U3319) );
  AOI22_X1 U12434 ( .A1(n10474), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n10424), .ZN(n9941) );
  OAI21_X1 U12435 ( .B1(n9945), .B2(n14327), .A(n9941), .ZN(P1_U3346) );
  INV_X1 U12436 ( .A(n9942), .ZN(n9943) );
  OAI222_X1 U12437 ( .A1(n12900), .A2(n9944), .B1(n12903), .B2(n9943), .C1(
        P3_U3151), .C2(n12388), .ZN(P3_U3282) );
  INV_X1 U12438 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9946) );
  INV_X1 U12439 ( .A(n10020), .ZN(n14946) );
  OAI222_X1 U12440 ( .A1(n13599), .A2(n9946), .B1(n14946), .B2(P2_U3088), .C1(
        n13597), .C2(n9945), .ZN(P2_U3318) );
  OAI222_X1 U12441 ( .A1(P3_U3151), .A2(n12436), .B1(n12900), .B2(n9948), .C1(
        n12903), .C2(n9947), .ZN(P3_U3281) );
  OR2_X1 U12442 ( .A1(n10175), .A2(P1_U3086), .ZN(n12157) );
  INV_X1 U12443 ( .A(n12157), .ZN(n9949) );
  OR2_X1 U12444 ( .A1(n10192), .A2(n9949), .ZN(n10075) );
  AOI21_X1 U12445 ( .B1(n11943), .B2(n10175), .A(n9950), .ZN(n10074) );
  INV_X1 U12446 ( .A(n10074), .ZN(n9951) );
  AND2_X1 U12447 ( .A1(n10075), .A2(n9951), .ZN(n14673) );
  NOR2_X1 U12448 ( .A1(n14673), .A2(P1_U4016), .ZN(P1_U3085) );
  AOI22_X1 U12449 ( .A1(n11033), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10424), .ZN(n9952) );
  OAI21_X1 U12450 ( .B1(n9961), .B2(n14327), .A(n9952), .ZN(P1_U3345) );
  NAND2_X2 U12451 ( .A1(n10192), .A2(n9953), .ZN(n14855) );
  INV_X1 U12452 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9956) );
  INV_X1 U12453 ( .A(n9954), .ZN(n9955) );
  AOI22_X1 U12454 ( .A1(n14855), .A2(n9956), .B1(n9958), .B2(n9955), .ZN(
        P1_U3446) );
  INV_X1 U12455 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9960) );
  INV_X1 U12456 ( .A(n9957), .ZN(n9959) );
  AOI22_X1 U12457 ( .A1(n14855), .A2(n9960), .B1(n9959), .B2(n9958), .ZN(
        P1_U3445) );
  INV_X1 U12458 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9963) );
  INV_X1 U12459 ( .A(n14973), .ZN(n9962) );
  OAI222_X1 U12460 ( .A1(n13599), .A2(n9963), .B1(n9962), .B2(P2_U3088), .C1(
        n13597), .C2(n9961), .ZN(P2_U3317) );
  INV_X1 U12461 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9965) );
  NAND2_X1 U12462 ( .A1(P1_U4016), .A2(n10342), .ZN(n9964) );
  OAI21_X1 U12463 ( .B1(P1_U4016), .B2(n9965), .A(n9964), .ZN(P1_U3560) );
  NAND2_X1 U12464 ( .A1(n6475), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n9970) );
  NAND2_X1 U12465 ( .A1(n9966), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9969) );
  NAND2_X1 U12466 ( .A1(n9967), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9968) );
  NAND3_X1 U12467 ( .A1(n9970), .A2(n9969), .A3(n9968), .ZN(n13935) );
  NAND2_X1 U12468 ( .A1(P1_U4016), .A2(n13935), .ZN(n9971) );
  OAI21_X1 U12469 ( .B1(P1_U4016), .B2(n9972), .A(n9971), .ZN(P1_U3591) );
  INV_X1 U12470 ( .A(n9973), .ZN(n10031) );
  AOI22_X1 U12471 ( .A1(n14680), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10424), .ZN(n9974) );
  OAI21_X1 U12472 ( .B1(n10031), .B2(n14327), .A(n9974), .ZN(P1_U3344) );
  INV_X1 U12473 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n9975) );
  MUX2_X1 U12474 ( .A(n9975), .B(P2_REG2_REG_11__SCAN_IN), .S(n10241), .Z(
        n9995) );
  XNOR2_X1 U12475 ( .A(n10006), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n13096) );
  AND2_X1 U12476 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n13095) );
  NAND2_X1 U12477 ( .A1(n13096), .A2(n13095), .ZN(n13094) );
  INV_X1 U12478 ( .A(n10006), .ZN(n13093) );
  NAND2_X1 U12479 ( .A1(n13093), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9976) );
  NAND2_X1 U12480 ( .A1(n13094), .A2(n9976), .ZN(n14925) );
  XNOR2_X1 U12481 ( .A(n14929), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n14926) );
  NAND2_X1 U12482 ( .A1(n14925), .A2(n14926), .ZN(n14924) );
  INV_X1 U12483 ( .A(n14929), .ZN(n10008) );
  NAND2_X1 U12484 ( .A1(n10008), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9977) );
  NAND2_X1 U12485 ( .A1(n14924), .A2(n9977), .ZN(n13112) );
  XNOR2_X1 U12486 ( .A(n13103), .B(P2_REG2_REG_3__SCAN_IN), .ZN(n13113) );
  NAND2_X1 U12487 ( .A1(n13112), .A2(n13113), .ZN(n13111) );
  INV_X1 U12488 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9978) );
  OR2_X1 U12489 ( .A1(n13103), .A2(n9978), .ZN(n9979) );
  NAND2_X1 U12490 ( .A1(n13111), .A2(n9979), .ZN(n13124) );
  XNOR2_X1 U12491 ( .A(n10012), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n13125) );
  NAND2_X1 U12492 ( .A1(n13124), .A2(n13125), .ZN(n13123) );
  INV_X1 U12493 ( .A(n10012), .ZN(n13119) );
  NAND2_X1 U12494 ( .A1(n13119), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9980) );
  NAND2_X1 U12495 ( .A1(n13123), .A2(n9980), .ZN(n13137) );
  INV_X1 U12496 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9981) );
  XNOR2_X1 U12497 ( .A(n13132), .B(n9981), .ZN(n13138) );
  NAND2_X1 U12498 ( .A1(n13137), .A2(n13138), .ZN(n13136) );
  NAND2_X1 U12499 ( .A1(n13132), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9982) );
  NAND2_X1 U12500 ( .A1(n13136), .A2(n9982), .ZN(n13149) );
  INV_X1 U12501 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n9983) );
  MUX2_X1 U12502 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n9983), .S(n13144), .Z(
        n13150) );
  NAND2_X1 U12503 ( .A1(n13149), .A2(n13150), .ZN(n13148) );
  NAND2_X1 U12504 ( .A1(n13144), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9984) );
  NAND2_X1 U12505 ( .A1(n13148), .A2(n9984), .ZN(n13158) );
  INV_X1 U12506 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9985) );
  MUX2_X1 U12507 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9985), .S(n13156), .Z(
        n13159) );
  NAND2_X1 U12508 ( .A1(n13158), .A2(n13159), .ZN(n13157) );
  NAND2_X1 U12509 ( .A1(n13156), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9986) );
  NAND2_X1 U12510 ( .A1(n13157), .A2(n9986), .ZN(n14937) );
  INV_X1 U12511 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9987) );
  XNOR2_X1 U12512 ( .A(n10018), .B(n9987), .ZN(n14938) );
  NAND2_X1 U12513 ( .A1(n14937), .A2(n14938), .ZN(n14936) );
  NAND2_X1 U12514 ( .A1(n10018), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9988) );
  NAND2_X1 U12515 ( .A1(n14936), .A2(n9988), .ZN(n14951) );
  XNOR2_X1 U12516 ( .A(n10020), .B(P2_REG2_REG_9__SCAN_IN), .ZN(n14952) );
  OR2_X1 U12517 ( .A1(n14951), .A2(n14952), .ZN(n14949) );
  INV_X1 U12518 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9989) );
  NAND2_X1 U12519 ( .A1(n14946), .A2(n9989), .ZN(n9990) );
  NAND2_X1 U12520 ( .A1(n14949), .A2(n9990), .ZN(n14969) );
  INV_X1 U12521 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9991) );
  MUX2_X1 U12522 ( .A(n9991), .B(P2_REG2_REG_10__SCAN_IN), .S(n14973), .Z(
        n14970) );
  OR2_X1 U12523 ( .A1(n14969), .A2(n14970), .ZN(n14967) );
  NAND2_X1 U12524 ( .A1(n14973), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9992) );
  NAND2_X1 U12525 ( .A1(n14967), .A2(n9992), .ZN(n9994) );
  INV_X1 U12526 ( .A(n10237), .ZN(n9993) );
  AOI21_X1 U12527 ( .B1(n9995), .B2(n9994), .A(n9993), .ZN(n10029) );
  NAND2_X1 U12528 ( .A1(n9997), .A2(n9996), .ZN(n9998) );
  AND2_X1 U12529 ( .A1(n9290), .A2(n9998), .ZN(n9999) );
  OR2_X1 U12530 ( .A1(n10000), .A2(n9999), .ZN(n10002) );
  NOR2_X1 U12531 ( .A1(n9825), .A2(P2_U3088), .ZN(n13579) );
  NAND2_X1 U12532 ( .A1(n10002), .A2(n13579), .ZN(n10024) );
  INV_X1 U12533 ( .A(n10024), .ZN(n10001) );
  INV_X1 U12534 ( .A(n13584), .ZN(n13196) );
  AND2_X1 U12535 ( .A1(n10001), .A2(n13196), .ZN(n15043) );
  NAND2_X1 U12536 ( .A1(n10002), .A2(n9825), .ZN(n14947) );
  INV_X1 U12537 ( .A(n10241), .ZN(n10030) );
  INV_X1 U12538 ( .A(n15046), .ZN(n14920) );
  NAND2_X1 U12539 ( .A1(n14920), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n10004) );
  NAND2_X1 U12540 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n10003)
         );
  OAI211_X1 U12541 ( .C1(n15037), .C2(n10030), .A(n10004), .B(n10003), .ZN(
        n10005) );
  INV_X1 U12542 ( .A(n10005), .ZN(n10028) );
  XNOR2_X1 U12543 ( .A(n10006), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n13099) );
  AND2_X1 U12544 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n13098) );
  NAND2_X1 U12545 ( .A1(n13099), .A2(n13098), .ZN(n13097) );
  NAND2_X1 U12546 ( .A1(n13093), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10007) );
  NAND2_X1 U12547 ( .A1(n13097), .A2(n10007), .ZN(n14922) );
  XNOR2_X1 U12548 ( .A(n14929), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n14923) );
  NAND2_X1 U12549 ( .A1(n14922), .A2(n14923), .ZN(n14921) );
  NAND2_X1 U12550 ( .A1(n10008), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10009) );
  NAND2_X1 U12551 ( .A1(n14921), .A2(n10009), .ZN(n13109) );
  XNOR2_X1 U12552 ( .A(n13103), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n13110) );
  NAND2_X1 U12553 ( .A1(n13109), .A2(n13110), .ZN(n13108) );
  INV_X1 U12554 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10010) );
  OR2_X1 U12555 ( .A1(n13103), .A2(n10010), .ZN(n10011) );
  NAND2_X1 U12556 ( .A1(n13108), .A2(n10011), .ZN(n13121) );
  XNOR2_X1 U12557 ( .A(n10012), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n13122) );
  NAND2_X1 U12558 ( .A1(n13121), .A2(n13122), .ZN(n13120) );
  NAND2_X1 U12559 ( .A1(n13119), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10013) );
  NAND2_X1 U12560 ( .A1(n13120), .A2(n10013), .ZN(n13134) );
  INV_X1 U12561 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10014) );
  XNOR2_X1 U12562 ( .A(n13132), .B(n10014), .ZN(n13135) );
  NAND2_X1 U12563 ( .A1(n13134), .A2(n13135), .ZN(n13133) );
  NAND2_X1 U12564 ( .A1(n13132), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10015) );
  NAND2_X1 U12565 ( .A1(n13133), .A2(n10015), .ZN(n13146) );
  INV_X1 U12566 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10764) );
  MUX2_X1 U12567 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10764), .S(n13144), .Z(
        n13147) );
  NAND2_X1 U12568 ( .A1(n13146), .A2(n13147), .ZN(n13145) );
  NAND2_X1 U12569 ( .A1(n13144), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10016) );
  NAND2_X1 U12570 ( .A1(n13145), .A2(n10016), .ZN(n13161) );
  INV_X1 U12571 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n11007) );
  MUX2_X1 U12572 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n11007), .S(n13156), .Z(
        n13162) );
  NAND2_X1 U12573 ( .A1(n13161), .A2(n13162), .ZN(n13160) );
  NAND2_X1 U12574 ( .A1(n13156), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10017) );
  NAND2_X1 U12575 ( .A1(n13160), .A2(n10017), .ZN(n14934) );
  INV_X1 U12576 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n15140) );
  MUX2_X1 U12577 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n15140), .S(n10018), .Z(
        n14935) );
  NAND2_X1 U12578 ( .A1(n14934), .A2(n14935), .ZN(n14933) );
  NAND2_X1 U12579 ( .A1(n10018), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10019) );
  NAND2_X1 U12580 ( .A1(n14933), .A2(n10019), .ZN(n14955) );
  INV_X1 U12581 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n11279) );
  MUX2_X1 U12582 ( .A(n11279), .B(P2_REG1_REG_9__SCAN_IN), .S(n10020), .Z(
        n14956) );
  OR2_X1 U12583 ( .A1(n14955), .A2(n14956), .ZN(n14953) );
  NAND2_X1 U12584 ( .A1(n14946), .A2(n11279), .ZN(n10021) );
  NAND2_X1 U12585 ( .A1(n14953), .A2(n10021), .ZN(n14965) );
  INV_X1 U12586 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10022) );
  MUX2_X1 U12587 ( .A(n10022), .B(P2_REG1_REG_10__SCAN_IN), .S(n14973), .Z(
        n14966) );
  OR2_X1 U12588 ( .A1(n14965), .A2(n14966), .ZN(n14963) );
  NAND2_X1 U12589 ( .A1(n14973), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10023) );
  NAND2_X1 U12590 ( .A1(n14963), .A2(n10023), .ZN(n10026) );
  INV_X1 U12591 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n15143) );
  MUX2_X1 U12592 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n15143), .S(n10241), .Z(
        n10025) );
  NAND2_X1 U12593 ( .A1(n10026), .A2(n10025), .ZN(n10243) );
  OR2_X1 U12594 ( .A1(n10024), .A2(n13196), .ZN(n15022) );
  OAI211_X1 U12595 ( .C1(n10026), .C2(n10025), .A(n10243), .B(n15035), .ZN(
        n10027) );
  OAI211_X1 U12596 ( .C1(n10029), .C2(n15008), .A(n10028), .B(n10027), .ZN(
        P2_U3225) );
  INV_X1 U12597 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10032) );
  OAI222_X1 U12598 ( .A1(n13599), .A2(n10032), .B1(n13597), .B2(n10031), .C1(
        P2_U3088), .C2(n10030), .ZN(P2_U3316) );
  NOR2_X1 U12599 ( .A1(n10033), .A2(n12881), .ZN(n10035) );
  INV_X1 U12600 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10034) );
  NOR2_X1 U12601 ( .A1(n10051), .A2(n10034), .ZN(P3_U3262) );
  CLKBUF_X1 U12602 ( .A(n10035), .Z(n10051) );
  INV_X1 U12603 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10036) );
  NOR2_X1 U12604 ( .A1(n10051), .A2(n10036), .ZN(P3_U3263) );
  INV_X1 U12605 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10037) );
  NOR2_X1 U12606 ( .A1(n10051), .A2(n10037), .ZN(P3_U3261) );
  INV_X1 U12607 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10038) );
  NOR2_X1 U12608 ( .A1(n10035), .A2(n10038), .ZN(P3_U3260) );
  INV_X1 U12609 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10039) );
  NOR2_X1 U12610 ( .A1(n10051), .A2(n10039), .ZN(P3_U3259) );
  INV_X1 U12611 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10040) );
  NOR2_X1 U12612 ( .A1(n10035), .A2(n10040), .ZN(P3_U3258) );
  INV_X1 U12613 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10041) );
  NOR2_X1 U12614 ( .A1(n10051), .A2(n10041), .ZN(P3_U3257) );
  INV_X1 U12615 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10042) );
  NOR2_X1 U12616 ( .A1(n10051), .A2(n10042), .ZN(P3_U3256) );
  INV_X1 U12617 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10043) );
  NOR2_X1 U12618 ( .A1(n10051), .A2(n10043), .ZN(P3_U3255) );
  INV_X1 U12619 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10044) );
  NOR2_X1 U12620 ( .A1(n10051), .A2(n10044), .ZN(P3_U3254) );
  INV_X1 U12621 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n15283) );
  NOR2_X1 U12622 ( .A1(n10051), .A2(n15283), .ZN(P3_U3253) );
  INV_X1 U12623 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10045) );
  NOR2_X1 U12624 ( .A1(n10051), .A2(n10045), .ZN(P3_U3252) );
  INV_X1 U12625 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n15401) );
  NOR2_X1 U12626 ( .A1(n10051), .A2(n15401), .ZN(P3_U3251) );
  INV_X1 U12627 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10046) );
  NOR2_X1 U12628 ( .A1(n10051), .A2(n10046), .ZN(P3_U3250) );
  INV_X1 U12629 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n15427) );
  NOR2_X1 U12630 ( .A1(n10051), .A2(n15427), .ZN(P3_U3249) );
  INV_X1 U12631 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10047) );
  NOR2_X1 U12632 ( .A1(n10051), .A2(n10047), .ZN(P3_U3248) );
  INV_X1 U12633 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10048) );
  NOR2_X1 U12634 ( .A1(n10035), .A2(n10048), .ZN(P3_U3240) );
  INV_X1 U12635 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10049) );
  NOR2_X1 U12636 ( .A1(n10051), .A2(n10049), .ZN(P3_U3247) );
  INV_X1 U12637 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10050) );
  NOR2_X1 U12638 ( .A1(n10051), .A2(n10050), .ZN(P3_U3246) );
  INV_X1 U12639 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10052) );
  NOR2_X1 U12640 ( .A1(n10035), .A2(n10052), .ZN(P3_U3245) );
  INV_X1 U12641 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10053) );
  NOR2_X1 U12642 ( .A1(n10035), .A2(n10053), .ZN(P3_U3244) );
  INV_X1 U12643 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10054) );
  NOR2_X1 U12644 ( .A1(n10035), .A2(n10054), .ZN(P3_U3243) );
  INV_X1 U12645 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10055) );
  NOR2_X1 U12646 ( .A1(n10035), .A2(n10055), .ZN(P3_U3242) );
  INV_X1 U12647 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10056) );
  NOR2_X1 U12648 ( .A1(n10035), .A2(n10056), .ZN(P3_U3241) );
  INV_X1 U12649 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10057) );
  NOR2_X1 U12650 ( .A1(n10035), .A2(n10057), .ZN(P3_U3234) );
  INV_X1 U12651 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10058) );
  NOR2_X1 U12652 ( .A1(n10035), .A2(n10058), .ZN(P3_U3239) );
  INV_X1 U12653 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10059) );
  NOR2_X1 U12654 ( .A1(n10035), .A2(n10059), .ZN(P3_U3238) );
  INV_X1 U12655 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10060) );
  NOR2_X1 U12656 ( .A1(n10051), .A2(n10060), .ZN(P3_U3237) );
  INV_X1 U12657 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n15290) );
  NOR2_X1 U12658 ( .A1(n10051), .A2(n15290), .ZN(P3_U3236) );
  INV_X1 U12659 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10061) );
  NOR2_X1 U12660 ( .A1(n10051), .A2(n10061), .ZN(P3_U3235) );
  INV_X1 U12661 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10062) );
  NAND2_X1 U12662 ( .A1(n15043), .A2(n10062), .ZN(n10063) );
  OAI211_X1 U12663 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n15022), .A(n10063), .B(
        n15037), .ZN(n10065) );
  INV_X1 U12664 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n15135) );
  OAI22_X1 U12665 ( .A1(n15008), .A2(n10062), .B1(n15135), .B2(n15022), .ZN(
        n10064) );
  MUX2_X1 U12666 ( .A(n10065), .B(n10064), .S(n7397), .Z(n10067) );
  INV_X1 U12667 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15448) );
  INV_X1 U12668 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n15069) );
  OAI22_X1 U12669 ( .A1(n15046), .A2(n15448), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15069), .ZN(n10066) );
  OR2_X1 U12670 ( .A1(n10067), .A2(n10066), .ZN(P2_U3214) );
  INV_X1 U12671 ( .A(n10068), .ZN(n10069) );
  OAI222_X1 U12672 ( .A1(P3_U3151), .A2(n12440), .B1(n12900), .B2(n15386), 
        .C1(n12903), .C2(n10069), .ZN(P3_U3280) );
  OAI222_X1 U12673 ( .A1(n12900), .A2(n10071), .B1(n12903), .B2(n10070), .C1(
        P3_U3151), .C2(n12483), .ZN(P3_U3279) );
  INV_X1 U12674 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n15256) );
  NAND2_X1 U12675 ( .A1(n10960), .A2(P3_U3897), .ZN(n10072) );
  OAI21_X1 U12676 ( .B1(P3_U3897), .B2(n15256), .A(n10072), .ZN(P3_U3494) );
  INV_X1 U12677 ( .A(n10073), .ZN(n10101) );
  INV_X1 U12678 ( .A(n13913), .ZN(n11030) );
  OAI222_X1 U12679 ( .A1(n14347), .A2(n7533), .B1(n14327), .B2(n10101), .C1(
        n11030), .C2(P1_U3086), .ZN(P1_U3343) );
  NAND2_X1 U12680 ( .A1(n10075), .A2(n10074), .ZN(n14675) );
  INV_X1 U12681 ( .A(n6487), .ZN(n14671) );
  XOR2_X1 U12682 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10124), .Z(n10080) );
  INV_X1 U12683 ( .A(n10087), .ZN(n10103) );
  INV_X1 U12684 ( .A(n10310), .ZN(n10086) );
  AND3_X1 U12685 ( .A1(n10146), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG1_REG_0__SCAN_IN), .ZN(n10147) );
  AOI21_X1 U12686 ( .B1(n10084), .B2(P1_REG1_REG_1__SCAN_IN), .A(n10147), .ZN(
        n10308) );
  INV_X1 U12687 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10076) );
  MUX2_X1 U12688 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10076), .S(n10310), .Z(
        n10307) );
  NOR2_X1 U12689 ( .A1(n10308), .A2(n10307), .ZN(n10306) );
  INV_X1 U12690 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10077) );
  MUX2_X1 U12691 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10077), .S(n10087), .Z(
        n10108) );
  NOR2_X1 U12692 ( .A1(n10109), .A2(n10108), .ZN(n10107) );
  INV_X1 U12693 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10078) );
  MUX2_X1 U12694 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10078), .S(n10321), .Z(
        n10315) );
  NOR2_X1 U12695 ( .A1(n10316), .A2(n10315), .ZN(n10314) );
  AOI21_X1 U12696 ( .B1(n10092), .B2(P1_REG1_REG_4__SCAN_IN), .A(n10314), .ZN(
        n10079) );
  NAND2_X1 U12697 ( .A1(n10079), .A2(n10080), .ZN(n10123) );
  OAI21_X1 U12698 ( .B1(n10080), .B2(n10079), .A(n10123), .ZN(n10099) );
  INV_X1 U12699 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10083) );
  NAND2_X1 U12700 ( .A1(n14778), .A2(n10124), .ZN(n10082) );
  NAND2_X1 U12701 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n10081) );
  OAI211_X1 U12702 ( .C1(n10083), .C2(n14781), .A(n10082), .B(n10081), .ZN(
        n10098) );
  NAND2_X1 U12703 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10296) );
  NOR2_X1 U12704 ( .A1(n10151), .A2(n10296), .ZN(n10150) );
  AOI21_X1 U12705 ( .B1(n10084), .B2(P1_REG2_REG_1__SCAN_IN), .A(n10150), .ZN(
        n10305) );
  INV_X1 U12706 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10085) );
  MUX2_X1 U12707 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10085), .S(n10310), .Z(
        n10304) );
  NOR2_X1 U12708 ( .A1(n10305), .A2(n10304), .ZN(n10303) );
  AOI21_X1 U12709 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n10086), .A(n10303), .ZN(
        n10112) );
  INV_X1 U12710 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10088) );
  MUX2_X1 U12711 ( .A(n10088), .B(P1_REG2_REG_3__SCAN_IN), .S(n10087), .Z(
        n10089) );
  INV_X1 U12712 ( .A(n10089), .ZN(n10111) );
  NOR2_X1 U12713 ( .A1(n10112), .A2(n10111), .ZN(n10110) );
  AOI21_X1 U12714 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n10103), .A(n10110), .ZN(
        n10319) );
  INV_X1 U12715 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10090) );
  MUX2_X1 U12716 ( .A(n10090), .B(P1_REG2_REG_4__SCAN_IN), .S(n10321), .Z(
        n10091) );
  INV_X1 U12717 ( .A(n10091), .ZN(n10318) );
  NOR2_X1 U12718 ( .A1(n10319), .A2(n10318), .ZN(n10317) );
  AOI21_X1 U12719 ( .B1(n10092), .B2(P1_REG2_REG_4__SCAN_IN), .A(n10317), .ZN(
        n10096) );
  XNOR2_X1 U12720 ( .A(n10124), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n10095) );
  INV_X1 U12721 ( .A(n14675), .ZN(n10094) );
  NOR2_X1 U12722 ( .A1(n14331), .A2(n6487), .ZN(n10093) );
  NOR2_X1 U12723 ( .A1(n10096), .A2(n10095), .ZN(n10116) );
  AOI211_X1 U12724 ( .C1(n10096), .C2(n10095), .A(n14767), .B(n10116), .ZN(
        n10097) );
  AOI211_X1 U12725 ( .C1(n14749), .C2(n10099), .A(n10098), .B(n10097), .ZN(
        n10100) );
  INV_X1 U12726 ( .A(n10100), .ZN(P1_U3248) );
  INV_X1 U12727 ( .A(n10244), .ZN(n14981) );
  OAI222_X1 U12728 ( .A1(n13599), .A2(n10102), .B1(n14981), .B2(P2_U3088), 
        .C1(n13597), .C2(n10101), .ZN(P2_U3315) );
  INV_X1 U12729 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10106) );
  NAND2_X1 U12730 ( .A1(n14778), .A2(n10103), .ZN(n10105) );
  NAND2_X1 U12731 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n10104) );
  OAI211_X1 U12732 ( .C1(n10106), .C2(n14781), .A(n10105), .B(n10104), .ZN(
        n10115) );
  AOI211_X1 U12733 ( .C1(n10109), .C2(n10108), .A(n10107), .B(n14772), .ZN(
        n10114) );
  AOI211_X1 U12734 ( .C1(n10112), .C2(n10111), .A(n10110), .B(n14767), .ZN(
        n10113) );
  OR3_X1 U12735 ( .A1(n10115), .A2(n10114), .A3(n10113), .ZN(P1_U3246) );
  AOI21_X1 U12736 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n10124), .A(n10116), .ZN(
        n10120) );
  INV_X1 U12737 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10117) );
  MUX2_X1 U12738 ( .A(n10117), .B(P1_REG2_REG_6__SCAN_IN), .S(n10121), .Z(
        n10118) );
  INV_X1 U12739 ( .A(n10118), .ZN(n10119) );
  NOR2_X1 U12740 ( .A1(n10120), .A2(n10119), .ZN(n10132) );
  AOI211_X1 U12741 ( .C1(n10120), .C2(n10119), .A(n14767), .B(n10132), .ZN(
        n10131) );
  INV_X1 U12742 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10122) );
  MUX2_X1 U12743 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10122), .S(n10121), .Z(
        n10126) );
  AOI211_X1 U12744 ( .C1(n10126), .C2(n10125), .A(n14772), .B(n10136), .ZN(
        n10130) );
  INV_X1 U12745 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14362) );
  NAND2_X1 U12746 ( .A1(n14778), .A2(n10137), .ZN(n10128) );
  NAND2_X1 U12747 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n10127) );
  OAI211_X1 U12748 ( .C1(n14362), .C2(n14781), .A(n10128), .B(n10127), .ZN(
        n10129) );
  OR3_X1 U12749 ( .A1(n10131), .A2(n10130), .A3(n10129), .ZN(P1_U3249) );
  INV_X1 U12750 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10133) );
  MUX2_X1 U12751 ( .A(n10133), .B(P1_REG2_REG_7__SCAN_IN), .S(n10164), .Z(
        n10134) );
  AOI211_X1 U12752 ( .C1(n10135), .C2(n10134), .A(n14767), .B(n10163), .ZN(
        n10145) );
  INV_X1 U12753 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10138) );
  MUX2_X1 U12754 ( .A(n10138), .B(P1_REG1_REG_7__SCAN_IN), .S(n10164), .Z(
        n10139) );
  NOR2_X1 U12755 ( .A1(n10140), .A2(n10139), .ZN(n10157) );
  AOI211_X1 U12756 ( .C1(n10140), .C2(n10139), .A(n14772), .B(n10157), .ZN(
        n10144) );
  INV_X1 U12757 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14366) );
  NAND2_X1 U12758 ( .A1(n14778), .A2(n10164), .ZN(n10142) );
  NAND2_X1 U12759 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n10141) );
  OAI211_X1 U12760 ( .C1(n14366), .C2(n14781), .A(n10142), .B(n10141), .ZN(
        n10143) );
  OR3_X1 U12761 ( .A1(n10145), .A2(n10144), .A3(n10143), .ZN(P1_U3250) );
  INV_X1 U12762 ( .A(n14778), .ZN(n14752) );
  NAND2_X1 U12763 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n10149) );
  INV_X1 U12764 ( .A(n10146), .ZN(n10148) );
  AOI211_X1 U12765 ( .C1(n10149), .C2(n10148), .A(n10147), .B(n14772), .ZN(
        n10153) );
  AOI211_X1 U12766 ( .C1(n10296), .C2(n10151), .A(n10150), .B(n14767), .ZN(
        n10152) );
  NOR2_X1 U12767 ( .A1(n10153), .A2(n10152), .ZN(n10155) );
  AOI22_X1 U12768 ( .A1(n14673), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n10154) );
  OAI211_X1 U12769 ( .C1(n10156), .C2(n14752), .A(n10155), .B(n10154), .ZN(
        P1_U3244) );
  INV_X1 U12770 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10158) );
  MUX2_X1 U12771 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10158), .S(n10287), .Z(
        n10159) );
  NAND2_X1 U12772 ( .A1(n10160), .A2(n10159), .ZN(n10281) );
  OAI21_X1 U12773 ( .B1(n10160), .B2(n10159), .A(n10281), .ZN(n10170) );
  INV_X1 U12774 ( .A(n10287), .ZN(n10162) );
  AND2_X1 U12775 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11522) );
  AOI21_X1 U12776 ( .B1(n14673), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n11522), .ZN(
        n10161) );
  OAI21_X1 U12777 ( .B1(n14752), .B2(n10162), .A(n10161), .ZN(n10169) );
  INV_X1 U12778 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10165) );
  MUX2_X1 U12779 ( .A(n10165), .B(P1_REG2_REG_8__SCAN_IN), .S(n10287), .Z(
        n10166) );
  AOI211_X1 U12780 ( .C1(n10167), .C2(n10166), .A(n14767), .B(n10286), .ZN(
        n10168) );
  AOI211_X1 U12781 ( .C1(n14749), .C2(n10170), .A(n10169), .B(n10168), .ZN(
        n10171) );
  INV_X1 U12782 ( .A(n10171), .ZN(P1_U3251) );
  AND2_X1 U12783 ( .A1(n10256), .A2(n10850), .ZN(n10197) );
  NAND2_X1 U12784 ( .A1(n10197), .A2(n10172), .ZN(n10174) );
  NAND2_X1 U12785 ( .A1(n10174), .A2(n10173), .ZN(n10181) );
  AND3_X1 U12786 ( .A1(n10185), .A2(n10176), .A3(n10175), .ZN(n12154) );
  NAND2_X1 U12787 ( .A1(n10181), .A2(n12154), .ZN(n10791) );
  NOR2_X1 U12788 ( .A1(n10791), .A2(P1_U3086), .ZN(n10279) );
  INV_X1 U12789 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10882) );
  NAND2_X1 U12790 ( .A1(n10192), .A2(n10178), .ZN(n10179) );
  NAND2_X1 U12791 ( .A1(n14831), .A2(n10179), .ZN(n10180) );
  AND2_X1 U12792 ( .A1(n13897), .A2(n14149), .ZN(n10885) );
  AOI22_X1 U12793 ( .A1(n14621), .A2(n10259), .B1(n14625), .B2(n10885), .ZN(
        n10199) );
  INV_X1 U12794 ( .A(n13615), .ZN(n10184) );
  INV_X1 U12795 ( .A(n10185), .ZN(n10188) );
  AOI22_X1 U12796 ( .A1(n10220), .A2(n10259), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n10188), .ZN(n10186) );
  NAND2_X1 U12797 ( .A1(n10188), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10189) );
  OAI211_X1 U12798 ( .C1(n13687), .C2(n10888), .A(n10190), .B(n10189), .ZN(
        n10222) );
  XNOR2_X1 U12799 ( .A(n10221), .B(n10222), .ZN(n10297) );
  NAND2_X1 U12800 ( .A1(n10192), .A2(n10191), .ZN(n10195) );
  INV_X1 U12801 ( .A(n11943), .ZN(n10193) );
  NAND2_X1 U12802 ( .A1(n14872), .A2(n10193), .ZN(n10194) );
  AOI21_X1 U12803 ( .B1(n14855), .B2(n10195), .A(n10194), .ZN(n10196) );
  NAND2_X1 U12804 ( .A1(n10297), .A2(n14623), .ZN(n10198) );
  OAI211_X1 U12805 ( .C1(n10279), .C2(n10882), .A(n10199), .B(n10198), .ZN(
        P1_U3232) );
  NOR2_X1 U12806 ( .A1(n9247), .A2(n10202), .ZN(n10201) );
  NAND2_X1 U12807 ( .A1(n10201), .A2(n9248), .ZN(n15107) );
  XOR2_X1 U12808 ( .A(n10505), .B(n10328), .Z(n10564) );
  AOI21_X1 U12809 ( .B1(n10200), .B2(n15107), .A(n10564), .ZN(n10207) );
  XNOR2_X1 U12810 ( .A(n10328), .B(n10327), .ZN(n10205) );
  NAND2_X1 U12811 ( .A1(n9747), .A2(n10202), .ZN(n10203) );
  AOI22_X1 U12812 ( .A1(n13049), .A2(n9782), .B1(n9784), .B2(n13198), .ZN(
        n10501) );
  OAI21_X1 U12813 ( .B1(n10205), .B2(n15127), .A(n10501), .ZN(n10563) );
  NOR3_X1 U12814 ( .A1(n10207), .A2(n10563), .A3(n10206), .ZN(n15093) );
  AND2_X1 U12815 ( .A1(n15082), .A2(n10208), .ZN(n10209) );
  AND2_X1 U12816 ( .A1(n10210), .A2(n10209), .ZN(n10621) );
  NOR2_X1 U12817 ( .A1(n10618), .A2(n15081), .ZN(n10211) );
  NAND2_X1 U12818 ( .A1(n15142), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10212) );
  OAI21_X1 U12819 ( .B1(n15093), .B2(n15142), .A(n10212), .ZN(P2_U3500) );
  INV_X1 U12820 ( .A(n10213), .ZN(n10232) );
  INV_X1 U12821 ( .A(n14699), .ZN(n10214) );
  OAI222_X1 U12822 ( .A1(n14347), .A2(n10215), .B1(n14327), .B2(n10232), .C1(
        n10214), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U12823 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10231) );
  NAND2_X1 U12824 ( .A1(n10342), .A2(n13861), .ZN(n10346) );
  INV_X1 U12825 ( .A(n14149), .ZN(n13806) );
  NOR2_X1 U12826 ( .A1(n10267), .A2(n13806), .ZN(n10348) );
  INV_X1 U12827 ( .A(n10348), .ZN(n10216) );
  AOI21_X1 U12828 ( .B1(n10346), .B2(n10216), .A(n13846), .ZN(n10217) );
  AOI21_X1 U12829 ( .B1(n14621), .B2(n7060), .A(n10217), .ZN(n10230) );
  XNOR2_X1 U12830 ( .A(n10269), .B(n10268), .ZN(n10227) );
  NAND2_X1 U12831 ( .A1(n10225), .A2(n10224), .ZN(n10226) );
  OAI21_X1 U12832 ( .B1(n10227), .B2(n10226), .A(n10272), .ZN(n10228) );
  NAND2_X1 U12833 ( .A1(n10228), .A2(n14623), .ZN(n10229) );
  OAI211_X1 U12834 ( .C1(n10279), .C2(n10231), .A(n10230), .B(n10229), .ZN(
        P1_U3222) );
  INV_X1 U12835 ( .A(n10583), .ZN(n10249) );
  OAI222_X1 U12836 ( .A1(n13599), .A2(n10233), .B1(n10249), .B2(P2_U3088), 
        .C1(n13597), .C2(n10232), .ZN(P2_U3314) );
  INV_X1 U12837 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10234) );
  MUX2_X1 U12838 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n10234), .S(n10583), .Z(
        n10235) );
  INV_X1 U12839 ( .A(n10235), .ZN(n10239) );
  OR2_X1 U12840 ( .A1(n10241), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10236) );
  XNOR2_X1 U12841 ( .A(n10244), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n14984) );
  OAI22_X1 U12842 ( .A1(n14985), .A2(n14984), .B1(n10244), .B2(
        P2_REG2_REG_12__SCAN_IN), .ZN(n10238) );
  NOR2_X1 U12843 ( .A1(n10238), .A2(n10239), .ZN(n10577) );
  AOI211_X1 U12844 ( .C1(n10239), .C2(n10238), .A(n15008), .B(n10577), .ZN(
        n10252) );
  INV_X1 U12845 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10240) );
  MUX2_X1 U12846 ( .A(n10240), .B(P2_REG1_REG_13__SCAN_IN), .S(n10583), .Z(
        n10246) );
  NAND2_X1 U12847 ( .A1(n10241), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10242) );
  NAND2_X1 U12848 ( .A1(n10243), .A2(n10242), .ZN(n14978) );
  INV_X1 U12849 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14587) );
  MUX2_X1 U12850 ( .A(n14587), .B(P2_REG1_REG_12__SCAN_IN), .S(n10244), .Z(
        n14977) );
  OAI21_X1 U12851 ( .B1(n10244), .B2(P2_REG1_REG_12__SCAN_IN), .A(n14980), 
        .ZN(n10245) );
  NOR2_X1 U12852 ( .A1(n10245), .A2(n10246), .ZN(n10582) );
  AOI211_X1 U12853 ( .C1(n10246), .C2(n10245), .A(n15022), .B(n10582), .ZN(
        n10251) );
  NAND2_X1 U12854 ( .A1(n14920), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n10248) );
  NAND2_X1 U12855 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n10247)
         );
  OAI211_X1 U12856 ( .C1(n15037), .C2(n10249), .A(n10248), .B(n10247), .ZN(
        n10250) );
  OR3_X1 U12857 ( .A1(n10252), .A2(n10251), .A3(n10250), .ZN(P2_U3227) );
  INV_X1 U12858 ( .A(n10253), .ZN(n10254) );
  OAI222_X1 U12859 ( .A1(P3_U3151), .A2(n12509), .B1(n12900), .B2(n10255), 
        .C1(n12903), .C2(n10254), .ZN(P3_U3278) );
  AND2_X1 U12860 ( .A1(n10342), .A2(n10888), .ZN(n10258) );
  OAI21_X1 U12861 ( .B1(n14887), .B2(n14269), .A(n12118), .ZN(n10263) );
  AND2_X1 U12862 ( .A1(n10259), .A2(n10260), .ZN(n10261) );
  NOR2_X1 U12863 ( .A1(n10885), .A2(n10261), .ZN(n10262) );
  AND2_X1 U12864 ( .A1(n10263), .A2(n10262), .ZN(n14857) );
  NAND2_X1 U12865 ( .A1(n14894), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10264) );
  OAI21_X1 U12866 ( .B1(n14894), .B2(n14857), .A(n10264), .ZN(P1_U3528) );
  INV_X1 U12867 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14830) );
  NAND2_X1 U12868 ( .A1(n10220), .A2(n13895), .ZN(n10265) );
  OAI22_X1 U12869 ( .A1(n13615), .A2(n10267), .B1(n14861), .B2(n13686), .ZN(
        n10793) );
  XNOR2_X1 U12870 ( .A(n10794), .B(n10793), .ZN(n10274) );
  INV_X1 U12871 ( .A(n10268), .ZN(n10270) );
  NAND2_X1 U12872 ( .A1(n10270), .A2(n10269), .ZN(n10271) );
  OAI21_X1 U12873 ( .B1(n10274), .B2(n10273), .A(n10797), .ZN(n10275) );
  NAND2_X1 U12874 ( .A1(n10275), .A2(n14623), .ZN(n10278) );
  OAI22_X1 U12875 ( .A1(n10341), .A2(n13804), .B1(n10801), .B2(n13806), .ZN(
        n14829) );
  AOI22_X1 U12876 ( .A1(n14621), .A2(n10276), .B1(n14625), .B2(n14829), .ZN(
        n10277) );
  OAI211_X1 U12877 ( .C1(n10279), .C2(n14830), .A(n10278), .B(n10277), .ZN(
        P1_U3237) );
  INV_X1 U12878 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10280) );
  MUX2_X1 U12879 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10280), .S(n10474), .Z(
        n10283) );
  OAI21_X1 U12880 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n10287), .A(n10281), .ZN(
        n10282) );
  NAND2_X1 U12881 ( .A1(n10282), .A2(n10283), .ZN(n10473) );
  OAI21_X1 U12882 ( .B1(n10283), .B2(n10282), .A(n10473), .ZN(n10294) );
  INV_X1 U12883 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14371) );
  NAND2_X1 U12884 ( .A1(n14778), .A2(n10474), .ZN(n10285) );
  NAND2_X1 U12885 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n10284) );
  OAI211_X1 U12886 ( .C1(n14371), .C2(n14781), .A(n10285), .B(n10284), .ZN(
        n10293) );
  AOI21_X1 U12887 ( .B1(n10287), .B2(P1_REG2_REG_8__SCAN_IN), .A(n10286), .ZN(
        n10291) );
  INV_X1 U12888 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10288) );
  MUX2_X1 U12889 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10288), .S(n10474), .Z(
        n10289) );
  INV_X1 U12890 ( .A(n10289), .ZN(n10290) );
  NOR2_X1 U12891 ( .A1(n10291), .A2(n10290), .ZN(n10468) );
  AOI211_X1 U12892 ( .C1(n10291), .C2(n10290), .A(n14767), .B(n10468), .ZN(
        n10292) );
  AOI211_X1 U12893 ( .C1(n14749), .C2(n10294), .A(n10293), .B(n10292), .ZN(
        n10295) );
  INV_X1 U12894 ( .A(n10295), .ZN(P1_U3252) );
  INV_X1 U12895 ( .A(n10296), .ZN(n10299) );
  INV_X1 U12896 ( .A(n10297), .ZN(n10298) );
  MUX2_X1 U12897 ( .A(n10299), .B(n10298), .S(n6487), .Z(n10302) );
  INV_X1 U12898 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10883) );
  AOI21_X1 U12899 ( .B1(n14671), .B2(n10883), .A(n14331), .ZN(n14670) );
  OAI21_X1 U12900 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n14670), .A(P1_U4016), .ZN(
        n10300) );
  AOI21_X1 U12901 ( .B1(n10302), .B2(n10301), .A(n10300), .ZN(n10325) );
  AOI211_X1 U12902 ( .C1(n10305), .C2(n10304), .A(n10303), .B(n14767), .ZN(
        n10313) );
  AOI211_X1 U12903 ( .C1(n10308), .C2(n10307), .A(n10306), .B(n14772), .ZN(
        n10312) );
  AOI22_X1 U12904 ( .A1(n14673), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n10309) );
  OAI21_X1 U12905 ( .B1(n14752), .B2(n10310), .A(n10309), .ZN(n10311) );
  OR4_X1 U12906 ( .A1(n10325), .A2(n10313), .A3(n10312), .A4(n10311), .ZN(
        P1_U3245) );
  AOI211_X1 U12907 ( .C1(n10316), .C2(n10315), .A(n10314), .B(n14772), .ZN(
        n10324) );
  AOI211_X1 U12908 ( .C1(n10319), .C2(n10318), .A(n10317), .B(n14767), .ZN(
        n10323) );
  NAND2_X1 U12909 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10814) );
  NAND2_X1 U12910 ( .A1(n14673), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n10320) );
  OAI211_X1 U12911 ( .C1(n14752), .C2(n10321), .A(n10814), .B(n10320), .ZN(
        n10322) );
  OR4_X1 U12912 ( .A1(n10325), .A2(n10324), .A3(n10323), .A4(n10322), .ZN(
        P1_U3247) );
  INV_X1 U12913 ( .A(n9833), .ZN(n10334) );
  INV_X1 U12914 ( .A(n14576), .ZN(n14570) );
  INV_X1 U12915 ( .A(n10327), .ZN(n10329) );
  NAND2_X1 U12916 ( .A1(n10329), .A2(n10328), .ZN(n10331) );
  NAND2_X1 U12917 ( .A1(n10334), .A2(n10502), .ZN(n10330) );
  NAND2_X1 U12918 ( .A1(n10333), .A2(n10332), .ZN(n10433) );
  OAI21_X1 U12919 ( .B1(n10333), .B2(n10332), .A(n10433), .ZN(n10335) );
  INV_X1 U12920 ( .A(n9780), .ZN(n10638) );
  OAI22_X1 U12921 ( .A1(n10334), .A2(n14541), .B1(n10638), .B2(n14539), .ZN(
        n14915) );
  AOI21_X1 U12922 ( .B1(n10335), .B2(n14579), .A(n14915), .ZN(n10704) );
  OAI211_X1 U12923 ( .C1(n7184), .C2(n9786), .A(n14562), .B(n10437), .ZN(
        n10698) );
  OAI211_X1 U12924 ( .C1(n9786), .C2(n15114), .A(n10704), .B(n10698), .ZN(
        n10337) );
  AOI21_X1 U12925 ( .B1(n10701), .B2(n14570), .A(n10337), .ZN(n15095) );
  NAND2_X1 U12926 ( .A1(n15142), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10338) );
  OAI21_X1 U12927 ( .B1(n15095), .B2(n15142), .A(n10338), .ZN(P2_U3501) );
  INV_X1 U12928 ( .A(n14868), .ZN(n14866) );
  XNOR2_X1 U12929 ( .A(n12117), .B(n10339), .ZN(n14850) );
  OAI21_X1 U12930 ( .B1(n10888), .B2(n14844), .A(n14835), .ZN(n10340) );
  OR2_X1 U12931 ( .A1(n10340), .A2(n10182), .ZN(n14847) );
  OAI21_X1 U12932 ( .B1(n14844), .B2(n14872), .A(n14847), .ZN(n10350) );
  INV_X1 U12933 ( .A(n11427), .ZN(n14877) );
  XNOR2_X1 U12934 ( .A(n10341), .B(n10340), .ZN(n10344) );
  NOR2_X1 U12935 ( .A1(n12117), .A2(n13861), .ZN(n10343) );
  MUX2_X1 U12936 ( .A(n10344), .B(n10343), .S(n10342), .Z(n10345) );
  AOI21_X1 U12937 ( .B1(n14885), .B2(n10346), .A(n10345), .ZN(n10347) );
  AOI211_X1 U12938 ( .C1(n14877), .C2(n14850), .A(n10348), .B(n10347), .ZN(
        n14854) );
  INV_X1 U12939 ( .A(n14854), .ZN(n10349) );
  AOI211_X1 U12940 ( .C1(n14866), .C2(n14850), .A(n10350), .B(n10349), .ZN(
        n14859) );
  NAND2_X1 U12941 ( .A1(n14894), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10351) );
  OAI21_X1 U12942 ( .B1(n14859), .B2(n14894), .A(n10351), .ZN(P1_U3529) );
  INV_X1 U12943 ( .A(n10352), .ZN(n10353) );
  OAI222_X1 U12944 ( .A1(P3_U3151), .A2(n12520), .B1(n12900), .B2(n10354), 
        .C1(n12903), .C2(n10353), .ZN(P3_U3277) );
  INV_X2 U12945 ( .A(P3_U3897), .ZN(n12375) );
  INV_X1 U12946 ( .A(n10688), .ZN(n10355) );
  NAND2_X1 U12947 ( .A1(n10355), .A2(n11303), .ZN(n10373) );
  NAND2_X1 U12948 ( .A1(n8307), .A2(n10672), .ZN(n10357) );
  NAND2_X1 U12949 ( .A1(n10357), .A2(n10356), .ZN(n10372) );
  INV_X1 U12950 ( .A(n10372), .ZN(n10358) );
  NAND2_X1 U12951 ( .A1(n10373), .A2(n10358), .ZN(n10365) );
  MUX2_X1 U12952 ( .A(n12375), .B(n10365), .S(n8450), .Z(n15147) );
  INV_X1 U12953 ( .A(n15162), .ZN(n12431) );
  XNOR2_X1 U12954 ( .A(n10406), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n10364) );
  NAND2_X1 U12955 ( .A1(n7016), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10362) );
  INV_X1 U12956 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15212) );
  NAND2_X1 U12957 ( .A1(n10533), .A2(n10362), .ZN(n10363) );
  NAND2_X1 U12958 ( .A1(n10364), .A2(n10363), .ZN(n10408) );
  OAI21_X1 U12959 ( .B1(n10364), .B2(n10363), .A(n10408), .ZN(n10377) );
  INV_X1 U12960 ( .A(n10365), .ZN(n10366) );
  NAND2_X1 U12961 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n7522), .ZN(n10367) );
  OR2_X1 U12962 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10367), .ZN(n10368) );
  OAI21_X1 U12963 ( .B1(n10370), .B2(n10369), .A(n10401), .ZN(n10371) );
  AND2_X1 U12964 ( .A1(n12547), .A2(n10371), .ZN(n10376) );
  INV_X1 U12965 ( .A(n15168), .ZN(n15156) );
  INV_X1 U12966 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10374) );
  OAI22_X1 U12967 ( .A1(n15156), .A2(n10374), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10733), .ZN(n10375) );
  AOI211_X1 U12968 ( .C1(n12431), .C2(n10377), .A(n10376), .B(n10375), .ZN(
        n10388) );
  MUX2_X1 U12969 ( .A(n15212), .B(n10378), .S(n12539), .Z(n10383) );
  XNOR2_X1 U12970 ( .A(n10383), .B(n10382), .ZN(n10530) );
  OR2_X1 U12971 ( .A1(n12539), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10381) );
  NAND2_X1 U12972 ( .A1(n12539), .A2(n7791), .ZN(n10380) );
  NAND2_X1 U12973 ( .A1(n10381), .A2(n10380), .ZN(n15149) );
  INV_X1 U12974 ( .A(n10382), .ZN(n10542) );
  AOI22_X1 U12975 ( .A1(n10530), .A2(n15153), .B1(n10542), .B2(n10383), .ZN(
        n10392) );
  OR2_X1 U12976 ( .A1(n12539), .A2(n10405), .ZN(n10385) );
  NAND2_X1 U12977 ( .A1(n12539), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10384) );
  NAND2_X1 U12978 ( .A1(n10385), .A2(n10384), .ZN(n10389) );
  XOR2_X1 U12979 ( .A(n10406), .B(n10389), .Z(n10391) );
  XNOR2_X1 U12980 ( .A(n10392), .B(n10391), .ZN(n10386) );
  NAND2_X1 U12981 ( .A1(P3_U3897), .A2(n8450), .ZN(n15150) );
  NAND2_X1 U12982 ( .A1(n10386), .A2(n15173), .ZN(n10387) );
  OAI211_X1 U12983 ( .C1(n15147), .C2(n10390), .A(n10388), .B(n10387), .ZN(
        P3_U3184) );
  OAI22_X1 U12984 ( .A1(n10392), .A2(n10391), .B1(n10390), .B2(n10389), .ZN(
        n10545) );
  MUX2_X1 U12985 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12539), .Z(n10393) );
  XNOR2_X1 U12986 ( .A(n10393), .B(n10558), .ZN(n10546) );
  INV_X1 U12987 ( .A(n10393), .ZN(n10394) );
  MUX2_X1 U12988 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12539), .Z(n10395) );
  XNOR2_X1 U12989 ( .A(n10395), .B(n10412), .ZN(n10513) );
  MUX2_X1 U12990 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12539), .Z(n10592) );
  XNOR2_X1 U12991 ( .A(n10592), .B(n10413), .ZN(n10396) );
  NAND2_X1 U12992 ( .A1(n10396), .A2(n10397), .ZN(n10593) );
  OAI21_X1 U12993 ( .B1(n10397), .B2(n10396), .A(n10593), .ZN(n10398) );
  NAND2_X1 U12994 ( .A1(n10398), .A2(n15173), .ZN(n10422) );
  OR2_X1 U12995 ( .A1(n10406), .A2(n10399), .ZN(n10400) );
  NAND2_X1 U12996 ( .A1(n10401), .A2(n10400), .ZN(n10402) );
  NAND2_X1 U12997 ( .A1(n10402), .A2(n10409), .ZN(n10514) );
  OR2_X1 U12998 ( .A1(n10402), .A2(n10409), .ZN(n10403) );
  XNOR2_X1 U12999 ( .A(n10412), .B(P3_REG1_REG_4__SCAN_IN), .ZN(n10515) );
  NOR2_X1 U13000 ( .A1(n10404), .A2(n10413), .ZN(n10602) );
  OAI21_X1 U13001 ( .B1(n6673), .B2(P3_REG1_REG_5__SCAN_IN), .A(n6523), .ZN(
        n10420) );
  OR2_X1 U13002 ( .A1(n10406), .A2(n10405), .ZN(n10407) );
  NAND2_X1 U13003 ( .A1(n10408), .A2(n10407), .ZN(n10410) );
  NAND2_X1 U13004 ( .A1(n10410), .A2(n10409), .ZN(n10518) );
  OR2_X1 U13005 ( .A1(n10410), .A2(n10409), .ZN(n10411) );
  NAND2_X1 U13006 ( .A1(n10518), .A2(n10411), .ZN(n10551) );
  XNOR2_X1 U13007 ( .A(n10412), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n10519) );
  NOR2_X1 U13008 ( .A1(n7863), .A2(n10415), .ZN(n10597) );
  AOI21_X1 U13009 ( .B1(n10415), .B2(n7863), .A(n10597), .ZN(n10418) );
  NOR2_X1 U13010 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10416), .ZN(n11214) );
  AOI21_X1 U13011 ( .B1(n15168), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11214), .ZN(
        n10417) );
  OAI21_X1 U13012 ( .B1(n10418), .B2(n15162), .A(n10417), .ZN(n10419) );
  AOI21_X1 U13013 ( .B1(n12547), .B2(n10420), .A(n10419), .ZN(n10421) );
  OAI211_X1 U13014 ( .C1(n15147), .C2(n7218), .A(n10422), .B(n10421), .ZN(
        P3_U3187) );
  INV_X1 U13015 ( .A(n10423), .ZN(n10444) );
  AOI22_X1 U13016 ( .A1(n14708), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n10424), .ZN(n10425) );
  OAI21_X1 U13017 ( .B1(n10444), .B2(n14327), .A(n10425), .ZN(P1_U3341) );
  OAI222_X1 U13018 ( .A1(n12903), .A2(n10427), .B1(n12900), .B2(n10426), .C1(
        P3_U3151), .C2(n12545), .ZN(P3_U3276) );
  INV_X1 U13019 ( .A(n9784), .ZN(n10431) );
  NAND2_X1 U13020 ( .A1(n10431), .A2(n9786), .ZN(n10429) );
  NAND2_X1 U13021 ( .A1(n10430), .A2(n10429), .ZN(n10635) );
  INV_X1 U13022 ( .A(n10636), .ZN(n10435) );
  XNOR2_X1 U13023 ( .A(n10635), .B(n10435), .ZN(n10634) );
  NAND2_X1 U13024 ( .A1(n10431), .A2(n9785), .ZN(n10432) );
  OAI21_X1 U13025 ( .B1(n10435), .B2(n10434), .A(n10647), .ZN(n10436) );
  AND2_X1 U13026 ( .A1(n10436), .A2(n14579), .ZN(n10630) );
  NAND2_X1 U13027 ( .A1(n10437), .A2(n10631), .ZN(n10438) );
  NAND2_X1 U13028 ( .A1(n10438), .A2(n14562), .ZN(n10439) );
  NOR2_X1 U13029 ( .A1(n10641), .A2(n10439), .ZN(n10625) );
  OAI21_X1 U13030 ( .B1(n10637), .B2(n15114), .A(n10627), .ZN(n10440) );
  NOR3_X1 U13031 ( .A1(n10630), .A2(n10625), .A3(n10440), .ZN(n10441) );
  OAI21_X1 U13032 ( .B1(n14576), .B2(n10634), .A(n10441), .ZN(n10622) );
  NAND2_X1 U13033 ( .A1(n10622), .A2(n15145), .ZN(n10442) );
  OAI21_X1 U13034 ( .B1(n15145), .B2(n10010), .A(n10442), .ZN(P2_U3502) );
  INV_X1 U13035 ( .A(n13180), .ZN(n10588) );
  OAI222_X1 U13036 ( .A1(n13597), .A2(n10444), .B1(n10588), .B2(P2_U3088), 
        .C1(n10443), .C2(n13599), .ZN(P2_U3313) );
  INV_X1 U13037 ( .A(n10445), .ZN(n10463) );
  OAI222_X1 U13038 ( .A1(n14347), .A2(n10446), .B1(n14327), .B2(n10463), .C1(
        n14744), .C2(P1_U3086), .ZN(P1_U3339) );
  XNOR2_X1 U13039 ( .A(n10657), .B(n12968), .ZN(n10449) );
  NAND2_X1 U13040 ( .A1(n13088), .A2(n10457), .ZN(n10450) );
  XNOR2_X1 U13041 ( .A(n10449), .B(n10450), .ZN(n10484) );
  AND2_X1 U13042 ( .A1(n10484), .A2(n10447), .ZN(n10448) );
  INV_X1 U13043 ( .A(n10449), .ZN(n10458) );
  NAND2_X1 U13044 ( .A1(n10450), .A2(n10458), .ZN(n10451) );
  XNOR2_X1 U13045 ( .A(n15105), .B(n12968), .ZN(n10823) );
  NAND2_X1 U13046 ( .A1(n13087), .A2(n10457), .ZN(n10824) );
  XNOR2_X1 U13047 ( .A(n10823), .B(n10824), .ZN(n10456) );
  NOR2_X1 U13048 ( .A1(n12998), .A2(n10756), .ZN(n10455) );
  AOI22_X1 U13049 ( .A1(n13049), .A2(n13088), .B1(n13086), .B2(n13198), .ZN(
        n10662) );
  OAI22_X1 U13050 ( .A1(n13038), .A2(n10662), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10453), .ZN(n10454) );
  AOI211_X1 U13051 ( .C1(n13007), .C2(n10665), .A(n10455), .B(n10454), .ZN(
        n10462) );
  INV_X1 U13052 ( .A(n10456), .ZN(n10460) );
  NOR2_X1 U13053 ( .A1(n14903), .A2(n11062), .ZN(n13068) );
  INV_X1 U13054 ( .A(n13068), .ZN(n13012) );
  INV_X1 U13055 ( .A(n13088), .ZN(n10658) );
  OAI22_X1 U13056 ( .A1(n13012), .A2(n10658), .B1(n10458), .B2(n14903), .ZN(
        n10459) );
  NAND3_X1 U13057 ( .A1(n10482), .A2(n10460), .A3(n10459), .ZN(n10461) );
  OAI211_X1 U13058 ( .C1(n10827), .C2(n14903), .A(n10462), .B(n10461), .ZN(
        P2_U3199) );
  OAI222_X1 U13059 ( .A1(n13599), .A2(n10464), .B1(n13171), .B2(P2_U3088), 
        .C1(n13597), .C2(n10463), .ZN(P2_U3311) );
  INV_X1 U13060 ( .A(n10465), .ZN(n10498) );
  INV_X1 U13061 ( .A(n15027), .ZN(n10467) );
  OAI222_X1 U13062 ( .A1(n13597), .A2(n10498), .B1(n10467), .B2(P2_U3088), 
        .C1(n10466), .C2(n13599), .ZN(P2_U3310) );
  INV_X1 U13063 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10469) );
  MUX2_X1 U13064 ( .A(n10469), .B(P1_REG2_REG_10__SCAN_IN), .S(n11033), .Z(
        n10470) );
  AOI211_X1 U13065 ( .C1(n10471), .C2(n10470), .A(n14767), .B(n11032), .ZN(
        n10481) );
  INV_X1 U13066 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10472) );
  MUX2_X1 U13067 ( .A(n10472), .B(P1_REG1_REG_10__SCAN_IN), .S(n11033), .Z(
        n10476) );
  OAI21_X1 U13068 ( .B1(n10474), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10473), .ZN(
        n10475) );
  NOR2_X1 U13069 ( .A1(n10475), .A2(n10476), .ZN(n11023) );
  AOI211_X1 U13070 ( .C1(n10476), .C2(n10475), .A(n14772), .B(n11023), .ZN(
        n10480) );
  INV_X1 U13071 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10478) );
  NAND2_X1 U13072 ( .A1(n14778), .A2(n11033), .ZN(n10477) );
  NAND2_X1 U13073 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11783)
         );
  OAI211_X1 U13074 ( .C1(n10478), .C2(n14781), .A(n10477), .B(n11783), .ZN(
        n10479) );
  OR3_X1 U13075 ( .A1(n10481), .A2(n10480), .A3(n10479), .ZN(P1_U3253) );
  OAI21_X1 U13076 ( .B1(n10484), .B2(n10483), .A(n10482), .ZN(n10494) );
  INV_X1 U13077 ( .A(n10484), .ZN(n10486) );
  AND4_X1 U13078 ( .A1(n13068), .A2(n10486), .A3(n9780), .A4(n10485), .ZN(
        n10493) );
  NAND2_X1 U13079 ( .A1(n9780), .A2(n13049), .ZN(n10488) );
  NAND2_X1 U13080 ( .A1(n13087), .A2(n13198), .ZN(n10487) );
  NAND2_X1 U13081 ( .A1(n10488), .A2(n10487), .ZN(n10649) );
  AOI22_X1 U13082 ( .A1(n14914), .A2(n10649), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10490) );
  NAND2_X1 U13083 ( .A1(n14916), .A2(n10657), .ZN(n10489) );
  OAI211_X1 U13084 ( .C1(n14551), .C2(n10491), .A(n10490), .B(n10489), .ZN(
        n10492) );
  AOI211_X1 U13085 ( .C1(n10494), .C2(n14912), .A(n10493), .B(n10492), .ZN(
        n10495) );
  INV_X1 U13086 ( .A(n10495), .ZN(P2_U3202) );
  INV_X1 U13087 ( .A(n10496), .ZN(n10511) );
  OAI222_X1 U13088 ( .A1(n13597), .A2(n10511), .B1(n13181), .B2(P2_U3088), 
        .C1(n10497), .C2(n13599), .ZN(P2_U3312) );
  INV_X1 U13089 ( .A(n13922), .ZN(n14753) );
  OAI222_X1 U13090 ( .A1(n14347), .A2(n7093), .B1(n14327), .B2(n10498), .C1(
        n14753), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U13091 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n13090) );
  NOR2_X1 U13092 ( .A1(n10500), .A2(P2_U3088), .ZN(n14919) );
  INV_X1 U13093 ( .A(n10501), .ZN(n10503) );
  AOI22_X1 U13094 ( .A1(n14914), .A2(n10503), .B1(n14916), .B2(n10502), .ZN(
        n10504) );
  OAI21_X1 U13095 ( .B1(n13090), .B2(n14919), .A(n10504), .ZN(n10508) );
  INV_X1 U13096 ( .A(n10505), .ZN(n10506) );
  AOI211_X1 U13097 ( .C1(n14912), .C2(n10509), .A(n10508), .B(n10507), .ZN(
        n10510) );
  INV_X1 U13098 ( .A(n10510), .ZN(P2_U3194) );
  OAI222_X1 U13099 ( .A1(n14347), .A2(n7095), .B1(n14327), .B2(n10511), .C1(
        n13917), .C2(P1_U3086), .ZN(P1_U3340) );
  XOR2_X1 U13100 ( .A(n10513), .B(n10512), .Z(n10529) );
  AND3_X1 U13101 ( .A1(n10547), .A2(n10515), .A3(n10514), .ZN(n10516) );
  OAI21_X1 U13102 ( .B1(n10517), .B2(n10516), .A(n12547), .ZN(n10525) );
  AND3_X1 U13103 ( .A1(n10553), .A2(n10519), .A3(n10518), .ZN(n10520) );
  OAI21_X1 U13104 ( .B1(n10521), .B2(n10520), .A(n12431), .ZN(n10524) );
  INV_X1 U13105 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10522) );
  NOR2_X1 U13106 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10522), .ZN(n10968) );
  AOI21_X1 U13107 ( .B1(n15168), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n10968), .ZN(
        n10523) );
  NAND3_X1 U13108 ( .A1(n10525), .A2(n10524), .A3(n10523), .ZN(n10526) );
  AOI21_X1 U13109 ( .B1(n10527), .B2(n15175), .A(n10526), .ZN(n10528) );
  OAI21_X1 U13110 ( .B1(n10529), .B2(n15150), .A(n10528), .ZN(P3_U3186) );
  XOR2_X1 U13111 ( .A(n15153), .B(n10530), .Z(n10544) );
  NAND2_X1 U13112 ( .A1(n10531), .A2(n15212), .ZN(n10532) );
  AND2_X1 U13113 ( .A1(n10533), .A2(n10532), .ZN(n10540) );
  NAND2_X1 U13114 ( .A1(n10534), .A2(n10378), .ZN(n10535) );
  NAND2_X1 U13115 ( .A1(n10536), .A2(n10535), .ZN(n10537) );
  NAND2_X1 U13116 ( .A1(n12547), .A2(n10537), .ZN(n10539) );
  AOI22_X1 U13117 ( .A1(n15168), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10538) );
  OAI211_X1 U13118 ( .C1(n10540), .C2(n15162), .A(n10539), .B(n10538), .ZN(
        n10541) );
  AOI21_X1 U13119 ( .B1(n10542), .B2(n15175), .A(n10541), .ZN(n10543) );
  OAI21_X1 U13120 ( .B1(n10544), .B2(n15150), .A(n10543), .ZN(P3_U3183) );
  XOR2_X1 U13121 ( .A(n10546), .B(n10545), .Z(n10560) );
  INV_X1 U13122 ( .A(n10547), .ZN(n10548) );
  AOI21_X1 U13123 ( .B1(n7828), .B2(n10549), .A(n10548), .ZN(n10556) );
  INV_X1 U13124 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10550) );
  NOR2_X1 U13125 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10550), .ZN(n10957) );
  NAND2_X1 U13126 ( .A1(n10551), .A2(n7827), .ZN(n10552) );
  AOI21_X1 U13127 ( .B1(n10553), .B2(n10552), .A(n15162), .ZN(n10554) );
  AOI211_X1 U13128 ( .C1(n15168), .C2(P3_ADDR_REG_3__SCAN_IN), .A(n10957), .B(
        n10554), .ZN(n10555) );
  OAI21_X1 U13129 ( .B1(n10556), .B2(n15164), .A(n10555), .ZN(n10557) );
  AOI21_X1 U13130 ( .B1(n10558), .B2(n15175), .A(n10557), .ZN(n10559) );
  OAI21_X1 U13131 ( .B1(n10560), .B2(n15150), .A(n10559), .ZN(P3_U3185) );
  AND2_X1 U13132 ( .A1(n15081), .A2(n10561), .ZN(n10562) );
  NAND2_X1 U13133 ( .A1(n10621), .A2(n10562), .ZN(n10568) );
  INV_X4 U13134 ( .A(n13446), .ZN(n15076) );
  INV_X1 U13135 ( .A(n10563), .ZN(n10576) );
  INV_X1 U13136 ( .A(n10564), .ZN(n10574) );
  INV_X1 U13137 ( .A(n10565), .ZN(n10566) );
  OR2_X1 U13138 ( .A1(n15076), .A2(n10200), .ZN(n10567) );
  NOR2_X2 U13139 ( .A1(n10568), .A2(n9550), .ZN(n15049) );
  INV_X1 U13140 ( .A(n10569), .ZN(n10570) );
  INV_X1 U13141 ( .A(n15070), .ZN(n15051) );
  AOI22_X1 U13142 ( .A1(n15049), .A2(n10570), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n15051), .ZN(n10572) );
  NAND2_X1 U13143 ( .A1(n15076), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10571) );
  AOI21_X1 U13144 ( .B1(n10574), .B2(n15059), .A(n10573), .ZN(n10575) );
  OAI21_X1 U13145 ( .B1(n15076), .B2(n10576), .A(n10575), .ZN(P2_U3264) );
  INV_X1 U13146 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n10581) );
  AOI21_X1 U13147 ( .B1(n10583), .B2(P2_REG2_REG_13__SCAN_IN), .A(n10577), 
        .ZN(n10578) );
  NOR2_X1 U13148 ( .A1(n10578), .A2(n10588), .ZN(n13167) );
  AOI21_X1 U13149 ( .B1(n10578), .B2(n10588), .A(n13167), .ZN(n10579) );
  INV_X1 U13150 ( .A(n10579), .ZN(n10580) );
  NOR2_X1 U13151 ( .A1(n10580), .A2(n10581), .ZN(n13166) );
  AOI211_X1 U13152 ( .C1(n10581), .C2(n10580), .A(n15008), .B(n13166), .ZN(
        n10591) );
  AOI21_X1 U13153 ( .B1(n10583), .B2(P2_REG1_REG_13__SCAN_IN), .A(n10582), 
        .ZN(n10586) );
  INV_X1 U13154 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10584) );
  MUX2_X1 U13155 ( .A(n10584), .B(P2_REG1_REG_14__SCAN_IN), .S(n13180), .Z(
        n10585) );
  NOR2_X1 U13156 ( .A1(n10586), .A2(n10585), .ZN(n13179) );
  AOI211_X1 U13157 ( .C1(n10586), .C2(n10585), .A(n15022), .B(n13179), .ZN(
        n10590) );
  NAND2_X1 U13158 ( .A1(n14920), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n10587) );
  NAND2_X1 U13159 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14548)
         );
  OAI211_X1 U13160 ( .C1(n15037), .C2(n10588), .A(n10587), .B(n14548), .ZN(
        n10589) );
  OR3_X1 U13161 ( .A1(n10591), .A2(n10590), .A3(n10589), .ZN(P2_U3228) );
  MUX2_X1 U13162 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12539), .Z(n10773) );
  XOR2_X1 U13163 ( .A(n10780), .B(n10773), .Z(n10596) );
  OR2_X1 U13164 ( .A1(n10592), .A2(n7218), .ZN(n10594) );
  NAND2_X1 U13165 ( .A1(n10594), .A2(n10593), .ZN(n10595) );
  NAND2_X1 U13166 ( .A1(n10596), .A2(n10595), .ZN(n10774) );
  OAI21_X1 U13167 ( .B1(n10596), .B2(n10595), .A(n10774), .ZN(n10613) );
  NOR2_X1 U13168 ( .A1(n15147), .A2(n10780), .ZN(n10612) );
  NOR2_X1 U13169 ( .A1(n10598), .A2(n10597), .ZN(n10601) );
  NAND2_X1 U13170 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n10780), .ZN(n10599) );
  OAI21_X1 U13171 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n10780), .A(n10599), .ZN(
        n10600) );
  NOR2_X1 U13172 ( .A1(n10601), .A2(n10600), .ZN(n10782) );
  AOI21_X1 U13173 ( .B1(n10601), .B2(n10600), .A(n10782), .ZN(n10610) );
  NAND2_X1 U13174 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(n10780), .ZN(n10603) );
  OAI21_X1 U13175 ( .B1(P3_REG1_REG_6__SCAN_IN), .B2(n10780), .A(n10603), .ZN(
        n10604) );
  NOR2_X1 U13176 ( .A1(n10605), .A2(n10604), .ZN(n10769) );
  AOI21_X1 U13177 ( .B1(n10605), .B2(n10604), .A(n10769), .ZN(n10606) );
  INV_X1 U13178 ( .A(n10606), .ZN(n10607) );
  NAND2_X1 U13179 ( .A1(n12547), .A2(n10607), .ZN(n10609) );
  AND2_X1 U13180 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n11501) );
  AOI21_X1 U13181 ( .B1(n15168), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n11501), .ZN(
        n10608) );
  OAI211_X1 U13182 ( .C1(n10610), .C2(n15162), .A(n10609), .B(n10608), .ZN(
        n10611) );
  AOI211_X1 U13183 ( .C1(n15173), .C2(n10613), .A(n10612), .B(n10611), .ZN(
        n10614) );
  INV_X1 U13184 ( .A(n10614), .ZN(P3_U3188) );
  NOR3_X1 U13185 ( .A1(n10686), .A2(n15188), .A3(n10615), .ZN(n10616) );
  AOI21_X1 U13186 ( .B1(n15200), .B2(n12374), .A(n10616), .ZN(n11193) );
  MUX2_X1 U13187 ( .A(n7791), .B(n11193), .S(n15254), .Z(n10617) );
  OAI21_X1 U13188 ( .B1(n10694), .B2(n12829), .A(n10617), .ZN(P3_U3459) );
  NOR2_X1 U13189 ( .A1(n10619), .A2(n10618), .ZN(n10620) );
  INV_X1 U13190 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10624) );
  NAND2_X1 U13191 ( .A1(n10622), .A2(n15134), .ZN(n10623) );
  OAI21_X1 U13192 ( .B1(n15134), .B2(n10624), .A(n10623), .ZN(P2_U3439) );
  INV_X1 U13193 ( .A(n10625), .ZN(n10628) );
  NAND2_X1 U13194 ( .A1(n15051), .A2(n9305), .ZN(n10626) );
  OAI211_X1 U13195 ( .C1(n10628), .C2(n9550), .A(n10627), .B(n10626), .ZN(
        n10629) );
  OAI21_X1 U13196 ( .B1(n10630), .B2(n10629), .A(n13446), .ZN(n10633) );
  AOI22_X1 U13197 ( .A1(n14556), .A2(n10631), .B1(P2_REG2_REG_3__SCAN_IN), 
        .B2(n15076), .ZN(n10632) );
  OAI211_X1 U13198 ( .C1(n13448), .C2(n10634), .A(n10633), .B(n10632), .ZN(
        P2_U3262) );
  NAND2_X1 U13199 ( .A1(n10636), .A2(n10635), .ZN(n10640) );
  NAND2_X1 U13200 ( .A1(n10638), .A2(n10637), .ZN(n10639) );
  INV_X1 U13201 ( .A(n10654), .ZN(n10644) );
  XNOR2_X1 U13202 ( .A(n10655), .B(n10644), .ZN(n15096) );
  INV_X1 U13203 ( .A(n15049), .ZN(n13444) );
  NAND2_X1 U13204 ( .A1(n10641), .A2(n15099), .ZN(n10664) );
  OAI211_X1 U13205 ( .C1(n10641), .C2(n15099), .A(n14562), .B(n10664), .ZN(
        n15097) );
  AOI22_X1 U13206 ( .A1(n15076), .A2(P2_REG2_REG_4__SCAN_IN), .B1(n10642), 
        .B2(n15051), .ZN(n10643) );
  OAI21_X1 U13207 ( .B1(n13444), .B2(n15097), .A(n10643), .ZN(n10652) );
  NAND2_X1 U13208 ( .A1(n10647), .A2(n10646), .ZN(n10645) );
  NAND3_X1 U13209 ( .A1(n10647), .A2(n10654), .A3(n10646), .ZN(n10648) );
  AOI21_X1 U13210 ( .B1(n10660), .B2(n10648), .A(n15127), .ZN(n10650) );
  NOR2_X1 U13211 ( .A1(n10650), .A2(n10649), .ZN(n15098) );
  NOR2_X1 U13212 ( .A1(n15098), .A2(n15076), .ZN(n10651) );
  AOI211_X1 U13213 ( .C1(n14556), .C2(n10657), .A(n10652), .B(n10651), .ZN(
        n10653) );
  OAI21_X1 U13214 ( .B1(n13448), .B2(n15096), .A(n10653), .ZN(P2_U3261) );
  NAND2_X1 U13215 ( .A1(n10658), .A2(n15099), .ZN(n10656) );
  XOR2_X1 U13216 ( .A(n10661), .B(n10749), .Z(n15108) );
  NAND2_X1 U13217 ( .A1(n10658), .A2(n10657), .ZN(n10659) );
  XNOR2_X1 U13218 ( .A(n10758), .B(n10661), .ZN(n10663) );
  OAI21_X1 U13219 ( .B1(n10663), .B2(n15127), .A(n10662), .ZN(n15110) );
  NAND2_X1 U13220 ( .A1(n15110), .A2(n13446), .ZN(n10669) );
  AOI211_X1 U13221 ( .C1(n15105), .C2(n10664), .A(n13459), .B(n6803), .ZN(
        n15104) );
  AOI22_X1 U13222 ( .A1(n15076), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n10665), 
        .B2(n15051), .ZN(n10666) );
  OAI21_X1 U13223 ( .B1(n15055), .B2(n10756), .A(n10666), .ZN(n10667) );
  AOI21_X1 U13224 ( .B1(n15104), .B2(n15049), .A(n10667), .ZN(n10668) );
  OAI211_X1 U13225 ( .C1(n15108), .C2(n13448), .A(n10669), .B(n10668), .ZN(
        P2_U3260) );
  INV_X1 U13226 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10670) );
  MUX2_X1 U13227 ( .A(n10670), .B(n11193), .S(n15246), .Z(n10671) );
  OAI21_X1 U13228 ( .B1(n10694), .B2(n12880), .A(n10671), .ZN(P3_U3390) );
  INV_X1 U13229 ( .A(n10681), .ZN(n10677) );
  INV_X1 U13230 ( .A(n10692), .ZN(n10679) );
  NAND3_X1 U13231 ( .A1(n10674), .A2(n10673), .A3(n10672), .ZN(n10675) );
  AOI21_X1 U13232 ( .B1(n10679), .B2(n10682), .A(n10675), .ZN(n10676) );
  OAI21_X1 U13233 ( .B1(n10677), .B2(n10687), .A(n10676), .ZN(n10680) );
  INV_X1 U13234 ( .A(n10678), .ZN(n10691) );
  INV_X1 U13235 ( .A(n12332), .ZN(n12297) );
  NOR2_X1 U13236 ( .A1(n12297), .A2(P3_U3151), .ZN(n10734) );
  NAND3_X1 U13237 ( .A1(n10687), .A2(n10681), .A3(n15195), .ZN(n10684) );
  NAND2_X1 U13238 ( .A1(n10692), .A2(n10682), .ZN(n10683) );
  NAND2_X1 U13239 ( .A1(n10684), .A2(n10683), .ZN(n10685) );
  INV_X1 U13240 ( .A(n10686), .ZN(n10696) );
  INV_X1 U13241 ( .A(n10687), .ZN(n10690) );
  INV_X1 U13242 ( .A(n15190), .ZN(n15208) );
  INV_X1 U13243 ( .A(n11192), .ZN(n10689) );
  INV_X1 U13244 ( .A(n12334), .ZN(n12347) );
  AND2_X1 U13245 ( .A1(n10692), .A2(n10691), .ZN(n10706) );
  INV_X1 U13246 ( .A(n10706), .ZN(n10693) );
  OAI22_X1 U13247 ( .A1(n12347), .A2(n10694), .B1(n7815), .B2(n12328), .ZN(
        n10695) );
  AOI21_X1 U13248 ( .B1(n12340), .B2(n10696), .A(n10695), .ZN(n10697) );
  OAI21_X1 U13249 ( .B1(n10734), .B2(n15146), .A(n10697), .ZN(P3_U3172) );
  NOR2_X1 U13250 ( .A1(n15055), .A2(n9786), .ZN(n10700) );
  INV_X1 U13251 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n14918) );
  OAI22_X1 U13252 ( .A1(n13444), .A2(n10698), .B1(n14918), .B2(n15070), .ZN(
        n10699) );
  AOI211_X1 U13253 ( .C1(n15076), .C2(P2_REG2_REG_2__SCAN_IN), .A(n10700), .B(
        n10699), .ZN(n10703) );
  NAND2_X1 U13254 ( .A1(n15059), .A2(n10701), .ZN(n10702) );
  OAI211_X1 U13255 ( .C1(n15076), .C2(n10704), .A(n10703), .B(n10702), .ZN(
        P2_U3263) );
  INV_X1 U13256 ( .A(n12328), .ZN(n12354) );
  INV_X1 U13257 ( .A(n15202), .ZN(n10707) );
  OAI22_X1 U13258 ( .A1(n12347), .A2(n15196), .B1(n12351), .B2(n10707), .ZN(
        n10708) );
  AOI21_X1 U13259 ( .B1(n12354), .B2(n15201), .A(n10708), .ZN(n10722) );
  NAND2_X1 U13260 ( .A1(n11084), .A2(n12531), .ZN(n10710) );
  NAND2_X1 U13261 ( .A1(n10710), .A2(n10977), .ZN(n10711) );
  NOR3_X1 U13262 ( .A1(n7815), .A2(n15196), .A3(n10712), .ZN(n10714) );
  XNOR2_X1 U13263 ( .A(n10712), .B(n15196), .ZN(n10713) );
  NOR2_X1 U13264 ( .A1(n10713), .A2(n12374), .ZN(n10726) );
  NOR2_X1 U13265 ( .A1(n10714), .A2(n10726), .ZN(n10719) );
  INV_X1 U13266 ( .A(n10718), .ZN(n15197) );
  OAI21_X1 U13267 ( .B1(n15197), .B2(n10712), .A(n10715), .ZN(n10716) );
  NAND2_X1 U13268 ( .A1(n10716), .A2(n10719), .ZN(n10728) );
  NAND3_X1 U13269 ( .A1(n8482), .A2(n15198), .A3(n10712), .ZN(n10717) );
  OAI211_X1 U13270 ( .C1(n10719), .C2(n10718), .A(n10728), .B(n10717), .ZN(
        n10720) );
  NAND2_X1 U13271 ( .A1(n10720), .A2(n12340), .ZN(n10721) );
  OAI211_X1 U13272 ( .C1(n10734), .C2(n10723), .A(n10722), .B(n10721), .ZN(
        P3_U3162) );
  OAI22_X1 U13273 ( .A1(n12347), .A2(n10724), .B1(n12351), .B2(n7815), .ZN(
        n10725) );
  AOI21_X1 U13274 ( .B1(n12354), .B2(n10960), .A(n10725), .ZN(n10732) );
  XNOR2_X1 U13275 ( .A(n10712), .B(n15189), .ZN(n10950) );
  INV_X1 U13276 ( .A(n10726), .ZN(n10727) );
  NAND2_X1 U13277 ( .A1(n10728), .A2(n10727), .ZN(n10729) );
  NAND2_X1 U13278 ( .A1(n10730), .A2(n12340), .ZN(n10731) );
  OAI211_X1 U13279 ( .C1(n10734), .C2(n10733), .A(n10732), .B(n10731), .ZN(
        P3_U3177) );
  OAI21_X1 U13280 ( .B1(n10736), .B2(n10738), .A(n10735), .ZN(n11644) );
  NAND2_X1 U13281 ( .A1(n10737), .A2(n10738), .ZN(n10739) );
  NAND3_X1 U13282 ( .A1(n10740), .A2(n14499), .A3(n10739), .ZN(n10742) );
  AOI22_X1 U13283 ( .A1(n15203), .A2(n15201), .B1(n12373), .B2(n15200), .ZN(
        n10741) );
  NAND2_X1 U13284 ( .A1(n10742), .A2(n10741), .ZN(n11641) );
  AOI21_X1 U13285 ( .B1(n8531), .B2(n11644), .A(n11641), .ZN(n10748) );
  OAI22_X1 U13286 ( .A1(n12829), .A2(n11640), .B1(n15254), .B2(n7828), .ZN(
        n10743) );
  INV_X1 U13287 ( .A(n10743), .ZN(n10744) );
  OAI21_X1 U13288 ( .B1(n10748), .B2(n12766), .A(n10744), .ZN(P3_U3462) );
  INV_X1 U13289 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n10745) );
  OAI22_X1 U13290 ( .A1(n11640), .A2(n12880), .B1(n15246), .B2(n10745), .ZN(
        n10746) );
  INV_X1 U13291 ( .A(n10746), .ZN(n10747) );
  OAI21_X1 U13292 ( .B1(n10748), .B2(n15244), .A(n10747), .ZN(P3_U3399) );
  NAND2_X1 U13293 ( .A1(n13087), .A2(n15105), .ZN(n10750) );
  XOR2_X1 U13294 ( .A(n10994), .B(n10991), .Z(n10984) );
  NAND2_X1 U13295 ( .A1(n13087), .A2(n13049), .ZN(n10753) );
  NAND2_X1 U13296 ( .A1(n13085), .A2(n13198), .ZN(n10752) );
  NAND2_X1 U13297 ( .A1(n10753), .A2(n10752), .ZN(n10979) );
  AOI21_X1 U13298 ( .B1(n10754), .B2(n10997), .A(n13459), .ZN(n10755) );
  AND2_X1 U13299 ( .A1(n11003), .A2(n10755), .ZN(n10987) );
  AOI211_X1 U13300 ( .C1(n15123), .C2(n10997), .A(n10979), .B(n10987), .ZN(
        n10762) );
  NAND2_X1 U13301 ( .A1(n10756), .A2(n13087), .ZN(n10757) );
  INV_X1 U13302 ( .A(n13087), .ZN(n10759) );
  NAND2_X1 U13303 ( .A1(n10759), .A2(n15105), .ZN(n10760) );
  XNOR2_X1 U13304 ( .A(n10995), .B(n10994), .ZN(n10978) );
  NAND2_X1 U13305 ( .A1(n10978), .A2(n14579), .ZN(n10761) );
  OAI211_X1 U13306 ( .C1(n10984), .C2(n14576), .A(n10762), .B(n10761), .ZN(
        n10765) );
  NAND2_X1 U13307 ( .A1(n10765), .A2(n15145), .ZN(n10763) );
  OAI21_X1 U13308 ( .B1(n15145), .B2(n10764), .A(n10763), .ZN(P2_U3505) );
  INV_X1 U13309 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10767) );
  NAND2_X1 U13310 ( .A1(n10765), .A2(n15134), .ZN(n10766) );
  OAI21_X1 U13311 ( .B1(n15134), .B2(n10767), .A(n10766), .ZN(P2_U3448) );
  AND2_X1 U13312 ( .A1(n10780), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10768) );
  NAND2_X1 U13313 ( .A1(n10770), .A2(n11159), .ZN(n11144) );
  AOI21_X1 U13314 ( .B1(n10771), .B2(n7901), .A(n11145), .ZN(n10790) );
  MUX2_X1 U13315 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12539), .Z(n11160) );
  XNOR2_X1 U13316 ( .A(n11160), .B(n10772), .ZN(n10777) );
  OR2_X1 U13317 ( .A1(n10773), .A2(n10780), .ZN(n10775) );
  NAND2_X1 U13318 ( .A1(n10775), .A2(n10774), .ZN(n10776) );
  NAND2_X1 U13319 ( .A1(n10777), .A2(n10776), .ZN(n11161) );
  OAI21_X1 U13320 ( .B1(n10777), .B2(n10776), .A(n11161), .ZN(n10788) );
  INV_X1 U13321 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n10778) );
  NOR2_X1 U13322 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10778), .ZN(n11605) );
  AOI21_X1 U13323 ( .B1(n15168), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11605), .ZN(
        n10779) );
  OAI21_X1 U13324 ( .B1(n15147), .B2(n11159), .A(n10779), .ZN(n10787) );
  AND2_X1 U13325 ( .A1(n10780), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10781) );
  NAND2_X1 U13326 ( .A1(n10783), .A2(n11159), .ZN(n11149) );
  AOI21_X1 U13327 ( .B1(n10784), .B2(n7898), .A(n11150), .ZN(n10785) );
  NOR2_X1 U13328 ( .A1(n10785), .A2(n15162), .ZN(n10786) );
  AOI211_X1 U13329 ( .C1(n15173), .C2(n10788), .A(n10787), .B(n10786), .ZN(
        n10789) );
  OAI21_X1 U13330 ( .B1(n10790), .B2(n15164), .A(n10789), .ZN(P3_U3189) );
  INV_X1 U13331 ( .A(n10792), .ZN(n10933) );
  INV_X1 U13332 ( .A(n10793), .ZN(n10795) );
  NAND2_X1 U13333 ( .A1(n10795), .A2(n10794), .ZN(n10796) );
  NAND2_X1 U13334 ( .A1(n10799), .A2(n10798), .ZN(n10800) );
  XNOR2_X1 U13335 ( .A(n10800), .B(n13604), .ZN(n10803) );
  OAI22_X1 U13336 ( .A1(n13615), .A2(n10801), .B1(n14873), .B2(n13686), .ZN(
        n10802) );
  NAND2_X1 U13337 ( .A1(n10803), .A2(n10802), .ZN(n10805) );
  OAI22_X1 U13338 ( .A1(n13615), .A2(n10929), .B1(n10928), .B2(n13686), .ZN(
        n10806) );
  NAND2_X1 U13339 ( .A1(n10807), .A2(n10806), .ZN(n10891) );
  INV_X1 U13340 ( .A(n10891), .ZN(n10808) );
  NOR2_X1 U13341 ( .A1(n10890), .A2(n10808), .ZN(n10810) );
  AOI22_X1 U13342 ( .A1(n10183), .A2(n14882), .B1(n10220), .B2(n7571), .ZN(
        n10809) );
  XNOR2_X1 U13343 ( .A(n10809), .B(n13604), .ZN(n10892) );
  XNOR2_X1 U13344 ( .A(n10810), .B(n10892), .ZN(n10811) );
  NAND2_X1 U13345 ( .A1(n10811), .A2(n14623), .ZN(n10818) );
  NAND2_X1 U13346 ( .A1(n13894), .A2(n13861), .ZN(n10813) );
  NAND2_X1 U13347 ( .A1(n13893), .A2(n14149), .ZN(n10812) );
  NAND2_X1 U13348 ( .A1(n10813), .A2(n10812), .ZN(n14880) );
  NAND2_X1 U13349 ( .A1(n14625), .A2(n14880), .ZN(n10815) );
  NAND2_X1 U13350 ( .A1(n10815), .A2(n10814), .ZN(n10816) );
  AOI21_X1 U13351 ( .B1(n14621), .B2(n14882), .A(n10816), .ZN(n10817) );
  OAI211_X1 U13352 ( .C1(n14629), .C2(n10933), .A(n10818), .B(n10817), .ZN(
        P1_U3230) );
  XNOR2_X1 U13353 ( .A(n10997), .B(n12968), .ZN(n11103) );
  AND2_X1 U13354 ( .A1(n13086), .A2(n10457), .ZN(n10819) );
  NAND2_X1 U13355 ( .A1(n11103), .A2(n10819), .ZN(n11063) );
  INV_X1 U13356 ( .A(n11103), .ZN(n10821) );
  INV_X1 U13357 ( .A(n10819), .ZN(n10820) );
  NAND2_X1 U13358 ( .A1(n10821), .A2(n10820), .ZN(n10822) );
  NAND2_X1 U13359 ( .A1(n11063), .A2(n10822), .ZN(n10830) );
  INV_X1 U13360 ( .A(n10823), .ZN(n10825) );
  NAND2_X1 U13361 ( .A1(n10825), .A2(n10824), .ZN(n10826) );
  AOI211_X1 U13362 ( .C1(n10830), .C2(n10829), .A(n14903), .B(n6656), .ZN(
        n10835) );
  INV_X1 U13363 ( .A(n10831), .ZN(n10983) );
  AOI22_X1 U13364 ( .A1(n14914), .A2(n10979), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10833) );
  NAND2_X1 U13365 ( .A1(n14916), .A2(n10997), .ZN(n10832) );
  OAI211_X1 U13366 ( .C1(n14551), .C2(n10983), .A(n10833), .B(n10832), .ZN(
        n10834) );
  OR2_X1 U13367 ( .A1(n10835), .A2(n10834), .ZN(P2_U3211) );
  OAI21_X1 U13368 ( .B1(n10838), .B2(n10837), .A(n10836), .ZN(n11631) );
  OAI211_X1 U13369 ( .C1(n10841), .C2(n10840), .A(n10839), .B(n14499), .ZN(
        n10843) );
  AOI22_X1 U13370 ( .A1(n15203), .A2(n10960), .B1(n12372), .B2(n15200), .ZN(
        n10842) );
  NAND2_X1 U13371 ( .A1(n10843), .A2(n10842), .ZN(n11628) );
  AOI21_X1 U13372 ( .B1(n8531), .B2(n11631), .A(n11628), .ZN(n10849) );
  INV_X1 U13373 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n10844) );
  OAI22_X1 U13374 ( .A1(n11627), .A2(n12880), .B1(n15246), .B2(n10844), .ZN(
        n10845) );
  INV_X1 U13375 ( .A(n10845), .ZN(n10846) );
  OAI21_X1 U13376 ( .B1(n10849), .B2(n15244), .A(n10846), .ZN(P3_U3402) );
  OAI22_X1 U13377 ( .A1(n12829), .A2(n11627), .B1(n15254), .B2(n7848), .ZN(
        n10847) );
  INV_X1 U13378 ( .A(n10847), .ZN(n10848) );
  OAI21_X1 U13379 ( .B1(n10849), .B2(n12766), .A(n10848), .ZN(P3_U3463) );
  NAND3_X1 U13380 ( .A1(n10852), .A2(n10851), .A3(n10850), .ZN(n13950) );
  INV_X4 U13381 ( .A(n14165), .ZN(n14842) );
  INV_X1 U13382 ( .A(n10853), .ZN(n10854) );
  XNOR2_X1 U13383 ( .A(n10855), .B(n11961), .ZN(n14869) );
  INV_X1 U13384 ( .A(n14836), .ZN(n10858) );
  INV_X1 U13385 ( .A(n10857), .ZN(n10932) );
  OAI211_X1 U13386 ( .C1(n14873), .C2(n10858), .A(n10932), .B(n14837), .ZN(
        n14870) );
  OAI22_X1 U13387 ( .A1(n14818), .A2(n14870), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14831), .ZN(n10859) );
  AOI21_X1 U13388 ( .B1(n14814), .B2(n13742), .A(n10859), .ZN(n10865) );
  XNOR2_X1 U13389 ( .A(n10860), .B(n11961), .ZN(n10863) );
  OR2_X1 U13390 ( .A1(n13806), .A2(n10929), .ZN(n10862) );
  NAND2_X1 U13391 ( .A1(n13895), .A2(n13861), .ZN(n10861) );
  NAND2_X1 U13392 ( .A1(n10862), .A2(n10861), .ZN(n13741) );
  AOI21_X1 U13393 ( .B1(n10863), .B2(n14269), .A(n13741), .ZN(n14871) );
  MUX2_X1 U13394 ( .A(n10088), .B(n14871), .S(n14165), .Z(n10864) );
  OAI211_X1 U13395 ( .C1(n14161), .C2(n14869), .A(n10865), .B(n10864), .ZN(
        P1_U3290) );
  OAI21_X1 U13396 ( .B1(n10867), .B2(n12125), .A(n10866), .ZN(n10924) );
  INV_X1 U13397 ( .A(n10924), .ZN(n10881) );
  NAND2_X1 U13398 ( .A1(n10943), .A2(n11982), .ZN(n10868) );
  NAND2_X1 U13399 ( .A1(n10868), .A2(n14837), .ZN(n10869) );
  OR2_X1 U13400 ( .A1(n10869), .A2(n11421), .ZN(n10920) );
  AOI21_X1 U13401 ( .B1(n10870), .B2(n12125), .A(n14885), .ZN(n10872) );
  NAND2_X1 U13402 ( .A1(n10872), .A2(n10871), .ZN(n10922) );
  INV_X1 U13403 ( .A(n14831), .ZN(n14841) );
  NAND2_X1 U13404 ( .A1(n13891), .A2(n13861), .ZN(n10874) );
  NAND2_X1 U13405 ( .A1(n13889), .A2(n14149), .ZN(n10873) );
  NAND2_X1 U13406 ( .A1(n10874), .A2(n10873), .ZN(n11523) );
  AOI21_X1 U13407 ( .B1(n14841), .B2(n10875), .A(n11523), .ZN(n10876) );
  OAI211_X1 U13408 ( .C1(n14818), .C2(n10920), .A(n10922), .B(n10876), .ZN(
        n10879) );
  INV_X1 U13409 ( .A(n11982), .ZN(n10877) );
  OAI22_X1 U13410 ( .A1(n10877), .A2(n14845), .B1(n14165), .B2(n10165), .ZN(
        n10878) );
  AOI21_X1 U13411 ( .B1(n10879), .B2(n14165), .A(n10878), .ZN(n10880) );
  OAI21_X1 U13412 ( .B1(n10881), .B2(n14161), .A(n10880), .ZN(P1_U3285) );
  NOR2_X1 U13413 ( .A1(n14842), .A2(n13930), .ZN(n14104) );
  AOI21_X1 U13414 ( .B1(n14837), .B2(n14104), .A(n14814), .ZN(n10889) );
  OAI22_X1 U13415 ( .A1(n14165), .A2(n10883), .B1(n10882), .B2(n14831), .ZN(
        n10884) );
  AOI21_X1 U13416 ( .B1(n10885), .B2(n14165), .A(n10884), .ZN(n10887) );
  INV_X1 U13417 ( .A(n14161), .ZN(n14789) );
  OAI21_X1 U13418 ( .B1(n14789), .B2(n14146), .A(n12118), .ZN(n10886) );
  OAI211_X1 U13419 ( .C1(n10889), .C2(n10888), .A(n10887), .B(n10886), .ZN(
        P1_U3293) );
  INV_X1 U13420 ( .A(n14815), .ZN(n10903) );
  AOI22_X1 U13421 ( .A1(n10183), .A2(n14813), .B1(n7054), .B2(n13893), .ZN(
        n10893) );
  XOR2_X1 U13422 ( .A(n13604), .B(n10893), .Z(n11043) );
  AOI22_X1 U13423 ( .A1(n13759), .A2(n13893), .B1(n7054), .B2(n14813), .ZN(
        n11040) );
  INV_X1 U13424 ( .A(n11040), .ZN(n11042) );
  XNOR2_X1 U13425 ( .A(n11043), .B(n11042), .ZN(n10894) );
  XNOR2_X1 U13426 ( .A(n11045), .B(n10894), .ZN(n10895) );
  NAND2_X1 U13427 ( .A1(n10895), .A2(n14623), .ZN(n10902) );
  OR2_X1 U13428 ( .A1(n13804), .A2(n10929), .ZN(n10897) );
  NAND2_X1 U13429 ( .A1(n13892), .A2(n14149), .ZN(n10896) );
  NAND2_X1 U13430 ( .A1(n10897), .A2(n10896), .ZN(n10909) );
  NAND2_X1 U13431 ( .A1(n14625), .A2(n10909), .ZN(n10898) );
  OAI21_X1 U13432 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n10899), .A(n10898), .ZN(
        n10900) );
  AOI21_X1 U13433 ( .B1(n14621), .B2(n14813), .A(n10900), .ZN(n10901) );
  OAI211_X1 U13434 ( .C1(n14629), .C2(n10903), .A(n10902), .B(n10901), .ZN(
        P1_U3227) );
  INV_X1 U13435 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10915) );
  INV_X1 U13436 ( .A(n10904), .ZN(n10905) );
  AOI21_X1 U13437 ( .B1(n12120), .B2(n10906), .A(n10905), .ZN(n14812) );
  XOR2_X1 U13438 ( .A(n12120), .B(n10907), .Z(n10910) );
  NOR2_X1 U13439 ( .A1(n14812), .A2(n11427), .ZN(n10908) );
  AOI211_X1 U13440 ( .C1(n10910), .C2(n14269), .A(n10909), .B(n10908), .ZN(
        n14823) );
  INV_X1 U13441 ( .A(n10911), .ZN(n11090) );
  OAI211_X1 U13442 ( .C1(n10912), .C2(n10931), .A(n11090), .B(n14837), .ZN(
        n14819) );
  OAI211_X1 U13443 ( .C1(n14812), .C2(n14868), .A(n14823), .B(n14819), .ZN(
        n10916) );
  NAND2_X1 U13444 ( .A1(n10916), .A2(n14891), .ZN(n10914) );
  NAND2_X1 U13445 ( .A1(n14306), .A2(n14813), .ZN(n10913) );
  OAI211_X1 U13446 ( .C1(n14891), .C2(n10915), .A(n10914), .B(n10913), .ZN(
        P1_U3474) );
  INV_X1 U13447 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10919) );
  NAND2_X1 U13448 ( .A1(n10916), .A2(n14896), .ZN(n10918) );
  NAND2_X1 U13449 ( .A1(n14230), .A2(n14813), .ZN(n10917) );
  OAI211_X1 U13450 ( .C1(n14896), .C2(n10919), .A(n10918), .B(n10917), .ZN(
        P1_U3533) );
  INV_X1 U13451 ( .A(n11523), .ZN(n10921) );
  NAND3_X1 U13452 ( .A1(n10922), .A2(n10921), .A3(n10920), .ZN(n10923) );
  AOI21_X1 U13453 ( .B1(n10924), .B2(n14887), .A(n10923), .ZN(n10927) );
  AOI22_X1 U13454 ( .A1(n14306), .A2(n11982), .B1(n14889), .B2(
        P1_REG0_REG_8__SCAN_IN), .ZN(n10925) );
  OAI21_X1 U13455 ( .B1(n10927), .B2(n14889), .A(n10925), .ZN(P1_U3483) );
  AOI22_X1 U13456 ( .A1(n14230), .A2(n11982), .B1(n14894), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n10926) );
  OAI21_X1 U13457 ( .B1(n10927), .B2(n14894), .A(n10926), .ZN(P1_U3536) );
  XNOR2_X1 U13458 ( .A(n10929), .B(n10928), .ZN(n12119) );
  XOR2_X1 U13459 ( .A(n10930), .B(n12119), .Z(n14884) );
  MUX2_X1 U13460 ( .A(n14880), .B(P1_REG2_REG_4__SCAN_IN), .S(n14842), .Z(
        n10937) );
  AOI211_X1 U13461 ( .C1(n14882), .C2(n10932), .A(n10182), .B(n10931), .ZN(
        n14879) );
  INV_X1 U13462 ( .A(n14879), .ZN(n10935) );
  INV_X1 U13463 ( .A(n14104), .ZN(n10934) );
  OAI22_X1 U13464 ( .A1(n10935), .A2(n10934), .B1(n10933), .B2(n14831), .ZN(
        n10936) );
  AOI211_X1 U13465 ( .C1(n14814), .C2(n14882), .A(n10937), .B(n10936), .ZN(
        n10940) );
  XOR2_X1 U13466 ( .A(n12119), .B(n10938), .Z(n14888) );
  NAND2_X1 U13467 ( .A1(n14888), .A2(n14789), .ZN(n10939) );
  OAI211_X1 U13468 ( .C1(n14884), .C2(n14143), .A(n10940), .B(n10939), .ZN(
        P1_U3289) );
  OAI21_X1 U13469 ( .B1(n10942), .B2(n12124), .A(n10941), .ZN(n11016) );
  AOI21_X1 U13470 ( .B1(n11089), .B2(n11979), .A(n10182), .ZN(n10944) );
  AND2_X1 U13471 ( .A1(n10944), .A2(n10943), .ZN(n11015) );
  XNOR2_X1 U13472 ( .A(n10945), .B(n12124), .ZN(n10946) );
  AOI22_X1 U13473 ( .A1(n14149), .A2(n13890), .B1(n13892), .B2(n13861), .ZN(
        n11120) );
  OAI21_X1 U13474 ( .B1(n10946), .B2(n14885), .A(n11120), .ZN(n11011) );
  AOI211_X1 U13475 ( .C1(n14887), .C2(n11016), .A(n11015), .B(n11011), .ZN(
        n10949) );
  AOI22_X1 U13476 ( .A1(n14306), .A2(n11979), .B1(n14889), .B2(
        P1_REG0_REG_7__SCAN_IN), .ZN(n10947) );
  OAI21_X1 U13477 ( .B1(n10949), .B2(n14889), .A(n10947), .ZN(P1_U3480) );
  AOI22_X1 U13478 ( .A1(n14230), .A2(n11979), .B1(n14894), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n10948) );
  OAI21_X1 U13479 ( .B1(n10949), .B2(n14894), .A(n10948), .ZN(P1_U3535) );
  INV_X1 U13480 ( .A(n15201), .ZN(n10955) );
  NAND2_X1 U13481 ( .A1(n10950), .A2(n10955), .ZN(n10951) );
  AND2_X1 U13482 ( .A1(n10952), .A2(n10951), .ZN(n10954) );
  XNOR2_X1 U13483 ( .A(n10712), .B(n6968), .ZN(n10962) );
  XNOR2_X1 U13484 ( .A(n10962), .B(n10960), .ZN(n10953) );
  OAI211_X1 U13485 ( .C1(n10954), .C2(n10953), .A(n12340), .B(n10961), .ZN(
        n10959) );
  INV_X1 U13486 ( .A(n12373), .ZN(n11212) );
  OAI22_X1 U13487 ( .A1(n12351), .A2(n10955), .B1(n11212), .B2(n12328), .ZN(
        n10956) );
  AOI211_X1 U13488 ( .C1(n12358), .C2(n6968), .A(n10957), .B(n10956), .ZN(
        n10958) );
  OAI211_X1 U13489 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12356), .A(n10959), .B(
        n10958), .ZN(P3_U3158) );
  XNOR2_X1 U13490 ( .A(n10712), .B(n10969), .ZN(n10964) );
  NAND2_X1 U13491 ( .A1(n10964), .A2(n11212), .ZN(n11207) );
  OAI21_X1 U13492 ( .B1(n10964), .B2(n11212), .A(n11207), .ZN(n10965) );
  AOI21_X1 U13493 ( .B1(n10966), .B2(n10965), .A(n11209), .ZN(n10973) );
  OAI22_X1 U13494 ( .A1(n12351), .A2(n6969), .B1(n6690), .B2(n12328), .ZN(
        n10967) );
  AOI211_X1 U13495 ( .C1(n12358), .C2(n10969), .A(n10968), .B(n10967), .ZN(
        n10972) );
  INV_X1 U13496 ( .A(n11626), .ZN(n10970) );
  NAND2_X1 U13497 ( .A1(n12297), .A2(n10970), .ZN(n10971) );
  OAI211_X1 U13498 ( .C1(n10973), .C2(n12360), .A(n10972), .B(n10971), .ZN(
        P3_U3170) );
  INV_X1 U13499 ( .A(n10974), .ZN(n10976) );
  OAI222_X1 U13500 ( .A1(P3_U3151), .A2(n10977), .B1(n12903), .B2(n10976), 
        .C1(n10975), .C2(n12900), .ZN(P3_U3275) );
  INV_X1 U13501 ( .A(n10978), .ZN(n10989) );
  NAND2_X1 U13502 ( .A1(n13446), .A2(n14579), .ZN(n13310) );
  NAND2_X1 U13503 ( .A1(n14556), .A2(n10997), .ZN(n10982) );
  INV_X1 U13504 ( .A(n10979), .ZN(n10980) );
  MUX2_X1 U13505 ( .A(n10980), .B(n9983), .S(n15076), .Z(n10981) );
  OAI211_X1 U13506 ( .C1(n15070), .C2(n10983), .A(n10982), .B(n10981), .ZN(
        n10986) );
  NOR2_X1 U13507 ( .A1(n10984), .A2(n13448), .ZN(n10985) );
  AOI211_X1 U13508 ( .C1(n10987), .C2(n15049), .A(n10986), .B(n10985), .ZN(
        n10988) );
  OAI21_X1 U13509 ( .B1(n10989), .B2(n13310), .A(n10988), .ZN(P2_U3259) );
  INV_X1 U13510 ( .A(n10990), .ZN(n11020) );
  INV_X1 U13511 ( .A(n14777), .ZN(n13923) );
  OAI222_X1 U13512 ( .A1(n14347), .A2(n7090), .B1(n14327), .B2(n11020), .C1(
        n13923), .C2(P1_U3086), .ZN(P1_U3337) );
  INV_X1 U13513 ( .A(n10999), .ZN(n10992) );
  OAI21_X1 U13514 ( .B1(n10993), .B2(n10992), .A(n11129), .ZN(n15058) );
  INV_X1 U13515 ( .A(n15058), .ZN(n11005) );
  NAND2_X1 U13516 ( .A1(n10997), .A2(n10996), .ZN(n10998) );
  XNOR2_X1 U13517 ( .A(n11127), .B(n10999), .ZN(n11002) );
  NAND2_X1 U13518 ( .A1(n13086), .A2(n13049), .ZN(n11001) );
  NAND2_X1 U13519 ( .A1(n13084), .A2(n13198), .ZN(n11000) );
  NAND2_X1 U13520 ( .A1(n11001), .A2(n11000), .ZN(n11100) );
  AOI21_X1 U13521 ( .B1(n11002), .B2(n14579), .A(n11100), .ZN(n15061) );
  AOI211_X1 U13522 ( .C1(n15048), .C2(n11003), .A(n13459), .B(n11137), .ZN(
        n15050) );
  AOI21_X1 U13523 ( .B1(n15123), .B2(n15048), .A(n15050), .ZN(n11004) );
  OAI211_X1 U13524 ( .C1(n11005), .C2(n14576), .A(n15061), .B(n11004), .ZN(
        n11008) );
  NAND2_X1 U13525 ( .A1(n11008), .A2(n15145), .ZN(n11006) );
  OAI21_X1 U13526 ( .B1(n15145), .B2(n11007), .A(n11006), .ZN(P2_U3506) );
  INV_X1 U13527 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n11010) );
  NAND2_X1 U13528 ( .A1(n11008), .A2(n15134), .ZN(n11009) );
  OAI21_X1 U13529 ( .B1(n15134), .B2(n11010), .A(n11009), .ZN(P2_U3451) );
  INV_X1 U13530 ( .A(n11011), .ZN(n11019) );
  NOR2_X1 U13531 ( .A1(n14845), .A2(n7227), .ZN(n11014) );
  INV_X1 U13532 ( .A(n11122), .ZN(n11012) );
  OAI22_X1 U13533 ( .A1(n14165), .A2(n10133), .B1(n11012), .B2(n14831), .ZN(
        n11013) );
  AOI211_X1 U13534 ( .C1(n11015), .C2(n14849), .A(n11014), .B(n11013), .ZN(
        n11018) );
  NAND2_X1 U13535 ( .A1(n11016), .A2(n14789), .ZN(n11017) );
  OAI211_X1 U13536 ( .C1(n11019), .C2(n14842), .A(n11018), .B(n11017), .ZN(
        P1_U3286) );
  INV_X1 U13537 ( .A(n13175), .ZN(n15038) );
  OAI222_X1 U13538 ( .A1(n13599), .A2(n11021), .B1(n15038), .B2(P2_U3088), 
        .C1(n13597), .C2(n11020), .ZN(P2_U3309) );
  INV_X1 U13539 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11022) );
  AOI22_X1 U13540 ( .A1(n13913), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n11022), 
        .B2(n11030), .ZN(n11026) );
  INV_X1 U13541 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11024) );
  MUX2_X1 U13542 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n11024), .S(n14680), .Z(
        n14678) );
  NAND2_X1 U13543 ( .A1(n14679), .A2(n14678), .ZN(n14677) );
  OAI21_X1 U13544 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n14680), .A(n14677), 
        .ZN(n11025) );
  OAI21_X1 U13545 ( .B1(n11026), .B2(n11025), .A(n13912), .ZN(n11029) );
  NAND2_X1 U13546 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n13783)
         );
  NAND2_X1 U13547 ( .A1(n14673), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n11027) );
  OAI211_X1 U13548 ( .C1(n14752), .C2(n11030), .A(n13783), .B(n11027), .ZN(
        n11028) );
  AOI21_X1 U13549 ( .B1(n11029), .B2(n14749), .A(n11028), .ZN(n11039) );
  INV_X1 U13550 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11031) );
  AOI22_X1 U13551 ( .A1(n13913), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n11031), 
        .B2(n11030), .ZN(n11036) );
  INV_X1 U13552 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11034) );
  MUX2_X1 U13553 ( .A(n11034), .B(P1_REG2_REG_11__SCAN_IN), .S(n14680), .Z(
        n14683) );
  AOI21_X1 U13554 ( .B1(n14680), .B2(P1_REG2_REG_11__SCAN_IN), .A(n14682), 
        .ZN(n11035) );
  NAND2_X1 U13555 ( .A1(n11036), .A2(n11035), .ZN(n13900) );
  OAI21_X1 U13556 ( .B1(n11036), .B2(n11035), .A(n13900), .ZN(n11037) );
  INV_X1 U13557 ( .A(n14767), .ZN(n14757) );
  NAND2_X1 U13558 ( .A1(n11037), .A2(n14757), .ZN(n11038) );
  NAND2_X1 U13559 ( .A1(n11039), .A2(n11038), .ZN(P1_U3255) );
  INV_X1 U13560 ( .A(n11043), .ZN(n11041) );
  NAND2_X1 U13561 ( .A1(n11041), .A2(n11040), .ZN(n11044) );
  NAND2_X1 U13562 ( .A1(n11976), .A2(n10183), .ZN(n11047) );
  NAND2_X1 U13563 ( .A1(n7054), .A2(n13892), .ZN(n11046) );
  NAND2_X1 U13564 ( .A1(n11047), .A2(n11046), .ZN(n11049) );
  XNOR2_X1 U13565 ( .A(n11049), .B(n11048), .ZN(n11051) );
  AOI22_X1 U13566 ( .A1(n11976), .A2(n7054), .B1(n13759), .B2(n13892), .ZN(
        n11050) );
  OR2_X1 U13567 ( .A1(n11051), .A2(n11050), .ZN(n11112) );
  INV_X1 U13568 ( .A(n11112), .ZN(n11052) );
  AND2_X1 U13569 ( .A1(n11051), .A2(n11050), .ZN(n11111) );
  NOR2_X1 U13570 ( .A1(n11052), .A2(n11111), .ZN(n11053) );
  XNOR2_X1 U13571 ( .A(n11113), .B(n11053), .ZN(n11060) );
  INV_X1 U13572 ( .A(n11054), .ZN(n14802) );
  NAND2_X1 U13573 ( .A1(n13893), .A2(n13861), .ZN(n11056) );
  NAND2_X1 U13574 ( .A1(n13891), .A2(n14149), .ZN(n11055) );
  NAND2_X1 U13575 ( .A1(n11056), .A2(n11055), .ZN(n11095) );
  AOI22_X1 U13576 ( .A1(n14625), .A2(n11095), .B1(P1_REG3_REG_6__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11058) );
  NAND2_X1 U13577 ( .A1(n14621), .A2(n11976), .ZN(n11057) );
  OAI211_X1 U13578 ( .C1(n14629), .C2(n14802), .A(n11058), .B(n11057), .ZN(
        n11059) );
  AOI21_X1 U13579 ( .B1(n11060), .B2(n14623), .A(n11059), .ZN(n11061) );
  INV_X1 U13580 ( .A(n11061), .ZN(P1_U3239) );
  XNOR2_X1 U13581 ( .A(n11222), .B(n12968), .ZN(n11179) );
  NAND2_X1 U13582 ( .A1(n13084), .A2(n10457), .ZN(n11172) );
  XNOR2_X1 U13583 ( .A(n11179), .B(n11172), .ZN(n11077) );
  INV_X1 U13584 ( .A(n11077), .ZN(n11071) );
  XNOR2_X1 U13585 ( .A(n15048), .B(n12968), .ZN(n11064) );
  AND2_X1 U13586 ( .A1(n13085), .A2(n10457), .ZN(n11065) );
  NAND2_X1 U13587 ( .A1(n11064), .A2(n11065), .ZN(n11068) );
  INV_X1 U13588 ( .A(n11064), .ZN(n11076) );
  INV_X1 U13589 ( .A(n11065), .ZN(n11066) );
  NAND2_X1 U13590 ( .A1(n11076), .A2(n11066), .ZN(n11067) );
  AND2_X1 U13591 ( .A1(n11068), .A2(n11067), .ZN(n11104) );
  INV_X1 U13592 ( .A(n11070), .ZN(n11105) );
  AND2_X1 U13593 ( .A1(n11077), .A2(n11068), .ZN(n11069) );
  INV_X1 U13594 ( .A(n11175), .ZN(n11182) );
  AOI21_X1 U13595 ( .B1(n11071), .B2(n11105), .A(n11182), .ZN(n11081) );
  NAND2_X1 U13596 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n14943) );
  NAND2_X1 U13597 ( .A1(n13085), .A2(n13049), .ZN(n11073) );
  NAND2_X1 U13598 ( .A1(n13082), .A2(n13198), .ZN(n11072) );
  NAND2_X1 U13599 ( .A1(n11073), .A2(n11072), .ZN(n11134) );
  NAND2_X1 U13600 ( .A1(n14914), .A2(n11134), .ZN(n11074) );
  OAI211_X1 U13601 ( .C1(n14551), .C2(n11075), .A(n14943), .B(n11074), .ZN(
        n11079) );
  NOR4_X1 U13602 ( .A1(n11077), .A2(n11125), .A3(n11076), .A4(n13012), .ZN(
        n11078) );
  AOI211_X1 U13603 ( .C1(n11222), .C2(n14916), .A(n11079), .B(n11078), .ZN(
        n11080) );
  OAI21_X1 U13604 ( .B1(n11081), .B2(n14903), .A(n11080), .ZN(P2_U3193) );
  NAND2_X1 U13605 ( .A1(n12375), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n11082) );
  OAI21_X1 U13606 ( .B1(n12205), .B2(n12375), .A(n11082), .ZN(P3_U3520) );
  INV_X1 U13607 ( .A(n11083), .ZN(n11086) );
  OAI222_X1 U13608 ( .A1(n12903), .A2(n11086), .B1(n12900), .B2(n11085), .C1(
        P3_U3151), .C2(n11084), .ZN(P3_U3274) );
  OAI21_X1 U13609 ( .B1(n11088), .B2(n11091), .A(n11087), .ZN(n14808) );
  AOI211_X1 U13610 ( .C1(n11976), .C2(n11090), .A(n10182), .B(n7228), .ZN(
        n14807) );
  XNOR2_X1 U13611 ( .A(n11092), .B(n11091), .ZN(n11093) );
  NOR2_X1 U13612 ( .A1(n11093), .A2(n14885), .ZN(n11094) );
  AOI211_X1 U13613 ( .C1(n14877), .C2(n14808), .A(n11095), .B(n11094), .ZN(
        n14811) );
  INV_X1 U13614 ( .A(n14811), .ZN(n11096) );
  AOI211_X1 U13615 ( .C1(n14866), .C2(n14808), .A(n14807), .B(n11096), .ZN(
        n11099) );
  AOI22_X1 U13616 ( .A1(n14230), .A2(n11976), .B1(n14894), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n11097) );
  OAI21_X1 U13617 ( .B1(n11099), .B2(n14894), .A(n11097), .ZN(P1_U3534) );
  AOI22_X1 U13618 ( .A1(n14306), .A2(n11976), .B1(n14889), .B2(
        P1_REG0_REG_6__SCAN_IN), .ZN(n11098) );
  OAI21_X1 U13619 ( .B1(n11099), .B2(n14889), .A(n11098), .ZN(P1_U3477) );
  INV_X1 U13620 ( .A(n15052), .ZN(n11102) );
  NAND2_X1 U13621 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n13154) );
  NAND2_X1 U13622 ( .A1(n14914), .A2(n11100), .ZN(n11101) );
  OAI211_X1 U13623 ( .C1(n14551), .C2(n11102), .A(n13154), .B(n11101), .ZN(
        n11109) );
  NAND3_X1 U13624 ( .A1(n13068), .A2(n13086), .A3(n11103), .ZN(n11107) );
  OAI21_X1 U13625 ( .B1(n6656), .B2(n11104), .A(n14912), .ZN(n11106) );
  AOI21_X1 U13626 ( .B1(n11107), .B2(n11106), .A(n11105), .ZN(n11108) );
  AOI211_X1 U13627 ( .C1(n15048), .C2(n14916), .A(n11109), .B(n11108), .ZN(
        n11110) );
  INV_X1 U13628 ( .A(n11110), .ZN(P2_U3185) );
  INV_X1 U13629 ( .A(n14621), .ZN(n13851) );
  NOR2_X1 U13630 ( .A1(n13615), .A2(n11114), .ZN(n11115) );
  AOI21_X1 U13631 ( .B1(n11979), .B2(n7054), .A(n11115), .ZN(n11531) );
  AOI22_X1 U13632 ( .A1(n11979), .A2(n10183), .B1(n7054), .B2(n13891), .ZN(
        n11116) );
  XNOR2_X1 U13633 ( .A(n11116), .B(n13604), .ZN(n11530) );
  XOR2_X1 U13634 ( .A(n11531), .B(n11530), .Z(n11117) );
  OAI211_X1 U13635 ( .C1(n11118), .C2(n11117), .A(n11529), .B(n14623), .ZN(
        n11124) );
  INV_X1 U13636 ( .A(n14629), .ZN(n13848) );
  OAI22_X1 U13637 ( .A1(n13846), .A2(n11120), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11119), .ZN(n11121) );
  AOI21_X1 U13638 ( .B1(n13848), .B2(n11122), .A(n11121), .ZN(n11123) );
  OAI211_X1 U13639 ( .C1(n7227), .C2(n13851), .A(n11124), .B(n11123), .ZN(
        P1_U3213) );
  AND2_X1 U13640 ( .A1(n15048), .A2(n11125), .ZN(n11126) );
  XNOR2_X1 U13641 ( .A(n11224), .B(n11131), .ZN(n11136) );
  OR2_X1 U13642 ( .A1(n15048), .A2(n13085), .ZN(n11128) );
  NAND2_X1 U13643 ( .A1(n11132), .A2(n11131), .ZN(n11133) );
  INV_X1 U13644 ( .A(n10200), .ZN(n15131) );
  AOI21_X1 U13645 ( .B1(n15118), .B2(n15131), .A(n11134), .ZN(n11135) );
  OAI21_X1 U13646 ( .B1(n15127), .B2(n11136), .A(n11135), .ZN(n15116) );
  INV_X1 U13647 ( .A(n15116), .ZN(n11143) );
  INV_X1 U13648 ( .A(n13427), .ZN(n15073) );
  INV_X1 U13649 ( .A(n11222), .ZN(n15115) );
  OAI211_X1 U13650 ( .C1(n11137), .C2(n15115), .A(n11229), .B(n14562), .ZN(
        n15113) );
  AOI22_X1 U13651 ( .A1(n15076), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n11138), 
        .B2(n15051), .ZN(n11140) );
  NAND2_X1 U13652 ( .A1(n14556), .A2(n11222), .ZN(n11139) );
  OAI211_X1 U13653 ( .C1(n15113), .C2(n13444), .A(n11140), .B(n11139), .ZN(
        n11141) );
  AOI21_X1 U13654 ( .B1(n15118), .B2(n15073), .A(n11141), .ZN(n11142) );
  OAI21_X1 U13655 ( .B1(n11143), .B2(n15076), .A(n11142), .ZN(P2_U3257) );
  INV_X1 U13656 ( .A(n11144), .ZN(n11146) );
  NAND2_X1 U13657 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n11406), .ZN(n11147) );
  OAI21_X1 U13658 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n11406), .A(n11147), .ZN(
        n11148) );
  AOI21_X1 U13659 ( .B1(n6675), .B2(n11148), .A(n11384), .ZN(n11171) );
  INV_X1 U13660 ( .A(n11149), .ZN(n11151) );
  NAND2_X1 U13661 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n11406), .ZN(n11152) );
  OAI21_X1 U13662 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n11406), .A(n11152), .ZN(
        n11153) );
  AOI21_X1 U13663 ( .B1(n6661), .B2(n11153), .A(n11390), .ZN(n11154) );
  NOR2_X1 U13664 ( .A1(n11154), .A2(n15162), .ZN(n11169) );
  AND2_X1 U13665 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n11669) );
  AOI21_X1 U13666 ( .B1(n15168), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11669), .ZN(
        n11167) );
  OR2_X1 U13667 ( .A1(n12539), .A2(n11155), .ZN(n11157) );
  NAND2_X1 U13668 ( .A1(n12539), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n11156) );
  NAND2_X1 U13669 ( .A1(n11157), .A2(n11156), .ZN(n11405) );
  INV_X1 U13670 ( .A(n11406), .ZN(n11158) );
  XNOR2_X1 U13671 ( .A(n11405), .B(n11158), .ZN(n11164) );
  OR2_X1 U13672 ( .A1(n11160), .A2(n11159), .ZN(n11162) );
  NAND2_X1 U13673 ( .A1(n11162), .A2(n11161), .ZN(n11163) );
  NAND2_X1 U13674 ( .A1(n11164), .A2(n11163), .ZN(n11407) );
  OAI21_X1 U13675 ( .B1(n11164), .B2(n11163), .A(n11407), .ZN(n11165) );
  NAND2_X1 U13676 ( .A1(n15173), .A2(n11165), .ZN(n11166) );
  OAI211_X1 U13677 ( .C1(n15147), .C2(n11406), .A(n11167), .B(n11166), .ZN(
        n11168) );
  NOR2_X1 U13678 ( .A1(n11169), .A2(n11168), .ZN(n11170) );
  OAI21_X1 U13679 ( .B1(n11171), .B2(n15164), .A(n11170), .ZN(P3_U3190) );
  INV_X1 U13680 ( .A(n11179), .ZN(n11173) );
  NAND2_X1 U13681 ( .A1(n11173), .A2(n11172), .ZN(n11174) );
  NAND2_X1 U13682 ( .A1(n11175), .A2(n11174), .ZN(n11176) );
  XNOR2_X1 U13683 ( .A(n11274), .B(n12968), .ZN(n11347) );
  NAND2_X1 U13684 ( .A1(n13082), .A2(n10457), .ZN(n11348) );
  XNOR2_X1 U13685 ( .A(n11347), .B(n11348), .ZN(n11180) );
  NAND2_X1 U13686 ( .A1(n11176), .A2(n11180), .ZN(n11351) );
  INV_X1 U13687 ( .A(n11231), .ZN(n11178) );
  INV_X1 U13688 ( .A(n13084), .ZN(n11221) );
  OAI22_X1 U13689 ( .A1(n11356), .A2(n14539), .B1(n11221), .B2(n14541), .ZN(
        n11227) );
  AOI22_X1 U13690 ( .A1(n14914), .A2(n11227), .B1(P2_REG3_REG_9__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11177) );
  OAI21_X1 U13691 ( .B1(n11178), .B2(n14551), .A(n11177), .ZN(n11184) );
  AOI22_X1 U13692 ( .A1(n11179), .A2(n14912), .B1(n13068), .B2(n13084), .ZN(
        n11181) );
  NOR3_X1 U13693 ( .A1(n11182), .A2(n11181), .A3(n11180), .ZN(n11183) );
  AOI211_X1 U13694 ( .C1(n11274), .C2(n14916), .A(n11184), .B(n11183), .ZN(
        n11185) );
  OAI21_X1 U13695 ( .B1(n11351), .B2(n14903), .A(n11185), .ZN(P2_U3203) );
  NAND2_X1 U13696 ( .A1(n12882), .A2(n11186), .ZN(n11187) );
  OAI21_X1 U13697 ( .B1(n12882), .B2(n11188), .A(n11187), .ZN(n11189) );
  INV_X1 U13698 ( .A(n11189), .ZN(n11190) );
  NAND2_X1 U13699 ( .A1(n11191), .A2(n11190), .ZN(n11195) );
  INV_X1 U13700 ( .A(n11193), .ZN(n11194) );
  AOI22_X1 U13701 ( .A1(n11194), .A2(n12749), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(n15209), .ZN(n11198) );
  OR2_X1 U13702 ( .A1(n11195), .A2(n15190), .ZN(n11806) );
  NAND2_X1 U13703 ( .A1(n12660), .A2(n11196), .ZN(n11197) );
  OAI211_X1 U13704 ( .C1(n10360), .C2(n12749), .A(n11198), .B(n11197), .ZN(
        P3_U3233) );
  NOR2_X1 U13705 ( .A1(n12900), .A2(SI_22_), .ZN(n11199) );
  AOI21_X1 U13706 ( .B1(n11200), .B2(P3_STATE_REG_SCAN_IN), .A(n11199), .ZN(
        n11201) );
  OAI21_X1 U13707 ( .B1(n11202), .B2(n12903), .A(n11201), .ZN(n11203) );
  INV_X1 U13708 ( .A(n11203), .ZN(P3_U3273) );
  INV_X1 U13709 ( .A(n11204), .ZN(n11206) );
  OAI222_X1 U13710 ( .A1(n13599), .A2(n11205), .B1(n13597), .B2(n11206), .C1(
        P2_U3088), .C2(n9247), .ZN(P2_U3308) );
  OAI222_X1 U13711 ( .A1(n14347), .A2(n7005), .B1(n14327), .B2(n11206), .C1(
        P1_U3086), .C2(n14138), .ZN(P1_U3336) );
  INV_X1 U13712 ( .A(n11207), .ZN(n11208) );
  AOI21_X1 U13713 ( .B1(n6659), .B2(n11211), .A(n11684), .ZN(n11218) );
  INV_X1 U13714 ( .A(n12371), .ZN(n11603) );
  OAI22_X1 U13715 ( .A1(n12351), .A2(n11212), .B1(n11603), .B2(n12328), .ZN(
        n11213) );
  AOI211_X1 U13716 ( .C1(n12334), .C2(n6691), .A(n11214), .B(n11213), .ZN(
        n11217) );
  INV_X1 U13717 ( .A(n11312), .ZN(n11215) );
  NAND2_X1 U13718 ( .A1(n12297), .A2(n11215), .ZN(n11216) );
  OAI211_X1 U13719 ( .C1(n11218), .C2(n12360), .A(n11217), .B(n11216), .ZN(
        P3_U3167) );
  NAND2_X1 U13720 ( .A1(n11222), .A2(n13084), .ZN(n11219) );
  XNOR2_X1 U13721 ( .A(n11253), .B(n11252), .ZN(n11277) );
  NOR2_X1 U13722 ( .A1(n11222), .A2(n11221), .ZN(n11223) );
  AOI21_X1 U13723 ( .B1(n11225), .B2(n11252), .A(n15127), .ZN(n11228) );
  INV_X1 U13724 ( .A(n11252), .ZN(n11226) );
  AOI21_X1 U13725 ( .B1(n11228), .B2(n11258), .A(n11227), .ZN(n11276) );
  INV_X1 U13726 ( .A(n11276), .ZN(n11236) );
  INV_X1 U13727 ( .A(n11274), .ZN(n11234) );
  AOI21_X1 U13728 ( .B1(n11229), .B2(n11274), .A(n13459), .ZN(n11230) );
  AND2_X1 U13729 ( .A1(n11230), .A2(n11260), .ZN(n11273) );
  NAND2_X1 U13730 ( .A1(n11273), .A2(n15049), .ZN(n11233) );
  AOI22_X1 U13731 ( .A1(n15076), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n11231), 
        .B2(n15051), .ZN(n11232) );
  OAI211_X1 U13732 ( .C1(n11234), .C2(n15055), .A(n11233), .B(n11232), .ZN(
        n11235) );
  AOI21_X1 U13733 ( .B1(n11236), .B2(n13446), .A(n11235), .ZN(n11237) );
  OAI21_X1 U13734 ( .B1(n13448), .B2(n11277), .A(n11237), .ZN(P2_U3256) );
  OAI21_X1 U13735 ( .B1(n11240), .B2(n11239), .A(n11238), .ZN(n11651) );
  OAI211_X1 U13736 ( .C1(n11243), .C2(n11242), .A(n11241), .B(n14499), .ZN(
        n11245) );
  AOI22_X1 U13737 ( .A1(n15203), .A2(n12372), .B1(n12370), .B2(n15200), .ZN(
        n11244) );
  NAND2_X1 U13738 ( .A1(n11245), .A2(n11244), .ZN(n11648) );
  AOI21_X1 U13739 ( .B1(n8531), .B2(n11651), .A(n11648), .ZN(n11251) );
  OAI22_X1 U13740 ( .A1(n12829), .A2(n11647), .B1(n15254), .B2(n7882), .ZN(
        n11246) );
  INV_X1 U13741 ( .A(n11246), .ZN(n11247) );
  OAI21_X1 U13742 ( .B1(n11251), .B2(n12766), .A(n11247), .ZN(P3_U3465) );
  INV_X1 U13743 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n11248) );
  OAI22_X1 U13744 ( .A1(n11647), .A2(n12880), .B1(n15246), .B2(n11248), .ZN(
        n11249) );
  INV_X1 U13745 ( .A(n11249), .ZN(n11250) );
  OAI21_X1 U13746 ( .B1(n11251), .B2(n15244), .A(n11250), .ZN(P3_U3408) );
  NAND2_X1 U13747 ( .A1(n11274), .A2(n13082), .ZN(n11254) );
  XNOR2_X1 U13748 ( .A(n11343), .B(n11259), .ZN(n11300) );
  OR2_X1 U13749 ( .A1(n11274), .A2(n11256), .ZN(n11257) );
  XNOR2_X1 U13750 ( .A(n11330), .B(n11259), .ZN(n11297) );
  NAND2_X1 U13751 ( .A1(n11297), .A2(n13384), .ZN(n11272) );
  NAND2_X1 U13752 ( .A1(n11260), .A2(n11465), .ZN(n11261) );
  NAND2_X1 U13753 ( .A1(n11261), .A2(n14562), .ZN(n11262) );
  NOR2_X1 U13754 ( .A1(n11335), .A2(n11262), .ZN(n11296) );
  INV_X1 U13755 ( .A(n11465), .ZN(n11269) );
  NAND2_X1 U13756 ( .A1(n13082), .A2(n13049), .ZN(n11264) );
  NAND2_X1 U13757 ( .A1(n13080), .A2(n13198), .ZN(n11263) );
  NAND2_X1 U13758 ( .A1(n11264), .A2(n11263), .ZN(n11456) );
  INV_X1 U13759 ( .A(n11456), .ZN(n11266) );
  INV_X1 U13760 ( .A(n11265), .ZN(n11458) );
  OAI22_X1 U13761 ( .A1(n15076), .A2(n11266), .B1(n11458), .B2(n15070), .ZN(
        n11267) );
  AOI21_X1 U13762 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n15076), .A(n11267), 
        .ZN(n11268) );
  OAI21_X1 U13763 ( .B1(n11269), .B2(n15055), .A(n11268), .ZN(n11270) );
  AOI21_X1 U13764 ( .B1(n11296), .B2(n15049), .A(n11270), .ZN(n11271) );
  OAI211_X1 U13765 ( .C1(n11300), .C2(n13448), .A(n11272), .B(n11271), .ZN(
        P2_U3255) );
  AOI21_X1 U13766 ( .B1(n15123), .B2(n11274), .A(n11273), .ZN(n11275) );
  OAI211_X1 U13767 ( .C1(n11277), .C2(n14576), .A(n11276), .B(n11275), .ZN(
        n11280) );
  NAND2_X1 U13768 ( .A1(n11280), .A2(n15145), .ZN(n11278) );
  OAI21_X1 U13769 ( .B1(n15145), .B2(n11279), .A(n11278), .ZN(P2_U3508) );
  INV_X1 U13770 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11282) );
  NAND2_X1 U13771 ( .A1(n11280), .A2(n15134), .ZN(n11281) );
  OAI21_X1 U13772 ( .B1(n15134), .B2(n11282), .A(n11281), .ZN(P2_U3457) );
  OAI21_X1 U13773 ( .B1(n11285), .B2(n11284), .A(n11283), .ZN(n11638) );
  OAI211_X1 U13774 ( .C1(n11287), .C2(n11599), .A(n11286), .B(n14499), .ZN(
        n11289) );
  AOI22_X1 U13775 ( .A1(n15203), .A2(n12371), .B1(n12369), .B2(n15200), .ZN(
        n11288) );
  NAND2_X1 U13776 ( .A1(n11289), .A2(n11288), .ZN(n11635) );
  AOI21_X1 U13777 ( .B1(n8531), .B2(n11638), .A(n11635), .ZN(n11295) );
  INV_X1 U13778 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n11290) );
  OAI22_X1 U13779 ( .A1(n11634), .A2(n12880), .B1(n15246), .B2(n11290), .ZN(
        n11291) );
  INV_X1 U13780 ( .A(n11291), .ZN(n11292) );
  OAI21_X1 U13781 ( .B1(n11295), .B2(n15244), .A(n11292), .ZN(P3_U3411) );
  OAI22_X1 U13782 ( .A1(n12829), .A2(n11634), .B1(n15254), .B2(n7901), .ZN(
        n11293) );
  INV_X1 U13783 ( .A(n11293), .ZN(n11294) );
  OAI21_X1 U13784 ( .B1(n11295), .B2(n12766), .A(n11294), .ZN(P3_U3466) );
  AOI211_X1 U13785 ( .C1(n15123), .C2(n11465), .A(n11456), .B(n11296), .ZN(
        n11299) );
  NAND2_X1 U13786 ( .A1(n11297), .A2(n14579), .ZN(n11298) );
  OAI211_X1 U13787 ( .C1(n11300), .C2(n14576), .A(n11299), .B(n11298), .ZN(
        n11306) );
  NAND2_X1 U13788 ( .A1(n11306), .A2(n15145), .ZN(n11301) );
  OAI21_X1 U13789 ( .B1(n15145), .B2(n10022), .A(n11301), .ZN(P2_U3509) );
  NAND2_X1 U13790 ( .A1(n11302), .A2(n12889), .ZN(n11304) );
  OAI211_X1 U13791 ( .C1(n11305), .C2(n12900), .A(n11304), .B(n11303), .ZN(
        P3_U3272) );
  INV_X1 U13792 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11308) );
  NAND2_X1 U13793 ( .A1(n11306), .A2(n15134), .ZN(n11307) );
  OAI21_X1 U13794 ( .B1(n15134), .B2(n11308), .A(n11307), .ZN(P2_U3460) );
  XNOR2_X1 U13795 ( .A(n11309), .B(n11314), .ZN(n15228) );
  NAND2_X1 U13796 ( .A1(n11310), .A2(n15190), .ZN(n15191) );
  INV_X1 U13797 ( .A(n15191), .ZN(n11311) );
  NAND2_X1 U13798 ( .A1(n12749), .A2(n11311), .ZN(n12593) );
  INV_X1 U13799 ( .A(n12593), .ZN(n15210) );
  NAND2_X1 U13800 ( .A1(n6691), .A2(n15188), .ZN(n15225) );
  OAI22_X1 U13801 ( .A1(n11806), .A2(n15225), .B1(n11312), .B2(n12746), .ZN(
        n11324) );
  OR2_X1 U13802 ( .A1(n11313), .A2(n11314), .ZN(n11316) );
  NAND2_X1 U13803 ( .A1(n11313), .A2(n11314), .ZN(n11315) );
  NAND2_X1 U13804 ( .A1(n11316), .A2(n11315), .ZN(n11320) );
  NAND2_X1 U13805 ( .A1(n12373), .A2(n15203), .ZN(n11318) );
  NAND2_X1 U13806 ( .A1(n12371), .A2(n15200), .ZN(n11317) );
  NAND2_X1 U13807 ( .A1(n11318), .A2(n11317), .ZN(n11319) );
  AOI21_X1 U13808 ( .B1(n11320), .B2(n14499), .A(n11319), .ZN(n11322) );
  INV_X1 U13809 ( .A(n12586), .ZN(n15199) );
  NAND2_X1 U13810 ( .A1(n15228), .A2(n15199), .ZN(n11321) );
  NAND2_X1 U13811 ( .A1(n11322), .A2(n11321), .ZN(n15226) );
  MUX2_X1 U13812 ( .A(n15226), .B(P3_REG2_REG_5__SCAN_IN), .S(n15214), .Z(
        n11323) );
  AOI211_X1 U13813 ( .C1(n15228), .C2(n15210), .A(n11324), .B(n11323), .ZN(
        n11325) );
  INV_X1 U13814 ( .A(n11325), .ZN(P3_U3228) );
  INV_X1 U13815 ( .A(n11326), .ZN(n11368) );
  OAI222_X1 U13816 ( .A1(n13597), .A2(n11368), .B1(n11328), .B2(P2_U3088), 
        .C1(n11327), .C2(n13599), .ZN(P2_U3307) );
  NAND2_X1 U13817 ( .A1(n11465), .A2(n11356), .ZN(n11329) );
  OR2_X1 U13818 ( .A1(n11465), .A2(n11356), .ZN(n11331) );
  INV_X1 U13819 ( .A(n11344), .ZN(n11332) );
  INV_X1 U13820 ( .A(n11614), .ZN(n11333) );
  AOI21_X1 U13821 ( .B1(n11344), .B2(n11334), .A(n11333), .ZN(n15128) );
  INV_X1 U13822 ( .A(n11335), .ZN(n11336) );
  INV_X1 U13823 ( .A(n15122), .ZN(n11367) );
  AOI211_X1 U13824 ( .C1(n15122), .C2(n11336), .A(n13459), .B(n11620), .ZN(
        n15120) );
  NAND2_X1 U13825 ( .A1(n13081), .A2(n13049), .ZN(n11338) );
  NAND2_X1 U13826 ( .A1(n13079), .A2(n13198), .ZN(n11337) );
  NAND2_X1 U13827 ( .A1(n11338), .A2(n11337), .ZN(n15121) );
  AOI22_X1 U13828 ( .A1(n13446), .A2(n15121), .B1(n11364), .B2(n15051), .ZN(
        n11340) );
  NAND2_X1 U13829 ( .A1(n15076), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n11339) );
  OAI211_X1 U13830 ( .C1(n11367), .C2(n15055), .A(n11340), .B(n11339), .ZN(
        n11341) );
  AOI21_X1 U13831 ( .B1(n15120), .B2(n15049), .A(n11341), .ZN(n11346) );
  AND2_X1 U13832 ( .A1(n11465), .A2(n13081), .ZN(n11342) );
  XNOR2_X1 U13833 ( .A(n11609), .B(n11344), .ZN(n15130) );
  NAND2_X1 U13834 ( .A1(n15130), .A2(n15059), .ZN(n11345) );
  OAI211_X1 U13835 ( .C1(n15128), .C2(n13310), .A(n11346), .B(n11345), .ZN(
        P2_U3254) );
  INV_X1 U13836 ( .A(n11347), .ZN(n11349) );
  NAND2_X1 U13837 ( .A1(n11349), .A2(n11348), .ZN(n11350) );
  XNOR2_X1 U13838 ( .A(n11465), .B(n12968), .ZN(n11352) );
  AND2_X1 U13839 ( .A1(n13081), .A2(n10457), .ZN(n11353) );
  NAND2_X1 U13840 ( .A1(n11352), .A2(n11353), .ZN(n11358) );
  INV_X1 U13841 ( .A(n11352), .ZN(n11357) );
  INV_X1 U13842 ( .A(n11353), .ZN(n11354) );
  NAND2_X1 U13843 ( .A1(n11357), .A2(n11354), .ZN(n11355) );
  NAND2_X1 U13844 ( .A1(n11358), .A2(n11355), .ZN(n11462) );
  XNOR2_X1 U13845 ( .A(n15122), .B(n12968), .ZN(n11511) );
  NAND2_X1 U13846 ( .A1(n13080), .A2(n10457), .ZN(n11509) );
  AOI21_X1 U13847 ( .B1(n11459), .B2(n6657), .A(n14903), .ZN(n11360) );
  NOR3_X1 U13848 ( .A1(n11357), .A2(n11356), .A3(n13012), .ZN(n11359) );
  OAI21_X1 U13849 ( .B1(n11360), .B2(n11359), .A(n11513), .ZN(n11366) );
  INV_X1 U13850 ( .A(n15121), .ZN(n11362) );
  OAI22_X1 U13851 ( .A1(n13038), .A2(n11362), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11361), .ZN(n11363) );
  AOI21_X1 U13852 ( .B1(n11364), .B2(n13007), .A(n11363), .ZN(n11365) );
  OAI211_X1 U13853 ( .C1(n11367), .C2(n12998), .A(n11366), .B(n11365), .ZN(
        P2_U3208) );
  OAI222_X1 U13854 ( .A1(n14347), .A2(n11369), .B1(n14327), .B2(n11368), .C1(
        n12085), .C2(P1_U3086), .ZN(P1_U3335) );
  OAI21_X1 U13855 ( .B1(n11372), .B2(n11371), .A(n11370), .ZN(n14790) );
  NAND2_X1 U13856 ( .A1(n13887), .A2(n14149), .ZN(n11784) );
  NAND2_X1 U13857 ( .A1(n11373), .A2(n11784), .ZN(n14783) );
  OAI211_X1 U13858 ( .C1(n11375), .C2(n12127), .A(n11374), .B(n14269), .ZN(
        n11376) );
  NAND2_X1 U13859 ( .A1(n13889), .A2(n13861), .ZN(n11785) );
  AND2_X1 U13860 ( .A1(n11376), .A2(n11785), .ZN(n14792) );
  INV_X1 U13861 ( .A(n14792), .ZN(n11377) );
  AOI211_X1 U13862 ( .C1(n14887), .C2(n14790), .A(n14783), .B(n11377), .ZN(
        n11382) );
  AOI22_X1 U13863 ( .A1(n11995), .A2(n14230), .B1(n14894), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n11378) );
  OAI21_X1 U13864 ( .B1(n11382), .B2(n14894), .A(n11378), .ZN(P1_U3538) );
  INV_X1 U13865 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n11379) );
  OAI22_X1 U13866 ( .A1(n14787), .A2(n14297), .B1(n14891), .B2(n11379), .ZN(
        n11380) );
  INV_X1 U13867 ( .A(n11380), .ZN(n11381) );
  OAI21_X1 U13868 ( .B1(n11382), .B2(n14889), .A(n11381), .ZN(P1_U3489) );
  AND2_X1 U13869 ( .A1(n11406), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n11383) );
  INV_X1 U13870 ( .A(n11385), .ZN(n11387) );
  NAND2_X1 U13871 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n11587), .ZN(n11388) );
  OAI21_X1 U13872 ( .B1(P3_REG1_REG_10__SCAN_IN), .B2(n11587), .A(n11388), 
        .ZN(n11389) );
  AOI21_X1 U13873 ( .B1(n6662), .B2(n11389), .A(n11573), .ZN(n11418) );
  INV_X1 U13874 ( .A(n11391), .ZN(n11393) );
  NAND2_X1 U13875 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n11587), .ZN(n11394) );
  OAI21_X1 U13876 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n11587), .A(n11394), 
        .ZN(n11395) );
  AOI21_X1 U13877 ( .B1(n6660), .B2(n11395), .A(n11577), .ZN(n11396) );
  NOR2_X1 U13878 ( .A1(n11396), .A2(n15162), .ZN(n11416) );
  AND2_X1 U13879 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n11744) );
  AOI21_X1 U13880 ( .B1(n15168), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11744), 
        .ZN(n11414) );
  OR2_X1 U13881 ( .A1(n12539), .A2(n11397), .ZN(n11399) );
  NAND2_X1 U13882 ( .A1(n6488), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n11398) );
  NAND2_X1 U13883 ( .A1(n11399), .A2(n11398), .ZN(n11586) );
  XNOR2_X1 U13884 ( .A(n11586), .B(n11400), .ZN(n11411) );
  MUX2_X1 U13885 ( .A(n11402), .B(n11401), .S(n12539), .Z(n11404) );
  NAND2_X1 U13886 ( .A1(n15174), .A2(n11404), .ZN(n11409) );
  XNOR2_X1 U13887 ( .A(n11404), .B(n11403), .ZN(n15171) );
  OR2_X1 U13888 ( .A1(n11406), .A2(n11405), .ZN(n11408) );
  NAND2_X1 U13889 ( .A1(n11408), .A2(n11407), .ZN(n15170) );
  NAND2_X1 U13890 ( .A1(n15171), .A2(n15170), .ZN(n15169) );
  NAND2_X1 U13891 ( .A1(n11409), .A2(n15169), .ZN(n11410) );
  NAND2_X1 U13892 ( .A1(n11411), .A2(n11410), .ZN(n11588) );
  OAI21_X1 U13893 ( .B1(n11411), .B2(n11410), .A(n11588), .ZN(n11412) );
  NAND2_X1 U13894 ( .A1(n15173), .A2(n11412), .ZN(n11413) );
  OAI211_X1 U13895 ( .C1(n15147), .C2(n11587), .A(n11414), .B(n11413), .ZN(
        n11415) );
  NOR2_X1 U13896 ( .A1(n11416), .A2(n11415), .ZN(n11417) );
  OAI21_X1 U13897 ( .B1(n11418), .B2(n15164), .A(n11417), .ZN(P3_U3192) );
  OAI21_X1 U13898 ( .B1(n11420), .B2(n12126), .A(n11419), .ZN(n14799) );
  XNOR2_X1 U13899 ( .A(n11421), .B(n14797), .ZN(n11422) );
  NOR2_X1 U13900 ( .A1(n11422), .A2(n10182), .ZN(n14793) );
  OAI21_X1 U13901 ( .B1(n6670), .B2(n11424), .A(n11423), .ZN(n11430) );
  NAND2_X1 U13902 ( .A1(n13890), .A2(n13861), .ZN(n11426) );
  NAND2_X1 U13903 ( .A1(n13888), .A2(n14149), .ZN(n11425) );
  NAND2_X1 U13904 ( .A1(n11426), .A2(n11425), .ZN(n11548) );
  INV_X1 U13905 ( .A(n14799), .ZN(n11428) );
  NOR2_X1 U13906 ( .A1(n11428), .A2(n11427), .ZN(n11429) );
  AOI211_X1 U13907 ( .C1(n14269), .C2(n11430), .A(n11548), .B(n11429), .ZN(
        n14801) );
  INV_X1 U13908 ( .A(n14801), .ZN(n11431) );
  AOI211_X1 U13909 ( .C1(n14866), .C2(n14799), .A(n14793), .B(n11431), .ZN(
        n11436) );
  AOI22_X1 U13910 ( .A1(n14230), .A2(n11991), .B1(n14894), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n11432) );
  OAI21_X1 U13911 ( .B1(n11436), .B2(n14894), .A(n11432), .ZN(P1_U3537) );
  INV_X1 U13912 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11433) );
  OAI22_X1 U13913 ( .A1(n14297), .A2(n14797), .B1(n14891), .B2(n11433), .ZN(
        n11434) );
  INV_X1 U13914 ( .A(n11434), .ZN(n11435) );
  OAI21_X1 U13915 ( .B1(n11436), .B2(n14889), .A(n11435), .ZN(P1_U3486) );
  INV_X1 U13916 ( .A(n11437), .ZN(n11440) );
  OAI222_X1 U13917 ( .A1(n14347), .A2(n11438), .B1(n14327), .B2(n11440), .C1(
        P1_U3086), .C2(n12100), .ZN(P1_U3334) );
  OAI222_X1 U13918 ( .A1(n13599), .A2(n11441), .B1(n13597), .B2(n11440), .C1(
        P2_U3088), .C2(n11439), .ZN(P2_U3306) );
  OAI211_X1 U13919 ( .C1(n11443), .C2(n12130), .A(n11442), .B(n14269), .ZN(
        n11446) );
  NAND2_X1 U13920 ( .A1(n13887), .A2(n13861), .ZN(n11445) );
  NAND2_X1 U13921 ( .A1(n13885), .A2(n14149), .ZN(n11444) );
  AND2_X1 U13922 ( .A1(n11445), .A2(n11444), .ZN(n13785) );
  NAND2_X1 U13923 ( .A1(n11446), .A2(n13785), .ZN(n11695) );
  INV_X1 U13924 ( .A(n11695), .ZN(n11455) );
  OAI21_X1 U13925 ( .B1(n11449), .B2(n11448), .A(n11447), .ZN(n11697) );
  INV_X1 U13926 ( .A(n13791), .ZN(n11452) );
  AOI211_X1 U13927 ( .C1(n13791), .C2(n11556), .A(n10182), .B(n11472), .ZN(
        n11696) );
  NAND2_X1 U13928 ( .A1(n11696), .A2(n14849), .ZN(n11451) );
  AOI22_X1 U13929 ( .A1(n14842), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n13782), 
        .B2(n14841), .ZN(n11450) );
  OAI211_X1 U13930 ( .C1(n11452), .C2(n14845), .A(n11451), .B(n11450), .ZN(
        n11453) );
  AOI21_X1 U13931 ( .B1(n11697), .B2(n14789), .A(n11453), .ZN(n11454) );
  OAI21_X1 U13932 ( .B1(n11455), .B2(n14842), .A(n11454), .ZN(P1_U3281) );
  AOI22_X1 U13933 ( .A1(n14914), .A2(n11456), .B1(P2_REG3_REG_10__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11457) );
  OAI21_X1 U13934 ( .B1(n11458), .B2(n14551), .A(n11457), .ZN(n11464) );
  INV_X1 U13935 ( .A(n11459), .ZN(n11460) );
  AOI211_X1 U13936 ( .C1(n11462), .C2(n11461), .A(n14903), .B(n11460), .ZN(
        n11463) );
  AOI211_X1 U13937 ( .C1(n11465), .C2(n14916), .A(n11464), .B(n11463), .ZN(
        n11466) );
  INV_X1 U13938 ( .A(n11466), .ZN(P2_U3189) );
  OAI21_X1 U13939 ( .B1(n11469), .B2(n11468), .A(n11467), .ZN(n14643) );
  OAI21_X1 U13940 ( .B1(n11471), .B2(n12132), .A(n11470), .ZN(n14646) );
  NAND2_X1 U13941 ( .A1(n14646), .A2(n14789), .ZN(n11481) );
  OAI211_X1 U13942 ( .C1(n14642), .C2(n11472), .A(n14837), .B(n11853), .ZN(
        n14641) );
  INV_X1 U13943 ( .A(n14641), .ZN(n11479) );
  NAND2_X1 U13944 ( .A1(n13886), .A2(n13861), .ZN(n11474) );
  NAND2_X1 U13945 ( .A1(n13884), .A2(n14149), .ZN(n11473) );
  AND2_X1 U13946 ( .A1(n11474), .A2(n11473), .ZN(n14640) );
  INV_X1 U13947 ( .A(n13830), .ZN(n11475) );
  OAI22_X1 U13948 ( .A1(n14842), .A2(n14640), .B1(n11475), .B2(n14831), .ZN(
        n11476) );
  AOI21_X1 U13949 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n14842), .A(n11476), 
        .ZN(n11477) );
  OAI21_X1 U13950 ( .B1(n14642), .B2(n14845), .A(n11477), .ZN(n11478) );
  AOI21_X1 U13951 ( .B1(n11479), .B2(n14849), .A(n11478), .ZN(n11480) );
  OAI211_X1 U13952 ( .C1(n14643), .C2(n14143), .A(n11481), .B(n11480), .ZN(
        P1_U3280) );
  INV_X1 U13953 ( .A(n11482), .ZN(n11483) );
  AOI21_X1 U13954 ( .B1(n11485), .B2(n11484), .A(n11483), .ZN(n11489) );
  AOI22_X1 U13955 ( .A1(n15200), .A2(n12368), .B1(n12370), .B2(n15203), .ZN(
        n11488) );
  XNOR2_X1 U13956 ( .A(n11486), .B(n11485), .ZN(n15232) );
  NAND2_X1 U13957 ( .A1(n15232), .A2(n15199), .ZN(n11487) );
  OAI211_X1 U13958 ( .C1(n11489), .C2(n15206), .A(n11488), .B(n11487), .ZN(
        n15230) );
  INV_X1 U13959 ( .A(n15230), .ZN(n11494) );
  INV_X1 U13960 ( .A(n11806), .ZN(n14508) );
  NOR2_X1 U13961 ( .A1(n11664), .A2(n15195), .ZN(n15231) );
  AOI22_X1 U13962 ( .A1(n14508), .A2(n15231), .B1(n15209), .B2(n11490), .ZN(
        n11491) );
  OAI21_X1 U13963 ( .B1(n11155), .B2(n12718), .A(n11491), .ZN(n11492) );
  AOI21_X1 U13964 ( .B1(n15232), .B2(n15210), .A(n11492), .ZN(n11493) );
  OAI21_X1 U13965 ( .B1(n11494), .B2(n15194), .A(n11493), .ZN(P3_U3225) );
  XNOR2_X1 U13966 ( .A(n10712), .B(n11647), .ZN(n11681) );
  XNOR2_X1 U13967 ( .A(n11681), .B(n12371), .ZN(n11498) );
  INV_X1 U13968 ( .A(n11684), .ZN(n11496) );
  NAND2_X1 U13969 ( .A1(n11495), .A2(n6690), .ZN(n11680) );
  NAND2_X1 U13970 ( .A1(n11496), .A2(n11680), .ZN(n11497) );
  NOR2_X1 U13971 ( .A1(n11497), .A2(n11498), .ZN(n11601) );
  AOI211_X1 U13972 ( .C1(n11498), .C2(n11497), .A(n12360), .B(n11601), .ZN(
        n11499) );
  INV_X1 U13973 ( .A(n11499), .ZN(n11504) );
  INV_X1 U13974 ( .A(n12370), .ZN(n11667) );
  OAI22_X1 U13975 ( .A1(n12351), .A2(n6690), .B1(n11667), .B2(n12328), .ZN(
        n11500) );
  AOI211_X1 U13976 ( .C1(n12358), .C2(n11502), .A(n11501), .B(n11500), .ZN(
        n11503) );
  OAI211_X1 U13977 ( .C1(n11646), .C2(n12332), .A(n11504), .B(n11503), .ZN(
        P3_U3179) );
  XNOR2_X1 U13978 ( .A(n11722), .B(n12937), .ZN(n11505) );
  NAND2_X1 U13979 ( .A1(n13079), .A2(n10457), .ZN(n11506) );
  NAND2_X1 U13980 ( .A1(n11505), .A2(n11506), .ZN(n11653) );
  INV_X1 U13981 ( .A(n11505), .ZN(n11508) );
  INV_X1 U13982 ( .A(n11506), .ZN(n11507) );
  NAND2_X1 U13983 ( .A1(n11508), .A2(n11507), .ZN(n11655) );
  NAND2_X1 U13984 ( .A1(n11653), .A2(n11655), .ZN(n11514) );
  INV_X1 U13985 ( .A(n11509), .ZN(n11510) );
  NAND2_X1 U13986 ( .A1(n11511), .A2(n11510), .ZN(n11512) );
  XOR2_X1 U13987 ( .A(n11514), .B(n11654), .Z(n11521) );
  INV_X1 U13988 ( .A(n11621), .ZN(n11518) );
  NAND2_X1 U13989 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n14989)
         );
  NAND2_X1 U13990 ( .A1(n13080), .A2(n13049), .ZN(n11516) );
  NAND2_X1 U13991 ( .A1(n13078), .A2(n13198), .ZN(n11515) );
  NAND2_X1 U13992 ( .A1(n11516), .A2(n11515), .ZN(n11616) );
  NAND2_X1 U13993 ( .A1(n14914), .A2(n11616), .ZN(n11517) );
  OAI211_X1 U13994 ( .C1(n14551), .C2(n11518), .A(n14989), .B(n11517), .ZN(
        n11519) );
  AOI21_X1 U13995 ( .B1(n11722), .B2(n14916), .A(n11519), .ZN(n11520) );
  OAI21_X1 U13996 ( .B1(n11521), .B2(n14903), .A(n11520), .ZN(P2_U3196) );
  AOI21_X1 U13997 ( .B1(n14625), .B2(n11523), .A(n11522), .ZN(n11524) );
  OAI21_X1 U13998 ( .B1(n14629), .B2(n11525), .A(n11524), .ZN(n11536) );
  AOI22_X1 U13999 ( .A1(n11982), .A2(n7054), .B1(n13759), .B2(n13890), .ZN(
        n11539) );
  NAND2_X1 U14000 ( .A1(n11982), .A2(n10183), .ZN(n11527) );
  NAND2_X1 U14001 ( .A1(n7054), .A2(n13890), .ZN(n11526) );
  NAND2_X1 U14002 ( .A1(n11527), .A2(n11526), .ZN(n11528) );
  XNOR2_X1 U14003 ( .A(n11528), .B(n13604), .ZN(n11538) );
  XOR2_X1 U14004 ( .A(n11539), .B(n11538), .Z(n11533) );
  AOI21_X1 U14005 ( .B1(n11533), .B2(n11532), .A(n11541), .ZN(n11534) );
  NOR2_X1 U14006 ( .A1(n11534), .A2(n13868), .ZN(n11535) );
  AOI211_X1 U14007 ( .C1(n14621), .C2(n11982), .A(n11536), .B(n11535), .ZN(
        n11537) );
  INV_X1 U14008 ( .A(n11537), .ZN(P1_U3221) );
  INV_X1 U14009 ( .A(n11538), .ZN(n11540) );
  NAND2_X1 U14010 ( .A1(n11991), .A2(n10183), .ZN(n11543) );
  NAND2_X1 U14011 ( .A1(n7054), .A2(n13889), .ZN(n11542) );
  NAND2_X1 U14012 ( .A1(n11543), .A2(n11542), .ZN(n11544) );
  XNOR2_X1 U14013 ( .A(n11544), .B(n13604), .ZN(n11775) );
  NOR2_X1 U14014 ( .A1(n13615), .A2(n11545), .ZN(n11546) );
  AOI21_X1 U14015 ( .B1(n11991), .B2(n7054), .A(n11546), .ZN(n11777) );
  XNOR2_X1 U14016 ( .A(n11775), .B(n11777), .ZN(n11547) );
  OAI211_X1 U14017 ( .C1(n6669), .C2(n11547), .A(n11776), .B(n14623), .ZN(
        n11553) );
  INV_X1 U14018 ( .A(n14794), .ZN(n11550) );
  AOI22_X1 U14019 ( .A1(n14625), .A2(n11548), .B1(P1_REG3_REG_9__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11549) );
  OAI21_X1 U14020 ( .B1(n14629), .B2(n11550), .A(n11549), .ZN(n11551) );
  INV_X1 U14021 ( .A(n11551), .ZN(n11552) );
  OAI211_X1 U14022 ( .C1(n14797), .C2(n13851), .A(n11553), .B(n11552), .ZN(
        P1_U3231) );
  OAI21_X1 U14023 ( .B1(n11555), .B2(n11560), .A(n11554), .ZN(n14637) );
  INV_X1 U14024 ( .A(n11556), .ZN(n11557) );
  AOI211_X1 U14025 ( .C1(n14630), .C2(n11558), .A(n10182), .B(n11557), .ZN(
        n14631) );
  INV_X1 U14026 ( .A(n11559), .ZN(n11561) );
  AOI21_X1 U14027 ( .B1(n11561), .B2(n11560), .A(n14885), .ZN(n11565) );
  NAND2_X1 U14028 ( .A1(n13888), .A2(n13861), .ZN(n11563) );
  NAND2_X1 U14029 ( .A1(n13886), .A2(n14149), .ZN(n11562) );
  NAND2_X1 U14030 ( .A1(n11563), .A2(n11562), .ZN(n14615) );
  AOI21_X1 U14031 ( .B1(n11565), .B2(n11564), .A(n14615), .ZN(n14639) );
  INV_X1 U14032 ( .A(n14639), .ZN(n11566) );
  AOI211_X1 U14033 ( .C1(n14887), .C2(n14637), .A(n14631), .B(n11566), .ZN(
        n11571) );
  AOI22_X1 U14034 ( .A1(n14630), .A2(n14230), .B1(n14894), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n11567) );
  OAI21_X1 U14035 ( .B1(n11571), .B2(n14894), .A(n11567), .ZN(P1_U3539) );
  INV_X1 U14036 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11568) );
  NOR2_X1 U14037 ( .A1(n14891), .A2(n11568), .ZN(n11569) );
  AOI21_X1 U14038 ( .B1(n14630), .B2(n14306), .A(n11569), .ZN(n11570) );
  OAI21_X1 U14039 ( .B1(n11571), .B2(n14889), .A(n11570), .ZN(P1_U3492) );
  AND2_X1 U14040 ( .A1(n11587), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n11572) );
  NAND2_X1 U14041 ( .A1(n11574), .A2(n11762), .ZN(n11748) );
  AOI21_X1 U14042 ( .B1(n11575), .B2(n7967), .A(n11749), .ZN(n11598) );
  AND2_X1 U14043 ( .A1(n11587), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n11576) );
  NAND2_X1 U14044 ( .A1(n11578), .A2(n11762), .ZN(n11752) );
  OAI21_X1 U14045 ( .B1(n11578), .B2(n11762), .A(n11752), .ZN(n11579) );
  AOI21_X1 U14046 ( .B1(n11579), .B2(n11582), .A(n11753), .ZN(n11580) );
  NOR2_X1 U14047 ( .A1(n11580), .A2(n15162), .ZN(n11596) );
  INV_X1 U14048 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11581) );
  NOR2_X1 U14049 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11581), .ZN(n11872) );
  AOI21_X1 U14050 ( .B1(n15168), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11872), 
        .ZN(n11594) );
  OR2_X1 U14051 ( .A1(n12506), .A2(n11582), .ZN(n11584) );
  NAND2_X1 U14052 ( .A1(n12506), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n11583) );
  NAND2_X1 U14053 ( .A1(n11584), .A2(n11583), .ZN(n11761) );
  XNOR2_X1 U14054 ( .A(n11761), .B(n11585), .ZN(n11591) );
  OR2_X1 U14055 ( .A1(n11587), .A2(n11586), .ZN(n11589) );
  NAND2_X1 U14056 ( .A1(n11589), .A2(n11588), .ZN(n11590) );
  NAND2_X1 U14057 ( .A1(n11591), .A2(n11590), .ZN(n11763) );
  OAI21_X1 U14058 ( .B1(n11591), .B2(n11590), .A(n11763), .ZN(n11592) );
  NAND2_X1 U14059 ( .A1(n15173), .A2(n11592), .ZN(n11593) );
  OAI211_X1 U14060 ( .C1(n15147), .C2(n11762), .A(n11594), .B(n11593), .ZN(
        n11595) );
  NOR2_X1 U14061 ( .A1(n11596), .A2(n11595), .ZN(n11597) );
  OAI21_X1 U14062 ( .B1(n11598), .B2(n15164), .A(n11597), .ZN(P3_U3193) );
  XNOR2_X1 U14063 ( .A(n11599), .B(n10712), .ZN(n11682) );
  INV_X1 U14064 ( .A(n11681), .ZN(n11600) );
  NOR2_X1 U14065 ( .A1(n11600), .A2(n11603), .ZN(n11674) );
  NOR2_X1 U14066 ( .A1(n11601), .A2(n11674), .ZN(n11663) );
  XOR2_X1 U14067 ( .A(n11682), .B(n11663), .Z(n11602) );
  NAND2_X1 U14068 ( .A1(n11602), .A2(n12340), .ZN(n11608) );
  OAI22_X1 U14069 ( .A1(n12351), .A2(n11603), .B1(n7085), .B2(n12328), .ZN(
        n11604) );
  AOI211_X1 U14070 ( .C1(n12358), .C2(n11606), .A(n11605), .B(n11604), .ZN(
        n11607) );
  OAI211_X1 U14071 ( .C1(n11633), .C2(n12332), .A(n11608), .B(n11607), .ZN(
        P3_U3153) );
  NAND2_X1 U14072 ( .A1(n15122), .A2(n13080), .ZN(n11610) );
  INV_X1 U14073 ( .A(n11718), .ZN(n11611) );
  XNOR2_X1 U14074 ( .A(n11719), .B(n11611), .ZN(n14584) );
  NAND2_X1 U14075 ( .A1(n14584), .A2(n15131), .ZN(n11619) );
  NAND2_X1 U14076 ( .A1(n15122), .A2(n11612), .ZN(n11613) );
  AOI21_X1 U14077 ( .B1(n11615), .B2(n11718), .A(n15127), .ZN(n11617) );
  AOI21_X1 U14078 ( .B1(n11617), .B2(n11724), .A(n11616), .ZN(n11618) );
  INV_X1 U14079 ( .A(n11722), .ZN(n14582) );
  OAI211_X1 U14080 ( .C1(n14582), .C2(n11620), .A(n14562), .B(n11726), .ZN(
        n14581) );
  AOI22_X1 U14081 ( .A1(n15076), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n11621), 
        .B2(n15051), .ZN(n11623) );
  NAND2_X1 U14082 ( .A1(n11722), .A2(n14556), .ZN(n11622) );
  OAI211_X1 U14083 ( .C1(n14581), .C2(n13444), .A(n11623), .B(n11622), .ZN(
        n11624) );
  AOI21_X1 U14084 ( .B1(n14584), .B2(n15073), .A(n11624), .ZN(n11625) );
  OAI21_X1 U14085 ( .B1(n14586), .B2(n15076), .A(n11625), .ZN(P2_U3253) );
  NAND2_X1 U14086 ( .A1(n12586), .A2(n15191), .ZN(n14489) );
  OAI22_X1 U14087 ( .A1(n12761), .A2(n11627), .B1(n11626), .B2(n12746), .ZN(
        n11630) );
  MUX2_X1 U14088 ( .A(n11628), .B(P3_REG2_REG_4__SCAN_IN), .S(n15214), .Z(
        n11629) );
  AOI211_X1 U14089 ( .C1(n14509), .C2(n11631), .A(n11630), .B(n11629), .ZN(
        n11632) );
  INV_X1 U14090 ( .A(n11632), .ZN(P3_U3229) );
  OAI22_X1 U14091 ( .A1(n12761), .A2(n11634), .B1(n11633), .B2(n12746), .ZN(
        n11637) );
  MUX2_X1 U14092 ( .A(n11635), .B(P3_REG2_REG_7__SCAN_IN), .S(n15194), .Z(
        n11636) );
  AOI211_X1 U14093 ( .C1(n14509), .C2(n11638), .A(n11637), .B(n11636), .ZN(
        n11639) );
  INV_X1 U14094 ( .A(n11639), .ZN(P3_U3226) );
  OAI22_X1 U14095 ( .A1(n12761), .A2(n11640), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n12746), .ZN(n11643) );
  MUX2_X1 U14096 ( .A(n11641), .B(P3_REG2_REG_3__SCAN_IN), .S(n15214), .Z(
        n11642) );
  AOI211_X1 U14097 ( .C1(n14509), .C2(n11644), .A(n11643), .B(n11642), .ZN(
        n11645) );
  INV_X1 U14098 ( .A(n11645), .ZN(P3_U3230) );
  OAI22_X1 U14099 ( .A1(n12761), .A2(n11647), .B1(n11646), .B2(n12746), .ZN(
        n11650) );
  MUX2_X1 U14100 ( .A(n11648), .B(P3_REG2_REG_6__SCAN_IN), .S(n15214), .Z(
        n11649) );
  AOI211_X1 U14101 ( .C1(n14509), .C2(n11651), .A(n11650), .B(n11649), .ZN(
        n11652) );
  INV_X1 U14102 ( .A(n11652), .ZN(P3_U3227) );
  XNOR2_X1 U14103 ( .A(n14573), .B(n12968), .ZN(n11830) );
  NAND2_X1 U14104 ( .A1(n13078), .A2(n10457), .ZN(n11828) );
  XNOR2_X1 U14105 ( .A(n11830), .B(n11828), .ZN(n11832) );
  XNOR2_X1 U14106 ( .A(n11833), .B(n11832), .ZN(n11662) );
  INV_X1 U14107 ( .A(n11656), .ZN(n11728) );
  NAND2_X1 U14108 ( .A1(n13077), .A2(n13198), .ZN(n11658) );
  NAND2_X1 U14109 ( .A1(n13079), .A2(n13049), .ZN(n11657) );
  NAND2_X1 U14110 ( .A1(n11658), .A2(n11657), .ZN(n14572) );
  AOI22_X1 U14111 ( .A1(n14914), .A2(n14572), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11659) );
  OAI21_X1 U14112 ( .B1(n11728), .B2(n14551), .A(n11659), .ZN(n11660) );
  AOI21_X1 U14113 ( .B1(n14573), .B2(n14916), .A(n11660), .ZN(n11661) );
  OAI21_X1 U14114 ( .B1(n11662), .B2(n14903), .A(n11661), .ZN(P2_U3206) );
  MUX2_X1 U14115 ( .A(n11663), .B(n11667), .S(n11682), .Z(n11665) );
  XNOR2_X1 U14116 ( .A(n11665), .B(n11673), .ZN(n11666) );
  NAND2_X1 U14117 ( .A1(n11666), .A2(n12340), .ZN(n11671) );
  INV_X1 U14118 ( .A(n12368), .ZN(n11742) );
  OAI22_X1 U14119 ( .A1(n12351), .A2(n11667), .B1(n11742), .B2(n12328), .ZN(
        n11668) );
  AOI211_X1 U14120 ( .C1(n12358), .C2(n7086), .A(n11669), .B(n11668), .ZN(
        n11670) );
  OAI211_X1 U14121 ( .C1(n11672), .C2(n12356), .A(n11671), .B(n11670), .ZN(
        P3_U3161) );
  XNOR2_X1 U14122 ( .A(n10712), .B(n11692), .ZN(n11737) );
  XNOR2_X1 U14123 ( .A(n11737), .B(n12368), .ZN(n11688) );
  NAND2_X1 U14124 ( .A1(n11673), .A2(n12370), .ZN(n11676) );
  AOI21_X1 U14125 ( .B1(n11674), .B2(n11673), .A(n11682), .ZN(n11675) );
  AOI21_X1 U14126 ( .B1(n11682), .B2(n11676), .A(n11675), .ZN(n11679) );
  AND2_X1 U14127 ( .A1(n11677), .A2(n12369), .ZN(n11678) );
  OAI21_X1 U14128 ( .B1(n11688), .B2(n11687), .A(n11739), .ZN(n11689) );
  NAND2_X1 U14129 ( .A1(n11689), .A2(n12340), .ZN(n11694) );
  NOR2_X1 U14130 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11690), .ZN(n15167) );
  INV_X1 U14131 ( .A(n14496), .ZN(n11870) );
  OAI22_X1 U14132 ( .A1(n12351), .A2(n7085), .B1(n11870), .B2(n12328), .ZN(
        n11691) );
  AOI211_X1 U14133 ( .C1(n12334), .C2(n11692), .A(n15167), .B(n11691), .ZN(
        n11693) );
  OAI211_X1 U14134 ( .C1(n11710), .C2(n12356), .A(n11694), .B(n11693), .ZN(
        P3_U3171) );
  AOI211_X1 U14135 ( .C1(n14887), .C2(n11697), .A(n11696), .B(n11695), .ZN(
        n11702) );
  AOI22_X1 U14136 ( .A1(n13791), .A2(n14230), .B1(n14894), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n11698) );
  OAI21_X1 U14137 ( .B1(n11702), .B2(n14894), .A(n11698), .ZN(P1_U3540) );
  INV_X1 U14138 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11699) );
  NOR2_X1 U14139 ( .A1(n14891), .A2(n11699), .ZN(n11700) );
  AOI21_X1 U14140 ( .B1(n13791), .B2(n14306), .A(n11700), .ZN(n11701) );
  OAI21_X1 U14141 ( .B1(n11702), .B2(n14889), .A(n11701), .ZN(P1_U3495) );
  XNOR2_X1 U14142 ( .A(n11703), .B(n11705), .ZN(n15234) );
  OAI211_X1 U14143 ( .C1(n11706), .C2(n11705), .A(n11704), .B(n14499), .ZN(
        n11708) );
  AOI22_X1 U14144 ( .A1(n15200), .A2(n14496), .B1(n12369), .B2(n15203), .ZN(
        n11707) );
  OAI211_X1 U14145 ( .C1(n12586), .C2(n15234), .A(n11708), .B(n11707), .ZN(
        n15235) );
  NAND2_X1 U14146 ( .A1(n15235), .A2(n12718), .ZN(n11714) );
  NOR2_X1 U14147 ( .A1(n11709), .A2(n15195), .ZN(n15236) );
  INV_X1 U14148 ( .A(n15236), .ZN(n11711) );
  OAI22_X1 U14149 ( .A1(n11806), .A2(n11711), .B1(n11710), .B2(n12746), .ZN(
        n11712) );
  AOI21_X1 U14150 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n15214), .A(n11712), .ZN(
        n11713) );
  OAI211_X1 U14151 ( .C1(n15234), .C2(n12593), .A(n11714), .B(n11713), .ZN(
        P3_U3224) );
  INV_X1 U14152 ( .A(n11715), .ZN(n11716) );
  OAI222_X1 U14153 ( .A1(n13599), .A2(n11717), .B1(n13597), .B2(n11716), .C1(
        P2_U3088), .C2(n9248), .ZN(P2_U3305) );
  NAND2_X1 U14154 ( .A1(n11722), .A2(n13079), .ZN(n11720) );
  XNOR2_X1 U14155 ( .A(n11878), .B(n11725), .ZN(n14577) );
  OR2_X1 U14156 ( .A1(n11722), .A2(n11721), .ZN(n11723) );
  XNOR2_X1 U14157 ( .A(n11880), .B(n11725), .ZN(n14580) );
  NAND2_X1 U14158 ( .A1(n14580), .A2(n13384), .ZN(n11736) );
  AOI21_X1 U14159 ( .B1(n11726), .B2(n14573), .A(n13459), .ZN(n11727) );
  NAND2_X1 U14160 ( .A1(n11727), .A2(n14560), .ZN(n14574) );
  INV_X1 U14161 ( .A(n14574), .ZN(n11734) );
  INV_X1 U14162 ( .A(n14573), .ZN(n11732) );
  INV_X1 U14163 ( .A(n14572), .ZN(n11729) );
  OAI22_X1 U14164 ( .A1(n15076), .A2(n11729), .B1(n11728), .B2(n15070), .ZN(
        n11730) );
  AOI21_X1 U14165 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n15076), .A(n11730), 
        .ZN(n11731) );
  OAI21_X1 U14166 ( .B1(n11732), .B2(n15055), .A(n11731), .ZN(n11733) );
  AOI21_X1 U14167 ( .B1(n11734), .B2(n15049), .A(n11733), .ZN(n11735) );
  OAI211_X1 U14168 ( .C1(n13448), .C2(n14577), .A(n11736), .B(n11735), .ZN(
        P2_U3252) );
  NAND2_X1 U14169 ( .A1(n11737), .A2(n11742), .ZN(n11738) );
  AND2_X1 U14170 ( .A1(n11739), .A2(n11738), .ZN(n11741) );
  XNOR2_X1 U14171 ( .A(n10712), .B(n11745), .ZN(n11868) );
  XNOR2_X1 U14172 ( .A(n11868), .B(n14496), .ZN(n11740) );
  OAI211_X1 U14173 ( .C1(n11741), .C2(n11740), .A(n12340), .B(n11867), .ZN(
        n11747) );
  INV_X1 U14174 ( .A(n12367), .ZN(n11897) );
  OAI22_X1 U14175 ( .A1(n12351), .A2(n11742), .B1(n11897), .B2(n12328), .ZN(
        n11743) );
  AOI211_X1 U14176 ( .C1(n12334), .C2(n11745), .A(n11744), .B(n11743), .ZN(
        n11746) );
  OAI211_X1 U14177 ( .C1(n11804), .C2(n12356), .A(n11747), .B(n11746), .ZN(
        P3_U3157) );
  INV_X1 U14178 ( .A(n11748), .ZN(n11750) );
  AOI22_X1 U14179 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n12377), .B1(n12382), 
        .B2(n12376), .ZN(n11751) );
  AOI21_X1 U14180 ( .B1(n6663), .B2(n11751), .A(n12379), .ZN(n11774) );
  AOI22_X1 U14181 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n12377), .B1(n12382), 
        .B2(n11898), .ZN(n11756) );
  INV_X1 U14182 ( .A(n11752), .ZN(n11754) );
  AOI21_X1 U14183 ( .B1(n11756), .B2(n11755), .A(n6653), .ZN(n11771) );
  AND2_X1 U14184 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n11910) );
  AOI21_X1 U14185 ( .B1(n15168), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n11910), 
        .ZN(n11770) );
  OR2_X1 U14186 ( .A1(n12506), .A2(n11898), .ZN(n11758) );
  NAND2_X1 U14187 ( .A1(n12506), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n11757) );
  NAND2_X1 U14188 ( .A1(n11758), .A2(n11757), .ZN(n11759) );
  AND2_X1 U14189 ( .A1(n11759), .A2(n12382), .ZN(n12390) );
  NOR2_X1 U14190 ( .A1(n11759), .A2(n12382), .ZN(n11760) );
  OR2_X1 U14191 ( .A1(n12390), .A2(n11760), .ZN(n11765) );
  OR2_X1 U14192 ( .A1(n11762), .A2(n11761), .ZN(n11764) );
  NAND2_X1 U14193 ( .A1(n11764), .A2(n11763), .ZN(n11766) );
  NAND2_X1 U14194 ( .A1(n11765), .A2(n11766), .ZN(n11768) );
  INV_X1 U14195 ( .A(n12389), .ZN(n11767) );
  NAND3_X1 U14196 ( .A1(n15173), .A2(n11768), .A3(n11767), .ZN(n11769) );
  OAI211_X1 U14197 ( .C1(n11771), .C2(n15162), .A(n11770), .B(n11769), .ZN(
        n11772) );
  AOI21_X1 U14198 ( .B1(n12377), .B2(n15175), .A(n11772), .ZN(n11773) );
  OAI21_X1 U14199 ( .B1(n11774), .B2(n15164), .A(n11773), .ZN(P3_U3194) );
  NOR2_X1 U14200 ( .A1(n13615), .A2(n11778), .ZN(n11779) );
  AOI21_X1 U14201 ( .B1(n11995), .B2(n7054), .A(n11779), .ZN(n13622) );
  AOI22_X1 U14202 ( .A1(n11995), .A2(n10183), .B1(n7054), .B2(n13888), .ZN(
        n11780) );
  XNOR2_X1 U14203 ( .A(n11780), .B(n13604), .ZN(n13621) );
  XOR2_X1 U14204 ( .A(n13622), .B(n13621), .Z(n11781) );
  OAI211_X1 U14205 ( .C1(n11782), .C2(n11781), .A(n14610), .B(n14623), .ZN(
        n11789) );
  INV_X1 U14206 ( .A(n11783), .ZN(n11787) );
  AOI21_X1 U14207 ( .B1(n11785), .B2(n11784), .A(n13846), .ZN(n11786) );
  AOI211_X1 U14208 ( .C1(n13848), .C2(n14784), .A(n11787), .B(n11786), .ZN(
        n11788) );
  OAI211_X1 U14209 ( .C1(n14787), .C2(n13851), .A(n11789), .B(n11788), .ZN(
        P1_U3217) );
  NAND2_X1 U14210 ( .A1(n11793), .A2(n14322), .ZN(n11790) );
  OAI211_X1 U14211 ( .C1(n11791), .C2(n14347), .A(n11790), .B(n12157), .ZN(
        P1_U3332) );
  NAND2_X1 U14212 ( .A1(n11793), .A2(n11792), .ZN(n11795) );
  OAI211_X1 U14213 ( .C1(n11796), .C2(n13599), .A(n11795), .B(n11794), .ZN(
        P2_U3304) );
  OAI21_X1 U14214 ( .B1(n6642), .B2(n11797), .A(n14501), .ZN(n15239) );
  AOI22_X1 U14215 ( .A1(n15203), .A2(n12368), .B1(n12367), .B2(n15200), .ZN(
        n11802) );
  OAI211_X1 U14216 ( .C1(n11800), .C2(n11799), .A(n11798), .B(n14499), .ZN(
        n11801) );
  OAI211_X1 U14217 ( .C1(n15239), .C2(n12586), .A(n11802), .B(n11801), .ZN(
        n15240) );
  NAND2_X1 U14218 ( .A1(n15240), .A2(n12718), .ZN(n11809) );
  NOR2_X1 U14219 ( .A1(n11803), .A2(n15195), .ZN(n15241) );
  INV_X1 U14220 ( .A(n15241), .ZN(n11805) );
  OAI22_X1 U14221 ( .A1(n11806), .A2(n11805), .B1(n11804), .B2(n12746), .ZN(
        n11807) );
  AOI21_X1 U14222 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n15214), .A(n11807), 
        .ZN(n11808) );
  OAI211_X1 U14223 ( .C1(n15239), .C2(n12593), .A(n11809), .B(n11808), .ZN(
        P3_U3223) );
  OAI21_X1 U14224 ( .B1(n11811), .B2(n12134), .A(n11810), .ZN(n14279) );
  OAI21_X1 U14225 ( .B1(n6654), .B2(n8831), .A(n11812), .ZN(n14275) );
  AOI21_X1 U14226 ( .B1(n14622), .B2(n6517), .A(n10182), .ZN(n11813) );
  AND2_X1 U14227 ( .A1(n11813), .A2(n14148), .ZN(n14276) );
  NAND2_X1 U14228 ( .A1(n14276), .A2(n14849), .ZN(n11819) );
  NAND2_X1 U14229 ( .A1(n13883), .A2(n14149), .ZN(n11815) );
  NAND2_X1 U14230 ( .A1(n13884), .A2(n13861), .ZN(n11814) );
  NAND2_X1 U14231 ( .A1(n11815), .A2(n11814), .ZN(n14626) );
  INV_X1 U14232 ( .A(n14626), .ZN(n11816) );
  OAI22_X1 U14233 ( .A1(n14842), .A2(n11816), .B1(n14628), .B2(n14831), .ZN(
        n11817) );
  AOI21_X1 U14234 ( .B1(n14842), .B2(P1_REG2_REG_15__SCAN_IN), .A(n11817), 
        .ZN(n11818) );
  OAI211_X1 U14235 ( .C1(n7233), .C2(n14845), .A(n11819), .B(n11818), .ZN(
        n11820) );
  AOI21_X1 U14236 ( .B1(n14275), .B2(n14789), .A(n11820), .ZN(n11821) );
  OAI21_X1 U14237 ( .B1(n14143), .B2(n14279), .A(n11821), .ZN(P1_U3278) );
  INV_X1 U14238 ( .A(n11822), .ZN(n11823) );
  OAI222_X1 U14239 ( .A1(P3_U3151), .A2(n11825), .B1(n12900), .B2(n11824), 
        .C1(n12903), .C2(n11823), .ZN(P3_U3271) );
  XNOR2_X1 U14240 ( .A(n13538), .B(n12937), .ZN(n11827) );
  NAND2_X1 U14241 ( .A1(n13233), .A2(n10457), .ZN(n11826) );
  NAND2_X1 U14242 ( .A1(n11827), .A2(n11826), .ZN(n12906) );
  OAI21_X1 U14243 ( .B1(n11827), .B2(n11826), .A(n12906), .ZN(n11843) );
  INV_X1 U14244 ( .A(n11828), .ZN(n11829) );
  AND2_X1 U14245 ( .A1(n11830), .A2(n11829), .ZN(n11831) );
  XNOR2_X1 U14246 ( .A(n14559), .B(n12937), .ZN(n11834) );
  NAND2_X1 U14247 ( .A1(n13077), .A2(n10457), .ZN(n11835) );
  NAND2_X1 U14248 ( .A1(n11834), .A2(n11835), .ZN(n13061) );
  INV_X1 U14249 ( .A(n11834), .ZN(n11837) );
  INV_X1 U14250 ( .A(n11835), .ZN(n11836) );
  NAND2_X1 U14251 ( .A1(n11837), .A2(n11836), .ZN(n11838) );
  AND2_X1 U14252 ( .A1(n13061), .A2(n11838), .ZN(n14546) );
  XNOR2_X1 U14253 ( .A(n13546), .B(n12968), .ZN(n11839) );
  AND2_X1 U14254 ( .A1(n13076), .A2(n10457), .ZN(n13065) );
  OAI21_X1 U14255 ( .B1(n11839), .B2(n13065), .A(n13061), .ZN(n11841) );
  INV_X1 U14256 ( .A(n11839), .ZN(n13063) );
  INV_X1 U14257 ( .A(n13065), .ZN(n11840) );
  AOI21_X1 U14258 ( .B1(n11843), .B2(n11842), .A(n12907), .ZN(n11849) );
  NAND2_X1 U14259 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n15014)
         );
  NAND2_X1 U14260 ( .A1(n13236), .A2(n13198), .ZN(n11845) );
  NAND2_X1 U14261 ( .A1(n13076), .A2(n13049), .ZN(n11844) );
  NAND2_X1 U14262 ( .A1(n11845), .A2(n11844), .ZN(n13537) );
  NAND2_X1 U14263 ( .A1(n14914), .A2(n13537), .ZN(n11846) );
  OAI211_X1 U14264 ( .C1(n14551), .C2(n11927), .A(n15014), .B(n11846), .ZN(
        n11847) );
  AOI21_X1 U14265 ( .B1(n13538), .B2(n14916), .A(n11847), .ZN(n11848) );
  OAI21_X1 U14266 ( .B1(n11849), .B2(n14903), .A(n11848), .ZN(P2_U3198) );
  INV_X1 U14267 ( .A(n14597), .ZN(n11866) );
  INV_X1 U14268 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11861) );
  INV_X1 U14269 ( .A(n11850), .ZN(n11851) );
  AOI21_X1 U14270 ( .B1(n12133), .B2(n11852), .A(n11851), .ZN(n14162) );
  AOI21_X1 U14271 ( .B1(n14597), .B2(n11853), .A(n10182), .ZN(n11854) );
  AND2_X1 U14272 ( .A1(n11854), .A2(n6517), .ZN(n14167) );
  OAI211_X1 U14273 ( .C1(n11856), .C2(n12133), .A(n11855), .B(n14269), .ZN(
        n11860) );
  NAND2_X1 U14274 ( .A1(n14151), .A2(n14149), .ZN(n11858) );
  NAND2_X1 U14275 ( .A1(n13885), .A2(n13861), .ZN(n11857) );
  NAND2_X1 U14276 ( .A1(n11858), .A2(n11857), .ZN(n14599) );
  INV_X1 U14277 ( .A(n14599), .ZN(n11859) );
  NAND2_X1 U14278 ( .A1(n11860), .A2(n11859), .ZN(n14166) );
  AOI211_X1 U14279 ( .C1(n14162), .C2(n14887), .A(n14167), .B(n14166), .ZN(
        n11863) );
  MUX2_X1 U14280 ( .A(n11861), .B(n11863), .S(n14896), .Z(n11862) );
  OAI21_X1 U14281 ( .B1(n11866), .B2(n14210), .A(n11862), .ZN(P1_U3542) );
  INV_X1 U14282 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n11864) );
  MUX2_X1 U14283 ( .A(n11864), .B(n11863), .S(n14891), .Z(n11865) );
  OAI21_X1 U14284 ( .B1(n11866), .B2(n14297), .A(n11865), .ZN(P1_U3501) );
  XNOR2_X1 U14285 ( .A(n10712), .B(n11873), .ZN(n11903) );
  XNOR2_X1 U14286 ( .A(n11906), .B(n11897), .ZN(n11869) );
  NAND2_X1 U14287 ( .A1(n11869), .A2(n12340), .ZN(n11875) );
  INV_X1 U14288 ( .A(n14497), .ZN(n14487) );
  OAI22_X1 U14289 ( .A1(n12351), .A2(n11870), .B1(n14487), .B2(n12328), .ZN(
        n11871) );
  AOI211_X1 U14290 ( .C1(n12358), .C2(n11873), .A(n11872), .B(n11871), .ZN(
        n11874) );
  OAI211_X1 U14291 ( .C1(n11876), .C2(n12332), .A(n11875), .B(n11874), .ZN(
        P3_U3176) );
  AND2_X1 U14292 ( .A1(n14573), .A2(n13078), .ZN(n11877) );
  NAND2_X1 U14293 ( .A1(n14559), .A2(n13077), .ZN(n11879) );
  XNOR2_X1 U14294 ( .A(n11918), .B(n11920), .ZN(n13549) );
  AND2_X1 U14295 ( .A1(n14559), .A2(n11881), .ZN(n11882) );
  INV_X1 U14296 ( .A(n11883), .ZN(n11884) );
  OAI21_X1 U14297 ( .B1(n11884), .B2(n11919), .A(n11934), .ZN(n13543) );
  INV_X1 U14298 ( .A(n11924), .ZN(n11885) );
  AOI211_X1 U14299 ( .C1(n13546), .C2(n14561), .A(n13459), .B(n11885), .ZN(
        n13544) );
  NAND2_X1 U14300 ( .A1(n13233), .A2(n13198), .ZN(n11887) );
  NAND2_X1 U14301 ( .A1(n13077), .A2(n13049), .ZN(n11886) );
  NAND2_X1 U14302 ( .A1(n11887), .A2(n11886), .ZN(n13545) );
  AOI21_X1 U14303 ( .B1(n13544), .B2(n9247), .A(n13545), .ZN(n11890) );
  AOI22_X1 U14304 ( .A1(n15076), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n13058), 
        .B2(n15051), .ZN(n11889) );
  NAND2_X1 U14305 ( .A1(n13546), .A2(n14556), .ZN(n11888) );
  OAI211_X1 U14306 ( .C1(n11890), .C2(n15076), .A(n11889), .B(n11888), .ZN(
        n11891) );
  AOI21_X1 U14307 ( .B1(n13543), .B2(n13384), .A(n11891), .ZN(n11892) );
  OAI21_X1 U14308 ( .B1(n13448), .B2(n13549), .A(n11892), .ZN(P2_U3250) );
  XNOR2_X1 U14309 ( .A(n11893), .B(n11895), .ZN(n14522) );
  XNOR2_X1 U14310 ( .A(n11894), .B(n11895), .ZN(n11896) );
  OAI222_X1 U14311 ( .A1(n15182), .A2(n11912), .B1(n15183), .B2(n11897), .C1(
        n11896), .C2(n15206), .ZN(n14524) );
  NAND2_X1 U14312 ( .A1(n14524), .A2(n12718), .ZN(n11901) );
  OAI22_X1 U14313 ( .A1(n12718), .A2(n11898), .B1(n11917), .B2(n12746), .ZN(
        n11899) );
  AOI21_X1 U14314 ( .B1(n12660), .B2(n11914), .A(n11899), .ZN(n11900) );
  OAI211_X1 U14315 ( .C1(n12663), .C2(n14522), .A(n11901), .B(n11900), .ZN(
        P3_U3221) );
  XNOR2_X1 U14316 ( .A(n10712), .B(n14520), .ZN(n11902) );
  NOR2_X1 U14317 ( .A1(n11902), .A2(n14497), .ZN(n12161) );
  AOI21_X1 U14318 ( .B1(n11902), .B2(n14497), .A(n12161), .ZN(n11908) );
  INV_X1 U14319 ( .A(n11903), .ZN(n11904) );
  OAI21_X1 U14320 ( .B1(n11908), .B2(n11907), .A(n12163), .ZN(n11909) );
  NAND2_X1 U14321 ( .A1(n11909), .A2(n12340), .ZN(n11916) );
  AOI21_X1 U14322 ( .B1(n12330), .B2(n12367), .A(n11910), .ZN(n11911) );
  OAI21_X1 U14323 ( .B1(n11912), .B2(n12328), .A(n11911), .ZN(n11913) );
  AOI21_X1 U14324 ( .B1(n12334), .B2(n11914), .A(n11913), .ZN(n11915) );
  OAI211_X1 U14325 ( .C1(n11917), .C2(n12356), .A(n11916), .B(n11915), .ZN(
        P3_U3164) );
  INV_X1 U14326 ( .A(n11922), .ZN(n11935) );
  OAI21_X1 U14327 ( .B1(n11923), .B2(n11922), .A(n13235), .ZN(n13542) );
  NAND2_X1 U14328 ( .A1(n11924), .A2(n13538), .ZN(n11925) );
  NAND2_X1 U14329 ( .A1(n11925), .A2(n14562), .ZN(n11926) );
  NOR2_X1 U14330 ( .A1(n13437), .A2(n11926), .ZN(n13536) );
  INV_X1 U14331 ( .A(n13538), .ZN(n11931) );
  INV_X1 U14332 ( .A(n13537), .ZN(n11928) );
  OAI22_X1 U14333 ( .A1(n15076), .A2(n11928), .B1(n11927), .B2(n15070), .ZN(
        n11929) );
  AOI21_X1 U14334 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n15076), .A(n11929), 
        .ZN(n11930) );
  OAI21_X1 U14335 ( .B1(n11931), .B2(n15055), .A(n11930), .ZN(n11932) );
  AOI21_X1 U14336 ( .B1(n13536), .B2(n15049), .A(n11932), .ZN(n11937) );
  INV_X1 U14337 ( .A(n13076), .ZN(n14540) );
  NAND2_X1 U14338 ( .A1(n13546), .A2(n14540), .ZN(n11933) );
  XNOR2_X1 U14339 ( .A(n13212), .B(n11935), .ZN(n13539) );
  NAND2_X1 U14340 ( .A1(n13539), .A2(n13384), .ZN(n11936) );
  OAI211_X1 U14341 ( .C1(n13542), .C2(n13448), .A(n11937), .B(n11936), .ZN(
        P2_U3249) );
  NAND2_X1 U14342 ( .A1(n14323), .A2(n12087), .ZN(n11940) );
  OR2_X1 U14343 ( .A1(n12088), .A2(n14318), .ZN(n11939) );
  NAND2_X1 U14344 ( .A1(n11940), .A2(n11939), .ZN(n12107) );
  INV_X1 U14345 ( .A(n13935), .ZN(n12105) );
  XNOR2_X1 U14346 ( .A(n12107), .B(n12105), .ZN(n12144) );
  NAND2_X1 U14347 ( .A1(n11941), .A2(n13930), .ZN(n13987) );
  OAI21_X1 U14348 ( .B1(n11943), .B2(n11942), .A(n13987), .ZN(n12102) );
  NAND2_X1 U14349 ( .A1(n11946), .A2(n12100), .ZN(n12093) );
  INV_X1 U14350 ( .A(n12085), .ZN(n12101) );
  NAND2_X1 U14351 ( .A1(n11947), .A2(n12101), .ZN(n11948) );
  MUX2_X1 U14352 ( .A(n13871), .B(n14180), .S(n6476), .Z(n12097) );
  MUX2_X1 U14353 ( .A(n14221), .B(n13877), .S(n12002), .Z(n12056) );
  XNOR2_X1 U14354 ( .A(n11950), .B(n12002), .ZN(n11951) );
  INV_X1 U14355 ( .A(n11953), .ZN(n11955) );
  AOI21_X1 U14356 ( .B1(n11955), .B2(n11954), .A(n14825), .ZN(n11956) );
  MUX2_X1 U14357 ( .A(n11959), .B(n11958), .S(n12002), .Z(n11960) );
  NAND2_X1 U14358 ( .A1(n11962), .A2(n11961), .ZN(n11966) );
  MUX2_X1 U14359 ( .A(n11964), .B(n11963), .S(n12002), .Z(n11965) );
  MUX2_X1 U14360 ( .A(n14882), .B(n7571), .S(n12002), .Z(n11969) );
  NAND2_X1 U14361 ( .A1(n11970), .A2(n11969), .ZN(n11968) );
  MUX2_X1 U14362 ( .A(n7571), .B(n14882), .S(n12002), .Z(n11967) );
  NAND2_X1 U14363 ( .A1(n11968), .A2(n11967), .ZN(n11972) );
  MUX2_X1 U14364 ( .A(n13893), .B(n14813), .S(n12002), .Z(n11974) );
  MUX2_X1 U14365 ( .A(n14813), .B(n13893), .S(n12002), .Z(n11973) );
  INV_X1 U14366 ( .A(n11974), .ZN(n11975) );
  MUX2_X1 U14367 ( .A(n11976), .B(n13892), .S(n12002), .Z(n11978) );
  MUX2_X1 U14368 ( .A(n13892), .B(n11976), .S(n12002), .Z(n11977) );
  MUX2_X1 U14369 ( .A(n13891), .B(n11979), .S(n12002), .Z(n11981) );
  MUX2_X1 U14370 ( .A(n13891), .B(n11979), .S(n6476), .Z(n11980) );
  MUX2_X1 U14371 ( .A(n13890), .B(n11982), .S(n6476), .Z(n11986) );
  NAND2_X1 U14372 ( .A1(n11985), .A2(n11986), .ZN(n11984) );
  MUX2_X1 U14373 ( .A(n13890), .B(n11982), .S(n12002), .Z(n11983) );
  NAND2_X1 U14374 ( .A1(n11984), .A2(n11983), .ZN(n11990) );
  INV_X1 U14375 ( .A(n11985), .ZN(n11988) );
  INV_X1 U14376 ( .A(n11986), .ZN(n11987) );
  NAND2_X1 U14377 ( .A1(n11988), .A2(n11987), .ZN(n11989) );
  NAND2_X1 U14378 ( .A1(n11990), .A2(n11989), .ZN(n11993) );
  MUX2_X1 U14379 ( .A(n13889), .B(n11991), .S(n12002), .Z(n11994) );
  MUX2_X1 U14380 ( .A(n13889), .B(n11991), .S(n6476), .Z(n11992) );
  MUX2_X1 U14381 ( .A(n13888), .B(n11995), .S(n6476), .Z(n11999) );
  MUX2_X1 U14382 ( .A(n13888), .B(n11995), .S(n12002), .Z(n11996) );
  NAND2_X1 U14383 ( .A1(n11997), .A2(n11996), .ZN(n12001) );
  MUX2_X1 U14384 ( .A(n13887), .B(n14630), .S(n12002), .Z(n12004) );
  MUX2_X1 U14385 ( .A(n13887), .B(n14630), .S(n6476), .Z(n12003) );
  MUX2_X1 U14386 ( .A(n13886), .B(n13791), .S(n6476), .Z(n12006) );
  MUX2_X1 U14387 ( .A(n13886), .B(n13791), .S(n12002), .Z(n12005) );
  INV_X1 U14388 ( .A(n12006), .ZN(n12007) );
  AND2_X1 U14389 ( .A1(n12026), .A2(n12008), .ZN(n12017) );
  MUX2_X1 U14390 ( .A(n13885), .B(n13837), .S(n12002), .Z(n12013) );
  NAND2_X1 U14391 ( .A1(n12002), .A2(n13885), .ZN(n12012) );
  NAND2_X1 U14392 ( .A1(n13837), .A2(n6476), .ZN(n12011) );
  NAND3_X1 U14393 ( .A1(n12013), .A2(n12012), .A3(n12011), .ZN(n12009) );
  OAI21_X1 U14394 ( .B1(n12013), .B2(n12011), .A(n12133), .ZN(n12016) );
  OR2_X1 U14395 ( .A1(n12013), .A2(n12012), .ZN(n12014) );
  OAI211_X1 U14396 ( .C1(n12133), .C2(n6476), .A(n12014), .B(n12020), .ZN(
        n12015) );
  AOI21_X1 U14397 ( .B1(n12017), .B2(n12016), .A(n12015), .ZN(n12018) );
  NAND2_X1 U14398 ( .A1(n12020), .A2(n12019), .ZN(n12022) );
  AND2_X1 U14399 ( .A1(n12023), .A2(n12021), .ZN(n12027) );
  INV_X1 U14400 ( .A(n14604), .ZN(n14157) );
  OAI22_X1 U14401 ( .A1(n12115), .A2(n14150), .B1(n14157), .B2(n12023), .ZN(
        n12029) );
  OR2_X1 U14402 ( .A1(n12023), .A2(n13805), .ZN(n12024) );
  OAI211_X1 U14403 ( .C1(n12027), .C2(n12026), .A(n12025), .B(n12024), .ZN(
        n12028) );
  NOR2_X1 U14404 ( .A1(n14264), .A2(n12002), .ZN(n12034) );
  AND2_X1 U14405 ( .A1(n14264), .A2(n12002), .ZN(n12033) );
  MUX2_X1 U14406 ( .A(n12034), .B(n12033), .S(n12032), .Z(n12035) );
  NAND2_X1 U14407 ( .A1(n13882), .A2(n6476), .ZN(n12037) );
  OR2_X1 U14408 ( .A1(n6476), .A2(n13882), .ZN(n12036) );
  MUX2_X1 U14409 ( .A(n12037), .B(n12036), .S(n14257), .Z(n12038) );
  MUX2_X1 U14410 ( .A(n12040), .B(n12039), .S(n12002), .Z(n12041) );
  MUX2_X1 U14411 ( .A(n13880), .B(n14240), .S(n12002), .Z(n12045) );
  MUX2_X1 U14412 ( .A(n13880), .B(n14240), .S(n6476), .Z(n12042) );
  NAND2_X1 U14413 ( .A1(n12043), .A2(n12042), .ZN(n12049) );
  INV_X1 U14414 ( .A(n12044), .ZN(n12047) );
  INV_X1 U14415 ( .A(n12045), .ZN(n12046) );
  MUX2_X1 U14416 ( .A(n13879), .B(n14076), .S(n6476), .Z(n12051) );
  MUX2_X1 U14417 ( .A(n13879), .B(n14076), .S(n12002), .Z(n12050) );
  MUX2_X1 U14418 ( .A(n13878), .B(n14305), .S(n12002), .Z(n12053) );
  MUX2_X1 U14419 ( .A(n13774), .B(n14065), .S(n6476), .Z(n12052) );
  MUX2_X1 U14420 ( .A(n13877), .B(n14221), .S(n12002), .Z(n12055) );
  MUX2_X1 U14421 ( .A(n13876), .B(n14211), .S(n12002), .Z(n12060) );
  NAND2_X1 U14422 ( .A1(n12059), .A2(n12060), .ZN(n12058) );
  MUX2_X1 U14423 ( .A(n13876), .B(n14211), .S(n6476), .Z(n12057) );
  NAND2_X1 U14424 ( .A1(n12058), .A2(n12057), .ZN(n12064) );
  INV_X1 U14425 ( .A(n12059), .ZN(n12062) );
  INV_X1 U14426 ( .A(n12060), .ZN(n12061) );
  MUX2_X1 U14427 ( .A(n13875), .B(n14201), .S(n6476), .Z(n12066) );
  MUX2_X1 U14428 ( .A(n13875), .B(n14201), .S(n12002), .Z(n12065) );
  MUX2_X1 U14429 ( .A(n13874), .B(n13866), .S(n12002), .Z(n12068) );
  MUX2_X1 U14430 ( .A(n13874), .B(n13866), .S(n6476), .Z(n12067) );
  INV_X1 U14431 ( .A(n12068), .ZN(n12069) );
  MUX2_X1 U14432 ( .A(n13873), .B(n13988), .S(n6476), .Z(n12073) );
  NAND2_X1 U14433 ( .A1(n12072), .A2(n12073), .ZN(n12071) );
  MUX2_X1 U14434 ( .A(n13873), .B(n13988), .S(n12002), .Z(n12070) );
  NAND2_X1 U14435 ( .A1(n12071), .A2(n12070), .ZN(n12077) );
  INV_X1 U14436 ( .A(n12072), .ZN(n12075) );
  INV_X1 U14437 ( .A(n12073), .ZN(n12074) );
  NAND2_X1 U14438 ( .A1(n12075), .A2(n12074), .ZN(n12076) );
  MUX2_X1 U14439 ( .A(n13872), .B(n14288), .S(n12002), .Z(n12081) );
  NAND2_X1 U14440 ( .A1(n12080), .A2(n12081), .ZN(n12079) );
  MUX2_X1 U14441 ( .A(n13872), .B(n14288), .S(n6476), .Z(n12078) );
  INV_X1 U14442 ( .A(n12080), .ZN(n12083) );
  INV_X1 U14443 ( .A(n12081), .ZN(n12082) );
  MUX2_X1 U14444 ( .A(n13871), .B(n14180), .S(n12002), .Z(n12084) );
  OAI21_X1 U14445 ( .B1(n13935), .B2(n12085), .A(n13870), .ZN(n12086) );
  INV_X1 U14446 ( .A(n12086), .ZN(n12091) );
  NAND2_X1 U14447 ( .A1(n13573), .A2(n12087), .ZN(n12090) );
  OR2_X1 U14448 ( .A1(n12088), .A2(n14328), .ZN(n12089) );
  MUX2_X1 U14449 ( .A(n12091), .B(n13942), .S(n12002), .Z(n12099) );
  NAND2_X1 U14450 ( .A1(n12002), .A2(n13935), .ZN(n12094) );
  INV_X1 U14451 ( .A(n13870), .ZN(n12092) );
  AOI21_X1 U14452 ( .B1(n12094), .B2(n12093), .A(n12092), .ZN(n12095) );
  AOI21_X1 U14453 ( .B1(n13942), .B2(n6476), .A(n12095), .ZN(n12098) );
  NAND2_X1 U14454 ( .A1(n12099), .A2(n12098), .ZN(n12096) );
  INV_X1 U14455 ( .A(n12149), .ZN(n12152) );
  INV_X1 U14456 ( .A(n12102), .ZN(n12109) );
  INV_X1 U14457 ( .A(n12144), .ZN(n12104) );
  NAND2_X1 U14458 ( .A1(n12101), .A2(n12100), .ZN(n12147) );
  AND2_X1 U14459 ( .A1(n12102), .A2(n12147), .ZN(n12111) );
  INV_X1 U14460 ( .A(n12111), .ZN(n12103) );
  NOR2_X1 U14461 ( .A1(n12104), .A2(n12103), .ZN(n12108) );
  MUX2_X1 U14462 ( .A(n14282), .B(n12105), .S(n12002), .Z(n12106) );
  OAI21_X1 U14463 ( .B1(n12107), .B2(n13935), .A(n12106), .ZN(n12112) );
  MUX2_X1 U14464 ( .A(n12109), .B(n12108), .S(n12112), .Z(n12110) );
  INV_X1 U14465 ( .A(n12110), .ZN(n12151) );
  NAND2_X1 U14466 ( .A1(n12112), .A2(n12111), .ZN(n12148) );
  XOR2_X1 U14467 ( .A(n13870), .B(n13942), .Z(n12143) );
  INV_X1 U14468 ( .A(n12113), .ZN(n12114) );
  NOR2_X1 U14469 ( .A1(n12115), .A2(n12114), .ZN(n14133) );
  NOR4_X1 U14470 ( .A1(n12118), .A2(n12117), .A3(n12116), .A4(n14825), .ZN(
        n12122) );
  NAND4_X1 U14471 ( .A1(n12122), .A2(n12121), .A3(n12120), .A4(n12119), .ZN(
        n12123) );
  NOR4_X1 U14472 ( .A1(n12126), .A2(n12125), .A3(n12124), .A4(n12123), .ZN(
        n12129) );
  NAND4_X1 U14473 ( .A1(n12130), .A2(n12129), .A3(n12128), .A4(n12127), .ZN(
        n12131) );
  NOR3_X1 U14474 ( .A1(n14133), .A2(n12132), .A3(n12131), .ZN(n12135) );
  NAND4_X1 U14475 ( .A1(n12135), .A2(n12134), .A3(n12133), .A4(n6514), .ZN(
        n12136) );
  NOR4_X1 U14476 ( .A1(n8922), .A2(n7483), .A3(n12137), .A4(n12136), .ZN(
        n12138) );
  NAND4_X1 U14477 ( .A1(n14066), .A2(n12138), .A3(n14045), .A4(n14073), .ZN(
        n12139) );
  NOR4_X1 U14478 ( .A1(n13996), .A2(n14020), .A3(n14025), .A4(n12139), .ZN(
        n12140) );
  INV_X1 U14479 ( .A(n13971), .ZN(n13962) );
  NAND4_X1 U14480 ( .A1(n12141), .A2(n12140), .A3(n13962), .A4(n13981), .ZN(
        n12142) );
  NOR3_X1 U14481 ( .A1(n12144), .A2(n12143), .A3(n12142), .ZN(n12145) );
  XNOR2_X1 U14482 ( .A(n12145), .B(n13930), .ZN(n12146) );
  OAI22_X1 U14483 ( .A1(n12149), .A2(n12148), .B1(n12147), .B2(n12146), .ZN(
        n12150) );
  NOR2_X1 U14484 ( .A1(n6487), .A2(P1_U3086), .ZN(n12153) );
  NAND3_X1 U14485 ( .A1(n12154), .A2(n13861), .A3(n12153), .ZN(n12155) );
  OAI211_X1 U14486 ( .C1(n14348), .C2(n12157), .A(n12155), .B(P1_B_REG_SCAN_IN), .ZN(n12156) );
  INV_X1 U14487 ( .A(n12158), .ZN(n12160) );
  OAI222_X1 U14488 ( .A1(n12903), .A2(n12160), .B1(n12900), .B2(n12159), .C1(
        P3_U3151), .C2(n12506), .ZN(P3_U3268) );
  INV_X1 U14489 ( .A(n12161), .ZN(n12162) );
  XNOR2_X1 U14490 ( .A(n14490), .B(n10963), .ZN(n12164) );
  NAND2_X1 U14491 ( .A1(n12164), .A2(n12755), .ZN(n12308) );
  XNOR2_X1 U14492 ( .A(n12879), .B(n10712), .ZN(n12165) );
  XNOR2_X1 U14493 ( .A(n12165), .B(n14488), .ZN(n12231) );
  NAND2_X1 U14494 ( .A1(n12165), .A2(n12737), .ZN(n12166) );
  XNOR2_X1 U14495 ( .A(n12745), .B(n10963), .ZN(n12348) );
  NAND2_X1 U14496 ( .A1(n12348), .A2(n12726), .ZN(n12167) );
  INV_X1 U14497 ( .A(n12348), .ZN(n12168) );
  NAND2_X1 U14498 ( .A1(n12168), .A2(n12754), .ZN(n12169) );
  XNOR2_X1 U14499 ( .A(n12729), .B(n10712), .ZN(n12170) );
  XNOR2_X1 U14500 ( .A(n12170), .B(n12353), .ZN(n12273) );
  INV_X1 U14501 ( .A(n12170), .ZN(n12171) );
  XNOR2_X1 U14502 ( .A(n12715), .B(n10712), .ZN(n12172) );
  XNOR2_X1 U14503 ( .A(n12172), .B(n12725), .ZN(n12280) );
  NAND2_X1 U14504 ( .A1(n12172), .A2(n12691), .ZN(n12173) );
  XNOR2_X1 U14505 ( .A(n12699), .B(n10712), .ZN(n12175) );
  XNOR2_X1 U14506 ( .A(n12175), .B(n12366), .ZN(n12325) );
  INV_X1 U14507 ( .A(n12175), .ZN(n12176) );
  NAND2_X1 U14508 ( .A1(n12176), .A2(n12366), .ZN(n12177) );
  XNOR2_X1 U14509 ( .A(n12249), .B(n10712), .ZN(n12178) );
  XNOR2_X1 U14510 ( .A(n12178), .B(n12692), .ZN(n12244) );
  INV_X1 U14511 ( .A(n12178), .ZN(n12179) );
  XNOR2_X1 U14512 ( .A(n12855), .B(n10712), .ZN(n12180) );
  XNOR2_X1 U14513 ( .A(n12180), .B(n12679), .ZN(n12300) );
  NAND2_X1 U14514 ( .A1(n12180), .A2(n12365), .ZN(n12181) );
  XNOR2_X1 U14515 ( .A(n12792), .B(n10712), .ZN(n12182) );
  NAND2_X1 U14516 ( .A1(n12182), .A2(n12667), .ZN(n12183) );
  OAI21_X1 U14517 ( .B1(n12182), .B2(n12667), .A(n12183), .ZN(n12255) );
  XNOR2_X1 U14518 ( .A(n12646), .B(n10712), .ZN(n12184) );
  XNOR2_X1 U14519 ( .A(n12633), .B(n10712), .ZN(n12186) );
  XNOR2_X1 U14520 ( .A(n12841), .B(n10963), .ZN(n12188) );
  NAND2_X1 U14521 ( .A1(n12188), .A2(n12187), .ZN(n12267) );
  INV_X1 U14522 ( .A(n12188), .ZN(n12189) );
  NAND2_X1 U14523 ( .A1(n12189), .A2(n12626), .ZN(n12190) );
  NAND2_X1 U14524 ( .A1(n12191), .A2(n12289), .ZN(n12264) );
  NAND2_X1 U14525 ( .A1(n12264), .A2(n12267), .ZN(n12195) );
  XNOR2_X1 U14526 ( .A(n12776), .B(n10712), .ZN(n12192) );
  NAND2_X1 U14527 ( .A1(n12192), .A2(n12614), .ZN(n12196) );
  INV_X1 U14528 ( .A(n12192), .ZN(n12193) );
  NAND2_X1 U14529 ( .A1(n12193), .A2(n12582), .ZN(n12194) );
  AND2_X1 U14530 ( .A1(n12196), .A2(n12194), .ZN(n12265) );
  NAND2_X1 U14531 ( .A1(n12195), .A2(n12265), .ZN(n12269) );
  NAND2_X1 U14532 ( .A1(n12269), .A2(n12196), .ZN(n12338) );
  XNOR2_X1 U14533 ( .A(n12836), .B(n10712), .ZN(n12197) );
  NOR2_X1 U14534 ( .A1(n12197), .A2(n12597), .ZN(n12198) );
  AOI21_X1 U14535 ( .B1(n12197), .B2(n12597), .A(n12198), .ZN(n12339) );
  INV_X1 U14536 ( .A(n12198), .ZN(n12199) );
  XNOR2_X1 U14537 ( .A(n12575), .B(n10963), .ZN(n12200) );
  NOR2_X1 U14538 ( .A1(n12200), .A2(n12583), .ZN(n12201) );
  AOI21_X1 U14539 ( .B1(n12200), .B2(n12583), .A(n12201), .ZN(n12224) );
  XNOR2_X1 U14540 ( .A(n12202), .B(n10712), .ZN(n12203) );
  NOR2_X1 U14541 ( .A1(n12356), .A2(n12557), .ZN(n12207) );
  AOI22_X1 U14542 ( .A1(n12330), .A2(n12583), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12204) );
  OAI21_X1 U14543 ( .B1(n12205), .B2(n12328), .A(n12204), .ZN(n12206) );
  AOI211_X1 U14544 ( .C1(n12767), .C2(n12334), .A(n12207), .B(n12206), .ZN(
        n12208) );
  OAI21_X1 U14545 ( .B1(n12209), .B2(n12360), .A(n12208), .ZN(P3_U3160) );
  INV_X1 U14546 ( .A(n12210), .ZN(n12211) );
  OAI222_X1 U14547 ( .A1(n12900), .A2(n12212), .B1(n12903), .B2(n12211), .C1(
        n8450), .C2(P3_U3151), .ZN(P3_U3267) );
  OAI22_X1 U14548 ( .A1(n12749), .A2(n15272), .B1(n12213), .B2(n12746), .ZN(
        n12216) );
  NOR2_X1 U14549 ( .A1(n12214), .A2(n12663), .ZN(n12215) );
  AOI211_X1 U14550 ( .C1(n12660), .C2(n12217), .A(n12216), .B(n12215), .ZN(
        n12218) );
  OAI21_X1 U14551 ( .B1(n12219), .B2(n15194), .A(n12218), .ZN(P3_U3204) );
  INV_X1 U14552 ( .A(n12220), .ZN(n12221) );
  OAI222_X1 U14553 ( .A1(n12223), .A2(P3_U3151), .B1(n12900), .B2(n12222), 
        .C1(n12903), .C2(n12221), .ZN(P3_U3265) );
  INV_X1 U14554 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n12225) );
  OAI22_X1 U14555 ( .A1(n12328), .A2(n12226), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12225), .ZN(n12228) );
  NOR2_X1 U14556 ( .A1(n12356), .A2(n12572), .ZN(n12227) );
  AOI211_X1 U14557 ( .C1(n12330), .C2(n12597), .A(n12228), .B(n12227), .ZN(
        n12229) );
  OAI211_X1 U14558 ( .C1(n12232), .C2(n12231), .A(n12230), .B(n12340), .ZN(
        n12236) );
  AND2_X1 U14559 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12408) );
  AOI21_X1 U14560 ( .B1(n12330), .B2(n12755), .A(n12408), .ZN(n12233) );
  OAI21_X1 U14561 ( .B1(n12726), .B2(n12328), .A(n12233), .ZN(n12234) );
  AOI21_X1 U14562 ( .B1(n12297), .B2(n12759), .A(n12234), .ZN(n12235) );
  OAI211_X1 U14563 ( .C1(n12347), .C2(n12879), .A(n12236), .B(n12235), .ZN(
        P3_U3155) );
  INV_X1 U14564 ( .A(n12237), .ZN(n12291) );
  AOI21_X1 U14565 ( .B1(n12363), .B2(n12238), .A(n12291), .ZN(n12243) );
  AOI22_X1 U14566 ( .A1(n12330), .A2(n12627), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12240) );
  NAND2_X1 U14567 ( .A1(n12354), .A2(n12626), .ZN(n12239) );
  OAI211_X1 U14568 ( .C1(n12356), .C2(n12630), .A(n12240), .B(n12239), .ZN(
        n12241) );
  AOI21_X1 U14569 ( .B1(n12633), .B2(n12358), .A(n12241), .ZN(n12242) );
  OAI21_X1 U14570 ( .B1(n12243), .B2(n12360), .A(n12242), .ZN(P3_U3156) );
  XNOR2_X1 U14571 ( .A(n12245), .B(n12244), .ZN(n12251) );
  AND2_X1 U14572 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12543) );
  NOR2_X1 U14573 ( .A1(n12328), .A2(n12679), .ZN(n12246) );
  AOI211_X1 U14574 ( .C1(n12330), .C2(n12366), .A(n12543), .B(n12246), .ZN(
        n12247) );
  OAI21_X1 U14575 ( .B1(n12682), .B2(n12332), .A(n12247), .ZN(n12248) );
  AOI21_X1 U14576 ( .B1(n12249), .B2(n12358), .A(n12248), .ZN(n12250) );
  OAI21_X1 U14577 ( .B1(n12251), .B2(n12360), .A(n12250), .ZN(P3_U3159) );
  INV_X1 U14578 ( .A(n12252), .ZN(n12253) );
  AOI21_X1 U14579 ( .B1(n12255), .B2(n12254), .A(n12253), .ZN(n12261) );
  OAI22_X1 U14580 ( .A1(n12351), .A2(n12679), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12256), .ZN(n12257) );
  AOI21_X1 U14581 ( .B1(n12354), .B2(n12627), .A(n12257), .ZN(n12258) );
  OAI21_X1 U14582 ( .B1(n12657), .B2(n12356), .A(n12258), .ZN(n12259) );
  AOI21_X1 U14583 ( .B1(n12792), .B2(n12334), .A(n12259), .ZN(n12260) );
  OAI21_X1 U14584 ( .B1(n12261), .B2(n12360), .A(n12260), .ZN(P3_U3163) );
  AOI22_X1 U14585 ( .A1(n12330), .A2(n12626), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12263) );
  NAND2_X1 U14586 ( .A1(n12354), .A2(n12597), .ZN(n12262) );
  OAI211_X1 U14587 ( .C1(n12356), .C2(n12600), .A(n12263), .B(n12262), .ZN(
        n12271) );
  INV_X1 U14588 ( .A(n12265), .ZN(n12266) );
  NAND3_X1 U14589 ( .A1(n12264), .A2(n12267), .A3(n12266), .ZN(n12268) );
  AOI21_X1 U14590 ( .B1(n12269), .B2(n12268), .A(n12360), .ZN(n12270) );
  AOI211_X1 U14591 ( .C1(n12334), .C2(n12776), .A(n12271), .B(n12270), .ZN(
        n12272) );
  INV_X1 U14592 ( .A(n12272), .ZN(P3_U3165) );
  XNOR2_X1 U14593 ( .A(n12274), .B(n12273), .ZN(n12279) );
  AND2_X1 U14594 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12463) );
  NOR2_X1 U14595 ( .A1(n12328), .A2(n12725), .ZN(n12275) );
  AOI211_X1 U14596 ( .C1(n12330), .C2(n12754), .A(n12463), .B(n12275), .ZN(
        n12276) );
  OAI21_X1 U14597 ( .B1(n12730), .B2(n12356), .A(n12276), .ZN(n12277) );
  AOI21_X1 U14598 ( .B1(n12729), .B2(n12334), .A(n12277), .ZN(n12278) );
  OAI21_X1 U14599 ( .B1(n12279), .B2(n12360), .A(n12278), .ZN(P3_U3166) );
  XNOR2_X1 U14600 ( .A(n12281), .B(n12280), .ZN(n12287) );
  INV_X1 U14601 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n12282) );
  NOR2_X1 U14602 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12282), .ZN(n12487) );
  NOR2_X1 U14603 ( .A1(n12328), .A2(n12707), .ZN(n12283) );
  AOI211_X1 U14604 ( .C1(n12330), .C2(n12353), .A(n12487), .B(n12283), .ZN(
        n12284) );
  OAI21_X1 U14605 ( .B1(n12716), .B2(n12356), .A(n12284), .ZN(n12285) );
  AOI21_X1 U14606 ( .B1(n12866), .B2(n12358), .A(n12285), .ZN(n12286) );
  OAI21_X1 U14607 ( .B1(n12287), .B2(n12360), .A(n12286), .ZN(P3_U3168) );
  INV_X1 U14608 ( .A(n12288), .ZN(n12290) );
  NOR3_X1 U14609 ( .A1(n12291), .A2(n12290), .A3(n12289), .ZN(n12293) );
  INV_X1 U14610 ( .A(n12264), .ZN(n12292) );
  OAI21_X1 U14611 ( .B1(n12293), .B2(n12292), .A(n12340), .ZN(n12299) );
  AOI22_X1 U14612 ( .A1(n12330), .A2(n12363), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12294) );
  OAI21_X1 U14613 ( .B1(n12614), .B2(n12328), .A(n12294), .ZN(n12295) );
  AOI21_X1 U14614 ( .B1(n12297), .B2(n12296), .A(n12295), .ZN(n12298) );
  OAI211_X1 U14615 ( .C1(n12841), .C2(n12347), .A(n12299), .B(n12298), .ZN(
        P3_U3169) );
  XNOR2_X1 U14616 ( .A(n12301), .B(n12300), .ZN(n12307) );
  AOI22_X1 U14617 ( .A1(n12330), .A2(n12692), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12303) );
  NAND2_X1 U14618 ( .A1(n12354), .A2(n12364), .ZN(n12302) );
  OAI211_X1 U14619 ( .C1(n12332), .C2(n12672), .A(n12303), .B(n12302), .ZN(
        n12304) );
  AOI21_X1 U14620 ( .B1(n12305), .B2(n12358), .A(n12304), .ZN(n12306) );
  OAI21_X1 U14621 ( .B1(n12307), .B2(n12360), .A(n12306), .ZN(P3_U3173) );
  NAND2_X1 U14622 ( .A1(n6672), .A2(n12308), .ZN(n12309) );
  XNOR2_X1 U14623 ( .A(n12310), .B(n12309), .ZN(n12316) );
  NOR2_X1 U14624 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15429), .ZN(n12384) );
  NOR2_X1 U14625 ( .A1(n12328), .A2(n14488), .ZN(n12311) );
  AOI211_X1 U14626 ( .C1(n12330), .C2(n14497), .A(n12384), .B(n12311), .ZN(
        n12312) );
  OAI21_X1 U14627 ( .B1(n12313), .B2(n12356), .A(n12312), .ZN(n12314) );
  AOI21_X1 U14628 ( .B1(n12358), .B2(n14490), .A(n12314), .ZN(n12315) );
  OAI21_X1 U14629 ( .B1(n12316), .B2(n12360), .A(n12315), .ZN(P3_U3174) );
  AOI21_X1 U14630 ( .B1(n12627), .B2(n12318), .A(n7079), .ZN(n12324) );
  OAI22_X1 U14631 ( .A1(n12351), .A2(n12667), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12319), .ZN(n12320) );
  AOI21_X1 U14632 ( .B1(n12354), .B2(n12363), .A(n12320), .ZN(n12321) );
  OAI21_X1 U14633 ( .B1(n12643), .B2(n12356), .A(n12321), .ZN(n12322) );
  AOI21_X1 U14634 ( .B1(n12646), .B2(n12358), .A(n12322), .ZN(n12323) );
  OAI21_X1 U14635 ( .B1(n12324), .B2(n12360), .A(n12323), .ZN(P3_U3175) );
  XNOR2_X1 U14636 ( .A(n12326), .B(n12325), .ZN(n12336) );
  AND2_X1 U14637 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12514) );
  NOR2_X1 U14638 ( .A1(n12328), .A2(n12327), .ZN(n12329) );
  AOI211_X1 U14639 ( .C1(n12330), .C2(n12691), .A(n12514), .B(n12329), .ZN(
        n12331) );
  OAI21_X1 U14640 ( .B1(n12700), .B2(n12332), .A(n12331), .ZN(n12333) );
  AOI21_X1 U14641 ( .B1(n12699), .B2(n12334), .A(n12333), .ZN(n12335) );
  OAI21_X1 U14642 ( .B1(n12336), .B2(n12360), .A(n12335), .ZN(P3_U3178) );
  OAI21_X1 U14643 ( .B1(n12339), .B2(n12338), .A(n12337), .ZN(n12341) );
  NAND2_X1 U14644 ( .A1(n12341), .A2(n12340), .ZN(n12346) );
  OAI22_X1 U14645 ( .A1(n12351), .A2(n12614), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12342), .ZN(n12344) );
  NOR2_X1 U14646 ( .A1(n12356), .A2(n12587), .ZN(n12343) );
  AOI211_X1 U14647 ( .C1(n12354), .C2(n12583), .A(n12344), .B(n12343), .ZN(
        n12345) );
  OAI211_X1 U14648 ( .C1(n12836), .C2(n12347), .A(n12346), .B(n12345), .ZN(
        P3_U3180) );
  XNOR2_X1 U14649 ( .A(n12348), .B(n12754), .ZN(n12349) );
  XNOR2_X1 U14650 ( .A(n12350), .B(n12349), .ZN(n12361) );
  OR2_X1 U14651 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15410), .ZN(n12433) );
  OAI21_X1 U14652 ( .B1(n12351), .B2(n14488), .A(n12433), .ZN(n12352) );
  AOI21_X1 U14653 ( .B1(n12354), .B2(n12353), .A(n12352), .ZN(n12355) );
  OAI21_X1 U14654 ( .B1(n12747), .B2(n12356), .A(n12355), .ZN(n12357) );
  AOI21_X1 U14655 ( .B1(n12873), .B2(n12358), .A(n12357), .ZN(n12359) );
  OAI21_X1 U14656 ( .B1(n12361), .B2(n12360), .A(n12359), .ZN(P3_U3181) );
  MUX2_X1 U14657 ( .A(n12552), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12375), .Z(
        P3_U3522) );
  MUX2_X1 U14658 ( .A(n12362), .B(P3_DATAO_REG_30__SCAN_IN), .S(n12375), .Z(
        P3_U3521) );
  MUX2_X1 U14659 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12570), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14660 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12583), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14661 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12597), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14662 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12582), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14663 ( .A(n12626), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12375), .Z(
        P3_U3515) );
  MUX2_X1 U14664 ( .A(n12363), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12375), .Z(
        P3_U3514) );
  MUX2_X1 U14665 ( .A(n12627), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12375), .Z(
        P3_U3513) );
  MUX2_X1 U14666 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12364), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14667 ( .A(n12365), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12375), .Z(
        P3_U3511) );
  MUX2_X1 U14668 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12692), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14669 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12366), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14670 ( .A(n12691), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12375), .Z(
        P3_U3508) );
  MUX2_X1 U14671 ( .A(n12754), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12375), .Z(
        P3_U3506) );
  MUX2_X1 U14672 ( .A(n12737), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12375), .Z(
        P3_U3505) );
  MUX2_X1 U14673 ( .A(n12755), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12375), .Z(
        P3_U3504) );
  MUX2_X1 U14674 ( .A(n14497), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12375), .Z(
        P3_U3503) );
  MUX2_X1 U14675 ( .A(n12367), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12375), .Z(
        P3_U3502) );
  MUX2_X1 U14676 ( .A(n14496), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12375), .Z(
        P3_U3501) );
  MUX2_X1 U14677 ( .A(n12368), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12375), .Z(
        P3_U3500) );
  MUX2_X1 U14678 ( .A(n12369), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12375), .Z(
        P3_U3499) );
  MUX2_X1 U14679 ( .A(n12370), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12375), .Z(
        P3_U3498) );
  MUX2_X1 U14680 ( .A(n12371), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12375), .Z(
        P3_U3497) );
  MUX2_X1 U14681 ( .A(n12372), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12375), .Z(
        P3_U3496) );
  MUX2_X1 U14682 ( .A(n12373), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12375), .Z(
        P3_U3495) );
  MUX2_X1 U14683 ( .A(n15201), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12375), .Z(
        P3_U3493) );
  MUX2_X1 U14684 ( .A(n12374), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12375), .Z(
        P3_U3492) );
  MUX2_X1 U14685 ( .A(n15202), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12375), .Z(
        P3_U3491) );
  NOR2_X1 U14686 ( .A1(n12377), .A2(n12376), .ZN(n12378) );
  NAND2_X1 U14687 ( .A1(n12380), .A2(n12388), .ZN(n12400) );
  AOI21_X1 U14688 ( .B1(n12381), .B2(n8014), .A(n12401), .ZN(n12399) );
  INV_X1 U14689 ( .A(n12388), .ZN(n12414) );
  AOI21_X1 U14690 ( .B1(n12383), .B2(n12385), .A(n12405), .ZN(n12396) );
  AOI21_X1 U14691 ( .B1(n15168), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12384), 
        .ZN(n12395) );
  OR2_X1 U14692 ( .A1(n12506), .A2(n12385), .ZN(n12387) );
  NAND2_X1 U14693 ( .A1(n12506), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n12386) );
  AND2_X1 U14694 ( .A1(n12387), .A2(n12386), .ZN(n12415) );
  XNOR2_X1 U14695 ( .A(n12415), .B(n12388), .ZN(n12392) );
  NOR2_X1 U14696 ( .A1(n12390), .A2(n12389), .ZN(n12391) );
  NAND2_X1 U14697 ( .A1(n12392), .A2(n12391), .ZN(n12412) );
  OAI21_X1 U14698 ( .B1(n12392), .B2(n12391), .A(n12412), .ZN(n12393) );
  NAND2_X1 U14699 ( .A1(n15173), .A2(n12393), .ZN(n12394) );
  OAI211_X1 U14700 ( .C1(n12396), .C2(n15162), .A(n12395), .B(n12394), .ZN(
        n12397) );
  AOI21_X1 U14701 ( .B1(n12414), .B2(n15175), .A(n12397), .ZN(n12398) );
  OAI21_X1 U14702 ( .B1(n12399), .B2(n15164), .A(n12398), .ZN(P3_U3195) );
  INV_X1 U14703 ( .A(n12400), .ZN(n12402) );
  XNOR2_X1 U14704 ( .A(n12436), .B(n12827), .ZN(n12410) );
  INV_X1 U14705 ( .A(n12410), .ZN(n12403) );
  AOI21_X1 U14706 ( .B1(n12404), .B2(n12403), .A(n12425), .ZN(n12424) );
  XNOR2_X1 U14707 ( .A(n12436), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n12409) );
  NOR2_X1 U14708 ( .A1(n12406), .A2(n12405), .ZN(n12407) );
  AOI21_X1 U14709 ( .B1(n12409), .B2(n12407), .A(n12428), .ZN(n12420) );
  AOI21_X1 U14710 ( .B1(n15168), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12408), 
        .ZN(n12419) );
  INV_X1 U14711 ( .A(n12409), .ZN(n12411) );
  MUX2_X1 U14712 ( .A(n12411), .B(n12410), .S(n12506), .Z(n12417) );
  INV_X1 U14713 ( .A(n12412), .ZN(n12413) );
  NAND2_X1 U14714 ( .A1(n12416), .A2(n12417), .ZN(n12439) );
  OAI211_X1 U14715 ( .C1(n12417), .C2(n12416), .A(n15173), .B(n12439), .ZN(
        n12418) );
  OAI211_X1 U14716 ( .C1(n12420), .C2(n15162), .A(n12419), .B(n12418), .ZN(
        n12421) );
  AOI21_X1 U14717 ( .B1(n12422), .B2(n15175), .A(n12421), .ZN(n12423) );
  OAI21_X1 U14718 ( .B1(n12424), .B2(n15164), .A(n12423), .ZN(P3_U3196) );
  AOI21_X1 U14719 ( .B1(n12427), .B2(n12426), .A(n12451), .ZN(n12449) );
  INV_X1 U14720 ( .A(n12430), .ZN(n12429) );
  NOR2_X1 U14721 ( .A1(n12429), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n12432) );
  OAI21_X1 U14722 ( .B1(n12432), .B2(n12457), .A(n12431), .ZN(n12448) );
  INV_X1 U14723 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14385) );
  OAI21_X1 U14724 ( .B1(n15156), .B2(n14385), .A(n12433), .ZN(n12446) );
  OR2_X1 U14725 ( .A1(n12506), .A2(n12748), .ZN(n12435) );
  NAND2_X1 U14726 ( .A1(n12506), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n12434) );
  AND2_X1 U14727 ( .A1(n12435), .A2(n12434), .ZN(n12444) );
  NAND2_X1 U14728 ( .A1(n12506), .A2(n12827), .ZN(n12437) );
  OAI211_X1 U14729 ( .C1(n12506), .C2(P3_REG2_REG_14__SCAN_IN), .A(n12437), 
        .B(n12436), .ZN(n12438) );
  NAND2_X1 U14730 ( .A1(n12439), .A2(n12438), .ZN(n12441) );
  AND2_X1 U14731 ( .A1(n12441), .A2(n12440), .ZN(n12469) );
  NOR2_X1 U14732 ( .A1(n12441), .A2(n12440), .ZN(n12442) );
  AOI211_X1 U14733 ( .C1(n12444), .C2(n12443), .A(n15150), .B(n12468), .ZN(
        n12445) );
  AOI211_X1 U14734 ( .C1(n15175), .C2(n12456), .A(n12446), .B(n12445), .ZN(
        n12447) );
  OAI211_X1 U14735 ( .C1(n12449), .C2(n15164), .A(n12448), .B(n12447), .ZN(
        P3_U3197) );
  NOR2_X1 U14736 ( .A1(n12456), .A2(n12450), .ZN(n12452) );
  AOI22_X1 U14737 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12459), .B1(n12483), 
        .B2(n12817), .ZN(n12453) );
  AOI21_X1 U14738 ( .B1(n12454), .B2(n12453), .A(n12482), .ZN(n12479) );
  NOR2_X1 U14739 ( .A1(n12456), .A2(n12455), .ZN(n12458) );
  AOI22_X1 U14740 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12459), .B1(n12483), 
        .B2(n12731), .ZN(n12460) );
  AOI21_X1 U14741 ( .B1(n12461), .B2(n12460), .A(n12480), .ZN(n12462) );
  NOR2_X1 U14742 ( .A1(n12462), .A2(n15162), .ZN(n12477) );
  AOI21_X1 U14743 ( .B1(n15168), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n12463), 
        .ZN(n12475) );
  OR2_X1 U14744 ( .A1(n12506), .A2(n12731), .ZN(n12465) );
  NAND2_X1 U14745 ( .A1(n12506), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n12464) );
  NAND2_X1 U14746 ( .A1(n12465), .A2(n12464), .ZN(n12466) );
  AND2_X1 U14747 ( .A1(n12466), .A2(n12483), .ZN(n12489) );
  NOR2_X1 U14748 ( .A1(n12466), .A2(n12483), .ZN(n12467) );
  OR2_X1 U14749 ( .A1(n12489), .A2(n12467), .ZN(n12470) );
  NOR2_X1 U14750 ( .A1(n12469), .A2(n12468), .ZN(n12471) );
  NAND2_X1 U14751 ( .A1(n12470), .A2(n12471), .ZN(n12473) );
  INV_X1 U14752 ( .A(n12488), .ZN(n12472) );
  NAND3_X1 U14753 ( .A1(n15173), .A2(n12473), .A3(n12472), .ZN(n12474) );
  OAI211_X1 U14754 ( .C1(n15147), .C2(n12483), .A(n12475), .B(n12474), .ZN(
        n12476) );
  NOR2_X1 U14755 ( .A1(n12477), .A2(n12476), .ZN(n12478) );
  OAI21_X1 U14756 ( .B1(n12479), .B2(n15164), .A(n12478), .ZN(P3_U3198) );
  AOI21_X1 U14757 ( .B1(n12481), .B2(n12717), .A(n12502), .ZN(n12500) );
  NOR2_X1 U14758 ( .A1(n12485), .A2(n12484), .ZN(n12518) );
  AOI21_X1 U14759 ( .B1(n12485), .B2(n12484), .A(n12518), .ZN(n12486) );
  NOR2_X1 U14760 ( .A1(n12486), .A2(n15164), .ZN(n12498) );
  AOI21_X1 U14761 ( .B1(n15168), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n12487), 
        .ZN(n12496) );
  NOR2_X1 U14762 ( .A1(n12489), .A2(n12488), .ZN(n12492) );
  OR2_X1 U14763 ( .A1(n12506), .A2(n12717), .ZN(n12491) );
  NAND2_X1 U14764 ( .A1(n12506), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n12490) );
  NAND2_X1 U14765 ( .A1(n12491), .A2(n12490), .ZN(n12510) );
  XNOR2_X1 U14766 ( .A(n12510), .B(n12509), .ZN(n12493) );
  NAND2_X1 U14767 ( .A1(n12493), .A2(n12492), .ZN(n12494) );
  NAND3_X1 U14768 ( .A1(n15173), .A2(n6531), .A3(n12494), .ZN(n12495) );
  OAI211_X1 U14769 ( .C1(n15147), .C2(n12509), .A(n12496), .B(n12495), .ZN(
        n12497) );
  NOR2_X1 U14770 ( .A1(n12498), .A2(n12497), .ZN(n12499) );
  OAI21_X1 U14771 ( .B1(n12500), .B2(n15162), .A(n12499), .ZN(P3_U3199) );
  NOR2_X1 U14772 ( .A1(n12517), .A2(n12501), .ZN(n12503) );
  NAND2_X1 U14773 ( .A1(n12520), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12527) );
  OAI21_X1 U14774 ( .B1(n12520), .B2(P3_REG2_REG_18__SCAN_IN), .A(n12527), 
        .ZN(n12504) );
  AOI21_X1 U14775 ( .B1(n12505), .B2(n12504), .A(n12529), .ZN(n12526) );
  OR2_X1 U14776 ( .A1(n12506), .A2(n12701), .ZN(n12508) );
  NAND2_X1 U14777 ( .A1(n12506), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n12507) );
  AND2_X1 U14778 ( .A1(n12508), .A2(n12507), .ZN(n12513) );
  NAND2_X1 U14779 ( .A1(n12510), .A2(n12509), .ZN(n12511) );
  NAND2_X1 U14780 ( .A1(n12511), .A2(n6531), .ZN(n12532) );
  INV_X1 U14781 ( .A(n12520), .ZN(n12533) );
  XNOR2_X1 U14782 ( .A(n12532), .B(n12533), .ZN(n12512) );
  NAND2_X1 U14783 ( .A1(n12512), .A2(n12513), .ZN(n12536) );
  OAI21_X1 U14784 ( .B1(n12513), .B2(n12512), .A(n12536), .ZN(n12524) );
  AOI21_X1 U14785 ( .B1(n15168), .B2(P3_ADDR_REG_18__SCAN_IN), .A(n12514), 
        .ZN(n12515) );
  OAI21_X1 U14786 ( .B1(n15147), .B2(n12520), .A(n12515), .ZN(n12523) );
  NOR2_X1 U14787 ( .A1(n12517), .A2(n12516), .ZN(n12519) );
  NOR2_X1 U14788 ( .A1(n12519), .A2(n12518), .ZN(n12522) );
  NAND2_X1 U14789 ( .A1(n12520), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n12530) );
  OAI21_X1 U14790 ( .B1(n12520), .B2(P3_REG1_REG_18__SCAN_IN), .A(n12530), 
        .ZN(n12521) );
  OAI21_X1 U14791 ( .B1(n12526), .B2(n15162), .A(n12525), .ZN(P3_U3200) );
  INV_X1 U14792 ( .A(n12527), .ZN(n12528) );
  MUX2_X1 U14793 ( .A(n12683), .B(P3_REG2_REG_19__SCAN_IN), .S(n12531), .Z(
        n12540) );
  XNOR2_X1 U14794 ( .A(n12531), .B(n12803), .ZN(n12537) );
  INV_X1 U14795 ( .A(n12532), .ZN(n12534) );
  NAND2_X1 U14796 ( .A1(n12534), .A2(n12533), .ZN(n12535) );
  NAND2_X1 U14797 ( .A1(n12536), .A2(n12535), .ZN(n12542) );
  NAND2_X1 U14798 ( .A1(n12506), .A2(n12537), .ZN(n12538) );
  OAI21_X1 U14799 ( .B1(n12540), .B2(n12506), .A(n12538), .ZN(n12541) );
  AOI21_X1 U14800 ( .B1(n15168), .B2(P3_ADDR_REG_19__SCAN_IN), .A(n12543), 
        .ZN(n12544) );
  OAI21_X1 U14801 ( .B1(n15147), .B2(n12545), .A(n12544), .ZN(n12546) );
  NAND2_X1 U14802 ( .A1(n12549), .A2(n15209), .ZN(n12553) );
  INV_X1 U14803 ( .A(n12550), .ZN(n12551) );
  NAND2_X1 U14804 ( .A1(n12552), .A2(n12551), .ZN(n14514) );
  AOI21_X1 U14805 ( .B1(n12553), .B2(n14514), .A(n15214), .ZN(n12556) );
  AOI21_X1 U14806 ( .B1(P3_REG2_REG_31__SCAN_IN), .B2(n15214), .A(n12556), 
        .ZN(n12554) );
  OAI21_X1 U14807 ( .B1(n14512), .B2(n12761), .A(n12554), .ZN(P3_U3202) );
  OAI22_X1 U14808 ( .A1(n12761), .A2(n14515), .B1(n15412), .B2(n12749), .ZN(
        n12555) );
  OR2_X1 U14809 ( .A1(n12556), .A2(n12555), .ZN(P3_U3203) );
  OAI22_X1 U14810 ( .A1(n12749), .A2(n12558), .B1(n12557), .B2(n12746), .ZN(
        n12561) );
  NOR2_X1 U14811 ( .A1(n12559), .A2(n12663), .ZN(n12560) );
  AOI211_X1 U14812 ( .C1(n12660), .C2(n12767), .A(n12561), .B(n12560), .ZN(
        n12562) );
  OAI21_X1 U14813 ( .B1(n12563), .B2(n15194), .A(n12562), .ZN(P3_U3205) );
  AOI21_X1 U14814 ( .B1(n12565), .B2(n12567), .A(n12564), .ZN(n12768) );
  OAI21_X1 U14815 ( .B1(n12568), .B2(n12567), .A(n12566), .ZN(n12569) );
  AOI22_X1 U14816 ( .A1(n15203), .A2(n12597), .B1(n12570), .B2(n15200), .ZN(
        n12571) );
  NAND2_X1 U14817 ( .A1(n12769), .A2(n12749), .ZN(n12577) );
  OAI22_X1 U14818 ( .A1(n12718), .A2(n12573), .B1(n12572), .B2(n12746), .ZN(
        n12574) );
  AOI21_X1 U14819 ( .B1(n12575), .B2(n12660), .A(n12574), .ZN(n12576) );
  OAI211_X1 U14820 ( .C1(n12768), .C2(n12593), .A(n12577), .B(n12576), .ZN(
        P3_U3206) );
  XOR2_X1 U14821 ( .A(n12579), .B(n12578), .Z(n12771) );
  XNOR2_X1 U14822 ( .A(n12580), .B(n12579), .ZN(n12581) );
  NAND2_X1 U14823 ( .A1(n12581), .A2(n14499), .ZN(n12585) );
  AOI22_X1 U14824 ( .A1(n15200), .A2(n12583), .B1(n12582), .B2(n15203), .ZN(
        n12584) );
  OAI211_X1 U14825 ( .C1(n12586), .C2(n12771), .A(n12585), .B(n12584), .ZN(
        n12772) );
  NAND2_X1 U14826 ( .A1(n12772), .A2(n12749), .ZN(n12592) );
  OAI22_X1 U14827 ( .A1(n12718), .A2(n12588), .B1(n12587), .B2(n12746), .ZN(
        n12589) );
  AOI21_X1 U14828 ( .B1(n12590), .B2(n12660), .A(n12589), .ZN(n12591) );
  OAI211_X1 U14829 ( .C1(n12771), .C2(n12593), .A(n12592), .B(n12591), .ZN(
        P3_U3207) );
  OAI211_X1 U14830 ( .C1(n12596), .C2(n12595), .A(n12594), .B(n14499), .ZN(
        n12599) );
  AOI22_X1 U14831 ( .A1(n12597), .A2(n15200), .B1(n15203), .B2(n12626), .ZN(
        n12598) );
  OAI22_X1 U14832 ( .A1(n12718), .A2(n12601), .B1(n12600), .B2(n12746), .ZN(
        n12605) );
  XNOR2_X1 U14833 ( .A(n12603), .B(n12602), .ZN(n12779) );
  NOR2_X1 U14834 ( .A1(n12779), .A2(n12663), .ZN(n12604) );
  AOI211_X1 U14835 ( .C1(n12660), .C2(n12776), .A(n12605), .B(n12604), .ZN(
        n12606) );
  OAI21_X1 U14836 ( .B1(n12778), .B2(n15214), .A(n12606), .ZN(P3_U3208) );
  AOI21_X1 U14837 ( .B1(n12609), .B2(n12608), .A(n12607), .ZN(n12780) );
  AOI21_X1 U14838 ( .B1(n12612), .B2(n12611), .A(n12610), .ZN(n12613) );
  OAI222_X1 U14839 ( .A1(n15182), .A2(n12614), .B1(n15183), .B2(n12642), .C1(
        n15206), .C2(n12613), .ZN(n12781) );
  NAND2_X1 U14840 ( .A1(n12781), .A2(n12718), .ZN(n12620) );
  OAI22_X1 U14841 ( .A1(n12718), .A2(n12616), .B1(n12615), .B2(n12746), .ZN(
        n12617) );
  AOI21_X1 U14842 ( .B1(n12618), .B2(n12660), .A(n12617), .ZN(n12619) );
  OAI211_X1 U14843 ( .C1(n12780), .C2(n12663), .A(n12620), .B(n12619), .ZN(
        P3_U3209) );
  XNOR2_X1 U14844 ( .A(n12622), .B(n12621), .ZN(n12786) );
  INV_X1 U14845 ( .A(n12786), .ZN(n12636) );
  OAI211_X1 U14846 ( .C1(n12625), .C2(n12624), .A(n12623), .B(n14499), .ZN(
        n12629) );
  AOI22_X1 U14847 ( .A1(n15203), .A2(n12627), .B1(n12626), .B2(n15200), .ZN(
        n12628) );
  NAND2_X1 U14848 ( .A1(n12629), .A2(n12628), .ZN(n12785) );
  NAND2_X1 U14849 ( .A1(n12785), .A2(n12718), .ZN(n12635) );
  OAI22_X1 U14850 ( .A1(n12718), .A2(n12631), .B1(n12630), .B2(n12746), .ZN(
        n12632) );
  AOI21_X1 U14851 ( .B1(n12633), .B2(n12660), .A(n12632), .ZN(n12634) );
  OAI211_X1 U14852 ( .C1(n12663), .C2(n12636), .A(n12635), .B(n12634), .ZN(
        P3_U3210) );
  XNOR2_X1 U14853 ( .A(n12638), .B(n12637), .ZN(n12789) );
  INV_X1 U14854 ( .A(n12789), .ZN(n12649) );
  XNOR2_X1 U14855 ( .A(n12639), .B(n12640), .ZN(n12641) );
  OAI222_X1 U14856 ( .A1(n15183), .A2(n12667), .B1(n15182), .B2(n12642), .C1(
        n15206), .C2(n12641), .ZN(n12788) );
  NAND2_X1 U14857 ( .A1(n12788), .A2(n12718), .ZN(n12648) );
  OAI22_X1 U14858 ( .A1(n12718), .A2(n12644), .B1(n12643), .B2(n12746), .ZN(
        n12645) );
  AOI21_X1 U14859 ( .B1(n12646), .B2(n12660), .A(n12645), .ZN(n12647) );
  OAI211_X1 U14860 ( .C1(n12649), .C2(n12663), .A(n12648), .B(n12647), .ZN(
        P3_U3211) );
  XNOR2_X1 U14861 ( .A(n12650), .B(n12654), .ZN(n12794) );
  INV_X1 U14862 ( .A(n12794), .ZN(n12664) );
  AOI21_X1 U14863 ( .B1(n12654), .B2(n12651), .A(n12653), .ZN(n12655) );
  OAI222_X1 U14864 ( .A1(n15182), .A2(n12656), .B1(n15183), .B2(n12679), .C1(
        n15206), .C2(n12655), .ZN(n12793) );
  NAND2_X1 U14865 ( .A1(n12793), .A2(n12749), .ZN(n12662) );
  OAI22_X1 U14866 ( .A1(n12718), .A2(n12658), .B1(n12657), .B2(n12746), .ZN(
        n12659) );
  AOI21_X1 U14867 ( .B1(n12792), .B2(n12660), .A(n12659), .ZN(n12661) );
  OAI211_X1 U14868 ( .C1(n12664), .C2(n12663), .A(n12662), .B(n12661), .ZN(
        P3_U3212) );
  XNOR2_X1 U14869 ( .A(n12665), .B(n12670), .ZN(n12669) );
  NAND2_X1 U14870 ( .A1(n12692), .A2(n15203), .ZN(n12666) );
  OAI21_X1 U14871 ( .B1(n12667), .B2(n15182), .A(n12666), .ZN(n12668) );
  AOI21_X1 U14872 ( .B1(n12669), .B2(n14499), .A(n12668), .ZN(n12799) );
  XNOR2_X1 U14873 ( .A(n12671), .B(n12670), .ZN(n12797) );
  NOR2_X1 U14874 ( .A1(n12855), .A2(n12761), .ZN(n12675) );
  OAI22_X1 U14875 ( .A1(n12718), .A2(n12673), .B1(n12672), .B2(n12746), .ZN(
        n12674) );
  AOI211_X1 U14876 ( .C1(n12797), .C2(n14509), .A(n12675), .B(n12674), .ZN(
        n12676) );
  OAI21_X1 U14877 ( .B1(n12799), .B2(n15214), .A(n12676), .ZN(P3_U3213) );
  XNOR2_X1 U14878 ( .A(n12677), .B(n12680), .ZN(n12678) );
  OAI222_X1 U14879 ( .A1(n15182), .A2(n12679), .B1(n15183), .B2(n12707), .C1(
        n12678), .C2(n15206), .ZN(n12801) );
  INV_X1 U14880 ( .A(n12801), .ZN(n12687) );
  XNOR2_X1 U14881 ( .A(n12681), .B(n12680), .ZN(n12802) );
  NOR2_X1 U14882 ( .A1(n12859), .A2(n12761), .ZN(n12685) );
  OAI22_X1 U14883 ( .A1(n12718), .A2(n12683), .B1(n12682), .B2(n12746), .ZN(
        n12684) );
  AOI211_X1 U14884 ( .C1(n12802), .C2(n14509), .A(n12685), .B(n12684), .ZN(
        n12686) );
  OAI21_X1 U14885 ( .B1(n12687), .B2(n15214), .A(n12686), .ZN(P3_U3214) );
  OAI21_X1 U14886 ( .B1(n12690), .B2(n12689), .A(n12688), .ZN(n12693) );
  AOI222_X1 U14887 ( .A1(n14499), .A2(n12693), .B1(n12692), .B2(n15200), .C1(
        n12691), .C2(n15203), .ZN(n12805) );
  INV_X1 U14888 ( .A(n12694), .ZN(n12698) );
  AOI21_X1 U14889 ( .B1(n12714), .B2(n12696), .A(n12695), .ZN(n12697) );
  NOR2_X1 U14890 ( .A1(n12698), .A2(n12697), .ZN(n12807) );
  INV_X1 U14891 ( .A(n12699), .ZN(n12863) );
  NOR2_X1 U14892 ( .A1(n12863), .A2(n12761), .ZN(n12703) );
  OAI22_X1 U14893 ( .A1(n12718), .A2(n12701), .B1(n12700), .B2(n12746), .ZN(
        n12702) );
  AOI211_X1 U14894 ( .C1(n12807), .C2(n14509), .A(n12703), .B(n12702), .ZN(
        n12704) );
  OAI21_X1 U14895 ( .B1(n12805), .B2(n15214), .A(n12704), .ZN(P3_U3215) );
  NAND2_X1 U14896 ( .A1(n12705), .A2(n12711), .ZN(n12706) );
  NAND3_X1 U14897 ( .A1(n6650), .A2(n14499), .A3(n12706), .ZN(n12710) );
  OAI22_X1 U14898 ( .A1(n15441), .A2(n15183), .B1(n12707), .B2(n15182), .ZN(
        n12708) );
  INV_X1 U14899 ( .A(n12708), .ZN(n12709) );
  AND2_X1 U14900 ( .A1(n12710), .A2(n12709), .ZN(n12812) );
  OR2_X1 U14901 ( .A1(n12712), .A2(n12711), .ZN(n12713) );
  NAND2_X1 U14902 ( .A1(n12714), .A2(n12713), .ZN(n12810) );
  NOR2_X1 U14903 ( .A1(n12715), .A2(n12761), .ZN(n12720) );
  OAI22_X1 U14904 ( .A1(n12718), .A2(n12717), .B1(n12716), .B2(n12746), .ZN(
        n12719) );
  AOI211_X1 U14905 ( .C1(n12810), .C2(n14509), .A(n12720), .B(n12719), .ZN(
        n12721) );
  OAI21_X1 U14906 ( .B1(n12812), .B2(n15214), .A(n12721), .ZN(P3_U3216) );
  XNOR2_X1 U14907 ( .A(n12723), .B(n12722), .ZN(n12724) );
  OAI222_X1 U14908 ( .A1(n15183), .A2(n12726), .B1(n15182), .B2(n12725), .C1(
        n12724), .C2(n15206), .ZN(n12815) );
  INV_X1 U14909 ( .A(n12815), .ZN(n12735) );
  XNOR2_X1 U14910 ( .A(n12728), .B(n12727), .ZN(n12816) );
  NOR2_X1 U14911 ( .A1(n7672), .A2(n12761), .ZN(n12733) );
  OAI22_X1 U14912 ( .A1(n12749), .A2(n12731), .B1(n12730), .B2(n12746), .ZN(
        n12732) );
  AOI211_X1 U14913 ( .C1(n12816), .C2(n14509), .A(n12733), .B(n12732), .ZN(
        n12734) );
  OAI21_X1 U14914 ( .B1(n12735), .B2(n15214), .A(n12734), .ZN(P3_U3217) );
  XNOR2_X1 U14915 ( .A(n12736), .B(n12741), .ZN(n12740) );
  NAND2_X1 U14916 ( .A1(n12737), .A2(n15203), .ZN(n12738) );
  OAI21_X1 U14917 ( .B1(n15441), .B2(n15182), .A(n12738), .ZN(n12739) );
  AOI21_X1 U14918 ( .B1(n12740), .B2(n14499), .A(n12739), .ZN(n12821) );
  OR2_X1 U14919 ( .A1(n12742), .A2(n12741), .ZN(n12743) );
  NAND2_X1 U14920 ( .A1(n12744), .A2(n12743), .ZN(n12819) );
  NOR2_X1 U14921 ( .A1(n12745), .A2(n12761), .ZN(n12751) );
  OAI22_X1 U14922 ( .A1(n12749), .A2(n12748), .B1(n12747), .B2(n12746), .ZN(
        n12750) );
  AOI211_X1 U14923 ( .C1(n12819), .C2(n14509), .A(n12751), .B(n12750), .ZN(
        n12752) );
  OAI21_X1 U14924 ( .B1(n12821), .B2(n15194), .A(n12752), .ZN(P3_U3218) );
  OAI211_X1 U14925 ( .C1(n6646), .C2(n6515), .A(n14499), .B(n12753), .ZN(
        n12757) );
  AOI22_X1 U14926 ( .A1(n15203), .A2(n12755), .B1(n12754), .B2(n15200), .ZN(
        n12756) );
  NAND2_X1 U14927 ( .A1(n12757), .A2(n12756), .ZN(n12825) );
  INV_X1 U14928 ( .A(n12825), .ZN(n12764) );
  XNOR2_X1 U14929 ( .A(n12758), .B(n6515), .ZN(n12826) );
  AOI22_X1 U14930 ( .A1(n15214), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15209), 
        .B2(n12759), .ZN(n12760) );
  OAI21_X1 U14931 ( .B1(n12879), .B2(n12761), .A(n12760), .ZN(n12762) );
  AOI21_X1 U14932 ( .B1(n12826), .B2(n14509), .A(n12762), .ZN(n12763) );
  OAI21_X1 U14933 ( .B1(n12764), .B2(n15214), .A(n12763), .ZN(P3_U3219) );
  INV_X1 U14934 ( .A(n12829), .ZN(n12823) );
  INV_X1 U14935 ( .A(n15254), .ZN(n12766) );
  OAI21_X1 U14936 ( .B1(n12832), .B2(n12829), .A(n12770), .ZN(P3_U3486) );
  INV_X1 U14937 ( .A(n12771), .ZN(n12773) );
  AOI21_X1 U14938 ( .B1(n15242), .B2(n12773), .A(n12772), .ZN(n12833) );
  MUX2_X1 U14939 ( .A(n12774), .B(n12833), .S(n15254), .Z(n12775) );
  OAI21_X1 U14940 ( .B1(n12836), .B2(n12829), .A(n12775), .ZN(P3_U3485) );
  NAND2_X1 U14941 ( .A1(n12776), .A2(n15188), .ZN(n12777) );
  OAI211_X1 U14942 ( .C1(n14521), .C2(n12779), .A(n12778), .B(n12777), .ZN(
        n12837) );
  MUX2_X1 U14943 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n12837), .S(n15254), .Z(
        P3_U3484) );
  INV_X1 U14944 ( .A(n12780), .ZN(n12782) );
  AOI21_X1 U14945 ( .B1(n8531), .B2(n12782), .A(n12781), .ZN(n12838) );
  MUX2_X1 U14946 ( .A(n12783), .B(n12838), .S(n15254), .Z(n12784) );
  OAI21_X1 U14947 ( .B1(n12841), .B2(n12829), .A(n12784), .ZN(P3_U3483) );
  AOI21_X1 U14948 ( .B1(n12786), .B2(n8531), .A(n12785), .ZN(n12842) );
  MUX2_X1 U14949 ( .A(n15390), .B(n12842), .S(n15254), .Z(n12787) );
  OAI21_X1 U14950 ( .B1(n12845), .B2(n12829), .A(n12787), .ZN(P3_U3482) );
  AOI21_X1 U14951 ( .B1(n8531), .B2(n12789), .A(n12788), .ZN(n12846) );
  MUX2_X1 U14952 ( .A(n12790), .B(n12846), .S(n15254), .Z(n12791) );
  OAI21_X1 U14953 ( .B1(n12849), .B2(n12829), .A(n12791), .ZN(P3_U3481) );
  AOI21_X1 U14954 ( .B1(n8531), .B2(n12794), .A(n12793), .ZN(n12850) );
  MUX2_X1 U14955 ( .A(n12795), .B(n12850), .S(n15254), .Z(n12796) );
  OAI21_X1 U14956 ( .B1(n8512), .B2(n12829), .A(n12796), .ZN(P3_U3480) );
  NAND2_X1 U14957 ( .A1(n12797), .A2(n8531), .ZN(n12798) );
  AND2_X1 U14958 ( .A1(n12799), .A2(n12798), .ZN(n12853) );
  MUX2_X1 U14959 ( .A(n15280), .B(n12853), .S(n15254), .Z(n12800) );
  OAI21_X1 U14960 ( .B1(n12855), .B2(n12829), .A(n12800), .ZN(P3_U3479) );
  AOI21_X1 U14961 ( .B1(n12802), .B2(n8531), .A(n12801), .ZN(n12856) );
  MUX2_X1 U14962 ( .A(n12803), .B(n12856), .S(n15254), .Z(n12804) );
  OAI21_X1 U14963 ( .B1(n12829), .B2(n12859), .A(n12804), .ZN(P3_U3478) );
  INV_X1 U14964 ( .A(n12805), .ZN(n12806) );
  AOI21_X1 U14965 ( .B1(n12807), .B2(n8531), .A(n12806), .ZN(n12860) );
  MUX2_X1 U14966 ( .A(n12808), .B(n12860), .S(n15254), .Z(n12809) );
  OAI21_X1 U14967 ( .B1(n12863), .B2(n12829), .A(n12809), .ZN(P3_U3477) );
  NAND2_X1 U14968 ( .A1(n12810), .A2(n8531), .ZN(n12811) );
  NAND2_X1 U14969 ( .A1(n12812), .A2(n12811), .ZN(n12864) );
  MUX2_X1 U14970 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n12864), .S(n15254), .Z(
        n12813) );
  AOI21_X1 U14971 ( .B1(n12823), .B2(n12866), .A(n12813), .ZN(n12814) );
  INV_X1 U14972 ( .A(n12814), .ZN(P3_U3476) );
  AOI21_X1 U14973 ( .B1(n12816), .B2(n8531), .A(n12815), .ZN(n12868) );
  MUX2_X1 U14974 ( .A(n12817), .B(n12868), .S(n15254), .Z(n12818) );
  OAI21_X1 U14975 ( .B1(n7672), .B2(n12829), .A(n12818), .ZN(P3_U3475) );
  NAND2_X1 U14976 ( .A1(n12819), .A2(n8531), .ZN(n12820) );
  NAND2_X1 U14977 ( .A1(n12821), .A2(n12820), .ZN(n12871) );
  MUX2_X1 U14978 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n12871), .S(n15254), .Z(
        n12822) );
  AOI21_X1 U14979 ( .B1(n12823), .B2(n12873), .A(n12822), .ZN(n12824) );
  INV_X1 U14980 ( .A(n12824), .ZN(P3_U3474) );
  AOI21_X1 U14981 ( .B1(n8531), .B2(n12826), .A(n12825), .ZN(n12876) );
  MUX2_X1 U14982 ( .A(n12827), .B(n12876), .S(n15254), .Z(n12828) );
  OAI21_X1 U14983 ( .B1(n12829), .B2(n12879), .A(n12828), .ZN(P3_U3473) );
  INV_X1 U14984 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12831) );
  INV_X1 U14985 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12834) );
  MUX2_X1 U14986 ( .A(n12834), .B(n12833), .S(n15246), .Z(n12835) );
  OAI21_X1 U14987 ( .B1(n12836), .B2(n12880), .A(n12835), .ZN(P3_U3453) );
  MUX2_X1 U14988 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n12837), .S(n15246), .Z(
        P3_U3452) );
  INV_X1 U14989 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12839) );
  MUX2_X1 U14990 ( .A(n12839), .B(n12838), .S(n15246), .Z(n12840) );
  OAI21_X1 U14991 ( .B1(n12841), .B2(n12880), .A(n12840), .ZN(P3_U3451) );
  INV_X1 U14992 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12843) );
  MUX2_X1 U14993 ( .A(n12843), .B(n12842), .S(n15246), .Z(n12844) );
  OAI21_X1 U14994 ( .B1(n12845), .B2(n12880), .A(n12844), .ZN(P3_U3450) );
  INV_X1 U14995 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12847) );
  MUX2_X1 U14996 ( .A(n12847), .B(n12846), .S(n15246), .Z(n12848) );
  OAI21_X1 U14997 ( .B1(n12849), .B2(n12880), .A(n12848), .ZN(P3_U3449) );
  INV_X1 U14998 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12851) );
  MUX2_X1 U14999 ( .A(n12851), .B(n12850), .S(n15246), .Z(n12852) );
  OAI21_X1 U15000 ( .B1(n8512), .B2(n12880), .A(n12852), .ZN(P3_U3448) );
  INV_X1 U15001 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n15399) );
  MUX2_X1 U15002 ( .A(n15399), .B(n12853), .S(n15246), .Z(n12854) );
  OAI21_X1 U15003 ( .B1(n12855), .B2(n12880), .A(n12854), .ZN(P3_U3447) );
  INV_X1 U15004 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12857) );
  MUX2_X1 U15005 ( .A(n12857), .B(n12856), .S(n15246), .Z(n12858) );
  OAI21_X1 U15006 ( .B1(n12880), .B2(n12859), .A(n12858), .ZN(P3_U3446) );
  INV_X1 U15007 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12861) );
  MUX2_X1 U15008 ( .A(n12861), .B(n12860), .S(n15246), .Z(n12862) );
  OAI21_X1 U15009 ( .B1(n12863), .B2(n12880), .A(n12862), .ZN(P3_U3444) );
  INV_X1 U15010 ( .A(n12880), .ZN(n12874) );
  MUX2_X1 U15011 ( .A(n12864), .B(P3_REG0_REG_17__SCAN_IN), .S(n15244), .Z(
        n12865) );
  AOI21_X1 U15012 ( .B1(n12874), .B2(n12866), .A(n12865), .ZN(n12867) );
  INV_X1 U15013 ( .A(n12867), .ZN(P3_U3441) );
  INV_X1 U15014 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12869) );
  MUX2_X1 U15015 ( .A(n12869), .B(n12868), .S(n15246), .Z(n12870) );
  OAI21_X1 U15016 ( .B1(n7672), .B2(n12880), .A(n12870), .ZN(P3_U3438) );
  MUX2_X1 U15017 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n12871), .S(n15246), .Z(
        n12872) );
  AOI21_X1 U15018 ( .B1(n12874), .B2(n12873), .A(n12872), .ZN(n12875) );
  INV_X1 U15019 ( .A(n12875), .ZN(P3_U3435) );
  INV_X1 U15020 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12877) );
  MUX2_X1 U15021 ( .A(n12877), .B(n12876), .S(n15246), .Z(n12878) );
  OAI21_X1 U15022 ( .B1(n12880), .B2(n12879), .A(n12878), .ZN(P3_U3432) );
  MUX2_X1 U15023 ( .A(n12882), .B(P3_D_REG_1__SCAN_IN), .S(n12881), .Z(
        P3_U3377) );
  MUX2_X1 U15024 ( .A(P3_D_REG_0__SCAN_IN), .B(n12884), .S(n12883), .Z(
        P3_U3376) );
  NAND4_X1 U15025 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_STATE_REG_SCAN_IN), 
        .A3(n7786), .A4(n7784), .ZN(n12887) );
  OAI22_X1 U15026 ( .A1(n12885), .A2(n12887), .B1(n12886), .B2(n12900), .ZN(
        n12888) );
  AOI21_X1 U15027 ( .B1(n12890), .B2(n12889), .A(n12888), .ZN(n12891) );
  INV_X1 U15028 ( .A(n12891), .ZN(P3_U3264) );
  INV_X1 U15029 ( .A(n12892), .ZN(n12894) );
  OAI222_X1 U15030 ( .A1(P3_U3151), .A2(n12895), .B1(n12903), .B2(n12894), 
        .C1(n12893), .C2(n12900), .ZN(P3_U3266) );
  INV_X1 U15031 ( .A(n12896), .ZN(n12898) );
  OAI222_X1 U15032 ( .A1(n7017), .A2(P3_U3151), .B1(n12903), .B2(n12898), .C1(
        n12897), .C2(n12900), .ZN(P3_U3269) );
  INV_X1 U15033 ( .A(n12899), .ZN(n12902) );
  OAI222_X1 U15034 ( .A1(n12904), .A2(P3_U3151), .B1(n12903), .B2(n12902), 
        .C1(n12901), .C2(n12900), .ZN(P3_U3270) );
  MUX2_X1 U15035 ( .A(n12905), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  XNOR2_X1 U15036 ( .A(n13375), .B(n12968), .ZN(n12917) );
  NAND2_X1 U15037 ( .A1(n13247), .A2(n10457), .ZN(n12918) );
  XNOR2_X1 U15038 ( .A(n13387), .B(n12937), .ZN(n12916) );
  NAND2_X1 U15039 ( .A1(n13245), .A2(n10457), .ZN(n12915) );
  NOR2_X1 U15040 ( .A1(n13218), .A2(n11062), .ZN(n12960) );
  XNOR2_X1 U15041 ( .A(n13533), .B(n12937), .ZN(n12909) );
  NAND2_X1 U15042 ( .A1(n13236), .A2(n10457), .ZN(n12908) );
  NAND2_X1 U15043 ( .A1(n12909), .A2(n12908), .ZN(n12910) );
  OAI21_X1 U15044 ( .B1(n12909), .B2(n12908), .A(n12910), .ZN(n12999) );
  INV_X1 U15045 ( .A(n12910), .ZN(n12911) );
  XNOR2_X1 U15046 ( .A(n13424), .B(n12968), .ZN(n12913) );
  NAND2_X1 U15047 ( .A1(n13239), .A2(n10457), .ZN(n12912) );
  XNOR2_X1 U15048 ( .A(n12913), .B(n12912), .ZN(n13035) );
  INV_X1 U15049 ( .A(n12912), .ZN(n12914) );
  XNOR2_X1 U15050 ( .A(n12916), .B(n12915), .ZN(n13016) );
  XNOR2_X1 U15051 ( .A(n13518), .B(n12968), .ZN(n12959) );
  NAND2_X1 U15052 ( .A1(n12959), .A2(n12960), .ZN(n12958) );
  XNOR2_X1 U15053 ( .A(n12917), .B(n12918), .ZN(n12980) );
  INV_X1 U15054 ( .A(n12919), .ZN(n12920) );
  XNOR2_X1 U15055 ( .A(n13494), .B(n12968), .ZN(n12924) );
  XNOR2_X1 U15056 ( .A(n12923), .B(n12924), .ZN(n12949) );
  NOR2_X1 U15057 ( .A1(n12921), .A2(n11062), .ZN(n12922) );
  INV_X1 U15058 ( .A(n12923), .ZN(n12925) );
  NAND2_X1 U15059 ( .A1(n12948), .A2(n6561), .ZN(n13005) );
  XNOR2_X1 U15060 ( .A(n13488), .B(n12937), .ZN(n12988) );
  NAND2_X1 U15061 ( .A1(n13074), .A2(n10457), .ZN(n12926) );
  NOR2_X1 U15062 ( .A1(n12988), .A2(n12926), .ZN(n12931) );
  AOI21_X1 U15063 ( .B1(n12988), .B2(n12926), .A(n12931), .ZN(n13006) );
  XNOR2_X1 U15064 ( .A(n13482), .B(n12968), .ZN(n13043) );
  AND2_X1 U15065 ( .A1(n13252), .A2(n10457), .ZN(n12927) );
  NAND2_X1 U15066 ( .A1(n13043), .A2(n12927), .ZN(n12932) );
  INV_X1 U15067 ( .A(n13043), .ZN(n12929) );
  INV_X1 U15068 ( .A(n12927), .ZN(n12928) );
  NAND2_X1 U15069 ( .A1(n12929), .A2(n12928), .ZN(n12930) );
  AND2_X1 U15070 ( .A1(n12932), .A2(n12930), .ZN(n12986) );
  XNOR2_X1 U15071 ( .A(n13476), .B(n12968), .ZN(n12933) );
  NAND2_X1 U15072 ( .A1(n13256), .A2(n10457), .ZN(n12934) );
  XNOR2_X1 U15073 ( .A(n12933), .B(n12934), .ZN(n13046) );
  INV_X1 U15074 ( .A(n12933), .ZN(n12935) );
  NAND2_X1 U15075 ( .A1(n12935), .A2(n12934), .ZN(n12936) );
  XNOR2_X1 U15076 ( .A(n13469), .B(n12937), .ZN(n12939) );
  NAND2_X1 U15077 ( .A1(n13227), .A2(n10457), .ZN(n12938) );
  NOR2_X1 U15078 ( .A1(n12939), .A2(n12938), .ZN(n12966) );
  AOI21_X1 U15079 ( .B1(n12939), .B2(n12938), .A(n12966), .ZN(n12940) );
  OAI211_X1 U15080 ( .C1(n12941), .C2(n12940), .A(n12967), .B(n14912), .ZN(
        n12947) );
  NAND2_X1 U15081 ( .A1(n13229), .A2(n13198), .ZN(n12943) );
  NAND2_X1 U15082 ( .A1(n13256), .A2(n13049), .ZN(n12942) );
  NAND2_X1 U15083 ( .A1(n12943), .A2(n12942), .ZN(n13468) );
  INV_X1 U15084 ( .A(n13468), .ZN(n13292) );
  OAI22_X1 U15085 ( .A1(n13038), .A2(n13292), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12944), .ZN(n12945) );
  AOI21_X1 U15086 ( .B1(n13290), .B2(n13007), .A(n12945), .ZN(n12946) );
  INV_X1 U15087 ( .A(n12948), .ZN(n12957) );
  AOI22_X1 U15088 ( .A1(n12949), .A2(n14912), .B1(n13068), .B2(n13226), .ZN(
        n12956) );
  NAND2_X1 U15089 ( .A1(n13248), .A2(n13049), .ZN(n12951) );
  NAND2_X1 U15090 ( .A1(n13074), .A2(n13198), .ZN(n12950) );
  NAND2_X1 U15091 ( .A1(n12951), .A2(n12950), .ZN(n13343) );
  AOI22_X1 U15092 ( .A1(n13343), .A2(n14914), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12952) );
  OAI21_X1 U15093 ( .B1(n12953), .B2(n14551), .A(n12952), .ZN(n12954) );
  AOI21_X1 U15094 ( .B1(n13225), .B2(n14916), .A(n12954), .ZN(n12955) );
  OAI21_X1 U15095 ( .B1(n12957), .B2(n12956), .A(n12955), .ZN(P2_U3188) );
  OAI21_X1 U15096 ( .B1(n12960), .B2(n12959), .A(n12958), .ZN(n12961) );
  XNOR2_X1 U15097 ( .A(n13013), .B(n12961), .ZN(n12965) );
  INV_X1 U15098 ( .A(n13239), .ZN(n13215) );
  OAI22_X1 U15099 ( .A1(n13221), .A2(n14539), .B1(n13215), .B2(n14541), .ZN(
        n13396) );
  NAND2_X1 U15100 ( .A1(n13396), .A2(n14914), .ZN(n12962) );
  NAND2_X1 U15101 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13193)
         );
  OAI211_X1 U15102 ( .C1(n14551), .C2(n13401), .A(n12962), .B(n13193), .ZN(
        n12963) );
  AOI21_X1 U15103 ( .B1(n13518), .B2(n14916), .A(n12963), .ZN(n12964) );
  OAI21_X1 U15104 ( .B1(n12965), .B2(n14903), .A(n12964), .ZN(P2_U3191) );
  NAND2_X1 U15105 ( .A1(n13229), .A2(n10457), .ZN(n12969) );
  XNOR2_X1 U15106 ( .A(n12969), .B(n12968), .ZN(n12970) );
  XNOR2_X1 U15107 ( .A(n13282), .B(n12970), .ZN(n12971) );
  XNOR2_X1 U15108 ( .A(n12972), .B(n12971), .ZN(n12978) );
  INV_X1 U15109 ( .A(n12973), .ZN(n13279) );
  OAI22_X1 U15110 ( .A1(n12974), .A2(n14539), .B1(n13258), .B2(n14541), .ZN(
        n13276) );
  AOI22_X1 U15111 ( .A1(n14914), .A2(n13276), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12975) );
  OAI21_X1 U15112 ( .B1(n13279), .B2(n14551), .A(n12975), .ZN(n12976) );
  AOI21_X1 U15113 ( .B1(n13282), .B2(n14916), .A(n12976), .ZN(n12977) );
  OAI21_X1 U15114 ( .B1(n12978), .B2(n14903), .A(n12977), .ZN(P2_U3192) );
  OAI211_X1 U15115 ( .C1(n12981), .C2(n12980), .A(n12979), .B(n14912), .ZN(
        n12985) );
  AOI22_X1 U15116 ( .A1(n13248), .A2(n13198), .B1(n13245), .B2(n13049), .ZN(
        n13368) );
  INV_X1 U15117 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12982) );
  OAI22_X1 U15118 ( .A1(n13368), .A2(n13038), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12982), .ZN(n12983) );
  AOI21_X1 U15119 ( .B1(n13374), .B2(n13007), .A(n12983), .ZN(n12984) );
  OAI211_X1 U15120 ( .C1(n6818), .C2(n12998), .A(n12985), .B(n12984), .ZN(
        P2_U3195) );
  INV_X1 U15121 ( .A(n12986), .ZN(n12987) );
  AOI21_X1 U15122 ( .B1(n6530), .B2(n12987), .A(n14903), .ZN(n12990) );
  NOR3_X1 U15123 ( .A1(n12988), .A2(n13251), .A3(n13012), .ZN(n12989) );
  OAI21_X1 U15124 ( .B1(n12990), .B2(n12989), .A(n13045), .ZN(n12997) );
  NAND2_X1 U15125 ( .A1(n13074), .A2(n13049), .ZN(n12992) );
  NAND2_X1 U15126 ( .A1(n13256), .A2(n13198), .ZN(n12991) );
  NAND2_X1 U15127 ( .A1(n12992), .A2(n12991), .ZN(n13481) );
  INV_X1 U15128 ( .A(n13481), .ZN(n12994) );
  OAI22_X1 U15129 ( .A1(n13038), .A2(n12994), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12993), .ZN(n12995) );
  AOI21_X1 U15130 ( .B1(n13314), .B2(n13007), .A(n12995), .ZN(n12996) );
  OAI211_X1 U15131 ( .C1(n13317), .C2(n12998), .A(n12997), .B(n12996), .ZN(
        P2_U3197) );
  AOI21_X1 U15132 ( .B1(n13000), .B2(n12999), .A(n6645), .ZN(n13004) );
  NOR2_X1 U15133 ( .A1(n14551), .A2(n13441), .ZN(n13002) );
  AOI22_X1 U15134 ( .A1(n13239), .A2(n13198), .B1(n13049), .B2(n13233), .ZN(
        n13434) );
  NAND2_X1 U15135 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n15029)
         );
  OAI21_X1 U15136 ( .B1(n13038), .B2(n13434), .A(n15029), .ZN(n13001) );
  AOI211_X1 U15137 ( .C1(n13533), .C2(n14916), .A(n13002), .B(n13001), .ZN(
        n13003) );
  OAI21_X1 U15138 ( .B1(n13004), .B2(n14903), .A(n13003), .ZN(P2_U3200) );
  OAI211_X1 U15139 ( .C1(n13006), .C2(n13005), .A(n6530), .B(n14912), .ZN(
        n13011) );
  OAI22_X1 U15140 ( .A1(n12921), .A2(n14541), .B1(n13254), .B2(n14539), .ZN(
        n13325) );
  AOI22_X1 U15141 ( .A1(n14914), .A2(n13325), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13010) );
  NAND2_X1 U15142 ( .A1(n13488), .A2(n14916), .ZN(n13009) );
  NAND2_X1 U15143 ( .A1(n13007), .A2(n13332), .ZN(n13008) );
  NAND4_X1 U15144 ( .A1(n13011), .A2(n13010), .A3(n13009), .A4(n13008), .ZN(
        P2_U3201) );
  NOR3_X1 U15145 ( .A1(n13013), .A2(n13218), .A3(n13012), .ZN(n13014) );
  AOI21_X1 U15146 ( .B1(n14912), .B2(n13015), .A(n13014), .ZN(n13025) );
  INV_X1 U15147 ( .A(n13016), .ZN(n13024) );
  NAND2_X1 U15148 ( .A1(n13017), .A2(n14912), .ZN(n13023) );
  INV_X1 U15149 ( .A(n13018), .ZN(n13388) );
  NOR2_X1 U15150 ( .A1(n14551), .A2(n13388), .ZN(n13021) );
  AOI22_X1 U15151 ( .A1(n13247), .A2(n13198), .B1(n13049), .B2(n13075), .ZN(
        n13510) );
  OAI22_X1 U15152 ( .A1(n13510), .A2(n13038), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13019), .ZN(n13020) );
  AOI211_X1 U15153 ( .C1(n13387), .C2(n14916), .A(n13021), .B(n13020), .ZN(
        n13022) );
  OAI211_X1 U15154 ( .C1(n13025), .C2(n13024), .A(n13023), .B(n13022), .ZN(
        P2_U3205) );
  AOI22_X1 U15155 ( .A1(n13026), .A2(n14912), .B1(n13068), .B2(n13248), .ZN(
        n13034) );
  INV_X1 U15156 ( .A(n13027), .ZN(n13033) );
  NAND2_X1 U15157 ( .A1(n13247), .A2(n13049), .ZN(n13029) );
  NAND2_X1 U15158 ( .A1(n13226), .A2(n13198), .ZN(n13028) );
  NAND2_X1 U15159 ( .A1(n13029), .A2(n13028), .ZN(n13351) );
  AOI22_X1 U15160 ( .A1(n13351), .A2(n14914), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13030) );
  OAI21_X1 U15161 ( .B1(n13358), .B2(n14551), .A(n13030), .ZN(n13031) );
  AOI21_X1 U15162 ( .B1(n13501), .B2(n14916), .A(n13031), .ZN(n13032) );
  OAI21_X1 U15163 ( .B1(n13034), .B2(n13033), .A(n13032), .ZN(P2_U3207) );
  XNOR2_X1 U15164 ( .A(n13036), .B(n13035), .ZN(n13042) );
  NOR2_X1 U15165 ( .A1(n14551), .A2(n13419), .ZN(n13040) );
  AND2_X1 U15166 ( .A1(n13236), .A2(n13049), .ZN(n13037) );
  AOI21_X1 U15167 ( .B1(n13075), .B2(n13198), .A(n13037), .ZN(n13417) );
  NAND2_X1 U15168 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n15044)
         );
  OAI21_X1 U15169 ( .B1(n13417), .B2(n13038), .A(n15044), .ZN(n13039) );
  AOI211_X1 U15170 ( .C1(n13424), .C2(n14916), .A(n13040), .B(n13039), .ZN(
        n13041) );
  OAI21_X1 U15171 ( .B1(n13042), .B2(n14903), .A(n13041), .ZN(P2_U3210) );
  NAND3_X1 U15172 ( .A1(n13043), .A2(n13068), .A3(n13252), .ZN(n13044) );
  OAI21_X1 U15173 ( .B1(n13045), .B2(n14903), .A(n13044), .ZN(n13048) );
  INV_X1 U15174 ( .A(n13046), .ZN(n13047) );
  NAND2_X1 U15175 ( .A1(n13048), .A2(n13047), .ZN(n13056) );
  INV_X1 U15176 ( .A(n13303), .ZN(n13053) );
  NAND2_X1 U15177 ( .A1(n13252), .A2(n13049), .ZN(n13051) );
  NAND2_X1 U15178 ( .A1(n13227), .A2(n13198), .ZN(n13050) );
  NAND2_X1 U15179 ( .A1(n13051), .A2(n13050), .ZN(n13475) );
  AOI22_X1 U15180 ( .A1(n14914), .A2(n13475), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13052) );
  OAI21_X1 U15181 ( .B1(n13053), .B2(n14551), .A(n13052), .ZN(n13054) );
  AOI21_X1 U15182 ( .B1(n13476), .B2(n14916), .A(n13054), .ZN(n13055) );
  OAI211_X1 U15183 ( .C1(n14903), .C2(n13057), .A(n13056), .B(n13055), .ZN(
        P2_U3212) );
  INV_X1 U15184 ( .A(n13058), .ZN(n13060) );
  AOI22_X1 U15185 ( .A1(n14914), .A2(n13545), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13059) );
  OAI21_X1 U15186 ( .B1(n13060), .B2(n14551), .A(n13059), .ZN(n13067) );
  INV_X1 U15187 ( .A(n13061), .ZN(n13062) );
  OR2_X1 U15188 ( .A1(n14543), .A2(n13062), .ZN(n13064) );
  XNOR2_X1 U15189 ( .A(n13064), .B(n13063), .ZN(n13069) );
  NOR3_X1 U15190 ( .A1(n13069), .A2(n13065), .A3(n14903), .ZN(n13066) );
  AOI211_X1 U15191 ( .C1(n13546), .C2(n14916), .A(n13067), .B(n13066), .ZN(
        n13071) );
  NAND3_X1 U15192 ( .A1(n13069), .A2(n13068), .A3(n13076), .ZN(n13070) );
  NAND2_X1 U15193 ( .A1(n13071), .A2(n13070), .ZN(P2_U3213) );
  MUX2_X1 U15194 ( .A(n13200), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13083), .Z(
        P2_U3562) );
  MUX2_X1 U15195 ( .A(n13072), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13083), .Z(
        P2_U3561) );
  MUX2_X1 U15196 ( .A(n13073), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13083), .Z(
        P2_U3560) );
  MUX2_X1 U15197 ( .A(n13229), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13083), .Z(
        P2_U3559) );
  MUX2_X1 U15198 ( .A(n13227), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13083), .Z(
        P2_U3558) );
  MUX2_X1 U15199 ( .A(n13256), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13083), .Z(
        P2_U3557) );
  MUX2_X1 U15200 ( .A(n13252), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13083), .Z(
        P2_U3556) );
  MUX2_X1 U15201 ( .A(n13074), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13083), .Z(
        P2_U3555) );
  MUX2_X1 U15202 ( .A(n13226), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13083), .Z(
        P2_U3554) );
  MUX2_X1 U15203 ( .A(n13248), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13083), .Z(
        P2_U3553) );
  MUX2_X1 U15204 ( .A(n13247), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13083), .Z(
        P2_U3552) );
  MUX2_X1 U15205 ( .A(n13245), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13083), .Z(
        P2_U3551) );
  INV_X1 U15206 ( .A(P2_U3947), .ZN(n13089) );
  MUX2_X1 U15207 ( .A(n13075), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13089), .Z(
        P2_U3550) );
  MUX2_X1 U15208 ( .A(n13239), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13083), .Z(
        P2_U3549) );
  MUX2_X1 U15209 ( .A(n13236), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13083), .Z(
        P2_U3548) );
  MUX2_X1 U15210 ( .A(n13233), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13089), .Z(
        P2_U3547) );
  MUX2_X1 U15211 ( .A(n13076), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13083), .Z(
        P2_U3546) );
  MUX2_X1 U15212 ( .A(n13077), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13083), .Z(
        P2_U3545) );
  MUX2_X1 U15213 ( .A(n13078), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13089), .Z(
        P2_U3544) );
  MUX2_X1 U15214 ( .A(n13079), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13083), .Z(
        P2_U3543) );
  MUX2_X1 U15215 ( .A(n13080), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13083), .Z(
        P2_U3542) );
  MUX2_X1 U15216 ( .A(n13081), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13089), .Z(
        P2_U3541) );
  MUX2_X1 U15217 ( .A(n13082), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13083), .Z(
        P2_U3540) );
  MUX2_X1 U15218 ( .A(n13084), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13083), .Z(
        P2_U3539) );
  MUX2_X1 U15219 ( .A(n13085), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13089), .Z(
        P2_U3538) );
  MUX2_X1 U15220 ( .A(n13086), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13089), .Z(
        P2_U3537) );
  MUX2_X1 U15221 ( .A(n13087), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13089), .Z(
        P2_U3536) );
  MUX2_X1 U15222 ( .A(n13088), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13089), .Z(
        P2_U3535) );
  MUX2_X1 U15223 ( .A(n9780), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13089), .Z(
        P2_U3534) );
  MUX2_X1 U15224 ( .A(n9784), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13089), .Z(
        P2_U3533) );
  MUX2_X1 U15225 ( .A(n9833), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13089), .Z(
        P2_U3532) );
  MUX2_X1 U15226 ( .A(n9782), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13089), .Z(
        P2_U3531) );
  INV_X1 U15227 ( .A(n15037), .ZN(n15028) );
  INV_X1 U15228 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n13091) );
  OAI22_X1 U15229 ( .A1(n15046), .A2(n13091), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13090), .ZN(n13092) );
  AOI21_X1 U15230 ( .B1(n13093), .B2(n15028), .A(n13092), .ZN(n13102) );
  OAI211_X1 U15231 ( .C1(n13096), .C2(n13095), .A(n15043), .B(n13094), .ZN(
        n13101) );
  OAI211_X1 U15232 ( .C1(n13099), .C2(n13098), .A(n15035), .B(n13097), .ZN(
        n13100) );
  NAND3_X1 U15233 ( .A1(n13102), .A2(n13101), .A3(n13100), .ZN(P2_U3215) );
  INV_X1 U15234 ( .A(n13103), .ZN(n13107) );
  INV_X1 U15235 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n13105) );
  NAND2_X1 U15236 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n13104) );
  OAI21_X1 U15237 ( .B1(n15046), .B2(n13105), .A(n13104), .ZN(n13106) );
  AOI21_X1 U15238 ( .B1(n13107), .B2(n15028), .A(n13106), .ZN(n13116) );
  OAI211_X1 U15239 ( .C1(n13110), .C2(n13109), .A(n15035), .B(n13108), .ZN(
        n13115) );
  OAI211_X1 U15240 ( .C1(n13113), .C2(n13112), .A(n15043), .B(n13111), .ZN(
        n13114) );
  NAND3_X1 U15241 ( .A1(n13116), .A2(n13115), .A3(n13114), .ZN(P2_U3217) );
  INV_X1 U15242 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14399) );
  NAND2_X1 U15243 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n13117) );
  OAI21_X1 U15244 ( .B1(n15046), .B2(n14399), .A(n13117), .ZN(n13118) );
  AOI21_X1 U15245 ( .B1(n13119), .B2(n15028), .A(n13118), .ZN(n13128) );
  OAI211_X1 U15246 ( .C1(n13122), .C2(n13121), .A(n15035), .B(n13120), .ZN(
        n13127) );
  OAI211_X1 U15247 ( .C1(n13125), .C2(n13124), .A(n15043), .B(n13123), .ZN(
        n13126) );
  NAND3_X1 U15248 ( .A1(n13128), .A2(n13127), .A3(n13126), .ZN(P2_U3218) );
  INV_X1 U15249 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n13130) );
  NAND2_X1 U15250 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n13129) );
  OAI21_X1 U15251 ( .B1(n15046), .B2(n13130), .A(n13129), .ZN(n13131) );
  AOI21_X1 U15252 ( .B1(n13132), .B2(n15028), .A(n13131), .ZN(n13141) );
  OAI211_X1 U15253 ( .C1(n13135), .C2(n13134), .A(n15035), .B(n13133), .ZN(
        n13140) );
  OAI211_X1 U15254 ( .C1(n13138), .C2(n13137), .A(n15043), .B(n13136), .ZN(
        n13139) );
  NAND3_X1 U15255 ( .A1(n13141), .A2(n13140), .A3(n13139), .ZN(P2_U3219) );
  NAND2_X1 U15256 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n13142) );
  OAI21_X1 U15257 ( .B1(n15046), .B2(n7515), .A(n13142), .ZN(n13143) );
  AOI21_X1 U15258 ( .B1(n13144), .B2(n15028), .A(n13143), .ZN(n13153) );
  OAI211_X1 U15259 ( .C1(n13147), .C2(n13146), .A(n15035), .B(n13145), .ZN(
        n13152) );
  OAI211_X1 U15260 ( .C1(n13150), .C2(n13149), .A(n15043), .B(n13148), .ZN(
        n13151) );
  NAND3_X1 U15261 ( .A1(n13153), .A2(n13152), .A3(n13151), .ZN(P2_U3220) );
  OAI21_X1 U15262 ( .B1(n15046), .B2(n7066), .A(n13154), .ZN(n13155) );
  AOI21_X1 U15263 ( .B1(n13156), .B2(n15028), .A(n13155), .ZN(n13165) );
  OAI211_X1 U15264 ( .C1(n13159), .C2(n13158), .A(n15043), .B(n13157), .ZN(
        n13164) );
  OAI211_X1 U15265 ( .C1(n13162), .C2(n13161), .A(n15035), .B(n13160), .ZN(
        n13163) );
  NAND3_X1 U15266 ( .A1(n13165), .A2(n13164), .A3(n13163), .ZN(P2_U3221) );
  NOR2_X1 U15267 ( .A1(n13167), .A2(n13166), .ZN(n13168) );
  NOR2_X1 U15268 ( .A1(n13168), .A2(n13181), .ZN(n13169) );
  INV_X1 U15269 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n14992) );
  XNOR2_X1 U15270 ( .A(n13181), .B(n13168), .ZN(n14993) );
  NOR2_X1 U15271 ( .A1(n14992), .A2(n14993), .ZN(n14991) );
  NOR2_X1 U15272 ( .A1(n13169), .A2(n14991), .ZN(n15010) );
  INV_X1 U15273 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13170) );
  XNOR2_X1 U15274 ( .A(n13171), .B(n13170), .ZN(n15009) );
  NAND2_X1 U15275 ( .A1(n15013), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n13172) );
  NAND2_X1 U15276 ( .A1(n15006), .A2(n13172), .ZN(n15019) );
  OR2_X1 U15277 ( .A1(n15027), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13173) );
  NAND2_X1 U15278 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n15027), .ZN(n13174) );
  AND2_X1 U15279 ( .A1(n13173), .A2(n13174), .ZN(n15018) );
  NAND2_X1 U15280 ( .A1(n15019), .A2(n15018), .ZN(n15017) );
  NAND2_X1 U15281 ( .A1(n15017), .A2(n13174), .ZN(n13176) );
  XOR2_X1 U15282 ( .A(n13175), .B(n13176), .Z(n15033) );
  INV_X1 U15283 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n15034) );
  NAND2_X1 U15284 ( .A1(n15033), .A2(n15034), .ZN(n15032) );
  OR2_X1 U15285 ( .A1(n13176), .A2(n13175), .ZN(n13177) );
  NAND2_X1 U15286 ( .A1(n15032), .A2(n13177), .ZN(n13178) );
  XNOR2_X1 U15287 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13178), .ZN(n13190) );
  INV_X1 U15288 ( .A(n13190), .ZN(n13188) );
  AOI21_X1 U15289 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n13180), .A(n13179), 
        .ZN(n13182) );
  NOR2_X1 U15290 ( .A1(n13182), .A2(n13181), .ZN(n13183) );
  INV_X1 U15291 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14995) );
  XNOR2_X1 U15292 ( .A(n13182), .B(n13181), .ZN(n14996) );
  NOR2_X1 U15293 ( .A1(n14995), .A2(n14996), .ZN(n14994) );
  NOR2_X1 U15294 ( .A1(n13183), .A2(n14994), .ZN(n15005) );
  XNOR2_X1 U15295 ( .A(n15013), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n15004) );
  NOR2_X1 U15296 ( .A1(n15005), .A2(n15004), .ZN(n15003) );
  AOI21_X1 U15297 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n15013), .A(n15003), 
        .ZN(n15024) );
  XNOR2_X1 U15298 ( .A(n15027), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15023) );
  NOR2_X1 U15299 ( .A1(n15024), .A2(n15023), .ZN(n15021) );
  AOI21_X1 U15300 ( .B1(n15027), .B2(P2_REG1_REG_17__SCAN_IN), .A(n15021), 
        .ZN(n13184) );
  NOR2_X1 U15301 ( .A1(n13184), .A2(n15038), .ZN(n13185) );
  AOI21_X1 U15302 ( .B1(n13184), .B2(n15038), .A(n13185), .ZN(n15036) );
  AND2_X1 U15303 ( .A1(n15036), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n15039) );
  NOR2_X1 U15304 ( .A1(n15039), .A2(n13185), .ZN(n13186) );
  XNOR2_X1 U15305 ( .A(n13186), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13189) );
  OAI21_X1 U15306 ( .B1(n13189), .B2(n15022), .A(n15037), .ZN(n13187) );
  AOI21_X1 U15307 ( .B1(n13188), .B2(n15043), .A(n13187), .ZN(n13192) );
  AOI22_X1 U15308 ( .A1(n13190), .A2(n15043), .B1(n15035), .B2(n13189), .ZN(
        n13191) );
  MUX2_X1 U15309 ( .A(n13192), .B(n13191), .S(n9247), .Z(n13194) );
  OAI211_X1 U15310 ( .C1(n6795), .C2(n15046), .A(n13194), .B(n13193), .ZN(
        P2_U3233) );
  INV_X1 U15311 ( .A(n13454), .ZN(n13267) );
  INV_X1 U15312 ( .A(n13533), .ZN(n13436) );
  INV_X1 U15313 ( .A(n13424), .ZN(n13525) );
  INV_X1 U15314 ( .A(n13518), .ZN(n13404) );
  NAND2_X1 U15315 ( .A1(n13195), .A2(n14562), .ZN(n13449) );
  NAND2_X1 U15316 ( .A1(n13196), .A2(P2_B_REG_SCAN_IN), .ZN(n13197) );
  NAND2_X1 U15317 ( .A1(n13198), .A2(n13197), .ZN(n13232) );
  INV_X1 U15318 ( .A(n13232), .ZN(n13199) );
  NAND2_X1 U15319 ( .A1(n13200), .A2(n13199), .ZN(n13451) );
  NOR2_X1 U15320 ( .A1(n15076), .A2(n13451), .ZN(n13208) );
  INV_X1 U15321 ( .A(n13201), .ZN(n13450) );
  NOR2_X1 U15322 ( .A1(n13450), .A2(n15055), .ZN(n13202) );
  AOI211_X1 U15323 ( .C1(n15076), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13208), 
        .B(n13202), .ZN(n13203) );
  OAI21_X1 U15324 ( .B1(n13449), .B2(n13444), .A(n13203), .ZN(P2_U3234) );
  INV_X1 U15325 ( .A(n13263), .ZN(n13206) );
  NOR2_X1 U15326 ( .A1(n13453), .A2(n15055), .ZN(n13207) );
  AOI211_X1 U15327 ( .C1(n15076), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13208), 
        .B(n13207), .ZN(n13209) );
  OAI21_X1 U15328 ( .B1(n13444), .B2(n13452), .A(n13209), .ZN(P2_U3235) );
  INV_X1 U15329 ( .A(n13282), .ZN(n13458) );
  AND2_X1 U15330 ( .A1(n13538), .A2(n13210), .ZN(n13211) );
  INV_X1 U15331 ( .A(n13429), .ZN(n13432) );
  NAND2_X1 U15332 ( .A1(n13424), .A2(n13215), .ZN(n13214) );
  OR2_X1 U15333 ( .A1(n13424), .A2(n13215), .ZN(n13216) );
  NAND2_X1 U15334 ( .A1(n13518), .A2(n13218), .ZN(n13219) );
  AND2_X1 U15335 ( .A1(n13387), .A2(n13221), .ZN(n13222) );
  OAI21_X1 U15336 ( .B1(n6818), .B2(n13247), .A(n13366), .ZN(n13223) );
  INV_X1 U15337 ( .A(n13501), .ZN(n13362) );
  INV_X1 U15338 ( .A(n13328), .ZN(n13323) );
  INV_X1 U15339 ( .A(n13298), .ZN(n13300) );
  INV_X1 U15340 ( .A(n13229), .ZN(n13230) );
  INV_X1 U15341 ( .A(n13476), .ZN(n13306) );
  INV_X1 U15342 ( .A(n13488), .ZN(n13335) );
  NAND2_X1 U15343 ( .A1(n13538), .A2(n13233), .ZN(n13234) );
  AND2_X1 U15344 ( .A1(n13533), .A2(n13236), .ZN(n13237) );
  NAND2_X1 U15345 ( .A1(n13410), .A2(n13413), .ZN(n13412) );
  OR2_X1 U15346 ( .A1(n13424), .A2(n13239), .ZN(n13240) );
  NAND2_X1 U15347 ( .A1(n13406), .A2(n13241), .ZN(n13243) );
  NOR2_X1 U15348 ( .A1(n13387), .A2(n13245), .ZN(n13244) );
  NAND2_X1 U15349 ( .A1(n13387), .A2(n13245), .ZN(n13246) );
  NAND2_X1 U15350 ( .A1(n13311), .A2(n13253), .ZN(n13255) );
  NAND2_X1 U15351 ( .A1(n13255), .A2(n7754), .ZN(n13301) );
  INV_X1 U15352 ( .A(n13277), .ZN(n13261) );
  AOI21_X1 U15353 ( .B1(n13454), .B2(n13261), .A(n13459), .ZN(n13262) );
  AND2_X1 U15354 ( .A1(n13263), .A2(n13262), .ZN(n13456) );
  NAND2_X1 U15355 ( .A1(n13456), .A2(n15049), .ZN(n13266) );
  AOI22_X1 U15356 ( .A1(n15076), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n13264), 
        .B2(n15051), .ZN(n13265) );
  OAI211_X1 U15357 ( .C1(n13267), .C2(n15055), .A(n13266), .B(n13265), .ZN(
        n13268) );
  AOI21_X1 U15358 ( .B1(n13269), .B2(n15059), .A(n13268), .ZN(n13270) );
  OAI21_X1 U15359 ( .B1(n13271), .B2(n15076), .A(n13270), .ZN(P2_U3236) );
  OAI21_X1 U15360 ( .B1(n13273), .B2(n13275), .A(n13272), .ZN(n13464) );
  INV_X1 U15361 ( .A(n13463), .ZN(n13281) );
  AND2_X1 U15362 ( .A1(n13282), .A2(n13288), .ZN(n13278) );
  OR2_X1 U15363 ( .A1(n13278), .A2(n13277), .ZN(n13460) );
  OAI22_X1 U15364 ( .A1(n13460), .A2(n10457), .B1(n13279), .B2(n15070), .ZN(
        n13280) );
  OAI21_X1 U15365 ( .B1(n13281), .B2(n13280), .A(n13446), .ZN(n13284) );
  AOI22_X1 U15366 ( .A1(n13282), .A2(n14556), .B1(n15076), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n13283) );
  OAI211_X1 U15367 ( .C1(n13448), .C2(n13464), .A(n13284), .B(n13283), .ZN(
        P2_U3237) );
  XOR2_X1 U15368 ( .A(n13286), .B(n13285), .Z(n13472) );
  OR2_X1 U15369 ( .A1(n13287), .A2(n13286), .ZN(n13466) );
  NAND3_X1 U15370 ( .A1(n13466), .A2(n13465), .A3(n15059), .ZN(n13297) );
  AOI21_X1 U15371 ( .B1(n13469), .B2(n13302), .A(n13459), .ZN(n13289) );
  AND2_X1 U15372 ( .A1(n13289), .A2(n13288), .ZN(n13467) );
  INV_X1 U15373 ( .A(n13290), .ZN(n13291) );
  OAI22_X1 U15374 ( .A1(n15076), .A2(n13292), .B1(n13291), .B2(n15070), .ZN(
        n13293) );
  AOI21_X1 U15375 ( .B1(P2_REG2_REG_27__SCAN_IN), .B2(n15076), .A(n13293), 
        .ZN(n13294) );
  OAI21_X1 U15376 ( .B1(n7185), .B2(n15055), .A(n13294), .ZN(n13295) );
  AOI21_X1 U15377 ( .B1(n15049), .B2(n13467), .A(n13295), .ZN(n13296) );
  OAI211_X1 U15378 ( .C1(n13472), .C2(n13310), .A(n13297), .B(n13296), .ZN(
        P2_U3238) );
  XNOR2_X1 U15379 ( .A(n13299), .B(n13298), .ZN(n13479) );
  XNOR2_X1 U15380 ( .A(n13301), .B(n13300), .ZN(n13473) );
  NAND2_X1 U15381 ( .A1(n13473), .A2(n15059), .ZN(n13309) );
  AOI211_X1 U15382 ( .C1(n13476), .C2(n13312), .A(n13459), .B(n7186), .ZN(
        n13474) );
  AOI22_X1 U15383 ( .A1(n13446), .A2(n13475), .B1(n13303), .B2(n15051), .ZN(
        n13305) );
  NAND2_X1 U15384 ( .A1(n15076), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n13304) );
  OAI211_X1 U15385 ( .C1(n13306), .C2(n15055), .A(n13305), .B(n13304), .ZN(
        n13307) );
  AOI21_X1 U15386 ( .B1(n13474), .B2(n15049), .A(n13307), .ZN(n13308) );
  OAI211_X1 U15387 ( .C1(n13479), .C2(n13310), .A(n13309), .B(n13308), .ZN(
        P2_U3239) );
  XNOR2_X1 U15388 ( .A(n13311), .B(n13319), .ZN(n13486) );
  INV_X1 U15389 ( .A(n13312), .ZN(n13313) );
  AOI211_X1 U15390 ( .C1(n13482), .C2(n13330), .A(n13459), .B(n13313), .ZN(
        n13480) );
  AOI22_X1 U15391 ( .A1(n13446), .A2(n13481), .B1(n13314), .B2(n15051), .ZN(
        n13316) );
  NAND2_X1 U15392 ( .A1(n15076), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n13315) );
  OAI211_X1 U15393 ( .C1(n13317), .C2(n15055), .A(n13316), .B(n13315), .ZN(
        n13318) );
  AOI21_X1 U15394 ( .B1(n13480), .B2(n15049), .A(n13318), .ZN(n13322) );
  XNOR2_X1 U15395 ( .A(n13320), .B(n13319), .ZN(n13483) );
  NAND2_X1 U15396 ( .A1(n13483), .A2(n13384), .ZN(n13321) );
  OAI211_X1 U15397 ( .C1(n13486), .C2(n13448), .A(n13322), .B(n13321), .ZN(
        P2_U3240) );
  XNOR2_X1 U15398 ( .A(n13324), .B(n13323), .ZN(n13326) );
  AOI21_X1 U15399 ( .B1(n13326), .B2(n14579), .A(n13325), .ZN(n13490) );
  OAI21_X1 U15400 ( .B1(n13329), .B2(n13328), .A(n13327), .ZN(n13491) );
  INV_X1 U15401 ( .A(n13491), .ZN(n13337) );
  AOI21_X1 U15402 ( .B1(n13488), .B2(n13342), .A(n13459), .ZN(n13331) );
  AND2_X1 U15403 ( .A1(n13331), .A2(n13330), .ZN(n13487) );
  NAND2_X1 U15404 ( .A1(n13487), .A2(n15049), .ZN(n13334) );
  AOI22_X1 U15405 ( .A1(n15076), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n13332), 
        .B2(n15051), .ZN(n13333) );
  OAI211_X1 U15406 ( .C1(n13335), .C2(n15055), .A(n13334), .B(n13333), .ZN(
        n13336) );
  AOI21_X1 U15407 ( .B1(n13337), .B2(n15059), .A(n13336), .ZN(n13338) );
  OAI21_X1 U15408 ( .B1(n15076), .B2(n13490), .A(n13338), .ZN(P2_U3241) );
  XNOR2_X1 U15409 ( .A(n13339), .B(n13340), .ZN(n13498) );
  XNOR2_X1 U15410 ( .A(n13341), .B(n13340), .ZN(n13496) );
  OAI211_X1 U15411 ( .C1(n13357), .C2(n13494), .A(n14562), .B(n13342), .ZN(
        n13493) );
  INV_X1 U15412 ( .A(n13343), .ZN(n13492) );
  OAI21_X1 U15413 ( .B1(n13493), .B2(n9550), .A(n13492), .ZN(n13344) );
  NAND2_X1 U15414 ( .A1(n13344), .A2(n13446), .ZN(n13347) );
  AOI22_X1 U15415 ( .A1(n15076), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n13345), 
        .B2(n15051), .ZN(n13346) );
  OAI211_X1 U15416 ( .C1(n13494), .C2(n15055), .A(n13347), .B(n13346), .ZN(
        n13348) );
  AOI21_X1 U15417 ( .B1(n13496), .B2(n13384), .A(n13348), .ZN(n13349) );
  OAI21_X1 U15418 ( .B1(n13498), .B2(n13448), .A(n13349), .ZN(P2_U3242) );
  XOR2_X1 U15419 ( .A(n13350), .B(n13354), .Z(n13352) );
  AOI21_X1 U15420 ( .B1(n13352), .B2(n14579), .A(n13351), .ZN(n13503) );
  AOI21_X1 U15421 ( .B1(n13354), .B2(n13353), .A(n6543), .ZN(n13499) );
  NAND2_X1 U15422 ( .A1(n13373), .A2(n13501), .ZN(n13355) );
  NAND2_X1 U15423 ( .A1(n13355), .A2(n14562), .ZN(n13356) );
  NOR2_X1 U15424 ( .A1(n13357), .A2(n13356), .ZN(n13500) );
  NAND2_X1 U15425 ( .A1(n13500), .A2(n15049), .ZN(n13361) );
  INV_X1 U15426 ( .A(n13358), .ZN(n13359) );
  AOI22_X1 U15427 ( .A1(P2_REG2_REG_22__SCAN_IN), .A2(n15076), .B1(n13359), 
        .B2(n15051), .ZN(n13360) );
  OAI211_X1 U15428 ( .C1(n13362), .C2(n15055), .A(n13361), .B(n13360), .ZN(
        n13363) );
  AOI21_X1 U15429 ( .B1(n13499), .B2(n15059), .A(n13363), .ZN(n13364) );
  OAI21_X1 U15430 ( .B1(n13503), .B2(n15076), .A(n13364), .ZN(P2_U3243) );
  INV_X1 U15431 ( .A(n13370), .ZN(n13365) );
  XNOR2_X1 U15432 ( .A(n13366), .B(n13365), .ZN(n13367) );
  NAND2_X1 U15433 ( .A1(n13367), .A2(n14579), .ZN(n13369) );
  NAND2_X1 U15434 ( .A1(n13369), .A2(n13368), .ZN(n13509) );
  INV_X1 U15435 ( .A(n13509), .ZN(n13380) );
  XNOR2_X1 U15436 ( .A(n13371), .B(n13370), .ZN(n13505) );
  NAND2_X1 U15437 ( .A1(n13375), .A2(n13385), .ZN(n13372) );
  NAND3_X1 U15438 ( .A1(n13373), .A2(n14562), .A3(n13372), .ZN(n13506) );
  AOI22_X1 U15439 ( .A1(n15076), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13374), 
        .B2(n15051), .ZN(n13377) );
  NAND2_X1 U15440 ( .A1(n13375), .A2(n14556), .ZN(n13376) );
  OAI211_X1 U15441 ( .C1(n13506), .C2(n13444), .A(n13377), .B(n13376), .ZN(
        n13378) );
  AOI21_X1 U15442 ( .B1(n13505), .B2(n15059), .A(n13378), .ZN(n13379) );
  OAI21_X1 U15443 ( .B1(n13380), .B2(n15076), .A(n13379), .ZN(P2_U3244) );
  XNOR2_X1 U15444 ( .A(n13381), .B(n13382), .ZN(n13516) );
  XNOR2_X1 U15445 ( .A(n13383), .B(n13382), .ZN(n13514) );
  NAND2_X1 U15446 ( .A1(n13514), .A2(n13384), .ZN(n13394) );
  AOI21_X1 U15447 ( .B1(n13387), .B2(n13398), .A(n13459), .ZN(n13386) );
  NAND2_X1 U15448 ( .A1(n13386), .A2(n13385), .ZN(n13511) );
  INV_X1 U15449 ( .A(n13511), .ZN(n13392) );
  INV_X1 U15450 ( .A(n13387), .ZN(n13512) );
  OAI22_X1 U15451 ( .A1(n13510), .A2(n15076), .B1(n13388), .B2(n15070), .ZN(
        n13389) );
  AOI21_X1 U15452 ( .B1(P2_REG2_REG_20__SCAN_IN), .B2(n15076), .A(n13389), 
        .ZN(n13390) );
  OAI21_X1 U15453 ( .B1(n13512), .B2(n15055), .A(n13390), .ZN(n13391) );
  AOI21_X1 U15454 ( .B1(n13392), .B2(n15049), .A(n13391), .ZN(n13393) );
  OAI211_X1 U15455 ( .C1(n13448), .C2(n13516), .A(n13394), .B(n13393), .ZN(
        P2_U3245) );
  XOR2_X1 U15456 ( .A(n13395), .B(n13405), .Z(n13397) );
  AOI21_X1 U15457 ( .B1(n13397), .B2(n14579), .A(n13396), .ZN(n13520) );
  INV_X1 U15458 ( .A(n13421), .ZN(n13400) );
  INV_X1 U15459 ( .A(n13398), .ZN(n13399) );
  AOI211_X1 U15460 ( .C1(n13518), .C2(n13400), .A(n13459), .B(n13399), .ZN(
        n13517) );
  INV_X1 U15461 ( .A(n13401), .ZN(n13402) );
  AOI22_X1 U15462 ( .A1(n15076), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13402), 
        .B2(n15051), .ZN(n13403) );
  OAI21_X1 U15463 ( .B1(n13404), .B2(n15055), .A(n13403), .ZN(n13408) );
  XNOR2_X1 U15464 ( .A(n13406), .B(n13405), .ZN(n13521) );
  NOR2_X1 U15465 ( .A1(n13521), .A2(n13448), .ZN(n13407) );
  AOI211_X1 U15466 ( .C1(n13517), .C2(n15049), .A(n13408), .B(n13407), .ZN(
        n13409) );
  OAI21_X1 U15467 ( .B1(n15076), .B2(n13520), .A(n13409), .ZN(P2_U3246) );
  OR2_X1 U15468 ( .A1(n13410), .A2(n13413), .ZN(n13411) );
  NAND2_X1 U15469 ( .A1(n13412), .A2(n13411), .ZN(n13522) );
  INV_X1 U15470 ( .A(n13522), .ZN(n13428) );
  XNOR2_X1 U15471 ( .A(n13414), .B(n13413), .ZN(n13415) );
  NAND2_X1 U15472 ( .A1(n13415), .A2(n14579), .ZN(n13418) );
  NAND2_X1 U15473 ( .A1(n13522), .A2(n15131), .ZN(n13416) );
  NAND3_X1 U15474 ( .A1(n13418), .A2(n13417), .A3(n13416), .ZN(n13527) );
  NAND2_X1 U15475 ( .A1(n13527), .A2(n13446), .ZN(n13426) );
  OAI22_X1 U15476 ( .A1(n13446), .A2(n15034), .B1(n13419), .B2(n15070), .ZN(
        n13423) );
  OAI21_X1 U15477 ( .B1(n13438), .B2(n13525), .A(n14562), .ZN(n13420) );
  OR2_X1 U15478 ( .A1(n13421), .A2(n13420), .ZN(n13523) );
  NOR2_X1 U15479 ( .A1(n13523), .A2(n13444), .ZN(n13422) );
  AOI211_X1 U15480 ( .C1(n14556), .C2(n13424), .A(n13423), .B(n13422), .ZN(
        n13425) );
  OAI211_X1 U15481 ( .C1(n13428), .C2(n13427), .A(n13426), .B(n13425), .ZN(
        P2_U3247) );
  XNOR2_X1 U15482 ( .A(n13430), .B(n13429), .ZN(n13535) );
  OAI211_X1 U15483 ( .C1(n13433), .C2(n13432), .A(n13431), .B(n14579), .ZN(
        n13435) );
  NAND2_X1 U15484 ( .A1(n13435), .A2(n13434), .ZN(n13531) );
  OAI21_X1 U15485 ( .B1(n13437), .B2(n13436), .A(n14562), .ZN(n13439) );
  OR2_X1 U15486 ( .A1(n13439), .A2(n13438), .ZN(n13530) );
  NAND2_X1 U15487 ( .A1(n15076), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13440) );
  OAI21_X1 U15488 ( .B1(n15070), .B2(n13441), .A(n13440), .ZN(n13442) );
  AOI21_X1 U15489 ( .B1(n13533), .B2(n14556), .A(n13442), .ZN(n13443) );
  OAI21_X1 U15490 ( .B1(n13530), .B2(n13444), .A(n13443), .ZN(n13445) );
  AOI21_X1 U15491 ( .B1(n13531), .B2(n13446), .A(n13445), .ZN(n13447) );
  OAI21_X1 U15492 ( .B1(n13448), .B2(n13535), .A(n13447), .ZN(P2_U3248) );
  OAI211_X1 U15493 ( .C1(n13450), .C2(n15114), .A(n13449), .B(n13451), .ZN(
        n13550) );
  MUX2_X1 U15494 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13550), .S(n15145), .Z(
        P2_U3530) );
  MUX2_X1 U15495 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13551), .S(n15145), .Z(
        P2_U3529) );
  OAI22_X1 U15496 ( .A1(n13460), .A2(n13459), .B1(n13458), .B2(n15114), .ZN(
        n13461) );
  INV_X1 U15497 ( .A(n13461), .ZN(n13462) );
  OAI211_X1 U15498 ( .C1(n14576), .C2(n13464), .A(n13463), .B(n13462), .ZN(
        n13553) );
  MUX2_X1 U15499 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13553), .S(n15145), .Z(
        P2_U3527) );
  NAND3_X1 U15500 ( .A1(n13466), .A2(n13465), .A3(n14570), .ZN(n13471) );
  AOI211_X1 U15501 ( .C1(n15123), .C2(n13469), .A(n13468), .B(n13467), .ZN(
        n13470) );
  OAI211_X1 U15502 ( .C1(n15127), .C2(n13472), .A(n13471), .B(n13470), .ZN(
        n13554) );
  MUX2_X1 U15503 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13554), .S(n15145), .Z(
        P2_U3526) );
  NAND2_X1 U15504 ( .A1(n13473), .A2(n14570), .ZN(n13478) );
  AOI211_X1 U15505 ( .C1(n15123), .C2(n13476), .A(n13475), .B(n13474), .ZN(
        n13477) );
  OAI211_X1 U15506 ( .C1(n15127), .C2(n13479), .A(n13478), .B(n13477), .ZN(
        n13555) );
  MUX2_X1 U15507 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13555), .S(n15145), .Z(
        P2_U3525) );
  AOI211_X1 U15508 ( .C1(n15123), .C2(n13482), .A(n13481), .B(n13480), .ZN(
        n13485) );
  NAND2_X1 U15509 ( .A1(n13483), .A2(n14579), .ZN(n13484) );
  OAI211_X1 U15510 ( .C1(n13486), .C2(n14576), .A(n13485), .B(n13484), .ZN(
        n13556) );
  MUX2_X1 U15511 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13556), .S(n15145), .Z(
        P2_U3524) );
  AOI21_X1 U15512 ( .B1(n15123), .B2(n13488), .A(n13487), .ZN(n13489) );
  OAI211_X1 U15513 ( .C1(n13491), .C2(n14576), .A(n13490), .B(n13489), .ZN(
        n13557) );
  MUX2_X1 U15514 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13557), .S(n15145), .Z(
        P2_U3523) );
  OAI211_X1 U15515 ( .C1(n13494), .C2(n15114), .A(n13493), .B(n13492), .ZN(
        n13495) );
  AOI21_X1 U15516 ( .B1(n13496), .B2(n14579), .A(n13495), .ZN(n13497) );
  OAI21_X1 U15517 ( .B1(n13498), .B2(n14576), .A(n13497), .ZN(n13558) );
  MUX2_X1 U15518 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13558), .S(n15145), .Z(
        P2_U3522) );
  INV_X1 U15519 ( .A(n13499), .ZN(n13504) );
  AOI21_X1 U15520 ( .B1(n15123), .B2(n13501), .A(n13500), .ZN(n13502) );
  OAI211_X1 U15521 ( .C1(n13504), .C2(n14576), .A(n13503), .B(n13502), .ZN(
        n13559) );
  MUX2_X1 U15522 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13559), .S(n15145), .Z(
        P2_U3521) );
  NAND2_X1 U15523 ( .A1(n13505), .A2(n14570), .ZN(n13507) );
  OAI211_X1 U15524 ( .C1(n6818), .C2(n15114), .A(n13507), .B(n13506), .ZN(
        n13508) );
  MUX2_X1 U15525 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13560), .S(n15145), .Z(
        P2_U3520) );
  OAI211_X1 U15526 ( .C1(n13512), .C2(n15114), .A(n13511), .B(n13510), .ZN(
        n13513) );
  AOI21_X1 U15527 ( .B1(n13514), .B2(n14579), .A(n13513), .ZN(n13515) );
  OAI21_X1 U15528 ( .B1(n14576), .B2(n13516), .A(n13515), .ZN(n13561) );
  MUX2_X1 U15529 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13561), .S(n15145), .Z(
        P2_U3519) );
  AOI21_X1 U15530 ( .B1(n15123), .B2(n13518), .A(n13517), .ZN(n13519) );
  OAI211_X1 U15531 ( .C1(n14576), .C2(n13521), .A(n13520), .B(n13519), .ZN(
        n13562) );
  MUX2_X1 U15532 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13562), .S(n15145), .Z(
        P2_U3518) );
  INV_X1 U15533 ( .A(n15107), .ZN(n15124) );
  NAND2_X1 U15534 ( .A1(n13522), .A2(n15124), .ZN(n13524) );
  OAI211_X1 U15535 ( .C1(n13525), .C2(n15114), .A(n13524), .B(n13523), .ZN(
        n13526) );
  NOR2_X1 U15536 ( .A1(n13527), .A2(n13526), .ZN(n13563) );
  MUX2_X1 U15537 ( .A(n13528), .B(n13563), .S(n15145), .Z(n13529) );
  INV_X1 U15538 ( .A(n13529), .ZN(P2_U3517) );
  INV_X1 U15539 ( .A(n13530), .ZN(n13532) );
  AOI211_X1 U15540 ( .C1(n15123), .C2(n13533), .A(n13532), .B(n13531), .ZN(
        n13534) );
  OAI21_X1 U15541 ( .B1(n14576), .B2(n13535), .A(n13534), .ZN(n13566) );
  MUX2_X1 U15542 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13566), .S(n15145), .Z(
        P2_U3516) );
  AOI211_X1 U15543 ( .C1(n15123), .C2(n13538), .A(n13537), .B(n13536), .ZN(
        n13541) );
  NAND2_X1 U15544 ( .A1(n13539), .A2(n14579), .ZN(n13540) );
  OAI211_X1 U15545 ( .C1(n13542), .C2(n14576), .A(n13541), .B(n13540), .ZN(
        n13567) );
  MUX2_X1 U15546 ( .A(n13567), .B(P2_REG1_REG_16__SCAN_IN), .S(n15142), .Z(
        P2_U3515) );
  NAND2_X1 U15547 ( .A1(n13543), .A2(n14579), .ZN(n13548) );
  AOI211_X1 U15548 ( .C1(n15123), .C2(n13546), .A(n13545), .B(n13544), .ZN(
        n13547) );
  OAI211_X1 U15549 ( .C1(n14576), .C2(n13549), .A(n13548), .B(n13547), .ZN(
        n13568) );
  MUX2_X1 U15550 ( .A(n13568), .B(P2_REG1_REG_15__SCAN_IN), .S(n15142), .Z(
        P2_U3514) );
  MUX2_X1 U15551 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13550), .S(n15134), .Z(
        P2_U3498) );
  MUX2_X1 U15552 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13551), .S(n15134), .Z(
        P2_U3497) );
  MUX2_X1 U15553 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13553), .S(n15134), .Z(
        P2_U3495) );
  MUX2_X1 U15554 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13554), .S(n15134), .Z(
        P2_U3494) );
  MUX2_X1 U15555 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13555), .S(n15134), .Z(
        P2_U3493) );
  MUX2_X1 U15556 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13556), .S(n15134), .Z(
        P2_U3492) );
  MUX2_X1 U15557 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13557), .S(n15134), .Z(
        P2_U3491) );
  MUX2_X1 U15558 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13558), .S(n15134), .Z(
        P2_U3490) );
  MUX2_X1 U15559 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13559), .S(n15134), .Z(
        P2_U3489) );
  MUX2_X1 U15560 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13560), .S(n15134), .Z(
        P2_U3488) );
  MUX2_X1 U15561 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13561), .S(n15134), .Z(
        P2_U3487) );
  MUX2_X1 U15562 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13562), .S(n15134), .Z(
        P2_U3486) );
  INV_X1 U15563 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n13564) );
  MUX2_X1 U15564 ( .A(n13564), .B(n13563), .S(n15134), .Z(n13565) );
  INV_X1 U15565 ( .A(n13565), .ZN(P2_U3484) );
  MUX2_X1 U15566 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13566), .S(n15134), .Z(
        P2_U3481) );
  MUX2_X1 U15567 ( .A(n13567), .B(P2_REG0_REG_16__SCAN_IN), .S(n15132), .Z(
        P2_U3478) );
  MUX2_X1 U15568 ( .A(n13568), .B(P2_REG0_REG_15__SCAN_IN), .S(n15132), .Z(
        P2_U3475) );
  INV_X1 U15569 ( .A(n14323), .ZN(n13572) );
  NOR4_X1 U15570 ( .A1(n13569), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3088), 
        .A4(n9208), .ZN(n13570) );
  AOI21_X1 U15571 ( .B1(n13580), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13570), 
        .ZN(n13571) );
  OAI21_X1 U15572 ( .B1(n13572), .B2(n13597), .A(n13571), .ZN(P2_U3296) );
  INV_X1 U15573 ( .A(n13573), .ZN(n14326) );
  OAI222_X1 U15574 ( .A1(n13597), .A2(n14326), .B1(n9240), .B2(P2_U3088), .C1(
        n13574), .C2(n13599), .ZN(P2_U3297) );
  INV_X1 U15575 ( .A(n13575), .ZN(n14329) );
  OAI222_X1 U15576 ( .A1(n13597), .A2(n14329), .B1(n13577), .B2(P2_U3088), 
        .C1(n13576), .C2(n13599), .ZN(P2_U3298) );
  INV_X1 U15577 ( .A(n13578), .ZN(n14332) );
  AOI21_X1 U15578 ( .B1(n13580), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13579), 
        .ZN(n13581) );
  OAI21_X1 U15579 ( .B1(n14332), .B2(n13597), .A(n13581), .ZN(P2_U3299) );
  INV_X1 U15580 ( .A(n13582), .ZN(n14335) );
  OAI222_X1 U15581 ( .A1(n13597), .A2(n14335), .B1(n13584), .B2(P2_U3088), 
        .C1(n13583), .C2(n13599), .ZN(P2_U3300) );
  INV_X1 U15582 ( .A(n13585), .ZN(n14338) );
  INV_X1 U15583 ( .A(n13586), .ZN(n13588) );
  OAI222_X1 U15584 ( .A1(n13597), .A2(n14338), .B1(P2_U3088), .B2(n13588), 
        .C1(n13587), .C2(n13599), .ZN(P2_U3301) );
  INV_X1 U15585 ( .A(n13590), .ZN(n14341) );
  INV_X1 U15586 ( .A(n13591), .ZN(n13592) );
  OAI222_X1 U15587 ( .A1(n13599), .A2(n13593), .B1(n13597), .B2(n14341), .C1(
        n13592), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U15588 ( .A(n13594), .ZN(n14345) );
  INV_X1 U15589 ( .A(n13595), .ZN(n13596) );
  OAI222_X1 U15590 ( .A1(n13599), .A2(n13598), .B1(n13597), .B2(n14345), .C1(
        n13596), .C2(P2_U3088), .ZN(P2_U3303) );
  INV_X1 U15591 ( .A(n13600), .ZN(n13601) );
  MUX2_X1 U15592 ( .A(n13601), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NAND2_X1 U15593 ( .A1(n13988), .A2(n10183), .ZN(n13603) );
  NAND2_X1 U15594 ( .A1(n10220), .A2(n13873), .ZN(n13602) );
  NAND2_X1 U15595 ( .A1(n13603), .A2(n13602), .ZN(n13605) );
  XNOR2_X1 U15596 ( .A(n13605), .B(n13604), .ZN(n13754) );
  AOI22_X1 U15597 ( .A1(n13988), .A2(n10220), .B1(n13759), .B2(n13873), .ZN(
        n13755) );
  XNOR2_X1 U15598 ( .A(n13754), .B(n13755), .ZN(n13757) );
  NOR2_X1 U15599 ( .A1(n13615), .A2(n13606), .ZN(n13607) );
  AOI21_X1 U15600 ( .B1(n13837), .B2(n7054), .A(n13607), .ZN(n13631) );
  INV_X1 U15601 ( .A(n13631), .ZN(n13634) );
  AOI22_X1 U15602 ( .A1(n13837), .A2(n10183), .B1(n7054), .B2(n13885), .ZN(
        n13608) );
  XNOR2_X1 U15603 ( .A(n13608), .B(n13604), .ZN(n13632) );
  INV_X1 U15604 ( .A(n13632), .ZN(n13633) );
  NOR2_X1 U15605 ( .A1(n13615), .A2(n13609), .ZN(n13610) );
  AOI21_X1 U15606 ( .B1(n13791), .B2(n7054), .A(n13610), .ZN(n13628) );
  INV_X1 U15607 ( .A(n13628), .ZN(n13630) );
  NAND2_X1 U15608 ( .A1(n13791), .A2(n10183), .ZN(n13612) );
  NAND2_X1 U15609 ( .A1(n7054), .A2(n13886), .ZN(n13611) );
  NAND2_X1 U15610 ( .A1(n13612), .A2(n13611), .ZN(n13613) );
  XNOR2_X1 U15611 ( .A(n13613), .B(n13604), .ZN(n13629) );
  NOR2_X1 U15612 ( .A1(n13615), .A2(n13614), .ZN(n13616) );
  AOI21_X1 U15613 ( .B1(n14630), .B2(n7054), .A(n13616), .ZN(n13620) );
  INV_X1 U15614 ( .A(n13620), .ZN(n13627) );
  NAND2_X1 U15615 ( .A1(n14630), .A2(n10183), .ZN(n13618) );
  NAND2_X1 U15616 ( .A1(n7054), .A2(n13887), .ZN(n13617) );
  NAND2_X1 U15617 ( .A1(n13618), .A2(n13617), .ZN(n13619) );
  XNOR2_X1 U15618 ( .A(n13619), .B(n13604), .ZN(n13626) );
  XNOR2_X1 U15619 ( .A(n13626), .B(n13620), .ZN(n14612) );
  INV_X1 U15620 ( .A(n13621), .ZN(n13624) );
  INV_X1 U15621 ( .A(n13622), .ZN(n13623) );
  NAND2_X1 U15622 ( .A1(n13624), .A2(n13623), .ZN(n14609) );
  XOR2_X1 U15623 ( .A(n13628), .B(n13629), .Z(n13788) );
  XNOR2_X1 U15624 ( .A(n13632), .B(n13631), .ZN(n13833) );
  NAND2_X1 U15625 ( .A1(n14597), .A2(n10183), .ZN(n13636) );
  NAND2_X1 U15626 ( .A1(n7054), .A2(n13884), .ZN(n13635) );
  NAND2_X1 U15627 ( .A1(n13636), .A2(n13635), .ZN(n13637) );
  XNOR2_X1 U15628 ( .A(n13637), .B(n13604), .ZN(n13640) );
  AOI22_X1 U15629 ( .A1(n14597), .A2(n7054), .B1(n13759), .B2(n13884), .ZN(
        n13638) );
  XNOR2_X1 U15630 ( .A(n13640), .B(n13638), .ZN(n14596) );
  INV_X1 U15631 ( .A(n13638), .ZN(n13639) );
  NAND2_X1 U15632 ( .A1(n14622), .A2(n10183), .ZN(n13643) );
  NAND2_X1 U15633 ( .A1(n7054), .A2(n14151), .ZN(n13642) );
  NAND2_X1 U15634 ( .A1(n13643), .A2(n13642), .ZN(n13644) );
  XNOR2_X1 U15635 ( .A(n13644), .B(n13604), .ZN(n13646) );
  AOI22_X1 U15636 ( .A1(n14622), .A2(n7054), .B1(n13759), .B2(n14151), .ZN(
        n14620) );
  INV_X1 U15637 ( .A(n13646), .ZN(n13647) );
  NAND2_X1 U15638 ( .A1(n14604), .A2(n10183), .ZN(n13650) );
  NAND2_X1 U15639 ( .A1(n7054), .A2(n13883), .ZN(n13649) );
  NAND2_X1 U15640 ( .A1(n13650), .A2(n13649), .ZN(n13651) );
  XNOR2_X1 U15641 ( .A(n13651), .B(n13604), .ZN(n13654) );
  AOI22_X1 U15642 ( .A1(n14604), .A2(n7054), .B1(n13759), .B2(n13883), .ZN(
        n13652) );
  XNOR2_X1 U15643 ( .A(n13654), .B(n13652), .ZN(n14602) );
  INV_X1 U15644 ( .A(n13652), .ZN(n13653) );
  NAND2_X1 U15645 ( .A1(n14264), .A2(n10183), .ZN(n13657) );
  NAND2_X1 U15646 ( .A1(n14150), .A2(n7054), .ZN(n13656) );
  NAND2_X1 U15647 ( .A1(n13657), .A2(n13656), .ZN(n13658) );
  XNOR2_X1 U15648 ( .A(n13658), .B(n13604), .ZN(n13659) );
  AOI22_X1 U15649 ( .A1(n14264), .A2(n7054), .B1(n13759), .B2(n14150), .ZN(
        n13660) );
  XNOR2_X1 U15650 ( .A(n13659), .B(n13660), .ZN(n13803) );
  INV_X1 U15651 ( .A(n13659), .ZN(n13661) );
  NAND2_X1 U15652 ( .A1(n13661), .A2(n13660), .ZN(n13662) );
  NAND2_X1 U15653 ( .A1(n14257), .A2(n10183), .ZN(n13664) );
  NAND2_X1 U15654 ( .A1(n13882), .A2(n7054), .ZN(n13663) );
  NAND2_X1 U15655 ( .A1(n13664), .A2(n13663), .ZN(n13665) );
  XNOR2_X1 U15656 ( .A(n13665), .B(n13604), .ZN(n13668) );
  AOI22_X1 U15657 ( .A1(n14257), .A2(n7054), .B1(n13759), .B2(n13882), .ZN(
        n13666) );
  XNOR2_X1 U15658 ( .A(n13668), .B(n13666), .ZN(n13853) );
  INV_X1 U15659 ( .A(n13666), .ZN(n13667) );
  AOI22_X1 U15660 ( .A1(n14251), .A2(n7054), .B1(n13759), .B2(n13881), .ZN(
        n13671) );
  AOI22_X1 U15661 ( .A1(n14251), .A2(n10183), .B1(n7054), .B2(n13881), .ZN(
        n13669) );
  XNOR2_X1 U15662 ( .A(n13669), .B(n13604), .ZN(n13670) );
  XOR2_X1 U15663 ( .A(n13671), .B(n13670), .Z(n13747) );
  INV_X1 U15664 ( .A(n13670), .ZN(n13673) );
  INV_X1 U15665 ( .A(n13671), .ZN(n13672) );
  AND2_X1 U15666 ( .A1(n13880), .A2(n13759), .ZN(n13674) );
  AOI21_X1 U15667 ( .B1(n14240), .B2(n10220), .A(n13674), .ZN(n13677) );
  AOI22_X1 U15668 ( .A1(n14240), .A2(n10183), .B1(n10220), .B2(n13880), .ZN(
        n13675) );
  XNOR2_X1 U15669 ( .A(n13675), .B(n13604), .ZN(n13676) );
  XOR2_X1 U15670 ( .A(n13677), .B(n13676), .Z(n13822) );
  INV_X1 U15671 ( .A(n13676), .ZN(n13679) );
  INV_X1 U15672 ( .A(n13677), .ZN(n13678) );
  NAND2_X1 U15673 ( .A1(n13679), .A2(n13678), .ZN(n13680) );
  AOI22_X1 U15674 ( .A1(n14076), .A2(n10183), .B1(n10220), .B2(n13879), .ZN(
        n13681) );
  XNOR2_X1 U15675 ( .A(n13681), .B(n13604), .ZN(n13684) );
  AOI22_X1 U15676 ( .A1(n14076), .A2(n7054), .B1(n13759), .B2(n13879), .ZN(
        n13683) );
  XNOR2_X1 U15677 ( .A(n13684), .B(n13683), .ZN(n13773) );
  NAND2_X1 U15678 ( .A1(n13684), .A2(n13683), .ZN(n13685) );
  OAI22_X1 U15679 ( .A1(n14065), .A2(n13687), .B1(n13774), .B2(n13686), .ZN(
        n13688) );
  XNOR2_X1 U15680 ( .A(n13688), .B(n13604), .ZN(n13689) );
  AOI22_X1 U15681 ( .A1(n14305), .A2(n7054), .B1(n13759), .B2(n13878), .ZN(
        n13690) );
  XNOR2_X1 U15682 ( .A(n13689), .B(n13690), .ZN(n13841) );
  INV_X1 U15683 ( .A(n13689), .ZN(n13691) );
  NAND2_X1 U15684 ( .A1(n13691), .A2(n13690), .ZN(n13692) );
  NAND2_X1 U15685 ( .A1(n14221), .A2(n10183), .ZN(n13694) );
  NAND2_X1 U15686 ( .A1(n10220), .A2(n13877), .ZN(n13693) );
  NAND2_X1 U15687 ( .A1(n13694), .A2(n13693), .ZN(n13695) );
  XNOR2_X1 U15688 ( .A(n13695), .B(n13604), .ZN(n13696) );
  AOI22_X1 U15689 ( .A1(n14221), .A2(n7054), .B1(n13759), .B2(n13877), .ZN(
        n13697) );
  XNOR2_X1 U15690 ( .A(n13696), .B(n13697), .ZN(n13729) );
  INV_X1 U15691 ( .A(n13696), .ZN(n13698) );
  NAND2_X1 U15692 ( .A1(n14211), .A2(n10183), .ZN(n13700) );
  NAND2_X1 U15693 ( .A1(n10220), .A2(n13876), .ZN(n13699) );
  NAND2_X1 U15694 ( .A1(n13700), .A2(n13699), .ZN(n13701) );
  XNOR2_X1 U15695 ( .A(n13701), .B(n13604), .ZN(n13702) );
  AOI22_X1 U15696 ( .A1(n14211), .A2(n7054), .B1(n13759), .B2(n13876), .ZN(
        n13703) );
  XNOR2_X1 U15697 ( .A(n13702), .B(n13703), .ZN(n13813) );
  INV_X1 U15698 ( .A(n13702), .ZN(n13704) );
  NAND2_X1 U15699 ( .A1(n13704), .A2(n13703), .ZN(n13705) );
  NAND2_X1 U15700 ( .A1(n14201), .A2(n10183), .ZN(n13708) );
  NAND2_X1 U15701 ( .A1(n10220), .A2(n13875), .ZN(n13707) );
  NAND2_X1 U15702 ( .A1(n13708), .A2(n13707), .ZN(n13709) );
  XNOR2_X1 U15703 ( .A(n13709), .B(n13604), .ZN(n13710) );
  AOI22_X1 U15704 ( .A1(n14201), .A2(n7054), .B1(n13759), .B2(n13875), .ZN(
        n13711) );
  XNOR2_X1 U15705 ( .A(n13710), .B(n13711), .ZN(n13794) );
  INV_X1 U15706 ( .A(n13710), .ZN(n13712) );
  NAND2_X1 U15707 ( .A1(n13712), .A2(n13711), .ZN(n13713) );
  NAND2_X1 U15708 ( .A1(n13866), .A2(n10183), .ZN(n13715) );
  NAND2_X1 U15709 ( .A1(n10220), .A2(n13874), .ZN(n13714) );
  NAND2_X1 U15710 ( .A1(n13715), .A2(n13714), .ZN(n13717) );
  XNOR2_X1 U15711 ( .A(n13717), .B(n13604), .ZN(n13718) );
  AOI22_X1 U15712 ( .A1(n13866), .A2(n7054), .B1(n13759), .B2(n13874), .ZN(
        n13719) );
  XNOR2_X1 U15713 ( .A(n13718), .B(n13719), .ZN(n13859) );
  INV_X1 U15714 ( .A(n13718), .ZN(n13720) );
  XOR2_X1 U15715 ( .A(n13757), .B(n13758), .Z(n13727) );
  INV_X1 U15716 ( .A(n13991), .ZN(n13724) );
  NAND2_X1 U15717 ( .A1(n13874), .A2(n13861), .ZN(n13722) );
  NAND2_X1 U15718 ( .A1(n13872), .A2(n14149), .ZN(n13721) );
  NAND2_X1 U15719 ( .A1(n13722), .A2(n13721), .ZN(n13979) );
  AOI22_X1 U15720 ( .A1(n14625), .A2(n13979), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13723) );
  OAI21_X1 U15721 ( .B1(n14629), .B2(n13724), .A(n13723), .ZN(n13725) );
  AOI21_X1 U15722 ( .B1(n13988), .B2(n14621), .A(n13725), .ZN(n13726) );
  OAI21_X1 U15723 ( .B1(n13727), .B2(n13868), .A(n13726), .ZN(P1_U3214) );
  XOR2_X1 U15724 ( .A(n13729), .B(n13728), .Z(n13736) );
  INV_X1 U15725 ( .A(n14049), .ZN(n13733) );
  OR2_X1 U15726 ( .A1(n13804), .A2(n13774), .ZN(n13731) );
  NAND2_X1 U15727 ( .A1(n13876), .A2(n14149), .ZN(n13730) );
  NAND2_X1 U15728 ( .A1(n13731), .A2(n13730), .ZN(n14220) );
  AOI22_X1 U15729 ( .A1(n14625), .A2(n14220), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13732) );
  OAI21_X1 U15730 ( .B1(n14629), .B2(n13733), .A(n13732), .ZN(n13734) );
  AOI21_X1 U15731 ( .B1(n14221), .B2(n14621), .A(n13734), .ZN(n13735) );
  OAI21_X1 U15732 ( .B1(n13736), .B2(n13868), .A(n13735), .ZN(P1_U3216) );
  AOI21_X1 U15733 ( .B1(n13738), .B2(n13737), .A(n13868), .ZN(n13740) );
  NAND2_X1 U15734 ( .A1(n13740), .A2(n13739), .ZN(n13745) );
  AOI22_X1 U15735 ( .A1(n14621), .A2(n13742), .B1(n14625), .B2(n13741), .ZN(
        n13744) );
  MUX2_X1 U15736 ( .A(n14629), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n13743) );
  NAND3_X1 U15737 ( .A1(n13745), .A2(n13744), .A3(n13743), .ZN(P1_U3218) );
  INV_X1 U15738 ( .A(n14251), .ZN(n14110) );
  OAI211_X1 U15739 ( .C1(n13748), .C2(n13747), .A(n13746), .B(n14623), .ZN(
        n13753) );
  NAND2_X1 U15740 ( .A1(n13880), .A2(n14149), .ZN(n13750) );
  NAND2_X1 U15741 ( .A1(n13882), .A2(n13861), .ZN(n13749) );
  NAND2_X1 U15742 ( .A1(n13750), .A2(n13749), .ZN(n14250) );
  AND2_X1 U15743 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13932) );
  NOR2_X1 U15744 ( .A1(n14629), .A2(n14105), .ZN(n13751) );
  AOI211_X1 U15745 ( .C1(n14625), .C2(n14250), .A(n13932), .B(n13751), .ZN(
        n13752) );
  OAI211_X1 U15746 ( .C1(n14110), .C2(n13851), .A(n13753), .B(n13752), .ZN(
        P1_U3219) );
  INV_X1 U15747 ( .A(n13754), .ZN(n13756) );
  AOI22_X1 U15748 ( .A1(n14288), .A2(n10220), .B1(n13759), .B2(n13872), .ZN(
        n13762) );
  AOI22_X1 U15749 ( .A1(n14288), .A2(n10183), .B1(n10220), .B2(n13872), .ZN(
        n13760) );
  XNOR2_X1 U15750 ( .A(n13760), .B(n13604), .ZN(n13761) );
  XOR2_X1 U15751 ( .A(n13762), .B(n13761), .Z(n13763) );
  INV_X1 U15752 ( .A(n13764), .ZN(n13966) );
  NAND2_X1 U15753 ( .A1(n13871), .A2(n14149), .ZN(n13766) );
  NAND2_X1 U15754 ( .A1(n13873), .A2(n13861), .ZN(n13765) );
  NAND2_X1 U15755 ( .A1(n13766), .A2(n13765), .ZN(n13965) );
  AOI22_X1 U15756 ( .A1(n14625), .A2(n13965), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13767) );
  OAI21_X1 U15757 ( .B1(n14629), .B2(n13966), .A(n13767), .ZN(n13768) );
  AOI21_X1 U15758 ( .B1(n14288), .B2(n14621), .A(n13768), .ZN(n13769) );
  INV_X1 U15759 ( .A(n13770), .ZN(n13771) );
  AOI21_X1 U15760 ( .B1(n13773), .B2(n13772), .A(n13771), .ZN(n13781) );
  NAND2_X1 U15761 ( .A1(n13880), .A2(n13861), .ZN(n13776) );
  OR2_X1 U15762 ( .A1(n13806), .A2(n13774), .ZN(n13775) );
  AND2_X1 U15763 ( .A1(n13776), .A2(n13775), .ZN(n14232) );
  OAI22_X1 U15764 ( .A1(n13846), .A2(n14232), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13777), .ZN(n13778) );
  AOI21_X1 U15765 ( .B1(n13848), .B2(n14077), .A(n13778), .ZN(n13780) );
  NAND2_X1 U15766 ( .A1(n14076), .A2(n14621), .ZN(n13779) );
  OAI211_X1 U15767 ( .C1(n13781), .C2(n13868), .A(n13780), .B(n13779), .ZN(
        P1_U3223) );
  NAND2_X1 U15768 ( .A1(n13848), .A2(n13782), .ZN(n13784) );
  OAI211_X1 U15769 ( .C1(n13785), .C2(n13846), .A(n13784), .B(n13783), .ZN(
        n13790) );
  AOI211_X1 U15770 ( .C1(n13788), .C2(n13787), .A(n13868), .B(n13786), .ZN(
        n13789) );
  AOI211_X1 U15771 ( .C1(n14621), .C2(n13791), .A(n13790), .B(n13789), .ZN(
        n13792) );
  INV_X1 U15772 ( .A(n13792), .ZN(P1_U3224) );
  XOR2_X1 U15773 ( .A(n13794), .B(n13793), .Z(n13801) );
  INV_X1 U15774 ( .A(n13795), .ZN(n14014) );
  NAND2_X1 U15775 ( .A1(n13876), .A2(n13861), .ZN(n13797) );
  NAND2_X1 U15776 ( .A1(n13874), .A2(n14149), .ZN(n13796) );
  NAND2_X1 U15777 ( .A1(n13797), .A2(n13796), .ZN(n14013) );
  AOI22_X1 U15778 ( .A1(n14625), .A2(n14013), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13798) );
  OAI21_X1 U15779 ( .B1(n14629), .B2(n14014), .A(n13798), .ZN(n13799) );
  AOI21_X1 U15780 ( .B1(n14201), .B2(n14621), .A(n13799), .ZN(n13800) );
  OAI21_X1 U15781 ( .B1(n13801), .B2(n13868), .A(n13800), .ZN(P1_U3225) );
  XOR2_X1 U15782 ( .A(n13803), .B(n13802), .Z(n13811) );
  NAND2_X1 U15783 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14763)
         );
  OAI22_X1 U15784 ( .A1(n13807), .A2(n13806), .B1(n13805), .B2(n13804), .ZN(
        n14263) );
  NAND2_X1 U15785 ( .A1(n14625), .A2(n14263), .ZN(n13808) );
  OAI211_X1 U15786 ( .C1(n14629), .C2(n14136), .A(n14763), .B(n13808), .ZN(
        n13809) );
  AOI21_X1 U15787 ( .B1(n14264), .B2(n14621), .A(n13809), .ZN(n13810) );
  OAI21_X1 U15788 ( .B1(n13811), .B2(n13868), .A(n13810), .ZN(P1_U3228) );
  XOR2_X1 U15789 ( .A(n13813), .B(n13812), .Z(n13820) );
  INV_X1 U15790 ( .A(n14037), .ZN(n13817) );
  NAND2_X1 U15791 ( .A1(n13877), .A2(n13861), .ZN(n13815) );
  NAND2_X1 U15792 ( .A1(n13875), .A2(n14149), .ZN(n13814) );
  NAND2_X1 U15793 ( .A1(n13815), .A2(n13814), .ZN(n14027) );
  AOI22_X1 U15794 ( .A1(n14625), .A2(n14027), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13816) );
  OAI21_X1 U15795 ( .B1(n14629), .B2(n13817), .A(n13816), .ZN(n13818) );
  AOI21_X1 U15796 ( .B1(n14211), .B2(n14621), .A(n13818), .ZN(n13819) );
  OAI21_X1 U15797 ( .B1(n13820), .B2(n13868), .A(n13819), .ZN(P1_U3229) );
  OAI211_X1 U15798 ( .C1(n13823), .C2(n13822), .A(n13821), .B(n14623), .ZN(
        n13829) );
  INV_X1 U15799 ( .A(n13824), .ZN(n14091) );
  AND2_X1 U15800 ( .A1(n13879), .A2(n14149), .ZN(n13825) );
  AOI21_X1 U15801 ( .B1(n13881), .B2(n13861), .A(n13825), .ZN(n14087) );
  OAI22_X1 U15802 ( .A1(n13846), .A2(n14087), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13826), .ZN(n13827) );
  AOI21_X1 U15803 ( .B1(n13848), .B2(n14091), .A(n13827), .ZN(n13828) );
  OAI211_X1 U15804 ( .C1(n6829), .C2(n13851), .A(n13829), .B(n13828), .ZN(
        P1_U3233) );
  NAND2_X1 U15805 ( .A1(n13848), .A2(n13830), .ZN(n13831) );
  NAND2_X1 U15806 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14700)
         );
  OAI211_X1 U15807 ( .C1(n14640), .C2(n13846), .A(n13831), .B(n14700), .ZN(
        n13836) );
  AOI211_X1 U15808 ( .C1(n13834), .C2(n13833), .A(n13868), .B(n13832), .ZN(
        n13835) );
  AOI211_X1 U15809 ( .C1(n14621), .C2(n13837), .A(n13836), .B(n13835), .ZN(
        n13838) );
  INV_X1 U15810 ( .A(n13838), .ZN(P1_U3234) );
  OAI21_X1 U15811 ( .B1(n13841), .B2(n13840), .A(n13839), .ZN(n13842) );
  NAND2_X1 U15812 ( .A1(n13842), .A2(n14623), .ZN(n13850) );
  NAND2_X1 U15813 ( .A1(n13879), .A2(n13861), .ZN(n13844) );
  NAND2_X1 U15814 ( .A1(n13877), .A2(n14149), .ZN(n13843) );
  AND2_X1 U15815 ( .A1(n13844), .A2(n13843), .ZN(n14057) );
  OAI22_X1 U15816 ( .A1(n13846), .A2(n14057), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13845), .ZN(n13847) );
  AOI21_X1 U15817 ( .B1(n13848), .B2(n14063), .A(n13847), .ZN(n13849) );
  OAI211_X1 U15818 ( .C1(n13851), .C2(n14065), .A(n13850), .B(n13849), .ZN(
        P1_U3235) );
  XOR2_X1 U15819 ( .A(n13852), .B(n13853), .Z(n13857) );
  NAND2_X1 U15820 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14779)
         );
  AND2_X1 U15821 ( .A1(n13881), .A2(n14149), .ZN(n14256) );
  AND2_X1 U15822 ( .A1(n14150), .A2(n13861), .ZN(n14118) );
  OAI21_X1 U15823 ( .B1(n14256), .B2(n14118), .A(n14625), .ZN(n13854) );
  OAI211_X1 U15824 ( .C1(n14629), .C2(n14124), .A(n14779), .B(n13854), .ZN(
        n13855) );
  AOI21_X1 U15825 ( .B1(n14257), .B2(n14621), .A(n13855), .ZN(n13856) );
  OAI21_X1 U15826 ( .B1(n13857), .B2(n13868), .A(n13856), .ZN(P1_U3238) );
  XOR2_X1 U15827 ( .A(n13859), .B(n13858), .Z(n13869) );
  INV_X1 U15828 ( .A(n13860), .ZN(n14003) );
  NAND2_X1 U15829 ( .A1(n13875), .A2(n13861), .ZN(n13863) );
  NAND2_X1 U15830 ( .A1(n13873), .A2(n14149), .ZN(n13862) );
  NAND2_X1 U15831 ( .A1(n13863), .A2(n13862), .ZN(n14002) );
  AOI22_X1 U15832 ( .A1(n14625), .A2(n14002), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13864) );
  OAI21_X1 U15833 ( .B1(n14629), .B2(n14003), .A(n13864), .ZN(n13865) );
  AOI21_X1 U15834 ( .B1(n13866), .B2(n14621), .A(n13865), .ZN(n13867) );
  OAI21_X1 U15835 ( .B1(n13869), .B2(n13868), .A(n13867), .ZN(P1_U3240) );
  MUX2_X1 U15836 ( .A(n13870), .B(P1_DATAO_REG_30__SCAN_IN), .S(n13896), .Z(
        P1_U3590) );
  MUX2_X1 U15837 ( .A(n13871), .B(P1_DATAO_REG_29__SCAN_IN), .S(n13896), .Z(
        P1_U3589) );
  MUX2_X1 U15838 ( .A(n13872), .B(P1_DATAO_REG_28__SCAN_IN), .S(n13896), .Z(
        P1_U3588) );
  MUX2_X1 U15839 ( .A(n13873), .B(P1_DATAO_REG_27__SCAN_IN), .S(n13896), .Z(
        P1_U3587) );
  MUX2_X1 U15840 ( .A(n13874), .B(P1_DATAO_REG_26__SCAN_IN), .S(n13896), .Z(
        P1_U3586) );
  MUX2_X1 U15841 ( .A(n13875), .B(P1_DATAO_REG_25__SCAN_IN), .S(n13896), .Z(
        P1_U3585) );
  MUX2_X1 U15842 ( .A(n13876), .B(P1_DATAO_REG_24__SCAN_IN), .S(n13896), .Z(
        P1_U3584) );
  MUX2_X1 U15843 ( .A(n13877), .B(P1_DATAO_REG_23__SCAN_IN), .S(n13896), .Z(
        P1_U3583) );
  MUX2_X1 U15844 ( .A(n13878), .B(P1_DATAO_REG_22__SCAN_IN), .S(n13896), .Z(
        P1_U3582) );
  MUX2_X1 U15845 ( .A(n13879), .B(P1_DATAO_REG_21__SCAN_IN), .S(n13896), .Z(
        P1_U3581) );
  MUX2_X1 U15846 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13880), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15847 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13881), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15848 ( .A(n13882), .B(P1_DATAO_REG_18__SCAN_IN), .S(n13896), .Z(
        P1_U3578) );
  MUX2_X1 U15849 ( .A(n14150), .B(P1_DATAO_REG_17__SCAN_IN), .S(n13896), .Z(
        P1_U3577) );
  MUX2_X1 U15850 ( .A(n13883), .B(P1_DATAO_REG_16__SCAN_IN), .S(n13896), .Z(
        P1_U3576) );
  MUX2_X1 U15851 ( .A(n14151), .B(P1_DATAO_REG_15__SCAN_IN), .S(n13896), .Z(
        P1_U3575) );
  MUX2_X1 U15852 ( .A(n13884), .B(P1_DATAO_REG_14__SCAN_IN), .S(n13896), .Z(
        P1_U3574) );
  MUX2_X1 U15853 ( .A(n13885), .B(P1_DATAO_REG_13__SCAN_IN), .S(n13896), .Z(
        P1_U3573) );
  MUX2_X1 U15854 ( .A(n13886), .B(P1_DATAO_REG_12__SCAN_IN), .S(n13896), .Z(
        P1_U3572) );
  MUX2_X1 U15855 ( .A(n13887), .B(P1_DATAO_REG_11__SCAN_IN), .S(n13896), .Z(
        P1_U3571) );
  MUX2_X1 U15856 ( .A(n13888), .B(P1_DATAO_REG_10__SCAN_IN), .S(n13896), .Z(
        P1_U3570) );
  MUX2_X1 U15857 ( .A(n13889), .B(P1_DATAO_REG_9__SCAN_IN), .S(n13896), .Z(
        P1_U3569) );
  MUX2_X1 U15858 ( .A(n13890), .B(P1_DATAO_REG_8__SCAN_IN), .S(n13896), .Z(
        P1_U3568) );
  MUX2_X1 U15859 ( .A(n13891), .B(P1_DATAO_REG_7__SCAN_IN), .S(n13896), .Z(
        P1_U3567) );
  MUX2_X1 U15860 ( .A(n13892), .B(P1_DATAO_REG_6__SCAN_IN), .S(n13896), .Z(
        P1_U3566) );
  MUX2_X1 U15861 ( .A(n13893), .B(P1_DATAO_REG_5__SCAN_IN), .S(n13896), .Z(
        P1_U3565) );
  MUX2_X1 U15862 ( .A(n7571), .B(P1_DATAO_REG_4__SCAN_IN), .S(n13896), .Z(
        P1_U3564) );
  MUX2_X1 U15863 ( .A(n13894), .B(P1_DATAO_REG_3__SCAN_IN), .S(n13896), .Z(
        P1_U3563) );
  MUX2_X1 U15864 ( .A(n13895), .B(P1_DATAO_REG_2__SCAN_IN), .S(n13896), .Z(
        P1_U3562) );
  MUX2_X1 U15865 ( .A(n13897), .B(P1_DATAO_REG_1__SCAN_IN), .S(n13896), .Z(
        P1_U3561) );
  INV_X1 U15866 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n13898) );
  MUX2_X1 U15867 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n13898), .S(n14699), .Z(
        n13899) );
  INV_X1 U15868 ( .A(n13899), .ZN(n14695) );
  OAI21_X1 U15869 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n13913), .A(n13900), 
        .ZN(n14696) );
  NOR2_X1 U15870 ( .A1(n14695), .A2(n14696), .ZN(n14694) );
  INV_X1 U15871 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n13901) );
  MUX2_X1 U15872 ( .A(n13901), .B(P1_REG2_REG_14__SCAN_IN), .S(n14708), .Z(
        n14704) );
  NAND2_X1 U15873 ( .A1(n13902), .A2(n13917), .ZN(n13904) );
  XNOR2_X1 U15874 ( .A(n13917), .B(n13903), .ZN(n14722) );
  INV_X1 U15875 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n14721) );
  NAND2_X1 U15876 ( .A1(n14722), .A2(n14721), .ZN(n14720) );
  XNOR2_X1 U15877 ( .A(n14744), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n14737) );
  NAND2_X1 U15878 ( .A1(n14738), .A2(n14737), .ZN(n14736) );
  NAND2_X1 U15879 ( .A1(n13919), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n13905) );
  NAND2_X1 U15880 ( .A1(n14736), .A2(n13905), .ZN(n14760) );
  OR2_X1 U15881 ( .A1(n13922), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n13906) );
  NAND2_X1 U15882 ( .A1(n13922), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n13907) );
  AND2_X1 U15883 ( .A1(n13906), .A2(n13907), .ZN(n14759) );
  NAND2_X1 U15884 ( .A1(n14760), .A2(n14759), .ZN(n14758) );
  NAND2_X1 U15885 ( .A1(n14758), .A2(n13907), .ZN(n13908) );
  NOR2_X1 U15886 ( .A1(n13908), .A2(n14777), .ZN(n13909) );
  INV_X1 U15887 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14769) );
  NOR2_X1 U15888 ( .A1(n14768), .A2(n14769), .ZN(n14766) );
  NOR2_X1 U15889 ( .A1(n13910), .A2(n14766), .ZN(n13911) );
  XNOR2_X1 U15890 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n13911), .ZN(n13928) );
  MUX2_X1 U15891 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n11861), .S(n14708), .Z(
        n14711) );
  INV_X1 U15892 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n13914) );
  MUX2_X1 U15893 ( .A(n13914), .B(P1_REG1_REG_13__SCAN_IN), .S(n14699), .Z(
        n14692) );
  NOR2_X1 U15894 ( .A1(n14693), .A2(n14692), .ZN(n14691) );
  NAND2_X1 U15895 ( .A1(n14711), .A2(n14710), .ZN(n14709) );
  OAI21_X1 U15896 ( .B1(n14708), .B2(P1_REG1_REG_14__SCAN_IN), .A(n14709), 
        .ZN(n13915) );
  NAND2_X1 U15897 ( .A1(n13917), .A2(n13915), .ZN(n13918) );
  INV_X1 U15898 ( .A(n13915), .ZN(n13916) );
  INV_X1 U15899 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14726) );
  NAND2_X1 U15900 ( .A1(n14727), .A2(n14726), .ZN(n14725) );
  AND2_X2 U15901 ( .A1(n13918), .A2(n14725), .ZN(n14741) );
  XNOR2_X1 U15902 ( .A(n14744), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n14740) );
  NAND2_X1 U15903 ( .A1(n13919), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n13920) );
  NAND2_X1 U15904 ( .A1(n14739), .A2(n13920), .ZN(n14751) );
  INV_X1 U15905 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n13921) );
  XNOR2_X1 U15906 ( .A(n13922), .B(n13921), .ZN(n14750) );
  NOR2_X1 U15907 ( .A1(n13924), .A2(n13923), .ZN(n13925) );
  AOI21_X1 U15908 ( .B1(n13924), .B2(n13923), .A(n13925), .ZN(n14770) );
  AND2_X1 U15909 ( .A1(n14770), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n14771) );
  NOR2_X1 U15910 ( .A1(n14771), .A2(n13925), .ZN(n13926) );
  AOI22_X1 U15911 ( .A1(n13928), .A2(n14757), .B1(n14749), .B2(n13927), .ZN(
        n13931) );
  INV_X1 U15912 ( .A(n13927), .ZN(n13929) );
  INV_X1 U15913 ( .A(n13932), .ZN(n13933) );
  XNOR2_X1 U15914 ( .A(n13940), .B(n14282), .ZN(n13934) );
  NAND2_X1 U15915 ( .A1(n14172), .A2(n14849), .ZN(n13939) );
  AND2_X1 U15916 ( .A1(n13936), .A2(n13935), .ZN(n14174) );
  INV_X1 U15917 ( .A(n14174), .ZN(n13937) );
  NOR2_X1 U15918 ( .A1(n14842), .A2(n13937), .ZN(n13944) );
  AOI21_X1 U15919 ( .B1(n14842), .B2(P1_REG2_REG_31__SCAN_IN), .A(n13944), 
        .ZN(n13938) );
  OAI211_X1 U15920 ( .C1(n14282), .C2(n14845), .A(n13939), .B(n13938), .ZN(
        P1_U3263) );
  AOI211_X1 U15921 ( .C1(n13942), .C2(n13941), .A(n10182), .B(n13940), .ZN(
        n14175) );
  NAND2_X1 U15922 ( .A1(n14175), .A2(n14849), .ZN(n13946) );
  AND2_X1 U15923 ( .A1(n14842), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n13943) );
  NOR2_X1 U15924 ( .A1(n13944), .A2(n13943), .ZN(n13945) );
  OAI211_X1 U15925 ( .C1(n14286), .C2(n14845), .A(n13946), .B(n13945), .ZN(
        P1_U3264) );
  INV_X1 U15926 ( .A(n13947), .ZN(n13960) );
  OAI22_X1 U15927 ( .A1(n13950), .A2(n13949), .B1(n13948), .B2(n14831), .ZN(
        n13953) );
  NOR2_X1 U15928 ( .A1(n14842), .A2(n13951), .ZN(n13952) );
  AOI211_X1 U15929 ( .C1(n14842), .C2(P1_REG2_REG_29__SCAN_IN), .A(n13953), 
        .B(n13952), .ZN(n13955) );
  NAND2_X1 U15930 ( .A1(n14180), .A2(n14814), .ZN(n13954) );
  OAI211_X1 U15931 ( .C1(n13956), .C2(n14818), .A(n13955), .B(n13954), .ZN(
        n13957) );
  AOI21_X1 U15932 ( .B1(n13958), .B2(n14146), .A(n13957), .ZN(n13959) );
  OAI21_X1 U15933 ( .B1(n13960), .B2(n14161), .A(n13959), .ZN(P1_U3356) );
  XNOR2_X1 U15934 ( .A(n13961), .B(n13962), .ZN(n14181) );
  AOI21_X1 U15935 ( .B1(n14288), .B2(n13989), .A(n10182), .ZN(n13964) );
  NAND2_X1 U15936 ( .A1(n13964), .A2(n13963), .ZN(n14183) );
  INV_X1 U15937 ( .A(n13965), .ZN(n14182) );
  NAND2_X1 U15938 ( .A1(n14842), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n13968) );
  OR2_X1 U15939 ( .A1(n14831), .A2(n13966), .ZN(n13967) );
  OAI211_X1 U15940 ( .C1(n14842), .C2(n14182), .A(n13968), .B(n13967), .ZN(
        n13969) );
  AOI21_X1 U15941 ( .B1(n14288), .B2(n14814), .A(n13969), .ZN(n13970) );
  OAI21_X1 U15942 ( .B1(n14183), .B2(n14818), .A(n13970), .ZN(n13975) );
  OR2_X2 U15943 ( .A1(n6620), .A2(n13971), .ZN(n13972) );
  NOR2_X1 U15944 ( .A1(n14185), .A2(n14161), .ZN(n13974) );
  INV_X1 U15945 ( .A(n13976), .ZN(P1_U3265) );
  OAI21_X1 U15946 ( .B1(n13978), .B2(n13981), .A(n13977), .ZN(n13980) );
  AOI21_X1 U15947 ( .B1(n13980), .B2(n14269), .A(n13979), .ZN(n13986) );
  NAND2_X1 U15948 ( .A1(n13982), .A2(n13981), .ZN(n13983) );
  NAND2_X1 U15949 ( .A1(n13984), .A2(n13983), .ZN(n14189) );
  NAND2_X1 U15950 ( .A1(n14189), .A2(n14877), .ZN(n13985) );
  NOR2_X1 U15951 ( .A1(n14842), .A2(n13987), .ZN(n14851) );
  INV_X1 U15952 ( .A(n13988), .ZN(n14292) );
  AOI21_X1 U15953 ( .B1(n13988), .B2(n14001), .A(n10182), .ZN(n13990) );
  AND2_X1 U15954 ( .A1(n13990), .A2(n13989), .ZN(n14188) );
  NAND2_X1 U15955 ( .A1(n14188), .A2(n14849), .ZN(n13993) );
  AOI22_X1 U15956 ( .A1(n14842), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n13991), 
        .B2(n14841), .ZN(n13992) );
  OAI211_X1 U15957 ( .C1(n14292), .C2(n14845), .A(n13993), .B(n13992), .ZN(
        n13994) );
  AOI21_X1 U15958 ( .B1(n14189), .B2(n14851), .A(n13994), .ZN(n13995) );
  OAI21_X1 U15959 ( .B1(n14191), .B2(n14842), .A(n13995), .ZN(P1_U3266) );
  XNOR2_X1 U15960 ( .A(n13997), .B(n13996), .ZN(n14200) );
  OAI21_X1 U15961 ( .B1(n14000), .B2(n13999), .A(n13998), .ZN(n14198) );
  OAI211_X1 U15962 ( .C1(n14196), .C2(n14012), .A(n14837), .B(n14001), .ZN(
        n14195) );
  INV_X1 U15963 ( .A(n14002), .ZN(n14194) );
  OAI22_X1 U15964 ( .A1(n14842), .A2(n14194), .B1(n14003), .B2(n14831), .ZN(
        n14005) );
  NOR2_X1 U15965 ( .A1(n14196), .A2(n14845), .ZN(n14004) );
  AOI211_X1 U15966 ( .C1(n14842), .C2(P1_REG2_REG_26__SCAN_IN), .A(n14005), 
        .B(n14004), .ZN(n14006) );
  OAI21_X1 U15967 ( .B1(n14818), .B2(n14195), .A(n14006), .ZN(n14007) );
  AOI21_X1 U15968 ( .B1(n14198), .B2(n14146), .A(n14007), .ZN(n14008) );
  OAI21_X1 U15969 ( .B1(n14200), .B2(n14161), .A(n14008), .ZN(P1_U3267) );
  XNOR2_X1 U15970 ( .A(n14009), .B(n14020), .ZN(n14204) );
  NAND2_X1 U15971 ( .A1(n14201), .A2(n14035), .ZN(n14010) );
  NAND2_X1 U15972 ( .A1(n14010), .A2(n14837), .ZN(n14011) );
  OR2_X1 U15973 ( .A1(n14012), .A2(n14011), .ZN(n14203) );
  INV_X1 U15974 ( .A(n14013), .ZN(n14202) );
  NAND2_X1 U15975 ( .A1(n14842), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n14016) );
  OR2_X1 U15976 ( .A1(n14831), .A2(n14014), .ZN(n14015) );
  OAI211_X1 U15977 ( .C1(n14842), .C2(n14202), .A(n14016), .B(n14015), .ZN(
        n14017) );
  AOI21_X1 U15978 ( .B1(n14201), .B2(n14814), .A(n14017), .ZN(n14018) );
  OAI21_X1 U15979 ( .B1(n14203), .B2(n14818), .A(n14018), .ZN(n14023) );
  OAI21_X1 U15980 ( .B1(n14021), .B2(n14020), .A(n14019), .ZN(n14207) );
  NOR2_X1 U15981 ( .A1(n14207), .A2(n14161), .ZN(n14022) );
  AOI211_X1 U15982 ( .C1(n14204), .C2(n14146), .A(n14023), .B(n14022), .ZN(
        n14024) );
  INV_X1 U15983 ( .A(n14024), .ZN(P1_U3268) );
  AOI21_X1 U15984 ( .B1(n14026), .B2(n14025), .A(n14885), .ZN(n14029) );
  AOI21_X1 U15985 ( .B1(n14029), .B2(n14028), .A(n14027), .ZN(n14034) );
  NAND2_X1 U15986 ( .A1(n14031), .A2(n14030), .ZN(n14032) );
  NAND2_X1 U15987 ( .A1(n6596), .A2(n14032), .ZN(n14212) );
  NAND2_X1 U15988 ( .A1(n14212), .A2(n14877), .ZN(n14033) );
  NAND2_X1 U15989 ( .A1(n14034), .A2(n14033), .ZN(n14216) );
  INV_X1 U15990 ( .A(n14216), .ZN(n14042) );
  AOI21_X1 U15991 ( .B1(n14211), .B2(n14047), .A(n10182), .ZN(n14036) );
  NAND2_X1 U15992 ( .A1(n14036), .A2(n14035), .ZN(n14213) );
  AOI22_X1 U15993 ( .A1(n14842), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14037), 
        .B2(n14841), .ZN(n14039) );
  NAND2_X1 U15994 ( .A1(n14211), .A2(n14814), .ZN(n14038) );
  OAI211_X1 U15995 ( .C1(n14213), .C2(n14818), .A(n14039), .B(n14038), .ZN(
        n14040) );
  AOI21_X1 U15996 ( .B1(n14212), .B2(n14851), .A(n14040), .ZN(n14041) );
  OAI21_X1 U15997 ( .B1(n14042), .B2(n14842), .A(n14041), .ZN(P1_U3269) );
  XNOR2_X1 U15998 ( .A(n14043), .B(n14045), .ZN(n14225) );
  OAI21_X1 U15999 ( .B1(n14046), .B2(n14045), .A(n14044), .ZN(n14222) );
  NAND2_X1 U16000 ( .A1(n14222), .A2(n14146), .ZN(n14055) );
  INV_X1 U16001 ( .A(n14047), .ZN(n14048) );
  AOI211_X1 U16002 ( .C1(n14221), .C2(n14061), .A(n10182), .B(n14048), .ZN(
        n14219) );
  AOI22_X1 U16003 ( .A1(n14165), .A2(n14220), .B1(n14049), .B2(n14841), .ZN(
        n14051) );
  NAND2_X1 U16004 ( .A1(n14842), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n14050) );
  OAI211_X1 U16005 ( .C1(n14052), .C2(n14845), .A(n14051), .B(n14050), .ZN(
        n14053) );
  AOI21_X1 U16006 ( .B1(n14219), .B2(n14849), .A(n14053), .ZN(n14054) );
  OAI211_X1 U16007 ( .C1(n14225), .C2(n14161), .A(n14055), .B(n14054), .ZN(
        P1_U3270) );
  XNOR2_X1 U16008 ( .A(n14056), .B(n14066), .ZN(n14059) );
  INV_X1 U16009 ( .A(n14057), .ZN(n14058) );
  AOI21_X1 U16010 ( .B1(n14059), .B2(n14269), .A(n14058), .ZN(n14227) );
  AOI21_X1 U16011 ( .B1(n14305), .B2(n14075), .A(n10182), .ZN(n14062) );
  NAND2_X1 U16012 ( .A1(n14062), .A2(n14061), .ZN(n14226) );
  INV_X1 U16013 ( .A(n14226), .ZN(n14070) );
  AOI22_X1 U16014 ( .A1(n14842), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n14063), 
        .B2(n14841), .ZN(n14064) );
  OAI21_X1 U16015 ( .B1(n14065), .B2(n14845), .A(n14064), .ZN(n14069) );
  XNOR2_X1 U16016 ( .A(n14067), .B(n14066), .ZN(n14228) );
  NOR2_X1 U16017 ( .A1(n14228), .A2(n14161), .ZN(n14068) );
  AOI211_X1 U16018 ( .C1(n14070), .C2(n14849), .A(n14069), .B(n14068), .ZN(
        n14071) );
  OAI21_X1 U16019 ( .B1(n14842), .B2(n14227), .A(n14071), .ZN(P1_U3271) );
  XNOR2_X1 U16020 ( .A(n14072), .B(n14073), .ZN(n14238) );
  OAI21_X1 U16021 ( .B1(n6623), .B2(n8937), .A(n14074), .ZN(n14236) );
  INV_X1 U16022 ( .A(n14076), .ZN(n14233) );
  AOI211_X1 U16023 ( .C1(n14076), .C2(n14089), .A(n10182), .B(n14060), .ZN(
        n14235) );
  NAND2_X1 U16024 ( .A1(n14235), .A2(n14849), .ZN(n14081) );
  INV_X1 U16025 ( .A(n14077), .ZN(n14078) );
  OAI22_X1 U16026 ( .A1(n14842), .A2(n14232), .B1(n14078), .B2(n14831), .ZN(
        n14079) );
  AOI21_X1 U16027 ( .B1(P1_REG2_REG_21__SCAN_IN), .B2(n14842), .A(n14079), 
        .ZN(n14080) );
  OAI211_X1 U16028 ( .C1(n14233), .C2(n14845), .A(n14081), .B(n14080), .ZN(
        n14082) );
  AOI21_X1 U16029 ( .B1(n14236), .B2(n14789), .A(n14082), .ZN(n14083) );
  OAI21_X1 U16030 ( .B1(n14143), .B2(n14238), .A(n14083), .ZN(P1_U3272) );
  NAND2_X1 U16031 ( .A1(n14084), .A2(n8922), .ZN(n14085) );
  NAND3_X1 U16032 ( .A1(n14086), .A2(n14269), .A3(n14085), .ZN(n14088) );
  NAND2_X1 U16033 ( .A1(n14088), .A2(n14087), .ZN(n14245) );
  INV_X1 U16034 ( .A(n14245), .ZN(n14100) );
  AOI21_X1 U16035 ( .B1(n14240), .B2(n14103), .A(n10182), .ZN(n14090) );
  NAND2_X1 U16036 ( .A1(n14090), .A2(n14089), .ZN(n14241) );
  INV_X1 U16037 ( .A(n14241), .ZN(n14094) );
  AOI22_X1 U16038 ( .A1(n14842), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14091), 
        .B2(n14841), .ZN(n14092) );
  OAI21_X1 U16039 ( .B1(n6829), .B2(n14845), .A(n14092), .ZN(n14093) );
  AOI21_X1 U16040 ( .B1(n14094), .B2(n14849), .A(n14093), .ZN(n14099) );
  NAND2_X1 U16041 ( .A1(n14097), .A2(n14096), .ZN(n14239) );
  NAND3_X1 U16042 ( .A1(n14095), .A2(n14239), .A3(n14789), .ZN(n14098) );
  OAI211_X1 U16043 ( .C1(n14100), .C2(n14842), .A(n14099), .B(n14098), .ZN(
        P1_U3273) );
  XNOR2_X1 U16044 ( .A(n14101), .B(n6960), .ZN(n14254) );
  OAI21_X1 U16045 ( .B1(n6640), .B2(n6960), .A(n14102), .ZN(n14248) );
  AOI211_X1 U16046 ( .C1(n14251), .C2(n14121), .A(n10182), .B(n6830), .ZN(
        n14249) );
  NAND2_X1 U16047 ( .A1(n14249), .A2(n14104), .ZN(n14109) );
  INV_X1 U16048 ( .A(n14250), .ZN(n14106) );
  OAI22_X1 U16049 ( .A1(n14842), .A2(n14106), .B1(n14105), .B2(n14831), .ZN(
        n14107) );
  AOI21_X1 U16050 ( .B1(P1_REG2_REG_19__SCAN_IN), .B2(n14842), .A(n14107), 
        .ZN(n14108) );
  OAI211_X1 U16051 ( .C1(n14110), .C2(n14845), .A(n14109), .B(n14108), .ZN(
        n14111) );
  AOI21_X1 U16052 ( .B1(n14248), .B2(n14146), .A(n14111), .ZN(n14112) );
  OAI21_X1 U16053 ( .B1(n14254), .B2(n14161), .A(n14112), .ZN(P1_U3274) );
  XNOR2_X1 U16054 ( .A(n14113), .B(n14115), .ZN(n14119) );
  INV_X1 U16055 ( .A(n14119), .ZN(n14260) );
  INV_X1 U16056 ( .A(n14851), .ZN(n14131) );
  XNOR2_X1 U16057 ( .A(n14114), .B(n14115), .ZN(n14116) );
  NOR2_X1 U16058 ( .A1(n14116), .A2(n14885), .ZN(n14117) );
  AOI211_X1 U16059 ( .C1(n14877), .C2(n14119), .A(n14118), .B(n14117), .ZN(
        n14259) );
  INV_X1 U16060 ( .A(n14259), .ZN(n14120) );
  OAI21_X1 U16061 ( .B1(n14120), .B2(n14256), .A(n14165), .ZN(n14130) );
  INV_X1 U16062 ( .A(n14135), .ZN(n14123) );
  INV_X1 U16063 ( .A(n14121), .ZN(n14122) );
  AOI211_X1 U16064 ( .C1(n14257), .C2(n14123), .A(n10182), .B(n14122), .ZN(
        n14255) );
  INV_X1 U16065 ( .A(n14124), .ZN(n14125) );
  AOI22_X1 U16066 ( .A1(n14842), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14125), 
        .B2(n14841), .ZN(n14126) );
  OAI21_X1 U16067 ( .B1(n14127), .B2(n14845), .A(n14126), .ZN(n14128) );
  AOI21_X1 U16068 ( .B1(n14255), .B2(n14849), .A(n14128), .ZN(n14129) );
  OAI211_X1 U16069 ( .C1(n14260), .C2(n14131), .A(n14130), .B(n14129), .ZN(
        P1_U3275) );
  XNOR2_X1 U16070 ( .A(n14132), .B(n14133), .ZN(n14267) );
  XNOR2_X1 U16071 ( .A(n14134), .B(n14133), .ZN(n14261) );
  AOI211_X1 U16072 ( .C1(n14264), .C2(n14147), .A(n10182), .B(n14135), .ZN(
        n14262) );
  NOR2_X1 U16073 ( .A1(n14831), .A2(n14136), .ZN(n14137) );
  AOI211_X1 U16074 ( .C1(n14262), .C2(n14138), .A(n14137), .B(n14263), .ZN(
        n14140) );
  AOI22_X1 U16075 ( .A1(n14264), .A2(n14814), .B1(n14842), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n14139) );
  OAI21_X1 U16076 ( .B1(n14140), .B2(n14842), .A(n14139), .ZN(n14141) );
  AOI21_X1 U16077 ( .B1(n14789), .B2(n14261), .A(n14141), .ZN(n14142) );
  OAI21_X1 U16078 ( .B1(n14267), .B2(n14143), .A(n14142), .ZN(P1_U3276) );
  XNOR2_X1 U16079 ( .A(n14144), .B(n6514), .ZN(n14274) );
  OAI21_X1 U16080 ( .B1(n6641), .B2(n6514), .A(n14145), .ZN(n14270) );
  NAND2_X1 U16081 ( .A1(n14270), .A2(n14146), .ZN(n14160) );
  AOI211_X1 U16082 ( .C1(n14604), .C2(n14148), .A(n10182), .B(n7232), .ZN(
        n14268) );
  NAND2_X1 U16083 ( .A1(n14150), .A2(n14149), .ZN(n14153) );
  NAND2_X1 U16084 ( .A1(n14151), .A2(n13861), .ZN(n14152) );
  NAND2_X1 U16085 ( .A1(n14153), .A2(n14152), .ZN(n14606) );
  AOI22_X1 U16086 ( .A1(n14165), .A2(n14606), .B1(n14154), .B2(n14841), .ZN(
        n14156) );
  NAND2_X1 U16087 ( .A1(n14842), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n14155) );
  OAI211_X1 U16088 ( .C1(n14157), .C2(n14845), .A(n14156), .B(n14155), .ZN(
        n14158) );
  AOI21_X1 U16089 ( .B1(n14268), .B2(n14849), .A(n14158), .ZN(n14159) );
  OAI211_X1 U16090 ( .C1(n14274), .C2(n14161), .A(n14160), .B(n14159), .ZN(
        P1_U3277) );
  NAND2_X1 U16091 ( .A1(n14162), .A2(n14789), .ZN(n14171) );
  NAND2_X1 U16092 ( .A1(n14842), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n14163) );
  OAI21_X1 U16093 ( .B1(n14831), .B2(n14601), .A(n14163), .ZN(n14164) );
  AOI21_X1 U16094 ( .B1(n14597), .B2(n14814), .A(n14164), .ZN(n14170) );
  NAND2_X1 U16095 ( .A1(n14166), .A2(n14165), .ZN(n14169) );
  NAND2_X1 U16096 ( .A1(n14167), .A2(n14849), .ZN(n14168) );
  NAND4_X1 U16097 ( .A1(n14171), .A2(n14170), .A3(n14169), .A4(n14168), .ZN(
        P1_U3279) );
  INV_X1 U16098 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14173) );
  INV_X1 U16099 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n14176) );
  NOR2_X1 U16100 ( .A1(n14175), .A2(n14174), .ZN(n14283) );
  MUX2_X1 U16101 ( .A(n14176), .B(n14283), .S(n14896), .Z(n14177) );
  OAI21_X1 U16102 ( .B1(n14286), .B2(n14210), .A(n14177), .ZN(P1_U3558) );
  AND2_X1 U16103 ( .A1(n14183), .A2(n14182), .ZN(n14184) );
  INV_X1 U16104 ( .A(n14187), .ZN(P1_U3556) );
  AOI21_X1 U16105 ( .B1(n14189), .B2(n14866), .A(n14188), .ZN(n14190) );
  AND2_X2 U16106 ( .A1(n14191), .A2(n14190), .ZN(n14290) );
  INV_X1 U16107 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n14192) );
  MUX2_X1 U16108 ( .A(n14290), .B(n14192), .S(n14894), .Z(n14193) );
  OAI21_X1 U16109 ( .B1(n14292), .B2(n14210), .A(n14193), .ZN(P1_U3555) );
  OAI211_X1 U16110 ( .C1(n14196), .C2(n14872), .A(n14195), .B(n14194), .ZN(
        n14197) );
  AOI21_X1 U16111 ( .B1(n14198), .B2(n14269), .A(n14197), .ZN(n14199) );
  OAI21_X1 U16112 ( .B1(n14200), .B2(n14273), .A(n14199), .ZN(n14293) );
  MUX2_X1 U16113 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14293), .S(n14896), .Z(
        P1_U3554) );
  INV_X1 U16114 ( .A(n14201), .ZN(n14298) );
  AND2_X1 U16115 ( .A1(n14203), .A2(n14202), .ZN(n14206) );
  NAND2_X1 U16116 ( .A1(n14204), .A2(n14269), .ZN(n14205) );
  OAI211_X1 U16117 ( .C1(n14207), .C2(n14273), .A(n14206), .B(n14205), .ZN(
        n14294) );
  MUX2_X1 U16118 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14294), .S(n14896), .Z(
        n14208) );
  INV_X1 U16119 ( .A(n14208), .ZN(n14209) );
  OAI21_X1 U16120 ( .B1(n14298), .B2(n14210), .A(n14209), .ZN(P1_U3553) );
  INV_X1 U16121 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n14217) );
  NAND2_X1 U16122 ( .A1(n14212), .A2(n14866), .ZN(n14214) );
  OAI211_X1 U16123 ( .C1(n7230), .C2(n14872), .A(n14214), .B(n14213), .ZN(
        n14215) );
  NOR2_X1 U16124 ( .A1(n14216), .A2(n14215), .ZN(n14299) );
  MUX2_X1 U16125 ( .A(n14217), .B(n14299), .S(n14896), .Z(n14218) );
  INV_X1 U16126 ( .A(n14218), .ZN(P1_U3552) );
  AOI211_X1 U16127 ( .C1(n14221), .C2(n14881), .A(n14220), .B(n14219), .ZN(
        n14224) );
  NAND2_X1 U16128 ( .A1(n14222), .A2(n14269), .ZN(n14223) );
  OAI211_X1 U16129 ( .C1(n14225), .C2(n14273), .A(n14224), .B(n14223), .ZN(
        n14302) );
  MUX2_X1 U16130 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14302), .S(n14896), .Z(
        P1_U3551) );
  OAI211_X1 U16131 ( .C1(n14273), .C2(n14228), .A(n14227), .B(n14226), .ZN(
        n14303) );
  MUX2_X1 U16132 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14303), .S(n14896), .Z(
        n14229) );
  AOI21_X1 U16133 ( .B1(n14230), .B2(n14305), .A(n14229), .ZN(n14231) );
  INV_X1 U16134 ( .A(n14231), .ZN(P1_U3550) );
  OAI21_X1 U16135 ( .B1(n14233), .B2(n14872), .A(n14232), .ZN(n14234) );
  AOI211_X1 U16136 ( .C1(n14236), .C2(n14887), .A(n14235), .B(n14234), .ZN(
        n14237) );
  OAI21_X1 U16137 ( .B1(n14885), .B2(n14238), .A(n14237), .ZN(n14308) );
  MUX2_X1 U16138 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14308), .S(n14896), .Z(
        P1_U3549) );
  NAND3_X1 U16139 ( .A1(n14095), .A2(n14239), .A3(n14887), .ZN(n14243) );
  NAND2_X1 U16140 ( .A1(n14240), .A2(n14881), .ZN(n14242) );
  NAND3_X1 U16141 ( .A1(n14243), .A2(n14242), .A3(n14241), .ZN(n14244) );
  NOR2_X1 U16142 ( .A1(n14245), .A2(n14244), .ZN(n14309) );
  MUX2_X1 U16143 ( .A(n14246), .B(n14309), .S(n14896), .Z(n14247) );
  INV_X1 U16144 ( .A(n14247), .ZN(P1_U3548) );
  NAND2_X1 U16145 ( .A1(n14248), .A2(n14269), .ZN(n14253) );
  AOI211_X1 U16146 ( .C1(n14251), .C2(n14881), .A(n14250), .B(n14249), .ZN(
        n14252) );
  OAI211_X1 U16147 ( .C1(n14254), .C2(n14273), .A(n14253), .B(n14252), .ZN(
        n14312) );
  MUX2_X1 U16148 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14312), .S(n14896), .Z(
        P1_U3547) );
  AOI211_X1 U16149 ( .C1(n14257), .C2(n14881), .A(n14256), .B(n14255), .ZN(
        n14258) );
  OAI211_X1 U16150 ( .C1(n14260), .C2(n14868), .A(n14259), .B(n14258), .ZN(
        n14313) );
  MUX2_X1 U16151 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14313), .S(n14896), .Z(
        P1_U3546) );
  NAND2_X1 U16152 ( .A1(n14261), .A2(n14887), .ZN(n14266) );
  AOI211_X1 U16153 ( .C1(n14264), .C2(n14881), .A(n14263), .B(n14262), .ZN(
        n14265) );
  OAI211_X1 U16154 ( .C1(n14267), .C2(n14885), .A(n14266), .B(n14265), .ZN(
        n14314) );
  MUX2_X1 U16155 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14314), .S(n14896), .Z(
        P1_U3545) );
  AOI211_X1 U16156 ( .C1(n14604), .C2(n14881), .A(n14606), .B(n14268), .ZN(
        n14272) );
  NAND2_X1 U16157 ( .A1(n14270), .A2(n14269), .ZN(n14271) );
  OAI211_X1 U16158 ( .C1(n14274), .C2(n14273), .A(n14272), .B(n14271), .ZN(
        n14315) );
  MUX2_X1 U16159 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14315), .S(n14896), .Z(
        P1_U3544) );
  NAND2_X1 U16160 ( .A1(n14275), .A2(n14887), .ZN(n14278) );
  AOI211_X1 U16161 ( .C1(n14622), .C2(n14881), .A(n14626), .B(n14276), .ZN(
        n14277) );
  OAI211_X1 U16162 ( .C1(n14885), .C2(n14279), .A(n14278), .B(n14277), .ZN(
        n14316) );
  MUX2_X1 U16163 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n14316), .S(n14896), .Z(
        P1_U3543) );
  INV_X1 U16164 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n14281) );
  INV_X1 U16165 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n14284) );
  MUX2_X1 U16166 ( .A(n14284), .B(n14283), .S(n14891), .Z(n14285) );
  OAI21_X1 U16167 ( .B1(n14286), .B2(n14297), .A(n14285), .ZN(P1_U3526) );
  INV_X1 U16168 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n14289) );
  MUX2_X1 U16169 ( .A(n14290), .B(n14289), .S(n14889), .Z(n14291) );
  OAI21_X1 U16170 ( .B1(n14292), .B2(n14297), .A(n14291), .ZN(P1_U3523) );
  MUX2_X1 U16171 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14293), .S(n14891), .Z(
        P1_U3522) );
  MUX2_X1 U16172 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14294), .S(n14891), .Z(
        n14295) );
  INV_X1 U16173 ( .A(n14295), .ZN(n14296) );
  OAI21_X1 U16174 ( .B1(n14298), .B2(n14297), .A(n14296), .ZN(P1_U3521) );
  INV_X1 U16175 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n14300) );
  MUX2_X1 U16176 ( .A(n14300), .B(n14299), .S(n14891), .Z(n14301) );
  INV_X1 U16177 ( .A(n14301), .ZN(P1_U3520) );
  MUX2_X1 U16178 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14302), .S(n14891), .Z(
        P1_U3519) );
  MUX2_X1 U16179 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14303), .S(n14891), .Z(
        n14304) );
  AOI21_X1 U16180 ( .B1(n14306), .B2(n14305), .A(n14304), .ZN(n14307) );
  INV_X1 U16181 ( .A(n14307), .ZN(P1_U3518) );
  MUX2_X1 U16182 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14308), .S(n14891), .Z(
        P1_U3517) );
  INV_X1 U16183 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n14310) );
  MUX2_X1 U16184 ( .A(n14310), .B(n14309), .S(n14891), .Z(n14311) );
  INV_X1 U16185 ( .A(n14311), .ZN(P1_U3516) );
  MUX2_X1 U16186 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14312), .S(n14891), .Z(
        P1_U3515) );
  MUX2_X1 U16187 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14313), .S(n14891), .Z(
        P1_U3513) );
  MUX2_X1 U16188 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14314), .S(n14891), .Z(
        P1_U3510) );
  MUX2_X1 U16189 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14315), .S(n14891), .Z(
        P1_U3507) );
  MUX2_X1 U16190 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n14316), .S(n14891), .Z(
        P1_U3504) );
  INV_X1 U16191 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n14317) );
  NAND3_X1 U16192 ( .A1(n14317), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n14319) );
  OAI22_X1 U16193 ( .A1(n14320), .A2(n14319), .B1(n14318), .B2(n14347), .ZN(
        n14321) );
  AOI21_X1 U16194 ( .B1(n14323), .B2(n14322), .A(n14321), .ZN(n14324) );
  INV_X1 U16195 ( .A(n14324), .ZN(P1_U3324) );
  OAI222_X1 U16196 ( .A1(n14347), .A2(n14328), .B1(n14327), .B2(n14326), .C1(
        n14325), .C2(P1_U3086), .ZN(P1_U3325) );
  OAI222_X1 U16197 ( .A1(n14347), .A2(n14330), .B1(n14327), .B2(n14329), .C1(
        n8549), .C2(P1_U3086), .ZN(P1_U3326) );
  OAI222_X1 U16198 ( .A1(n14347), .A2(n14333), .B1(n14327), .B2(n14332), .C1(
        P1_U3086), .C2(n14331), .ZN(P1_U3327) );
  OAI222_X1 U16199 ( .A1(n14347), .A2(n14336), .B1(n14327), .B2(n14335), .C1(
        n6487), .C2(P1_U3086), .ZN(P1_U3328) );
  OAI222_X1 U16200 ( .A1(n14339), .A2(P1_U3086), .B1(n14327), .B2(n14338), 
        .C1(n14337), .C2(n14347), .ZN(P1_U3329) );
  OAI222_X1 U16201 ( .A1(n14347), .A2(n14342), .B1(n14327), .B2(n14341), .C1(
        n14340), .C2(P1_U3086), .ZN(P1_U3330) );
  OAI222_X1 U16202 ( .A1(n14347), .A2(n14346), .B1(n14327), .B2(n14345), .C1(
        n14344), .C2(P1_U3086), .ZN(P1_U3331) );
  MUX2_X1 U16203 ( .A(n14349), .B(n14348), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U16204 ( .A(n14350), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16205 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14765) );
  INV_X1 U16206 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14381) );
  INV_X1 U16207 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14379) );
  INV_X1 U16208 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14376) );
  INV_X1 U16209 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14374) );
  XNOR2_X1 U16210 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(P3_ADDR_REG_9__SCAN_IN), 
        .ZN(n14425) );
  NOR2_X1 U16211 ( .A1(n14352), .A2(n14353), .ZN(n14355) );
  NOR2_X1 U16212 ( .A1(n14358), .A2(n14359), .ZN(n14361) );
  NOR2_X1 U16213 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14362), .ZN(n14364) );
  NOR2_X1 U16214 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14365), .ZN(n14368) );
  XNOR2_X1 U16215 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n14365), .ZN(n14418) );
  XNOR2_X1 U16216 ( .A(n15398), .B(P1_ADDR_REG_8__SCAN_IN), .ZN(n14396) );
  INV_X1 U16217 ( .A(n14395), .ZN(n14372) );
  XOR2_X1 U16218 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n14394) );
  INV_X1 U16219 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14690) );
  XOR2_X1 U16220 ( .A(n14376), .B(n14690), .Z(n14392) );
  INV_X1 U16221 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14377) );
  NAND2_X1 U16222 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(n14377), .ZN(n14378) );
  INV_X1 U16223 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14702) );
  NOR2_X1 U16224 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14702), .ZN(n14380) );
  INV_X1 U16225 ( .A(n14436), .ZN(n14384) );
  INV_X1 U16226 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14719) );
  NAND2_X1 U16227 ( .A1(P3_ADDR_REG_14__SCAN_IN), .A2(n14719), .ZN(n14383) );
  INV_X1 U16228 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14382) );
  NAND2_X1 U16229 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14385), .ZN(n14386) );
  INV_X1 U16230 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14735) );
  AOI22_X1 U16231 ( .A1(n14440), .A2(n14386), .B1(P3_ADDR_REG_15__SCAN_IN), 
        .B2(n14735), .ZN(n14444) );
  INV_X1 U16232 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14748) );
  NAND2_X1 U16233 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n14748), .ZN(n14387) );
  INV_X1 U16234 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14443) );
  AOI22_X1 U16235 ( .A1(n14444), .A2(n14387), .B1(P1_ADDR_REG_16__SCAN_IN), 
        .B2(n14443), .ZN(n14388) );
  AND2_X1 U16236 ( .A1(n14765), .A2(n14388), .ZN(n14390) );
  XNOR2_X1 U16237 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14388), .ZN(n14447) );
  AND2_X1 U16238 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14447), .ZN(n14389) );
  INV_X1 U16239 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14474) );
  NOR2_X1 U16240 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n14474), .ZN(n14391) );
  AOI21_X1 U16241 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n14474), .A(n14391), 
        .ZN(n14472) );
  XNOR2_X1 U16242 ( .A(n14471), .B(n14472), .ZN(n14479) );
  INV_X1 U16243 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15031) );
  INV_X1 U16244 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15016) );
  INV_X1 U16245 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15002) );
  INV_X1 U16246 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15387) );
  XOR2_X1 U16247 ( .A(n14393), .B(n14392), .Z(n14428) );
  INV_X1 U16248 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14976) );
  XNOR2_X1 U16249 ( .A(n14395), .B(n14394), .ZN(n14465) );
  XOR2_X1 U16250 ( .A(n14397), .B(n14396), .Z(n14422) );
  OR2_X1 U16251 ( .A1(n14399), .A2(n14400), .ZN(n14410) );
  INV_X1 U16252 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14454) );
  XNOR2_X1 U16253 ( .A(n6547), .B(n14401), .ZN(n14452) );
  NAND2_X1 U16254 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14404), .ZN(n14406) );
  AOI21_X1 U16255 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n15157), .A(n14403), .ZN(
        n15449) );
  NOR2_X1 U16256 ( .A1(n15449), .A2(n15448), .ZN(n15457) );
  XOR2_X1 U16257 ( .A(n14404), .B(P2_ADDR_REG_1__SCAN_IN), .Z(n15456) );
  NAND2_X1 U16258 ( .A1(n15457), .A2(n15456), .ZN(n14405) );
  NAND2_X1 U16259 ( .A1(n14452), .A2(n14453), .ZN(n14407) );
  NOR2_X1 U16260 ( .A1(n14452), .A2(n14453), .ZN(n14451) );
  XNOR2_X1 U16261 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14408), .ZN(n15454) );
  NOR2_X1 U16262 ( .A1(n15453), .A2(n15454), .ZN(n14409) );
  NAND2_X1 U16263 ( .A1(n15453), .A2(n15454), .ZN(n15452) );
  XNOR2_X1 U16264 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n14411), .ZN(n14412) );
  NAND2_X1 U16265 ( .A1(n14414), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14417) );
  XNOR2_X1 U16266 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n14416) );
  XOR2_X1 U16267 ( .A(n14416), .B(n14415), .Z(n14456) );
  NAND2_X1 U16268 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14419), .ZN(n14420) );
  XNOR2_X1 U16269 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14418), .ZN(n15451) );
  NOR2_X1 U16270 ( .A1(n14422), .A2(n14421), .ZN(n14423) );
  XNOR2_X1 U16271 ( .A(n14425), .B(n14424), .ZN(n14461) );
  INV_X1 U16272 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14962) );
  NAND2_X1 U16273 ( .A1(n14460), .A2(n14461), .ZN(n14459) );
  NAND2_X1 U16274 ( .A1(n14465), .A2(n14464), .ZN(n14426) );
  NOR2_X1 U16275 ( .A1(n14465), .A2(n14464), .ZN(n14463) );
  NOR2_X1 U16276 ( .A1(n14428), .A2(n14427), .ZN(n14650) );
  NOR2_X1 U16277 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n14649), .ZN(n14429) );
  XNOR2_X1 U16278 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n14431) );
  XNOR2_X1 U16279 ( .A(n14431), .B(n14430), .ZN(n14653) );
  XOR2_X1 U16280 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .Z(n14432) );
  XOR2_X1 U16281 ( .A(n14433), .B(n14432), .Z(n14434) );
  XNOR2_X1 U16282 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n14437) );
  XNOR2_X1 U16283 ( .A(n14437), .B(n14436), .ZN(n14438) );
  XNOR2_X1 U16284 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n14441) );
  XNOR2_X1 U16285 ( .A(n14441), .B(n14440), .ZN(n14663) );
  NAND2_X1 U16286 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14443), .ZN(n14442) );
  OAI21_X1 U16287 ( .B1(n14443), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n14442), 
        .ZN(n14445) );
  XNOR2_X1 U16288 ( .A(n14445), .B(n14444), .ZN(n14668) );
  NAND2_X1 U16289 ( .A1(n14667), .A2(n14668), .ZN(n14446) );
  XNOR2_X1 U16290 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14447), .ZN(n14468) );
  NAND2_X1 U16291 ( .A1(n14469), .A2(n14468), .ZN(n14448) );
  XNOR2_X1 U16292 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14481), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16293 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14449) );
  OAI21_X1 U16294 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14449), 
        .ZN(U28) );
  AOI21_X1 U16295 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14450) );
  OAI21_X1 U16296 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14450), 
        .ZN(U29) );
  AOI21_X1 U16297 ( .B1(n14453), .B2(n14452), .A(n14451), .ZN(n14455) );
  XNOR2_X1 U16298 ( .A(n14455), .B(n14454), .ZN(SUB_1596_U61) );
  XOR2_X1 U16299 ( .A(n14457), .B(n14456), .Z(SUB_1596_U57) );
  XNOR2_X1 U16300 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14458), .ZN(SUB_1596_U55)
         );
  OAI21_X1 U16301 ( .B1(n14461), .B2(n14460), .A(n14459), .ZN(n14462) );
  XNOR2_X1 U16302 ( .A(n14462), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(SUB_1596_U54)
         );
  AOI21_X1 U16303 ( .B1(n14465), .B2(n14464), .A(n14463), .ZN(n14466) );
  XNOR2_X1 U16304 ( .A(n14466), .B(n14976), .ZN(SUB_1596_U70) );
  AOI21_X1 U16305 ( .B1(n14469), .B2(n14468), .A(n14467), .ZN(n14470) );
  XNOR2_X1 U16306 ( .A(n14470), .B(n15031), .ZN(SUB_1596_U63) );
  NAND2_X1 U16307 ( .A1(n14472), .A2(n14471), .ZN(n14473) );
  OAI21_X1 U16308 ( .B1(n14474), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n14473), 
        .ZN(n14478) );
  XNOR2_X1 U16309 ( .A(n14475), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n14476) );
  XNOR2_X1 U16310 ( .A(n14476), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n14477) );
  XNOR2_X1 U16311 ( .A(n14478), .B(n14477), .ZN(n14482) );
  XOR2_X1 U16312 ( .A(n14483), .B(n14484), .Z(n14519) );
  XNOR2_X1 U16313 ( .A(n14485), .B(n14484), .ZN(n14486) );
  OAI222_X1 U16314 ( .A1(n15182), .A2(n14488), .B1(n15183), .B2(n14487), .C1(
        n14486), .C2(n15206), .ZN(n14517) );
  AOI21_X1 U16315 ( .B1(n14519), .B2(n14489), .A(n14517), .ZN(n14493) );
  AND2_X1 U16316 ( .A1(n14490), .A2(n15188), .ZN(n14518) );
  AOI22_X1 U16317 ( .A1(n14518), .A2(n14508), .B1(n15209), .B2(n14491), .ZN(
        n14492) );
  OAI221_X1 U16318 ( .B1(n15214), .B2(n14493), .C1(n12749), .C2(n12385), .A(
        n14492), .ZN(P3_U3220) );
  XNOR2_X1 U16319 ( .A(n14495), .B(n14494), .ZN(n14498) );
  AOI222_X1 U16320 ( .A1(n14499), .A2(n14498), .B1(n14497), .B2(n15200), .C1(
        n14496), .C2(n15203), .ZN(n14525) );
  AOI22_X1 U16321 ( .A1(n15214), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n15209), 
        .B2(n14500), .ZN(n14511) );
  INV_X1 U16322 ( .A(n14501), .ZN(n14504) );
  OAI21_X1 U16323 ( .B1(n14504), .B2(n14503), .A(n14502), .ZN(n14506) );
  NAND2_X1 U16324 ( .A1(n14506), .A2(n14505), .ZN(n14528) );
  NOR2_X1 U16325 ( .A1(n14507), .A2(n15195), .ZN(n14527) );
  AOI22_X1 U16326 ( .A1(n14528), .A2(n14509), .B1(n14508), .B2(n14527), .ZN(
        n14510) );
  OAI211_X1 U16327 ( .C1(n15214), .C2(n14525), .A(n14511), .B(n14510), .ZN(
        P3_U3222) );
  OR2_X1 U16328 ( .A1(n14512), .A2(n15195), .ZN(n14513) );
  AOI22_X1 U16329 ( .A1(n15254), .A2(n14530), .B1(n8226), .B2(n12766), .ZN(
        P3_U3490) );
  OAI21_X1 U16330 ( .B1(n14515), .B2(n15195), .A(n14514), .ZN(n14531) );
  OAI22_X1 U16331 ( .A1(n12766), .A2(n14531), .B1(P3_REG1_REG_30__SCAN_IN), 
        .B2(n15254), .ZN(n14516) );
  INV_X1 U16332 ( .A(n14516), .ZN(P3_U3489) );
  AOI211_X1 U16333 ( .C1(n14519), .C2(n8531), .A(n14518), .B(n14517), .ZN(
        n14534) );
  AOI22_X1 U16334 ( .A1(n15254), .A2(n14534), .B1(n8014), .B2(n12766), .ZN(
        P3_U3472) );
  OAI22_X1 U16335 ( .A1(n14522), .A2(n14521), .B1(n14520), .B2(n15195), .ZN(
        n14523) );
  NOR2_X1 U16336 ( .A1(n14524), .A2(n14523), .ZN(n14536) );
  AOI22_X1 U16337 ( .A1(n15254), .A2(n14536), .B1(n12376), .B2(n12766), .ZN(
        P3_U3471) );
  INV_X1 U16338 ( .A(n14525), .ZN(n14526) );
  AOI211_X1 U16339 ( .C1(n8531), .C2(n14528), .A(n14527), .B(n14526), .ZN(
        n14538) );
  AOI22_X1 U16340 ( .A1(n15254), .A2(n14538), .B1(n7967), .B2(n12766), .ZN(
        P3_U3470) );
  INV_X1 U16341 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n14529) );
  AOI22_X1 U16342 ( .A1(n15246), .A2(n14530), .B1(n14529), .B2(n15244), .ZN(
        P3_U3458) );
  OAI22_X1 U16343 ( .A1(n15244), .A2(n14531), .B1(P3_REG0_REG_30__SCAN_IN), 
        .B2(n15246), .ZN(n14532) );
  INV_X1 U16344 ( .A(n14532), .ZN(P3_U3457) );
  INV_X1 U16345 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14533) );
  AOI22_X1 U16346 ( .A1(n15246), .A2(n14534), .B1(n14533), .B2(n15244), .ZN(
        P3_U3429) );
  INV_X1 U16347 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14535) );
  AOI22_X1 U16348 ( .A1(n15246), .A2(n14536), .B1(n14535), .B2(n15244), .ZN(
        P3_U3426) );
  INV_X1 U16349 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14537) );
  AOI22_X1 U16350 ( .A1(n15246), .A2(n14538), .B1(n14537), .B2(n15244), .ZN(
        P3_U3423) );
  OAI22_X1 U16351 ( .A1(n14542), .A2(n14541), .B1(n14540), .B2(n14539), .ZN(
        n14553) );
  INV_X1 U16352 ( .A(n14543), .ZN(n14544) );
  OAI21_X1 U16353 ( .B1(n14546), .B2(n14545), .A(n14544), .ZN(n14547) );
  AOI222_X1 U16354 ( .A1(n14916), .A2(n14559), .B1(n14553), .B2(n14914), .C1(
        n14547), .C2(n14912), .ZN(n14549) );
  OAI211_X1 U16355 ( .C1(n14551), .C2(n14550), .A(n14549), .B(n14548), .ZN(
        P2_U3187) );
  XOR2_X1 U16356 ( .A(n14557), .B(n14552), .Z(n14554) );
  AOI21_X1 U16357 ( .B1(n14554), .B2(n14579), .A(n14553), .ZN(n14567) );
  AOI222_X1 U16358 ( .A1(n14559), .A2(n14556), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n15076), .C1(n15051), .C2(n14555), .ZN(n14565) );
  XNOR2_X1 U16359 ( .A(n14558), .B(n14557), .ZN(n14571) );
  OAI211_X1 U16360 ( .C1(n7182), .C2(n7183), .A(n14562), .B(n14561), .ZN(
        n14566) );
  INV_X1 U16361 ( .A(n14566), .ZN(n14563) );
  AOI22_X1 U16362 ( .A1(n14571), .A2(n15059), .B1(n14563), .B2(n15049), .ZN(
        n14564) );
  OAI211_X1 U16363 ( .C1(n15076), .C2(n14567), .A(n14565), .B(n14564), .ZN(
        P2_U3251) );
  OAI21_X1 U16364 ( .B1(n7182), .B2(n15114), .A(n14566), .ZN(n14569) );
  INV_X1 U16365 ( .A(n14567), .ZN(n14568) );
  AOI211_X1 U16366 ( .C1(n14571), .C2(n14570), .A(n14569), .B(n14568), .ZN(
        n14589) );
  AOI22_X1 U16367 ( .A1(n15145), .A2(n14589), .B1(n10584), .B2(n15142), .ZN(
        P2_U3513) );
  AOI21_X1 U16368 ( .B1(n14573), .B2(n15123), .A(n14572), .ZN(n14575) );
  OAI211_X1 U16369 ( .C1(n14577), .C2(n14576), .A(n14575), .B(n14574), .ZN(
        n14578) );
  AOI21_X1 U16370 ( .B1(n14580), .B2(n14579), .A(n14578), .ZN(n14591) );
  AOI22_X1 U16371 ( .A1(n15145), .A2(n14591), .B1(n10240), .B2(n15142), .ZN(
        P2_U3512) );
  OAI21_X1 U16372 ( .B1(n14582), .B2(n15114), .A(n14581), .ZN(n14583) );
  AOI21_X1 U16373 ( .B1(n14584), .B2(n15124), .A(n14583), .ZN(n14585) );
  AOI22_X1 U16374 ( .A1(n15145), .A2(n14593), .B1(n14587), .B2(n15142), .ZN(
        P2_U3511) );
  INV_X1 U16375 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14588) );
  AOI22_X1 U16376 ( .A1(n15134), .A2(n14589), .B1(n14588), .B2(n15132), .ZN(
        P2_U3472) );
  INV_X1 U16377 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14590) );
  AOI22_X1 U16378 ( .A1(n15134), .A2(n14591), .B1(n14590), .B2(n15132), .ZN(
        P2_U3469) );
  INV_X1 U16379 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14592) );
  AOI22_X1 U16380 ( .A1(n15134), .A2(n14593), .B1(n14592), .B2(n15132), .ZN(
        P2_U3466) );
  OAI21_X1 U16381 ( .B1(n14596), .B2(n14595), .A(n14594), .ZN(n14598) );
  AOI222_X1 U16382 ( .A1(n14599), .A2(n14625), .B1(n14598), .B2(n14623), .C1(
        n14597), .C2(n14621), .ZN(n14600) );
  NAND2_X1 U16383 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14717)
         );
  OAI211_X1 U16384 ( .C1(n14629), .C2(n14601), .A(n14600), .B(n14717), .ZN(
        P1_U3215) );
  XNOR2_X1 U16385 ( .A(n14603), .B(n14602), .ZN(n14605) );
  AOI222_X1 U16386 ( .A1(n14606), .A2(n14625), .B1(n14623), .B2(n14605), .C1(
        n14604), .C2(n14621), .ZN(n14607) );
  NAND2_X1 U16387 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n14746)
         );
  OAI211_X1 U16388 ( .C1(n14629), .C2(n14608), .A(n14607), .B(n14746), .ZN(
        P1_U3226) );
  AND2_X1 U16389 ( .A1(n14610), .A2(n14609), .ZN(n14613) );
  OAI21_X1 U16390 ( .B1(n14613), .B2(n14612), .A(n14611), .ZN(n14614) );
  AOI222_X1 U16391 ( .A1(n14615), .A2(n14625), .B1(n14614), .B2(n14623), .C1(
        n14630), .C2(n14621), .ZN(n14616) );
  NAND2_X1 U16392 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14688)
         );
  OAI211_X1 U16393 ( .C1(n14629), .C2(n14617), .A(n14616), .B(n14688), .ZN(
        P1_U3236) );
  OAI21_X1 U16394 ( .B1(n14620), .B2(n14619), .A(n14618), .ZN(n14624) );
  AOI222_X1 U16395 ( .A1(n14626), .A2(n14625), .B1(n14624), .B2(n14623), .C1(
        n14622), .C2(n14621), .ZN(n14627) );
  NAND2_X1 U16396 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14733)
         );
  OAI211_X1 U16397 ( .C1(n14629), .C2(n14628), .A(n14627), .B(n14733), .ZN(
        P1_U3241) );
  INV_X1 U16398 ( .A(n14630), .ZN(n14635) );
  NAND2_X1 U16399 ( .A1(n14631), .A2(n14849), .ZN(n14634) );
  AOI22_X1 U16400 ( .A1(n14842), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n14632), 
        .B2(n14841), .ZN(n14633) );
  OAI211_X1 U16401 ( .C1(n14635), .C2(n14845), .A(n14634), .B(n14633), .ZN(
        n14636) );
  AOI21_X1 U16402 ( .B1(n14637), .B2(n14789), .A(n14636), .ZN(n14638) );
  OAI21_X1 U16403 ( .B1(n14842), .B2(n14639), .A(n14638), .ZN(P1_U3282) );
  OAI211_X1 U16404 ( .C1(n14642), .C2(n14872), .A(n14641), .B(n14640), .ZN(
        n14645) );
  NOR2_X1 U16405 ( .A1(n14643), .A2(n14885), .ZN(n14644) );
  AOI211_X1 U16406 ( .C1(n14887), .C2(n14646), .A(n14645), .B(n14644), .ZN(
        n14648) );
  AOI22_X1 U16407 ( .A1(n14896), .A2(n14648), .B1(n13914), .B2(n14894), .ZN(
        P1_U3541) );
  INV_X1 U16408 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14647) );
  AOI22_X1 U16409 ( .A1(n14891), .A2(n14648), .B1(n14647), .B2(n14889), .ZN(
        P1_U3498) );
  NOR2_X1 U16410 ( .A1(n14650), .A2(n14649), .ZN(n14651) );
  XOR2_X1 U16411 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n14651), .Z(SUB_1596_U69)
         );
  AOI21_X1 U16412 ( .B1(n14654), .B2(n14653), .A(n14652), .ZN(n14655) );
  XNOR2_X1 U16413 ( .A(n14655), .B(n15387), .ZN(SUB_1596_U68) );
  NOR2_X1 U16414 ( .A1(n14657), .A2(n14656), .ZN(n14658) );
  XOR2_X1 U16415 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n14658), .Z(SUB_1596_U67)
         );
  NOR2_X1 U16416 ( .A1(n14660), .A2(n14659), .ZN(n14661) );
  XOR2_X1 U16417 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n14661), .Z(SUB_1596_U66)
         );
  AOI21_X1 U16418 ( .B1(n14664), .B2(n14663), .A(n14662), .ZN(n14665) );
  XNOR2_X1 U16419 ( .A(n14665), .B(n15002), .ZN(SUB_1596_U65) );
  AOI21_X1 U16420 ( .B1(n14668), .B2(n14667), .A(n14666), .ZN(n14669) );
  XNOR2_X1 U16421 ( .A(n14669), .B(n15016), .ZN(SUB_1596_U64) );
  OAI21_X1 U16422 ( .B1(n14671), .B2(P1_REG1_REG_0__SCAN_IN), .A(n14670), .ZN(
        n14672) );
  XOR2_X1 U16423 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14672), .Z(n14676) );
  AOI22_X1 U16424 ( .A1(n14673), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14674) );
  OAI21_X1 U16425 ( .B1(n14676), .B2(n14675), .A(n14674), .ZN(P1_U3243) );
  OAI21_X1 U16426 ( .B1(n14679), .B2(n14678), .A(n14677), .ZN(n14687) );
  INV_X1 U16427 ( .A(n14680), .ZN(n14681) );
  NOR2_X1 U16428 ( .A1(n14752), .A2(n14681), .ZN(n14686) );
  AOI211_X1 U16429 ( .C1(n14684), .C2(n14683), .A(n14767), .B(n14682), .ZN(
        n14685) );
  AOI211_X1 U16430 ( .C1(n14749), .C2(n14687), .A(n14686), .B(n14685), .ZN(
        n14689) );
  OAI211_X1 U16431 ( .C1(n14690), .C2(n14781), .A(n14689), .B(n14688), .ZN(
        P1_U3254) );
  AOI211_X1 U16432 ( .C1(n14693), .C2(n14692), .A(n14691), .B(n14772), .ZN(
        n14698) );
  AOI211_X1 U16433 ( .C1(n14696), .C2(n14695), .A(n14694), .B(n14767), .ZN(
        n14697) );
  AOI211_X1 U16434 ( .C1(n14778), .C2(n14699), .A(n14698), .B(n14697), .ZN(
        n14701) );
  OAI211_X1 U16435 ( .C1(n14702), .C2(n14781), .A(n14701), .B(n14700), .ZN(
        P1_U3256) );
  NAND2_X1 U16436 ( .A1(n14704), .A2(n14703), .ZN(n14707) );
  INV_X1 U16437 ( .A(n14705), .ZN(n14706) );
  NAND2_X1 U16438 ( .A1(n14707), .A2(n14706), .ZN(n14715) );
  NAND2_X1 U16439 ( .A1(n14778), .A2(n14708), .ZN(n14714) );
  OAI21_X1 U16440 ( .B1(n14711), .B2(n14710), .A(n14709), .ZN(n14712) );
  NAND2_X1 U16441 ( .A1(n14749), .A2(n14712), .ZN(n14713) );
  OAI211_X1 U16442 ( .C1(n14767), .C2(n14715), .A(n14714), .B(n14713), .ZN(
        n14716) );
  INV_X1 U16443 ( .A(n14716), .ZN(n14718) );
  OAI211_X1 U16444 ( .C1(n14719), .C2(n14781), .A(n14718), .B(n14717), .ZN(
        P1_U3257) );
  OAI21_X1 U16445 ( .B1(n14722), .B2(n14721), .A(n14720), .ZN(n14723) );
  INV_X1 U16446 ( .A(n14723), .ZN(n14731) );
  NAND2_X1 U16447 ( .A1(n14778), .A2(n14724), .ZN(n14730) );
  OAI21_X1 U16448 ( .B1(n14727), .B2(n14726), .A(n14725), .ZN(n14728) );
  NAND2_X1 U16449 ( .A1(n14749), .A2(n14728), .ZN(n14729) );
  OAI211_X1 U16450 ( .C1(n14767), .C2(n14731), .A(n14730), .B(n14729), .ZN(
        n14732) );
  INV_X1 U16451 ( .A(n14732), .ZN(n14734) );
  OAI211_X1 U16452 ( .C1(n14735), .C2(n14781), .A(n14734), .B(n14733), .ZN(
        P1_U3258) );
  OAI211_X1 U16453 ( .C1(n14738), .C2(n14737), .A(n14736), .B(n14757), .ZN(
        n14743) );
  OAI211_X1 U16454 ( .C1(n14741), .C2(n14740), .A(n14739), .B(n14749), .ZN(
        n14742) );
  OAI211_X1 U16455 ( .C1(n14752), .C2(n14744), .A(n14743), .B(n14742), .ZN(
        n14745) );
  INV_X1 U16456 ( .A(n14745), .ZN(n14747) );
  OAI211_X1 U16457 ( .C1(n14748), .C2(n14781), .A(n14747), .B(n14746), .ZN(
        P1_U3259) );
  OAI21_X1 U16458 ( .B1(n14751), .B2(n14750), .A(n14749), .ZN(n14755) );
  OAI22_X1 U16459 ( .A1(n14755), .A2(n14754), .B1(n14753), .B2(n14752), .ZN(
        n14756) );
  INV_X1 U16460 ( .A(n14756), .ZN(n14762) );
  OAI211_X1 U16461 ( .C1(n14760), .C2(n14759), .A(n14758), .B(n14757), .ZN(
        n14761) );
  AND2_X1 U16462 ( .A1(n14762), .A2(n14761), .ZN(n14764) );
  OAI211_X1 U16463 ( .C1(n14765), .C2(n14781), .A(n14764), .B(n14763), .ZN(
        P1_U3260) );
  INV_X1 U16464 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14782) );
  AOI211_X1 U16465 ( .C1(n14769), .C2(n14768), .A(n14767), .B(n14766), .ZN(
        n14776) );
  INV_X1 U16466 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14774) );
  INV_X1 U16467 ( .A(n14770), .ZN(n14773) );
  AOI211_X1 U16468 ( .C1(n14774), .C2(n14773), .A(n14772), .B(n14771), .ZN(
        n14775) );
  AOI211_X1 U16469 ( .C1(n14778), .C2(n14777), .A(n14776), .B(n14775), .ZN(
        n14780) );
  OAI211_X1 U16470 ( .C1(n14782), .C2(n14781), .A(n14780), .B(n14779), .ZN(
        P1_U3261) );
  NAND2_X1 U16471 ( .A1(n14783), .A2(n14849), .ZN(n14786) );
  AOI22_X1 U16472 ( .A1(n14842), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n14784), 
        .B2(n14841), .ZN(n14785) );
  OAI211_X1 U16473 ( .C1(n14787), .C2(n14845), .A(n14786), .B(n14785), .ZN(
        n14788) );
  AOI21_X1 U16474 ( .B1(n14790), .B2(n14789), .A(n14788), .ZN(n14791) );
  OAI21_X1 U16475 ( .B1(n14842), .B2(n14792), .A(n14791), .ZN(P1_U3283) );
  NAND2_X1 U16476 ( .A1(n14793), .A2(n14849), .ZN(n14796) );
  AOI22_X1 U16477 ( .A1(n14842), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n14794), 
        .B2(n14841), .ZN(n14795) );
  OAI211_X1 U16478 ( .C1(n14797), .C2(n14845), .A(n14796), .B(n14795), .ZN(
        n14798) );
  AOI21_X1 U16479 ( .B1(n14799), .B2(n14851), .A(n14798), .ZN(n14800) );
  OAI21_X1 U16480 ( .B1(n14842), .B2(n14801), .A(n14800), .ZN(P1_U3284) );
  NOR2_X1 U16481 ( .A1(n14831), .A2(n14802), .ZN(n14803) );
  AOI21_X1 U16482 ( .B1(n14842), .B2(P1_REG2_REG_6__SCAN_IN), .A(n14803), .ZN(
        n14804) );
  OAI21_X1 U16483 ( .B1(n14845), .B2(n14805), .A(n14804), .ZN(n14806) );
  INV_X1 U16484 ( .A(n14806), .ZN(n14810) );
  AOI22_X1 U16485 ( .A1(n14808), .A2(n14851), .B1(n14849), .B2(n14807), .ZN(
        n14809) );
  OAI211_X1 U16486 ( .C1(n14842), .C2(n14811), .A(n14810), .B(n14809), .ZN(
        P1_U3287) );
  INV_X1 U16487 ( .A(n14812), .ZN(n14821) );
  NAND2_X1 U16488 ( .A1(n14814), .A2(n14813), .ZN(n14817) );
  AOI22_X1 U16489 ( .A1(n14842), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n14815), 
        .B2(n14841), .ZN(n14816) );
  OAI211_X1 U16490 ( .C1(n14819), .C2(n14818), .A(n14817), .B(n14816), .ZN(
        n14820) );
  AOI21_X1 U16491 ( .B1(n14821), .B2(n14851), .A(n14820), .ZN(n14822) );
  OAI21_X1 U16492 ( .B1(n14842), .B2(n14823), .A(n14822), .ZN(P1_U3288) );
  XNOR2_X1 U16493 ( .A(n14824), .B(n14825), .ZN(n14865) );
  XNOR2_X1 U16494 ( .A(n14826), .B(n14825), .ZN(n14827) );
  NOR2_X1 U16495 ( .A1(n14827), .A2(n14885), .ZN(n14828) );
  AOI211_X1 U16496 ( .C1(n14877), .C2(n14865), .A(n14829), .B(n14828), .ZN(
        n14862) );
  NOR2_X1 U16497 ( .A1(n14831), .A2(n14830), .ZN(n14832) );
  AOI21_X1 U16498 ( .B1(n14842), .B2(P1_REG2_REG_2__SCAN_IN), .A(n14832), .ZN(
        n14833) );
  OAI21_X1 U16499 ( .B1(n14845), .B2(n14861), .A(n14833), .ZN(n14834) );
  INV_X1 U16500 ( .A(n14834), .ZN(n14840) );
  OAI211_X1 U16501 ( .C1(n6828), .C2(n14861), .A(n14837), .B(n14836), .ZN(
        n14860) );
  INV_X1 U16502 ( .A(n14860), .ZN(n14838) );
  AOI22_X1 U16503 ( .A1(n14851), .A2(n14865), .B1(n14849), .B2(n14838), .ZN(
        n14839) );
  OAI211_X1 U16504 ( .C1(n14842), .C2(n14862), .A(n14840), .B(n14839), .ZN(
        P1_U3291) );
  AOI22_X1 U16505 ( .A1(n14842), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n14841), .ZN(n14843) );
  OAI21_X1 U16506 ( .B1(n14845), .B2(n14844), .A(n14843), .ZN(n14846) );
  INV_X1 U16507 ( .A(n14846), .ZN(n14853) );
  INV_X1 U16508 ( .A(n14847), .ZN(n14848) );
  AOI22_X1 U16509 ( .A1(n14851), .A2(n14850), .B1(n14849), .B2(n14848), .ZN(
        n14852) );
  OAI211_X1 U16510 ( .C1(n14842), .C2(n14854), .A(n14853), .B(n14852), .ZN(
        P1_U3292) );
  AND2_X1 U16511 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14855), .ZN(P1_U3294) );
  AND2_X1 U16512 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14855), .ZN(P1_U3295) );
  AND2_X1 U16513 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14855), .ZN(P1_U3296) );
  AND2_X1 U16514 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14855), .ZN(P1_U3297) );
  AND2_X1 U16515 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14855), .ZN(P1_U3298) );
  AND2_X1 U16516 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14855), .ZN(P1_U3299) );
  AND2_X1 U16517 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14855), .ZN(P1_U3300) );
  AND2_X1 U16518 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14855), .ZN(P1_U3301) );
  AND2_X1 U16519 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14855), .ZN(P1_U3302) );
  AND2_X1 U16520 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14855), .ZN(P1_U3303) );
  AND2_X1 U16521 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14855), .ZN(P1_U3304) );
  AND2_X1 U16522 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14855), .ZN(P1_U3305) );
  AND2_X1 U16523 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14855), .ZN(P1_U3306) );
  AND2_X1 U16524 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14855), .ZN(P1_U3307) );
  AND2_X1 U16525 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14855), .ZN(P1_U3308) );
  AND2_X1 U16526 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14855), .ZN(P1_U3309) );
  AND2_X1 U16527 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14855), .ZN(P1_U3310) );
  AND2_X1 U16528 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14855), .ZN(P1_U3311) );
  AND2_X1 U16529 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14855), .ZN(P1_U3312) );
  AND2_X1 U16530 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14855), .ZN(P1_U3313) );
  AND2_X1 U16531 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14855), .ZN(P1_U3314) );
  AND2_X1 U16532 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14855), .ZN(P1_U3315) );
  AND2_X1 U16533 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14855), .ZN(P1_U3316) );
  AND2_X1 U16534 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14855), .ZN(P1_U3317) );
  AND2_X1 U16535 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14855), .ZN(P1_U3318) );
  AND2_X1 U16536 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14855), .ZN(P1_U3319) );
  AND2_X1 U16537 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14855), .ZN(P1_U3320) );
  AND2_X1 U16538 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14855), .ZN(P1_U3321) );
  AND2_X1 U16539 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14855), .ZN(P1_U3322) );
  AND2_X1 U16540 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14855), .ZN(P1_U3323) );
  INV_X1 U16541 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n14856) );
  AOI22_X1 U16542 ( .A1(n14891), .A2(n14857), .B1(n14856), .B2(n14889), .ZN(
        P1_U3459) );
  INV_X1 U16543 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14858) );
  AOI22_X1 U16544 ( .A1(n14891), .A2(n14859), .B1(n14858), .B2(n14889), .ZN(
        P1_U3462) );
  OAI21_X1 U16545 ( .B1(n14861), .B2(n14872), .A(n14860), .ZN(n14864) );
  INV_X1 U16546 ( .A(n14862), .ZN(n14863) );
  AOI211_X1 U16547 ( .C1(n14866), .C2(n14865), .A(n14864), .B(n14863), .ZN(
        n14892) );
  INV_X1 U16548 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n14867) );
  AOI22_X1 U16549 ( .A1(n14891), .A2(n14892), .B1(n14867), .B2(n14889), .ZN(
        P1_U3465) );
  INV_X1 U16550 ( .A(n14869), .ZN(n14876) );
  NOR2_X1 U16551 ( .A1(n14869), .A2(n14868), .ZN(n14875) );
  OAI211_X1 U16552 ( .C1(n14873), .C2(n14872), .A(n14871), .B(n14870), .ZN(
        n14874) );
  AOI211_X1 U16553 ( .C1(n14877), .C2(n14876), .A(n14875), .B(n14874), .ZN(
        n14893) );
  INV_X1 U16554 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14878) );
  AOI22_X1 U16555 ( .A1(n14891), .A2(n14893), .B1(n14878), .B2(n14889), .ZN(
        P1_U3468) );
  AOI211_X1 U16556 ( .C1(n14882), .C2(n14881), .A(n14880), .B(n14879), .ZN(
        n14883) );
  OAI21_X1 U16557 ( .B1(n14885), .B2(n14884), .A(n14883), .ZN(n14886) );
  AOI21_X1 U16558 ( .B1(n14888), .B2(n14887), .A(n14886), .ZN(n14895) );
  INV_X1 U16559 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14890) );
  AOI22_X1 U16560 ( .A1(n14891), .A2(n14895), .B1(n14890), .B2(n14889), .ZN(
        P1_U3471) );
  AOI22_X1 U16561 ( .A1(n14896), .A2(n14892), .B1(n10076), .B2(n14894), .ZN(
        P1_U3530) );
  AOI22_X1 U16562 ( .A1(n14896), .A2(n14893), .B1(n10077), .B2(n14894), .ZN(
        P1_U3531) );
  AOI22_X1 U16563 ( .A1(n14896), .A2(n14895), .B1(n10078), .B2(n14894), .ZN(
        P1_U3532) );
  NOR2_X1 U16564 ( .A1(n14920), .A2(P2_U3947), .ZN(P2_U3087) );
  NAND2_X1 U16565 ( .A1(n9782), .A2(n10457), .ZN(n14897) );
  NAND2_X1 U16566 ( .A1(n14897), .A2(n15067), .ZN(n14898) );
  NAND2_X1 U16567 ( .A1(n14899), .A2(n14898), .ZN(n14902) );
  NAND2_X1 U16568 ( .A1(n14916), .A2(n15089), .ZN(n14901) );
  AND2_X1 U16569 ( .A1(n9833), .A2(n13198), .ZN(n15063) );
  NAND2_X1 U16570 ( .A1(n14914), .A2(n15063), .ZN(n14900) );
  OAI211_X1 U16571 ( .C1(n14903), .C2(n14902), .A(n14901), .B(n14900), .ZN(
        n14904) );
  INV_X1 U16572 ( .A(n14904), .ZN(n14905) );
  OAI21_X1 U16573 ( .B1(n14919), .B2(n15069), .A(n14905), .ZN(P2_U3204) );
  INV_X1 U16574 ( .A(n14906), .ZN(n14908) );
  NAND3_X1 U16575 ( .A1(n14909), .A2(n14908), .A3(n14907), .ZN(n14910) );
  NAND2_X1 U16576 ( .A1(n14911), .A2(n14910), .ZN(n14913) );
  AOI222_X1 U16577 ( .A1(n14916), .A2(n9785), .B1(n14915), .B2(n14914), .C1(
        n14913), .C2(n14912), .ZN(n14917) );
  OAI21_X1 U16578 ( .B1(n14919), .B2(n14918), .A(n14917), .ZN(P2_U3209) );
  AOI22_X1 U16579 ( .A1(n14920), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n14932) );
  OAI211_X1 U16580 ( .C1(n14923), .C2(n14922), .A(n15035), .B(n14921), .ZN(
        n14928) );
  OAI211_X1 U16581 ( .C1(n14926), .C2(n14925), .A(n15043), .B(n14924), .ZN(
        n14927) );
  OAI211_X1 U16582 ( .C1(n15037), .C2(n14929), .A(n14928), .B(n14927), .ZN(
        n14930) );
  INV_X1 U16583 ( .A(n14930), .ZN(n14931) );
  NAND2_X1 U16584 ( .A1(n14932), .A2(n14931), .ZN(P2_U3216) );
  INV_X1 U16585 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14945) );
  OAI211_X1 U16586 ( .C1(n14935), .C2(n14934), .A(n15035), .B(n14933), .ZN(
        n14940) );
  OAI211_X1 U16587 ( .C1(n14938), .C2(n14937), .A(n15043), .B(n14936), .ZN(
        n14939) );
  OAI211_X1 U16588 ( .C1(n15037), .C2(n14941), .A(n14940), .B(n14939), .ZN(
        n14942) );
  INV_X1 U16589 ( .A(n14942), .ZN(n14944) );
  OAI211_X1 U16590 ( .C1(n14945), .C2(n15046), .A(n14944), .B(n14943), .ZN(
        P2_U3222) );
  OAI21_X1 U16591 ( .B1(n14947), .B2(n14946), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n14948) );
  OAI21_X1 U16592 ( .B1(P2_STATE_REG_SCAN_IN), .B2(P2_REG3_REG_9__SCAN_IN), 
        .A(n14948), .ZN(n14961) );
  INV_X1 U16593 ( .A(n14949), .ZN(n14950) );
  AOI21_X1 U16594 ( .B1(n14952), .B2(n14951), .A(n14950), .ZN(n14958) );
  INV_X1 U16595 ( .A(n14953), .ZN(n14954) );
  AOI21_X1 U16596 ( .B1(n14956), .B2(n14955), .A(n14954), .ZN(n14957) );
  OAI22_X1 U16597 ( .A1(n15008), .A2(n14958), .B1(n14957), .B2(n15022), .ZN(
        n14959) );
  INV_X1 U16598 ( .A(n14959), .ZN(n14960) );
  OAI211_X1 U16599 ( .C1(n14962), .C2(n15046), .A(n14961), .B(n14960), .ZN(
        P2_U3223) );
  INV_X1 U16600 ( .A(n14963), .ZN(n14964) );
  AOI211_X1 U16601 ( .C1(n14966), .C2(n14965), .A(n15022), .B(n14964), .ZN(
        n14972) );
  INV_X1 U16602 ( .A(n14967), .ZN(n14968) );
  AOI211_X1 U16603 ( .C1(n14970), .C2(n14969), .A(n14968), .B(n15008), .ZN(
        n14971) );
  AOI211_X1 U16604 ( .C1(n15028), .C2(n14973), .A(n14972), .B(n14971), .ZN(
        n14975) );
  NAND2_X1 U16605 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n14974)
         );
  OAI211_X1 U16606 ( .C1(n14976), .C2(n15046), .A(n14975), .B(n14974), .ZN(
        P2_U3224) );
  NAND2_X1 U16607 ( .A1(n14978), .A2(n14977), .ZN(n14979) );
  NAND2_X1 U16608 ( .A1(n14980), .A2(n14979), .ZN(n14983) );
  NOR2_X1 U16609 ( .A1(n15037), .A2(n14981), .ZN(n14982) );
  AOI21_X1 U16610 ( .B1(n14983), .B2(n15035), .A(n14982), .ZN(n14988) );
  XNOR2_X1 U16611 ( .A(n14985), .B(n14984), .ZN(n14986) );
  NAND2_X1 U16612 ( .A1(n14986), .A2(n15043), .ZN(n14987) );
  AND2_X1 U16613 ( .A1(n14988), .A2(n14987), .ZN(n14990) );
  OAI211_X1 U16614 ( .C1(n15387), .C2(n15046), .A(n14990), .B(n14989), .ZN(
        P2_U3226) );
  AOI211_X1 U16615 ( .C1(n14993), .C2(n14992), .A(n14991), .B(n15008), .ZN(
        n14998) );
  AOI211_X1 U16616 ( .C1(n14996), .C2(n14995), .A(n14994), .B(n15022), .ZN(
        n14997) );
  AOI211_X1 U16617 ( .C1(n15028), .C2(n14999), .A(n14998), .B(n14997), .ZN(
        n15001) );
  NAND2_X1 U16618 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n15000)
         );
  OAI211_X1 U16619 ( .C1(n15002), .C2(n15046), .A(n15001), .B(n15000), .ZN(
        P2_U3229) );
  AOI211_X1 U16620 ( .C1(n15005), .C2(n15004), .A(n15022), .B(n15003), .ZN(
        n15012) );
  INV_X1 U16621 ( .A(n15006), .ZN(n15007) );
  AOI211_X1 U16622 ( .C1(n15010), .C2(n15009), .A(n15008), .B(n15007), .ZN(
        n15011) );
  AOI211_X1 U16623 ( .C1(n15028), .C2(n15013), .A(n15012), .B(n15011), .ZN(
        n15015) );
  OAI211_X1 U16624 ( .C1(n15016), .C2(n15046), .A(n15015), .B(n15014), .ZN(
        P2_U3230) );
  OAI211_X1 U16625 ( .C1(n15019), .C2(n15018), .A(n15017), .B(n15043), .ZN(
        n15020) );
  INV_X1 U16626 ( .A(n15020), .ZN(n15026) );
  AOI211_X1 U16627 ( .C1(n15024), .C2(n15023), .A(n15022), .B(n15021), .ZN(
        n15025) );
  AOI211_X1 U16628 ( .C1(n15028), .C2(n15027), .A(n15026), .B(n15025), .ZN(
        n15030) );
  OAI211_X1 U16629 ( .C1(n15031), .C2(n15046), .A(n15030), .B(n15029), .ZN(
        P2_U3231) );
  INV_X1 U16630 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n15047) );
  OAI21_X1 U16631 ( .B1(n15034), .B2(n15033), .A(n15032), .ZN(n15042) );
  OAI21_X1 U16632 ( .B1(n15036), .B2(P2_REG1_REG_18__SCAN_IN), .A(n15035), 
        .ZN(n15040) );
  OAI22_X1 U16633 ( .A1(n15040), .A2(n15039), .B1(n15038), .B2(n15037), .ZN(
        n15041) );
  AOI21_X1 U16634 ( .B1(n15043), .B2(n15042), .A(n15041), .ZN(n15045) );
  OAI211_X1 U16635 ( .C1(n15047), .C2(n15046), .A(n15045), .B(n15044), .ZN(
        P2_U3232) );
  INV_X1 U16636 ( .A(n15048), .ZN(n15056) );
  NAND2_X1 U16637 ( .A1(n15050), .A2(n15049), .ZN(n15054) );
  AOI22_X1 U16638 ( .A1(n15076), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n15052), 
        .B2(n15051), .ZN(n15053) );
  OAI211_X1 U16639 ( .C1(n15056), .C2(n15055), .A(n15054), .B(n15053), .ZN(
        n15057) );
  AOI21_X1 U16640 ( .B1(n15059), .B2(n15058), .A(n15057), .ZN(n15060) );
  OAI21_X1 U16641 ( .B1(n15076), .B2(n15061), .A(n15060), .ZN(P2_U3258) );
  NAND2_X1 U16642 ( .A1(n10200), .A2(n15127), .ZN(n15062) );
  NAND2_X1 U16643 ( .A1(n15072), .A2(n15062), .ZN(n15065) );
  INV_X1 U16644 ( .A(n15063), .ZN(n15064) );
  NAND2_X1 U16645 ( .A1(n15065), .A2(n15064), .ZN(n15088) );
  AND2_X1 U16646 ( .A1(n10457), .A2(n15066), .ZN(n15068) );
  OAI22_X1 U16647 ( .A1(n15070), .A2(n15069), .B1(n15068), .B2(n15067), .ZN(
        n15071) );
  NOR2_X1 U16648 ( .A1(n15088), .A2(n15071), .ZN(n15075) );
  AOI22_X1 U16649 ( .A1(n15073), .A2(n15072), .B1(P2_REG2_REG_0__SCAN_IN), 
        .B2(n15076), .ZN(n15074) );
  OAI21_X1 U16650 ( .B1(n15076), .B2(n15075), .A(n15074), .ZN(P2_U3265) );
  INV_X1 U16651 ( .A(n15077), .ZN(n15078) );
  AND2_X1 U16652 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15080), .ZN(P2_U3266) );
  INV_X1 U16653 ( .A(n15080), .ZN(n15079) );
  INV_X1 U16654 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15323) );
  NOR2_X1 U16655 ( .A1(n15079), .A2(n15323), .ZN(P2_U3267) );
  INV_X1 U16656 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15281) );
  NOR2_X1 U16657 ( .A1(n15079), .A2(n15281), .ZN(P2_U3268) );
  AND2_X1 U16658 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15080), .ZN(P2_U3269) );
  AND2_X1 U16659 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15080), .ZN(P2_U3270) );
  INV_X1 U16660 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n15421) );
  NOR2_X1 U16661 ( .A1(n15079), .A2(n15421), .ZN(P2_U3271) );
  AND2_X1 U16662 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15080), .ZN(P2_U3272) );
  AND2_X1 U16663 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15080), .ZN(P2_U3273) );
  AND2_X1 U16664 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15080), .ZN(P2_U3274) );
  AND2_X1 U16665 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15080), .ZN(P2_U3275) );
  AND2_X1 U16666 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15080), .ZN(P2_U3276) );
  AND2_X1 U16667 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15080), .ZN(P2_U3277) );
  AND2_X1 U16668 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15080), .ZN(P2_U3278) );
  AND2_X1 U16669 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15080), .ZN(P2_U3279) );
  AND2_X1 U16670 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15080), .ZN(P2_U3280) );
  AND2_X1 U16671 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15080), .ZN(P2_U3281) );
  AND2_X1 U16672 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15080), .ZN(P2_U3282) );
  AND2_X1 U16673 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15080), .ZN(P2_U3283) );
  AND2_X1 U16674 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15080), .ZN(P2_U3284) );
  AND2_X1 U16675 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15080), .ZN(P2_U3285) );
  AND2_X1 U16676 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15080), .ZN(P2_U3286) );
  AND2_X1 U16677 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15080), .ZN(P2_U3287) );
  AND2_X1 U16678 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15080), .ZN(P2_U3288) );
  AND2_X1 U16679 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15080), .ZN(P2_U3289) );
  AND2_X1 U16680 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15080), .ZN(P2_U3290) );
  INV_X1 U16681 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15322) );
  NOR2_X1 U16682 ( .A1(n15079), .A2(n15322), .ZN(P2_U3291) );
  AND2_X1 U16683 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15080), .ZN(P2_U3292) );
  AND2_X1 U16684 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15080), .ZN(P2_U3293) );
  AND2_X1 U16685 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15080), .ZN(P2_U3294) );
  AND2_X1 U16686 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15080), .ZN(P2_U3295) );
  AOI22_X1 U16687 ( .A1(n15082), .A2(n15081), .B1(n9862), .B2(n15084), .ZN(
        P2_U3416) );
  AOI21_X1 U16688 ( .B1(P2_D_REG_1__SCAN_IN), .B2(n15084), .A(n15083), .ZN(
        n15085) );
  INV_X1 U16689 ( .A(n15085), .ZN(P2_U3417) );
  NOR2_X1 U16690 ( .A1(n15086), .A2(n15107), .ZN(n15087) );
  AOI211_X1 U16691 ( .C1(n15090), .C2(n15089), .A(n15088), .B(n15087), .ZN(
        n15136) );
  INV_X1 U16692 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15091) );
  AOI22_X1 U16693 ( .A1(n15134), .A2(n15136), .B1(n15091), .B2(n15132), .ZN(
        P2_U3430) );
  INV_X1 U16694 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n15092) );
  AOI22_X1 U16695 ( .A1(n15134), .A2(n15093), .B1(n15092), .B2(n15132), .ZN(
        P2_U3433) );
  INV_X1 U16696 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15094) );
  AOI22_X1 U16697 ( .A1(n15134), .A2(n15095), .B1(n15094), .B2(n15132), .ZN(
        P2_U3436) );
  INV_X1 U16698 ( .A(n15096), .ZN(n15102) );
  NOR2_X1 U16699 ( .A1(n15096), .A2(n15107), .ZN(n15101) );
  OAI211_X1 U16700 ( .C1(n15099), .C2(n15114), .A(n15098), .B(n15097), .ZN(
        n15100) );
  AOI211_X1 U16701 ( .C1(n15102), .C2(n15131), .A(n15101), .B(n15100), .ZN(
        n15138) );
  INV_X1 U16702 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15103) );
  AOI22_X1 U16703 ( .A1(n15134), .A2(n15138), .B1(n15103), .B2(n15132), .ZN(
        P2_U3442) );
  INV_X1 U16704 ( .A(n15108), .ZN(n15111) );
  AOI21_X1 U16705 ( .B1(n15123), .B2(n15105), .A(n15104), .ZN(n15106) );
  OAI21_X1 U16706 ( .B1(n15108), .B2(n15107), .A(n15106), .ZN(n15109) );
  AOI211_X1 U16707 ( .C1(n15131), .C2(n15111), .A(n15110), .B(n15109), .ZN(
        n15139) );
  INV_X1 U16708 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15112) );
  AOI22_X1 U16709 ( .A1(n15134), .A2(n15139), .B1(n15112), .B2(n15132), .ZN(
        P2_U3445) );
  OAI21_X1 U16710 ( .B1(n15115), .B2(n15114), .A(n15113), .ZN(n15117) );
  AOI211_X1 U16711 ( .C1(n15124), .C2(n15118), .A(n15117), .B(n15116), .ZN(
        n15141) );
  INV_X1 U16712 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15119) );
  AOI22_X1 U16713 ( .A1(n15134), .A2(n15141), .B1(n15119), .B2(n15132), .ZN(
        P2_U3454) );
  AOI211_X1 U16714 ( .C1(n15123), .C2(n15122), .A(n15121), .B(n15120), .ZN(
        n15126) );
  NAND2_X1 U16715 ( .A1(n15130), .A2(n15124), .ZN(n15125) );
  OAI211_X1 U16716 ( .C1(n15128), .C2(n15127), .A(n15126), .B(n15125), .ZN(
        n15129) );
  AOI21_X1 U16717 ( .B1(n15131), .B2(n15130), .A(n15129), .ZN(n15144) );
  INV_X1 U16718 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n15133) );
  AOI22_X1 U16719 ( .A1(n15134), .A2(n15144), .B1(n15133), .B2(n15132), .ZN(
        P2_U3463) );
  AOI22_X1 U16720 ( .A1(n15145), .A2(n15136), .B1(n15135), .B2(n15142), .ZN(
        P2_U3499) );
  INV_X1 U16721 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n15137) );
  AOI22_X1 U16722 ( .A1(n15145), .A2(n15138), .B1(n15137), .B2(n15142), .ZN(
        P2_U3503) );
  AOI22_X1 U16723 ( .A1(n15145), .A2(n15139), .B1(n10014), .B2(n15142), .ZN(
        P2_U3504) );
  AOI22_X1 U16724 ( .A1(n15145), .A2(n15141), .B1(n15140), .B2(n15142), .ZN(
        P2_U3507) );
  AOI22_X1 U16725 ( .A1(n15145), .A2(n15144), .B1(n15143), .B2(n15142), .ZN(
        P2_U3510) );
  NOR2_X1 U16726 ( .A1(P3_U3897), .A2(n15168), .ZN(P3_U3150) );
  OAI22_X1 U16727 ( .A1(n15147), .A2(n7522), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15146), .ZN(n15148) );
  INV_X1 U16728 ( .A(n15148), .ZN(n15155) );
  NOR2_X1 U16729 ( .A1(n15149), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15152) );
  NAND3_X1 U16730 ( .A1(n15164), .A2(n15162), .A3(n15150), .ZN(n15151) );
  OAI21_X1 U16731 ( .B1(n15153), .B2(n15152), .A(n15151), .ZN(n15154) );
  OAI211_X1 U16732 ( .C1(n15157), .C2(n15156), .A(n15155), .B(n15154), .ZN(
        P3_U3182) );
  AOI21_X1 U16733 ( .B1(n15159), .B2(n11401), .A(n15158), .ZN(n15165) );
  AOI21_X1 U16734 ( .B1(n15161), .B2(n11402), .A(n15160), .ZN(n15163) );
  OAI22_X1 U16735 ( .A1(n15165), .A2(n15164), .B1(n15163), .B2(n15162), .ZN(
        n15166) );
  AOI211_X1 U16736 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n15168), .A(n15167), .B(
        n15166), .ZN(n15177) );
  OAI21_X1 U16737 ( .B1(n15171), .B2(n15170), .A(n15169), .ZN(n15172) );
  AOI22_X1 U16738 ( .A1(n15175), .A2(n15174), .B1(n15173), .B2(n15172), .ZN(
        n15176) );
  NAND2_X1 U16739 ( .A1(n15177), .A2(n15176), .ZN(P3_U3191) );
  XNOR2_X1 U16740 ( .A(n15178), .B(n15180), .ZN(n15186) );
  OAI21_X1 U16741 ( .B1(n15181), .B2(n15180), .A(n15179), .ZN(n15187) );
  OAI22_X1 U16742 ( .A1(n7815), .A2(n15183), .B1(n6969), .B2(n15182), .ZN(
        n15184) );
  AOI21_X1 U16743 ( .B1(n15187), .B2(n15199), .A(n15184), .ZN(n15185) );
  OAI21_X1 U16744 ( .B1(n15206), .B2(n15186), .A(n15185), .ZN(n15219) );
  INV_X1 U16745 ( .A(n15187), .ZN(n15223) );
  NAND2_X1 U16746 ( .A1(n15189), .A2(n15188), .ZN(n15220) );
  OAI22_X1 U16747 ( .A1(n15223), .A2(n15191), .B1(n15190), .B2(n15220), .ZN(
        n15192) );
  AOI211_X1 U16748 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15209), .A(n15219), .B(
        n15192), .ZN(n15193) );
  AOI22_X1 U16749 ( .A1(n15194), .A2(n10405), .B1(n15193), .B2(n12718), .ZN(
        P3_U3231) );
  NOR2_X1 U16750 ( .A1(n15196), .A2(n15195), .ZN(n15216) );
  XNOR2_X1 U16751 ( .A(n8482), .B(n15197), .ZN(n15207) );
  XNOR2_X1 U16752 ( .A(n8482), .B(n15198), .ZN(n15217) );
  NAND2_X1 U16753 ( .A1(n15217), .A2(n15199), .ZN(n15205) );
  AOI22_X1 U16754 ( .A1(n15203), .A2(n15202), .B1(n15201), .B2(n15200), .ZN(
        n15204) );
  OAI211_X1 U16755 ( .C1(n15207), .C2(n15206), .A(n15205), .B(n15204), .ZN(
        n15215) );
  AOI21_X1 U16756 ( .B1(n15216), .B2(n15208), .A(n15215), .ZN(n15213) );
  AOI22_X1 U16757 ( .A1(n15210), .A2(n15217), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15209), .ZN(n15211) );
  OAI221_X1 U16758 ( .B1(n15214), .B2(n15213), .C1(n12749), .C2(n15212), .A(
        n15211), .ZN(P3_U3232) );
  AOI211_X1 U16759 ( .C1(n15242), .C2(n15217), .A(n15216), .B(n15215), .ZN(
        n15247) );
  INV_X1 U16760 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15218) );
  AOI22_X1 U16761 ( .A1(n15246), .A2(n15247), .B1(n15218), .B2(n15244), .ZN(
        P3_U3393) );
  INV_X1 U16762 ( .A(n15219), .ZN(n15221) );
  OAI211_X1 U16763 ( .C1(n15223), .C2(n15222), .A(n15221), .B(n15220), .ZN(
        n15248) );
  OAI22_X1 U16764 ( .A1(n15244), .A2(n15248), .B1(P3_REG0_REG_2__SCAN_IN), 
        .B2(n15246), .ZN(n15224) );
  INV_X1 U16765 ( .A(n15224), .ZN(P3_U3396) );
  INV_X1 U16766 ( .A(n15225), .ZN(n15227) );
  AOI211_X1 U16767 ( .C1(n15228), .C2(n15242), .A(n15227), .B(n15226), .ZN(
        n15250) );
  INV_X1 U16768 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15229) );
  AOI22_X1 U16769 ( .A1(n15246), .A2(n15250), .B1(n15229), .B2(n15244), .ZN(
        P3_U3405) );
  AOI211_X1 U16770 ( .C1(n15232), .C2(n15242), .A(n15231), .B(n15230), .ZN(
        n15251) );
  INV_X1 U16771 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15233) );
  AOI22_X1 U16772 ( .A1(n15246), .A2(n15251), .B1(n15233), .B2(n15244), .ZN(
        P3_U3414) );
  INV_X1 U16773 ( .A(n15234), .ZN(n15237) );
  AOI211_X1 U16774 ( .C1(n15237), .C2(n15242), .A(n15236), .B(n15235), .ZN(
        n15252) );
  INV_X1 U16775 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15238) );
  AOI22_X1 U16776 ( .A1(n15246), .A2(n15252), .B1(n15238), .B2(n15244), .ZN(
        P3_U3417) );
  INV_X1 U16777 ( .A(n15239), .ZN(n15243) );
  AOI211_X1 U16778 ( .C1(n15243), .C2(n15242), .A(n15241), .B(n15240), .ZN(
        n15253) );
  INV_X1 U16779 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15245) );
  AOI22_X1 U16780 ( .A1(n15246), .A2(n15253), .B1(n15245), .B2(n15244), .ZN(
        P3_U3420) );
  AOI22_X1 U16781 ( .A1(n15254), .A2(n15247), .B1(n10378), .B2(n12766), .ZN(
        P3_U3460) );
  OAI22_X1 U16782 ( .A1(n12766), .A2(n15248), .B1(P3_REG1_REG_2__SCAN_IN), 
        .B2(n15254), .ZN(n15249) );
  INV_X1 U16783 ( .A(n15249), .ZN(P3_U3461) );
  AOI22_X1 U16784 ( .A1(n15254), .A2(n15250), .B1(n7866), .B2(n12766), .ZN(
        P3_U3464) );
  AOI22_X1 U16785 ( .A1(n15254), .A2(n15251), .B1(n7919), .B2(n12766), .ZN(
        P3_U3467) );
  AOI22_X1 U16786 ( .A1(n15254), .A2(n15252), .B1(n11401), .B2(n12766), .ZN(
        P3_U3468) );
  AOI22_X1 U16787 ( .A1(n15254), .A2(n15253), .B1(n7955), .B2(n12766), .ZN(
        P3_U3469) );
  AOI22_X1 U16788 ( .A1(n15429), .A2(keyinput92), .B1(keyinput110), .B2(n15256), .ZN(n15255) );
  OAI221_X1 U16789 ( .B1(n15429), .B2(keyinput92), .C1(n15256), .C2(
        keyinput110), .A(n15255), .ZN(n15267) );
  INV_X1 U16790 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n15258) );
  AOI22_X1 U16791 ( .A1(n15259), .A2(keyinput99), .B1(keyinput84), .B2(n15258), 
        .ZN(n15257) );
  OAI221_X1 U16792 ( .B1(n15259), .B2(keyinput99), .C1(n15258), .C2(keyinput84), .A(n15257), .ZN(n15266) );
  AOI22_X1 U16793 ( .A1(n15261), .A2(keyinput118), .B1(keyinput87), .B2(n14179), .ZN(n15260) );
  OAI221_X1 U16794 ( .B1(n15261), .B2(keyinput118), .C1(n14179), .C2(
        keyinput87), .A(n15260), .ZN(n15265) );
  XOR2_X1 U16795 ( .A(n7898), .B(keyinput81), .Z(n15263) );
  XNOR2_X1 U16796 ( .A(P3_IR_REG_16__SCAN_IN), .B(keyinput103), .ZN(n15262) );
  NAND2_X1 U16797 ( .A1(n15263), .A2(n15262), .ZN(n15264) );
  NOR4_X1 U16798 ( .A1(n15267), .A2(n15266), .A3(n15265), .A4(n15264), .ZN(
        n15304) );
  INV_X1 U16799 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n15383) );
  AOI22_X1 U16800 ( .A1(n15383), .A2(keyinput71), .B1(keyinput89), .B2(n11034), 
        .ZN(n15268) );
  OAI221_X1 U16801 ( .B1(n15383), .B2(keyinput71), .C1(n11034), .C2(keyinput89), .A(n15268), .ZN(n15276) );
  AOI22_X1 U16802 ( .A1(n7786), .A2(keyinput127), .B1(keyinput112), .B2(n15421), .ZN(n15269) );
  OAI221_X1 U16803 ( .B1(n7786), .B2(keyinput127), .C1(n15421), .C2(
        keyinput112), .A(n15269), .ZN(n15275) );
  AOI22_X1 U16804 ( .A1(n15401), .A2(keyinput108), .B1(keyinput114), .B2(n7784), .ZN(n15270) );
  OAI221_X1 U16805 ( .B1(n15401), .B2(keyinput108), .C1(n7784), .C2(
        keyinput114), .A(n15270), .ZN(n15274) );
  AOI22_X1 U16806 ( .A1(n15272), .A2(keyinput86), .B1(keyinput121), .B2(n12673), .ZN(n15271) );
  OAI221_X1 U16807 ( .B1(n15272), .B2(keyinput86), .C1(n12673), .C2(
        keyinput121), .A(n15271), .ZN(n15273) );
  NOR4_X1 U16808 ( .A1(n15276), .A2(n15275), .A3(n15274), .A4(n15273), .ZN(
        n15303) );
  AOI22_X1 U16809 ( .A1(n15399), .A2(keyinput113), .B1(n11824), .B2(
        keyinput123), .ZN(n15277) );
  OAI221_X1 U16810 ( .B1(n15399), .B2(keyinput113), .C1(n11824), .C2(
        keyinput123), .A(n15277), .ZN(n15287) );
  INV_X1 U16811 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n15384) );
  AOI22_X1 U16812 ( .A1(n15384), .A2(keyinput67), .B1(n15389), .B2(keyinput94), 
        .ZN(n15278) );
  OAI221_X1 U16813 ( .B1(n15384), .B2(keyinput67), .C1(n15389), .C2(keyinput94), .A(n15278), .ZN(n15286) );
  AOI22_X1 U16814 ( .A1(n15281), .A2(keyinput77), .B1(n15280), .B2(keyinput106), .ZN(n15279) );
  OAI221_X1 U16815 ( .B1(n15281), .B2(keyinput77), .C1(n15280), .C2(
        keyinput106), .A(n15279), .ZN(n15285) );
  AOI22_X1 U16816 ( .A1(n15283), .A2(keyinput74), .B1(keyinput107), .B2(n15390), .ZN(n15282) );
  OAI221_X1 U16817 ( .B1(n15283), .B2(keyinput74), .C1(n15390), .C2(
        keyinput107), .A(n15282), .ZN(n15284) );
  NOR4_X1 U16818 ( .A1(n15287), .A2(n15286), .A3(n15285), .A4(n15284), .ZN(
        n15302) );
  INV_X1 U16819 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n15289) );
  AOI22_X1 U16820 ( .A1(n11155), .A2(keyinput69), .B1(keyinput91), .B2(n15289), 
        .ZN(n15288) );
  OAI221_X1 U16821 ( .B1(n11155), .B2(keyinput69), .C1(n15289), .C2(keyinput91), .A(n15288), .ZN(n15293) );
  XOR2_X1 U16822 ( .A(P3_IR_REG_5__SCAN_IN), .B(keyinput83), .Z(n15292) );
  XNOR2_X1 U16823 ( .A(n15290), .B(keyinput122), .ZN(n15291) );
  OR3_X1 U16824 ( .A1(n15293), .A2(n15292), .A3(n15291), .ZN(n15300) );
  AOI22_X1 U16825 ( .A1(n15387), .A2(keyinput70), .B1(n10158), .B2(keyinput115), .ZN(n15294) );
  OAI221_X1 U16826 ( .B1(n15387), .B2(keyinput70), .C1(n10158), .C2(
        keyinput115), .A(n15294), .ZN(n15299) );
  INV_X1 U16827 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n15297) );
  INV_X1 U16828 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n15296) );
  AOI22_X1 U16829 ( .A1(n15297), .A2(keyinput120), .B1(keyinput124), .B2(
        n15296), .ZN(n15295) );
  OAI221_X1 U16830 ( .B1(n15297), .B2(keyinput120), .C1(n15296), .C2(
        keyinput124), .A(n15295), .ZN(n15298) );
  NOR3_X1 U16831 ( .A1(n15300), .A2(n15299), .A3(n15298), .ZN(n15301) );
  AND4_X1 U16832 ( .A1(n15304), .A2(n15303), .A3(n15302), .A4(n15301), .ZN(
        n15440) );
  OAI22_X1 U16833 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(keyinput75), .B1(
        keyinput90), .B2(P2_IR_REG_21__SCAN_IN), .ZN(n15305) );
  AOI221_X1 U16834 ( .B1(P3_REG1_REG_6__SCAN_IN), .B2(keyinput75), .C1(
        P2_IR_REG_21__SCAN_IN), .C2(keyinput90), .A(n15305), .ZN(n15312) );
  OAI22_X1 U16835 ( .A1(P3_REG3_REG_15__SCAN_IN), .A2(keyinput66), .B1(
        P2_REG2_REG_29__SCAN_IN), .B2(keyinput117), .ZN(n15306) );
  AOI221_X1 U16836 ( .B1(P3_REG3_REG_15__SCAN_IN), .B2(keyinput66), .C1(
        keyinput117), .C2(P2_REG2_REG_29__SCAN_IN), .A(n15306), .ZN(n15311) );
  OAI22_X1 U16837 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(keyinput125), .B1(
        P2_REG0_REG_11__SCAN_IN), .B2(keyinput116), .ZN(n15307) );
  AOI221_X1 U16838 ( .B1(P1_DATAO_REG_16__SCAN_IN), .B2(keyinput125), .C1(
        keyinput116), .C2(P2_REG0_REG_11__SCAN_IN), .A(n15307), .ZN(n15310) );
  OAI22_X1 U16839 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(keyinput98), .B1(
        keyinput93), .B2(P2_REG0_REG_18__SCAN_IN), .ZN(n15308) );
  AOI221_X1 U16840 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(keyinput98), .C1(
        P2_REG0_REG_18__SCAN_IN), .C2(keyinput93), .A(n15308), .ZN(n15309) );
  NAND4_X1 U16841 ( .A1(n15312), .A2(n15311), .A3(n15310), .A4(n15309), .ZN(
        n15345) );
  OAI22_X1 U16842 ( .A1(P3_REG0_REG_11__SCAN_IN), .A2(keyinput80), .B1(
        keyinput105), .B2(P1_REG0_REG_27__SCAN_IN), .ZN(n15313) );
  AOI221_X1 U16843 ( .B1(P3_REG0_REG_11__SCAN_IN), .B2(keyinput80), .C1(
        P1_REG0_REG_27__SCAN_IN), .C2(keyinput105), .A(n15313), .ZN(n15320) );
  OAI22_X1 U16844 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(keyinput79), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(keyinput96), .ZN(n15314) );
  AOI221_X1 U16845 ( .B1(P2_IR_REG_22__SCAN_IN), .B2(keyinput79), .C1(
        keyinput96), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n15314), .ZN(n15319) );
  OAI22_X1 U16846 ( .A1(SI_15_), .A2(keyinput102), .B1(keyinput97), .B2(
        P3_REG2_REG_30__SCAN_IN), .ZN(n15315) );
  AOI221_X1 U16847 ( .B1(SI_15_), .B2(keyinput102), .C1(
        P3_REG2_REG_30__SCAN_IN), .C2(keyinput97), .A(n15315), .ZN(n15318) );
  OAI22_X1 U16848 ( .A1(P3_D_REG_16__SCAN_IN), .A2(keyinput72), .B1(
        P3_REG1_REG_17__SCAN_IN), .B2(keyinput73), .ZN(n15316) );
  AOI221_X1 U16849 ( .B1(P3_D_REG_16__SCAN_IN), .B2(keyinput72), .C1(
        keyinput73), .C2(P3_REG1_REG_17__SCAN_IN), .A(n15316), .ZN(n15317) );
  NAND4_X1 U16850 ( .A1(n15320), .A2(n15319), .A3(n15318), .A4(n15317), .ZN(
        n15344) );
  OAI22_X1 U16851 ( .A1(n15323), .A2(keyinput82), .B1(n15322), .B2(keyinput104), .ZN(n15321) );
  AOI221_X1 U16852 ( .B1(n15323), .B2(keyinput82), .C1(keyinput104), .C2(
        n15322), .A(n15321), .ZN(n15333) );
  OAI22_X1 U16853 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(keyinput65), .B1(
        keyinput100), .B2(P3_ADDR_REG_8__SCAN_IN), .ZN(n15324) );
  AOI221_X1 U16854 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(keyinput65), .C1(
        P3_ADDR_REG_8__SCAN_IN), .C2(keyinput100), .A(n15324), .ZN(n15332) );
  XNOR2_X1 U16855 ( .A(n15325), .B(keyinput126), .ZN(n15328) );
  INV_X1 U16856 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n15326) );
  XNOR2_X1 U16857 ( .A(keyinput76), .B(n15326), .ZN(n15327) );
  NOR2_X1 U16858 ( .A1(n15328), .A2(n15327), .ZN(n15331) );
  OAI22_X1 U16859 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(keyinput78), .B1(
        keyinput64), .B2(P2_IR_REG_27__SCAN_IN), .ZN(n15329) );
  AOI221_X1 U16860 ( .B1(P2_IR_REG_13__SCAN_IN), .B2(keyinput78), .C1(
        P2_IR_REG_27__SCAN_IN), .C2(keyinput64), .A(n15329), .ZN(n15330) );
  NAND4_X1 U16861 ( .A1(n15333), .A2(n15332), .A3(n15331), .A4(n15330), .ZN(
        n15343) );
  OAI22_X1 U16862 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput85), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(keyinput68), .ZN(n15334) );
  AOI221_X1 U16863 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput85), .C1(
        keyinput68), .C2(P1_DATAO_REG_3__SCAN_IN), .A(n15334), .ZN(n15341) );
  OAI22_X1 U16864 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput88), .B1(
        keyinput119), .B2(P1_REG2_REG_10__SCAN_IN), .ZN(n15335) );
  AOI221_X1 U16865 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput88), .C1(
        P1_REG2_REG_10__SCAN_IN), .C2(keyinput119), .A(n15335), .ZN(n15340) );
  OAI22_X1 U16866 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(keyinput109), .B1(
        keyinput111), .B2(P1_REG3_REG_15__SCAN_IN), .ZN(n15336) );
  AOI221_X1 U16867 ( .B1(P2_DATAO_REG_19__SCAN_IN), .B2(keyinput109), .C1(
        P1_REG3_REG_15__SCAN_IN), .C2(keyinput111), .A(n15336), .ZN(n15339) );
  OAI22_X1 U16868 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(keyinput95), .B1(
        keyinput101), .B2(P2_ADDR_REG_1__SCAN_IN), .ZN(n15337) );
  AOI221_X1 U16869 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(keyinput95), .C1(
        P2_ADDR_REG_1__SCAN_IN), .C2(keyinput101), .A(n15337), .ZN(n15338) );
  NAND4_X1 U16870 ( .A1(n15341), .A2(n15340), .A3(n15339), .A4(n15338), .ZN(
        n15342) );
  NOR4_X1 U16871 ( .A1(n15345), .A2(n15344), .A3(n15343), .A4(n15342), .ZN(
        n15439) );
  AOI22_X1 U16872 ( .A1(P3_REG0_REG_11__SCAN_IN), .A2(keyinput16), .B1(
        P3_D_REG_29__SCAN_IN), .B2(keyinput58), .ZN(n15346) );
  OAI221_X1 U16873 ( .B1(P3_REG0_REG_11__SCAN_IN), .B2(keyinput16), .C1(
        P3_D_REG_29__SCAN_IN), .C2(keyinput58), .A(n15346), .ZN(n15353) );
  AOI22_X1 U16874 ( .A1(P2_D_REG_29__SCAN_IN), .A2(keyinput13), .B1(
        P3_REG1_REG_27__SCAN_IN), .B2(keyinput35), .ZN(n15347) );
  OAI221_X1 U16875 ( .B1(P2_D_REG_29__SCAN_IN), .B2(keyinput13), .C1(
        P3_REG1_REG_27__SCAN_IN), .C2(keyinput35), .A(n15347), .ZN(n15352) );
  AOI22_X1 U16876 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(keyinput47), .B1(
        P2_REG0_REG_11__SCAN_IN), .B2(keyinput52), .ZN(n15348) );
  OAI221_X1 U16877 ( .B1(P1_REG3_REG_15__SCAN_IN), .B2(keyinput47), .C1(
        P2_REG0_REG_11__SCAN_IN), .C2(keyinput52), .A(n15348), .ZN(n15351) );
  AOI22_X1 U16878 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(keyinput37), .B1(
        P2_REG0_REG_23__SCAN_IN), .B2(keyinput27), .ZN(n15349) );
  OAI221_X1 U16879 ( .B1(P2_ADDR_REG_1__SCAN_IN), .B2(keyinput37), .C1(
        P2_REG0_REG_23__SCAN_IN), .C2(keyinput27), .A(n15349), .ZN(n15350) );
  NOR4_X1 U16880 ( .A1(n15353), .A2(n15352), .A3(n15351), .A4(n15350), .ZN(
        n15381) );
  AOI22_X1 U16881 ( .A1(P2_REG0_REG_18__SCAN_IN), .A2(keyinput29), .B1(
        P2_IR_REG_13__SCAN_IN), .B2(keyinput14), .ZN(n15354) );
  OAI221_X1 U16882 ( .B1(P2_REG0_REG_18__SCAN_IN), .B2(keyinput29), .C1(
        P2_IR_REG_13__SCAN_IN), .C2(keyinput14), .A(n15354), .ZN(n15361) );
  AOI22_X1 U16883 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(keyinput32), .B1(
        P3_D_REG_12__SCAN_IN), .B2(keyinput10), .ZN(n15355) );
  OAI221_X1 U16884 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(keyinput32), .C1(
        P3_D_REG_12__SCAN_IN), .C2(keyinput10), .A(n15355), .ZN(n15360) );
  AOI22_X1 U16885 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(keyinput31), .B1(
        P3_REG2_REG_20__SCAN_IN), .B2(keyinput57), .ZN(n15356) );
  OAI221_X1 U16886 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(keyinput31), .C1(
        P3_REG2_REG_20__SCAN_IN), .C2(keyinput57), .A(n15356), .ZN(n15359) );
  AOI22_X1 U16887 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(keyinput12), .B1(
        P2_IR_REG_21__SCAN_IN), .B2(keyinput26), .ZN(n15357) );
  OAI221_X1 U16888 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(keyinput12), .C1(
        P2_IR_REG_21__SCAN_IN), .C2(keyinput26), .A(n15357), .ZN(n15358) );
  NOR4_X1 U16889 ( .A1(n15361), .A2(n15360), .A3(n15359), .A4(n15358), .ZN(
        n15380) );
  AOI22_X1 U16890 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(keyinput62), .B1(
        P2_REG0_REG_21__SCAN_IN), .B2(keyinput54), .ZN(n15362) );
  OAI221_X1 U16891 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(keyinput62), .C1(
        P2_REG0_REG_21__SCAN_IN), .C2(keyinput54), .A(n15362), .ZN(n15369) );
  AOI22_X1 U16892 ( .A1(P2_REG2_REG_29__SCAN_IN), .A2(keyinput53), .B1(
        P3_REG1_REG_17__SCAN_IN), .B2(keyinput9), .ZN(n15363) );
  OAI221_X1 U16893 ( .B1(P2_REG2_REG_29__SCAN_IN), .B2(keyinput53), .C1(
        P3_REG1_REG_17__SCAN_IN), .C2(keyinput9), .A(n15363), .ZN(n15368) );
  AOI22_X1 U16894 ( .A1(P2_REG2_REG_27__SCAN_IN), .A2(keyinput20), .B1(
        P2_D_REG_30__SCAN_IN), .B2(keyinput18), .ZN(n15364) );
  OAI221_X1 U16895 ( .B1(P2_REG2_REG_27__SCAN_IN), .B2(keyinput20), .C1(
        P2_D_REG_30__SCAN_IN), .C2(keyinput18), .A(n15364), .ZN(n15367) );
  AOI22_X1 U16896 ( .A1(P1_REG0_REG_27__SCAN_IN), .A2(keyinput41), .B1(
        P2_DATAO_REG_31__SCAN_IN), .B2(keyinput24), .ZN(n15365) );
  OAI221_X1 U16897 ( .B1(P1_REG0_REG_27__SCAN_IN), .B2(keyinput41), .C1(
        P2_DATAO_REG_31__SCAN_IN), .C2(keyinput24), .A(n15365), .ZN(n15366) );
  NOR4_X1 U16898 ( .A1(n15369), .A2(n15368), .A3(n15367), .A4(n15366), .ZN(
        n15379) );
  AOI22_X1 U16899 ( .A1(P3_DATAO_REG_3__SCAN_IN), .A2(keyinput46), .B1(
        P2_REG1_REG_11__SCAN_IN), .B2(keyinput1), .ZN(n15370) );
  OAI221_X1 U16900 ( .B1(P3_DATAO_REG_3__SCAN_IN), .B2(keyinput46), .C1(
        P2_REG1_REG_11__SCAN_IN), .C2(keyinput1), .A(n15370), .ZN(n15377) );
  AOI22_X1 U16901 ( .A1(P3_REG2_REG_29__SCAN_IN), .A2(keyinput22), .B1(
        P3_IR_REG_29__SCAN_IN), .B2(keyinput63), .ZN(n15371) );
  OAI221_X1 U16902 ( .B1(P3_REG2_REG_29__SCAN_IN), .B2(keyinput22), .C1(
        P3_IR_REG_29__SCAN_IN), .C2(keyinput63), .A(n15371), .ZN(n15376) );
  AOI22_X1 U16903 ( .A1(P2_D_REG_6__SCAN_IN), .A2(keyinput40), .B1(
        P3_IR_REG_30__SCAN_IN), .B2(keyinput50), .ZN(n15372) );
  OAI221_X1 U16904 ( .B1(P2_D_REG_6__SCAN_IN), .B2(keyinput40), .C1(
        P3_IR_REG_30__SCAN_IN), .C2(keyinput50), .A(n15372), .ZN(n15375) );
  AOI22_X1 U16905 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(keyinput0), .B1(
        P3_REG2_REG_8__SCAN_IN), .B2(keyinput5), .ZN(n15373) );
  OAI221_X1 U16906 ( .B1(P2_IR_REG_27__SCAN_IN), .B2(keyinput0), .C1(
        P3_REG2_REG_8__SCAN_IN), .C2(keyinput5), .A(n15373), .ZN(n15374) );
  NOR4_X1 U16907 ( .A1(n15377), .A2(n15376), .A3(n15375), .A4(n15374), .ZN(
        n15378) );
  NAND4_X1 U16908 ( .A1(n15381), .A2(n15380), .A3(n15379), .A4(n15378), .ZN(
        n15438) );
  AOI22_X1 U16909 ( .A1(n15384), .A2(keyinput3), .B1(keyinput7), .B2(n15383), 
        .ZN(n15382) );
  OAI221_X1 U16910 ( .B1(n15384), .B2(keyinput3), .C1(n15383), .C2(keyinput7), 
        .A(n15382), .ZN(n15396) );
  AOI22_X1 U16911 ( .A1(n15387), .A2(keyinput6), .B1(n15386), .B2(keyinput38), 
        .ZN(n15385) );
  OAI221_X1 U16912 ( .B1(n15387), .B2(keyinput6), .C1(n15386), .C2(keyinput38), 
        .A(n15385), .ZN(n15395) );
  AOI22_X1 U16913 ( .A1(n15390), .A2(keyinput43), .B1(n15389), .B2(keyinput30), 
        .ZN(n15388) );
  OAI221_X1 U16914 ( .B1(n15390), .B2(keyinput43), .C1(n15389), .C2(keyinput30), .A(n15388), .ZN(n15394) );
  XOR2_X1 U16915 ( .A(n7882), .B(keyinput11), .Z(n15392) );
  XNOR2_X1 U16916 ( .A(P3_IR_REG_5__SCAN_IN), .B(keyinput19), .ZN(n15391) );
  NAND2_X1 U16917 ( .A1(n15392), .A2(n15391), .ZN(n15393) );
  NOR4_X1 U16918 ( .A1(n15396), .A2(n15395), .A3(n15394), .A4(n15393), .ZN(
        n15436) );
  AOI22_X1 U16919 ( .A1(n15399), .A2(keyinput49), .B1(keyinput36), .B2(n15398), 
        .ZN(n15397) );
  OAI221_X1 U16920 ( .B1(n15399), .B2(keyinput49), .C1(n15398), .C2(keyinput36), .A(n15397), .ZN(n15408) );
  AOI22_X1 U16921 ( .A1(P1_REG2_REG_31__SCAN_IN), .A2(keyinput60), .B1(
        P1_REG1_REG_25__SCAN_IN), .B2(keyinput56), .ZN(n15400) );
  OAI221_X1 U16922 ( .B1(P1_REG2_REG_31__SCAN_IN), .B2(keyinput60), .C1(
        P1_REG1_REG_25__SCAN_IN), .C2(keyinput56), .A(n15400), .ZN(n15407) );
  XNOR2_X1 U16923 ( .A(n15401), .B(keyinput44), .ZN(n15406) );
  XNOR2_X1 U16924 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput4), .ZN(n15404) );
  XNOR2_X1 U16925 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(keyinput61), .ZN(n15403)
         );
  XNOR2_X1 U16926 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput21), .ZN(n15402)
         );
  NAND3_X1 U16927 ( .A1(n15404), .A2(n15403), .A3(n15402), .ZN(n15405) );
  NOR4_X1 U16928 ( .A1(n15408), .A2(n15407), .A3(n15406), .A4(n15405), .ZN(
        n15435) );
  AOI22_X1 U16929 ( .A1(n15410), .A2(keyinput2), .B1(keyinput25), .B2(n11034), 
        .ZN(n15409) );
  OAI221_X1 U16930 ( .B1(n15410), .B2(keyinput2), .C1(n11034), .C2(keyinput25), 
        .A(n15409), .ZN(n15419) );
  AOI22_X1 U16931 ( .A1(n15412), .A2(keyinput33), .B1(n7898), .B2(keyinput17), 
        .ZN(n15411) );
  OAI221_X1 U16932 ( .B1(n15412), .B2(keyinput33), .C1(n7898), .C2(keyinput17), 
        .A(n15411), .ZN(n15418) );
  AOI22_X1 U16933 ( .A1(n7901), .A2(keyinput34), .B1(keyinput23), .B2(n14179), 
        .ZN(n15413) );
  OAI221_X1 U16934 ( .B1(n7901), .B2(keyinput34), .C1(n14179), .C2(keyinput23), 
        .A(n15413), .ZN(n15417) );
  XNOR2_X1 U16935 ( .A(P3_REG1_REG_20__SCAN_IN), .B(keyinput42), .ZN(n15415)
         );
  XNOR2_X1 U16936 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput15), .ZN(n15414) );
  NAND2_X1 U16937 ( .A1(n15415), .A2(n15414), .ZN(n15416) );
  NOR4_X1 U16938 ( .A1(n15419), .A2(n15418), .A3(n15417), .A4(n15416), .ZN(
        n15434) );
  AOI22_X1 U16939 ( .A1(n10469), .A2(keyinput55), .B1(n7005), .B2(keyinput45), 
        .ZN(n15420) );
  OAI221_X1 U16940 ( .B1(n10469), .B2(keyinput55), .C1(n7005), .C2(keyinput45), 
        .A(n15420), .ZN(n15425) );
  XNOR2_X1 U16941 ( .A(n15421), .B(keyinput48), .ZN(n15424) );
  XNOR2_X1 U16942 ( .A(n15422), .B(keyinput39), .ZN(n15423) );
  OR3_X1 U16943 ( .A1(n15425), .A2(n15424), .A3(n15423), .ZN(n15432) );
  AOI22_X1 U16944 ( .A1(n11824), .A2(keyinput59), .B1(n15427), .B2(keyinput8), 
        .ZN(n15426) );
  OAI221_X1 U16945 ( .B1(n11824), .B2(keyinput59), .C1(n15427), .C2(keyinput8), 
        .A(n15426), .ZN(n15431) );
  AOI22_X1 U16946 ( .A1(n10158), .A2(keyinput51), .B1(n15429), .B2(keyinput28), 
        .ZN(n15428) );
  OAI221_X1 U16947 ( .B1(n10158), .B2(keyinput51), .C1(n15429), .C2(keyinput28), .A(n15428), .ZN(n15430) );
  NOR3_X1 U16948 ( .A1(n15432), .A2(n15431), .A3(n15430), .ZN(n15433) );
  NAND4_X1 U16949 ( .A1(n15436), .A2(n15435), .A3(n15434), .A4(n15433), .ZN(
        n15437) );
  AOI211_X1 U16950 ( .C1(n15440), .C2(n15439), .A(n15438), .B(n15437), .ZN(
        n15444) );
  NAND2_X1 U16951 ( .A1(n15441), .A2(P3_U3897), .ZN(n15442) );
  OAI21_X1 U16952 ( .B1(P3_U3897), .B2(P3_DATAO_REG_16__SCAN_IN), .A(n15442), 
        .ZN(n15443) );
  XNOR2_X1 U16953 ( .A(n15444), .B(n15443), .ZN(P3_U3507) );
  XOR2_X1 U16954 ( .A(n15446), .B(n15445), .Z(SUB_1596_U59) );
  XNOR2_X1 U16955 ( .A(n15447), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16956 ( .B1(n15449), .B2(n15448), .A(n15457), .ZN(SUB_1596_U53) );
  XOR2_X1 U16957 ( .A(n15450), .B(n15451), .Z(SUB_1596_U56) );
  OAI21_X1 U16958 ( .B1(n15454), .B2(n15453), .A(n15452), .ZN(n15455) );
  XNOR2_X1 U16959 ( .A(n15455), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  XOR2_X1 U16960 ( .A(n15457), .B(n15456), .Z(SUB_1596_U5) );
  INV_X2 U8369 ( .A(n11048), .ZN(n13604) );
  CLKBUF_X1 U7225 ( .A(n7788), .Z(n12895) );
endmodule

